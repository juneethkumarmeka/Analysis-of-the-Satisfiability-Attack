module basic_2000_20000_2500_40_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1605,In_1939);
and U1 (N_1,In_539,In_110);
and U2 (N_2,In_1023,In_1957);
nor U3 (N_3,In_327,In_1751);
nor U4 (N_4,In_1064,In_441);
or U5 (N_5,In_1103,In_1268);
or U6 (N_6,In_1140,In_1386);
nor U7 (N_7,In_885,In_450);
or U8 (N_8,In_1501,In_147);
nand U9 (N_9,In_820,In_608);
or U10 (N_10,In_171,In_646);
nor U11 (N_11,In_266,In_1571);
nor U12 (N_12,In_1733,In_949);
or U13 (N_13,In_1104,In_1361);
nor U14 (N_14,In_1496,In_1639);
or U15 (N_15,In_332,In_619);
nor U16 (N_16,In_439,In_948);
or U17 (N_17,In_193,In_644);
or U18 (N_18,In_1875,In_1589);
and U19 (N_19,In_1973,In_1168);
nor U20 (N_20,In_1811,In_476);
or U21 (N_21,In_1247,In_1293);
and U22 (N_22,In_1926,In_1357);
nor U23 (N_23,In_497,In_1533);
nand U24 (N_24,In_1857,In_1102);
or U25 (N_25,In_1473,In_808);
and U26 (N_26,In_279,In_756);
or U27 (N_27,In_943,In_500);
and U28 (N_28,In_106,In_385);
xnor U29 (N_29,In_702,In_1414);
nand U30 (N_30,In_1925,In_1828);
and U31 (N_31,In_225,In_1931);
nor U32 (N_32,In_417,In_514);
and U33 (N_33,In_1792,In_1946);
and U34 (N_34,In_483,In_596);
and U35 (N_35,In_871,In_1777);
or U36 (N_36,In_980,In_1389);
nand U37 (N_37,In_945,In_1175);
nor U38 (N_38,In_1216,In_1056);
nand U39 (N_39,In_452,In_773);
and U40 (N_40,In_79,In_1853);
or U41 (N_41,In_669,In_1510);
nor U42 (N_42,In_70,In_531);
and U43 (N_43,In_757,In_1679);
xnor U44 (N_44,In_1930,In_334);
nand U45 (N_45,In_1830,In_992);
or U46 (N_46,In_1573,In_1222);
nand U47 (N_47,In_648,In_309);
nand U48 (N_48,In_1479,In_1036);
nand U49 (N_49,In_1328,In_1863);
nand U50 (N_50,In_523,In_1867);
nand U51 (N_51,In_84,In_1918);
and U52 (N_52,In_817,In_1518);
nand U53 (N_53,In_1452,In_1907);
or U54 (N_54,In_739,In_663);
or U55 (N_55,In_302,In_745);
nor U56 (N_56,In_616,In_335);
nor U57 (N_57,In_315,In_1537);
and U58 (N_58,In_1786,In_402);
nand U59 (N_59,In_546,In_113);
nand U60 (N_60,In_971,In_314);
nor U61 (N_61,In_738,In_1065);
nor U62 (N_62,In_1517,In_433);
or U63 (N_63,In_1026,In_120);
xor U64 (N_64,In_359,In_10);
or U65 (N_65,In_1581,In_1621);
nor U66 (N_66,In_1719,In_1669);
nand U67 (N_67,In_625,In_1705);
nor U68 (N_68,In_706,In_510);
nor U69 (N_69,In_1708,In_382);
nor U70 (N_70,In_1068,In_287);
or U71 (N_71,In_1538,In_190);
nor U72 (N_72,In_1506,In_1425);
nor U73 (N_73,In_1028,In_1338);
or U74 (N_74,In_1944,In_1618);
xor U75 (N_75,In_714,In_479);
xor U76 (N_76,In_1149,In_1720);
nor U77 (N_77,In_1539,In_379);
and U78 (N_78,In_277,In_1241);
or U79 (N_79,In_983,In_1730);
nor U80 (N_80,In_785,In_1316);
nand U81 (N_81,In_698,In_1782);
nor U82 (N_82,In_1834,In_563);
or U83 (N_83,In_1963,In_1291);
or U84 (N_84,In_1899,In_1344);
and U85 (N_85,In_164,In_1864);
and U86 (N_86,In_291,In_1100);
nand U87 (N_87,In_1673,In_770);
nand U88 (N_88,In_1655,In_1549);
nor U89 (N_89,In_435,In_65);
and U90 (N_90,In_261,In_1649);
nand U91 (N_91,In_955,In_478);
nor U92 (N_92,In_244,In_428);
or U93 (N_93,In_1121,In_1002);
nor U94 (N_94,In_654,In_1732);
xnor U95 (N_95,In_1996,In_1094);
and U96 (N_96,In_605,In_1415);
nand U97 (N_97,In_683,In_1844);
or U98 (N_98,In_606,In_1681);
or U99 (N_99,In_519,In_867);
and U100 (N_100,In_1833,In_668);
and U101 (N_101,In_636,In_281);
nor U102 (N_102,In_73,In_722);
nor U103 (N_103,In_1579,In_1279);
nor U104 (N_104,In_656,In_1147);
and U105 (N_105,In_525,In_1006);
nor U106 (N_106,In_456,In_1876);
nand U107 (N_107,In_787,In_1166);
or U108 (N_108,In_1296,In_8);
nor U109 (N_109,In_1157,In_1628);
and U110 (N_110,In_484,In_251);
nand U111 (N_111,In_628,In_1155);
nor U112 (N_112,In_348,In_1896);
or U113 (N_113,In_1472,In_235);
nor U114 (N_114,In_1362,In_1829);
nor U115 (N_115,In_836,In_140);
nand U116 (N_116,In_13,In_1210);
nor U117 (N_117,In_1982,In_1892);
nand U118 (N_118,In_1053,In_445);
and U119 (N_119,In_587,In_117);
nand U120 (N_120,In_1906,In_1608);
and U121 (N_121,In_301,In_1770);
and U122 (N_122,In_1738,In_969);
and U123 (N_123,In_1968,In_1237);
nor U124 (N_124,In_1215,In_783);
nand U125 (N_125,In_517,In_394);
and U126 (N_126,In_200,In_1230);
nand U127 (N_127,In_1756,In_39);
nor U128 (N_128,In_1909,In_1250);
and U129 (N_129,In_1904,In_568);
and U130 (N_130,In_845,In_1635);
or U131 (N_131,In_1272,In_1124);
nor U132 (N_132,In_583,In_1118);
and U133 (N_133,In_1242,In_432);
nor U134 (N_134,In_552,In_1612);
or U135 (N_135,In_1217,In_135);
or U136 (N_136,In_1000,In_1278);
nor U137 (N_137,In_1716,In_1596);
nand U138 (N_138,In_473,In_96);
or U139 (N_139,In_1662,In_812);
and U140 (N_140,In_1249,In_1312);
or U141 (N_141,In_1275,In_901);
nor U142 (N_142,In_1895,In_1757);
and U143 (N_143,In_1183,In_60);
nor U144 (N_144,In_1526,In_710);
and U145 (N_145,In_1727,In_151);
nor U146 (N_146,In_1841,In_933);
nand U147 (N_147,In_1475,In_1873);
nand U148 (N_148,In_99,In_612);
and U149 (N_149,In_1880,In_1810);
or U150 (N_150,In_1602,In_138);
nor U151 (N_151,In_701,In_51);
nand U152 (N_152,In_797,In_127);
nor U153 (N_153,In_1041,In_838);
or U154 (N_154,In_1209,In_589);
or U155 (N_155,In_979,In_1342);
xnor U156 (N_156,In_290,In_639);
nand U157 (N_157,In_1910,In_1191);
or U158 (N_158,In_1771,In_1014);
or U159 (N_159,In_1504,In_310);
nor U160 (N_160,In_582,In_280);
nand U161 (N_161,In_565,In_278);
nor U162 (N_162,In_1185,In_32);
and U163 (N_163,In_900,In_796);
nor U164 (N_164,In_143,In_1154);
and U165 (N_165,In_803,In_726);
or U166 (N_166,In_1928,In_64);
nor U167 (N_167,In_1848,In_821);
or U168 (N_168,In_1158,In_1435);
nor U169 (N_169,In_1831,In_376);
or U170 (N_170,In_1260,In_1043);
nand U171 (N_171,In_666,In_371);
nor U172 (N_172,In_960,In_34);
or U173 (N_173,In_720,In_273);
and U174 (N_174,In_1208,In_951);
nand U175 (N_175,In_819,In_1683);
and U176 (N_176,In_1647,In_643);
or U177 (N_177,In_931,In_1707);
nor U178 (N_178,In_1850,In_1265);
or U179 (N_179,In_630,In_1039);
or U180 (N_180,In_216,In_1574);
nor U181 (N_181,In_1687,In_1257);
or U182 (N_182,In_1544,In_547);
and U183 (N_183,In_363,In_1862);
nor U184 (N_184,In_1491,In_313);
and U185 (N_185,In_1013,In_88);
xnor U186 (N_186,In_1570,In_1214);
or U187 (N_187,In_711,In_161);
nor U188 (N_188,In_1128,In_48);
or U189 (N_189,In_317,In_1801);
and U190 (N_190,In_1430,In_573);
nor U191 (N_191,In_369,In_1685);
and U192 (N_192,In_386,In_1497);
nand U193 (N_193,In_1854,In_1045);
or U194 (N_194,In_1358,In_1311);
or U195 (N_195,In_1148,In_1093);
and U196 (N_196,In_1565,In_904);
nand U197 (N_197,In_1370,In_130);
nand U198 (N_198,In_139,In_1402);
and U199 (N_199,In_1972,In_1646);
nor U200 (N_200,In_1456,In_1108);
or U201 (N_201,In_31,In_1568);
nor U202 (N_202,In_1440,In_1998);
or U203 (N_203,In_1162,In_769);
or U204 (N_204,In_1404,In_700);
nor U205 (N_205,In_468,In_883);
nand U206 (N_206,In_1694,In_367);
and U207 (N_207,In_912,In_851);
and U208 (N_208,In_860,In_1697);
nand U209 (N_209,In_337,In_790);
and U210 (N_210,In_1165,In_1345);
nor U211 (N_211,In_1986,In_118);
or U212 (N_212,In_984,In_938);
nand U213 (N_213,In_749,In_1084);
nor U214 (N_214,In_543,In_1980);
nand U215 (N_215,In_356,In_249);
and U216 (N_216,In_509,In_1059);
nand U217 (N_217,In_1933,In_870);
nor U218 (N_218,In_176,In_1392);
or U219 (N_219,In_36,In_237);
nor U220 (N_220,In_196,In_908);
nor U221 (N_221,In_1700,In_1110);
and U222 (N_222,In_1835,In_1809);
or U223 (N_223,In_585,In_358);
and U224 (N_224,In_453,In_929);
nor U225 (N_225,In_530,In_688);
and U226 (N_226,In_1119,In_1469);
nand U227 (N_227,In_1758,In_325);
nor U228 (N_228,In_53,In_2);
or U229 (N_229,In_1228,In_1839);
nor U230 (N_230,In_14,In_221);
xor U231 (N_231,In_276,In_1805);
or U232 (N_232,In_897,In_1021);
or U233 (N_233,In_22,In_555);
and U234 (N_234,In_160,In_1781);
and U235 (N_235,In_1253,In_189);
nor U236 (N_236,In_1412,In_300);
and U237 (N_237,In_418,In_805);
and U238 (N_238,In_857,In_1726);
and U239 (N_239,In_1812,In_1535);
nand U240 (N_240,In_810,In_416);
xnor U241 (N_241,In_1636,In_1849);
nor U242 (N_242,In_1901,In_1027);
and U243 (N_243,In_575,In_384);
nor U244 (N_244,In_1586,In_1569);
and U245 (N_245,In_288,In_131);
nor U246 (N_246,In_111,In_1945);
and U247 (N_247,In_1150,In_374);
nand U248 (N_248,In_1037,In_1657);
or U249 (N_249,In_1753,In_446);
and U250 (N_250,In_1717,In_1785);
nand U251 (N_251,In_482,In_26);
xnor U252 (N_252,In_1317,In_434);
nor U253 (N_253,In_1122,In_696);
nor U254 (N_254,In_466,In_1252);
nor U255 (N_255,In_581,In_227);
xor U256 (N_256,In_1672,In_352);
nand U257 (N_257,In_1625,In_1207);
or U258 (N_258,In_1146,In_1519);
nand U259 (N_259,In_1285,In_1181);
and U260 (N_260,In_1992,In_1595);
nor U261 (N_261,In_1527,In_1225);
and U262 (N_262,In_1624,In_556);
and U263 (N_263,In_856,In_778);
nand U264 (N_264,In_1198,In_1838);
and U265 (N_265,In_753,In_1299);
nor U266 (N_266,In_1741,In_1195);
nand U267 (N_267,In_1351,In_1858);
or U268 (N_268,In_1085,In_1558);
nand U269 (N_269,In_35,In_206);
and U270 (N_270,In_613,In_1413);
or U271 (N_271,In_30,In_823);
nor U272 (N_272,In_329,In_932);
and U273 (N_273,In_881,In_1817);
or U274 (N_274,In_1714,In_615);
nor U275 (N_275,In_1057,In_1650);
and U276 (N_276,In_766,In_19);
and U277 (N_277,In_684,In_1547);
nand U278 (N_278,In_1474,In_217);
or U279 (N_279,In_444,In_1471);
nand U280 (N_280,In_1325,In_1224);
and U281 (N_281,In_1827,In_77);
or U282 (N_282,In_631,In_561);
or U283 (N_283,In_112,In_360);
and U284 (N_284,In_108,In_1302);
and U285 (N_285,In_295,In_1659);
and U286 (N_286,In_991,In_534);
and U287 (N_287,In_1555,In_889);
and U288 (N_288,In_768,In_1139);
and U289 (N_289,In_1403,In_1005);
nand U290 (N_290,In_737,In_734);
nor U291 (N_291,In_214,In_494);
or U292 (N_292,In_1609,In_1219);
nor U293 (N_293,In_1420,In_1642);
or U294 (N_294,In_1449,In_1613);
nand U295 (N_295,In_406,In_437);
or U296 (N_296,In_564,In_63);
nor U297 (N_297,In_1480,In_1453);
and U298 (N_298,In_1067,In_451);
nor U299 (N_299,In_1962,In_809);
nand U300 (N_300,In_802,In_1987);
or U301 (N_301,In_1914,In_1004);
nor U302 (N_302,In_846,In_1594);
nand U303 (N_303,In_318,In_1540);
and U304 (N_304,In_179,In_1090);
nor U305 (N_305,In_887,In_877);
and U306 (N_306,In_392,In_843);
and U307 (N_307,In_818,In_306);
nand U308 (N_308,In_1887,In_957);
nor U309 (N_309,In_307,In_849);
nor U310 (N_310,In_1330,In_1695);
and U311 (N_311,In_560,In_1578);
nand U312 (N_312,In_532,In_833);
or U313 (N_313,In_1176,In_1256);
or U314 (N_314,In_1346,In_209);
nor U315 (N_315,In_1395,In_1038);
or U316 (N_316,In_799,In_1706);
or U317 (N_317,In_1360,In_292);
nor U318 (N_318,In_1567,In_776);
and U319 (N_319,In_1840,In_1324);
or U320 (N_320,In_1137,In_41);
nand U321 (N_321,In_675,In_1514);
or U322 (N_322,In_7,In_1120);
and U323 (N_323,In_144,In_1096);
nor U324 (N_324,In_940,In_975);
nor U325 (N_325,In_1401,In_536);
nand U326 (N_326,In_1033,In_89);
nand U327 (N_327,In_1597,In_1665);
or U328 (N_328,In_1188,In_1097);
or U329 (N_329,In_1759,In_464);
or U330 (N_330,In_1600,In_562);
nor U331 (N_331,In_1190,In_1676);
nor U332 (N_332,In_966,In_1744);
and U333 (N_333,In_1276,In_173);
nor U334 (N_334,In_1932,In_1333);
and U335 (N_335,In_829,In_25);
or U336 (N_336,In_569,In_1463);
and U337 (N_337,In_1807,In_754);
nor U338 (N_338,In_1248,In_1677);
or U339 (N_339,In_1836,In_1787);
nand U340 (N_340,In_1699,In_1457);
nor U341 (N_341,In_1913,In_430);
nand U342 (N_342,In_1941,In_331);
nor U343 (N_343,In_840,In_37);
nor U344 (N_344,In_1294,In_1587);
and U345 (N_345,In_1794,In_471);
nand U346 (N_346,In_149,In_798);
and U347 (N_347,In_76,In_1866);
or U348 (N_348,In_375,In_1654);
and U349 (N_349,In_1375,In_1383);
nand U350 (N_350,In_1803,In_664);
and U351 (N_351,In_1800,In_1916);
nand U352 (N_352,In_1079,In_865);
nand U353 (N_353,In_80,In_1105);
and U354 (N_354,In_93,In_1825);
or U355 (N_355,In_467,In_642);
and U356 (N_356,In_199,In_1696);
nor U357 (N_357,In_1832,In_124);
nand U358 (N_358,In_158,In_1750);
nand U359 (N_359,In_1437,In_772);
or U360 (N_360,In_1981,In_740);
nand U361 (N_361,In_690,In_353);
xnor U362 (N_362,In_1194,In_529);
and U363 (N_363,In_213,In_988);
nor U364 (N_364,In_1365,In_863);
nor U365 (N_365,In_1572,In_1689);
or U366 (N_366,In_1490,In_647);
nor U367 (N_367,In_487,In_342);
or U368 (N_368,In_712,In_340);
and U369 (N_369,In_1485,In_421);
or U370 (N_370,In_259,In_289);
xor U371 (N_371,In_588,In_492);
or U372 (N_372,In_1025,In_218);
nor U373 (N_373,In_1731,In_634);
nor U374 (N_374,In_602,In_105);
nand U375 (N_375,In_990,In_66);
nor U376 (N_376,In_254,In_873);
nand U377 (N_377,In_1815,In_377);
or U378 (N_378,In_1381,In_792);
nor U379 (N_379,In_1979,In_1837);
nand U380 (N_380,In_758,In_1813);
nor U381 (N_381,In_1116,In_659);
or U382 (N_382,In_47,In_748);
or U383 (N_383,In_1368,In_1988);
or U384 (N_384,In_174,In_761);
or U385 (N_385,In_886,In_1016);
and U386 (N_386,In_515,In_389);
nand U387 (N_387,In_178,In_1274);
nor U388 (N_388,In_1948,In_516);
and U389 (N_389,In_308,In_1894);
xnor U390 (N_390,In_658,In_1077);
or U391 (N_391,In_157,In_633);
and U392 (N_392,In_312,In_297);
and U393 (N_393,In_1623,In_1416);
and U394 (N_394,In_286,In_501);
or U395 (N_395,In_1055,In_1106);
nor U396 (N_396,In_258,In_1993);
and U397 (N_397,In_1554,In_526);
nand U398 (N_398,In_640,In_858);
nand U399 (N_399,In_191,In_366);
nor U400 (N_400,In_9,In_226);
and U401 (N_401,In_17,In_1954);
nand U402 (N_402,In_142,In_114);
and U403 (N_403,In_299,In_1458);
nand U404 (N_404,In_1664,In_1890);
nand U405 (N_405,In_1995,In_207);
nor U406 (N_406,In_0,In_239);
nor U407 (N_407,In_717,In_879);
and U408 (N_408,In_1729,In_595);
and U409 (N_409,In_1728,In_201);
or U410 (N_410,In_848,In_1542);
nor U411 (N_411,In_1536,In_346);
and U412 (N_412,In_1952,In_103);
and U413 (N_413,In_62,In_1966);
or U414 (N_414,In_972,In_1049);
nor U415 (N_415,In_1483,In_1897);
nand U416 (N_416,In_1465,In_985);
and U417 (N_417,In_921,In_1804);
nand U418 (N_418,In_275,In_1454);
or U419 (N_419,In_220,In_1520);
xor U420 (N_420,In_665,In_1069);
nor U421 (N_421,In_1598,In_1975);
or U422 (N_422,In_645,In_1397);
xor U423 (N_423,In_1123,In_601);
nor U424 (N_424,In_61,In_1099);
and U425 (N_425,In_511,In_162);
nand U426 (N_426,In_994,In_973);
or U427 (N_427,In_101,In_952);
and U428 (N_428,In_383,In_660);
and U429 (N_429,In_123,In_1132);
or U430 (N_430,In_1640,In_1630);
nand U431 (N_431,In_283,In_78);
nor U432 (N_432,In_1436,In_1385);
and U433 (N_433,In_1444,In_1213);
nand U434 (N_434,In_146,In_1281);
or U435 (N_435,In_771,In_1289);
nor U436 (N_436,In_1445,In_1938);
and U437 (N_437,In_1318,In_705);
and U438 (N_438,In_284,In_1762);
nor U439 (N_439,In_1113,In_593);
nor U440 (N_440,In_1062,In_687);
and U441 (N_441,In_1797,In_524);
nor U442 (N_442,In_567,In_1799);
or U443 (N_443,In_1088,In_210);
or U444 (N_444,In_1791,In_811);
nand U445 (N_445,In_600,In_1160);
nand U446 (N_446,In_1703,In_1347);
or U447 (N_447,In_1192,In_641);
or U448 (N_448,In_1870,In_1236);
or U449 (N_449,In_1240,In_1845);
or U450 (N_450,In_731,In_319);
or U451 (N_451,In_528,In_1965);
or U452 (N_452,In_1882,In_1656);
and U453 (N_453,In_1488,In_1502);
and U454 (N_454,In_255,In_584);
nor U455 (N_455,In_744,In_372);
nor U456 (N_456,In_1243,In_1802);
nand U457 (N_457,In_695,In_362);
and U458 (N_458,In_1081,In_43);
nand U459 (N_459,In_880,In_1865);
or U460 (N_460,In_1020,In_350);
or U461 (N_461,In_815,In_128);
nand U462 (N_462,In_1307,In_1722);
and U463 (N_463,In_566,In_759);
and U464 (N_464,In_1396,In_1852);
or U465 (N_465,In_126,In_397);
xnor U466 (N_466,In_305,In_1545);
xnor U467 (N_467,In_1507,In_219);
and U468 (N_468,In_942,In_752);
and U469 (N_469,In_400,In_1564);
or U470 (N_470,In_1843,In_175);
nand U471 (N_471,In_1961,In_1203);
nor U472 (N_472,In_1199,In_1552);
xor U473 (N_473,In_1877,In_1284);
and U474 (N_474,In_1955,In_545);
and U475 (N_475,In_1789,In_1776);
nor U476 (N_476,In_1616,In_1143);
nor U477 (N_477,In_1127,In_1739);
xnor U478 (N_478,In_1737,In_429);
and U479 (N_479,In_703,In_793);
nand U480 (N_480,In_842,In_964);
and U481 (N_481,In_559,In_246);
or U482 (N_482,In_784,In_1262);
or U483 (N_483,In_1723,In_1713);
nand U484 (N_484,In_155,In_55);
nor U485 (N_485,In_1796,In_493);
and U486 (N_486,In_1363,In_1818);
nand U487 (N_487,In_747,In_937);
and U488 (N_488,In_1201,In_1267);
nor U489 (N_489,In_1888,In_1089);
nand U490 (N_490,In_1304,In_344);
nand U491 (N_491,In_203,In_326);
or U492 (N_492,In_764,In_1310);
and U493 (N_493,In_1513,In_1331);
and U494 (N_494,In_1806,In_629);
or U495 (N_495,In_495,In_1292);
or U496 (N_496,In_592,In_920);
nor U497 (N_497,In_1784,In_580);
or U498 (N_498,In_490,In_1305);
nor U499 (N_499,In_1748,In_1891);
and U500 (N_500,N_343,N_86);
or U501 (N_501,N_462,In_1384);
nand U502 (N_502,N_48,In_298);
and U503 (N_503,N_270,In_141);
or U504 (N_504,N_103,N_429);
and U505 (N_505,In_1651,In_1410);
nor U506 (N_506,In_1956,N_336);
and U507 (N_507,N_301,In_963);
xnor U508 (N_508,N_488,In_970);
nand U509 (N_509,In_742,N_226);
nand U510 (N_510,In_859,In_522);
nor U511 (N_511,In_1072,In_939);
and U512 (N_512,N_328,N_326);
or U513 (N_513,N_183,In_250);
or U514 (N_514,N_265,N_214);
xnor U515 (N_515,N_108,N_53);
nand U516 (N_516,In_607,In_553);
and U517 (N_517,N_466,In_736);
or U518 (N_518,N_101,N_107);
or U519 (N_519,In_1532,In_1476);
nand U520 (N_520,In_1522,In_304);
nor U521 (N_521,In_1071,In_458);
nor U522 (N_522,N_251,In_1138);
nor U523 (N_523,In_1238,In_650);
and U524 (N_524,N_266,N_352);
nand U525 (N_525,In_610,In_763);
nor U526 (N_526,In_725,N_496);
nand U527 (N_527,In_412,In_1283);
nand U528 (N_528,In_294,N_246);
nor U529 (N_529,In_370,In_618);
nor U530 (N_530,N_6,N_221);
or U531 (N_531,In_599,In_1277);
nand U532 (N_532,N_458,N_62);
and U533 (N_533,N_479,In_1969);
or U534 (N_534,In_52,In_488);
and U535 (N_535,In_1101,N_416);
and U536 (N_536,In_322,N_369);
nand U537 (N_537,In_1076,N_232);
nand U538 (N_538,N_436,In_263);
or U539 (N_539,In_459,In_1058);
nor U540 (N_540,N_84,N_51);
nand U541 (N_541,In_1369,In_426);
nand U542 (N_542,In_894,In_169);
or U543 (N_543,N_110,In_1117);
or U544 (N_544,In_1417,In_1761);
and U545 (N_545,In_674,N_345);
nand U546 (N_546,N_457,N_386);
and U547 (N_547,N_424,N_80);
nand U548 (N_548,In_586,N_421);
and U549 (N_549,In_1083,In_271);
nand U550 (N_550,N_82,In_1012);
nand U551 (N_551,In_572,In_11);
nor U552 (N_552,N_374,N_341);
or U553 (N_553,In_777,In_1273);
and U554 (N_554,In_1261,In_676);
nand U555 (N_555,In_204,N_315);
and U556 (N_556,In_1196,N_319);
nand U557 (N_557,N_7,N_308);
or U558 (N_558,In_67,In_1953);
or U559 (N_559,In_709,In_579);
nor U560 (N_560,N_159,N_60);
xor U561 (N_561,N_117,In_496);
nor U562 (N_562,N_16,N_401);
nand U563 (N_563,In_474,In_655);
and U564 (N_564,In_197,N_150);
nor U565 (N_565,In_623,N_15);
nand U566 (N_566,In_1001,In_730);
and U567 (N_567,N_178,N_302);
nor U568 (N_568,In_1411,In_1629);
or U569 (N_569,N_392,N_339);
or U570 (N_570,In_1715,In_1583);
nand U571 (N_571,In_686,In_1354);
nand U572 (N_572,In_145,N_426);
or U573 (N_573,N_448,In_1743);
and U574 (N_574,In_202,N_229);
and U575 (N_575,In_187,In_751);
nand U576 (N_576,In_1653,In_902);
nand U577 (N_577,In_234,In_533);
nor U578 (N_578,In_1167,In_1808);
nand U579 (N_579,In_1061,N_346);
nor U580 (N_580,N_160,N_112);
nand U581 (N_581,In_472,N_172);
nand U582 (N_582,In_913,In_729);
or U583 (N_583,N_454,N_152);
or U584 (N_584,In_1874,In_1034);
xor U585 (N_585,In_211,In_170);
nand U586 (N_586,N_202,In_956);
or U587 (N_587,In_550,In_243);
nor U588 (N_588,In_841,In_916);
or U589 (N_589,N_409,N_131);
and U590 (N_590,In_1134,In_391);
and U591 (N_591,In_109,In_1044);
and U592 (N_592,In_1446,In_981);
or U593 (N_593,N_428,N_434);
nor U594 (N_594,In_1477,In_1929);
and U595 (N_595,In_715,In_850);
and U596 (N_596,In_953,In_557);
and U597 (N_597,In_898,In_1611);
nand U598 (N_598,In_1467,In_447);
and U599 (N_599,In_333,In_1408);
nand U600 (N_600,In_1173,In_1821);
nor U601 (N_601,In_148,In_1764);
xnor U602 (N_602,N_72,N_365);
nand U603 (N_603,In_381,N_411);
or U604 (N_604,In_1371,N_321);
nand U605 (N_605,In_1182,In_713);
nand U606 (N_606,In_1712,N_247);
or U607 (N_607,In_95,N_227);
or U608 (N_608,In_962,In_508);
and U609 (N_609,In_125,In_837);
or U610 (N_610,In_339,N_4);
and U611 (N_611,In_152,In_1881);
nor U612 (N_612,In_1164,In_576);
nor U613 (N_613,In_465,N_235);
xnor U614 (N_614,In_1266,In_965);
xor U615 (N_615,In_775,N_288);
or U616 (N_616,In_1314,In_436);
nand U617 (N_617,In_1340,In_708);
nor U618 (N_618,In_1428,N_260);
nor U619 (N_619,In_1631,N_79);
nand U620 (N_620,N_205,In_1136);
nand U621 (N_621,In_1846,In_475);
and U622 (N_622,In_1429,In_1159);
nand U623 (N_623,In_590,In_1200);
or U624 (N_624,N_238,In_97);
nor U625 (N_625,N_177,In_1098);
or U626 (N_626,N_14,In_1823);
nand U627 (N_627,N_440,In_470);
nand U628 (N_628,N_388,In_924);
or U629 (N_629,In_390,In_311);
and U630 (N_630,N_196,N_19);
nand U631 (N_631,N_295,In_1329);
nand U632 (N_632,In_195,In_950);
nor U633 (N_633,In_230,In_1643);
nand U634 (N_634,N_360,In_274);
or U635 (N_635,In_967,In_1271);
or U636 (N_636,In_409,N_189);
and U637 (N_637,In_1336,N_252);
nand U638 (N_638,In_351,N_334);
nand U639 (N_639,In_1905,In_69);
or U640 (N_640,N_442,In_499);
and U641 (N_641,N_480,In_1978);
or U642 (N_642,In_1842,In_765);
and U643 (N_643,In_1235,In_1795);
or U644 (N_644,In_1290,In_653);
nand U645 (N_645,In_864,N_453);
nor U646 (N_646,In_1516,In_535);
and U647 (N_647,N_314,In_934);
and U648 (N_648,N_477,In_1652);
or U649 (N_649,In_923,In_1494);
nand U650 (N_650,N_151,In_1352);
nor U651 (N_651,N_37,N_176);
or U652 (N_652,In_1111,In_541);
and U653 (N_653,In_1161,In_1588);
nor U654 (N_654,In_993,In_1889);
nand U655 (N_655,In_1179,In_1353);
and U656 (N_656,In_1859,In_1633);
or U657 (N_657,In_82,N_487);
nor U658 (N_658,In_544,In_780);
and U659 (N_659,In_296,In_743);
nor U660 (N_660,In_892,In_282);
or U661 (N_661,In_1721,In_1432);
nand U662 (N_662,In_574,In_469);
nor U663 (N_663,N_350,In_1964);
nand U664 (N_664,N_206,In_941);
or U665 (N_665,In_83,N_464);
nor U666 (N_666,In_1295,N_42);
or U667 (N_667,N_277,In_477);
nand U668 (N_668,N_398,N_459);
and U669 (N_669,In_919,N_433);
nor U670 (N_670,In_380,In_1202);
and U671 (N_671,In_673,N_299);
and U672 (N_672,N_95,N_78);
and U673 (N_673,In_1919,In_1793);
nor U674 (N_674,N_407,In_537);
or U675 (N_675,N_121,N_220);
nor U676 (N_676,In_172,In_989);
nor U677 (N_677,N_354,N_342);
nand U678 (N_678,In_1011,In_293);
or U679 (N_679,In_1169,In_1212);
or U680 (N_680,In_1671,In_1251);
or U681 (N_681,In_661,N_300);
nor U682 (N_682,N_310,In_1421);
or U683 (N_683,N_38,In_205);
nor U684 (N_684,In_995,In_1320);
nor U685 (N_685,In_1967,In_1523);
nand U686 (N_686,In_1779,N_372);
nand U687 (N_687,In_460,N_165);
and U688 (N_688,N_30,In_1227);
nand U689 (N_689,In_1433,In_1790);
or U690 (N_690,In_718,In_1382);
or U691 (N_691,In_1580,N_18);
nor U692 (N_692,In_723,In_50);
or U693 (N_693,In_789,N_190);
and U694 (N_694,In_1701,N_470);
nor U695 (N_695,N_186,In_1019);
nor U696 (N_696,In_861,In_1617);
nand U697 (N_697,In_1372,In_1172);
nor U698 (N_698,In_1950,N_200);
nand U699 (N_699,In_1563,N_175);
nand U700 (N_700,N_154,In_100);
nand U701 (N_701,N_25,N_188);
xnor U702 (N_702,In_1915,In_1530);
or U703 (N_703,In_443,N_122);
or U704 (N_704,In_1912,In_520);
and U705 (N_705,N_253,In_1614);
nand U706 (N_706,In_1824,In_56);
nor U707 (N_707,In_594,In_1591);
or U708 (N_708,In_1622,In_1441);
nand U709 (N_709,In_548,N_420);
and U710 (N_710,N_381,In_598);
nand U711 (N_711,N_306,In_888);
or U712 (N_712,In_521,N_47);
nor U713 (N_713,In_1958,In_91);
and U714 (N_714,N_325,In_27);
or U715 (N_715,In_1074,In_1170);
nand U716 (N_716,In_253,In_248);
nor U717 (N_717,In_760,In_834);
nand U718 (N_718,In_44,N_298);
nand U719 (N_719,In_1999,In_672);
nand U720 (N_720,In_1724,In_341);
nor U721 (N_721,N_102,In_399);
and U722 (N_722,In_1080,In_875);
and U723 (N_723,In_262,N_282);
nor U724 (N_724,In_398,In_448);
nand U725 (N_725,In_878,N_410);
or U726 (N_726,N_437,In_264);
nor U727 (N_727,N_320,In_1985);
or U728 (N_728,N_363,In_506);
nand U729 (N_729,In_944,In_741);
nor U730 (N_730,In_1989,N_274);
and U731 (N_731,In_1187,In_677);
or U732 (N_732,In_252,In_1658);
and U733 (N_733,N_224,In_361);
nor U734 (N_734,N_243,N_245);
nand U735 (N_735,In_1760,In_1460);
nor U736 (N_736,In_163,In_611);
or U737 (N_737,N_181,N_187);
nand U738 (N_738,In_1585,N_168);
or U739 (N_739,In_455,N_338);
xor U740 (N_740,In_1604,In_231);
and U741 (N_741,In_1478,In_1335);
nand U742 (N_742,In_791,In_1112);
or U743 (N_743,N_67,N_362);
and U744 (N_744,N_173,N_468);
and U745 (N_745,In_996,In_75);
nor U746 (N_746,N_316,In_1615);
and U747 (N_747,In_1493,N_432);
or U748 (N_748,In_917,In_1607);
or U749 (N_749,N_8,N_104);
and U750 (N_750,N_2,In_1704);
or U751 (N_751,In_68,In_542);
nand U752 (N_752,In_419,N_368);
nor U753 (N_753,In_1220,In_1814);
and U754 (N_754,In_844,In_1400);
or U755 (N_755,In_1619,N_275);
nor U756 (N_756,In_1977,In_192);
and U757 (N_757,N_132,In_1561);
nor U758 (N_758,In_1702,N_441);
nand U759 (N_759,In_1500,In_1718);
nand U760 (N_760,N_134,N_127);
or U761 (N_761,N_161,In_1348);
nor U762 (N_762,In_876,In_1135);
xnor U763 (N_763,N_413,In_46);
nor U764 (N_764,In_1040,N_261);
or U765 (N_765,N_353,In_1847);
or U766 (N_766,In_1606,N_141);
nand U767 (N_767,N_228,In_1052);
and U768 (N_768,In_1070,In_498);
and U769 (N_769,In_852,In_1184);
nor U770 (N_770,In_85,In_71);
nand U771 (N_771,In_1984,In_828);
and U772 (N_772,In_727,N_248);
or U773 (N_773,In_1590,In_680);
nand U774 (N_774,N_136,In_1898);
and U775 (N_775,In_724,In_1603);
and U776 (N_776,In_186,In_1855);
nor U777 (N_777,In_1145,In_662);
nor U778 (N_778,In_373,In_4);
nor U779 (N_779,In_365,N_471);
nor U780 (N_780,In_1936,In_270);
or U781 (N_781,N_391,In_959);
nor U782 (N_782,In_1951,In_1778);
xor U783 (N_783,In_1745,In_503);
nand U784 (N_784,In_396,N_494);
xor U785 (N_785,N_491,In_1487);
and U786 (N_786,In_922,N_303);
nor U787 (N_787,N_318,In_1178);
and U788 (N_788,In_1455,In_198);
or U789 (N_789,In_1900,N_234);
or U790 (N_790,In_1991,N_99);
nor U791 (N_791,In_1922,In_1007);
and U792 (N_792,In_1675,In_268);
nand U793 (N_793,N_399,N_167);
nand U794 (N_794,In_728,In_338);
nor U795 (N_795,N_361,N_311);
and U796 (N_796,In_685,N_375);
or U797 (N_797,In_1774,In_1258);
xnor U798 (N_798,N_125,In_16);
nor U799 (N_799,In_1018,N_166);
and U800 (N_800,In_1379,In_637);
nand U801 (N_801,N_387,In_1551);
and U802 (N_802,In_364,In_1923);
nor U803 (N_803,In_1893,In_485);
nor U804 (N_804,N_126,In_1484);
and U805 (N_805,In_1498,In_29);
nor U806 (N_806,In_442,In_440);
nor U807 (N_807,In_1393,In_49);
nor U808 (N_808,In_911,N_484);
nand U809 (N_809,N_417,In_1131);
nor U810 (N_810,N_359,In_905);
nor U811 (N_811,In_121,In_853);
nor U812 (N_812,In_368,N_156);
and U813 (N_813,In_926,In_1339);
nand U814 (N_814,In_1620,In_1543);
and U815 (N_815,In_256,N_71);
nor U816 (N_816,N_218,In_72);
nand U817 (N_817,N_397,N_367);
and U818 (N_818,In_1601,N_358);
and U819 (N_819,N_406,In_1763);
nand U820 (N_820,In_1470,In_1990);
and U821 (N_821,N_317,N_83);
nand U822 (N_822,In_1691,In_1003);
nand U823 (N_823,In_999,In_987);
nand U824 (N_824,N_493,N_465);
nor U825 (N_825,N_46,In_678);
nand U826 (N_826,In_914,N_225);
nand U827 (N_827,In_153,N_313);
nor U828 (N_828,In_1627,In_597);
and U829 (N_829,In_814,In_513);
or U830 (N_830,In_257,N_330);
xor U831 (N_831,In_427,In_1766);
or U832 (N_832,In_58,In_1947);
and U833 (N_833,In_1754,In_1078);
nor U834 (N_834,In_621,In_869);
and U835 (N_835,In_1711,In_133);
nor U836 (N_836,In_438,In_1450);
nor U837 (N_837,N_394,In_1288);
nand U838 (N_838,N_431,N_400);
nand U839 (N_839,N_492,N_443);
or U840 (N_840,In_632,N_280);
or U841 (N_841,N_193,In_1503);
or U842 (N_842,In_1576,N_66);
and U843 (N_843,N_182,In_1046);
and U844 (N_844,In_657,In_1355);
nand U845 (N_845,In_694,N_142);
and U846 (N_846,In_425,N_192);
nand U847 (N_847,In_1130,In_733);
and U848 (N_848,In_181,N_268);
and U849 (N_849,In_1462,In_1851);
and U850 (N_850,N_114,In_481);
and U851 (N_851,In_1211,N_174);
nand U852 (N_852,N_219,In_183);
nor U853 (N_853,N_147,In_413);
nand U854 (N_854,In_167,In_1282);
nand U855 (N_855,In_824,In_1775);
nand U856 (N_856,In_1949,N_40);
nand U857 (N_857,N_143,In_1350);
or U858 (N_858,In_936,N_39);
or U859 (N_859,N_271,In_571);
nand U860 (N_860,N_153,In_423);
or U861 (N_861,In_1742,In_116);
or U862 (N_862,N_26,N_257);
and U863 (N_863,In_132,N_366);
and U864 (N_864,In_1788,In_1690);
nand U865 (N_865,In_233,In_1528);
nor U866 (N_866,In_461,N_45);
xnor U867 (N_867,In_1593,In_1254);
or U868 (N_868,In_1599,In_652);
nand U869 (N_869,In_927,In_236);
nor U870 (N_870,In_1826,N_304);
nor U871 (N_871,In_918,In_830);
nand U872 (N_872,N_290,N_3);
nand U873 (N_873,In_1734,In_1332);
nor U874 (N_874,N_59,In_1693);
and U875 (N_875,In_907,N_461);
and U876 (N_876,In_1525,N_28);
or U877 (N_877,In_1868,In_681);
nand U878 (N_878,In_1270,N_119);
and U879 (N_879,In_156,In_1343);
or U880 (N_880,In_1218,In_38);
xor U881 (N_881,In_671,In_1780);
and U882 (N_882,In_15,N_382);
and U883 (N_883,N_408,N_452);
nor U884 (N_884,In_1407,N_404);
nor U885 (N_885,In_240,In_1073);
or U886 (N_886,N_481,In_679);
and U887 (N_887,In_330,N_129);
nand U888 (N_888,In_903,In_1908);
nand U889 (N_889,In_401,In_767);
or U890 (N_890,In_928,In_855);
and U891 (N_891,N_116,In_486);
or U892 (N_892,In_424,In_558);
nand U893 (N_893,N_216,In_825);
or U894 (N_894,In_1193,In_1534);
nor U895 (N_895,In_229,In_1047);
nand U896 (N_896,In_1466,In_1548);
and U897 (N_897,N_17,N_415);
nand U898 (N_898,In_1531,In_982);
or U899 (N_899,In_242,In_1661);
or U900 (N_900,In_1075,In_910);
or U901 (N_901,In_622,N_430);
or U902 (N_902,In_154,In_1577);
nand U903 (N_903,In_1431,In_925);
and U904 (N_904,N_144,In_935);
nor U905 (N_905,N_356,In_208);
nor U906 (N_906,In_1767,N_292);
and U907 (N_907,N_35,N_133);
nor U908 (N_908,In_1009,In_977);
nand U909 (N_909,In_1246,In_1521);
nor U910 (N_910,In_847,N_43);
nand U911 (N_911,N_305,N_324);
nor U912 (N_912,N_283,N_63);
nand U913 (N_913,N_263,In_480);
or U914 (N_914,In_891,In_1575);
and U915 (N_915,In_1180,In_102);
nor U916 (N_916,N_473,N_85);
nor U917 (N_917,N_128,In_168);
and U918 (N_918,In_269,In_1107);
or U919 (N_919,N_55,In_355);
or U920 (N_920,N_162,In_285);
nor U921 (N_921,N_393,N_256);
or U922 (N_922,In_28,N_482);
and U923 (N_923,In_1032,In_1935);
or U924 (N_924,N_357,In_1066);
nor U925 (N_925,N_169,In_1783);
nand U926 (N_926,In_538,N_377);
nor U927 (N_927,In_395,In_357);
or U928 (N_928,N_148,In_1768);
and U929 (N_929,In_549,In_33);
nand U930 (N_930,In_1287,In_1321);
or U931 (N_931,In_303,In_1970);
or U932 (N_932,In_1313,In_816);
nand U933 (N_933,In_241,N_478);
nand U934 (N_934,In_1245,In_746);
nor U935 (N_935,N_64,N_262);
xor U936 (N_936,In_1223,N_106);
and U937 (N_937,N_109,N_447);
or U938 (N_938,N_233,In_349);
nand U939 (N_939,N_74,In_930);
nand U940 (N_940,In_1641,N_20);
or U941 (N_941,In_343,In_1709);
nor U942 (N_942,In_378,N_287);
nand U943 (N_943,N_204,In_1816);
nand U944 (N_944,N_333,In_1566);
and U945 (N_945,In_603,N_49);
nand U946 (N_946,N_396,In_1374);
or U947 (N_947,N_191,In_512);
nand U948 (N_948,In_1688,N_5);
or U949 (N_949,In_1423,In_635);
or U950 (N_950,In_1438,N_207);
nor U951 (N_951,In_947,In_788);
nor U952 (N_952,In_1637,N_370);
nand U953 (N_953,In_1736,In_1663);
nand U954 (N_954,In_1886,In_54);
or U955 (N_955,In_1327,In_1869);
nor U956 (N_956,N_412,In_1388);
or U957 (N_957,In_1298,In_716);
nor U958 (N_958,In_895,In_1226);
and U959 (N_959,N_9,In_5);
nand U960 (N_960,N_258,N_323);
or U961 (N_961,N_348,N_364);
nand U962 (N_962,N_65,In_807);
or U963 (N_963,N_239,In_946);
nor U964 (N_964,In_1322,In_1424);
nand U965 (N_965,In_504,In_1592);
and U966 (N_966,N_383,In_420);
nor U967 (N_967,In_806,In_1419);
or U968 (N_968,In_180,In_1684);
nand U969 (N_969,In_906,In_958);
nor U970 (N_970,In_1660,In_801);
and U971 (N_971,In_1060,In_755);
nor U972 (N_972,In_90,In_527);
nor U973 (N_973,In_578,In_1746);
or U974 (N_974,N_486,In_1405);
nor U975 (N_975,In_1878,In_92);
or U976 (N_976,In_1481,In_1434);
or U977 (N_977,N_29,In_1442);
or U978 (N_978,In_177,In_1391);
and U979 (N_979,N_371,In_1752);
or U980 (N_980,In_1,In_1174);
nor U981 (N_981,In_1482,N_322);
or U982 (N_982,In_1648,In_1819);
or U983 (N_983,N_340,In_862);
nor U984 (N_984,In_502,N_445);
nor U985 (N_985,N_69,In_1234);
nand U986 (N_986,In_1367,In_260);
nand U987 (N_987,In_463,In_215);
or U988 (N_988,N_425,In_1974);
nor U989 (N_989,N_118,In_150);
or U990 (N_990,N_427,In_540);
nor U991 (N_991,In_1115,N_460);
nor U992 (N_992,N_10,N_68);
or U993 (N_993,N_98,N_24);
nand U994 (N_994,In_45,N_52);
or U995 (N_995,N_120,In_1092);
and U996 (N_996,In_1670,In_1959);
nor U997 (N_997,N_93,N_490);
nand U998 (N_998,In_1303,In_554);
or U999 (N_999,In_1259,In_704);
nor U1000 (N_1000,In_1422,N_556);
and U1001 (N_1001,In_854,N_648);
nor U1002 (N_1002,In_1366,N_910);
nor U1003 (N_1003,N_621,N_76);
nor U1004 (N_1004,N_449,N_741);
or U1005 (N_1005,N_327,N_549);
nand U1006 (N_1006,N_987,In_1378);
nand U1007 (N_1007,In_974,N_586);
or U1008 (N_1008,N_896,N_222);
or U1009 (N_1009,N_504,N_866);
or U1010 (N_1010,In_1668,N_605);
nand U1011 (N_1011,N_242,N_928);
nand U1012 (N_1012,In_732,N_730);
or U1013 (N_1013,N_644,N_567);
nor U1014 (N_1014,In_1204,N_631);
nand U1015 (N_1015,N_273,N_670);
nand U1016 (N_1016,N_972,N_842);
nand U1017 (N_1017,N_870,N_763);
or U1018 (N_1018,In_1468,In_222);
or U1019 (N_1019,N_933,In_1680);
or U1020 (N_1020,N_998,N_718);
nor U1021 (N_1021,N_210,N_557);
and U1022 (N_1022,In_212,In_1323);
nand U1023 (N_1023,N_777,N_598);
or U1024 (N_1024,N_516,N_990);
and U1025 (N_1025,In_1772,N_934);
nor U1026 (N_1026,N_757,N_709);
and U1027 (N_1027,In_1156,N_668);
nor U1028 (N_1028,N_779,In_624);
nor U1029 (N_1029,N_943,N_627);
nor U1030 (N_1030,N_951,N_850);
nor U1031 (N_1031,In_1029,N_163);
nor U1032 (N_1032,N_989,N_878);
nor U1033 (N_1033,In_505,N_640);
xor U1034 (N_1034,N_563,N_510);
nor U1035 (N_1035,In_976,In_1940);
or U1036 (N_1036,In_839,In_1042);
nand U1037 (N_1037,In_1151,N_883);
nand U1038 (N_1038,N_872,N_145);
nor U1039 (N_1039,In_1153,N_231);
nand U1040 (N_1040,N_882,N_916);
and U1041 (N_1041,In_1769,In_1610);
or U1042 (N_1042,N_291,In_518);
nor U1043 (N_1043,N_619,In_896);
xnor U1044 (N_1044,N_799,N_965);
or U1045 (N_1045,N_180,In_1309);
or U1046 (N_1046,N_754,N_686);
and U1047 (N_1047,In_570,N_679);
xnor U1048 (N_1048,N_941,N_767);
nand U1049 (N_1049,N_570,In_1921);
or U1050 (N_1050,N_863,N_701);
or U1051 (N_1051,In_1319,N_776);
nor U1052 (N_1052,In_21,N_552);
or U1053 (N_1053,N_956,N_911);
xor U1054 (N_1054,N_968,N_981);
xnor U1055 (N_1055,In_682,N_89);
nor U1056 (N_1056,N_900,N_969);
and U1057 (N_1057,N_505,N_795);
and U1058 (N_1058,N_782,In_786);
or U1059 (N_1059,In_59,In_1010);
nor U1060 (N_1060,In_1280,N_285);
nor U1061 (N_1061,In_909,N_250);
and U1062 (N_1062,In_1903,In_1860);
and U1063 (N_1063,In_1562,N_543);
xor U1064 (N_1064,In_779,In_1994);
or U1065 (N_1065,N_562,In_986);
or U1066 (N_1066,In_1409,N_75);
and U1067 (N_1067,N_771,N_975);
nand U1068 (N_1068,N_497,In_119);
or U1069 (N_1069,N_34,In_1233);
or U1070 (N_1070,N_804,N_859);
nand U1071 (N_1071,N_545,N_736);
nor U1072 (N_1072,In_1186,N_211);
nor U1073 (N_1073,N_255,N_501);
nor U1074 (N_1074,In_336,In_1205);
or U1075 (N_1075,N_915,In_1447);
nor U1076 (N_1076,N_73,N_518);
nor U1077 (N_1077,In_272,In_316);
and U1078 (N_1078,N_615,In_1439);
and U1079 (N_1079,In_1141,N_685);
and U1080 (N_1080,N_0,N_700);
and U1081 (N_1081,N_772,N_574);
or U1082 (N_1082,N_790,N_959);
nand U1083 (N_1083,N_841,N_532);
or U1084 (N_1084,N_832,In_826);
nand U1085 (N_1085,N_750,N_659);
nand U1086 (N_1086,N_715,In_1308);
or U1087 (N_1087,N_661,N_476);
nand U1088 (N_1088,In_1394,N_653);
or U1089 (N_1089,N_704,N_61);
nor U1090 (N_1090,N_852,N_851);
nor U1091 (N_1091,In_1109,In_794);
nor U1092 (N_1092,In_782,In_1725);
nand U1093 (N_1093,In_74,N_703);
nand U1094 (N_1094,In_1221,In_1553);
nand U1095 (N_1095,In_1133,In_1356);
or U1096 (N_1096,N_419,In_1418);
or U1097 (N_1097,In_1035,N_138);
and U1098 (N_1098,N_784,N_822);
or U1099 (N_1099,N_713,In_1443);
nor U1100 (N_1100,In_1263,N_942);
nor U1101 (N_1101,N_569,In_1239);
and U1102 (N_1102,N_985,N_137);
or U1103 (N_1103,In_223,In_874);
nor U1104 (N_1104,N_711,N_678);
nor U1105 (N_1105,In_866,In_1927);
nor U1106 (N_1106,N_32,N_828);
nor U1107 (N_1107,In_1334,In_414);
nand U1108 (N_1108,N_762,In_94);
and U1109 (N_1109,N_833,N_797);
nor U1110 (N_1110,N_373,N_976);
and U1111 (N_1111,N_611,N_11);
nand U1112 (N_1112,N_885,In_491);
or U1113 (N_1113,N_115,N_652);
nor U1114 (N_1114,N_249,N_513);
nand U1115 (N_1115,N_694,N_939);
nor U1116 (N_1116,N_402,N_418);
nor U1117 (N_1117,N_815,N_618);
nor U1118 (N_1118,N_230,N_684);
and U1119 (N_1119,N_12,N_826);
and U1120 (N_1120,In_1883,N_843);
nor U1121 (N_1121,N_884,N_595);
or U1122 (N_1122,N_512,N_922);
nor U1123 (N_1123,N_675,In_1902);
nand U1124 (N_1124,N_597,N_240);
nor U1125 (N_1125,N_696,N_893);
and U1126 (N_1126,N_873,In_1017);
or U1127 (N_1127,N_874,N_502);
nand U1128 (N_1128,N_606,N_810);
nand U1129 (N_1129,N_522,N_806);
or U1130 (N_1130,N_525,In_134);
nand U1131 (N_1131,N_816,N_607);
nor U1132 (N_1132,N_444,In_1710);
nor U1133 (N_1133,In_238,N_717);
or U1134 (N_1134,N_719,N_599);
or U1135 (N_1135,N_467,N_707);
or U1136 (N_1136,N_337,In_577);
nand U1137 (N_1137,In_649,N_612);
nand U1138 (N_1138,N_739,N_895);
or U1139 (N_1139,N_680,In_1971);
and U1140 (N_1140,N_332,N_748);
nor U1141 (N_1141,N_721,N_984);
nand U1142 (N_1142,N_879,N_825);
nand U1143 (N_1143,N_785,N_728);
nor U1144 (N_1144,N_921,N_897);
nor U1145 (N_1145,N_913,N_583);
nor U1146 (N_1146,N_854,N_979);
or U1147 (N_1147,N_906,N_405);
or U1148 (N_1148,N_940,N_269);
or U1149 (N_1149,In_1559,N_550);
nor U1150 (N_1150,N_966,N_539);
nand U1151 (N_1151,N_839,N_974);
nor U1152 (N_1152,N_179,In_638);
and U1153 (N_1153,In_1464,N_656);
nand U1154 (N_1154,N_50,N_536);
nand U1155 (N_1155,N_201,N_860);
and U1156 (N_1156,N_614,N_809);
nor U1157 (N_1157,N_349,N_953);
nand U1158 (N_1158,N_977,N_743);
nand U1159 (N_1159,N_929,In_697);
nand U1160 (N_1160,N_592,N_546);
nor U1161 (N_1161,N_281,N_293);
nor U1162 (N_1162,N_744,N_111);
nand U1163 (N_1163,N_455,In_404);
or U1164 (N_1164,N_573,N_946);
and U1165 (N_1165,N_687,N_857);
nand U1166 (N_1166,N_665,N_438);
nand U1167 (N_1167,In_813,N_868);
nand U1168 (N_1168,N_520,N_716);
nand U1169 (N_1169,In_1269,N_824);
and U1170 (N_1170,N_203,N_676);
nand U1171 (N_1171,In_1798,In_324);
nor U1172 (N_1172,N_297,N_31);
nor U1173 (N_1173,In_20,N_813);
and U1174 (N_1174,In_1022,N_993);
nand U1175 (N_1175,N_914,N_814);
nor U1176 (N_1176,In_689,In_1678);
and U1177 (N_1177,In_978,In_431);
nor U1178 (N_1178,N_259,In_1560);
nand U1179 (N_1179,In_1924,N_628);
nor U1180 (N_1180,N_651,N_164);
nand U1181 (N_1181,N_389,N_517);
and U1182 (N_1182,In_1426,N_647);
nand U1183 (N_1183,N_664,N_209);
nand U1184 (N_1184,N_902,N_912);
and U1185 (N_1185,N_856,N_451);
or U1186 (N_1186,In_12,N_760);
or U1187 (N_1187,In_998,N_919);
or U1188 (N_1188,In_182,N_714);
nand U1189 (N_1189,In_691,N_90);
nor U1190 (N_1190,N_602,N_329);
nor U1191 (N_1191,N_636,In_1879);
nand U1192 (N_1192,N_279,N_740);
nand U1193 (N_1193,N_309,In_795);
and U1194 (N_1194,N_964,In_721);
nand U1195 (N_1195,In_719,In_1373);
nor U1196 (N_1196,In_1541,N_56);
or U1197 (N_1197,N_955,N_158);
nor U1198 (N_1198,In_551,N_997);
nand U1199 (N_1199,In_1638,N_877);
nand U1200 (N_1200,N_803,N_507);
and U1201 (N_1201,In_247,N_683);
and U1202 (N_1202,N_962,N_495);
and U1203 (N_1203,In_626,N_585);
or U1204 (N_1204,N_590,N_376);
nand U1205 (N_1205,N_645,In_1524);
nand U1206 (N_1206,N_880,N_197);
xor U1207 (N_1207,In_489,In_1820);
nand U1208 (N_1208,In_40,N_712);
or U1209 (N_1209,N_735,N_1);
and U1210 (N_1210,In_87,N_589);
or U1211 (N_1211,In_1054,In_1152);
or U1212 (N_1212,N_542,N_891);
nand U1213 (N_1213,N_580,In_403);
nand U1214 (N_1214,In_6,N_475);
nor U1215 (N_1215,In_1632,N_140);
or U1216 (N_1216,N_637,N_198);
and U1217 (N_1217,In_1177,N_385);
nor U1218 (N_1218,N_610,N_335);
nor U1219 (N_1219,N_94,In_1315);
or U1220 (N_1220,N_861,N_331);
and U1221 (N_1221,N_184,N_380);
and U1222 (N_1222,N_667,N_961);
nor U1223 (N_1223,N_830,N_731);
or U1224 (N_1224,N_931,N_617);
nand U1225 (N_1225,N_92,In_1050);
nor U1226 (N_1226,N_690,N_938);
nor U1227 (N_1227,N_742,N_547);
or U1228 (N_1228,N_541,N_576);
nor U1229 (N_1229,N_267,N_519);
and U1230 (N_1230,In_1822,N_738);
and U1231 (N_1231,N_13,N_677);
or U1232 (N_1232,In_884,In_750);
nand U1233 (N_1233,N_91,N_87);
nor U1234 (N_1234,N_849,N_633);
or U1235 (N_1235,In_1550,N_195);
or U1236 (N_1236,N_559,In_868);
nor U1237 (N_1237,N_758,In_699);
nor U1238 (N_1238,In_1512,N_768);
nor U1239 (N_1239,N_769,In_1492);
and U1240 (N_1240,N_871,N_970);
nand U1241 (N_1241,N_554,N_945);
and U1242 (N_1242,N_21,N_96);
nor U1243 (N_1243,N_575,N_528);
or U1244 (N_1244,N_529,In_320);
nor U1245 (N_1245,N_561,In_1546);
nor U1246 (N_1246,N_604,N_498);
and U1247 (N_1247,N_783,N_641);
nor U1248 (N_1248,In_1765,In_347);
or U1249 (N_1249,N_821,In_1459);
nor U1250 (N_1250,N_773,N_982);
nand U1251 (N_1251,In_831,In_232);
nor U1252 (N_1252,N_862,N_881);
or U1253 (N_1253,N_834,In_1461);
nand U1254 (N_1254,In_1171,N_568);
nor U1255 (N_1255,N_820,N_995);
nand U1256 (N_1256,N_105,N_571);
or U1257 (N_1257,In_228,N_626);
nand U1258 (N_1258,N_514,In_1024);
nor U1259 (N_1259,N_710,N_609);
or U1260 (N_1260,N_515,In_328);
and U1261 (N_1261,N_720,N_135);
nor U1262 (N_1262,N_759,N_199);
or U1263 (N_1263,N_212,N_70);
or U1264 (N_1264,In_1376,N_837);
and U1265 (N_1265,In_591,N_698);
and U1266 (N_1266,N_623,N_608);
and U1267 (N_1267,N_761,N_54);
nor U1268 (N_1268,In_42,N_77);
nand U1269 (N_1269,In_462,In_954);
nor U1270 (N_1270,In_1051,In_822);
and U1271 (N_1271,In_3,In_1626);
nor U1272 (N_1272,N_469,In_1509);
nor U1273 (N_1273,In_1337,N_789);
and U1274 (N_1274,N_625,In_1231);
nor U1275 (N_1275,In_1942,N_523);
and U1276 (N_1276,N_765,N_812);
or U1277 (N_1277,N_403,In_136);
nor U1278 (N_1278,In_1529,In_774);
nor U1279 (N_1279,N_185,N_905);
and U1280 (N_1280,In_323,N_947);
nand U1281 (N_1281,In_184,N_732);
and U1282 (N_1282,N_936,N_733);
or U1283 (N_1283,N_509,N_456);
nor U1284 (N_1284,In_23,N_639);
or U1285 (N_1285,N_892,In_614);
or U1286 (N_1286,N_904,N_994);
nand U1287 (N_1287,In_1861,In_1095);
or U1288 (N_1288,N_876,N_781);
or U1289 (N_1289,N_845,N_967);
nand U1290 (N_1290,N_572,In_224);
and U1291 (N_1291,N_603,N_622);
nor U1292 (N_1292,N_666,N_472);
and U1293 (N_1293,N_553,N_727);
or U1294 (N_1294,In_1300,In_1682);
nor U1295 (N_1295,N_838,N_926);
or U1296 (N_1296,In_651,N_450);
or U1297 (N_1297,In_1634,In_1872);
nor U1298 (N_1298,N_948,N_887);
nand U1299 (N_1299,N_766,In_1448);
and U1300 (N_1300,In_1911,In_18);
nand U1301 (N_1301,N_286,N_819);
and U1302 (N_1302,N_963,N_708);
and U1303 (N_1303,N_801,N_706);
nand U1304 (N_1304,N_296,N_867);
and U1305 (N_1305,In_57,N_786);
and U1306 (N_1306,In_165,N_672);
and U1307 (N_1307,N_903,N_593);
and U1308 (N_1308,N_775,In_185);
nor U1309 (N_1309,In_1129,N_794);
nor U1310 (N_1310,N_33,In_762);
or U1311 (N_1311,N_474,N_691);
nor U1312 (N_1312,In_387,In_1871);
nor U1313 (N_1313,N_688,N_802);
and U1314 (N_1314,In_1326,N_980);
nand U1315 (N_1315,In_1505,In_1359);
nand U1316 (N_1316,N_836,N_534);
nor U1317 (N_1317,In_86,In_1556);
nand U1318 (N_1318,N_194,N_620);
and U1319 (N_1319,In_1644,N_531);
and U1320 (N_1320,In_1451,N_751);
nor U1321 (N_1321,N_705,N_601);
and U1322 (N_1322,In_1499,N_829);
nor U1323 (N_1323,In_1341,N_702);
and U1324 (N_1324,N_662,N_787);
nor U1325 (N_1325,N_932,In_1582);
xor U1326 (N_1326,In_393,In_98);
nor U1327 (N_1327,In_265,N_500);
nand U1328 (N_1328,N_954,N_747);
and U1329 (N_1329,N_579,N_582);
and U1330 (N_1330,In_1125,N_650);
or U1331 (N_1331,In_1740,N_535);
nor U1332 (N_1332,In_1114,N_960);
or U1333 (N_1333,In_422,N_734);
and U1334 (N_1334,In_129,N_937);
or U1335 (N_1335,N_681,N_483);
nor U1336 (N_1336,In_1495,N_752);
nand U1337 (N_1337,N_898,N_807);
nand U1338 (N_1338,N_499,In_620);
nor U1339 (N_1339,In_997,N_655);
and U1340 (N_1340,N_489,N_792);
and U1341 (N_1341,N_530,N_663);
nor U1342 (N_1342,In_800,N_635);
or U1343 (N_1343,N_999,In_345);
and U1344 (N_1344,In_1390,N_996);
nand U1345 (N_1345,N_347,N_643);
and U1346 (N_1346,N_634,N_791);
or U1347 (N_1347,N_920,N_577);
nand U1348 (N_1348,In_159,In_872);
nor U1349 (N_1349,In_1508,N_81);
or U1350 (N_1350,N_737,N_699);
nand U1351 (N_1351,N_521,In_1349);
nor U1352 (N_1352,In_24,N_764);
nor U1353 (N_1353,N_800,In_667);
or U1354 (N_1354,N_890,N_889);
and U1355 (N_1355,N_564,N_755);
nand U1356 (N_1356,N_565,In_1511);
or U1357 (N_1357,N_749,In_781);
nand U1358 (N_1358,In_1399,N_538);
and U1359 (N_1359,N_855,N_689);
nand U1360 (N_1360,In_1885,N_798);
and U1361 (N_1361,N_508,N_146);
nand U1362 (N_1362,N_682,N_591);
or U1363 (N_1363,In_454,N_692);
or U1364 (N_1364,N_524,N_924);
or U1365 (N_1365,In_104,In_1091);
or U1366 (N_1366,N_865,N_894);
or U1367 (N_1367,N_446,N_254);
or U1368 (N_1368,N_726,In_1406);
and U1369 (N_1369,N_864,In_1163);
nand U1370 (N_1370,N_908,N_823);
or U1371 (N_1371,In_1264,N_558);
nor U1372 (N_1372,In_388,N_671);
nand U1373 (N_1373,N_673,N_869);
and U1374 (N_1374,N_796,In_1486);
nand U1375 (N_1375,In_407,N_22);
nand U1376 (N_1376,N_658,N_983);
nand U1377 (N_1377,N_463,N_213);
nand U1378 (N_1378,N_986,N_566);
nand U1379 (N_1379,N_378,In_1735);
nor U1380 (N_1380,In_1255,N_171);
or U1381 (N_1381,N_284,N_139);
or U1382 (N_1382,In_1686,In_1086);
nor U1383 (N_1383,N_927,N_971);
nand U1384 (N_1384,In_122,N_853);
nor U1385 (N_1385,In_1030,N_439);
and U1386 (N_1386,N_817,N_379);
and U1387 (N_1387,N_41,In_411);
nand U1388 (N_1388,N_847,In_890);
nand U1389 (N_1389,N_925,N_533);
nor U1390 (N_1390,In_1917,N_944);
nand U1391 (N_1391,In_1286,N_780);
or U1392 (N_1392,N_560,N_511);
or U1393 (N_1393,N_695,N_630);
nand U1394 (N_1394,N_241,N_395);
nor U1395 (N_1395,In_1297,In_1997);
and U1396 (N_1396,N_638,N_674);
nor U1397 (N_1397,In_670,N_208);
or U1398 (N_1398,In_1048,N_276);
or U1399 (N_1399,N_808,N_899);
nand U1400 (N_1400,N_918,In_408);
and U1401 (N_1401,In_961,N_835);
or U1402 (N_1402,In_1377,N_646);
or U1403 (N_1403,N_312,N_594);
nand U1404 (N_1404,In_1008,In_1666);
and U1405 (N_1405,In_1427,N_544);
nand U1406 (N_1406,N_724,N_588);
and U1407 (N_1407,N_756,In_1126);
and U1408 (N_1408,In_617,N_827);
and U1409 (N_1409,In_354,In_1934);
nor U1410 (N_1410,In_321,N_722);
nand U1411 (N_1411,In_1557,N_632);
or U1412 (N_1412,In_899,N_616);
and U1413 (N_1413,N_949,N_978);
nor U1414 (N_1414,In_609,N_307);
and U1415 (N_1415,In_1306,In_267);
nor U1416 (N_1416,In_835,N_113);
nand U1417 (N_1417,N_289,In_1206);
nand U1418 (N_1418,N_992,In_166);
and U1419 (N_1419,N_58,N_875);
and U1420 (N_1420,N_149,N_988);
nor U1421 (N_1421,N_264,In_507);
nor U1422 (N_1422,N_624,In_1960);
and U1423 (N_1423,In_245,In_449);
and U1424 (N_1424,In_1244,N_840);
nand U1425 (N_1425,In_1015,In_1698);
nand U1426 (N_1426,In_1197,In_1031);
nand U1427 (N_1427,N_745,In_832);
or U1428 (N_1428,N_551,In_1144);
nor U1429 (N_1429,In_1976,N_657);
nor U1430 (N_1430,In_1749,N_527);
and U1431 (N_1431,In_1755,In_410);
nand U1432 (N_1432,N_27,N_649);
or U1433 (N_1433,In_604,N_223);
nand U1434 (N_1434,N_917,N_753);
nor U1435 (N_1435,N_344,In_81);
and U1436 (N_1436,In_627,N_581);
or U1437 (N_1437,N_600,N_435);
nor U1438 (N_1438,In_1082,N_729);
nand U1439 (N_1439,N_44,In_415);
and U1440 (N_1440,In_1229,N_858);
nor U1441 (N_1441,In_1301,In_1692);
nor U1442 (N_1442,In_115,N_503);
nor U1443 (N_1443,N_957,N_57);
or U1444 (N_1444,N_909,In_804);
or U1445 (N_1445,N_950,N_237);
or U1446 (N_1446,In_1667,In_1364);
nor U1447 (N_1447,N_930,In_968);
nand U1448 (N_1448,In_1920,N_526);
and U1449 (N_1449,In_1856,In_1983);
and U1450 (N_1450,N_414,N_725);
or U1451 (N_1451,N_793,N_778);
or U1452 (N_1452,N_907,N_555);
and U1453 (N_1453,In_1943,In_1142);
and U1454 (N_1454,N_36,N_540);
and U1455 (N_1455,N_958,N_818);
nor U1456 (N_1456,N_215,N_901);
and U1457 (N_1457,N_923,In_915);
nand U1458 (N_1458,In_1380,N_485);
xnor U1459 (N_1459,N_886,N_423);
and U1460 (N_1460,In_457,In_405);
nor U1461 (N_1461,N_537,N_697);
or U1462 (N_1462,N_506,In_1087);
nand U1463 (N_1463,N_846,N_991);
nand U1464 (N_1464,N_584,N_693);
nand U1465 (N_1465,In_1645,N_294);
nor U1466 (N_1466,N_596,In_693);
or U1467 (N_1467,In_137,In_882);
or U1468 (N_1468,N_629,N_774);
nand U1469 (N_1469,N_23,N_130);
or U1470 (N_1470,N_272,N_654);
nor U1471 (N_1471,In_692,N_770);
nor U1472 (N_1472,N_888,N_848);
and U1473 (N_1473,N_642,N_244);
and U1474 (N_1474,N_952,N_548);
and U1475 (N_1475,In_1884,N_123);
xnor U1476 (N_1476,N_587,In_707);
nand U1477 (N_1477,N_660,In_1937);
and U1478 (N_1478,N_973,N_355);
nand U1479 (N_1479,In_107,N_613);
or U1480 (N_1480,N_88,In_1674);
nor U1481 (N_1481,In_194,In_1584);
nor U1482 (N_1482,N_236,In_1398);
nand U1483 (N_1483,N_788,N_351);
nor U1484 (N_1484,In_1232,N_669);
or U1485 (N_1485,In_1773,N_422);
nand U1486 (N_1486,N_157,N_831);
and U1487 (N_1487,In_1387,In_1189);
and U1488 (N_1488,In_735,N_97);
nand U1489 (N_1489,N_844,N_746);
nor U1490 (N_1490,N_384,In_1515);
or U1491 (N_1491,N_100,In_893);
or U1492 (N_1492,In_188,In_1063);
and U1493 (N_1493,N_805,N_278);
nor U1494 (N_1494,N_124,In_827);
and U1495 (N_1495,N_935,N_578);
or U1496 (N_1496,In_1489,N_390);
nor U1497 (N_1497,N_155,N_217);
or U1498 (N_1498,N_811,N_723);
and U1499 (N_1499,N_170,In_1747);
and U1500 (N_1500,N_1175,N_1193);
or U1501 (N_1501,N_1412,N_1491);
and U1502 (N_1502,N_1257,N_1423);
nand U1503 (N_1503,N_1203,N_1405);
nor U1504 (N_1504,N_1072,N_1101);
and U1505 (N_1505,N_1165,N_1221);
nor U1506 (N_1506,N_1071,N_1037);
nor U1507 (N_1507,N_1170,N_1451);
and U1508 (N_1508,N_1186,N_1105);
xor U1509 (N_1509,N_1212,N_1296);
nor U1510 (N_1510,N_1332,N_1301);
nand U1511 (N_1511,N_1152,N_1145);
nor U1512 (N_1512,N_1126,N_1441);
and U1513 (N_1513,N_1015,N_1137);
nand U1514 (N_1514,N_1245,N_1365);
or U1515 (N_1515,N_1172,N_1415);
nor U1516 (N_1516,N_1255,N_1469);
nand U1517 (N_1517,N_1486,N_1272);
nand U1518 (N_1518,N_1450,N_1166);
and U1519 (N_1519,N_1322,N_1223);
or U1520 (N_1520,N_1076,N_1096);
and U1521 (N_1521,N_1446,N_1147);
nor U1522 (N_1522,N_1463,N_1346);
nand U1523 (N_1523,N_1281,N_1409);
nor U1524 (N_1524,N_1133,N_1499);
nor U1525 (N_1525,N_1222,N_1014);
or U1526 (N_1526,N_1494,N_1237);
nor U1527 (N_1527,N_1164,N_1006);
nand U1528 (N_1528,N_1309,N_1473);
nand U1529 (N_1529,N_1016,N_1075);
or U1530 (N_1530,N_1369,N_1227);
or U1531 (N_1531,N_1178,N_1366);
nand U1532 (N_1532,N_1102,N_1114);
or U1533 (N_1533,N_1058,N_1158);
xnor U1534 (N_1534,N_1111,N_1263);
nor U1535 (N_1535,N_1236,N_1268);
nor U1536 (N_1536,N_1427,N_1032);
nor U1537 (N_1537,N_1080,N_1083);
nor U1538 (N_1538,N_1442,N_1122);
nor U1539 (N_1539,N_1431,N_1249);
xnor U1540 (N_1540,N_1398,N_1484);
or U1541 (N_1541,N_1031,N_1429);
or U1542 (N_1542,N_1224,N_1368);
nand U1543 (N_1543,N_1213,N_1480);
or U1544 (N_1544,N_1008,N_1397);
nor U1545 (N_1545,N_1399,N_1407);
nand U1546 (N_1546,N_1261,N_1449);
or U1547 (N_1547,N_1355,N_1470);
nor U1548 (N_1548,N_1460,N_1005);
nand U1549 (N_1549,N_1112,N_1344);
nand U1550 (N_1550,N_1271,N_1216);
nor U1551 (N_1551,N_1052,N_1201);
and U1552 (N_1552,N_1074,N_1033);
nand U1553 (N_1553,N_1455,N_1478);
nor U1554 (N_1554,N_1230,N_1483);
xnor U1555 (N_1555,N_1337,N_1079);
nand U1556 (N_1556,N_1490,N_1396);
nor U1557 (N_1557,N_1256,N_1444);
and U1558 (N_1558,N_1046,N_1240);
nor U1559 (N_1559,N_1289,N_1089);
or U1560 (N_1560,N_1043,N_1310);
nand U1561 (N_1561,N_1180,N_1000);
nor U1562 (N_1562,N_1466,N_1218);
nor U1563 (N_1563,N_1479,N_1424);
and U1564 (N_1564,N_1234,N_1282);
or U1565 (N_1565,N_1044,N_1188);
nor U1566 (N_1566,N_1010,N_1199);
or U1567 (N_1567,N_1348,N_1125);
or U1568 (N_1568,N_1150,N_1389);
and U1569 (N_1569,N_1247,N_1454);
nand U1570 (N_1570,N_1078,N_1476);
or U1571 (N_1571,N_1085,N_1035);
nand U1572 (N_1572,N_1232,N_1123);
or U1573 (N_1573,N_1377,N_1362);
nand U1574 (N_1574,N_1229,N_1493);
and U1575 (N_1575,N_1340,N_1302);
nand U1576 (N_1576,N_1023,N_1211);
or U1577 (N_1577,N_1445,N_1059);
or U1578 (N_1578,N_1204,N_1163);
or U1579 (N_1579,N_1195,N_1329);
nand U1580 (N_1580,N_1034,N_1130);
xor U1581 (N_1581,N_1251,N_1090);
and U1582 (N_1582,N_1269,N_1179);
and U1583 (N_1583,N_1065,N_1330);
and U1584 (N_1584,N_1182,N_1320);
nor U1585 (N_1585,N_1465,N_1134);
nand U1586 (N_1586,N_1081,N_1060);
nor U1587 (N_1587,N_1017,N_1262);
or U1588 (N_1588,N_1316,N_1390);
or U1589 (N_1589,N_1073,N_1385);
or U1590 (N_1590,N_1131,N_1144);
nor U1591 (N_1591,N_1202,N_1207);
xor U1592 (N_1592,N_1275,N_1359);
or U1593 (N_1593,N_1136,N_1420);
or U1594 (N_1594,N_1413,N_1238);
nand U1595 (N_1595,N_1228,N_1287);
nand U1596 (N_1596,N_1432,N_1048);
and U1597 (N_1597,N_1135,N_1443);
nor U1598 (N_1598,N_1384,N_1307);
and U1599 (N_1599,N_1321,N_1098);
or U1600 (N_1600,N_1472,N_1153);
or U1601 (N_1601,N_1438,N_1051);
and U1602 (N_1602,N_1378,N_1371);
nand U1603 (N_1603,N_1258,N_1194);
or U1604 (N_1604,N_1278,N_1056);
nand U1605 (N_1605,N_1082,N_1250);
nor U1606 (N_1606,N_1294,N_1298);
and U1607 (N_1607,N_1403,N_1115);
nor U1608 (N_1608,N_1091,N_1244);
nor U1609 (N_1609,N_1118,N_1217);
nand U1610 (N_1610,N_1143,N_1146);
and U1611 (N_1611,N_1200,N_1311);
nor U1612 (N_1612,N_1488,N_1099);
nor U1613 (N_1613,N_1127,N_1109);
or U1614 (N_1614,N_1038,N_1300);
nor U1615 (N_1615,N_1279,N_1459);
or U1616 (N_1616,N_1364,N_1024);
or U1617 (N_1617,N_1174,N_1057);
nor U1618 (N_1618,N_1283,N_1208);
and U1619 (N_1619,N_1132,N_1107);
nor U1620 (N_1620,N_1293,N_1456);
and U1621 (N_1621,N_1266,N_1264);
nor U1622 (N_1622,N_1406,N_1485);
and U1623 (N_1623,N_1428,N_1265);
or U1624 (N_1624,N_1372,N_1084);
or U1625 (N_1625,N_1387,N_1284);
nor U1626 (N_1626,N_1086,N_1018);
or U1627 (N_1627,N_1149,N_1425);
and U1628 (N_1628,N_1104,N_1343);
and U1629 (N_1629,N_1197,N_1350);
and U1630 (N_1630,N_1013,N_1339);
and U1631 (N_1631,N_1410,N_1108);
or U1632 (N_1632,N_1276,N_1070);
or U1633 (N_1633,N_1360,N_1181);
or U1634 (N_1634,N_1467,N_1253);
or U1635 (N_1635,N_1007,N_1435);
nand U1636 (N_1636,N_1342,N_1226);
nor U1637 (N_1637,N_1171,N_1295);
and U1638 (N_1638,N_1291,N_1292);
nor U1639 (N_1639,N_1430,N_1440);
nor U1640 (N_1640,N_1411,N_1347);
or U1641 (N_1641,N_1448,N_1317);
nand U1642 (N_1642,N_1219,N_1209);
nand U1643 (N_1643,N_1148,N_1011);
nor U1644 (N_1644,N_1333,N_1142);
xor U1645 (N_1645,N_1367,N_1028);
and U1646 (N_1646,N_1280,N_1205);
nor U1647 (N_1647,N_1094,N_1335);
xnor U1648 (N_1648,N_1419,N_1388);
nand U1649 (N_1649,N_1254,N_1119);
nand U1650 (N_1650,N_1285,N_1157);
or U1651 (N_1651,N_1439,N_1246);
or U1652 (N_1652,N_1358,N_1187);
xor U1653 (N_1653,N_1045,N_1354);
nand U1654 (N_1654,N_1482,N_1452);
nor U1655 (N_1655,N_1386,N_1416);
nand U1656 (N_1656,N_1129,N_1069);
xnor U1657 (N_1657,N_1259,N_1139);
and U1658 (N_1658,N_1277,N_1004);
nand U1659 (N_1659,N_1319,N_1433);
and U1660 (N_1660,N_1021,N_1026);
and U1661 (N_1661,N_1110,N_1477);
or U1662 (N_1662,N_1453,N_1029);
and U1663 (N_1663,N_1379,N_1050);
nor U1664 (N_1664,N_1155,N_1394);
and U1665 (N_1665,N_1375,N_1159);
nor U1666 (N_1666,N_1248,N_1496);
and U1667 (N_1667,N_1039,N_1312);
or U1668 (N_1668,N_1288,N_1192);
and U1669 (N_1669,N_1242,N_1189);
nand U1670 (N_1670,N_1220,N_1267);
or U1671 (N_1671,N_1383,N_1345);
and U1672 (N_1672,N_1184,N_1055);
or U1673 (N_1673,N_1349,N_1068);
nor U1674 (N_1674,N_1331,N_1049);
and U1675 (N_1675,N_1214,N_1012);
nor U1676 (N_1676,N_1231,N_1323);
nand U1677 (N_1677,N_1233,N_1417);
and U1678 (N_1678,N_1437,N_1092);
nand U1679 (N_1679,N_1003,N_1001);
nor U1680 (N_1680,N_1243,N_1401);
nor U1681 (N_1681,N_1270,N_1156);
nor U1682 (N_1682,N_1421,N_1273);
or U1683 (N_1683,N_1036,N_1315);
or U1684 (N_1684,N_1325,N_1471);
nor U1685 (N_1685,N_1128,N_1169);
or U1686 (N_1686,N_1299,N_1206);
nand U1687 (N_1687,N_1097,N_1373);
or U1688 (N_1688,N_1318,N_1492);
or U1689 (N_1689,N_1376,N_1009);
nor U1690 (N_1690,N_1363,N_1324);
nand U1691 (N_1691,N_1225,N_1464);
nand U1692 (N_1692,N_1370,N_1481);
and U1693 (N_1693,N_1168,N_1434);
and U1694 (N_1694,N_1357,N_1025);
nand U1695 (N_1695,N_1489,N_1374);
or U1696 (N_1696,N_1177,N_1381);
xnor U1697 (N_1697,N_1391,N_1426);
nand U1698 (N_1698,N_1041,N_1239);
and U1699 (N_1699,N_1124,N_1140);
nor U1700 (N_1700,N_1351,N_1022);
nor U1701 (N_1701,N_1487,N_1196);
nor U1702 (N_1702,N_1027,N_1341);
or U1703 (N_1703,N_1141,N_1334);
nand U1704 (N_1704,N_1047,N_1042);
xor U1705 (N_1705,N_1167,N_1095);
or U1706 (N_1706,N_1392,N_1393);
nor U1707 (N_1707,N_1303,N_1297);
or U1708 (N_1708,N_1382,N_1100);
nor U1709 (N_1709,N_1457,N_1495);
nand U1710 (N_1710,N_1067,N_1162);
and U1711 (N_1711,N_1290,N_1103);
and U1712 (N_1712,N_1062,N_1215);
nand U1713 (N_1713,N_1461,N_1154);
or U1714 (N_1714,N_1402,N_1116);
nand U1715 (N_1715,N_1306,N_1210);
or U1716 (N_1716,N_1408,N_1198);
nand U1717 (N_1717,N_1308,N_1462);
nand U1718 (N_1718,N_1422,N_1474);
nor U1719 (N_1719,N_1336,N_1087);
and U1720 (N_1720,N_1404,N_1113);
and U1721 (N_1721,N_1352,N_1066);
and U1722 (N_1722,N_1185,N_1160);
xnor U1723 (N_1723,N_1053,N_1338);
nor U1724 (N_1724,N_1190,N_1002);
or U1725 (N_1725,N_1327,N_1328);
or U1726 (N_1726,N_1241,N_1138);
or U1727 (N_1727,N_1497,N_1176);
or U1728 (N_1728,N_1400,N_1120);
nor U1729 (N_1729,N_1093,N_1286);
and U1730 (N_1730,N_1106,N_1458);
and U1731 (N_1731,N_1414,N_1019);
nor U1732 (N_1732,N_1020,N_1380);
and U1733 (N_1733,N_1353,N_1252);
or U1734 (N_1734,N_1313,N_1030);
xnor U1735 (N_1735,N_1121,N_1117);
xnor U1736 (N_1736,N_1361,N_1305);
nand U1737 (N_1737,N_1475,N_1151);
nor U1738 (N_1738,N_1326,N_1395);
nor U1739 (N_1739,N_1088,N_1304);
nand U1740 (N_1740,N_1436,N_1356);
nand U1741 (N_1741,N_1274,N_1077);
nand U1742 (N_1742,N_1418,N_1040);
nand U1743 (N_1743,N_1314,N_1235);
nand U1744 (N_1744,N_1183,N_1447);
nand U1745 (N_1745,N_1161,N_1054);
and U1746 (N_1746,N_1061,N_1173);
nand U1747 (N_1747,N_1260,N_1191);
nand U1748 (N_1748,N_1498,N_1063);
or U1749 (N_1749,N_1468,N_1064);
nor U1750 (N_1750,N_1379,N_1432);
xor U1751 (N_1751,N_1277,N_1443);
nor U1752 (N_1752,N_1060,N_1434);
or U1753 (N_1753,N_1027,N_1050);
or U1754 (N_1754,N_1426,N_1323);
and U1755 (N_1755,N_1423,N_1444);
or U1756 (N_1756,N_1181,N_1315);
or U1757 (N_1757,N_1116,N_1383);
nor U1758 (N_1758,N_1060,N_1386);
and U1759 (N_1759,N_1253,N_1053);
or U1760 (N_1760,N_1141,N_1478);
and U1761 (N_1761,N_1445,N_1370);
nor U1762 (N_1762,N_1239,N_1336);
nor U1763 (N_1763,N_1426,N_1389);
and U1764 (N_1764,N_1423,N_1212);
and U1765 (N_1765,N_1345,N_1048);
xor U1766 (N_1766,N_1367,N_1385);
and U1767 (N_1767,N_1347,N_1441);
nand U1768 (N_1768,N_1332,N_1445);
nand U1769 (N_1769,N_1487,N_1091);
or U1770 (N_1770,N_1254,N_1339);
or U1771 (N_1771,N_1319,N_1249);
nand U1772 (N_1772,N_1004,N_1119);
nor U1773 (N_1773,N_1429,N_1079);
nor U1774 (N_1774,N_1073,N_1293);
and U1775 (N_1775,N_1287,N_1142);
nor U1776 (N_1776,N_1486,N_1126);
or U1777 (N_1777,N_1122,N_1497);
or U1778 (N_1778,N_1436,N_1452);
nand U1779 (N_1779,N_1250,N_1166);
or U1780 (N_1780,N_1248,N_1103);
or U1781 (N_1781,N_1301,N_1471);
and U1782 (N_1782,N_1198,N_1184);
or U1783 (N_1783,N_1317,N_1056);
and U1784 (N_1784,N_1215,N_1464);
nand U1785 (N_1785,N_1361,N_1078);
and U1786 (N_1786,N_1125,N_1358);
and U1787 (N_1787,N_1360,N_1261);
or U1788 (N_1788,N_1085,N_1375);
nand U1789 (N_1789,N_1268,N_1020);
and U1790 (N_1790,N_1482,N_1201);
or U1791 (N_1791,N_1121,N_1165);
and U1792 (N_1792,N_1245,N_1308);
and U1793 (N_1793,N_1493,N_1440);
or U1794 (N_1794,N_1163,N_1436);
nand U1795 (N_1795,N_1041,N_1477);
nor U1796 (N_1796,N_1496,N_1263);
nand U1797 (N_1797,N_1033,N_1279);
xor U1798 (N_1798,N_1347,N_1122);
nor U1799 (N_1799,N_1398,N_1337);
nand U1800 (N_1800,N_1236,N_1030);
nor U1801 (N_1801,N_1147,N_1287);
nor U1802 (N_1802,N_1294,N_1279);
nor U1803 (N_1803,N_1279,N_1479);
nand U1804 (N_1804,N_1487,N_1303);
xnor U1805 (N_1805,N_1096,N_1396);
and U1806 (N_1806,N_1322,N_1358);
and U1807 (N_1807,N_1471,N_1087);
nand U1808 (N_1808,N_1076,N_1084);
nor U1809 (N_1809,N_1451,N_1124);
nand U1810 (N_1810,N_1493,N_1372);
and U1811 (N_1811,N_1474,N_1042);
or U1812 (N_1812,N_1197,N_1310);
and U1813 (N_1813,N_1289,N_1423);
and U1814 (N_1814,N_1375,N_1219);
nand U1815 (N_1815,N_1067,N_1289);
or U1816 (N_1816,N_1167,N_1125);
and U1817 (N_1817,N_1039,N_1421);
nand U1818 (N_1818,N_1497,N_1147);
nand U1819 (N_1819,N_1340,N_1053);
nor U1820 (N_1820,N_1335,N_1433);
nand U1821 (N_1821,N_1367,N_1338);
nor U1822 (N_1822,N_1170,N_1096);
or U1823 (N_1823,N_1246,N_1347);
or U1824 (N_1824,N_1341,N_1333);
or U1825 (N_1825,N_1312,N_1455);
and U1826 (N_1826,N_1391,N_1320);
nand U1827 (N_1827,N_1494,N_1398);
or U1828 (N_1828,N_1471,N_1454);
and U1829 (N_1829,N_1270,N_1483);
or U1830 (N_1830,N_1054,N_1060);
or U1831 (N_1831,N_1173,N_1046);
or U1832 (N_1832,N_1047,N_1112);
and U1833 (N_1833,N_1110,N_1403);
or U1834 (N_1834,N_1037,N_1185);
or U1835 (N_1835,N_1456,N_1216);
or U1836 (N_1836,N_1319,N_1081);
nor U1837 (N_1837,N_1197,N_1348);
and U1838 (N_1838,N_1487,N_1312);
or U1839 (N_1839,N_1015,N_1178);
xnor U1840 (N_1840,N_1302,N_1179);
xnor U1841 (N_1841,N_1044,N_1438);
nand U1842 (N_1842,N_1070,N_1385);
and U1843 (N_1843,N_1416,N_1373);
nand U1844 (N_1844,N_1474,N_1138);
nor U1845 (N_1845,N_1376,N_1416);
and U1846 (N_1846,N_1379,N_1357);
nor U1847 (N_1847,N_1100,N_1418);
nor U1848 (N_1848,N_1414,N_1304);
and U1849 (N_1849,N_1327,N_1286);
or U1850 (N_1850,N_1413,N_1404);
or U1851 (N_1851,N_1423,N_1147);
or U1852 (N_1852,N_1486,N_1459);
nand U1853 (N_1853,N_1167,N_1271);
nand U1854 (N_1854,N_1041,N_1355);
nand U1855 (N_1855,N_1237,N_1183);
nor U1856 (N_1856,N_1390,N_1056);
nand U1857 (N_1857,N_1440,N_1163);
nor U1858 (N_1858,N_1467,N_1488);
nor U1859 (N_1859,N_1077,N_1300);
or U1860 (N_1860,N_1471,N_1328);
or U1861 (N_1861,N_1473,N_1250);
nor U1862 (N_1862,N_1071,N_1033);
nor U1863 (N_1863,N_1189,N_1377);
or U1864 (N_1864,N_1433,N_1279);
nor U1865 (N_1865,N_1290,N_1200);
or U1866 (N_1866,N_1209,N_1455);
nor U1867 (N_1867,N_1416,N_1036);
nor U1868 (N_1868,N_1391,N_1252);
nand U1869 (N_1869,N_1014,N_1484);
xor U1870 (N_1870,N_1379,N_1040);
or U1871 (N_1871,N_1331,N_1089);
nand U1872 (N_1872,N_1168,N_1185);
xor U1873 (N_1873,N_1214,N_1343);
nor U1874 (N_1874,N_1324,N_1010);
or U1875 (N_1875,N_1020,N_1490);
and U1876 (N_1876,N_1174,N_1029);
nor U1877 (N_1877,N_1058,N_1323);
and U1878 (N_1878,N_1166,N_1287);
xnor U1879 (N_1879,N_1232,N_1333);
nand U1880 (N_1880,N_1456,N_1404);
nor U1881 (N_1881,N_1422,N_1005);
nand U1882 (N_1882,N_1233,N_1342);
or U1883 (N_1883,N_1419,N_1067);
nor U1884 (N_1884,N_1498,N_1163);
and U1885 (N_1885,N_1120,N_1053);
and U1886 (N_1886,N_1350,N_1007);
and U1887 (N_1887,N_1209,N_1388);
nand U1888 (N_1888,N_1011,N_1425);
nor U1889 (N_1889,N_1379,N_1466);
or U1890 (N_1890,N_1053,N_1422);
nand U1891 (N_1891,N_1390,N_1130);
or U1892 (N_1892,N_1261,N_1077);
and U1893 (N_1893,N_1366,N_1463);
or U1894 (N_1894,N_1166,N_1475);
and U1895 (N_1895,N_1035,N_1390);
and U1896 (N_1896,N_1362,N_1371);
or U1897 (N_1897,N_1324,N_1445);
and U1898 (N_1898,N_1108,N_1325);
or U1899 (N_1899,N_1176,N_1325);
nor U1900 (N_1900,N_1195,N_1147);
xnor U1901 (N_1901,N_1395,N_1056);
or U1902 (N_1902,N_1329,N_1157);
or U1903 (N_1903,N_1070,N_1250);
nand U1904 (N_1904,N_1340,N_1018);
and U1905 (N_1905,N_1385,N_1010);
and U1906 (N_1906,N_1072,N_1111);
nor U1907 (N_1907,N_1370,N_1171);
and U1908 (N_1908,N_1458,N_1425);
or U1909 (N_1909,N_1423,N_1357);
nor U1910 (N_1910,N_1471,N_1374);
or U1911 (N_1911,N_1030,N_1156);
nor U1912 (N_1912,N_1482,N_1335);
or U1913 (N_1913,N_1176,N_1010);
or U1914 (N_1914,N_1268,N_1150);
nor U1915 (N_1915,N_1209,N_1119);
and U1916 (N_1916,N_1189,N_1096);
and U1917 (N_1917,N_1005,N_1068);
and U1918 (N_1918,N_1193,N_1124);
xnor U1919 (N_1919,N_1457,N_1406);
and U1920 (N_1920,N_1005,N_1267);
nor U1921 (N_1921,N_1477,N_1457);
nor U1922 (N_1922,N_1160,N_1227);
and U1923 (N_1923,N_1337,N_1271);
and U1924 (N_1924,N_1457,N_1088);
nor U1925 (N_1925,N_1005,N_1325);
nand U1926 (N_1926,N_1067,N_1370);
and U1927 (N_1927,N_1154,N_1287);
and U1928 (N_1928,N_1106,N_1099);
nand U1929 (N_1929,N_1054,N_1320);
and U1930 (N_1930,N_1144,N_1230);
and U1931 (N_1931,N_1174,N_1048);
nand U1932 (N_1932,N_1256,N_1328);
nor U1933 (N_1933,N_1289,N_1355);
nand U1934 (N_1934,N_1377,N_1099);
nand U1935 (N_1935,N_1472,N_1167);
nor U1936 (N_1936,N_1132,N_1084);
or U1937 (N_1937,N_1436,N_1384);
or U1938 (N_1938,N_1036,N_1035);
nor U1939 (N_1939,N_1233,N_1262);
and U1940 (N_1940,N_1284,N_1123);
and U1941 (N_1941,N_1345,N_1300);
and U1942 (N_1942,N_1154,N_1247);
or U1943 (N_1943,N_1495,N_1191);
and U1944 (N_1944,N_1375,N_1242);
or U1945 (N_1945,N_1171,N_1108);
and U1946 (N_1946,N_1031,N_1252);
nand U1947 (N_1947,N_1434,N_1055);
nor U1948 (N_1948,N_1307,N_1042);
and U1949 (N_1949,N_1135,N_1375);
xnor U1950 (N_1950,N_1135,N_1232);
nor U1951 (N_1951,N_1494,N_1137);
and U1952 (N_1952,N_1352,N_1415);
xnor U1953 (N_1953,N_1407,N_1366);
or U1954 (N_1954,N_1369,N_1464);
nand U1955 (N_1955,N_1150,N_1104);
nor U1956 (N_1956,N_1470,N_1035);
and U1957 (N_1957,N_1002,N_1112);
xor U1958 (N_1958,N_1373,N_1183);
nand U1959 (N_1959,N_1026,N_1029);
or U1960 (N_1960,N_1052,N_1179);
xnor U1961 (N_1961,N_1162,N_1404);
xor U1962 (N_1962,N_1072,N_1321);
and U1963 (N_1963,N_1259,N_1390);
or U1964 (N_1964,N_1425,N_1307);
nor U1965 (N_1965,N_1474,N_1128);
nor U1966 (N_1966,N_1090,N_1415);
nand U1967 (N_1967,N_1114,N_1182);
or U1968 (N_1968,N_1372,N_1183);
and U1969 (N_1969,N_1365,N_1454);
nand U1970 (N_1970,N_1447,N_1177);
nand U1971 (N_1971,N_1497,N_1120);
or U1972 (N_1972,N_1389,N_1096);
and U1973 (N_1973,N_1304,N_1144);
xnor U1974 (N_1974,N_1125,N_1441);
nor U1975 (N_1975,N_1456,N_1427);
nand U1976 (N_1976,N_1442,N_1496);
or U1977 (N_1977,N_1094,N_1460);
nand U1978 (N_1978,N_1194,N_1074);
nor U1979 (N_1979,N_1241,N_1219);
nor U1980 (N_1980,N_1198,N_1461);
or U1981 (N_1981,N_1405,N_1317);
nor U1982 (N_1982,N_1156,N_1371);
or U1983 (N_1983,N_1348,N_1070);
nor U1984 (N_1984,N_1286,N_1002);
nor U1985 (N_1985,N_1352,N_1329);
or U1986 (N_1986,N_1064,N_1100);
or U1987 (N_1987,N_1433,N_1014);
and U1988 (N_1988,N_1078,N_1417);
nand U1989 (N_1989,N_1396,N_1299);
or U1990 (N_1990,N_1369,N_1216);
nor U1991 (N_1991,N_1298,N_1304);
nand U1992 (N_1992,N_1289,N_1364);
nor U1993 (N_1993,N_1282,N_1068);
and U1994 (N_1994,N_1432,N_1166);
and U1995 (N_1995,N_1015,N_1089);
nand U1996 (N_1996,N_1011,N_1164);
nand U1997 (N_1997,N_1143,N_1287);
nor U1998 (N_1998,N_1475,N_1201);
and U1999 (N_1999,N_1291,N_1079);
or U2000 (N_2000,N_1724,N_1595);
nand U2001 (N_2001,N_1771,N_1743);
and U2002 (N_2002,N_1605,N_1768);
or U2003 (N_2003,N_1702,N_1844);
or U2004 (N_2004,N_1654,N_1892);
or U2005 (N_2005,N_1804,N_1908);
nand U2006 (N_2006,N_1759,N_1564);
nand U2007 (N_2007,N_1829,N_1730);
or U2008 (N_2008,N_1741,N_1664);
nor U2009 (N_2009,N_1584,N_1708);
nor U2010 (N_2010,N_1976,N_1931);
nand U2011 (N_2011,N_1715,N_1933);
or U2012 (N_2012,N_1902,N_1573);
and U2013 (N_2013,N_1623,N_1524);
or U2014 (N_2014,N_1675,N_1577);
nor U2015 (N_2015,N_1587,N_1515);
nand U2016 (N_2016,N_1954,N_1533);
nand U2017 (N_2017,N_1549,N_1838);
or U2018 (N_2018,N_1793,N_1789);
nor U2019 (N_2019,N_1568,N_1596);
or U2020 (N_2020,N_1689,N_1751);
nor U2021 (N_2021,N_1792,N_1758);
nor U2022 (N_2022,N_1853,N_1643);
nor U2023 (N_2023,N_1574,N_1858);
nor U2024 (N_2024,N_1923,N_1508);
nor U2025 (N_2025,N_1728,N_1590);
or U2026 (N_2026,N_1502,N_1677);
or U2027 (N_2027,N_1993,N_1887);
or U2028 (N_2028,N_1613,N_1937);
nor U2029 (N_2029,N_1553,N_1952);
or U2030 (N_2030,N_1698,N_1714);
or U2031 (N_2031,N_1671,N_1622);
nor U2032 (N_2032,N_1755,N_1628);
nand U2033 (N_2033,N_1554,N_1523);
and U2034 (N_2034,N_1692,N_1944);
nand U2035 (N_2035,N_1682,N_1784);
nor U2036 (N_2036,N_1917,N_1879);
or U2037 (N_2037,N_1561,N_1669);
nand U2038 (N_2038,N_1722,N_1555);
nand U2039 (N_2039,N_1816,N_1990);
and U2040 (N_2040,N_1836,N_1802);
nand U2041 (N_2041,N_1935,N_1780);
nand U2042 (N_2042,N_1672,N_1712);
nor U2043 (N_2043,N_1635,N_1795);
or U2044 (N_2044,N_1960,N_1987);
nand U2045 (N_2045,N_1552,N_1537);
nor U2046 (N_2046,N_1786,N_1968);
and U2047 (N_2047,N_1504,N_1765);
and U2048 (N_2048,N_1681,N_1992);
nand U2049 (N_2049,N_1746,N_1773);
nor U2050 (N_2050,N_1875,N_1513);
or U2051 (N_2051,N_1897,N_1685);
or U2052 (N_2052,N_1785,N_1868);
or U2053 (N_2053,N_1687,N_1979);
or U2054 (N_2054,N_1831,N_1691);
nand U2055 (N_2055,N_1601,N_1866);
or U2056 (N_2056,N_1617,N_1857);
nor U2057 (N_2057,N_1840,N_1511);
nor U2058 (N_2058,N_1950,N_1860);
and U2059 (N_2059,N_1631,N_1646);
nor U2060 (N_2060,N_1713,N_1888);
and U2061 (N_2061,N_1794,N_1761);
nor U2062 (N_2062,N_1823,N_1727);
or U2063 (N_2063,N_1907,N_1556);
nor U2064 (N_2064,N_1753,N_1589);
nand U2065 (N_2065,N_1739,N_1750);
nor U2066 (N_2066,N_1567,N_1830);
nand U2067 (N_2067,N_1695,N_1690);
and U2068 (N_2068,N_1781,N_1859);
nor U2069 (N_2069,N_1930,N_1873);
and U2070 (N_2070,N_1565,N_1641);
or U2071 (N_2071,N_1890,N_1837);
and U2072 (N_2072,N_1655,N_1649);
or U2073 (N_2073,N_1704,N_1970);
and U2074 (N_2074,N_1865,N_1807);
or U2075 (N_2075,N_1606,N_1855);
nor U2076 (N_2076,N_1676,N_1774);
or U2077 (N_2077,N_1578,N_1763);
xnor U2078 (N_2078,N_1749,N_1877);
and U2079 (N_2079,N_1540,N_1534);
nor U2080 (N_2080,N_1788,N_1705);
or U2081 (N_2081,N_1921,N_1744);
or U2082 (N_2082,N_1583,N_1520);
and U2083 (N_2083,N_1949,N_1645);
xnor U2084 (N_2084,N_1965,N_1947);
and U2085 (N_2085,N_1633,N_1674);
nor U2086 (N_2086,N_1560,N_1500);
nand U2087 (N_2087,N_1599,N_1967);
nor U2088 (N_2088,N_1934,N_1754);
nand U2089 (N_2089,N_1847,N_1787);
nor U2090 (N_2090,N_1863,N_1939);
and U2091 (N_2091,N_1607,N_1512);
nand U2092 (N_2092,N_1963,N_1598);
nand U2093 (N_2093,N_1615,N_1521);
and U2094 (N_2094,N_1852,N_1946);
and U2095 (N_2095,N_1639,N_1706);
or U2096 (N_2096,N_1660,N_1725);
nor U2097 (N_2097,N_1919,N_1550);
nand U2098 (N_2098,N_1699,N_1679);
nor U2099 (N_2099,N_1911,N_1668);
or U2100 (N_2100,N_1642,N_1629);
or U2101 (N_2101,N_1618,N_1594);
or U2102 (N_2102,N_1572,N_1582);
and U2103 (N_2103,N_1527,N_1720);
nor U2104 (N_2104,N_1964,N_1586);
nor U2105 (N_2105,N_1718,N_1870);
nor U2106 (N_2106,N_1820,N_1841);
or U2107 (N_2107,N_1736,N_1834);
nand U2108 (N_2108,N_1542,N_1833);
or U2109 (N_2109,N_1878,N_1637);
nor U2110 (N_2110,N_1891,N_1723);
or U2111 (N_2111,N_1593,N_1581);
or U2112 (N_2112,N_1977,N_1528);
nor U2113 (N_2113,N_1899,N_1673);
and U2114 (N_2114,N_1592,N_1996);
or U2115 (N_2115,N_1544,N_1825);
nor U2116 (N_2116,N_1636,N_1822);
or U2117 (N_2117,N_1734,N_1536);
or U2118 (N_2118,N_1986,N_1576);
nand U2119 (N_2119,N_1651,N_1988);
nor U2120 (N_2120,N_1882,N_1700);
or U2121 (N_2121,N_1611,N_1980);
or U2122 (N_2122,N_1678,N_1849);
and U2123 (N_2123,N_1546,N_1747);
or U2124 (N_2124,N_1604,N_1703);
or U2125 (N_2125,N_1721,N_1925);
nand U2126 (N_2126,N_1969,N_1850);
nor U2127 (N_2127,N_1505,N_1588);
and U2128 (N_2128,N_1777,N_1731);
nor U2129 (N_2129,N_1740,N_1842);
nand U2130 (N_2130,N_1864,N_1693);
nor U2131 (N_2131,N_1506,N_1800);
or U2132 (N_2132,N_1883,N_1994);
xor U2133 (N_2133,N_1711,N_1627);
and U2134 (N_2134,N_1648,N_1958);
xnor U2135 (N_2135,N_1716,N_1936);
or U2136 (N_2136,N_1757,N_1610);
or U2137 (N_2137,N_1570,N_1770);
nor U2138 (N_2138,N_1748,N_1752);
nor U2139 (N_2139,N_1647,N_1558);
nor U2140 (N_2140,N_1983,N_1991);
and U2141 (N_2141,N_1885,N_1846);
or U2142 (N_2142,N_1719,N_1966);
or U2143 (N_2143,N_1955,N_1760);
or U2144 (N_2144,N_1798,N_1975);
or U2145 (N_2145,N_1898,N_1626);
or U2146 (N_2146,N_1501,N_1791);
nor U2147 (N_2147,N_1562,N_1707);
or U2148 (N_2148,N_1951,N_1656);
or U2149 (N_2149,N_1614,N_1808);
nand U2150 (N_2150,N_1625,N_1783);
nor U2151 (N_2151,N_1519,N_1906);
and U2152 (N_2152,N_1900,N_1959);
and U2153 (N_2153,N_1922,N_1518);
and U2154 (N_2154,N_1717,N_1904);
nor U2155 (N_2155,N_1545,N_1650);
or U2156 (N_2156,N_1597,N_1538);
nand U2157 (N_2157,N_1600,N_1799);
and U2158 (N_2158,N_1630,N_1978);
nand U2159 (N_2159,N_1805,N_1889);
nand U2160 (N_2160,N_1843,N_1810);
nand U2161 (N_2161,N_1827,N_1551);
xnor U2162 (N_2162,N_1943,N_1697);
nor U2163 (N_2163,N_1809,N_1973);
or U2164 (N_2164,N_1579,N_1894);
or U2165 (N_2165,N_1670,N_1517);
or U2166 (N_2166,N_1881,N_1522);
nand U2167 (N_2167,N_1856,N_1817);
or U2168 (N_2168,N_1998,N_1516);
and U2169 (N_2169,N_1608,N_1621);
or U2170 (N_2170,N_1624,N_1580);
nor U2171 (N_2171,N_1742,N_1880);
or U2172 (N_2172,N_1530,N_1938);
nor U2173 (N_2173,N_1945,N_1826);
nand U2174 (N_2174,N_1652,N_1814);
or U2175 (N_2175,N_1812,N_1926);
nand U2176 (N_2176,N_1709,N_1845);
or U2177 (N_2177,N_1912,N_1972);
or U2178 (N_2178,N_1920,N_1667);
nor U2179 (N_2179,N_1862,N_1575);
nand U2180 (N_2180,N_1957,N_1839);
or U2181 (N_2181,N_1948,N_1738);
nand U2182 (N_2182,N_1874,N_1941);
nor U2183 (N_2183,N_1927,N_1803);
nand U2184 (N_2184,N_1539,N_1818);
or U2185 (N_2185,N_1732,N_1884);
nor U2186 (N_2186,N_1526,N_1886);
nand U2187 (N_2187,N_1782,N_1851);
nor U2188 (N_2188,N_1811,N_1981);
and U2189 (N_2189,N_1871,N_1832);
and U2190 (N_2190,N_1796,N_1776);
or U2191 (N_2191,N_1547,N_1985);
and U2192 (N_2192,N_1801,N_1861);
nand U2193 (N_2193,N_1657,N_1971);
and U2194 (N_2194,N_1563,N_1916);
nor U2195 (N_2195,N_1543,N_1616);
or U2196 (N_2196,N_1525,N_1632);
or U2197 (N_2197,N_1733,N_1531);
nor U2198 (N_2198,N_1510,N_1901);
or U2199 (N_2199,N_1710,N_1835);
or U2200 (N_2200,N_1918,N_1932);
or U2201 (N_2201,N_1997,N_1984);
and U2202 (N_2202,N_1797,N_1696);
or U2203 (N_2203,N_1953,N_1790);
nor U2204 (N_2204,N_1683,N_1989);
nor U2205 (N_2205,N_1620,N_1680);
or U2206 (N_2206,N_1653,N_1766);
nand U2207 (N_2207,N_1914,N_1775);
nand U2208 (N_2208,N_1640,N_1619);
nor U2209 (N_2209,N_1602,N_1815);
or U2210 (N_2210,N_1828,N_1638);
and U2211 (N_2211,N_1999,N_1659);
or U2212 (N_2212,N_1658,N_1909);
nor U2213 (N_2213,N_1694,N_1735);
nand U2214 (N_2214,N_1701,N_1824);
nor U2215 (N_2215,N_1813,N_1571);
nor U2216 (N_2216,N_1905,N_1929);
and U2217 (N_2217,N_1569,N_1895);
nor U2218 (N_2218,N_1928,N_1982);
nor U2219 (N_2219,N_1854,N_1557);
nor U2220 (N_2220,N_1726,N_1661);
or U2221 (N_2221,N_1974,N_1872);
nand U2222 (N_2222,N_1896,N_1729);
nor U2223 (N_2223,N_1848,N_1924);
nand U2224 (N_2224,N_1819,N_1591);
nand U2225 (N_2225,N_1867,N_1644);
and U2226 (N_2226,N_1684,N_1903);
nand U2227 (N_2227,N_1913,N_1634);
and U2228 (N_2228,N_1806,N_1778);
nand U2229 (N_2229,N_1688,N_1514);
nor U2230 (N_2230,N_1609,N_1962);
nor U2231 (N_2231,N_1503,N_1910);
and U2232 (N_2232,N_1686,N_1772);
nand U2233 (N_2233,N_1956,N_1666);
or U2234 (N_2234,N_1779,N_1940);
nand U2235 (N_2235,N_1737,N_1745);
xor U2236 (N_2236,N_1915,N_1769);
or U2237 (N_2237,N_1764,N_1821);
nor U2238 (N_2238,N_1585,N_1509);
and U2239 (N_2239,N_1548,N_1869);
nand U2240 (N_2240,N_1541,N_1559);
or U2241 (N_2241,N_1663,N_1662);
or U2242 (N_2242,N_1532,N_1767);
or U2243 (N_2243,N_1876,N_1942);
nor U2244 (N_2244,N_1893,N_1665);
or U2245 (N_2245,N_1529,N_1762);
or U2246 (N_2246,N_1756,N_1995);
nand U2247 (N_2247,N_1535,N_1566);
nand U2248 (N_2248,N_1507,N_1961);
or U2249 (N_2249,N_1612,N_1603);
nand U2250 (N_2250,N_1820,N_1910);
nand U2251 (N_2251,N_1639,N_1896);
and U2252 (N_2252,N_1710,N_1847);
and U2253 (N_2253,N_1864,N_1787);
or U2254 (N_2254,N_1571,N_1720);
or U2255 (N_2255,N_1856,N_1569);
or U2256 (N_2256,N_1830,N_1949);
nand U2257 (N_2257,N_1696,N_1775);
or U2258 (N_2258,N_1514,N_1789);
and U2259 (N_2259,N_1561,N_1631);
or U2260 (N_2260,N_1882,N_1651);
and U2261 (N_2261,N_1590,N_1807);
and U2262 (N_2262,N_1883,N_1769);
nand U2263 (N_2263,N_1670,N_1767);
nand U2264 (N_2264,N_1545,N_1920);
and U2265 (N_2265,N_1582,N_1754);
nor U2266 (N_2266,N_1800,N_1942);
nand U2267 (N_2267,N_1814,N_1595);
or U2268 (N_2268,N_1695,N_1801);
or U2269 (N_2269,N_1988,N_1823);
nor U2270 (N_2270,N_1638,N_1603);
nand U2271 (N_2271,N_1685,N_1866);
and U2272 (N_2272,N_1593,N_1754);
nand U2273 (N_2273,N_1642,N_1605);
nor U2274 (N_2274,N_1720,N_1659);
nand U2275 (N_2275,N_1874,N_1937);
or U2276 (N_2276,N_1540,N_1937);
nor U2277 (N_2277,N_1626,N_1895);
nand U2278 (N_2278,N_1973,N_1588);
nand U2279 (N_2279,N_1975,N_1883);
and U2280 (N_2280,N_1647,N_1994);
nor U2281 (N_2281,N_1648,N_1520);
and U2282 (N_2282,N_1962,N_1882);
or U2283 (N_2283,N_1720,N_1940);
xnor U2284 (N_2284,N_1699,N_1921);
nor U2285 (N_2285,N_1502,N_1896);
or U2286 (N_2286,N_1566,N_1528);
nor U2287 (N_2287,N_1813,N_1686);
or U2288 (N_2288,N_1583,N_1841);
nand U2289 (N_2289,N_1962,N_1596);
nand U2290 (N_2290,N_1550,N_1740);
nand U2291 (N_2291,N_1715,N_1691);
and U2292 (N_2292,N_1611,N_1709);
nor U2293 (N_2293,N_1826,N_1978);
and U2294 (N_2294,N_1590,N_1688);
xnor U2295 (N_2295,N_1713,N_1716);
or U2296 (N_2296,N_1668,N_1504);
and U2297 (N_2297,N_1875,N_1941);
nand U2298 (N_2298,N_1979,N_1767);
and U2299 (N_2299,N_1916,N_1976);
or U2300 (N_2300,N_1761,N_1645);
nor U2301 (N_2301,N_1504,N_1818);
or U2302 (N_2302,N_1996,N_1787);
nand U2303 (N_2303,N_1828,N_1518);
and U2304 (N_2304,N_1586,N_1788);
and U2305 (N_2305,N_1986,N_1831);
and U2306 (N_2306,N_1924,N_1726);
or U2307 (N_2307,N_1935,N_1658);
nor U2308 (N_2308,N_1887,N_1863);
nor U2309 (N_2309,N_1693,N_1736);
nor U2310 (N_2310,N_1581,N_1769);
nand U2311 (N_2311,N_1927,N_1883);
and U2312 (N_2312,N_1897,N_1775);
nor U2313 (N_2313,N_1826,N_1714);
nand U2314 (N_2314,N_1940,N_1570);
or U2315 (N_2315,N_1951,N_1730);
or U2316 (N_2316,N_1659,N_1821);
and U2317 (N_2317,N_1843,N_1556);
nor U2318 (N_2318,N_1744,N_1507);
and U2319 (N_2319,N_1937,N_1609);
nor U2320 (N_2320,N_1917,N_1976);
and U2321 (N_2321,N_1553,N_1819);
nor U2322 (N_2322,N_1572,N_1863);
nand U2323 (N_2323,N_1754,N_1589);
and U2324 (N_2324,N_1878,N_1980);
nand U2325 (N_2325,N_1993,N_1542);
or U2326 (N_2326,N_1782,N_1552);
nand U2327 (N_2327,N_1515,N_1926);
and U2328 (N_2328,N_1850,N_1888);
nor U2329 (N_2329,N_1720,N_1508);
xor U2330 (N_2330,N_1632,N_1722);
nor U2331 (N_2331,N_1600,N_1755);
and U2332 (N_2332,N_1557,N_1653);
nor U2333 (N_2333,N_1814,N_1573);
or U2334 (N_2334,N_1986,N_1894);
or U2335 (N_2335,N_1517,N_1739);
and U2336 (N_2336,N_1887,N_1590);
and U2337 (N_2337,N_1966,N_1619);
nand U2338 (N_2338,N_1943,N_1624);
xor U2339 (N_2339,N_1630,N_1534);
and U2340 (N_2340,N_1931,N_1961);
nand U2341 (N_2341,N_1883,N_1667);
or U2342 (N_2342,N_1584,N_1923);
nor U2343 (N_2343,N_1629,N_1979);
and U2344 (N_2344,N_1700,N_1522);
nor U2345 (N_2345,N_1642,N_1816);
and U2346 (N_2346,N_1729,N_1775);
nor U2347 (N_2347,N_1991,N_1989);
nor U2348 (N_2348,N_1578,N_1672);
nor U2349 (N_2349,N_1823,N_1838);
nor U2350 (N_2350,N_1802,N_1910);
nand U2351 (N_2351,N_1746,N_1632);
nand U2352 (N_2352,N_1675,N_1976);
nand U2353 (N_2353,N_1882,N_1843);
or U2354 (N_2354,N_1792,N_1694);
or U2355 (N_2355,N_1842,N_1718);
nand U2356 (N_2356,N_1798,N_1500);
nand U2357 (N_2357,N_1559,N_1621);
or U2358 (N_2358,N_1998,N_1661);
nand U2359 (N_2359,N_1864,N_1789);
and U2360 (N_2360,N_1899,N_1520);
nor U2361 (N_2361,N_1580,N_1650);
nor U2362 (N_2362,N_1899,N_1952);
and U2363 (N_2363,N_1804,N_1907);
nand U2364 (N_2364,N_1533,N_1957);
nor U2365 (N_2365,N_1650,N_1524);
or U2366 (N_2366,N_1615,N_1513);
and U2367 (N_2367,N_1932,N_1922);
nor U2368 (N_2368,N_1625,N_1585);
or U2369 (N_2369,N_1619,N_1995);
or U2370 (N_2370,N_1548,N_1912);
or U2371 (N_2371,N_1977,N_1958);
nor U2372 (N_2372,N_1607,N_1727);
and U2373 (N_2373,N_1738,N_1626);
and U2374 (N_2374,N_1585,N_1647);
nand U2375 (N_2375,N_1877,N_1817);
or U2376 (N_2376,N_1819,N_1824);
or U2377 (N_2377,N_1606,N_1738);
nand U2378 (N_2378,N_1632,N_1833);
nor U2379 (N_2379,N_1611,N_1995);
and U2380 (N_2380,N_1987,N_1544);
or U2381 (N_2381,N_1874,N_1500);
nor U2382 (N_2382,N_1843,N_1676);
or U2383 (N_2383,N_1948,N_1974);
or U2384 (N_2384,N_1836,N_1817);
and U2385 (N_2385,N_1697,N_1563);
nand U2386 (N_2386,N_1900,N_1899);
and U2387 (N_2387,N_1579,N_1622);
or U2388 (N_2388,N_1657,N_1849);
or U2389 (N_2389,N_1790,N_1873);
nor U2390 (N_2390,N_1660,N_1673);
nor U2391 (N_2391,N_1874,N_1597);
and U2392 (N_2392,N_1551,N_1890);
and U2393 (N_2393,N_1705,N_1901);
nor U2394 (N_2394,N_1714,N_1829);
and U2395 (N_2395,N_1853,N_1519);
or U2396 (N_2396,N_1516,N_1773);
xnor U2397 (N_2397,N_1552,N_1715);
and U2398 (N_2398,N_1944,N_1842);
and U2399 (N_2399,N_1565,N_1987);
nand U2400 (N_2400,N_1502,N_1596);
nand U2401 (N_2401,N_1695,N_1670);
or U2402 (N_2402,N_1831,N_1510);
nand U2403 (N_2403,N_1598,N_1924);
nand U2404 (N_2404,N_1552,N_1947);
or U2405 (N_2405,N_1591,N_1929);
nor U2406 (N_2406,N_1964,N_1836);
nand U2407 (N_2407,N_1979,N_1936);
and U2408 (N_2408,N_1927,N_1773);
or U2409 (N_2409,N_1850,N_1655);
and U2410 (N_2410,N_1760,N_1603);
and U2411 (N_2411,N_1838,N_1729);
and U2412 (N_2412,N_1826,N_1739);
or U2413 (N_2413,N_1600,N_1848);
nand U2414 (N_2414,N_1852,N_1572);
and U2415 (N_2415,N_1646,N_1814);
or U2416 (N_2416,N_1538,N_1531);
nor U2417 (N_2417,N_1968,N_1598);
or U2418 (N_2418,N_1705,N_1752);
and U2419 (N_2419,N_1811,N_1911);
xnor U2420 (N_2420,N_1807,N_1556);
or U2421 (N_2421,N_1769,N_1744);
or U2422 (N_2422,N_1676,N_1582);
nor U2423 (N_2423,N_1831,N_1790);
nor U2424 (N_2424,N_1648,N_1729);
nand U2425 (N_2425,N_1748,N_1707);
nand U2426 (N_2426,N_1591,N_1909);
and U2427 (N_2427,N_1851,N_1691);
xnor U2428 (N_2428,N_1779,N_1706);
nor U2429 (N_2429,N_1652,N_1871);
nor U2430 (N_2430,N_1869,N_1653);
nand U2431 (N_2431,N_1833,N_1929);
and U2432 (N_2432,N_1782,N_1919);
or U2433 (N_2433,N_1524,N_1520);
nand U2434 (N_2434,N_1795,N_1716);
nand U2435 (N_2435,N_1625,N_1888);
nand U2436 (N_2436,N_1585,N_1715);
and U2437 (N_2437,N_1872,N_1573);
or U2438 (N_2438,N_1535,N_1704);
nand U2439 (N_2439,N_1894,N_1805);
nand U2440 (N_2440,N_1566,N_1639);
nand U2441 (N_2441,N_1632,N_1675);
nor U2442 (N_2442,N_1745,N_1522);
and U2443 (N_2443,N_1557,N_1600);
nor U2444 (N_2444,N_1944,N_1872);
xor U2445 (N_2445,N_1857,N_1848);
and U2446 (N_2446,N_1836,N_1652);
nand U2447 (N_2447,N_1719,N_1707);
or U2448 (N_2448,N_1541,N_1723);
nand U2449 (N_2449,N_1651,N_1535);
or U2450 (N_2450,N_1645,N_1969);
or U2451 (N_2451,N_1822,N_1536);
nor U2452 (N_2452,N_1983,N_1933);
and U2453 (N_2453,N_1631,N_1958);
or U2454 (N_2454,N_1744,N_1937);
and U2455 (N_2455,N_1836,N_1828);
nor U2456 (N_2456,N_1839,N_1797);
xnor U2457 (N_2457,N_1735,N_1766);
nand U2458 (N_2458,N_1873,N_1677);
or U2459 (N_2459,N_1519,N_1807);
and U2460 (N_2460,N_1733,N_1925);
nand U2461 (N_2461,N_1776,N_1671);
or U2462 (N_2462,N_1952,N_1914);
or U2463 (N_2463,N_1957,N_1766);
nor U2464 (N_2464,N_1690,N_1753);
nand U2465 (N_2465,N_1796,N_1506);
and U2466 (N_2466,N_1783,N_1850);
nand U2467 (N_2467,N_1689,N_1633);
xor U2468 (N_2468,N_1691,N_1871);
or U2469 (N_2469,N_1639,N_1575);
nand U2470 (N_2470,N_1520,N_1712);
nor U2471 (N_2471,N_1597,N_1836);
nand U2472 (N_2472,N_1899,N_1815);
nor U2473 (N_2473,N_1847,N_1777);
nor U2474 (N_2474,N_1626,N_1710);
nor U2475 (N_2475,N_1672,N_1934);
nor U2476 (N_2476,N_1985,N_1515);
nor U2477 (N_2477,N_1801,N_1908);
or U2478 (N_2478,N_1708,N_1531);
and U2479 (N_2479,N_1927,N_1648);
or U2480 (N_2480,N_1987,N_1514);
and U2481 (N_2481,N_1693,N_1703);
nand U2482 (N_2482,N_1563,N_1596);
or U2483 (N_2483,N_1692,N_1697);
and U2484 (N_2484,N_1649,N_1753);
nor U2485 (N_2485,N_1668,N_1656);
nor U2486 (N_2486,N_1934,N_1925);
and U2487 (N_2487,N_1990,N_1756);
or U2488 (N_2488,N_1744,N_1787);
nor U2489 (N_2489,N_1621,N_1597);
nor U2490 (N_2490,N_1655,N_1963);
or U2491 (N_2491,N_1599,N_1919);
nand U2492 (N_2492,N_1957,N_1657);
or U2493 (N_2493,N_1943,N_1508);
nor U2494 (N_2494,N_1728,N_1599);
nor U2495 (N_2495,N_1926,N_1778);
nand U2496 (N_2496,N_1911,N_1662);
nand U2497 (N_2497,N_1598,N_1951);
nand U2498 (N_2498,N_1826,N_1804);
nor U2499 (N_2499,N_1993,N_1868);
or U2500 (N_2500,N_2429,N_2268);
nor U2501 (N_2501,N_2065,N_2369);
and U2502 (N_2502,N_2491,N_2127);
nand U2503 (N_2503,N_2138,N_2171);
nor U2504 (N_2504,N_2010,N_2099);
nor U2505 (N_2505,N_2176,N_2359);
and U2506 (N_2506,N_2451,N_2348);
and U2507 (N_2507,N_2363,N_2011);
nand U2508 (N_2508,N_2102,N_2088);
and U2509 (N_2509,N_2421,N_2150);
or U2510 (N_2510,N_2175,N_2492);
nor U2511 (N_2511,N_2228,N_2391);
and U2512 (N_2512,N_2213,N_2202);
nor U2513 (N_2513,N_2301,N_2195);
nor U2514 (N_2514,N_2241,N_2459);
and U2515 (N_2515,N_2232,N_2427);
nand U2516 (N_2516,N_2340,N_2154);
or U2517 (N_2517,N_2333,N_2013);
or U2518 (N_2518,N_2172,N_2380);
nand U2519 (N_2519,N_2223,N_2186);
nand U2520 (N_2520,N_2394,N_2456);
and U2521 (N_2521,N_2418,N_2049);
nor U2522 (N_2522,N_2270,N_2033);
and U2523 (N_2523,N_2306,N_2239);
or U2524 (N_2524,N_2177,N_2317);
nand U2525 (N_2525,N_2260,N_2300);
nand U2526 (N_2526,N_2145,N_2471);
xor U2527 (N_2527,N_2080,N_2235);
nor U2528 (N_2528,N_2203,N_2252);
nor U2529 (N_2529,N_2346,N_2409);
nor U2530 (N_2530,N_2162,N_2225);
and U2531 (N_2531,N_2424,N_2056);
and U2532 (N_2532,N_2042,N_2321);
or U2533 (N_2533,N_2337,N_2255);
nor U2534 (N_2534,N_2237,N_2123);
xor U2535 (N_2535,N_2121,N_2018);
nand U2536 (N_2536,N_2478,N_2152);
nand U2537 (N_2537,N_2179,N_2373);
and U2538 (N_2538,N_2231,N_2496);
and U2539 (N_2539,N_2097,N_2227);
and U2540 (N_2540,N_2430,N_2111);
or U2541 (N_2541,N_2151,N_2081);
and U2542 (N_2542,N_2307,N_2417);
and U2543 (N_2543,N_2003,N_2262);
xnor U2544 (N_2544,N_2020,N_2000);
or U2545 (N_2545,N_2073,N_2328);
nand U2546 (N_2546,N_2170,N_2209);
nand U2547 (N_2547,N_2071,N_2050);
nand U2548 (N_2548,N_2182,N_2426);
nand U2549 (N_2549,N_2038,N_2113);
nand U2550 (N_2550,N_2057,N_2193);
or U2551 (N_2551,N_2083,N_2282);
or U2552 (N_2552,N_2105,N_2037);
or U2553 (N_2553,N_2462,N_2481);
nand U2554 (N_2554,N_2035,N_2469);
or U2555 (N_2555,N_2399,N_2324);
or U2556 (N_2556,N_2461,N_2101);
and U2557 (N_2557,N_2400,N_2008);
and U2558 (N_2558,N_2433,N_2410);
nor U2559 (N_2559,N_2398,N_2141);
nor U2560 (N_2560,N_2063,N_2485);
or U2561 (N_2561,N_2377,N_2210);
nor U2562 (N_2562,N_2201,N_2499);
nand U2563 (N_2563,N_2279,N_2070);
and U2564 (N_2564,N_2126,N_2115);
nor U2565 (N_2565,N_2079,N_2110);
or U2566 (N_2566,N_2293,N_2173);
nor U2567 (N_2567,N_2296,N_2072);
nor U2568 (N_2568,N_2207,N_2100);
nor U2569 (N_2569,N_2382,N_2303);
and U2570 (N_2570,N_2261,N_2157);
and U2571 (N_2571,N_2388,N_2124);
or U2572 (N_2572,N_2236,N_2197);
nand U2573 (N_2573,N_2187,N_2455);
or U2574 (N_2574,N_2159,N_2169);
or U2575 (N_2575,N_2017,N_2278);
xor U2576 (N_2576,N_2016,N_2449);
nor U2577 (N_2577,N_2158,N_2006);
nor U2578 (N_2578,N_2022,N_2474);
nand U2579 (N_2579,N_2198,N_2498);
nand U2580 (N_2580,N_2160,N_2423);
nand U2581 (N_2581,N_2224,N_2025);
nand U2582 (N_2582,N_2468,N_2392);
or U2583 (N_2583,N_2362,N_2036);
nand U2584 (N_2584,N_2336,N_2298);
nand U2585 (N_2585,N_2415,N_2411);
and U2586 (N_2586,N_2463,N_2047);
or U2587 (N_2587,N_2334,N_2311);
nor U2588 (N_2588,N_2167,N_2457);
or U2589 (N_2589,N_2351,N_2316);
xnor U2590 (N_2590,N_2387,N_2304);
or U2591 (N_2591,N_2078,N_2059);
xor U2592 (N_2592,N_2218,N_2275);
nor U2593 (N_2593,N_2092,N_2444);
or U2594 (N_2594,N_2386,N_2132);
nand U2595 (N_2595,N_2361,N_2133);
nand U2596 (N_2596,N_2031,N_2039);
or U2597 (N_2597,N_2299,N_2199);
or U2598 (N_2598,N_2030,N_2371);
xnor U2599 (N_2599,N_2318,N_2486);
nor U2600 (N_2600,N_2226,N_2453);
or U2601 (N_2601,N_2390,N_2314);
and U2602 (N_2602,N_2263,N_2289);
nand U2603 (N_2603,N_2470,N_2290);
nand U2604 (N_2604,N_2412,N_2434);
nor U2605 (N_2605,N_2479,N_2309);
nand U2606 (N_2606,N_2093,N_2122);
or U2607 (N_2607,N_2185,N_2165);
and U2608 (N_2608,N_2029,N_2229);
nor U2609 (N_2609,N_2295,N_2366);
nand U2610 (N_2610,N_2472,N_2385);
nand U2611 (N_2611,N_2403,N_2118);
and U2612 (N_2612,N_2266,N_2048);
and U2613 (N_2613,N_2054,N_2188);
or U2614 (N_2614,N_2082,N_2248);
or U2615 (N_2615,N_2383,N_2443);
and U2616 (N_2616,N_2393,N_2350);
or U2617 (N_2617,N_2490,N_2313);
and U2618 (N_2618,N_2024,N_2149);
or U2619 (N_2619,N_2086,N_2397);
and U2620 (N_2620,N_2040,N_2114);
nor U2621 (N_2621,N_2484,N_2445);
or U2622 (N_2622,N_2379,N_2352);
and U2623 (N_2623,N_2338,N_2108);
xnor U2624 (N_2624,N_2284,N_2436);
and U2625 (N_2625,N_2343,N_2005);
or U2626 (N_2626,N_2345,N_2422);
nor U2627 (N_2627,N_2137,N_2274);
nor U2628 (N_2628,N_2211,N_2161);
nand U2629 (N_2629,N_2208,N_2250);
or U2630 (N_2630,N_2358,N_2075);
and U2631 (N_2631,N_2001,N_2272);
nor U2632 (N_2632,N_2089,N_2367);
and U2633 (N_2633,N_2058,N_2032);
nand U2634 (N_2634,N_2251,N_2384);
or U2635 (N_2635,N_2117,N_2212);
nand U2636 (N_2636,N_2407,N_2319);
nand U2637 (N_2637,N_2476,N_2026);
xnor U2638 (N_2638,N_2448,N_2046);
or U2639 (N_2639,N_2045,N_2475);
or U2640 (N_2640,N_2204,N_2090);
or U2641 (N_2641,N_2192,N_2164);
or U2642 (N_2642,N_2220,N_2216);
or U2643 (N_2643,N_2104,N_2419);
nor U2644 (N_2644,N_2374,N_2437);
nand U2645 (N_2645,N_2023,N_2349);
nor U2646 (N_2646,N_2277,N_2327);
or U2647 (N_2647,N_2180,N_2254);
or U2648 (N_2648,N_2466,N_2068);
or U2649 (N_2649,N_2129,N_2473);
nand U2650 (N_2650,N_2420,N_2178);
or U2651 (N_2651,N_2458,N_2493);
and U2652 (N_2652,N_2215,N_2428);
and U2653 (N_2653,N_2431,N_2283);
and U2654 (N_2654,N_2087,N_2310);
and U2655 (N_2655,N_2134,N_2249);
nor U2656 (N_2656,N_2234,N_2253);
and U2657 (N_2657,N_2136,N_2246);
nand U2658 (N_2658,N_2294,N_2357);
nand U2659 (N_2659,N_2140,N_2495);
and U2660 (N_2660,N_2144,N_2214);
and U2661 (N_2661,N_2323,N_2480);
nor U2662 (N_2662,N_2244,N_2467);
nand U2663 (N_2663,N_2460,N_2389);
or U2664 (N_2664,N_2413,N_2406);
nand U2665 (N_2665,N_2009,N_2168);
nand U2666 (N_2666,N_2489,N_2191);
nand U2667 (N_2667,N_2146,N_2330);
nor U2668 (N_2668,N_2356,N_2265);
nand U2669 (N_2669,N_2217,N_2103);
or U2670 (N_2670,N_2256,N_2372);
nand U2671 (N_2671,N_2085,N_2014);
xnor U2672 (N_2672,N_2194,N_2242);
or U2673 (N_2673,N_2074,N_2095);
nand U2674 (N_2674,N_2130,N_2332);
nor U2675 (N_2675,N_2062,N_2452);
and U2676 (N_2676,N_2052,N_2286);
nand U2677 (N_2677,N_2408,N_2183);
nor U2678 (N_2678,N_2135,N_2401);
nor U2679 (N_2679,N_2028,N_2375);
nand U2680 (N_2680,N_2477,N_2106);
and U2681 (N_2681,N_2305,N_2331);
nor U2682 (N_2682,N_2432,N_2425);
and U2683 (N_2683,N_2271,N_2112);
and U2684 (N_2684,N_2076,N_2339);
nand U2685 (N_2685,N_2258,N_2354);
nor U2686 (N_2686,N_2219,N_2245);
and U2687 (N_2687,N_2240,N_2004);
nor U2688 (N_2688,N_2094,N_2405);
and U2689 (N_2689,N_2131,N_2053);
or U2690 (N_2690,N_2402,N_2497);
or U2691 (N_2691,N_2153,N_2494);
and U2692 (N_2692,N_2381,N_2291);
nor U2693 (N_2693,N_2320,N_2069);
and U2694 (N_2694,N_2007,N_2273);
or U2695 (N_2695,N_2055,N_2347);
and U2696 (N_2696,N_2044,N_2125);
or U2697 (N_2697,N_2483,N_2156);
nand U2698 (N_2698,N_2096,N_2155);
or U2699 (N_2699,N_2259,N_2163);
or U2700 (N_2700,N_2342,N_2285);
nor U2701 (N_2701,N_2378,N_2396);
or U2702 (N_2702,N_2465,N_2438);
xnor U2703 (N_2703,N_2308,N_2142);
and U2704 (N_2704,N_2190,N_2442);
or U2705 (N_2705,N_2454,N_2148);
nand U2706 (N_2706,N_2482,N_2368);
or U2707 (N_2707,N_2181,N_2435);
nor U2708 (N_2708,N_2002,N_2395);
nand U2709 (N_2709,N_2206,N_2109);
nor U2710 (N_2710,N_2404,N_2312);
or U2711 (N_2711,N_2064,N_2043);
nand U2712 (N_2712,N_2128,N_2416);
nor U2713 (N_2713,N_2267,N_2205);
and U2714 (N_2714,N_2264,N_2322);
nand U2715 (N_2715,N_2166,N_2370);
nor U2716 (N_2716,N_2439,N_2288);
or U2717 (N_2717,N_2200,N_2021);
or U2718 (N_2718,N_2184,N_2281);
nor U2719 (N_2719,N_2066,N_2341);
or U2720 (N_2720,N_2297,N_2287);
nand U2721 (N_2721,N_2143,N_2302);
xnor U2722 (N_2722,N_2139,N_2376);
nor U2723 (N_2723,N_2189,N_2441);
nand U2724 (N_2724,N_2326,N_2243);
or U2725 (N_2725,N_2067,N_2034);
and U2726 (N_2726,N_2488,N_2257);
or U2727 (N_2727,N_2091,N_2174);
nor U2728 (N_2728,N_2353,N_2450);
or U2729 (N_2729,N_2222,N_2051);
or U2730 (N_2730,N_2464,N_2447);
nand U2731 (N_2731,N_2027,N_2098);
and U2732 (N_2732,N_2233,N_2280);
and U2733 (N_2733,N_2355,N_2414);
nand U2734 (N_2734,N_2325,N_2292);
nand U2735 (N_2735,N_2147,N_2360);
or U2736 (N_2736,N_2060,N_2364);
nor U2737 (N_2737,N_2344,N_2315);
or U2738 (N_2738,N_2487,N_2440);
xnor U2739 (N_2739,N_2041,N_2276);
or U2740 (N_2740,N_2119,N_2077);
or U2741 (N_2741,N_2015,N_2107);
or U2742 (N_2742,N_2230,N_2116);
or U2743 (N_2743,N_2329,N_2061);
nor U2744 (N_2744,N_2084,N_2221);
nor U2745 (N_2745,N_2120,N_2269);
or U2746 (N_2746,N_2365,N_2019);
or U2747 (N_2747,N_2335,N_2196);
nand U2748 (N_2748,N_2446,N_2238);
and U2749 (N_2749,N_2247,N_2012);
or U2750 (N_2750,N_2339,N_2489);
and U2751 (N_2751,N_2008,N_2061);
nand U2752 (N_2752,N_2287,N_2461);
nor U2753 (N_2753,N_2020,N_2214);
nor U2754 (N_2754,N_2041,N_2420);
and U2755 (N_2755,N_2183,N_2411);
nor U2756 (N_2756,N_2262,N_2223);
or U2757 (N_2757,N_2257,N_2059);
nor U2758 (N_2758,N_2159,N_2235);
or U2759 (N_2759,N_2434,N_2257);
and U2760 (N_2760,N_2498,N_2302);
nor U2761 (N_2761,N_2335,N_2373);
nor U2762 (N_2762,N_2467,N_2473);
or U2763 (N_2763,N_2171,N_2477);
or U2764 (N_2764,N_2352,N_2025);
or U2765 (N_2765,N_2481,N_2327);
or U2766 (N_2766,N_2120,N_2270);
nor U2767 (N_2767,N_2187,N_2371);
nand U2768 (N_2768,N_2397,N_2304);
or U2769 (N_2769,N_2051,N_2167);
xor U2770 (N_2770,N_2264,N_2170);
nor U2771 (N_2771,N_2241,N_2344);
or U2772 (N_2772,N_2047,N_2484);
or U2773 (N_2773,N_2046,N_2126);
and U2774 (N_2774,N_2002,N_2140);
nor U2775 (N_2775,N_2284,N_2058);
and U2776 (N_2776,N_2389,N_2355);
xor U2777 (N_2777,N_2307,N_2496);
nand U2778 (N_2778,N_2309,N_2226);
or U2779 (N_2779,N_2103,N_2128);
and U2780 (N_2780,N_2215,N_2367);
xnor U2781 (N_2781,N_2425,N_2186);
and U2782 (N_2782,N_2145,N_2127);
or U2783 (N_2783,N_2138,N_2491);
and U2784 (N_2784,N_2115,N_2311);
nand U2785 (N_2785,N_2439,N_2277);
nor U2786 (N_2786,N_2437,N_2431);
nand U2787 (N_2787,N_2358,N_2476);
xnor U2788 (N_2788,N_2274,N_2159);
nand U2789 (N_2789,N_2347,N_2146);
nand U2790 (N_2790,N_2180,N_2030);
and U2791 (N_2791,N_2016,N_2203);
nor U2792 (N_2792,N_2264,N_2144);
nor U2793 (N_2793,N_2007,N_2016);
or U2794 (N_2794,N_2164,N_2263);
nand U2795 (N_2795,N_2011,N_2415);
nor U2796 (N_2796,N_2284,N_2064);
nor U2797 (N_2797,N_2250,N_2140);
nor U2798 (N_2798,N_2126,N_2094);
or U2799 (N_2799,N_2231,N_2493);
nand U2800 (N_2800,N_2204,N_2195);
nor U2801 (N_2801,N_2242,N_2365);
nor U2802 (N_2802,N_2000,N_2070);
nand U2803 (N_2803,N_2221,N_2497);
or U2804 (N_2804,N_2113,N_2292);
and U2805 (N_2805,N_2263,N_2056);
or U2806 (N_2806,N_2476,N_2005);
nor U2807 (N_2807,N_2165,N_2000);
and U2808 (N_2808,N_2475,N_2082);
or U2809 (N_2809,N_2258,N_2039);
nor U2810 (N_2810,N_2234,N_2348);
and U2811 (N_2811,N_2133,N_2207);
nor U2812 (N_2812,N_2451,N_2179);
nor U2813 (N_2813,N_2112,N_2423);
nand U2814 (N_2814,N_2421,N_2305);
nor U2815 (N_2815,N_2338,N_2181);
or U2816 (N_2816,N_2217,N_2014);
nand U2817 (N_2817,N_2101,N_2321);
nor U2818 (N_2818,N_2386,N_2474);
or U2819 (N_2819,N_2105,N_2331);
and U2820 (N_2820,N_2199,N_2142);
and U2821 (N_2821,N_2439,N_2318);
nand U2822 (N_2822,N_2404,N_2456);
xnor U2823 (N_2823,N_2065,N_2061);
or U2824 (N_2824,N_2079,N_2450);
nand U2825 (N_2825,N_2353,N_2483);
and U2826 (N_2826,N_2331,N_2124);
nand U2827 (N_2827,N_2231,N_2337);
and U2828 (N_2828,N_2361,N_2320);
nor U2829 (N_2829,N_2486,N_2045);
or U2830 (N_2830,N_2121,N_2189);
nand U2831 (N_2831,N_2028,N_2401);
nand U2832 (N_2832,N_2163,N_2406);
and U2833 (N_2833,N_2335,N_2053);
nand U2834 (N_2834,N_2403,N_2255);
nand U2835 (N_2835,N_2214,N_2282);
xor U2836 (N_2836,N_2249,N_2216);
nor U2837 (N_2837,N_2182,N_2049);
nand U2838 (N_2838,N_2113,N_2228);
nand U2839 (N_2839,N_2019,N_2096);
nand U2840 (N_2840,N_2104,N_2084);
or U2841 (N_2841,N_2068,N_2070);
nand U2842 (N_2842,N_2496,N_2386);
and U2843 (N_2843,N_2097,N_2457);
and U2844 (N_2844,N_2163,N_2131);
nor U2845 (N_2845,N_2355,N_2262);
nand U2846 (N_2846,N_2082,N_2107);
nor U2847 (N_2847,N_2458,N_2041);
nor U2848 (N_2848,N_2470,N_2161);
nor U2849 (N_2849,N_2224,N_2413);
or U2850 (N_2850,N_2354,N_2186);
nand U2851 (N_2851,N_2090,N_2154);
and U2852 (N_2852,N_2009,N_2057);
or U2853 (N_2853,N_2042,N_2180);
nor U2854 (N_2854,N_2163,N_2191);
nor U2855 (N_2855,N_2204,N_2002);
and U2856 (N_2856,N_2250,N_2435);
nor U2857 (N_2857,N_2208,N_2338);
nand U2858 (N_2858,N_2419,N_2433);
nand U2859 (N_2859,N_2269,N_2315);
nor U2860 (N_2860,N_2442,N_2218);
nor U2861 (N_2861,N_2128,N_2443);
or U2862 (N_2862,N_2303,N_2129);
nand U2863 (N_2863,N_2448,N_2151);
nor U2864 (N_2864,N_2160,N_2266);
nor U2865 (N_2865,N_2196,N_2265);
and U2866 (N_2866,N_2291,N_2156);
nor U2867 (N_2867,N_2328,N_2048);
nand U2868 (N_2868,N_2487,N_2041);
or U2869 (N_2869,N_2418,N_2301);
or U2870 (N_2870,N_2288,N_2033);
nor U2871 (N_2871,N_2078,N_2418);
and U2872 (N_2872,N_2215,N_2268);
or U2873 (N_2873,N_2349,N_2100);
or U2874 (N_2874,N_2073,N_2083);
nor U2875 (N_2875,N_2244,N_2030);
and U2876 (N_2876,N_2452,N_2046);
nor U2877 (N_2877,N_2012,N_2214);
and U2878 (N_2878,N_2365,N_2043);
and U2879 (N_2879,N_2461,N_2422);
and U2880 (N_2880,N_2142,N_2419);
or U2881 (N_2881,N_2246,N_2108);
or U2882 (N_2882,N_2056,N_2259);
or U2883 (N_2883,N_2102,N_2128);
and U2884 (N_2884,N_2024,N_2011);
nor U2885 (N_2885,N_2241,N_2247);
or U2886 (N_2886,N_2346,N_2474);
and U2887 (N_2887,N_2442,N_2458);
nor U2888 (N_2888,N_2314,N_2110);
and U2889 (N_2889,N_2213,N_2176);
nand U2890 (N_2890,N_2381,N_2490);
and U2891 (N_2891,N_2049,N_2152);
nor U2892 (N_2892,N_2480,N_2117);
nand U2893 (N_2893,N_2243,N_2345);
and U2894 (N_2894,N_2216,N_2132);
or U2895 (N_2895,N_2315,N_2008);
and U2896 (N_2896,N_2289,N_2300);
xnor U2897 (N_2897,N_2353,N_2478);
and U2898 (N_2898,N_2294,N_2148);
nand U2899 (N_2899,N_2099,N_2455);
or U2900 (N_2900,N_2430,N_2016);
nand U2901 (N_2901,N_2061,N_2040);
or U2902 (N_2902,N_2287,N_2277);
and U2903 (N_2903,N_2046,N_2266);
or U2904 (N_2904,N_2331,N_2125);
or U2905 (N_2905,N_2395,N_2397);
nor U2906 (N_2906,N_2439,N_2047);
or U2907 (N_2907,N_2262,N_2374);
and U2908 (N_2908,N_2429,N_2176);
nor U2909 (N_2909,N_2416,N_2403);
or U2910 (N_2910,N_2223,N_2236);
nand U2911 (N_2911,N_2075,N_2237);
and U2912 (N_2912,N_2078,N_2037);
nand U2913 (N_2913,N_2117,N_2299);
or U2914 (N_2914,N_2073,N_2399);
nand U2915 (N_2915,N_2471,N_2339);
nor U2916 (N_2916,N_2206,N_2215);
or U2917 (N_2917,N_2360,N_2313);
nand U2918 (N_2918,N_2057,N_2385);
and U2919 (N_2919,N_2317,N_2079);
or U2920 (N_2920,N_2220,N_2047);
or U2921 (N_2921,N_2342,N_2184);
nor U2922 (N_2922,N_2197,N_2300);
or U2923 (N_2923,N_2052,N_2155);
or U2924 (N_2924,N_2345,N_2280);
nand U2925 (N_2925,N_2437,N_2492);
nand U2926 (N_2926,N_2073,N_2138);
and U2927 (N_2927,N_2192,N_2009);
nand U2928 (N_2928,N_2263,N_2053);
nand U2929 (N_2929,N_2073,N_2313);
and U2930 (N_2930,N_2146,N_2129);
or U2931 (N_2931,N_2064,N_2480);
nor U2932 (N_2932,N_2165,N_2302);
nand U2933 (N_2933,N_2063,N_2174);
and U2934 (N_2934,N_2419,N_2410);
nand U2935 (N_2935,N_2144,N_2335);
xor U2936 (N_2936,N_2289,N_2026);
nor U2937 (N_2937,N_2087,N_2159);
or U2938 (N_2938,N_2100,N_2146);
nand U2939 (N_2939,N_2400,N_2131);
and U2940 (N_2940,N_2322,N_2147);
nor U2941 (N_2941,N_2184,N_2492);
nor U2942 (N_2942,N_2359,N_2206);
nand U2943 (N_2943,N_2316,N_2037);
nor U2944 (N_2944,N_2206,N_2380);
or U2945 (N_2945,N_2444,N_2234);
and U2946 (N_2946,N_2012,N_2126);
and U2947 (N_2947,N_2186,N_2114);
and U2948 (N_2948,N_2066,N_2069);
nor U2949 (N_2949,N_2003,N_2190);
xor U2950 (N_2950,N_2091,N_2191);
nand U2951 (N_2951,N_2154,N_2215);
nor U2952 (N_2952,N_2209,N_2403);
and U2953 (N_2953,N_2207,N_2254);
nor U2954 (N_2954,N_2344,N_2051);
nand U2955 (N_2955,N_2006,N_2186);
nor U2956 (N_2956,N_2263,N_2407);
and U2957 (N_2957,N_2288,N_2350);
and U2958 (N_2958,N_2224,N_2296);
nand U2959 (N_2959,N_2448,N_2296);
nand U2960 (N_2960,N_2027,N_2462);
and U2961 (N_2961,N_2371,N_2210);
and U2962 (N_2962,N_2462,N_2482);
nor U2963 (N_2963,N_2416,N_2094);
nand U2964 (N_2964,N_2269,N_2387);
and U2965 (N_2965,N_2105,N_2221);
and U2966 (N_2966,N_2452,N_2287);
or U2967 (N_2967,N_2011,N_2303);
and U2968 (N_2968,N_2439,N_2464);
nor U2969 (N_2969,N_2205,N_2216);
nand U2970 (N_2970,N_2104,N_2371);
and U2971 (N_2971,N_2115,N_2145);
nor U2972 (N_2972,N_2468,N_2465);
and U2973 (N_2973,N_2293,N_2308);
nand U2974 (N_2974,N_2423,N_2072);
nor U2975 (N_2975,N_2201,N_2119);
nand U2976 (N_2976,N_2461,N_2459);
and U2977 (N_2977,N_2340,N_2263);
nor U2978 (N_2978,N_2053,N_2341);
or U2979 (N_2979,N_2215,N_2056);
and U2980 (N_2980,N_2221,N_2483);
nor U2981 (N_2981,N_2465,N_2498);
nor U2982 (N_2982,N_2233,N_2130);
or U2983 (N_2983,N_2286,N_2011);
nor U2984 (N_2984,N_2167,N_2169);
or U2985 (N_2985,N_2460,N_2373);
and U2986 (N_2986,N_2217,N_2050);
xor U2987 (N_2987,N_2090,N_2121);
nand U2988 (N_2988,N_2097,N_2432);
or U2989 (N_2989,N_2008,N_2412);
xnor U2990 (N_2990,N_2247,N_2153);
nor U2991 (N_2991,N_2291,N_2468);
nor U2992 (N_2992,N_2149,N_2228);
or U2993 (N_2993,N_2406,N_2155);
nand U2994 (N_2994,N_2289,N_2292);
nand U2995 (N_2995,N_2316,N_2448);
or U2996 (N_2996,N_2051,N_2070);
nor U2997 (N_2997,N_2194,N_2342);
nand U2998 (N_2998,N_2385,N_2270);
nand U2999 (N_2999,N_2128,N_2118);
nand U3000 (N_3000,N_2996,N_2979);
and U3001 (N_3001,N_2754,N_2552);
nand U3002 (N_3002,N_2941,N_2923);
nor U3003 (N_3003,N_2859,N_2560);
or U3004 (N_3004,N_2890,N_2659);
nand U3005 (N_3005,N_2947,N_2800);
nor U3006 (N_3006,N_2879,N_2648);
nor U3007 (N_3007,N_2866,N_2954);
nor U3008 (N_3008,N_2785,N_2778);
or U3009 (N_3009,N_2522,N_2776);
xnor U3010 (N_3010,N_2672,N_2640);
or U3011 (N_3011,N_2874,N_2861);
or U3012 (N_3012,N_2862,N_2809);
and U3013 (N_3013,N_2703,N_2747);
and U3014 (N_3014,N_2674,N_2810);
xor U3015 (N_3015,N_2592,N_2614);
nor U3016 (N_3016,N_2515,N_2737);
nand U3017 (N_3017,N_2511,N_2799);
or U3018 (N_3018,N_2624,N_2895);
and U3019 (N_3019,N_2958,N_2847);
and U3020 (N_3020,N_2584,N_2792);
nor U3021 (N_3021,N_2568,N_2531);
and U3022 (N_3022,N_2977,N_2884);
or U3023 (N_3023,N_2639,N_2543);
or U3024 (N_3024,N_2671,N_2616);
xor U3025 (N_3025,N_2816,N_2535);
or U3026 (N_3026,N_2723,N_2811);
or U3027 (N_3027,N_2873,N_2601);
nor U3028 (N_3028,N_2902,N_2605);
nand U3029 (N_3029,N_2891,N_2542);
and U3030 (N_3030,N_2870,N_2677);
and U3031 (N_3031,N_2911,N_2719);
and U3032 (N_3032,N_2732,N_2538);
nand U3033 (N_3033,N_2507,N_2990);
or U3034 (N_3034,N_2618,N_2924);
nor U3035 (N_3035,N_2652,N_2899);
nand U3036 (N_3036,N_2520,N_2836);
nand U3037 (N_3037,N_2706,N_2527);
or U3038 (N_3038,N_2968,N_2602);
nand U3039 (N_3039,N_2794,N_2583);
nand U3040 (N_3040,N_2917,N_2757);
nand U3041 (N_3041,N_2819,N_2502);
nor U3042 (N_3042,N_2830,N_2815);
or U3043 (N_3043,N_2980,N_2608);
and U3044 (N_3044,N_2994,N_2738);
nand U3045 (N_3045,N_2506,N_2715);
xor U3046 (N_3046,N_2777,N_2982);
nand U3047 (N_3047,N_2629,N_2525);
nand U3048 (N_3048,N_2883,N_2972);
nand U3049 (N_3049,N_2988,N_2822);
nand U3050 (N_3050,N_2854,N_2554);
nor U3051 (N_3051,N_2651,N_2563);
nand U3052 (N_3052,N_2852,N_2936);
or U3053 (N_3053,N_2905,N_2995);
nand U3054 (N_3054,N_2653,N_2536);
nand U3055 (N_3055,N_2551,N_2686);
and U3056 (N_3056,N_2705,N_2570);
nand U3057 (N_3057,N_2864,N_2802);
or U3058 (N_3058,N_2576,N_2888);
nor U3059 (N_3059,N_2661,N_2760);
nand U3060 (N_3060,N_2635,N_2939);
nand U3061 (N_3061,N_2665,N_2832);
or U3062 (N_3062,N_2505,N_2914);
and U3063 (N_3063,N_2827,N_2998);
nor U3064 (N_3064,N_2935,N_2675);
nand U3065 (N_3065,N_2553,N_2817);
nor U3066 (N_3066,N_2634,N_2965);
nor U3067 (N_3067,N_2581,N_2750);
and U3068 (N_3068,N_2627,N_2893);
or U3069 (N_3069,N_2641,N_2532);
and U3070 (N_3070,N_2868,N_2956);
nand U3071 (N_3071,N_2730,N_2633);
nand U3072 (N_3072,N_2781,N_2828);
or U3073 (N_3073,N_2670,N_2805);
nand U3074 (N_3074,N_2673,N_2925);
or U3075 (N_3075,N_2518,N_2562);
nor U3076 (N_3076,N_2892,N_2882);
or U3077 (N_3077,N_2609,N_2840);
or U3078 (N_3078,N_2950,N_2790);
and U3079 (N_3079,N_2743,N_2758);
nor U3080 (N_3080,N_2697,N_2572);
and U3081 (N_3081,N_2603,N_2713);
nand U3082 (N_3082,N_2595,N_2636);
and U3083 (N_3083,N_2824,N_2896);
nand U3084 (N_3084,N_2787,N_2749);
nand U3085 (N_3085,N_2692,N_2717);
and U3086 (N_3086,N_2643,N_2751);
or U3087 (N_3087,N_2959,N_2718);
or U3088 (N_3088,N_2875,N_2877);
or U3089 (N_3089,N_2617,N_2843);
and U3090 (N_3090,N_2786,N_2638);
or U3091 (N_3091,N_2733,N_2529);
nor U3092 (N_3092,N_2669,N_2649);
or U3093 (N_3093,N_2849,N_2752);
and U3094 (N_3094,N_2565,N_2517);
nand U3095 (N_3095,N_2789,N_2782);
nor U3096 (N_3096,N_2928,N_2657);
nand U3097 (N_3097,N_2756,N_2764);
nand U3098 (N_3098,N_2807,N_2918);
nor U3099 (N_3099,N_2586,N_2545);
nand U3100 (N_3100,N_2944,N_2714);
nand U3101 (N_3101,N_2927,N_2773);
nand U3102 (N_3102,N_2772,N_2647);
nand U3103 (N_3103,N_2908,N_2966);
or U3104 (N_3104,N_2667,N_2838);
xnor U3105 (N_3105,N_2587,N_2779);
or U3106 (N_3106,N_2798,N_2567);
nand U3107 (N_3107,N_2682,N_2655);
or U3108 (N_3108,N_2526,N_2770);
or U3109 (N_3109,N_2516,N_2963);
and U3110 (N_3110,N_2912,N_2981);
and U3111 (N_3111,N_2933,N_2630);
or U3112 (N_3112,N_2556,N_2696);
nor U3113 (N_3113,N_2729,N_2625);
or U3114 (N_3114,N_2755,N_2753);
or U3115 (N_3115,N_2740,N_2955);
nor U3116 (N_3116,N_2626,N_2727);
and U3117 (N_3117,N_2559,N_2558);
or U3118 (N_3118,N_2801,N_2916);
nand U3119 (N_3119,N_2930,N_2704);
and U3120 (N_3120,N_2537,N_2897);
and U3121 (N_3121,N_2793,N_2622);
nand U3122 (N_3122,N_2698,N_2604);
nor U3123 (N_3123,N_2620,N_2984);
nand U3124 (N_3124,N_2865,N_2970);
nand U3125 (N_3125,N_2846,N_2668);
nand U3126 (N_3126,N_2783,N_2579);
and U3127 (N_3127,N_2837,N_2871);
and U3128 (N_3128,N_2654,N_2631);
nor U3129 (N_3129,N_2961,N_2742);
nand U3130 (N_3130,N_2937,N_2549);
xnor U3131 (N_3131,N_2589,N_2615);
or U3132 (N_3132,N_2685,N_2858);
or U3133 (N_3133,N_2681,N_2948);
or U3134 (N_3134,N_2528,N_2722);
or U3135 (N_3135,N_2833,N_2876);
nand U3136 (N_3136,N_2748,N_2872);
nand U3137 (N_3137,N_2569,N_2845);
xor U3138 (N_3138,N_2744,N_2943);
and U3139 (N_3139,N_2775,N_2663);
and U3140 (N_3140,N_2960,N_2967);
nand U3141 (N_3141,N_2857,N_2946);
or U3142 (N_3142,N_2978,N_2664);
and U3143 (N_3143,N_2546,N_2901);
nor U3144 (N_3144,N_2796,N_2702);
or U3145 (N_3145,N_2683,N_2716);
nand U3146 (N_3146,N_2728,N_2774);
or U3147 (N_3147,N_2588,N_2596);
or U3148 (N_3148,N_2539,N_2619);
nor U3149 (N_3149,N_2880,N_2564);
nand U3150 (N_3150,N_2594,N_2574);
nand U3151 (N_3151,N_2920,N_2650);
nor U3152 (N_3152,N_2646,N_2841);
nand U3153 (N_3153,N_2989,N_2869);
and U3154 (N_3154,N_2662,N_2621);
nand U3155 (N_3155,N_2761,N_2940);
and U3156 (N_3156,N_2745,N_2711);
and U3157 (N_3157,N_2831,N_2985);
and U3158 (N_3158,N_2544,N_2577);
and U3159 (N_3159,N_2964,N_2855);
or U3160 (N_3160,N_2500,N_2573);
nor U3161 (N_3161,N_2886,N_2679);
and U3162 (N_3162,N_2910,N_2839);
nand U3163 (N_3163,N_2942,N_2741);
or U3164 (N_3164,N_2898,N_2922);
and U3165 (N_3165,N_2746,N_2524);
nor U3166 (N_3166,N_2680,N_2707);
or U3167 (N_3167,N_2550,N_2637);
and U3168 (N_3168,N_2504,N_2987);
and U3169 (N_3169,N_2628,N_2700);
nor U3170 (N_3170,N_2509,N_2823);
nand U3171 (N_3171,N_2540,N_2523);
or U3172 (N_3172,N_2991,N_2571);
nor U3173 (N_3173,N_2885,N_2533);
and U3174 (N_3174,N_2736,N_2771);
nor U3175 (N_3175,N_2557,N_2934);
and U3176 (N_3176,N_2561,N_2580);
and U3177 (N_3177,N_2971,N_2945);
xnor U3178 (N_3178,N_2709,N_2720);
and U3179 (N_3179,N_2784,N_2521);
nor U3180 (N_3180,N_2708,N_2766);
nor U3181 (N_3181,N_2607,N_2835);
and U3182 (N_3182,N_2606,N_2863);
nand U3183 (N_3183,N_2642,N_2814);
or U3184 (N_3184,N_2689,N_2795);
nand U3185 (N_3185,N_2694,N_2599);
and U3186 (N_3186,N_2804,N_2818);
or U3187 (N_3187,N_2623,N_2999);
or U3188 (N_3188,N_2514,N_2949);
and U3189 (N_3189,N_2725,N_2578);
or U3190 (N_3190,N_2699,N_2889);
and U3191 (N_3191,N_2701,N_2519);
and U3192 (N_3192,N_2585,N_2530);
and U3193 (N_3193,N_2821,N_2860);
or U3194 (N_3194,N_2907,N_2566);
nand U3195 (N_3195,N_2887,N_2951);
or U3196 (N_3196,N_2510,N_2878);
nor U3197 (N_3197,N_2900,N_2903);
nor U3198 (N_3198,N_2508,N_2691);
and U3199 (N_3199,N_2929,N_2534);
nor U3200 (N_3200,N_2938,N_2610);
and U3201 (N_3201,N_2894,N_2803);
or U3202 (N_3202,N_2932,N_2768);
nor U3203 (N_3203,N_2762,N_2695);
and U3204 (N_3204,N_2829,N_2921);
or U3205 (N_3205,N_2731,N_2913);
and U3206 (N_3206,N_2974,N_2598);
and U3207 (N_3207,N_2848,N_2856);
and U3208 (N_3208,N_2597,N_2844);
and U3209 (N_3209,N_2842,N_2780);
or U3210 (N_3210,N_2724,N_2660);
or U3211 (N_3211,N_2666,N_2658);
nand U3212 (N_3212,N_2788,N_2992);
nand U3213 (N_3213,N_2644,N_2541);
or U3214 (N_3214,N_2739,N_2765);
or U3215 (N_3215,N_2986,N_2993);
or U3216 (N_3216,N_2813,N_2611);
nor U3217 (N_3217,N_2976,N_2645);
nor U3218 (N_3218,N_2926,N_2904);
or U3219 (N_3219,N_2881,N_2632);
and U3220 (N_3220,N_2726,N_2759);
and U3221 (N_3221,N_2688,N_2676);
and U3222 (N_3222,N_2593,N_2975);
and U3223 (N_3223,N_2825,N_2710);
nor U3224 (N_3224,N_2769,N_2656);
or U3225 (N_3225,N_2555,N_2952);
or U3226 (N_3226,N_2767,N_2820);
nand U3227 (N_3227,N_2612,N_2953);
nand U3228 (N_3228,N_2791,N_2983);
and U3229 (N_3229,N_2806,N_2501);
nor U3230 (N_3230,N_2690,N_2906);
and U3231 (N_3231,N_2735,N_2853);
or U3232 (N_3232,N_2797,N_2851);
and U3233 (N_3233,N_2763,N_2915);
and U3234 (N_3234,N_2548,N_2721);
and U3235 (N_3235,N_2850,N_2812);
or U3236 (N_3236,N_2957,N_2687);
or U3237 (N_3237,N_2590,N_2867);
nor U3238 (N_3238,N_2808,N_2834);
and U3239 (N_3239,N_2591,N_2513);
nor U3240 (N_3240,N_2909,N_2931);
or U3241 (N_3241,N_2547,N_2582);
and U3242 (N_3242,N_2693,N_2575);
nand U3243 (N_3243,N_2969,N_2962);
nand U3244 (N_3244,N_2600,N_2712);
nor U3245 (N_3245,N_2678,N_2684);
nand U3246 (N_3246,N_2919,N_2503);
or U3247 (N_3247,N_2613,N_2997);
nand U3248 (N_3248,N_2512,N_2734);
nor U3249 (N_3249,N_2973,N_2826);
nand U3250 (N_3250,N_2756,N_2630);
or U3251 (N_3251,N_2773,N_2894);
or U3252 (N_3252,N_2602,N_2932);
nand U3253 (N_3253,N_2877,N_2781);
and U3254 (N_3254,N_2587,N_2885);
nand U3255 (N_3255,N_2994,N_2931);
nand U3256 (N_3256,N_2677,N_2674);
or U3257 (N_3257,N_2954,N_2710);
nand U3258 (N_3258,N_2892,N_2731);
or U3259 (N_3259,N_2546,N_2684);
nand U3260 (N_3260,N_2517,N_2759);
nor U3261 (N_3261,N_2515,N_2668);
xnor U3262 (N_3262,N_2946,N_2964);
or U3263 (N_3263,N_2514,N_2586);
and U3264 (N_3264,N_2861,N_2573);
nand U3265 (N_3265,N_2806,N_2841);
or U3266 (N_3266,N_2656,N_2549);
nor U3267 (N_3267,N_2776,N_2595);
nor U3268 (N_3268,N_2502,N_2550);
nor U3269 (N_3269,N_2635,N_2515);
nor U3270 (N_3270,N_2791,N_2943);
nand U3271 (N_3271,N_2780,N_2623);
or U3272 (N_3272,N_2816,N_2671);
and U3273 (N_3273,N_2901,N_2878);
and U3274 (N_3274,N_2920,N_2874);
or U3275 (N_3275,N_2584,N_2765);
and U3276 (N_3276,N_2836,N_2605);
and U3277 (N_3277,N_2856,N_2585);
and U3278 (N_3278,N_2748,N_2801);
and U3279 (N_3279,N_2597,N_2923);
or U3280 (N_3280,N_2937,N_2771);
nor U3281 (N_3281,N_2595,N_2534);
or U3282 (N_3282,N_2626,N_2970);
and U3283 (N_3283,N_2938,N_2764);
and U3284 (N_3284,N_2764,N_2917);
and U3285 (N_3285,N_2689,N_2608);
nand U3286 (N_3286,N_2728,N_2715);
or U3287 (N_3287,N_2561,N_2966);
or U3288 (N_3288,N_2581,N_2713);
or U3289 (N_3289,N_2817,N_2759);
nor U3290 (N_3290,N_2881,N_2856);
nor U3291 (N_3291,N_2693,N_2613);
nand U3292 (N_3292,N_2726,N_2697);
nor U3293 (N_3293,N_2737,N_2928);
nand U3294 (N_3294,N_2876,N_2822);
nor U3295 (N_3295,N_2742,N_2518);
nor U3296 (N_3296,N_2985,N_2513);
or U3297 (N_3297,N_2785,N_2839);
or U3298 (N_3298,N_2854,N_2858);
and U3299 (N_3299,N_2706,N_2643);
and U3300 (N_3300,N_2579,N_2916);
nor U3301 (N_3301,N_2624,N_2659);
and U3302 (N_3302,N_2660,N_2613);
nand U3303 (N_3303,N_2693,N_2809);
nor U3304 (N_3304,N_2872,N_2787);
nand U3305 (N_3305,N_2769,N_2659);
xor U3306 (N_3306,N_2648,N_2921);
and U3307 (N_3307,N_2736,N_2602);
nand U3308 (N_3308,N_2745,N_2676);
or U3309 (N_3309,N_2545,N_2662);
nor U3310 (N_3310,N_2582,N_2664);
and U3311 (N_3311,N_2530,N_2983);
or U3312 (N_3312,N_2893,N_2977);
nand U3313 (N_3313,N_2586,N_2782);
and U3314 (N_3314,N_2895,N_2718);
xor U3315 (N_3315,N_2600,N_2893);
nor U3316 (N_3316,N_2508,N_2822);
nor U3317 (N_3317,N_2638,N_2769);
or U3318 (N_3318,N_2691,N_2699);
nand U3319 (N_3319,N_2512,N_2843);
and U3320 (N_3320,N_2751,N_2726);
nand U3321 (N_3321,N_2879,N_2636);
or U3322 (N_3322,N_2512,N_2559);
and U3323 (N_3323,N_2706,N_2801);
or U3324 (N_3324,N_2861,N_2864);
or U3325 (N_3325,N_2733,N_2874);
nand U3326 (N_3326,N_2556,N_2633);
or U3327 (N_3327,N_2588,N_2839);
nand U3328 (N_3328,N_2559,N_2616);
and U3329 (N_3329,N_2981,N_2867);
or U3330 (N_3330,N_2981,N_2895);
and U3331 (N_3331,N_2795,N_2745);
and U3332 (N_3332,N_2981,N_2991);
nand U3333 (N_3333,N_2741,N_2752);
xnor U3334 (N_3334,N_2795,N_2915);
nor U3335 (N_3335,N_2591,N_2694);
nor U3336 (N_3336,N_2552,N_2773);
or U3337 (N_3337,N_2707,N_2705);
or U3338 (N_3338,N_2704,N_2556);
nor U3339 (N_3339,N_2590,N_2633);
and U3340 (N_3340,N_2863,N_2788);
or U3341 (N_3341,N_2749,N_2816);
nand U3342 (N_3342,N_2583,N_2566);
nand U3343 (N_3343,N_2629,N_2773);
or U3344 (N_3344,N_2971,N_2942);
nor U3345 (N_3345,N_2775,N_2922);
and U3346 (N_3346,N_2679,N_2801);
nor U3347 (N_3347,N_2916,N_2587);
nand U3348 (N_3348,N_2956,N_2705);
nand U3349 (N_3349,N_2638,N_2720);
and U3350 (N_3350,N_2682,N_2753);
and U3351 (N_3351,N_2573,N_2665);
nand U3352 (N_3352,N_2733,N_2868);
nand U3353 (N_3353,N_2814,N_2678);
nand U3354 (N_3354,N_2717,N_2956);
nand U3355 (N_3355,N_2829,N_2691);
or U3356 (N_3356,N_2619,N_2634);
and U3357 (N_3357,N_2818,N_2581);
or U3358 (N_3358,N_2961,N_2691);
nand U3359 (N_3359,N_2798,N_2917);
nor U3360 (N_3360,N_2738,N_2854);
nor U3361 (N_3361,N_2774,N_2897);
nor U3362 (N_3362,N_2983,N_2537);
and U3363 (N_3363,N_2868,N_2971);
nand U3364 (N_3364,N_2550,N_2737);
and U3365 (N_3365,N_2857,N_2668);
and U3366 (N_3366,N_2791,N_2688);
or U3367 (N_3367,N_2837,N_2901);
or U3368 (N_3368,N_2687,N_2594);
nand U3369 (N_3369,N_2714,N_2644);
and U3370 (N_3370,N_2865,N_2885);
nand U3371 (N_3371,N_2946,N_2630);
or U3372 (N_3372,N_2710,N_2906);
or U3373 (N_3373,N_2978,N_2659);
or U3374 (N_3374,N_2690,N_2637);
nor U3375 (N_3375,N_2998,N_2842);
or U3376 (N_3376,N_2567,N_2719);
nand U3377 (N_3377,N_2575,N_2991);
or U3378 (N_3378,N_2522,N_2845);
or U3379 (N_3379,N_2590,N_2526);
or U3380 (N_3380,N_2733,N_2748);
and U3381 (N_3381,N_2936,N_2733);
nand U3382 (N_3382,N_2840,N_2529);
nand U3383 (N_3383,N_2597,N_2629);
or U3384 (N_3384,N_2534,N_2845);
nand U3385 (N_3385,N_2696,N_2848);
nand U3386 (N_3386,N_2727,N_2738);
nand U3387 (N_3387,N_2854,N_2956);
nor U3388 (N_3388,N_2784,N_2606);
and U3389 (N_3389,N_2722,N_2946);
and U3390 (N_3390,N_2614,N_2759);
and U3391 (N_3391,N_2945,N_2783);
nand U3392 (N_3392,N_2931,N_2875);
nor U3393 (N_3393,N_2629,N_2929);
and U3394 (N_3394,N_2800,N_2589);
xnor U3395 (N_3395,N_2992,N_2575);
nand U3396 (N_3396,N_2626,N_2763);
or U3397 (N_3397,N_2527,N_2513);
nand U3398 (N_3398,N_2911,N_2991);
nand U3399 (N_3399,N_2697,N_2620);
or U3400 (N_3400,N_2595,N_2746);
or U3401 (N_3401,N_2834,N_2587);
nand U3402 (N_3402,N_2765,N_2917);
nor U3403 (N_3403,N_2783,N_2510);
and U3404 (N_3404,N_2692,N_2923);
and U3405 (N_3405,N_2965,N_2615);
and U3406 (N_3406,N_2724,N_2846);
and U3407 (N_3407,N_2811,N_2824);
and U3408 (N_3408,N_2509,N_2750);
xor U3409 (N_3409,N_2652,N_2545);
and U3410 (N_3410,N_2648,N_2525);
nand U3411 (N_3411,N_2844,N_2787);
nor U3412 (N_3412,N_2668,N_2583);
nand U3413 (N_3413,N_2528,N_2639);
or U3414 (N_3414,N_2918,N_2525);
nand U3415 (N_3415,N_2538,N_2841);
nand U3416 (N_3416,N_2573,N_2698);
or U3417 (N_3417,N_2693,N_2775);
nand U3418 (N_3418,N_2675,N_2682);
nand U3419 (N_3419,N_2671,N_2631);
nand U3420 (N_3420,N_2910,N_2527);
nand U3421 (N_3421,N_2543,N_2771);
nand U3422 (N_3422,N_2578,N_2795);
or U3423 (N_3423,N_2588,N_2584);
nand U3424 (N_3424,N_2621,N_2665);
nor U3425 (N_3425,N_2654,N_2915);
or U3426 (N_3426,N_2532,N_2791);
xnor U3427 (N_3427,N_2836,N_2881);
or U3428 (N_3428,N_2733,N_2715);
nor U3429 (N_3429,N_2739,N_2695);
and U3430 (N_3430,N_2694,N_2792);
nor U3431 (N_3431,N_2928,N_2505);
and U3432 (N_3432,N_2934,N_2674);
nand U3433 (N_3433,N_2818,N_2562);
or U3434 (N_3434,N_2949,N_2605);
or U3435 (N_3435,N_2580,N_2553);
or U3436 (N_3436,N_2553,N_2526);
or U3437 (N_3437,N_2846,N_2867);
or U3438 (N_3438,N_2532,N_2790);
nor U3439 (N_3439,N_2560,N_2951);
nand U3440 (N_3440,N_2681,N_2679);
and U3441 (N_3441,N_2984,N_2695);
or U3442 (N_3442,N_2957,N_2657);
or U3443 (N_3443,N_2827,N_2684);
or U3444 (N_3444,N_2555,N_2608);
and U3445 (N_3445,N_2836,N_2926);
nand U3446 (N_3446,N_2769,N_2557);
or U3447 (N_3447,N_2998,N_2911);
nand U3448 (N_3448,N_2886,N_2691);
nor U3449 (N_3449,N_2621,N_2749);
nand U3450 (N_3450,N_2741,N_2854);
and U3451 (N_3451,N_2975,N_2894);
and U3452 (N_3452,N_2922,N_2770);
nor U3453 (N_3453,N_2808,N_2745);
nor U3454 (N_3454,N_2593,N_2566);
or U3455 (N_3455,N_2785,N_2533);
nand U3456 (N_3456,N_2721,N_2994);
nor U3457 (N_3457,N_2784,N_2568);
nand U3458 (N_3458,N_2552,N_2753);
nor U3459 (N_3459,N_2874,N_2757);
and U3460 (N_3460,N_2935,N_2725);
nand U3461 (N_3461,N_2867,N_2992);
or U3462 (N_3462,N_2876,N_2984);
nand U3463 (N_3463,N_2888,N_2636);
or U3464 (N_3464,N_2575,N_2892);
or U3465 (N_3465,N_2855,N_2795);
and U3466 (N_3466,N_2893,N_2505);
nand U3467 (N_3467,N_2781,N_2981);
nor U3468 (N_3468,N_2957,N_2903);
and U3469 (N_3469,N_2889,N_2585);
nor U3470 (N_3470,N_2932,N_2842);
or U3471 (N_3471,N_2811,N_2888);
and U3472 (N_3472,N_2562,N_2556);
and U3473 (N_3473,N_2879,N_2565);
and U3474 (N_3474,N_2914,N_2694);
nand U3475 (N_3475,N_2813,N_2956);
nand U3476 (N_3476,N_2959,N_2784);
and U3477 (N_3477,N_2661,N_2546);
nand U3478 (N_3478,N_2536,N_2866);
and U3479 (N_3479,N_2754,N_2529);
and U3480 (N_3480,N_2639,N_2736);
nand U3481 (N_3481,N_2953,N_2780);
nand U3482 (N_3482,N_2886,N_2827);
nor U3483 (N_3483,N_2704,N_2739);
and U3484 (N_3484,N_2894,N_2807);
nand U3485 (N_3485,N_2605,N_2698);
and U3486 (N_3486,N_2846,N_2859);
or U3487 (N_3487,N_2628,N_2580);
nand U3488 (N_3488,N_2658,N_2689);
nand U3489 (N_3489,N_2506,N_2904);
or U3490 (N_3490,N_2684,N_2952);
nor U3491 (N_3491,N_2992,N_2623);
nor U3492 (N_3492,N_2625,N_2528);
and U3493 (N_3493,N_2584,N_2698);
xor U3494 (N_3494,N_2650,N_2640);
and U3495 (N_3495,N_2923,N_2549);
or U3496 (N_3496,N_2729,N_2837);
nand U3497 (N_3497,N_2628,N_2781);
or U3498 (N_3498,N_2621,N_2744);
and U3499 (N_3499,N_2737,N_2725);
or U3500 (N_3500,N_3165,N_3210);
or U3501 (N_3501,N_3006,N_3254);
xnor U3502 (N_3502,N_3004,N_3031);
nor U3503 (N_3503,N_3183,N_3396);
and U3504 (N_3504,N_3371,N_3121);
nand U3505 (N_3505,N_3336,N_3224);
and U3506 (N_3506,N_3058,N_3249);
nand U3507 (N_3507,N_3172,N_3242);
or U3508 (N_3508,N_3496,N_3442);
and U3509 (N_3509,N_3331,N_3042);
nand U3510 (N_3510,N_3047,N_3448);
and U3511 (N_3511,N_3081,N_3474);
nand U3512 (N_3512,N_3404,N_3184);
nand U3513 (N_3513,N_3060,N_3278);
or U3514 (N_3514,N_3204,N_3239);
nor U3515 (N_3515,N_3392,N_3306);
or U3516 (N_3516,N_3037,N_3284);
nor U3517 (N_3517,N_3388,N_3300);
nand U3518 (N_3518,N_3492,N_3260);
nor U3519 (N_3519,N_3401,N_3114);
nand U3520 (N_3520,N_3145,N_3299);
or U3521 (N_3521,N_3132,N_3194);
nor U3522 (N_3522,N_3261,N_3480);
nor U3523 (N_3523,N_3197,N_3068);
and U3524 (N_3524,N_3432,N_3196);
nor U3525 (N_3525,N_3310,N_3164);
and U3526 (N_3526,N_3235,N_3153);
or U3527 (N_3527,N_3471,N_3486);
or U3528 (N_3528,N_3203,N_3276);
nor U3529 (N_3529,N_3352,N_3103);
xnor U3530 (N_3530,N_3315,N_3245);
nor U3531 (N_3531,N_3199,N_3307);
nor U3532 (N_3532,N_3086,N_3266);
or U3533 (N_3533,N_3303,N_3246);
or U3534 (N_3534,N_3441,N_3127);
nand U3535 (N_3535,N_3369,N_3157);
and U3536 (N_3536,N_3177,N_3309);
and U3537 (N_3537,N_3113,N_3061);
and U3538 (N_3538,N_3329,N_3370);
nor U3539 (N_3539,N_3105,N_3272);
nor U3540 (N_3540,N_3250,N_3312);
nand U3541 (N_3541,N_3039,N_3146);
nand U3542 (N_3542,N_3470,N_3407);
and U3543 (N_3543,N_3419,N_3138);
and U3544 (N_3544,N_3048,N_3390);
nor U3545 (N_3545,N_3195,N_3283);
nand U3546 (N_3546,N_3410,N_3359);
and U3547 (N_3547,N_3134,N_3355);
nor U3548 (N_3548,N_3200,N_3149);
nor U3549 (N_3549,N_3099,N_3161);
or U3550 (N_3550,N_3228,N_3137);
and U3551 (N_3551,N_3072,N_3301);
nor U3552 (N_3552,N_3043,N_3167);
nand U3553 (N_3553,N_3464,N_3232);
or U3554 (N_3554,N_3259,N_3148);
or U3555 (N_3555,N_3302,N_3001);
and U3556 (N_3556,N_3033,N_3364);
or U3557 (N_3557,N_3133,N_3330);
nor U3558 (N_3558,N_3215,N_3084);
and U3559 (N_3559,N_3322,N_3425);
or U3560 (N_3560,N_3490,N_3156);
nor U3561 (N_3561,N_3460,N_3285);
and U3562 (N_3562,N_3350,N_3237);
nor U3563 (N_3563,N_3489,N_3078);
and U3564 (N_3564,N_3187,N_3125);
and U3565 (N_3565,N_3162,N_3345);
and U3566 (N_3566,N_3214,N_3181);
nor U3567 (N_3567,N_3076,N_3354);
nand U3568 (N_3568,N_3434,N_3383);
nor U3569 (N_3569,N_3003,N_3339);
and U3570 (N_3570,N_3136,N_3440);
and U3571 (N_3571,N_3130,N_3038);
nor U3572 (N_3572,N_3473,N_3495);
or U3573 (N_3573,N_3362,N_3100);
nor U3574 (N_3574,N_3155,N_3377);
or U3575 (N_3575,N_3318,N_3051);
or U3576 (N_3576,N_3258,N_3211);
nor U3577 (N_3577,N_3064,N_3154);
and U3578 (N_3578,N_3485,N_3201);
or U3579 (N_3579,N_3433,N_3091);
or U3580 (N_3580,N_3202,N_3144);
nand U3581 (N_3581,N_3163,N_3281);
or U3582 (N_3582,N_3212,N_3421);
nor U3583 (N_3583,N_3188,N_3159);
nand U3584 (N_3584,N_3080,N_3169);
nor U3585 (N_3585,N_3192,N_3208);
xor U3586 (N_3586,N_3279,N_3358);
or U3587 (N_3587,N_3381,N_3207);
and U3588 (N_3588,N_3223,N_3296);
xor U3589 (N_3589,N_3252,N_3436);
and U3590 (N_3590,N_3349,N_3314);
and U3591 (N_3591,N_3240,N_3447);
and U3592 (N_3592,N_3221,N_3170);
or U3593 (N_3593,N_3041,N_3244);
nor U3594 (N_3594,N_3123,N_3124);
nand U3595 (N_3595,N_3182,N_3117);
nor U3596 (N_3596,N_3411,N_3400);
or U3597 (N_3597,N_3241,N_3055);
or U3598 (N_3598,N_3226,N_3189);
nand U3599 (N_3599,N_3217,N_3115);
nor U3600 (N_3600,N_3360,N_3096);
nand U3601 (N_3601,N_3319,N_3010);
xnor U3602 (N_3602,N_3040,N_3206);
nand U3603 (N_3603,N_3173,N_3367);
and U3604 (N_3604,N_3045,N_3393);
nor U3605 (N_3605,N_3427,N_3268);
nor U3606 (N_3606,N_3479,N_3482);
nand U3607 (N_3607,N_3093,N_3015);
nand U3608 (N_3608,N_3443,N_3158);
nor U3609 (N_3609,N_3294,N_3332);
nand U3610 (N_3610,N_3234,N_3147);
and U3611 (N_3611,N_3365,N_3229);
nor U3612 (N_3612,N_3009,N_3498);
or U3613 (N_3613,N_3243,N_3389);
or U3614 (N_3614,N_3449,N_3374);
and U3615 (N_3615,N_3414,N_3190);
nand U3616 (N_3616,N_3253,N_3112);
nor U3617 (N_3617,N_3325,N_3139);
and U3618 (N_3618,N_3487,N_3417);
or U3619 (N_3619,N_3067,N_3057);
and U3620 (N_3620,N_3311,N_3408);
or U3621 (N_3621,N_3263,N_3437);
and U3622 (N_3622,N_3152,N_3363);
or U3623 (N_3623,N_3021,N_3267);
or U3624 (N_3624,N_3368,N_3185);
nand U3625 (N_3625,N_3002,N_3450);
nand U3626 (N_3626,N_3451,N_3444);
and U3627 (N_3627,N_3028,N_3459);
or U3628 (N_3628,N_3036,N_3225);
nand U3629 (N_3629,N_3431,N_3012);
nand U3630 (N_3630,N_3366,N_3070);
or U3631 (N_3631,N_3483,N_3412);
or U3632 (N_3632,N_3373,N_3213);
nand U3633 (N_3633,N_3405,N_3085);
or U3634 (N_3634,N_3461,N_3439);
and U3635 (N_3635,N_3446,N_3288);
and U3636 (N_3636,N_3334,N_3230);
nand U3637 (N_3637,N_3357,N_3394);
nor U3638 (N_3638,N_3397,N_3101);
and U3639 (N_3639,N_3455,N_3000);
or U3640 (N_3640,N_3475,N_3337);
nor U3641 (N_3641,N_3292,N_3198);
or U3642 (N_3642,N_3052,N_3293);
and U3643 (N_3643,N_3494,N_3476);
and U3644 (N_3644,N_3484,N_3026);
or U3645 (N_3645,N_3290,N_3341);
or U3646 (N_3646,N_3472,N_3077);
and U3647 (N_3647,N_3297,N_3463);
and U3648 (N_3648,N_3110,N_3168);
nor U3649 (N_3649,N_3372,N_3375);
or U3650 (N_3650,N_3035,N_3320);
nand U3651 (N_3651,N_3273,N_3378);
xnor U3652 (N_3652,N_3324,N_3104);
nor U3653 (N_3653,N_3030,N_3017);
or U3654 (N_3654,N_3347,N_3291);
nor U3655 (N_3655,N_3346,N_3097);
nand U3656 (N_3656,N_3270,N_3452);
and U3657 (N_3657,N_3430,N_3326);
or U3658 (N_3658,N_3335,N_3088);
nand U3659 (N_3659,N_3106,N_3094);
nand U3660 (N_3660,N_3298,N_3071);
nand U3661 (N_3661,N_3219,N_3118);
nor U3662 (N_3662,N_3090,N_3174);
and U3663 (N_3663,N_3044,N_3049);
nand U3664 (N_3664,N_3415,N_3348);
or U3665 (N_3665,N_3423,N_3435);
nand U3666 (N_3666,N_3286,N_3287);
and U3667 (N_3667,N_3481,N_3422);
nand U3668 (N_3668,N_3166,N_3054);
nand U3669 (N_3669,N_3493,N_3108);
nand U3670 (N_3670,N_3499,N_3102);
and U3671 (N_3671,N_3274,N_3176);
nand U3672 (N_3672,N_3251,N_3128);
or U3673 (N_3673,N_3141,N_3340);
or U3674 (N_3674,N_3257,N_3059);
or U3675 (N_3675,N_3126,N_3066);
or U3676 (N_3676,N_3327,N_3063);
or U3677 (N_3677,N_3295,N_3328);
or U3678 (N_3678,N_3022,N_3020);
xor U3679 (N_3679,N_3338,N_3416);
nor U3680 (N_3680,N_3018,N_3008);
and U3681 (N_3681,N_3248,N_3247);
nor U3682 (N_3682,N_3316,N_3160);
or U3683 (N_3683,N_3264,N_3227);
and U3684 (N_3684,N_3395,N_3007);
nand U3685 (N_3685,N_3380,N_3438);
nor U3686 (N_3686,N_3409,N_3062);
nor U3687 (N_3687,N_3466,N_3075);
and U3688 (N_3688,N_3069,N_3098);
and U3689 (N_3689,N_3180,N_3356);
or U3690 (N_3690,N_3005,N_3135);
nor U3691 (N_3691,N_3317,N_3304);
nand U3692 (N_3692,N_3218,N_3426);
and U3693 (N_3693,N_3428,N_3175);
and U3694 (N_3694,N_3032,N_3398);
or U3695 (N_3695,N_3216,N_3420);
nand U3696 (N_3696,N_3457,N_3024);
nor U3697 (N_3697,N_3351,N_3379);
nand U3698 (N_3698,N_3083,N_3477);
or U3699 (N_3699,N_3491,N_3343);
or U3700 (N_3700,N_3387,N_3089);
nor U3701 (N_3701,N_3107,N_3150);
and U3702 (N_3702,N_3353,N_3313);
nand U3703 (N_3703,N_3478,N_3403);
and U3704 (N_3704,N_3342,N_3282);
nor U3705 (N_3705,N_3386,N_3344);
and U3706 (N_3706,N_3073,N_3361);
nor U3707 (N_3707,N_3178,N_3385);
nor U3708 (N_3708,N_3019,N_3011);
or U3709 (N_3709,N_3468,N_3333);
or U3710 (N_3710,N_3462,N_3458);
nor U3711 (N_3711,N_3467,N_3142);
or U3712 (N_3712,N_3143,N_3454);
nor U3713 (N_3713,N_3469,N_3238);
or U3714 (N_3714,N_3056,N_3120);
or U3715 (N_3715,N_3013,N_3384);
or U3716 (N_3716,N_3465,N_3140);
or U3717 (N_3717,N_3236,N_3193);
nand U3718 (N_3718,N_3382,N_3376);
or U3719 (N_3719,N_3087,N_3456);
or U3720 (N_3720,N_3053,N_3233);
xor U3721 (N_3721,N_3095,N_3453);
and U3722 (N_3722,N_3014,N_3029);
nand U3723 (N_3723,N_3222,N_3429);
nand U3724 (N_3724,N_3116,N_3151);
and U3725 (N_3725,N_3323,N_3256);
nand U3726 (N_3726,N_3079,N_3488);
or U3727 (N_3727,N_3065,N_3231);
and U3728 (N_3728,N_3122,N_3092);
nor U3729 (N_3729,N_3497,N_3082);
xnor U3730 (N_3730,N_3275,N_3179);
nand U3731 (N_3731,N_3119,N_3445);
or U3732 (N_3732,N_3321,N_3271);
and U3733 (N_3733,N_3027,N_3025);
nor U3734 (N_3734,N_3129,N_3023);
nor U3735 (N_3735,N_3399,N_3205);
or U3736 (N_3736,N_3413,N_3305);
nor U3737 (N_3737,N_3289,N_3191);
or U3738 (N_3738,N_3406,N_3131);
nand U3739 (N_3739,N_3418,N_3424);
nor U3740 (N_3740,N_3402,N_3050);
nand U3741 (N_3741,N_3308,N_3074);
or U3742 (N_3742,N_3034,N_3046);
nand U3743 (N_3743,N_3209,N_3109);
nor U3744 (N_3744,N_3220,N_3016);
and U3745 (N_3745,N_3280,N_3269);
or U3746 (N_3746,N_3186,N_3277);
nand U3747 (N_3747,N_3171,N_3111);
and U3748 (N_3748,N_3262,N_3255);
and U3749 (N_3749,N_3265,N_3391);
nand U3750 (N_3750,N_3030,N_3485);
nand U3751 (N_3751,N_3064,N_3494);
and U3752 (N_3752,N_3241,N_3180);
xnor U3753 (N_3753,N_3013,N_3132);
or U3754 (N_3754,N_3179,N_3486);
nand U3755 (N_3755,N_3082,N_3211);
or U3756 (N_3756,N_3356,N_3060);
nor U3757 (N_3757,N_3015,N_3019);
nor U3758 (N_3758,N_3316,N_3011);
nor U3759 (N_3759,N_3208,N_3454);
and U3760 (N_3760,N_3163,N_3076);
nand U3761 (N_3761,N_3328,N_3464);
nand U3762 (N_3762,N_3131,N_3297);
or U3763 (N_3763,N_3141,N_3128);
nor U3764 (N_3764,N_3328,N_3389);
nor U3765 (N_3765,N_3373,N_3044);
nand U3766 (N_3766,N_3486,N_3367);
nor U3767 (N_3767,N_3283,N_3021);
nand U3768 (N_3768,N_3225,N_3478);
nor U3769 (N_3769,N_3325,N_3216);
or U3770 (N_3770,N_3020,N_3265);
nand U3771 (N_3771,N_3078,N_3024);
nand U3772 (N_3772,N_3332,N_3060);
and U3773 (N_3773,N_3112,N_3306);
xnor U3774 (N_3774,N_3064,N_3365);
nand U3775 (N_3775,N_3049,N_3422);
or U3776 (N_3776,N_3248,N_3171);
or U3777 (N_3777,N_3307,N_3466);
nand U3778 (N_3778,N_3146,N_3451);
nor U3779 (N_3779,N_3332,N_3397);
and U3780 (N_3780,N_3110,N_3288);
nand U3781 (N_3781,N_3485,N_3000);
or U3782 (N_3782,N_3051,N_3169);
nand U3783 (N_3783,N_3418,N_3471);
or U3784 (N_3784,N_3056,N_3027);
or U3785 (N_3785,N_3337,N_3241);
nand U3786 (N_3786,N_3253,N_3308);
xor U3787 (N_3787,N_3465,N_3468);
xor U3788 (N_3788,N_3163,N_3373);
nand U3789 (N_3789,N_3459,N_3313);
nand U3790 (N_3790,N_3422,N_3088);
nor U3791 (N_3791,N_3433,N_3407);
nand U3792 (N_3792,N_3306,N_3397);
nand U3793 (N_3793,N_3102,N_3167);
nor U3794 (N_3794,N_3099,N_3357);
nand U3795 (N_3795,N_3260,N_3247);
or U3796 (N_3796,N_3362,N_3296);
or U3797 (N_3797,N_3059,N_3250);
or U3798 (N_3798,N_3264,N_3234);
or U3799 (N_3799,N_3407,N_3468);
nor U3800 (N_3800,N_3453,N_3202);
nor U3801 (N_3801,N_3237,N_3337);
and U3802 (N_3802,N_3440,N_3157);
or U3803 (N_3803,N_3291,N_3005);
nand U3804 (N_3804,N_3008,N_3341);
xnor U3805 (N_3805,N_3448,N_3465);
or U3806 (N_3806,N_3055,N_3217);
nand U3807 (N_3807,N_3226,N_3094);
or U3808 (N_3808,N_3274,N_3297);
and U3809 (N_3809,N_3418,N_3168);
nor U3810 (N_3810,N_3204,N_3323);
or U3811 (N_3811,N_3291,N_3268);
nand U3812 (N_3812,N_3186,N_3014);
nor U3813 (N_3813,N_3219,N_3047);
nand U3814 (N_3814,N_3447,N_3465);
or U3815 (N_3815,N_3377,N_3355);
nand U3816 (N_3816,N_3339,N_3268);
nor U3817 (N_3817,N_3466,N_3394);
nand U3818 (N_3818,N_3097,N_3108);
and U3819 (N_3819,N_3474,N_3298);
nor U3820 (N_3820,N_3181,N_3422);
and U3821 (N_3821,N_3077,N_3373);
and U3822 (N_3822,N_3003,N_3490);
nor U3823 (N_3823,N_3246,N_3428);
or U3824 (N_3824,N_3441,N_3237);
and U3825 (N_3825,N_3189,N_3153);
nand U3826 (N_3826,N_3251,N_3297);
and U3827 (N_3827,N_3023,N_3025);
nand U3828 (N_3828,N_3061,N_3109);
or U3829 (N_3829,N_3030,N_3057);
nand U3830 (N_3830,N_3307,N_3253);
and U3831 (N_3831,N_3457,N_3191);
nor U3832 (N_3832,N_3318,N_3086);
and U3833 (N_3833,N_3010,N_3047);
nor U3834 (N_3834,N_3325,N_3003);
and U3835 (N_3835,N_3075,N_3378);
nand U3836 (N_3836,N_3080,N_3149);
or U3837 (N_3837,N_3141,N_3205);
or U3838 (N_3838,N_3370,N_3156);
nor U3839 (N_3839,N_3203,N_3292);
nand U3840 (N_3840,N_3046,N_3425);
or U3841 (N_3841,N_3394,N_3483);
xnor U3842 (N_3842,N_3480,N_3281);
nand U3843 (N_3843,N_3165,N_3413);
or U3844 (N_3844,N_3215,N_3320);
nand U3845 (N_3845,N_3078,N_3109);
or U3846 (N_3846,N_3489,N_3142);
nor U3847 (N_3847,N_3324,N_3185);
and U3848 (N_3848,N_3253,N_3389);
and U3849 (N_3849,N_3193,N_3334);
and U3850 (N_3850,N_3452,N_3297);
nor U3851 (N_3851,N_3313,N_3087);
and U3852 (N_3852,N_3246,N_3213);
nor U3853 (N_3853,N_3099,N_3176);
nor U3854 (N_3854,N_3045,N_3487);
or U3855 (N_3855,N_3401,N_3452);
and U3856 (N_3856,N_3485,N_3466);
nor U3857 (N_3857,N_3061,N_3358);
nor U3858 (N_3858,N_3419,N_3202);
or U3859 (N_3859,N_3281,N_3290);
nor U3860 (N_3860,N_3307,N_3076);
nor U3861 (N_3861,N_3422,N_3186);
nand U3862 (N_3862,N_3450,N_3142);
nand U3863 (N_3863,N_3442,N_3470);
nor U3864 (N_3864,N_3311,N_3095);
nor U3865 (N_3865,N_3016,N_3177);
or U3866 (N_3866,N_3438,N_3221);
and U3867 (N_3867,N_3133,N_3115);
or U3868 (N_3868,N_3192,N_3498);
nand U3869 (N_3869,N_3141,N_3101);
nor U3870 (N_3870,N_3104,N_3166);
nor U3871 (N_3871,N_3492,N_3483);
or U3872 (N_3872,N_3278,N_3307);
nand U3873 (N_3873,N_3103,N_3108);
nor U3874 (N_3874,N_3040,N_3447);
or U3875 (N_3875,N_3277,N_3012);
nor U3876 (N_3876,N_3421,N_3087);
nor U3877 (N_3877,N_3353,N_3475);
nor U3878 (N_3878,N_3067,N_3004);
nand U3879 (N_3879,N_3077,N_3047);
nor U3880 (N_3880,N_3087,N_3150);
or U3881 (N_3881,N_3298,N_3462);
nor U3882 (N_3882,N_3311,N_3113);
and U3883 (N_3883,N_3401,N_3469);
or U3884 (N_3884,N_3059,N_3393);
or U3885 (N_3885,N_3457,N_3035);
nor U3886 (N_3886,N_3141,N_3494);
nor U3887 (N_3887,N_3386,N_3083);
nor U3888 (N_3888,N_3288,N_3264);
and U3889 (N_3889,N_3285,N_3153);
nand U3890 (N_3890,N_3375,N_3333);
and U3891 (N_3891,N_3175,N_3228);
nand U3892 (N_3892,N_3360,N_3148);
and U3893 (N_3893,N_3267,N_3198);
or U3894 (N_3894,N_3135,N_3308);
or U3895 (N_3895,N_3217,N_3341);
or U3896 (N_3896,N_3452,N_3409);
and U3897 (N_3897,N_3471,N_3152);
or U3898 (N_3898,N_3020,N_3276);
or U3899 (N_3899,N_3318,N_3026);
and U3900 (N_3900,N_3143,N_3323);
nand U3901 (N_3901,N_3234,N_3246);
nand U3902 (N_3902,N_3327,N_3070);
and U3903 (N_3903,N_3107,N_3141);
or U3904 (N_3904,N_3440,N_3474);
nor U3905 (N_3905,N_3053,N_3066);
and U3906 (N_3906,N_3374,N_3168);
and U3907 (N_3907,N_3362,N_3263);
nor U3908 (N_3908,N_3243,N_3316);
nor U3909 (N_3909,N_3057,N_3408);
nor U3910 (N_3910,N_3177,N_3035);
or U3911 (N_3911,N_3265,N_3485);
nand U3912 (N_3912,N_3150,N_3303);
nor U3913 (N_3913,N_3259,N_3470);
and U3914 (N_3914,N_3332,N_3165);
or U3915 (N_3915,N_3154,N_3499);
or U3916 (N_3916,N_3132,N_3120);
nand U3917 (N_3917,N_3451,N_3116);
nor U3918 (N_3918,N_3229,N_3364);
or U3919 (N_3919,N_3273,N_3156);
or U3920 (N_3920,N_3063,N_3287);
and U3921 (N_3921,N_3181,N_3434);
and U3922 (N_3922,N_3385,N_3309);
and U3923 (N_3923,N_3046,N_3413);
nor U3924 (N_3924,N_3355,N_3372);
nand U3925 (N_3925,N_3054,N_3371);
or U3926 (N_3926,N_3165,N_3491);
nor U3927 (N_3927,N_3051,N_3212);
nand U3928 (N_3928,N_3054,N_3051);
nand U3929 (N_3929,N_3323,N_3008);
nor U3930 (N_3930,N_3177,N_3440);
nor U3931 (N_3931,N_3221,N_3167);
nor U3932 (N_3932,N_3434,N_3011);
nand U3933 (N_3933,N_3418,N_3333);
nor U3934 (N_3934,N_3472,N_3163);
and U3935 (N_3935,N_3421,N_3052);
and U3936 (N_3936,N_3071,N_3325);
and U3937 (N_3937,N_3202,N_3459);
nor U3938 (N_3938,N_3283,N_3086);
or U3939 (N_3939,N_3096,N_3312);
nand U3940 (N_3940,N_3028,N_3066);
nor U3941 (N_3941,N_3439,N_3039);
and U3942 (N_3942,N_3448,N_3438);
and U3943 (N_3943,N_3320,N_3221);
and U3944 (N_3944,N_3172,N_3093);
or U3945 (N_3945,N_3422,N_3005);
and U3946 (N_3946,N_3068,N_3437);
nor U3947 (N_3947,N_3231,N_3096);
or U3948 (N_3948,N_3275,N_3116);
or U3949 (N_3949,N_3283,N_3141);
and U3950 (N_3950,N_3385,N_3122);
nand U3951 (N_3951,N_3464,N_3203);
or U3952 (N_3952,N_3135,N_3023);
and U3953 (N_3953,N_3268,N_3054);
or U3954 (N_3954,N_3143,N_3188);
nand U3955 (N_3955,N_3255,N_3412);
and U3956 (N_3956,N_3367,N_3189);
nor U3957 (N_3957,N_3085,N_3256);
or U3958 (N_3958,N_3321,N_3294);
or U3959 (N_3959,N_3287,N_3289);
and U3960 (N_3960,N_3054,N_3382);
and U3961 (N_3961,N_3383,N_3218);
nand U3962 (N_3962,N_3430,N_3145);
nor U3963 (N_3963,N_3390,N_3345);
nor U3964 (N_3964,N_3428,N_3412);
nor U3965 (N_3965,N_3396,N_3317);
and U3966 (N_3966,N_3472,N_3397);
and U3967 (N_3967,N_3031,N_3268);
or U3968 (N_3968,N_3327,N_3207);
or U3969 (N_3969,N_3288,N_3439);
and U3970 (N_3970,N_3427,N_3060);
or U3971 (N_3971,N_3291,N_3176);
nor U3972 (N_3972,N_3484,N_3125);
or U3973 (N_3973,N_3377,N_3363);
and U3974 (N_3974,N_3080,N_3229);
nand U3975 (N_3975,N_3120,N_3498);
nor U3976 (N_3976,N_3336,N_3114);
nand U3977 (N_3977,N_3009,N_3082);
and U3978 (N_3978,N_3361,N_3150);
and U3979 (N_3979,N_3414,N_3494);
nor U3980 (N_3980,N_3126,N_3327);
and U3981 (N_3981,N_3346,N_3396);
or U3982 (N_3982,N_3178,N_3372);
nor U3983 (N_3983,N_3074,N_3361);
and U3984 (N_3984,N_3406,N_3265);
xnor U3985 (N_3985,N_3371,N_3033);
or U3986 (N_3986,N_3486,N_3085);
and U3987 (N_3987,N_3104,N_3051);
nand U3988 (N_3988,N_3092,N_3321);
nor U3989 (N_3989,N_3380,N_3349);
or U3990 (N_3990,N_3095,N_3186);
nor U3991 (N_3991,N_3024,N_3386);
nor U3992 (N_3992,N_3235,N_3243);
and U3993 (N_3993,N_3301,N_3111);
or U3994 (N_3994,N_3238,N_3320);
and U3995 (N_3995,N_3394,N_3166);
or U3996 (N_3996,N_3110,N_3076);
and U3997 (N_3997,N_3223,N_3134);
and U3998 (N_3998,N_3072,N_3455);
nor U3999 (N_3999,N_3157,N_3271);
or U4000 (N_4000,N_3859,N_3986);
nand U4001 (N_4001,N_3695,N_3806);
and U4002 (N_4002,N_3895,N_3908);
and U4003 (N_4003,N_3547,N_3590);
nor U4004 (N_4004,N_3995,N_3709);
and U4005 (N_4005,N_3528,N_3651);
nor U4006 (N_4006,N_3565,N_3734);
nor U4007 (N_4007,N_3624,N_3999);
nand U4008 (N_4008,N_3967,N_3613);
and U4009 (N_4009,N_3523,N_3943);
or U4010 (N_4010,N_3681,N_3520);
nand U4011 (N_4011,N_3915,N_3625);
and U4012 (N_4012,N_3641,N_3955);
and U4013 (N_4013,N_3716,N_3822);
nor U4014 (N_4014,N_3530,N_3906);
or U4015 (N_4015,N_3803,N_3937);
or U4016 (N_4016,N_3932,N_3934);
or U4017 (N_4017,N_3997,N_3699);
nor U4018 (N_4018,N_3634,N_3790);
or U4019 (N_4019,N_3629,N_3774);
nor U4020 (N_4020,N_3797,N_3794);
or U4021 (N_4021,N_3686,N_3584);
nand U4022 (N_4022,N_3534,N_3777);
nand U4023 (N_4023,N_3996,N_3899);
and U4024 (N_4024,N_3741,N_3637);
or U4025 (N_4025,N_3704,N_3931);
or U4026 (N_4026,N_3974,N_3628);
or U4027 (N_4027,N_3820,N_3635);
nor U4028 (N_4028,N_3987,N_3732);
and U4029 (N_4029,N_3792,N_3655);
or U4030 (N_4030,N_3607,N_3860);
or U4031 (N_4031,N_3764,N_3516);
nand U4032 (N_4032,N_3731,N_3983);
or U4033 (N_4033,N_3621,N_3865);
nand U4034 (N_4034,N_3879,N_3562);
nand U4035 (N_4035,N_3990,N_3918);
or U4036 (N_4036,N_3919,N_3608);
and U4037 (N_4037,N_3927,N_3905);
and U4038 (N_4038,N_3500,N_3828);
or U4039 (N_4039,N_3855,N_3761);
nor U4040 (N_4040,N_3598,N_3599);
nor U4041 (N_4041,N_3907,N_3580);
and U4042 (N_4042,N_3617,N_3872);
or U4043 (N_4043,N_3532,N_3657);
or U4044 (N_4044,N_3810,N_3666);
nor U4045 (N_4045,N_3816,N_3964);
nand U4046 (N_4046,N_3750,N_3929);
nand U4047 (N_4047,N_3623,N_3642);
nand U4048 (N_4048,N_3900,N_3733);
or U4049 (N_4049,N_3705,N_3745);
nand U4050 (N_4050,N_3809,N_3756);
nor U4051 (N_4051,N_3744,N_3805);
or U4052 (N_4052,N_3798,N_3939);
and U4053 (N_4053,N_3891,N_3989);
or U4054 (N_4054,N_3721,N_3722);
and U4055 (N_4055,N_3930,N_3869);
or U4056 (N_4056,N_3982,N_3706);
and U4057 (N_4057,N_3845,N_3739);
nand U4058 (N_4058,N_3549,N_3852);
or U4059 (N_4059,N_3904,N_3848);
nor U4060 (N_4060,N_3522,N_3885);
and U4061 (N_4061,N_3842,N_3773);
and U4062 (N_4062,N_3707,N_3896);
and U4063 (N_4063,N_3515,N_3619);
nand U4064 (N_4064,N_3688,N_3597);
nor U4065 (N_4065,N_3938,N_3550);
nand U4066 (N_4066,N_3693,N_3600);
or U4067 (N_4067,N_3609,N_3627);
or U4068 (N_4068,N_3646,N_3540);
and U4069 (N_4069,N_3743,N_3768);
or U4070 (N_4070,N_3780,N_3779);
nand U4071 (N_4071,N_3763,N_3799);
and U4072 (N_4072,N_3873,N_3933);
or U4073 (N_4073,N_3740,N_3949);
or U4074 (N_4074,N_3793,N_3714);
and U4075 (N_4075,N_3563,N_3587);
nand U4076 (N_4076,N_3749,N_3804);
or U4077 (N_4077,N_3633,N_3573);
and U4078 (N_4078,N_3735,N_3593);
nor U4079 (N_4079,N_3993,N_3509);
and U4080 (N_4080,N_3874,N_3850);
or U4081 (N_4081,N_3977,N_3559);
nand U4082 (N_4082,N_3877,N_3753);
nor U4083 (N_4083,N_3514,N_3660);
and U4084 (N_4084,N_3862,N_3730);
or U4085 (N_4085,N_3647,N_3579);
nor U4086 (N_4086,N_3663,N_3759);
nor U4087 (N_4087,N_3962,N_3680);
or U4088 (N_4088,N_3829,N_3638);
nand U4089 (N_4089,N_3728,N_3992);
or U4090 (N_4090,N_3737,N_3970);
nor U4091 (N_4091,N_3594,N_3557);
nor U4092 (N_4092,N_3770,N_3687);
or U4093 (N_4093,N_3678,N_3653);
nand U4094 (N_4094,N_3917,N_3662);
or U4095 (N_4095,N_3781,N_3576);
nand U4096 (N_4096,N_3566,N_3656);
or U4097 (N_4097,N_3504,N_3630);
nor U4098 (N_4098,N_3672,N_3815);
nor U4099 (N_4099,N_3751,N_3881);
nand U4100 (N_4100,N_3808,N_3920);
and U4101 (N_4101,N_3615,N_3802);
nand U4102 (N_4102,N_3925,N_3851);
and U4103 (N_4103,N_3769,N_3512);
nor U4104 (N_4104,N_3531,N_3736);
nor U4105 (N_4105,N_3517,N_3632);
nor U4106 (N_4106,N_3618,N_3545);
nor U4107 (N_4107,N_3758,N_3585);
xor U4108 (N_4108,N_3571,N_3592);
nand U4109 (N_4109,N_3752,N_3772);
nor U4110 (N_4110,N_3928,N_3871);
or U4111 (N_4111,N_3813,N_3601);
nor U4112 (N_4112,N_3844,N_3708);
and U4113 (N_4113,N_3849,N_3510);
and U4114 (N_4114,N_3775,N_3575);
or U4115 (N_4115,N_3981,N_3711);
or U4116 (N_4116,N_3503,N_3880);
nand U4117 (N_4117,N_3991,N_3692);
nor U4118 (N_4118,N_3947,N_3664);
nor U4119 (N_4119,N_3537,N_3720);
and U4120 (N_4120,N_3696,N_3935);
or U4121 (N_4121,N_3833,N_3760);
and U4122 (N_4122,N_3723,N_3957);
or U4123 (N_4123,N_3645,N_3742);
nor U4124 (N_4124,N_3644,N_3971);
nor U4125 (N_4125,N_3538,N_3541);
nor U4126 (N_4126,N_3507,N_3972);
nor U4127 (N_4127,N_3924,N_3511);
and U4128 (N_4128,N_3786,N_3560);
nand U4129 (N_4129,N_3755,N_3643);
nand U4130 (N_4130,N_3694,N_3572);
xor U4131 (N_4131,N_3551,N_3564);
and U4132 (N_4132,N_3668,N_3856);
and U4133 (N_4133,N_3715,N_3703);
or U4134 (N_4134,N_3941,N_3506);
nand U4135 (N_4135,N_3554,N_3868);
nor U4136 (N_4136,N_3948,N_3836);
nand U4137 (N_4137,N_3544,N_3535);
nor U4138 (N_4138,N_3639,N_3909);
or U4139 (N_4139,N_3876,N_3835);
and U4140 (N_4140,N_3807,N_3866);
nor U4141 (N_4141,N_3719,N_3748);
or U4142 (N_4142,N_3826,N_3603);
nor U4143 (N_4143,N_3689,N_3713);
nor U4144 (N_4144,N_3819,N_3683);
nor U4145 (N_4145,N_3785,N_3976);
nor U4146 (N_4146,N_3953,N_3998);
and U4147 (N_4147,N_3596,N_3757);
nor U4148 (N_4148,N_3979,N_3595);
or U4149 (N_4149,N_3838,N_3832);
or U4150 (N_4150,N_3961,N_3913);
or U4151 (N_4151,N_3978,N_3926);
nand U4152 (N_4152,N_3670,N_3887);
and U4153 (N_4153,N_3529,N_3831);
or U4154 (N_4154,N_3543,N_3582);
or U4155 (N_4155,N_3667,N_3984);
nand U4156 (N_4156,N_3502,N_3602);
or U4157 (N_4157,N_3843,N_3898);
and U4158 (N_4158,N_3911,N_3766);
nand U4159 (N_4159,N_3654,N_3966);
and U4160 (N_4160,N_3508,N_3616);
and U4161 (N_4161,N_3944,N_3675);
nand U4162 (N_4162,N_3631,N_3903);
nor U4163 (N_4163,N_3589,N_3669);
xnor U4164 (N_4164,N_3969,N_3622);
and U4165 (N_4165,N_3568,N_3526);
or U4166 (N_4166,N_3676,N_3893);
nand U4167 (N_4167,N_3762,N_3837);
or U4168 (N_4168,N_3519,N_3727);
and U4169 (N_4169,N_3548,N_3821);
nand U4170 (N_4170,N_3536,N_3942);
nand U4171 (N_4171,N_3671,N_3814);
and U4172 (N_4172,N_3956,N_3890);
and U4173 (N_4173,N_3784,N_3945);
nand U4174 (N_4174,N_3700,N_3620);
nand U4175 (N_4175,N_3800,N_3677);
nor U4176 (N_4176,N_3542,N_3888);
nand U4177 (N_4177,N_3847,N_3724);
nor U4178 (N_4178,N_3747,N_3787);
and U4179 (N_4179,N_3701,N_3527);
nand U4180 (N_4180,N_3827,N_3994);
or U4181 (N_4181,N_3946,N_3611);
and U4182 (N_4182,N_3556,N_3988);
and U4183 (N_4183,N_3746,N_3658);
and U4184 (N_4184,N_3636,N_3682);
xnor U4185 (N_4185,N_3950,N_3659);
nand U4186 (N_4186,N_3717,N_3738);
nand U4187 (N_4187,N_3697,N_3782);
nand U4188 (N_4188,N_3652,N_3965);
or U4189 (N_4189,N_3846,N_3916);
and U4190 (N_4190,N_3910,N_3936);
or U4191 (N_4191,N_3754,N_3606);
nor U4192 (N_4192,N_3570,N_3854);
nor U4193 (N_4193,N_3959,N_3980);
or U4194 (N_4194,N_3922,N_3830);
nand U4195 (N_4195,N_3975,N_3569);
and U4196 (N_4196,N_3783,N_3857);
or U4197 (N_4197,N_3649,N_3778);
nand U4198 (N_4198,N_3889,N_3875);
xnor U4199 (N_4199,N_3533,N_3912);
nor U4200 (N_4200,N_3921,N_3870);
or U4201 (N_4201,N_3588,N_3546);
or U4202 (N_4202,N_3679,N_3840);
nand U4203 (N_4203,N_3818,N_3897);
or U4204 (N_4204,N_3789,N_3673);
nand U4205 (N_4205,N_3698,N_3525);
nor U4206 (N_4206,N_3882,N_3811);
nand U4207 (N_4207,N_3610,N_3513);
or U4208 (N_4208,N_3886,N_3726);
nor U4209 (N_4209,N_3552,N_3864);
nor U4210 (N_4210,N_3812,N_3940);
and U4211 (N_4211,N_3902,N_3914);
nor U4212 (N_4212,N_3674,N_3841);
nand U4213 (N_4213,N_3973,N_3958);
and U4214 (N_4214,N_3577,N_3858);
nor U4215 (N_4215,N_3801,N_3834);
nand U4216 (N_4216,N_3796,N_3853);
xnor U4217 (N_4217,N_3521,N_3963);
nand U4218 (N_4218,N_3867,N_3586);
or U4219 (N_4219,N_3518,N_3581);
and U4220 (N_4220,N_3901,N_3578);
or U4221 (N_4221,N_3884,N_3952);
nor U4222 (N_4222,N_3791,N_3684);
nor U4223 (N_4223,N_3825,N_3640);
and U4224 (N_4224,N_3883,N_3685);
or U4225 (N_4225,N_3718,N_3817);
nand U4226 (N_4226,N_3823,N_3725);
or U4227 (N_4227,N_3954,N_3960);
and U4228 (N_4228,N_3863,N_3691);
and U4229 (N_4229,N_3771,N_3648);
or U4230 (N_4230,N_3878,N_3729);
nor U4231 (N_4231,N_3985,N_3539);
or U4232 (N_4232,N_3839,N_3558);
xor U4233 (N_4233,N_3861,N_3501);
nand U4234 (N_4234,N_3788,N_3591);
nand U4235 (N_4235,N_3583,N_3892);
nand U4236 (N_4236,N_3795,N_3951);
or U4237 (N_4237,N_3555,N_3553);
nand U4238 (N_4238,N_3712,N_3604);
xnor U4239 (N_4239,N_3650,N_3612);
nor U4240 (N_4240,N_3894,N_3776);
or U4241 (N_4241,N_3614,N_3567);
or U4242 (N_4242,N_3665,N_3690);
nor U4243 (N_4243,N_3605,N_3767);
xor U4244 (N_4244,N_3574,N_3661);
or U4245 (N_4245,N_3968,N_3524);
or U4246 (N_4246,N_3923,N_3710);
and U4247 (N_4247,N_3702,N_3505);
or U4248 (N_4248,N_3765,N_3824);
and U4249 (N_4249,N_3626,N_3561);
nand U4250 (N_4250,N_3563,N_3952);
or U4251 (N_4251,N_3973,N_3893);
nand U4252 (N_4252,N_3559,N_3953);
nand U4253 (N_4253,N_3943,N_3886);
or U4254 (N_4254,N_3745,N_3701);
or U4255 (N_4255,N_3595,N_3546);
nor U4256 (N_4256,N_3616,N_3695);
nand U4257 (N_4257,N_3501,N_3644);
or U4258 (N_4258,N_3826,N_3507);
nand U4259 (N_4259,N_3893,N_3745);
nand U4260 (N_4260,N_3852,N_3674);
and U4261 (N_4261,N_3864,N_3827);
or U4262 (N_4262,N_3626,N_3805);
nor U4263 (N_4263,N_3820,N_3778);
and U4264 (N_4264,N_3555,N_3573);
nor U4265 (N_4265,N_3599,N_3708);
nor U4266 (N_4266,N_3954,N_3777);
nor U4267 (N_4267,N_3580,N_3824);
or U4268 (N_4268,N_3611,N_3731);
and U4269 (N_4269,N_3695,N_3733);
nand U4270 (N_4270,N_3758,N_3899);
and U4271 (N_4271,N_3923,N_3912);
nor U4272 (N_4272,N_3852,N_3524);
and U4273 (N_4273,N_3504,N_3529);
nor U4274 (N_4274,N_3890,N_3751);
and U4275 (N_4275,N_3517,N_3722);
and U4276 (N_4276,N_3629,N_3634);
nor U4277 (N_4277,N_3503,N_3789);
nor U4278 (N_4278,N_3958,N_3653);
and U4279 (N_4279,N_3668,N_3891);
nand U4280 (N_4280,N_3863,N_3909);
and U4281 (N_4281,N_3963,N_3726);
nor U4282 (N_4282,N_3676,N_3749);
xor U4283 (N_4283,N_3909,N_3739);
or U4284 (N_4284,N_3722,N_3789);
nor U4285 (N_4285,N_3730,N_3875);
nand U4286 (N_4286,N_3587,N_3901);
and U4287 (N_4287,N_3976,N_3579);
and U4288 (N_4288,N_3994,N_3817);
and U4289 (N_4289,N_3969,N_3702);
or U4290 (N_4290,N_3681,N_3887);
or U4291 (N_4291,N_3666,N_3587);
nand U4292 (N_4292,N_3721,N_3845);
and U4293 (N_4293,N_3840,N_3978);
and U4294 (N_4294,N_3710,N_3993);
nor U4295 (N_4295,N_3860,N_3618);
nand U4296 (N_4296,N_3834,N_3635);
nor U4297 (N_4297,N_3927,N_3851);
and U4298 (N_4298,N_3777,N_3871);
or U4299 (N_4299,N_3705,N_3971);
and U4300 (N_4300,N_3623,N_3504);
nand U4301 (N_4301,N_3945,N_3586);
and U4302 (N_4302,N_3689,N_3611);
nor U4303 (N_4303,N_3801,N_3833);
nand U4304 (N_4304,N_3662,N_3673);
nor U4305 (N_4305,N_3568,N_3896);
or U4306 (N_4306,N_3924,N_3642);
nand U4307 (N_4307,N_3697,N_3948);
nor U4308 (N_4308,N_3674,N_3940);
and U4309 (N_4309,N_3829,N_3866);
nand U4310 (N_4310,N_3707,N_3901);
nand U4311 (N_4311,N_3968,N_3595);
nor U4312 (N_4312,N_3513,N_3681);
nor U4313 (N_4313,N_3794,N_3867);
nor U4314 (N_4314,N_3741,N_3920);
and U4315 (N_4315,N_3785,N_3903);
and U4316 (N_4316,N_3608,N_3582);
or U4317 (N_4317,N_3594,N_3664);
or U4318 (N_4318,N_3768,N_3574);
and U4319 (N_4319,N_3653,N_3526);
and U4320 (N_4320,N_3707,N_3542);
or U4321 (N_4321,N_3768,N_3971);
or U4322 (N_4322,N_3586,N_3907);
nor U4323 (N_4323,N_3803,N_3928);
nand U4324 (N_4324,N_3958,N_3873);
nor U4325 (N_4325,N_3941,N_3885);
nand U4326 (N_4326,N_3889,N_3846);
nor U4327 (N_4327,N_3667,N_3854);
nand U4328 (N_4328,N_3518,N_3702);
nor U4329 (N_4329,N_3843,N_3951);
nand U4330 (N_4330,N_3731,N_3714);
nand U4331 (N_4331,N_3692,N_3643);
or U4332 (N_4332,N_3595,N_3640);
and U4333 (N_4333,N_3638,N_3870);
and U4334 (N_4334,N_3507,N_3596);
nand U4335 (N_4335,N_3733,N_3559);
nand U4336 (N_4336,N_3738,N_3903);
and U4337 (N_4337,N_3877,N_3774);
nor U4338 (N_4338,N_3771,N_3727);
nand U4339 (N_4339,N_3546,N_3885);
and U4340 (N_4340,N_3564,N_3891);
nor U4341 (N_4341,N_3935,N_3800);
and U4342 (N_4342,N_3900,N_3963);
nand U4343 (N_4343,N_3945,N_3846);
nor U4344 (N_4344,N_3782,N_3732);
and U4345 (N_4345,N_3548,N_3954);
or U4346 (N_4346,N_3708,N_3794);
nor U4347 (N_4347,N_3899,N_3616);
or U4348 (N_4348,N_3811,N_3533);
or U4349 (N_4349,N_3788,N_3983);
nor U4350 (N_4350,N_3733,N_3723);
nand U4351 (N_4351,N_3547,N_3596);
or U4352 (N_4352,N_3907,N_3834);
or U4353 (N_4353,N_3593,N_3847);
or U4354 (N_4354,N_3750,N_3891);
nand U4355 (N_4355,N_3898,N_3713);
or U4356 (N_4356,N_3874,N_3737);
nor U4357 (N_4357,N_3570,N_3522);
and U4358 (N_4358,N_3812,N_3572);
or U4359 (N_4359,N_3547,N_3611);
nand U4360 (N_4360,N_3655,N_3824);
nand U4361 (N_4361,N_3998,N_3917);
and U4362 (N_4362,N_3687,N_3598);
nand U4363 (N_4363,N_3806,N_3761);
nand U4364 (N_4364,N_3797,N_3859);
nand U4365 (N_4365,N_3562,N_3862);
nor U4366 (N_4366,N_3983,N_3759);
nand U4367 (N_4367,N_3903,N_3792);
or U4368 (N_4368,N_3614,N_3578);
and U4369 (N_4369,N_3961,N_3986);
nor U4370 (N_4370,N_3999,N_3679);
or U4371 (N_4371,N_3659,N_3930);
nand U4372 (N_4372,N_3816,N_3609);
or U4373 (N_4373,N_3544,N_3509);
xnor U4374 (N_4374,N_3861,N_3661);
nand U4375 (N_4375,N_3565,N_3841);
nand U4376 (N_4376,N_3636,N_3999);
and U4377 (N_4377,N_3780,N_3859);
nand U4378 (N_4378,N_3529,N_3798);
or U4379 (N_4379,N_3714,N_3586);
or U4380 (N_4380,N_3620,N_3798);
or U4381 (N_4381,N_3910,N_3854);
nand U4382 (N_4382,N_3591,N_3645);
nor U4383 (N_4383,N_3510,N_3500);
and U4384 (N_4384,N_3878,N_3510);
or U4385 (N_4385,N_3699,N_3662);
nand U4386 (N_4386,N_3685,N_3543);
and U4387 (N_4387,N_3746,N_3895);
and U4388 (N_4388,N_3822,N_3768);
nor U4389 (N_4389,N_3582,N_3900);
nand U4390 (N_4390,N_3957,N_3702);
nor U4391 (N_4391,N_3712,N_3732);
or U4392 (N_4392,N_3541,N_3913);
nand U4393 (N_4393,N_3723,N_3931);
or U4394 (N_4394,N_3624,N_3955);
nor U4395 (N_4395,N_3590,N_3672);
or U4396 (N_4396,N_3963,N_3885);
or U4397 (N_4397,N_3943,N_3852);
and U4398 (N_4398,N_3687,N_3582);
and U4399 (N_4399,N_3729,N_3578);
nor U4400 (N_4400,N_3711,N_3725);
nor U4401 (N_4401,N_3699,N_3660);
nand U4402 (N_4402,N_3965,N_3641);
nand U4403 (N_4403,N_3817,N_3950);
and U4404 (N_4404,N_3877,N_3645);
or U4405 (N_4405,N_3597,N_3881);
and U4406 (N_4406,N_3698,N_3844);
nor U4407 (N_4407,N_3995,N_3682);
or U4408 (N_4408,N_3997,N_3673);
or U4409 (N_4409,N_3564,N_3734);
nand U4410 (N_4410,N_3593,N_3586);
and U4411 (N_4411,N_3586,N_3798);
or U4412 (N_4412,N_3512,N_3926);
nand U4413 (N_4413,N_3955,N_3899);
nand U4414 (N_4414,N_3911,N_3618);
and U4415 (N_4415,N_3794,N_3691);
nor U4416 (N_4416,N_3534,N_3662);
or U4417 (N_4417,N_3785,N_3939);
and U4418 (N_4418,N_3748,N_3812);
or U4419 (N_4419,N_3763,N_3812);
nand U4420 (N_4420,N_3879,N_3605);
and U4421 (N_4421,N_3789,N_3617);
nor U4422 (N_4422,N_3694,N_3631);
or U4423 (N_4423,N_3940,N_3973);
nor U4424 (N_4424,N_3777,N_3576);
and U4425 (N_4425,N_3989,N_3529);
or U4426 (N_4426,N_3560,N_3687);
and U4427 (N_4427,N_3532,N_3704);
nor U4428 (N_4428,N_3757,N_3570);
or U4429 (N_4429,N_3807,N_3805);
nor U4430 (N_4430,N_3567,N_3710);
nand U4431 (N_4431,N_3628,N_3540);
nand U4432 (N_4432,N_3587,N_3990);
nand U4433 (N_4433,N_3946,N_3635);
nor U4434 (N_4434,N_3583,N_3971);
nand U4435 (N_4435,N_3500,N_3697);
or U4436 (N_4436,N_3539,N_3699);
nor U4437 (N_4437,N_3560,N_3718);
nand U4438 (N_4438,N_3851,N_3576);
and U4439 (N_4439,N_3759,N_3571);
nor U4440 (N_4440,N_3858,N_3788);
nand U4441 (N_4441,N_3859,N_3729);
and U4442 (N_4442,N_3683,N_3996);
or U4443 (N_4443,N_3613,N_3785);
xnor U4444 (N_4444,N_3818,N_3970);
and U4445 (N_4445,N_3731,N_3567);
xor U4446 (N_4446,N_3874,N_3849);
nor U4447 (N_4447,N_3526,N_3766);
and U4448 (N_4448,N_3689,N_3995);
or U4449 (N_4449,N_3918,N_3524);
and U4450 (N_4450,N_3940,N_3907);
or U4451 (N_4451,N_3883,N_3815);
and U4452 (N_4452,N_3786,N_3815);
or U4453 (N_4453,N_3861,N_3930);
nand U4454 (N_4454,N_3763,N_3923);
nor U4455 (N_4455,N_3878,N_3578);
nor U4456 (N_4456,N_3757,N_3953);
nor U4457 (N_4457,N_3972,N_3848);
nand U4458 (N_4458,N_3951,N_3936);
and U4459 (N_4459,N_3694,N_3651);
and U4460 (N_4460,N_3784,N_3694);
and U4461 (N_4461,N_3897,N_3537);
or U4462 (N_4462,N_3534,N_3788);
and U4463 (N_4463,N_3683,N_3709);
and U4464 (N_4464,N_3833,N_3776);
nor U4465 (N_4465,N_3817,N_3617);
or U4466 (N_4466,N_3876,N_3895);
and U4467 (N_4467,N_3743,N_3536);
and U4468 (N_4468,N_3659,N_3799);
or U4469 (N_4469,N_3723,N_3548);
and U4470 (N_4470,N_3866,N_3716);
nor U4471 (N_4471,N_3700,N_3634);
nor U4472 (N_4472,N_3802,N_3604);
nor U4473 (N_4473,N_3793,N_3556);
and U4474 (N_4474,N_3942,N_3648);
and U4475 (N_4475,N_3887,N_3734);
and U4476 (N_4476,N_3587,N_3798);
nor U4477 (N_4477,N_3936,N_3794);
and U4478 (N_4478,N_3763,N_3855);
or U4479 (N_4479,N_3579,N_3997);
or U4480 (N_4480,N_3925,N_3813);
or U4481 (N_4481,N_3558,N_3764);
nor U4482 (N_4482,N_3704,N_3766);
or U4483 (N_4483,N_3592,N_3738);
and U4484 (N_4484,N_3811,N_3888);
or U4485 (N_4485,N_3858,N_3551);
nand U4486 (N_4486,N_3501,N_3726);
nand U4487 (N_4487,N_3846,N_3894);
nor U4488 (N_4488,N_3997,N_3935);
nand U4489 (N_4489,N_3548,N_3775);
or U4490 (N_4490,N_3540,N_3672);
or U4491 (N_4491,N_3692,N_3624);
nor U4492 (N_4492,N_3620,N_3949);
and U4493 (N_4493,N_3739,N_3589);
and U4494 (N_4494,N_3881,N_3582);
nor U4495 (N_4495,N_3765,N_3602);
and U4496 (N_4496,N_3831,N_3766);
or U4497 (N_4497,N_3839,N_3659);
nand U4498 (N_4498,N_3566,N_3955);
nor U4499 (N_4499,N_3517,N_3504);
nor U4500 (N_4500,N_4167,N_4156);
and U4501 (N_4501,N_4077,N_4349);
nor U4502 (N_4502,N_4197,N_4394);
nor U4503 (N_4503,N_4292,N_4054);
and U4504 (N_4504,N_4201,N_4298);
nand U4505 (N_4505,N_4411,N_4308);
or U4506 (N_4506,N_4441,N_4109);
and U4507 (N_4507,N_4249,N_4198);
nand U4508 (N_4508,N_4439,N_4188);
or U4509 (N_4509,N_4141,N_4379);
and U4510 (N_4510,N_4242,N_4426);
nor U4511 (N_4511,N_4325,N_4177);
or U4512 (N_4512,N_4289,N_4313);
nor U4513 (N_4513,N_4029,N_4192);
or U4514 (N_4514,N_4027,N_4282);
nand U4515 (N_4515,N_4280,N_4068);
nor U4516 (N_4516,N_4438,N_4337);
or U4517 (N_4517,N_4346,N_4272);
nand U4518 (N_4518,N_4161,N_4030);
nor U4519 (N_4519,N_4266,N_4022);
or U4520 (N_4520,N_4045,N_4130);
and U4521 (N_4521,N_4191,N_4464);
and U4522 (N_4522,N_4255,N_4490);
and U4523 (N_4523,N_4224,N_4361);
and U4524 (N_4524,N_4305,N_4078);
nor U4525 (N_4525,N_4101,N_4344);
or U4526 (N_4526,N_4491,N_4055);
and U4527 (N_4527,N_4422,N_4137);
and U4528 (N_4528,N_4142,N_4367);
or U4529 (N_4529,N_4225,N_4442);
nor U4530 (N_4530,N_4237,N_4015);
nor U4531 (N_4531,N_4283,N_4395);
nor U4532 (N_4532,N_4258,N_4195);
or U4533 (N_4533,N_4063,N_4259);
nor U4534 (N_4534,N_4489,N_4475);
or U4535 (N_4535,N_4116,N_4342);
or U4536 (N_4536,N_4327,N_4217);
nand U4537 (N_4537,N_4113,N_4004);
or U4538 (N_4538,N_4302,N_4321);
or U4539 (N_4539,N_4414,N_4125);
nand U4540 (N_4540,N_4229,N_4157);
and U4541 (N_4541,N_4447,N_4200);
nand U4542 (N_4542,N_4139,N_4417);
nor U4543 (N_4543,N_4360,N_4136);
nand U4544 (N_4544,N_4383,N_4213);
and U4545 (N_4545,N_4042,N_4216);
or U4546 (N_4546,N_4455,N_4017);
and U4547 (N_4547,N_4482,N_4354);
nor U4548 (N_4548,N_4076,N_4187);
nor U4549 (N_4549,N_4485,N_4398);
and U4550 (N_4550,N_4276,N_4430);
nand U4551 (N_4551,N_4038,N_4037);
nor U4552 (N_4552,N_4173,N_4368);
and U4553 (N_4553,N_4215,N_4232);
nor U4554 (N_4554,N_4220,N_4124);
nand U4555 (N_4555,N_4051,N_4393);
or U4556 (N_4556,N_4285,N_4300);
and U4557 (N_4557,N_4218,N_4160);
nand U4558 (N_4558,N_4025,N_4243);
nor U4559 (N_4559,N_4102,N_4153);
or U4560 (N_4560,N_4370,N_4221);
nand U4561 (N_4561,N_4401,N_4081);
nor U4562 (N_4562,N_4031,N_4185);
or U4563 (N_4563,N_4330,N_4032);
nor U4564 (N_4564,N_4362,N_4089);
or U4565 (N_4565,N_4046,N_4159);
or U4566 (N_4566,N_4431,N_4115);
and U4567 (N_4567,N_4403,N_4207);
and U4568 (N_4568,N_4286,N_4408);
nor U4569 (N_4569,N_4412,N_4098);
nand U4570 (N_4570,N_4105,N_4110);
xor U4571 (N_4571,N_4180,N_4453);
nand U4572 (N_4572,N_4212,N_4470);
or U4573 (N_4573,N_4333,N_4168);
nand U4574 (N_4574,N_4070,N_4399);
nand U4575 (N_4575,N_4460,N_4497);
nor U4576 (N_4576,N_4021,N_4169);
or U4577 (N_4577,N_4114,N_4226);
or U4578 (N_4578,N_4176,N_4432);
nor U4579 (N_4579,N_4041,N_4165);
and U4580 (N_4580,N_4499,N_4445);
xnor U4581 (N_4581,N_4240,N_4372);
or U4582 (N_4582,N_4359,N_4118);
nor U4583 (N_4583,N_4483,N_4040);
nand U4584 (N_4584,N_4264,N_4448);
nor U4585 (N_4585,N_4026,N_4211);
nor U4586 (N_4586,N_4277,N_4146);
or U4587 (N_4587,N_4074,N_4481);
nand U4588 (N_4588,N_4091,N_4446);
nand U4589 (N_4589,N_4083,N_4099);
nand U4590 (N_4590,N_4376,N_4126);
and U4591 (N_4591,N_4248,N_4131);
nand U4592 (N_4592,N_4196,N_4143);
nor U4593 (N_4593,N_4246,N_4247);
and U4594 (N_4594,N_4477,N_4410);
nand U4595 (N_4595,N_4275,N_4092);
nor U4596 (N_4596,N_4100,N_4343);
nand U4597 (N_4597,N_4474,N_4381);
and U4598 (N_4598,N_4036,N_4375);
and U4599 (N_4599,N_4424,N_4230);
or U4600 (N_4600,N_4458,N_4340);
nand U4601 (N_4601,N_4095,N_4048);
nor U4602 (N_4602,N_4496,N_4402);
nand U4603 (N_4603,N_4338,N_4364);
and U4604 (N_4604,N_4009,N_4444);
nor U4605 (N_4605,N_4476,N_4005);
and U4606 (N_4606,N_4251,N_4443);
and U4607 (N_4607,N_4205,N_4303);
nor U4608 (N_4608,N_4479,N_4049);
and U4609 (N_4609,N_4382,N_4067);
or U4610 (N_4610,N_4179,N_4204);
and U4611 (N_4611,N_4210,N_4405);
or U4612 (N_4612,N_4064,N_4366);
nor U4613 (N_4613,N_4473,N_4466);
and U4614 (N_4614,N_4094,N_4365);
nand U4615 (N_4615,N_4181,N_4072);
nor U4616 (N_4616,N_4128,N_4059);
xnor U4617 (N_4617,N_4323,N_4409);
nand U4618 (N_4618,N_4271,N_4019);
or U4619 (N_4619,N_4384,N_4082);
nand U4620 (N_4620,N_4469,N_4011);
nand U4621 (N_4621,N_4468,N_4086);
or U4622 (N_4622,N_4075,N_4132);
nor U4623 (N_4623,N_4133,N_4208);
or U4624 (N_4624,N_4363,N_4149);
and U4625 (N_4625,N_4274,N_4163);
nor U4626 (N_4626,N_4016,N_4090);
or U4627 (N_4627,N_4106,N_4378);
nor U4628 (N_4628,N_4257,N_4087);
nor U4629 (N_4629,N_4209,N_4147);
or U4630 (N_4630,N_4241,N_4312);
nor U4631 (N_4631,N_4175,N_4206);
or U4632 (N_4632,N_4145,N_4413);
nor U4633 (N_4633,N_4415,N_4202);
and U4634 (N_4634,N_4425,N_4331);
nand U4635 (N_4635,N_4290,N_4385);
or U4636 (N_4636,N_4487,N_4315);
nand U4637 (N_4637,N_4096,N_4281);
or U4638 (N_4638,N_4267,N_4352);
nand U4639 (N_4639,N_4419,N_4449);
and U4640 (N_4640,N_4456,N_4339);
nand U4641 (N_4641,N_4158,N_4494);
or U4642 (N_4642,N_4459,N_4355);
nand U4643 (N_4643,N_4079,N_4214);
nor U4644 (N_4644,N_4461,N_4244);
and U4645 (N_4645,N_4463,N_4199);
or U4646 (N_4646,N_4073,N_4080);
nand U4647 (N_4647,N_4035,N_4127);
xor U4648 (N_4648,N_4471,N_4391);
or U4649 (N_4649,N_4278,N_4162);
nand U4650 (N_4650,N_4288,N_4033);
nor U4651 (N_4651,N_4052,N_4423);
nand U4652 (N_4652,N_4317,N_4034);
or U4653 (N_4653,N_4238,N_4390);
or U4654 (N_4654,N_4012,N_4299);
and U4655 (N_4655,N_4332,N_4150);
and U4656 (N_4656,N_4454,N_4043);
and U4657 (N_4657,N_4235,N_4002);
nand U4658 (N_4658,N_4231,N_4297);
and U4659 (N_4659,N_4223,N_4254);
nor U4660 (N_4660,N_4270,N_4164);
and U4661 (N_4661,N_4172,N_4301);
and U4662 (N_4662,N_4318,N_4097);
nand U4663 (N_4663,N_4154,N_4166);
or U4664 (N_4664,N_4252,N_4256);
or U4665 (N_4665,N_4138,N_4295);
nand U4666 (N_4666,N_4085,N_4347);
nand U4667 (N_4667,N_4400,N_4350);
nor U4668 (N_4668,N_4013,N_4062);
nor U4669 (N_4669,N_4152,N_4227);
nor U4670 (N_4670,N_4478,N_4486);
nor U4671 (N_4671,N_4324,N_4151);
nor U4672 (N_4672,N_4069,N_4000);
nand U4673 (N_4673,N_4122,N_4465);
nand U4674 (N_4674,N_4006,N_4261);
and U4675 (N_4675,N_4319,N_4358);
or U4676 (N_4676,N_4392,N_4388);
nor U4677 (N_4677,N_4234,N_4245);
nor U4678 (N_4678,N_4121,N_4291);
and U4679 (N_4679,N_4260,N_4320);
and U4680 (N_4680,N_4003,N_4129);
nand U4681 (N_4681,N_4493,N_4228);
and U4682 (N_4682,N_4386,N_4155);
or U4683 (N_4683,N_4189,N_4039);
nand U4684 (N_4684,N_4001,N_4287);
nand U4685 (N_4685,N_4488,N_4397);
nor U4686 (N_4686,N_4345,N_4296);
or U4687 (N_4687,N_4265,N_4023);
nor U4688 (N_4688,N_4307,N_4050);
or U4689 (N_4689,N_4007,N_4071);
nand U4690 (N_4690,N_4404,N_4348);
nand U4691 (N_4691,N_4111,N_4310);
and U4692 (N_4692,N_4322,N_4279);
and U4693 (N_4693,N_4269,N_4203);
and U4694 (N_4694,N_4356,N_4311);
nor U4695 (N_4695,N_4421,N_4429);
nor U4696 (N_4696,N_4066,N_4123);
and U4697 (N_4697,N_4434,N_4467);
or U4698 (N_4698,N_4057,N_4377);
and U4699 (N_4699,N_4184,N_4088);
nand U4700 (N_4700,N_4480,N_4452);
or U4701 (N_4701,N_4484,N_4058);
or U4702 (N_4702,N_4357,N_4472);
nor U4703 (N_4703,N_4250,N_4104);
nand U4704 (N_4704,N_4387,N_4406);
or U4705 (N_4705,N_4233,N_4428);
and U4706 (N_4706,N_4060,N_4140);
nand U4707 (N_4707,N_4047,N_4262);
and U4708 (N_4708,N_4273,N_4371);
nand U4709 (N_4709,N_4190,N_4144);
or U4710 (N_4710,N_4450,N_4020);
nor U4711 (N_4711,N_4263,N_4326);
nor U4712 (N_4712,N_4369,N_4028);
or U4713 (N_4713,N_4108,N_4457);
and U4714 (N_4714,N_4117,N_4380);
or U4715 (N_4715,N_4194,N_4440);
or U4716 (N_4716,N_4120,N_4024);
xor U4717 (N_4717,N_4341,N_4084);
or U4718 (N_4718,N_4353,N_4495);
nor U4719 (N_4719,N_4389,N_4433);
and U4720 (N_4720,N_4435,N_4407);
nand U4721 (N_4721,N_4134,N_4119);
and U4722 (N_4722,N_4293,N_4418);
and U4723 (N_4723,N_4492,N_4420);
or U4724 (N_4724,N_4416,N_4183);
nand U4725 (N_4725,N_4135,N_4284);
nor U4726 (N_4726,N_4328,N_4451);
or U4727 (N_4727,N_4112,N_4182);
or U4728 (N_4728,N_4239,N_4236);
or U4729 (N_4729,N_4268,N_4336);
or U4730 (N_4730,N_4193,N_4170);
nand U4731 (N_4731,N_4056,N_4314);
nand U4732 (N_4732,N_4396,N_4053);
nor U4733 (N_4733,N_4018,N_4103);
or U4734 (N_4734,N_4351,N_4010);
and U4735 (N_4735,N_4107,N_4436);
and U4736 (N_4736,N_4061,N_4373);
or U4737 (N_4737,N_4309,N_4178);
nor U4738 (N_4738,N_4253,N_4437);
and U4739 (N_4739,N_4093,N_4498);
and U4740 (N_4740,N_4008,N_4174);
xnor U4741 (N_4741,N_4306,N_4222);
nor U4742 (N_4742,N_4316,N_4329);
nor U4743 (N_4743,N_4374,N_4014);
and U4744 (N_4744,N_4171,N_4186);
and U4745 (N_4745,N_4294,N_4427);
and U4746 (N_4746,N_4462,N_4335);
xnor U4747 (N_4747,N_4334,N_4065);
and U4748 (N_4748,N_4148,N_4219);
nand U4749 (N_4749,N_4304,N_4044);
and U4750 (N_4750,N_4144,N_4196);
nand U4751 (N_4751,N_4003,N_4009);
nor U4752 (N_4752,N_4154,N_4031);
or U4753 (N_4753,N_4425,N_4359);
or U4754 (N_4754,N_4353,N_4284);
nand U4755 (N_4755,N_4250,N_4366);
nor U4756 (N_4756,N_4340,N_4186);
and U4757 (N_4757,N_4188,N_4045);
and U4758 (N_4758,N_4340,N_4264);
and U4759 (N_4759,N_4498,N_4239);
nor U4760 (N_4760,N_4194,N_4245);
nor U4761 (N_4761,N_4471,N_4007);
or U4762 (N_4762,N_4463,N_4440);
and U4763 (N_4763,N_4191,N_4325);
or U4764 (N_4764,N_4219,N_4126);
xor U4765 (N_4765,N_4151,N_4072);
and U4766 (N_4766,N_4081,N_4167);
nand U4767 (N_4767,N_4251,N_4456);
or U4768 (N_4768,N_4183,N_4280);
nor U4769 (N_4769,N_4475,N_4335);
nand U4770 (N_4770,N_4374,N_4489);
nand U4771 (N_4771,N_4185,N_4198);
nor U4772 (N_4772,N_4284,N_4066);
and U4773 (N_4773,N_4440,N_4185);
or U4774 (N_4774,N_4107,N_4359);
and U4775 (N_4775,N_4117,N_4074);
nor U4776 (N_4776,N_4260,N_4094);
nand U4777 (N_4777,N_4283,N_4316);
nor U4778 (N_4778,N_4266,N_4305);
or U4779 (N_4779,N_4462,N_4489);
nand U4780 (N_4780,N_4060,N_4314);
xnor U4781 (N_4781,N_4303,N_4364);
nor U4782 (N_4782,N_4472,N_4437);
nand U4783 (N_4783,N_4340,N_4494);
or U4784 (N_4784,N_4126,N_4413);
xnor U4785 (N_4785,N_4178,N_4155);
and U4786 (N_4786,N_4278,N_4021);
or U4787 (N_4787,N_4415,N_4408);
or U4788 (N_4788,N_4417,N_4205);
nand U4789 (N_4789,N_4318,N_4195);
nand U4790 (N_4790,N_4417,N_4160);
or U4791 (N_4791,N_4284,N_4283);
and U4792 (N_4792,N_4121,N_4162);
nor U4793 (N_4793,N_4018,N_4268);
nand U4794 (N_4794,N_4372,N_4016);
nor U4795 (N_4795,N_4038,N_4130);
nor U4796 (N_4796,N_4156,N_4454);
or U4797 (N_4797,N_4094,N_4339);
nand U4798 (N_4798,N_4474,N_4068);
nor U4799 (N_4799,N_4058,N_4001);
or U4800 (N_4800,N_4028,N_4150);
and U4801 (N_4801,N_4143,N_4395);
nor U4802 (N_4802,N_4431,N_4061);
nor U4803 (N_4803,N_4402,N_4483);
nand U4804 (N_4804,N_4065,N_4117);
nor U4805 (N_4805,N_4435,N_4071);
nand U4806 (N_4806,N_4064,N_4046);
nor U4807 (N_4807,N_4308,N_4208);
and U4808 (N_4808,N_4471,N_4380);
and U4809 (N_4809,N_4270,N_4294);
nor U4810 (N_4810,N_4117,N_4200);
nand U4811 (N_4811,N_4342,N_4049);
or U4812 (N_4812,N_4391,N_4287);
nor U4813 (N_4813,N_4197,N_4339);
nand U4814 (N_4814,N_4181,N_4310);
nand U4815 (N_4815,N_4308,N_4136);
or U4816 (N_4816,N_4217,N_4001);
nor U4817 (N_4817,N_4464,N_4332);
or U4818 (N_4818,N_4292,N_4203);
nor U4819 (N_4819,N_4063,N_4323);
nand U4820 (N_4820,N_4021,N_4235);
nand U4821 (N_4821,N_4449,N_4021);
nand U4822 (N_4822,N_4227,N_4466);
nor U4823 (N_4823,N_4137,N_4304);
and U4824 (N_4824,N_4301,N_4177);
and U4825 (N_4825,N_4169,N_4273);
nor U4826 (N_4826,N_4192,N_4296);
nor U4827 (N_4827,N_4297,N_4213);
or U4828 (N_4828,N_4268,N_4382);
nor U4829 (N_4829,N_4395,N_4396);
and U4830 (N_4830,N_4335,N_4451);
nor U4831 (N_4831,N_4389,N_4441);
nor U4832 (N_4832,N_4453,N_4301);
nand U4833 (N_4833,N_4214,N_4060);
and U4834 (N_4834,N_4488,N_4338);
or U4835 (N_4835,N_4045,N_4393);
and U4836 (N_4836,N_4085,N_4428);
nor U4837 (N_4837,N_4325,N_4389);
and U4838 (N_4838,N_4289,N_4441);
or U4839 (N_4839,N_4020,N_4211);
nand U4840 (N_4840,N_4186,N_4415);
or U4841 (N_4841,N_4038,N_4079);
or U4842 (N_4842,N_4141,N_4155);
nor U4843 (N_4843,N_4448,N_4411);
nor U4844 (N_4844,N_4268,N_4188);
and U4845 (N_4845,N_4322,N_4208);
nor U4846 (N_4846,N_4275,N_4376);
and U4847 (N_4847,N_4218,N_4352);
nor U4848 (N_4848,N_4132,N_4200);
and U4849 (N_4849,N_4433,N_4033);
or U4850 (N_4850,N_4034,N_4336);
xor U4851 (N_4851,N_4421,N_4171);
or U4852 (N_4852,N_4221,N_4289);
nor U4853 (N_4853,N_4192,N_4493);
or U4854 (N_4854,N_4343,N_4063);
nand U4855 (N_4855,N_4246,N_4459);
or U4856 (N_4856,N_4214,N_4091);
and U4857 (N_4857,N_4165,N_4002);
and U4858 (N_4858,N_4222,N_4330);
and U4859 (N_4859,N_4391,N_4094);
or U4860 (N_4860,N_4248,N_4276);
and U4861 (N_4861,N_4008,N_4164);
nand U4862 (N_4862,N_4010,N_4262);
and U4863 (N_4863,N_4207,N_4466);
nand U4864 (N_4864,N_4306,N_4264);
nand U4865 (N_4865,N_4361,N_4085);
nand U4866 (N_4866,N_4011,N_4117);
nor U4867 (N_4867,N_4370,N_4386);
and U4868 (N_4868,N_4013,N_4296);
or U4869 (N_4869,N_4176,N_4256);
or U4870 (N_4870,N_4097,N_4266);
nand U4871 (N_4871,N_4193,N_4414);
or U4872 (N_4872,N_4415,N_4401);
and U4873 (N_4873,N_4495,N_4008);
nand U4874 (N_4874,N_4203,N_4103);
nor U4875 (N_4875,N_4284,N_4461);
nor U4876 (N_4876,N_4055,N_4322);
or U4877 (N_4877,N_4432,N_4254);
and U4878 (N_4878,N_4485,N_4035);
nor U4879 (N_4879,N_4293,N_4408);
nand U4880 (N_4880,N_4357,N_4131);
or U4881 (N_4881,N_4231,N_4033);
or U4882 (N_4882,N_4304,N_4388);
nand U4883 (N_4883,N_4321,N_4421);
nand U4884 (N_4884,N_4016,N_4472);
and U4885 (N_4885,N_4497,N_4326);
and U4886 (N_4886,N_4485,N_4437);
or U4887 (N_4887,N_4189,N_4337);
nand U4888 (N_4888,N_4468,N_4023);
and U4889 (N_4889,N_4179,N_4184);
or U4890 (N_4890,N_4435,N_4417);
xnor U4891 (N_4891,N_4259,N_4203);
or U4892 (N_4892,N_4436,N_4214);
or U4893 (N_4893,N_4099,N_4293);
or U4894 (N_4894,N_4353,N_4472);
or U4895 (N_4895,N_4244,N_4095);
nand U4896 (N_4896,N_4284,N_4495);
or U4897 (N_4897,N_4375,N_4312);
nor U4898 (N_4898,N_4084,N_4165);
or U4899 (N_4899,N_4431,N_4222);
nor U4900 (N_4900,N_4377,N_4249);
nor U4901 (N_4901,N_4337,N_4236);
or U4902 (N_4902,N_4342,N_4005);
nor U4903 (N_4903,N_4022,N_4306);
nor U4904 (N_4904,N_4176,N_4429);
nand U4905 (N_4905,N_4380,N_4490);
nand U4906 (N_4906,N_4160,N_4328);
and U4907 (N_4907,N_4214,N_4076);
nor U4908 (N_4908,N_4469,N_4244);
and U4909 (N_4909,N_4119,N_4075);
nand U4910 (N_4910,N_4271,N_4232);
or U4911 (N_4911,N_4283,N_4263);
nor U4912 (N_4912,N_4474,N_4206);
and U4913 (N_4913,N_4184,N_4087);
and U4914 (N_4914,N_4230,N_4136);
or U4915 (N_4915,N_4241,N_4141);
and U4916 (N_4916,N_4440,N_4196);
nand U4917 (N_4917,N_4000,N_4090);
and U4918 (N_4918,N_4188,N_4198);
or U4919 (N_4919,N_4301,N_4140);
or U4920 (N_4920,N_4162,N_4181);
or U4921 (N_4921,N_4370,N_4396);
and U4922 (N_4922,N_4104,N_4074);
xnor U4923 (N_4923,N_4176,N_4318);
and U4924 (N_4924,N_4426,N_4117);
or U4925 (N_4925,N_4408,N_4024);
nand U4926 (N_4926,N_4409,N_4125);
nand U4927 (N_4927,N_4357,N_4046);
or U4928 (N_4928,N_4242,N_4140);
nor U4929 (N_4929,N_4205,N_4046);
and U4930 (N_4930,N_4485,N_4123);
nor U4931 (N_4931,N_4227,N_4061);
nand U4932 (N_4932,N_4343,N_4471);
or U4933 (N_4933,N_4446,N_4083);
or U4934 (N_4934,N_4083,N_4258);
or U4935 (N_4935,N_4107,N_4462);
or U4936 (N_4936,N_4383,N_4234);
nor U4937 (N_4937,N_4251,N_4496);
nand U4938 (N_4938,N_4488,N_4358);
or U4939 (N_4939,N_4457,N_4229);
or U4940 (N_4940,N_4256,N_4020);
and U4941 (N_4941,N_4219,N_4174);
nor U4942 (N_4942,N_4294,N_4460);
nor U4943 (N_4943,N_4361,N_4097);
nand U4944 (N_4944,N_4469,N_4391);
and U4945 (N_4945,N_4355,N_4410);
nor U4946 (N_4946,N_4105,N_4186);
nor U4947 (N_4947,N_4322,N_4242);
nand U4948 (N_4948,N_4162,N_4157);
nor U4949 (N_4949,N_4013,N_4226);
or U4950 (N_4950,N_4187,N_4036);
and U4951 (N_4951,N_4420,N_4228);
nor U4952 (N_4952,N_4488,N_4174);
nor U4953 (N_4953,N_4226,N_4186);
or U4954 (N_4954,N_4102,N_4408);
and U4955 (N_4955,N_4179,N_4051);
nand U4956 (N_4956,N_4430,N_4084);
or U4957 (N_4957,N_4203,N_4493);
and U4958 (N_4958,N_4472,N_4032);
xnor U4959 (N_4959,N_4251,N_4106);
nor U4960 (N_4960,N_4082,N_4372);
nor U4961 (N_4961,N_4123,N_4090);
nand U4962 (N_4962,N_4081,N_4363);
nor U4963 (N_4963,N_4480,N_4147);
and U4964 (N_4964,N_4220,N_4433);
nand U4965 (N_4965,N_4279,N_4102);
or U4966 (N_4966,N_4360,N_4377);
nor U4967 (N_4967,N_4129,N_4487);
and U4968 (N_4968,N_4473,N_4180);
or U4969 (N_4969,N_4217,N_4259);
and U4970 (N_4970,N_4081,N_4233);
nor U4971 (N_4971,N_4052,N_4096);
and U4972 (N_4972,N_4325,N_4137);
and U4973 (N_4973,N_4188,N_4304);
nand U4974 (N_4974,N_4419,N_4344);
nand U4975 (N_4975,N_4353,N_4055);
nand U4976 (N_4976,N_4443,N_4186);
and U4977 (N_4977,N_4440,N_4067);
nand U4978 (N_4978,N_4316,N_4317);
or U4979 (N_4979,N_4092,N_4427);
nor U4980 (N_4980,N_4227,N_4199);
nand U4981 (N_4981,N_4100,N_4017);
and U4982 (N_4982,N_4342,N_4186);
nand U4983 (N_4983,N_4498,N_4012);
and U4984 (N_4984,N_4020,N_4331);
nand U4985 (N_4985,N_4119,N_4174);
or U4986 (N_4986,N_4031,N_4363);
or U4987 (N_4987,N_4441,N_4118);
nand U4988 (N_4988,N_4085,N_4123);
or U4989 (N_4989,N_4472,N_4400);
and U4990 (N_4990,N_4012,N_4122);
or U4991 (N_4991,N_4391,N_4412);
nor U4992 (N_4992,N_4361,N_4359);
or U4993 (N_4993,N_4458,N_4464);
or U4994 (N_4994,N_4044,N_4032);
and U4995 (N_4995,N_4298,N_4438);
nor U4996 (N_4996,N_4064,N_4321);
or U4997 (N_4997,N_4148,N_4424);
or U4998 (N_4998,N_4279,N_4042);
nor U4999 (N_4999,N_4273,N_4391);
or U5000 (N_5000,N_4898,N_4727);
nand U5001 (N_5001,N_4575,N_4873);
nand U5002 (N_5002,N_4834,N_4584);
and U5003 (N_5003,N_4787,N_4555);
and U5004 (N_5004,N_4817,N_4528);
nor U5005 (N_5005,N_4815,N_4501);
nand U5006 (N_5006,N_4759,N_4965);
or U5007 (N_5007,N_4619,N_4832);
nor U5008 (N_5008,N_4559,N_4703);
and U5009 (N_5009,N_4944,N_4950);
nand U5010 (N_5010,N_4977,N_4953);
nor U5011 (N_5011,N_4734,N_4547);
nor U5012 (N_5012,N_4979,N_4598);
nor U5013 (N_5013,N_4949,N_4908);
nor U5014 (N_5014,N_4722,N_4512);
nand U5015 (N_5015,N_4629,N_4837);
or U5016 (N_5016,N_4566,N_4589);
or U5017 (N_5017,N_4620,N_4997);
nand U5018 (N_5018,N_4565,N_4931);
nand U5019 (N_5019,N_4884,N_4780);
nand U5020 (N_5020,N_4867,N_4503);
and U5021 (N_5021,N_4511,N_4593);
xnor U5022 (N_5022,N_4825,N_4536);
or U5023 (N_5023,N_4890,N_4641);
nand U5024 (N_5024,N_4693,N_4718);
or U5025 (N_5025,N_4752,N_4923);
nand U5026 (N_5026,N_4994,N_4645);
and U5027 (N_5027,N_4914,N_4828);
xnor U5028 (N_5028,N_4674,N_4863);
or U5029 (N_5029,N_4721,N_4982);
nand U5030 (N_5030,N_4657,N_4579);
nor U5031 (N_5031,N_4842,N_4713);
nor U5032 (N_5032,N_4646,N_4917);
and U5033 (N_5033,N_4580,N_4869);
nor U5034 (N_5034,N_4905,N_4519);
and U5035 (N_5035,N_4683,N_4918);
nand U5036 (N_5036,N_4983,N_4625);
or U5037 (N_5037,N_4790,N_4864);
nor U5038 (N_5038,N_4849,N_4880);
or U5039 (N_5039,N_4616,N_4577);
nor U5040 (N_5040,N_4609,N_4538);
and U5041 (N_5041,N_4690,N_4553);
and U5042 (N_5042,N_4604,N_4818);
and U5043 (N_5043,N_4866,N_4673);
nor U5044 (N_5044,N_4853,N_4699);
and U5045 (N_5045,N_4698,N_4529);
or U5046 (N_5046,N_4545,N_4899);
or U5047 (N_5047,N_4573,N_4719);
nor U5048 (N_5048,N_4938,N_4760);
nand U5049 (N_5049,N_4662,N_4981);
nor U5050 (N_5050,N_4875,N_4824);
nor U5051 (N_5051,N_4739,N_4618);
and U5052 (N_5052,N_4655,N_4877);
nand U5053 (N_5053,N_4562,N_4777);
and U5054 (N_5054,N_4996,N_4667);
nand U5055 (N_5055,N_4642,N_4986);
nand U5056 (N_5056,N_4906,N_4692);
nor U5057 (N_5057,N_4627,N_4883);
and U5058 (N_5058,N_4578,N_4596);
and U5059 (N_5059,N_4820,N_4804);
nor U5060 (N_5060,N_4518,N_4705);
and U5061 (N_5061,N_4821,N_4970);
or U5062 (N_5062,N_4819,N_4661);
or U5063 (N_5063,N_4791,N_4796);
nand U5064 (N_5064,N_4707,N_4812);
and U5065 (N_5065,N_4885,N_4505);
nor U5066 (N_5066,N_4521,N_4636);
or U5067 (N_5067,N_4751,N_4913);
xor U5068 (N_5068,N_4685,N_4639);
or U5069 (N_5069,N_4643,N_4992);
nand U5070 (N_5070,N_4606,N_4640);
nand U5071 (N_5071,N_4676,N_4856);
or U5072 (N_5072,N_4978,N_4850);
and U5073 (N_5073,N_4564,N_4909);
or U5074 (N_5074,N_4985,N_4717);
nand U5075 (N_5075,N_4581,N_4874);
or U5076 (N_5076,N_4767,N_4786);
nor U5077 (N_5077,N_4724,N_4915);
nor U5078 (N_5078,N_4628,N_4811);
nor U5079 (N_5079,N_4845,N_4907);
nand U5080 (N_5080,N_4858,N_4860);
or U5081 (N_5081,N_4813,N_4569);
nand U5082 (N_5082,N_4622,N_4653);
nand U5083 (N_5083,N_4847,N_4774);
nand U5084 (N_5084,N_4612,N_4762);
nand U5085 (N_5085,N_4998,N_4506);
nor U5086 (N_5086,N_4588,N_4967);
and U5087 (N_5087,N_4586,N_4988);
nor U5088 (N_5088,N_4689,N_4725);
or U5089 (N_5089,N_4525,N_4631);
nor U5090 (N_5090,N_4669,N_4556);
nor U5091 (N_5091,N_4697,N_4614);
or U5092 (N_5092,N_4870,N_4647);
nand U5093 (N_5093,N_4763,N_4814);
nor U5094 (N_5094,N_4781,N_4776);
or U5095 (N_5095,N_4865,N_4527);
and U5096 (N_5096,N_4783,N_4803);
nor U5097 (N_5097,N_4935,N_4753);
or U5098 (N_5098,N_4520,N_4857);
and U5099 (N_5099,N_4920,N_4746);
or U5100 (N_5100,N_4946,N_4543);
or U5101 (N_5101,N_4621,N_4792);
nor U5102 (N_5102,N_4966,N_4758);
or U5103 (N_5103,N_4859,N_4597);
nor U5104 (N_5104,N_4720,N_4749);
nand U5105 (N_5105,N_4663,N_4868);
nand U5106 (N_5106,N_4782,N_4648);
and U5107 (N_5107,N_4537,N_4638);
nor U5108 (N_5108,N_4954,N_4926);
nand U5109 (N_5109,N_4568,N_4633);
or U5110 (N_5110,N_4678,N_4700);
nand U5111 (N_5111,N_4708,N_4887);
nand U5112 (N_5112,N_4924,N_4879);
or U5113 (N_5113,N_4969,N_4583);
nand U5114 (N_5114,N_4740,N_4592);
or U5115 (N_5115,N_4761,N_4574);
nand U5116 (N_5116,N_4769,N_4947);
or U5117 (N_5117,N_4735,N_4927);
or U5118 (N_5118,N_4801,N_4770);
or U5119 (N_5119,N_4539,N_4710);
or U5120 (N_5120,N_4766,N_4823);
nand U5121 (N_5121,N_4535,N_4590);
nor U5122 (N_5122,N_4902,N_4534);
nand U5123 (N_5123,N_4549,N_4682);
nand U5124 (N_5124,N_4650,N_4962);
or U5125 (N_5125,N_4807,N_4838);
nor U5126 (N_5126,N_4896,N_4541);
or U5127 (N_5127,N_4798,N_4613);
and U5128 (N_5128,N_4702,N_4611);
nand U5129 (N_5129,N_4911,N_4548);
or U5130 (N_5130,N_4932,N_4972);
or U5131 (N_5131,N_4560,N_4973);
and U5132 (N_5132,N_4893,N_4844);
nor U5133 (N_5133,N_4773,N_4572);
or U5134 (N_5134,N_4610,N_4958);
or U5135 (N_5135,N_4743,N_4542);
nor U5136 (N_5136,N_4943,N_4582);
nor U5137 (N_5137,N_4848,N_4554);
nor U5138 (N_5138,N_4839,N_4933);
and U5139 (N_5139,N_4530,N_4993);
and U5140 (N_5140,N_4892,N_4715);
or U5141 (N_5141,N_4878,N_4855);
nand U5142 (N_5142,N_4779,N_4862);
and U5143 (N_5143,N_4665,N_4546);
nor U5144 (N_5144,N_4601,N_4513);
and U5145 (N_5145,N_4660,N_4889);
nor U5146 (N_5146,N_4936,N_4732);
xor U5147 (N_5147,N_4989,N_4654);
or U5148 (N_5148,N_4939,N_4659);
or U5149 (N_5149,N_4522,N_4594);
nor U5150 (N_5150,N_4726,N_4504);
or U5151 (N_5151,N_4833,N_4711);
and U5152 (N_5152,N_4681,N_4895);
and U5153 (N_5153,N_4608,N_4664);
nor U5154 (N_5154,N_4843,N_4772);
or U5155 (N_5155,N_4960,N_4778);
nor U5156 (N_5156,N_4649,N_4876);
nor U5157 (N_5157,N_4595,N_4615);
and U5158 (N_5158,N_4516,N_4937);
xnor U5159 (N_5159,N_4502,N_4658);
or U5160 (N_5160,N_4567,N_4644);
and U5161 (N_5161,N_4925,N_4836);
or U5162 (N_5162,N_4768,N_4540);
nand U5163 (N_5163,N_4775,N_4784);
or U5164 (N_5164,N_4872,N_4750);
nor U5165 (N_5165,N_4948,N_4532);
or U5166 (N_5166,N_4789,N_4716);
and U5167 (N_5167,N_4919,N_4809);
or U5168 (N_5168,N_4912,N_4687);
nor U5169 (N_5169,N_4861,N_4624);
or U5170 (N_5170,N_4846,N_4764);
nor U5171 (N_5171,N_4675,N_4921);
xor U5172 (N_5172,N_4508,N_4795);
nor U5173 (N_5173,N_4737,N_4617);
and U5174 (N_5174,N_4526,N_4765);
nand U5175 (N_5175,N_4696,N_4904);
and U5176 (N_5176,N_4805,N_4680);
nand U5177 (N_5177,N_4600,N_4688);
or U5178 (N_5178,N_4701,N_4558);
nor U5179 (N_5179,N_4882,N_4552);
and U5180 (N_5180,N_4999,N_4509);
nor U5181 (N_5181,N_4563,N_4799);
and U5182 (N_5182,N_4930,N_4964);
and U5183 (N_5183,N_4995,N_4738);
or U5184 (N_5184,N_4666,N_4771);
or U5185 (N_5185,N_4854,N_4852);
nand U5186 (N_5186,N_4668,N_4524);
or U5187 (N_5187,N_4788,N_4651);
and U5188 (N_5188,N_4888,N_4500);
nor U5189 (N_5189,N_4712,N_4956);
nand U5190 (N_5190,N_4975,N_4632);
nor U5191 (N_5191,N_4723,N_4951);
and U5192 (N_5192,N_4901,N_4968);
xor U5193 (N_5193,N_4980,N_4945);
or U5194 (N_5194,N_4955,N_4736);
nand U5195 (N_5195,N_4709,N_4797);
and U5196 (N_5196,N_4741,N_4742);
or U5197 (N_5197,N_4747,N_4748);
nand U5198 (N_5198,N_4652,N_4802);
and U5199 (N_5199,N_4974,N_4971);
and U5200 (N_5200,N_4599,N_4991);
nor U5201 (N_5201,N_4603,N_4677);
nor U5202 (N_5202,N_4557,N_4672);
and U5203 (N_5203,N_4634,N_4816);
nor U5204 (N_5204,N_4785,N_4886);
and U5205 (N_5205,N_4637,N_4510);
and U5206 (N_5206,N_4731,N_4656);
nor U5207 (N_5207,N_4695,N_4959);
nor U5208 (N_5208,N_4903,N_4730);
nand U5209 (N_5209,N_4835,N_4523);
nor U5210 (N_5210,N_4591,N_4794);
nand U5211 (N_5211,N_4756,N_4691);
nand U5212 (N_5212,N_4827,N_4829);
nor U5213 (N_5213,N_4987,N_4871);
or U5214 (N_5214,N_4757,N_4571);
nand U5215 (N_5215,N_4745,N_4830);
and U5216 (N_5216,N_4851,N_4585);
and U5217 (N_5217,N_4894,N_4990);
nor U5218 (N_5218,N_4607,N_4929);
nor U5219 (N_5219,N_4576,N_4800);
nor U5220 (N_5220,N_4754,N_4635);
nor U5221 (N_5221,N_4840,N_4934);
and U5222 (N_5222,N_4605,N_4963);
and U5223 (N_5223,N_4942,N_4729);
nand U5224 (N_5224,N_4507,N_4684);
nor U5225 (N_5225,N_4515,N_4928);
and U5226 (N_5226,N_4900,N_4686);
nand U5227 (N_5227,N_4984,N_4587);
nand U5228 (N_5228,N_4897,N_4679);
or U5229 (N_5229,N_4806,N_4517);
and U5230 (N_5230,N_4957,N_4961);
nor U5231 (N_5231,N_4755,N_4793);
and U5232 (N_5232,N_4544,N_4831);
nor U5233 (N_5233,N_4694,N_4531);
nor U5234 (N_5234,N_4551,N_4714);
nand U5235 (N_5235,N_4561,N_4514);
nor U5236 (N_5236,N_4881,N_4602);
and U5237 (N_5237,N_4533,N_4706);
or U5238 (N_5238,N_4728,N_4570);
nor U5239 (N_5239,N_4916,N_4671);
nor U5240 (N_5240,N_4733,N_4623);
or U5241 (N_5241,N_4744,N_4626);
nand U5242 (N_5242,N_4922,N_4941);
nor U5243 (N_5243,N_4630,N_4952);
and U5244 (N_5244,N_4808,N_4910);
nand U5245 (N_5245,N_4976,N_4550);
nand U5246 (N_5246,N_4826,N_4704);
or U5247 (N_5247,N_4822,N_4810);
and U5248 (N_5248,N_4841,N_4670);
nand U5249 (N_5249,N_4891,N_4940);
nor U5250 (N_5250,N_4838,N_4733);
or U5251 (N_5251,N_4516,N_4956);
nand U5252 (N_5252,N_4957,N_4780);
or U5253 (N_5253,N_4772,N_4680);
nand U5254 (N_5254,N_4876,N_4510);
nor U5255 (N_5255,N_4587,N_4512);
nand U5256 (N_5256,N_4925,N_4829);
xnor U5257 (N_5257,N_4633,N_4734);
nor U5258 (N_5258,N_4939,N_4592);
and U5259 (N_5259,N_4865,N_4565);
nor U5260 (N_5260,N_4893,N_4850);
or U5261 (N_5261,N_4971,N_4798);
nor U5262 (N_5262,N_4597,N_4634);
and U5263 (N_5263,N_4525,N_4768);
nand U5264 (N_5264,N_4768,N_4984);
xor U5265 (N_5265,N_4762,N_4651);
and U5266 (N_5266,N_4692,N_4835);
and U5267 (N_5267,N_4908,N_4838);
or U5268 (N_5268,N_4523,N_4509);
or U5269 (N_5269,N_4642,N_4998);
and U5270 (N_5270,N_4536,N_4533);
nand U5271 (N_5271,N_4873,N_4597);
nor U5272 (N_5272,N_4630,N_4766);
nor U5273 (N_5273,N_4743,N_4763);
nor U5274 (N_5274,N_4892,N_4755);
nor U5275 (N_5275,N_4908,N_4710);
or U5276 (N_5276,N_4551,N_4833);
nand U5277 (N_5277,N_4718,N_4809);
nor U5278 (N_5278,N_4872,N_4677);
or U5279 (N_5279,N_4654,N_4889);
or U5280 (N_5280,N_4872,N_4844);
or U5281 (N_5281,N_4763,N_4772);
nor U5282 (N_5282,N_4836,N_4691);
nor U5283 (N_5283,N_4866,N_4727);
or U5284 (N_5284,N_4983,N_4620);
or U5285 (N_5285,N_4513,N_4745);
nor U5286 (N_5286,N_4644,N_4519);
or U5287 (N_5287,N_4677,N_4996);
nor U5288 (N_5288,N_4909,N_4929);
nor U5289 (N_5289,N_4830,N_4992);
xor U5290 (N_5290,N_4574,N_4877);
nand U5291 (N_5291,N_4935,N_4739);
nor U5292 (N_5292,N_4801,N_4811);
nor U5293 (N_5293,N_4759,N_4566);
nor U5294 (N_5294,N_4886,N_4699);
and U5295 (N_5295,N_4854,N_4868);
nor U5296 (N_5296,N_4994,N_4682);
nand U5297 (N_5297,N_4540,N_4601);
or U5298 (N_5298,N_4850,N_4681);
nand U5299 (N_5299,N_4605,N_4846);
and U5300 (N_5300,N_4700,N_4505);
nand U5301 (N_5301,N_4647,N_4975);
and U5302 (N_5302,N_4938,N_4648);
or U5303 (N_5303,N_4895,N_4692);
and U5304 (N_5304,N_4696,N_4621);
nand U5305 (N_5305,N_4648,N_4892);
or U5306 (N_5306,N_4645,N_4899);
and U5307 (N_5307,N_4960,N_4503);
or U5308 (N_5308,N_4795,N_4780);
xnor U5309 (N_5309,N_4910,N_4550);
or U5310 (N_5310,N_4540,N_4851);
and U5311 (N_5311,N_4542,N_4655);
and U5312 (N_5312,N_4756,N_4685);
or U5313 (N_5313,N_4574,N_4758);
nor U5314 (N_5314,N_4774,N_4725);
nand U5315 (N_5315,N_4629,N_4960);
or U5316 (N_5316,N_4624,N_4696);
and U5317 (N_5317,N_4509,N_4874);
nand U5318 (N_5318,N_4877,N_4896);
and U5319 (N_5319,N_4787,N_4676);
nor U5320 (N_5320,N_4538,N_4876);
nor U5321 (N_5321,N_4919,N_4921);
nand U5322 (N_5322,N_4553,N_4874);
and U5323 (N_5323,N_4684,N_4792);
nand U5324 (N_5324,N_4794,N_4817);
or U5325 (N_5325,N_4703,N_4925);
or U5326 (N_5326,N_4640,N_4865);
nand U5327 (N_5327,N_4778,N_4555);
nand U5328 (N_5328,N_4908,N_4681);
and U5329 (N_5329,N_4581,N_4607);
and U5330 (N_5330,N_4660,N_4895);
nor U5331 (N_5331,N_4819,N_4969);
nand U5332 (N_5332,N_4876,N_4961);
and U5333 (N_5333,N_4980,N_4524);
nand U5334 (N_5334,N_4967,N_4946);
nand U5335 (N_5335,N_4946,N_4754);
nand U5336 (N_5336,N_4763,N_4565);
nand U5337 (N_5337,N_4633,N_4819);
and U5338 (N_5338,N_4643,N_4914);
and U5339 (N_5339,N_4533,N_4939);
and U5340 (N_5340,N_4675,N_4605);
nand U5341 (N_5341,N_4999,N_4936);
and U5342 (N_5342,N_4510,N_4622);
nand U5343 (N_5343,N_4555,N_4747);
xnor U5344 (N_5344,N_4708,N_4974);
and U5345 (N_5345,N_4637,N_4979);
nor U5346 (N_5346,N_4731,N_4562);
nor U5347 (N_5347,N_4787,N_4808);
and U5348 (N_5348,N_4636,N_4516);
nand U5349 (N_5349,N_4801,N_4917);
or U5350 (N_5350,N_4612,N_4938);
nand U5351 (N_5351,N_4796,N_4922);
nand U5352 (N_5352,N_4951,N_4598);
or U5353 (N_5353,N_4911,N_4927);
nor U5354 (N_5354,N_4792,N_4799);
or U5355 (N_5355,N_4730,N_4729);
and U5356 (N_5356,N_4556,N_4626);
or U5357 (N_5357,N_4818,N_4668);
nor U5358 (N_5358,N_4504,N_4623);
and U5359 (N_5359,N_4556,N_4806);
xor U5360 (N_5360,N_4596,N_4745);
and U5361 (N_5361,N_4981,N_4850);
and U5362 (N_5362,N_4982,N_4702);
or U5363 (N_5363,N_4710,N_4848);
nand U5364 (N_5364,N_4833,N_4865);
nand U5365 (N_5365,N_4749,N_4944);
nor U5366 (N_5366,N_4984,N_4573);
or U5367 (N_5367,N_4532,N_4671);
nand U5368 (N_5368,N_4612,N_4538);
nand U5369 (N_5369,N_4504,N_4952);
nor U5370 (N_5370,N_4871,N_4912);
and U5371 (N_5371,N_4733,N_4526);
nor U5372 (N_5372,N_4839,N_4850);
nand U5373 (N_5373,N_4948,N_4984);
nand U5374 (N_5374,N_4844,N_4854);
and U5375 (N_5375,N_4853,N_4655);
or U5376 (N_5376,N_4598,N_4605);
nand U5377 (N_5377,N_4648,N_4594);
nand U5378 (N_5378,N_4904,N_4743);
xor U5379 (N_5379,N_4932,N_4806);
and U5380 (N_5380,N_4619,N_4524);
and U5381 (N_5381,N_4738,N_4897);
nor U5382 (N_5382,N_4603,N_4534);
or U5383 (N_5383,N_4778,N_4981);
nand U5384 (N_5384,N_4802,N_4770);
nand U5385 (N_5385,N_4930,N_4616);
and U5386 (N_5386,N_4754,N_4776);
nand U5387 (N_5387,N_4954,N_4589);
or U5388 (N_5388,N_4524,N_4685);
nand U5389 (N_5389,N_4611,N_4710);
and U5390 (N_5390,N_4600,N_4755);
nor U5391 (N_5391,N_4532,N_4770);
and U5392 (N_5392,N_4866,N_4840);
or U5393 (N_5393,N_4803,N_4677);
and U5394 (N_5394,N_4722,N_4999);
nor U5395 (N_5395,N_4615,N_4770);
or U5396 (N_5396,N_4951,N_4990);
and U5397 (N_5397,N_4986,N_4632);
or U5398 (N_5398,N_4532,N_4709);
nor U5399 (N_5399,N_4972,N_4621);
and U5400 (N_5400,N_4696,N_4683);
or U5401 (N_5401,N_4958,N_4862);
or U5402 (N_5402,N_4842,N_4574);
nor U5403 (N_5403,N_4629,N_4673);
nand U5404 (N_5404,N_4629,N_4911);
nor U5405 (N_5405,N_4879,N_4520);
or U5406 (N_5406,N_4705,N_4957);
and U5407 (N_5407,N_4515,N_4503);
nor U5408 (N_5408,N_4742,N_4974);
and U5409 (N_5409,N_4992,N_4957);
or U5410 (N_5410,N_4717,N_4776);
nor U5411 (N_5411,N_4802,N_4701);
and U5412 (N_5412,N_4950,N_4680);
and U5413 (N_5413,N_4577,N_4802);
and U5414 (N_5414,N_4722,N_4877);
nor U5415 (N_5415,N_4860,N_4726);
and U5416 (N_5416,N_4684,N_4850);
nor U5417 (N_5417,N_4913,N_4597);
nand U5418 (N_5418,N_4911,N_4693);
or U5419 (N_5419,N_4704,N_4707);
nand U5420 (N_5420,N_4584,N_4607);
or U5421 (N_5421,N_4647,N_4530);
and U5422 (N_5422,N_4830,N_4770);
nand U5423 (N_5423,N_4811,N_4837);
nor U5424 (N_5424,N_4646,N_4932);
nor U5425 (N_5425,N_4931,N_4640);
nand U5426 (N_5426,N_4580,N_4790);
or U5427 (N_5427,N_4783,N_4589);
or U5428 (N_5428,N_4833,N_4898);
nand U5429 (N_5429,N_4722,N_4981);
nor U5430 (N_5430,N_4964,N_4590);
and U5431 (N_5431,N_4697,N_4834);
and U5432 (N_5432,N_4584,N_4997);
or U5433 (N_5433,N_4925,N_4774);
nor U5434 (N_5434,N_4755,N_4604);
and U5435 (N_5435,N_4602,N_4615);
and U5436 (N_5436,N_4960,N_4807);
nor U5437 (N_5437,N_4764,N_4552);
or U5438 (N_5438,N_4637,N_4793);
or U5439 (N_5439,N_4878,N_4635);
and U5440 (N_5440,N_4578,N_4916);
or U5441 (N_5441,N_4888,N_4513);
or U5442 (N_5442,N_4608,N_4990);
nand U5443 (N_5443,N_4736,N_4855);
or U5444 (N_5444,N_4995,N_4565);
nand U5445 (N_5445,N_4543,N_4716);
nor U5446 (N_5446,N_4905,N_4713);
nand U5447 (N_5447,N_4882,N_4645);
or U5448 (N_5448,N_4622,N_4812);
nor U5449 (N_5449,N_4710,N_4860);
xnor U5450 (N_5450,N_4693,N_4650);
nor U5451 (N_5451,N_4759,N_4574);
nand U5452 (N_5452,N_4840,N_4618);
nor U5453 (N_5453,N_4847,N_4659);
nor U5454 (N_5454,N_4528,N_4848);
or U5455 (N_5455,N_4652,N_4712);
nor U5456 (N_5456,N_4981,N_4766);
nand U5457 (N_5457,N_4772,N_4933);
nor U5458 (N_5458,N_4521,N_4662);
nand U5459 (N_5459,N_4965,N_4977);
and U5460 (N_5460,N_4842,N_4651);
and U5461 (N_5461,N_4889,N_4770);
and U5462 (N_5462,N_4920,N_4788);
or U5463 (N_5463,N_4512,N_4759);
or U5464 (N_5464,N_4972,N_4570);
nand U5465 (N_5465,N_4600,N_4959);
nor U5466 (N_5466,N_4638,N_4892);
nand U5467 (N_5467,N_4810,N_4873);
nand U5468 (N_5468,N_4958,N_4517);
nand U5469 (N_5469,N_4660,N_4965);
nand U5470 (N_5470,N_4794,N_4574);
xor U5471 (N_5471,N_4536,N_4660);
and U5472 (N_5472,N_4930,N_4702);
nor U5473 (N_5473,N_4546,N_4992);
or U5474 (N_5474,N_4773,N_4663);
nand U5475 (N_5475,N_4724,N_4767);
nand U5476 (N_5476,N_4774,N_4926);
nor U5477 (N_5477,N_4901,N_4616);
and U5478 (N_5478,N_4782,N_4693);
and U5479 (N_5479,N_4919,N_4819);
or U5480 (N_5480,N_4861,N_4994);
nand U5481 (N_5481,N_4851,N_4926);
nand U5482 (N_5482,N_4692,N_4535);
or U5483 (N_5483,N_4629,N_4636);
nor U5484 (N_5484,N_4882,N_4680);
and U5485 (N_5485,N_4566,N_4561);
nand U5486 (N_5486,N_4581,N_4530);
nand U5487 (N_5487,N_4646,N_4556);
xnor U5488 (N_5488,N_4889,N_4964);
nor U5489 (N_5489,N_4752,N_4890);
or U5490 (N_5490,N_4680,N_4730);
nand U5491 (N_5491,N_4924,N_4887);
and U5492 (N_5492,N_4971,N_4510);
and U5493 (N_5493,N_4973,N_4999);
nand U5494 (N_5494,N_4568,N_4555);
nor U5495 (N_5495,N_4858,N_4542);
or U5496 (N_5496,N_4917,N_4837);
and U5497 (N_5497,N_4929,N_4641);
nand U5498 (N_5498,N_4612,N_4662);
nor U5499 (N_5499,N_4981,N_4658);
nor U5500 (N_5500,N_5115,N_5455);
nand U5501 (N_5501,N_5394,N_5092);
or U5502 (N_5502,N_5047,N_5492);
or U5503 (N_5503,N_5320,N_5112);
nor U5504 (N_5504,N_5379,N_5341);
or U5505 (N_5505,N_5241,N_5045);
xor U5506 (N_5506,N_5421,N_5063);
or U5507 (N_5507,N_5037,N_5064);
or U5508 (N_5508,N_5058,N_5025);
nand U5509 (N_5509,N_5152,N_5444);
nor U5510 (N_5510,N_5287,N_5149);
or U5511 (N_5511,N_5384,N_5484);
nand U5512 (N_5512,N_5452,N_5436);
and U5513 (N_5513,N_5318,N_5263);
nor U5514 (N_5514,N_5148,N_5357);
nand U5515 (N_5515,N_5103,N_5479);
or U5516 (N_5516,N_5284,N_5162);
nor U5517 (N_5517,N_5191,N_5268);
or U5518 (N_5518,N_5186,N_5435);
nor U5519 (N_5519,N_5406,N_5293);
nor U5520 (N_5520,N_5105,N_5121);
or U5521 (N_5521,N_5294,N_5478);
and U5522 (N_5522,N_5317,N_5041);
nor U5523 (N_5523,N_5480,N_5381);
or U5524 (N_5524,N_5082,N_5091);
nor U5525 (N_5525,N_5183,N_5039);
nand U5526 (N_5526,N_5274,N_5044);
nor U5527 (N_5527,N_5368,N_5457);
or U5528 (N_5528,N_5032,N_5449);
nor U5529 (N_5529,N_5077,N_5342);
nor U5530 (N_5530,N_5225,N_5004);
nand U5531 (N_5531,N_5024,N_5173);
and U5532 (N_5532,N_5288,N_5218);
or U5533 (N_5533,N_5232,N_5249);
nor U5534 (N_5534,N_5314,N_5431);
or U5535 (N_5535,N_5494,N_5270);
or U5536 (N_5536,N_5476,N_5203);
nor U5537 (N_5537,N_5172,N_5206);
or U5538 (N_5538,N_5223,N_5151);
and U5539 (N_5539,N_5350,N_5062);
nor U5540 (N_5540,N_5427,N_5266);
and U5541 (N_5541,N_5482,N_5323);
or U5542 (N_5542,N_5193,N_5477);
or U5543 (N_5543,N_5168,N_5271);
nand U5544 (N_5544,N_5201,N_5345);
and U5545 (N_5545,N_5275,N_5154);
xnor U5546 (N_5546,N_5396,N_5362);
or U5547 (N_5547,N_5009,N_5185);
and U5548 (N_5548,N_5269,N_5461);
nand U5549 (N_5549,N_5158,N_5087);
or U5550 (N_5550,N_5034,N_5170);
nand U5551 (N_5551,N_5175,N_5391);
nand U5552 (N_5552,N_5367,N_5422);
nor U5553 (N_5553,N_5289,N_5131);
nand U5554 (N_5554,N_5013,N_5330);
nor U5555 (N_5555,N_5303,N_5048);
and U5556 (N_5556,N_5007,N_5003);
or U5557 (N_5557,N_5377,N_5408);
or U5558 (N_5558,N_5385,N_5414);
nand U5559 (N_5559,N_5182,N_5069);
nand U5560 (N_5560,N_5002,N_5160);
and U5561 (N_5561,N_5043,N_5205);
or U5562 (N_5562,N_5022,N_5207);
nand U5563 (N_5563,N_5051,N_5403);
nand U5564 (N_5564,N_5230,N_5277);
nor U5565 (N_5565,N_5420,N_5297);
or U5566 (N_5566,N_5358,N_5272);
and U5567 (N_5567,N_5417,N_5333);
or U5568 (N_5568,N_5176,N_5231);
or U5569 (N_5569,N_5397,N_5061);
nor U5570 (N_5570,N_5393,N_5008);
or U5571 (N_5571,N_5361,N_5080);
nor U5572 (N_5572,N_5120,N_5329);
nand U5573 (N_5573,N_5015,N_5111);
nor U5574 (N_5574,N_5295,N_5319);
nand U5575 (N_5575,N_5486,N_5095);
or U5576 (N_5576,N_5071,N_5059);
nand U5577 (N_5577,N_5456,N_5311);
and U5578 (N_5578,N_5215,N_5171);
or U5579 (N_5579,N_5369,N_5497);
or U5580 (N_5580,N_5038,N_5244);
nor U5581 (N_5581,N_5331,N_5286);
or U5582 (N_5582,N_5030,N_5363);
nor U5583 (N_5583,N_5247,N_5102);
and U5584 (N_5584,N_5260,N_5014);
nor U5585 (N_5585,N_5254,N_5267);
or U5586 (N_5586,N_5220,N_5027);
or U5587 (N_5587,N_5094,N_5138);
xnor U5588 (N_5588,N_5156,N_5219);
nor U5589 (N_5589,N_5181,N_5147);
or U5590 (N_5590,N_5150,N_5400);
or U5591 (N_5591,N_5387,N_5221);
or U5592 (N_5592,N_5125,N_5302);
nor U5593 (N_5593,N_5235,N_5439);
nor U5594 (N_5594,N_5113,N_5290);
nand U5595 (N_5595,N_5026,N_5285);
or U5596 (N_5596,N_5118,N_5140);
xnor U5597 (N_5597,N_5458,N_5093);
nand U5598 (N_5598,N_5401,N_5360);
and U5599 (N_5599,N_5243,N_5016);
or U5600 (N_5600,N_5465,N_5257);
and U5601 (N_5601,N_5386,N_5453);
or U5602 (N_5602,N_5473,N_5296);
and U5603 (N_5603,N_5169,N_5307);
and U5604 (N_5604,N_5259,N_5124);
or U5605 (N_5605,N_5432,N_5404);
nor U5606 (N_5606,N_5460,N_5495);
and U5607 (N_5607,N_5159,N_5264);
or U5608 (N_5608,N_5310,N_5141);
or U5609 (N_5609,N_5233,N_5145);
nand U5610 (N_5610,N_5212,N_5279);
and U5611 (N_5611,N_5142,N_5299);
xor U5612 (N_5612,N_5018,N_5445);
nor U5613 (N_5613,N_5190,N_5410);
nand U5614 (N_5614,N_5070,N_5312);
or U5615 (N_5615,N_5447,N_5119);
and U5616 (N_5616,N_5174,N_5443);
nand U5617 (N_5617,N_5122,N_5086);
and U5618 (N_5618,N_5129,N_5011);
or U5619 (N_5619,N_5356,N_5382);
nand U5620 (N_5620,N_5265,N_5315);
or U5621 (N_5621,N_5019,N_5425);
nor U5622 (N_5622,N_5472,N_5462);
or U5623 (N_5623,N_5348,N_5078);
and U5624 (N_5624,N_5165,N_5155);
and U5625 (N_5625,N_5338,N_5202);
nand U5626 (N_5626,N_5236,N_5208);
and U5627 (N_5627,N_5075,N_5245);
and U5628 (N_5628,N_5251,N_5390);
nor U5629 (N_5629,N_5237,N_5454);
nor U5630 (N_5630,N_5132,N_5375);
nor U5631 (N_5631,N_5413,N_5049);
and U5632 (N_5632,N_5372,N_5424);
nand U5633 (N_5633,N_5109,N_5389);
nor U5634 (N_5634,N_5446,N_5126);
nor U5635 (N_5635,N_5352,N_5136);
and U5636 (N_5636,N_5035,N_5128);
nor U5637 (N_5637,N_5180,N_5388);
nand U5638 (N_5638,N_5496,N_5110);
and U5639 (N_5639,N_5252,N_5184);
and U5640 (N_5640,N_5104,N_5199);
nand U5641 (N_5641,N_5485,N_5085);
and U5642 (N_5642,N_5426,N_5399);
nand U5643 (N_5643,N_5306,N_5336);
and U5644 (N_5644,N_5304,N_5281);
nand U5645 (N_5645,N_5050,N_5261);
and U5646 (N_5646,N_5209,N_5188);
or U5647 (N_5647,N_5239,N_5227);
nand U5648 (N_5648,N_5402,N_5409);
nor U5649 (N_5649,N_5380,N_5098);
and U5650 (N_5650,N_5346,N_5498);
or U5651 (N_5651,N_5166,N_5229);
nand U5652 (N_5652,N_5493,N_5434);
or U5653 (N_5653,N_5405,N_5052);
and U5654 (N_5654,N_5195,N_5090);
nand U5655 (N_5655,N_5114,N_5033);
or U5656 (N_5656,N_5471,N_5134);
nor U5657 (N_5657,N_5108,N_5029);
nand U5658 (N_5658,N_5468,N_5101);
nor U5659 (N_5659,N_5300,N_5097);
and U5660 (N_5660,N_5234,N_5353);
nor U5661 (N_5661,N_5242,N_5060);
nand U5662 (N_5662,N_5322,N_5343);
nand U5663 (N_5663,N_5433,N_5466);
and U5664 (N_5664,N_5163,N_5001);
and U5665 (N_5665,N_5258,N_5366);
or U5666 (N_5666,N_5339,N_5179);
nand U5667 (N_5667,N_5189,N_5351);
and U5668 (N_5668,N_5238,N_5328);
and U5669 (N_5669,N_5324,N_5076);
nand U5670 (N_5670,N_5450,N_5196);
or U5671 (N_5671,N_5255,N_5489);
nand U5672 (N_5672,N_5068,N_5423);
or U5673 (N_5673,N_5211,N_5475);
and U5674 (N_5674,N_5214,N_5240);
or U5675 (N_5675,N_5490,N_5084);
or U5676 (N_5676,N_5153,N_5056);
or U5677 (N_5677,N_5040,N_5398);
nand U5678 (N_5678,N_5481,N_5222);
and U5679 (N_5679,N_5276,N_5364);
nor U5680 (N_5680,N_5347,N_5415);
or U5681 (N_5681,N_5157,N_5074);
and U5682 (N_5682,N_5079,N_5020);
and U5683 (N_5683,N_5428,N_5370);
nand U5684 (N_5684,N_5010,N_5253);
or U5685 (N_5685,N_5135,N_5204);
nor U5686 (N_5686,N_5216,N_5292);
and U5687 (N_5687,N_5055,N_5117);
nand U5688 (N_5688,N_5349,N_5248);
or U5689 (N_5689,N_5213,N_5451);
and U5690 (N_5690,N_5187,N_5143);
nand U5691 (N_5691,N_5429,N_5441);
nor U5692 (N_5692,N_5066,N_5042);
nor U5693 (N_5693,N_5440,N_5072);
nand U5694 (N_5694,N_5392,N_5021);
nand U5695 (N_5695,N_5167,N_5028);
nor U5696 (N_5696,N_5407,N_5464);
nor U5697 (N_5697,N_5116,N_5430);
nor U5698 (N_5698,N_5096,N_5127);
nand U5699 (N_5699,N_5337,N_5133);
nor U5700 (N_5700,N_5335,N_5448);
nor U5701 (N_5701,N_5359,N_5365);
and U5702 (N_5702,N_5298,N_5228);
and U5703 (N_5703,N_5144,N_5470);
and U5704 (N_5704,N_5332,N_5067);
and U5705 (N_5705,N_5073,N_5419);
or U5706 (N_5706,N_5130,N_5226);
or U5707 (N_5707,N_5262,N_5474);
nor U5708 (N_5708,N_5469,N_5278);
or U5709 (N_5709,N_5194,N_5442);
or U5710 (N_5710,N_5418,N_5334);
and U5711 (N_5711,N_5099,N_5100);
or U5712 (N_5712,N_5054,N_5023);
nand U5713 (N_5713,N_5164,N_5107);
and U5714 (N_5714,N_5081,N_5467);
or U5715 (N_5715,N_5354,N_5313);
nor U5716 (N_5716,N_5005,N_5309);
or U5717 (N_5717,N_5210,N_5499);
nor U5718 (N_5718,N_5161,N_5411);
nor U5719 (N_5719,N_5316,N_5178);
nand U5720 (N_5720,N_5017,N_5283);
nand U5721 (N_5721,N_5177,N_5246);
or U5722 (N_5722,N_5373,N_5282);
or U5723 (N_5723,N_5378,N_5280);
or U5724 (N_5724,N_5291,N_5463);
or U5725 (N_5725,N_5437,N_5198);
nor U5726 (N_5726,N_5137,N_5301);
or U5727 (N_5727,N_5256,N_5344);
nand U5728 (N_5728,N_5491,N_5438);
or U5729 (N_5729,N_5326,N_5139);
and U5730 (N_5730,N_5273,N_5325);
nand U5731 (N_5731,N_5340,N_5488);
nand U5732 (N_5732,N_5371,N_5146);
nand U5733 (N_5733,N_5305,N_5192);
nand U5734 (N_5734,N_5065,N_5057);
nor U5735 (N_5735,N_5083,N_5321);
nand U5736 (N_5736,N_5416,N_5383);
and U5737 (N_5737,N_5197,N_5376);
or U5738 (N_5738,N_5006,N_5088);
nand U5739 (N_5739,N_5355,N_5327);
nand U5740 (N_5740,N_5012,N_5106);
and U5741 (N_5741,N_5046,N_5123);
nor U5742 (N_5742,N_5487,N_5483);
or U5743 (N_5743,N_5089,N_5395);
nor U5744 (N_5744,N_5031,N_5200);
nor U5745 (N_5745,N_5053,N_5308);
and U5746 (N_5746,N_5036,N_5000);
or U5747 (N_5747,N_5374,N_5459);
or U5748 (N_5748,N_5412,N_5217);
and U5749 (N_5749,N_5250,N_5224);
nor U5750 (N_5750,N_5488,N_5419);
and U5751 (N_5751,N_5048,N_5003);
nor U5752 (N_5752,N_5231,N_5161);
nor U5753 (N_5753,N_5143,N_5271);
nand U5754 (N_5754,N_5012,N_5455);
and U5755 (N_5755,N_5138,N_5496);
nand U5756 (N_5756,N_5060,N_5290);
xor U5757 (N_5757,N_5069,N_5164);
nor U5758 (N_5758,N_5159,N_5318);
and U5759 (N_5759,N_5170,N_5471);
and U5760 (N_5760,N_5200,N_5423);
nand U5761 (N_5761,N_5381,N_5212);
nand U5762 (N_5762,N_5432,N_5028);
nor U5763 (N_5763,N_5461,N_5420);
or U5764 (N_5764,N_5373,N_5433);
nand U5765 (N_5765,N_5169,N_5187);
or U5766 (N_5766,N_5023,N_5072);
nor U5767 (N_5767,N_5024,N_5151);
nor U5768 (N_5768,N_5098,N_5293);
nand U5769 (N_5769,N_5279,N_5012);
nor U5770 (N_5770,N_5211,N_5431);
or U5771 (N_5771,N_5332,N_5496);
or U5772 (N_5772,N_5324,N_5023);
xor U5773 (N_5773,N_5283,N_5118);
or U5774 (N_5774,N_5017,N_5020);
and U5775 (N_5775,N_5370,N_5409);
nand U5776 (N_5776,N_5034,N_5151);
or U5777 (N_5777,N_5104,N_5406);
and U5778 (N_5778,N_5161,N_5342);
nor U5779 (N_5779,N_5096,N_5469);
nand U5780 (N_5780,N_5278,N_5207);
and U5781 (N_5781,N_5357,N_5013);
nor U5782 (N_5782,N_5314,N_5103);
or U5783 (N_5783,N_5250,N_5472);
nand U5784 (N_5784,N_5102,N_5260);
nand U5785 (N_5785,N_5205,N_5059);
nand U5786 (N_5786,N_5060,N_5167);
or U5787 (N_5787,N_5347,N_5055);
or U5788 (N_5788,N_5480,N_5143);
and U5789 (N_5789,N_5292,N_5370);
or U5790 (N_5790,N_5090,N_5043);
nand U5791 (N_5791,N_5351,N_5238);
or U5792 (N_5792,N_5085,N_5288);
or U5793 (N_5793,N_5047,N_5417);
or U5794 (N_5794,N_5280,N_5310);
nor U5795 (N_5795,N_5449,N_5385);
and U5796 (N_5796,N_5220,N_5431);
or U5797 (N_5797,N_5487,N_5136);
and U5798 (N_5798,N_5496,N_5428);
and U5799 (N_5799,N_5224,N_5497);
or U5800 (N_5800,N_5038,N_5331);
and U5801 (N_5801,N_5041,N_5270);
nor U5802 (N_5802,N_5214,N_5202);
or U5803 (N_5803,N_5292,N_5483);
nor U5804 (N_5804,N_5325,N_5096);
nand U5805 (N_5805,N_5225,N_5381);
nor U5806 (N_5806,N_5338,N_5402);
or U5807 (N_5807,N_5179,N_5028);
xnor U5808 (N_5808,N_5362,N_5350);
nand U5809 (N_5809,N_5120,N_5304);
and U5810 (N_5810,N_5413,N_5483);
nand U5811 (N_5811,N_5478,N_5386);
nor U5812 (N_5812,N_5405,N_5278);
xnor U5813 (N_5813,N_5189,N_5194);
or U5814 (N_5814,N_5323,N_5388);
and U5815 (N_5815,N_5039,N_5396);
or U5816 (N_5816,N_5148,N_5045);
and U5817 (N_5817,N_5060,N_5359);
and U5818 (N_5818,N_5171,N_5139);
or U5819 (N_5819,N_5414,N_5116);
nand U5820 (N_5820,N_5024,N_5266);
nand U5821 (N_5821,N_5309,N_5491);
nand U5822 (N_5822,N_5293,N_5257);
or U5823 (N_5823,N_5150,N_5336);
nor U5824 (N_5824,N_5226,N_5063);
nor U5825 (N_5825,N_5463,N_5132);
nor U5826 (N_5826,N_5192,N_5165);
nor U5827 (N_5827,N_5212,N_5009);
or U5828 (N_5828,N_5406,N_5210);
nand U5829 (N_5829,N_5385,N_5128);
and U5830 (N_5830,N_5381,N_5120);
and U5831 (N_5831,N_5136,N_5428);
or U5832 (N_5832,N_5485,N_5043);
xnor U5833 (N_5833,N_5046,N_5473);
nand U5834 (N_5834,N_5120,N_5491);
nor U5835 (N_5835,N_5352,N_5393);
nor U5836 (N_5836,N_5189,N_5376);
or U5837 (N_5837,N_5240,N_5016);
and U5838 (N_5838,N_5292,N_5412);
nor U5839 (N_5839,N_5049,N_5081);
nand U5840 (N_5840,N_5160,N_5264);
or U5841 (N_5841,N_5127,N_5497);
and U5842 (N_5842,N_5247,N_5138);
nand U5843 (N_5843,N_5195,N_5254);
nor U5844 (N_5844,N_5074,N_5340);
or U5845 (N_5845,N_5310,N_5238);
and U5846 (N_5846,N_5117,N_5238);
and U5847 (N_5847,N_5116,N_5264);
or U5848 (N_5848,N_5159,N_5397);
and U5849 (N_5849,N_5290,N_5278);
or U5850 (N_5850,N_5093,N_5303);
or U5851 (N_5851,N_5071,N_5022);
or U5852 (N_5852,N_5390,N_5038);
nor U5853 (N_5853,N_5071,N_5498);
nor U5854 (N_5854,N_5296,N_5119);
or U5855 (N_5855,N_5000,N_5176);
and U5856 (N_5856,N_5305,N_5287);
or U5857 (N_5857,N_5173,N_5262);
or U5858 (N_5858,N_5271,N_5419);
nor U5859 (N_5859,N_5465,N_5090);
nand U5860 (N_5860,N_5211,N_5479);
nand U5861 (N_5861,N_5045,N_5304);
and U5862 (N_5862,N_5489,N_5168);
and U5863 (N_5863,N_5458,N_5128);
nor U5864 (N_5864,N_5121,N_5469);
and U5865 (N_5865,N_5234,N_5255);
nand U5866 (N_5866,N_5349,N_5275);
nor U5867 (N_5867,N_5263,N_5083);
or U5868 (N_5868,N_5071,N_5015);
nand U5869 (N_5869,N_5348,N_5041);
and U5870 (N_5870,N_5436,N_5471);
or U5871 (N_5871,N_5208,N_5369);
nor U5872 (N_5872,N_5009,N_5288);
nand U5873 (N_5873,N_5252,N_5079);
nand U5874 (N_5874,N_5386,N_5365);
nor U5875 (N_5875,N_5195,N_5196);
nand U5876 (N_5876,N_5319,N_5335);
nand U5877 (N_5877,N_5030,N_5039);
nor U5878 (N_5878,N_5217,N_5338);
and U5879 (N_5879,N_5128,N_5112);
and U5880 (N_5880,N_5424,N_5107);
and U5881 (N_5881,N_5408,N_5073);
nor U5882 (N_5882,N_5362,N_5427);
nand U5883 (N_5883,N_5340,N_5204);
nand U5884 (N_5884,N_5036,N_5416);
nand U5885 (N_5885,N_5412,N_5400);
and U5886 (N_5886,N_5329,N_5398);
and U5887 (N_5887,N_5336,N_5025);
nor U5888 (N_5888,N_5254,N_5362);
nor U5889 (N_5889,N_5377,N_5460);
nor U5890 (N_5890,N_5389,N_5373);
or U5891 (N_5891,N_5020,N_5144);
nand U5892 (N_5892,N_5231,N_5480);
nor U5893 (N_5893,N_5428,N_5066);
nor U5894 (N_5894,N_5302,N_5101);
nand U5895 (N_5895,N_5451,N_5034);
or U5896 (N_5896,N_5267,N_5155);
nor U5897 (N_5897,N_5324,N_5303);
nor U5898 (N_5898,N_5224,N_5122);
nand U5899 (N_5899,N_5173,N_5358);
and U5900 (N_5900,N_5145,N_5160);
or U5901 (N_5901,N_5351,N_5458);
nor U5902 (N_5902,N_5493,N_5121);
and U5903 (N_5903,N_5135,N_5473);
nand U5904 (N_5904,N_5478,N_5092);
nand U5905 (N_5905,N_5333,N_5033);
nand U5906 (N_5906,N_5091,N_5284);
nand U5907 (N_5907,N_5021,N_5075);
or U5908 (N_5908,N_5060,N_5341);
nor U5909 (N_5909,N_5484,N_5271);
and U5910 (N_5910,N_5276,N_5275);
or U5911 (N_5911,N_5441,N_5139);
and U5912 (N_5912,N_5181,N_5283);
or U5913 (N_5913,N_5394,N_5371);
nand U5914 (N_5914,N_5093,N_5030);
or U5915 (N_5915,N_5112,N_5184);
or U5916 (N_5916,N_5008,N_5045);
nand U5917 (N_5917,N_5426,N_5144);
and U5918 (N_5918,N_5328,N_5080);
or U5919 (N_5919,N_5154,N_5047);
and U5920 (N_5920,N_5118,N_5264);
and U5921 (N_5921,N_5226,N_5444);
xor U5922 (N_5922,N_5040,N_5436);
and U5923 (N_5923,N_5014,N_5440);
or U5924 (N_5924,N_5047,N_5062);
or U5925 (N_5925,N_5044,N_5019);
or U5926 (N_5926,N_5013,N_5000);
nand U5927 (N_5927,N_5063,N_5143);
and U5928 (N_5928,N_5432,N_5403);
nand U5929 (N_5929,N_5196,N_5283);
nor U5930 (N_5930,N_5477,N_5036);
nor U5931 (N_5931,N_5479,N_5306);
nor U5932 (N_5932,N_5130,N_5493);
and U5933 (N_5933,N_5145,N_5435);
nor U5934 (N_5934,N_5214,N_5406);
nand U5935 (N_5935,N_5415,N_5481);
nor U5936 (N_5936,N_5361,N_5417);
nor U5937 (N_5937,N_5000,N_5077);
and U5938 (N_5938,N_5445,N_5363);
nor U5939 (N_5939,N_5216,N_5104);
and U5940 (N_5940,N_5262,N_5430);
and U5941 (N_5941,N_5270,N_5157);
xnor U5942 (N_5942,N_5293,N_5022);
or U5943 (N_5943,N_5123,N_5062);
nor U5944 (N_5944,N_5360,N_5393);
and U5945 (N_5945,N_5448,N_5215);
nor U5946 (N_5946,N_5257,N_5158);
or U5947 (N_5947,N_5116,N_5269);
nor U5948 (N_5948,N_5242,N_5110);
or U5949 (N_5949,N_5229,N_5171);
and U5950 (N_5950,N_5361,N_5085);
nor U5951 (N_5951,N_5210,N_5126);
and U5952 (N_5952,N_5107,N_5122);
and U5953 (N_5953,N_5329,N_5025);
nand U5954 (N_5954,N_5158,N_5131);
nand U5955 (N_5955,N_5189,N_5146);
or U5956 (N_5956,N_5301,N_5400);
or U5957 (N_5957,N_5254,N_5253);
and U5958 (N_5958,N_5228,N_5290);
nor U5959 (N_5959,N_5323,N_5005);
and U5960 (N_5960,N_5377,N_5363);
xor U5961 (N_5961,N_5349,N_5432);
or U5962 (N_5962,N_5325,N_5192);
nand U5963 (N_5963,N_5274,N_5431);
nand U5964 (N_5964,N_5297,N_5146);
and U5965 (N_5965,N_5041,N_5194);
xnor U5966 (N_5966,N_5288,N_5496);
and U5967 (N_5967,N_5026,N_5156);
and U5968 (N_5968,N_5054,N_5213);
or U5969 (N_5969,N_5254,N_5164);
nand U5970 (N_5970,N_5320,N_5183);
or U5971 (N_5971,N_5264,N_5092);
nand U5972 (N_5972,N_5419,N_5097);
xor U5973 (N_5973,N_5200,N_5078);
or U5974 (N_5974,N_5190,N_5083);
nand U5975 (N_5975,N_5332,N_5108);
and U5976 (N_5976,N_5408,N_5329);
and U5977 (N_5977,N_5322,N_5232);
or U5978 (N_5978,N_5349,N_5069);
or U5979 (N_5979,N_5139,N_5285);
xnor U5980 (N_5980,N_5059,N_5038);
and U5981 (N_5981,N_5329,N_5306);
or U5982 (N_5982,N_5025,N_5230);
nor U5983 (N_5983,N_5184,N_5318);
and U5984 (N_5984,N_5490,N_5408);
nor U5985 (N_5985,N_5163,N_5363);
nand U5986 (N_5986,N_5481,N_5173);
nand U5987 (N_5987,N_5313,N_5059);
and U5988 (N_5988,N_5483,N_5331);
xor U5989 (N_5989,N_5256,N_5115);
and U5990 (N_5990,N_5039,N_5056);
nor U5991 (N_5991,N_5432,N_5459);
and U5992 (N_5992,N_5126,N_5473);
or U5993 (N_5993,N_5267,N_5160);
nand U5994 (N_5994,N_5121,N_5041);
nand U5995 (N_5995,N_5078,N_5144);
nand U5996 (N_5996,N_5442,N_5083);
or U5997 (N_5997,N_5233,N_5469);
nand U5998 (N_5998,N_5442,N_5114);
nor U5999 (N_5999,N_5345,N_5265);
and U6000 (N_6000,N_5999,N_5880);
or U6001 (N_6001,N_5670,N_5510);
nand U6002 (N_6002,N_5816,N_5676);
or U6003 (N_6003,N_5671,N_5612);
or U6004 (N_6004,N_5761,N_5511);
nand U6005 (N_6005,N_5754,N_5663);
or U6006 (N_6006,N_5698,N_5645);
nand U6007 (N_6007,N_5700,N_5956);
nand U6008 (N_6008,N_5689,N_5746);
or U6009 (N_6009,N_5872,N_5642);
and U6010 (N_6010,N_5686,N_5807);
nand U6011 (N_6011,N_5554,N_5934);
nor U6012 (N_6012,N_5734,N_5650);
nand U6013 (N_6013,N_5944,N_5602);
nor U6014 (N_6014,N_5531,N_5738);
or U6015 (N_6015,N_5742,N_5916);
or U6016 (N_6016,N_5898,N_5792);
or U6017 (N_6017,N_5727,N_5585);
or U6018 (N_6018,N_5767,N_5917);
or U6019 (N_6019,N_5955,N_5744);
or U6020 (N_6020,N_5803,N_5790);
and U6021 (N_6021,N_5566,N_5843);
or U6022 (N_6022,N_5993,N_5674);
nor U6023 (N_6023,N_5597,N_5827);
and U6024 (N_6024,N_5969,N_5682);
or U6025 (N_6025,N_5909,N_5977);
and U6026 (N_6026,N_5683,N_5929);
nor U6027 (N_6027,N_5756,N_5695);
nand U6028 (N_6028,N_5551,N_5813);
or U6029 (N_6029,N_5576,N_5802);
nand U6030 (N_6030,N_5693,N_5509);
nor U6031 (N_6031,N_5811,N_5637);
nor U6032 (N_6032,N_5945,N_5640);
nand U6033 (N_6033,N_5719,N_5728);
and U6034 (N_6034,N_5900,N_5873);
nand U6035 (N_6035,N_5829,N_5966);
and U6036 (N_6036,N_5610,N_5634);
or U6037 (N_6037,N_5992,N_5986);
nand U6038 (N_6038,N_5899,N_5621);
or U6039 (N_6039,N_5745,N_5548);
or U6040 (N_6040,N_5893,N_5623);
nand U6041 (N_6041,N_5948,N_5764);
nand U6042 (N_6042,N_5794,N_5501);
nor U6043 (N_6043,N_5889,N_5527);
nand U6044 (N_6044,N_5595,N_5523);
and U6045 (N_6045,N_5500,N_5841);
nand U6046 (N_6046,N_5903,N_5805);
nand U6047 (N_6047,N_5681,N_5517);
nand U6048 (N_6048,N_5839,N_5935);
nand U6049 (N_6049,N_5987,N_5796);
and U6050 (N_6050,N_5861,N_5836);
nor U6051 (N_6051,N_5776,N_5543);
or U6052 (N_6052,N_5658,N_5592);
nor U6053 (N_6053,N_5895,N_5562);
or U6054 (N_6054,N_5506,N_5743);
or U6055 (N_6055,N_5820,N_5518);
nand U6056 (N_6056,N_5897,N_5888);
or U6057 (N_6057,N_5582,N_5710);
or U6058 (N_6058,N_5636,N_5835);
nand U6059 (N_6059,N_5863,N_5546);
nor U6060 (N_6060,N_5782,N_5603);
or U6061 (N_6061,N_5516,N_5559);
xnor U6062 (N_6062,N_5971,N_5979);
xnor U6063 (N_6063,N_5780,N_5949);
or U6064 (N_6064,N_5750,N_5660);
nor U6065 (N_6065,N_5726,N_5923);
nand U6066 (N_6066,N_5731,N_5667);
nor U6067 (N_6067,N_5529,N_5706);
or U6068 (N_6068,N_5614,N_5959);
nand U6069 (N_6069,N_5797,N_5534);
nand U6070 (N_6070,N_5665,N_5618);
nor U6071 (N_6071,N_5646,N_5926);
and U6072 (N_6072,N_5675,N_5937);
nor U6073 (N_6073,N_5677,N_5608);
and U6074 (N_6074,N_5963,N_5615);
or U6075 (N_6075,N_5639,N_5910);
nand U6076 (N_6076,N_5657,N_5522);
and U6077 (N_6077,N_5870,N_5537);
nand U6078 (N_6078,N_5655,N_5564);
or U6079 (N_6079,N_5567,N_5672);
or U6080 (N_6080,N_5994,N_5584);
nor U6081 (N_6081,N_5775,N_5632);
and U6082 (N_6082,N_5881,N_5985);
nor U6083 (N_6083,N_5656,N_5882);
nand U6084 (N_6084,N_5644,N_5659);
nand U6085 (N_6085,N_5611,N_5749);
and U6086 (N_6086,N_5512,N_5707);
nor U6087 (N_6087,N_5814,N_5572);
or U6088 (N_6088,N_5856,N_5647);
nand U6089 (N_6089,N_5950,N_5624);
nor U6090 (N_6090,N_5730,N_5828);
or U6091 (N_6091,N_5840,N_5718);
nand U6092 (N_6092,N_5740,N_5823);
or U6093 (N_6093,N_5504,N_5515);
and U6094 (N_6094,N_5654,N_5855);
and U6095 (N_6095,N_5544,N_5942);
nor U6096 (N_6096,N_5673,N_5601);
nor U6097 (N_6097,N_5704,N_5692);
or U6098 (N_6098,N_5535,N_5765);
or U6099 (N_6099,N_5877,N_5806);
or U6100 (N_6100,N_5505,N_5625);
or U6101 (N_6101,N_5812,N_5968);
nand U6102 (N_6102,N_5555,N_5751);
or U6103 (N_6103,N_5715,N_5589);
nand U6104 (N_6104,N_5770,N_5653);
nand U6105 (N_6105,N_5894,N_5859);
or U6106 (N_6106,N_5778,N_5842);
nand U6107 (N_6107,N_5560,N_5561);
and U6108 (N_6108,N_5771,N_5834);
nor U6109 (N_6109,N_5911,N_5631);
nand U6110 (N_6110,N_5857,N_5540);
and U6111 (N_6111,N_5865,N_5871);
nand U6112 (N_6112,N_5789,N_5787);
nand U6113 (N_6113,N_5701,N_5846);
or U6114 (N_6114,N_5613,N_5581);
nor U6115 (N_6115,N_5599,N_5661);
and U6116 (N_6116,N_5961,N_5697);
xnor U6117 (N_6117,N_5586,N_5784);
nor U6118 (N_6118,N_5568,N_5924);
nor U6119 (N_6119,N_5801,N_5960);
or U6120 (N_6120,N_5606,N_5652);
and U6121 (N_6121,N_5616,N_5587);
nor U6122 (N_6122,N_5635,N_5884);
and U6123 (N_6123,N_5600,N_5702);
and U6124 (N_6124,N_5556,N_5574);
nand U6125 (N_6125,N_5521,N_5763);
and U6126 (N_6126,N_5699,N_5804);
nand U6127 (N_6127,N_5712,N_5970);
and U6128 (N_6128,N_5539,N_5541);
or U6129 (N_6129,N_5912,N_5902);
or U6130 (N_6130,N_5684,N_5844);
and U6131 (N_6131,N_5925,N_5837);
and U6132 (N_6132,N_5831,N_5641);
nand U6133 (N_6133,N_5685,N_5739);
nor U6134 (N_6134,N_5777,N_5988);
and U6135 (N_6135,N_5849,N_5799);
or U6136 (N_6136,N_5502,N_5946);
nand U6137 (N_6137,N_5668,N_5905);
and U6138 (N_6138,N_5896,N_5920);
and U6139 (N_6139,N_5536,N_5991);
nor U6140 (N_6140,N_5847,N_5533);
nand U6141 (N_6141,N_5547,N_5725);
and U6142 (N_6142,N_5818,N_5648);
or U6143 (N_6143,N_5591,N_5759);
and U6144 (N_6144,N_5891,N_5729);
nand U6145 (N_6145,N_5943,N_5957);
nor U6146 (N_6146,N_5976,N_5519);
and U6147 (N_6147,N_5952,N_5983);
nor U6148 (N_6148,N_5732,N_5679);
and U6149 (N_6149,N_5958,N_5760);
and U6150 (N_6150,N_5830,N_5542);
and U6151 (N_6151,N_5622,N_5904);
or U6152 (N_6152,N_5724,N_5965);
or U6153 (N_6153,N_5748,N_5810);
nand U6154 (N_6154,N_5680,N_5617);
nand U6155 (N_6155,N_5954,N_5953);
nand U6156 (N_6156,N_5705,N_5711);
nand U6157 (N_6157,N_5975,N_5577);
nor U6158 (N_6158,N_5703,N_5785);
nand U6159 (N_6159,N_5569,N_5620);
nand U6160 (N_6160,N_5514,N_5972);
nor U6161 (N_6161,N_5598,N_5793);
nor U6162 (N_6162,N_5850,N_5768);
nor U6163 (N_6163,N_5526,N_5919);
nand U6164 (N_6164,N_5908,N_5995);
nor U6165 (N_6165,N_5819,N_5821);
nand U6166 (N_6166,N_5688,N_5938);
or U6167 (N_6167,N_5552,N_5513);
xor U6168 (N_6168,N_5982,N_5575);
or U6169 (N_6169,N_5887,N_5753);
nand U6170 (N_6170,N_5538,N_5981);
nor U6171 (N_6171,N_5525,N_5503);
nor U6172 (N_6172,N_5878,N_5752);
nand U6173 (N_6173,N_5558,N_5716);
or U6174 (N_6174,N_5628,N_5978);
and U6175 (N_6175,N_5875,N_5845);
nor U6176 (N_6176,N_5666,N_5824);
or U6177 (N_6177,N_5858,N_5649);
or U6178 (N_6178,N_5741,N_5769);
nand U6179 (N_6179,N_5643,N_5713);
and U6180 (N_6180,N_5890,N_5973);
and U6181 (N_6181,N_5570,N_5723);
and U6182 (N_6182,N_5809,N_5596);
or U6183 (N_6183,N_5578,N_5867);
or U6184 (N_6184,N_5808,N_5918);
or U6185 (N_6185,N_5691,N_5879);
nand U6186 (N_6186,N_5930,N_5984);
nand U6187 (N_6187,N_5990,N_5951);
and U6188 (N_6188,N_5714,N_5530);
and U6189 (N_6189,N_5678,N_5662);
nor U6190 (N_6190,N_5694,N_5869);
nand U6191 (N_6191,N_5781,N_5866);
or U6192 (N_6192,N_5507,N_5573);
xnor U6193 (N_6193,N_5757,N_5996);
nor U6194 (N_6194,N_5579,N_5528);
and U6195 (N_6195,N_5580,N_5627);
and U6196 (N_6196,N_5874,N_5901);
nand U6197 (N_6197,N_5721,N_5928);
or U6198 (N_6198,N_5633,N_5669);
or U6199 (N_6199,N_5583,N_5594);
nor U6200 (N_6200,N_5520,N_5892);
and U6201 (N_6201,N_5974,N_5630);
or U6202 (N_6202,N_5876,N_5832);
xor U6203 (N_6203,N_5906,N_5779);
nor U6204 (N_6204,N_5860,N_5619);
nand U6205 (N_6205,N_5854,N_5788);
and U6206 (N_6206,N_5815,N_5549);
nor U6207 (N_6207,N_5800,N_5997);
xnor U6208 (N_6208,N_5914,N_5626);
nor U6209 (N_6209,N_5921,N_5588);
nand U6210 (N_6210,N_5629,N_5817);
nor U6211 (N_6211,N_5825,N_5696);
nor U6212 (N_6212,N_5786,N_5798);
and U6213 (N_6213,N_5593,N_5783);
nand U6214 (N_6214,N_5605,N_5931);
nand U6215 (N_6215,N_5720,N_5736);
or U6216 (N_6216,N_5795,N_5737);
nand U6217 (N_6217,N_5638,N_5563);
nor U6218 (N_6218,N_5651,N_5962);
nor U6219 (N_6219,N_5690,N_5709);
nand U6220 (N_6220,N_5885,N_5604);
nand U6221 (N_6221,N_5913,N_5758);
or U6222 (N_6222,N_5989,N_5853);
nor U6223 (N_6223,N_5833,N_5545);
xor U6224 (N_6224,N_5851,N_5571);
and U6225 (N_6225,N_5848,N_5941);
and U6226 (N_6226,N_5852,N_5557);
and U6227 (N_6227,N_5773,N_5927);
nand U6228 (N_6228,N_5947,N_5762);
nand U6229 (N_6229,N_5722,N_5862);
or U6230 (N_6230,N_5550,N_5964);
or U6231 (N_6231,N_5907,N_5607);
nor U6232 (N_6232,N_5967,N_5980);
nand U6233 (N_6233,N_5733,N_5936);
nand U6234 (N_6234,N_5932,N_5933);
or U6235 (N_6235,N_5524,N_5922);
and U6236 (N_6236,N_5717,N_5532);
and U6237 (N_6237,N_5998,N_5664);
and U6238 (N_6238,N_5590,N_5838);
or U6239 (N_6239,N_5708,N_5883);
and U6240 (N_6240,N_5826,N_5609);
and U6241 (N_6241,N_5508,N_5766);
and U6242 (N_6242,N_5791,N_5774);
nor U6243 (N_6243,N_5565,N_5735);
and U6244 (N_6244,N_5868,N_5864);
nand U6245 (N_6245,N_5747,N_5915);
and U6246 (N_6246,N_5940,N_5939);
nand U6247 (N_6247,N_5886,N_5822);
or U6248 (N_6248,N_5553,N_5687);
xor U6249 (N_6249,N_5755,N_5772);
or U6250 (N_6250,N_5878,N_5559);
nor U6251 (N_6251,N_5913,N_5786);
nand U6252 (N_6252,N_5709,N_5973);
nor U6253 (N_6253,N_5780,N_5609);
and U6254 (N_6254,N_5943,N_5898);
or U6255 (N_6255,N_5805,N_5528);
nand U6256 (N_6256,N_5698,N_5810);
nand U6257 (N_6257,N_5607,N_5711);
or U6258 (N_6258,N_5544,N_5641);
nor U6259 (N_6259,N_5903,N_5538);
or U6260 (N_6260,N_5631,N_5804);
nor U6261 (N_6261,N_5772,N_5577);
xor U6262 (N_6262,N_5665,N_5532);
nor U6263 (N_6263,N_5745,N_5797);
nor U6264 (N_6264,N_5860,N_5834);
nor U6265 (N_6265,N_5760,N_5875);
nor U6266 (N_6266,N_5657,N_5733);
nor U6267 (N_6267,N_5665,N_5543);
nand U6268 (N_6268,N_5560,N_5503);
and U6269 (N_6269,N_5894,N_5960);
nor U6270 (N_6270,N_5762,N_5865);
nand U6271 (N_6271,N_5580,N_5976);
nand U6272 (N_6272,N_5663,N_5715);
and U6273 (N_6273,N_5721,N_5651);
and U6274 (N_6274,N_5719,N_5759);
and U6275 (N_6275,N_5783,N_5771);
nand U6276 (N_6276,N_5769,N_5663);
or U6277 (N_6277,N_5762,N_5863);
or U6278 (N_6278,N_5573,N_5781);
nand U6279 (N_6279,N_5714,N_5556);
nand U6280 (N_6280,N_5743,N_5742);
nand U6281 (N_6281,N_5835,N_5820);
or U6282 (N_6282,N_5509,N_5901);
or U6283 (N_6283,N_5727,N_5884);
or U6284 (N_6284,N_5583,N_5816);
or U6285 (N_6285,N_5908,N_5741);
nand U6286 (N_6286,N_5637,N_5577);
or U6287 (N_6287,N_5560,N_5755);
nand U6288 (N_6288,N_5588,N_5603);
or U6289 (N_6289,N_5650,N_5502);
xnor U6290 (N_6290,N_5636,N_5727);
and U6291 (N_6291,N_5622,N_5627);
nand U6292 (N_6292,N_5897,N_5580);
or U6293 (N_6293,N_5777,N_5813);
nor U6294 (N_6294,N_5907,N_5734);
and U6295 (N_6295,N_5729,N_5804);
nor U6296 (N_6296,N_5890,N_5659);
nand U6297 (N_6297,N_5584,N_5503);
or U6298 (N_6298,N_5748,N_5970);
or U6299 (N_6299,N_5964,N_5693);
nand U6300 (N_6300,N_5523,N_5993);
and U6301 (N_6301,N_5802,N_5940);
and U6302 (N_6302,N_5754,N_5863);
or U6303 (N_6303,N_5935,N_5519);
xor U6304 (N_6304,N_5836,N_5906);
nor U6305 (N_6305,N_5582,N_5853);
nor U6306 (N_6306,N_5578,N_5655);
or U6307 (N_6307,N_5551,N_5956);
and U6308 (N_6308,N_5543,N_5996);
nor U6309 (N_6309,N_5759,N_5903);
or U6310 (N_6310,N_5650,N_5950);
or U6311 (N_6311,N_5879,N_5698);
and U6312 (N_6312,N_5713,N_5699);
or U6313 (N_6313,N_5842,N_5609);
and U6314 (N_6314,N_5968,N_5702);
nor U6315 (N_6315,N_5988,N_5674);
xnor U6316 (N_6316,N_5860,N_5666);
and U6317 (N_6317,N_5650,N_5934);
nand U6318 (N_6318,N_5604,N_5994);
nor U6319 (N_6319,N_5981,N_5773);
nand U6320 (N_6320,N_5877,N_5535);
nor U6321 (N_6321,N_5869,N_5986);
or U6322 (N_6322,N_5688,N_5713);
nor U6323 (N_6323,N_5859,N_5617);
or U6324 (N_6324,N_5880,N_5871);
and U6325 (N_6325,N_5946,N_5725);
and U6326 (N_6326,N_5728,N_5717);
nor U6327 (N_6327,N_5538,N_5549);
nor U6328 (N_6328,N_5610,N_5727);
and U6329 (N_6329,N_5991,N_5811);
and U6330 (N_6330,N_5566,N_5793);
or U6331 (N_6331,N_5532,N_5813);
and U6332 (N_6332,N_5717,N_5637);
or U6333 (N_6333,N_5537,N_5924);
nor U6334 (N_6334,N_5720,N_5524);
or U6335 (N_6335,N_5893,N_5941);
nand U6336 (N_6336,N_5871,N_5928);
nand U6337 (N_6337,N_5985,N_5860);
or U6338 (N_6338,N_5809,N_5814);
and U6339 (N_6339,N_5943,N_5833);
nand U6340 (N_6340,N_5677,N_5526);
nor U6341 (N_6341,N_5988,N_5924);
nor U6342 (N_6342,N_5726,N_5706);
or U6343 (N_6343,N_5702,N_5764);
nand U6344 (N_6344,N_5655,N_5758);
nor U6345 (N_6345,N_5878,N_5881);
nand U6346 (N_6346,N_5565,N_5827);
nand U6347 (N_6347,N_5502,N_5606);
xor U6348 (N_6348,N_5610,N_5510);
nand U6349 (N_6349,N_5631,N_5975);
nand U6350 (N_6350,N_5695,N_5740);
nand U6351 (N_6351,N_5713,N_5604);
nor U6352 (N_6352,N_5639,N_5832);
and U6353 (N_6353,N_5907,N_5623);
and U6354 (N_6354,N_5936,N_5515);
nand U6355 (N_6355,N_5977,N_5983);
and U6356 (N_6356,N_5757,N_5594);
or U6357 (N_6357,N_5737,N_5763);
nor U6358 (N_6358,N_5634,N_5872);
nand U6359 (N_6359,N_5616,N_5643);
xnor U6360 (N_6360,N_5660,N_5949);
nor U6361 (N_6361,N_5649,N_5993);
and U6362 (N_6362,N_5523,N_5937);
nand U6363 (N_6363,N_5933,N_5714);
or U6364 (N_6364,N_5745,N_5895);
nor U6365 (N_6365,N_5719,N_5795);
nand U6366 (N_6366,N_5558,N_5764);
nand U6367 (N_6367,N_5975,N_5672);
nand U6368 (N_6368,N_5773,N_5623);
nor U6369 (N_6369,N_5779,N_5766);
nand U6370 (N_6370,N_5664,N_5777);
or U6371 (N_6371,N_5809,N_5505);
nor U6372 (N_6372,N_5652,N_5650);
or U6373 (N_6373,N_5786,N_5683);
nand U6374 (N_6374,N_5795,N_5874);
and U6375 (N_6375,N_5791,N_5514);
nand U6376 (N_6376,N_5976,N_5935);
nor U6377 (N_6377,N_5609,N_5991);
nand U6378 (N_6378,N_5950,N_5899);
nand U6379 (N_6379,N_5852,N_5906);
nor U6380 (N_6380,N_5821,N_5695);
or U6381 (N_6381,N_5718,N_5517);
nand U6382 (N_6382,N_5945,N_5830);
xor U6383 (N_6383,N_5748,N_5566);
or U6384 (N_6384,N_5764,N_5858);
nor U6385 (N_6385,N_5621,N_5664);
and U6386 (N_6386,N_5980,N_5998);
or U6387 (N_6387,N_5618,N_5746);
xnor U6388 (N_6388,N_5853,N_5706);
nor U6389 (N_6389,N_5946,N_5904);
nor U6390 (N_6390,N_5665,N_5668);
nor U6391 (N_6391,N_5663,N_5698);
and U6392 (N_6392,N_5814,N_5962);
and U6393 (N_6393,N_5809,N_5566);
or U6394 (N_6394,N_5672,N_5528);
or U6395 (N_6395,N_5590,N_5604);
xor U6396 (N_6396,N_5969,N_5689);
nand U6397 (N_6397,N_5787,N_5973);
and U6398 (N_6398,N_5511,N_5806);
or U6399 (N_6399,N_5891,N_5908);
nor U6400 (N_6400,N_5722,N_5724);
nor U6401 (N_6401,N_5838,N_5812);
nand U6402 (N_6402,N_5565,N_5622);
nand U6403 (N_6403,N_5821,N_5783);
or U6404 (N_6404,N_5872,N_5896);
or U6405 (N_6405,N_5609,N_5793);
nand U6406 (N_6406,N_5763,N_5782);
and U6407 (N_6407,N_5920,N_5784);
or U6408 (N_6408,N_5950,N_5891);
and U6409 (N_6409,N_5688,N_5764);
and U6410 (N_6410,N_5728,N_5876);
xnor U6411 (N_6411,N_5513,N_5534);
or U6412 (N_6412,N_5579,N_5749);
nor U6413 (N_6413,N_5580,N_5805);
or U6414 (N_6414,N_5990,N_5919);
nor U6415 (N_6415,N_5850,N_5668);
or U6416 (N_6416,N_5663,N_5977);
nand U6417 (N_6417,N_5934,N_5958);
nand U6418 (N_6418,N_5811,N_5876);
and U6419 (N_6419,N_5557,N_5565);
nor U6420 (N_6420,N_5681,N_5819);
and U6421 (N_6421,N_5679,N_5941);
and U6422 (N_6422,N_5689,N_5518);
and U6423 (N_6423,N_5695,N_5896);
nand U6424 (N_6424,N_5627,N_5620);
nor U6425 (N_6425,N_5922,N_5552);
nor U6426 (N_6426,N_5513,N_5726);
or U6427 (N_6427,N_5887,N_5534);
and U6428 (N_6428,N_5785,N_5797);
and U6429 (N_6429,N_5517,N_5635);
or U6430 (N_6430,N_5556,N_5842);
nor U6431 (N_6431,N_5686,N_5942);
and U6432 (N_6432,N_5515,N_5718);
nor U6433 (N_6433,N_5889,N_5810);
or U6434 (N_6434,N_5648,N_5872);
and U6435 (N_6435,N_5590,N_5638);
or U6436 (N_6436,N_5838,N_5995);
nor U6437 (N_6437,N_5686,N_5675);
nand U6438 (N_6438,N_5846,N_5572);
nand U6439 (N_6439,N_5733,N_5983);
or U6440 (N_6440,N_5646,N_5997);
nand U6441 (N_6441,N_5620,N_5749);
or U6442 (N_6442,N_5526,N_5782);
and U6443 (N_6443,N_5990,N_5509);
or U6444 (N_6444,N_5657,N_5768);
nand U6445 (N_6445,N_5952,N_5683);
or U6446 (N_6446,N_5911,N_5560);
or U6447 (N_6447,N_5678,N_5889);
nand U6448 (N_6448,N_5568,N_5828);
nand U6449 (N_6449,N_5882,N_5568);
nand U6450 (N_6450,N_5947,N_5940);
nand U6451 (N_6451,N_5898,N_5731);
nor U6452 (N_6452,N_5977,N_5563);
nand U6453 (N_6453,N_5605,N_5822);
nand U6454 (N_6454,N_5651,N_5573);
or U6455 (N_6455,N_5991,N_5737);
nand U6456 (N_6456,N_5750,N_5719);
or U6457 (N_6457,N_5561,N_5726);
nor U6458 (N_6458,N_5966,N_5520);
or U6459 (N_6459,N_5686,N_5599);
or U6460 (N_6460,N_5786,N_5541);
nand U6461 (N_6461,N_5730,N_5804);
or U6462 (N_6462,N_5829,N_5890);
and U6463 (N_6463,N_5925,N_5543);
nand U6464 (N_6464,N_5745,N_5543);
nor U6465 (N_6465,N_5875,N_5548);
nand U6466 (N_6466,N_5663,N_5747);
nor U6467 (N_6467,N_5589,N_5704);
nor U6468 (N_6468,N_5834,N_5878);
nor U6469 (N_6469,N_5755,N_5870);
and U6470 (N_6470,N_5751,N_5845);
nand U6471 (N_6471,N_5971,N_5839);
or U6472 (N_6472,N_5507,N_5896);
or U6473 (N_6473,N_5924,N_5955);
nand U6474 (N_6474,N_5896,N_5581);
and U6475 (N_6475,N_5742,N_5724);
and U6476 (N_6476,N_5613,N_5632);
or U6477 (N_6477,N_5591,N_5578);
xor U6478 (N_6478,N_5802,N_5509);
nor U6479 (N_6479,N_5568,N_5981);
and U6480 (N_6480,N_5768,N_5909);
and U6481 (N_6481,N_5572,N_5797);
nand U6482 (N_6482,N_5852,N_5946);
nand U6483 (N_6483,N_5960,N_5937);
or U6484 (N_6484,N_5631,N_5732);
nand U6485 (N_6485,N_5729,N_5661);
xnor U6486 (N_6486,N_5752,N_5994);
or U6487 (N_6487,N_5736,N_5876);
nand U6488 (N_6488,N_5593,N_5722);
nand U6489 (N_6489,N_5836,N_5865);
nor U6490 (N_6490,N_5632,N_5822);
nor U6491 (N_6491,N_5836,N_5910);
nor U6492 (N_6492,N_5590,N_5911);
nand U6493 (N_6493,N_5660,N_5894);
and U6494 (N_6494,N_5637,N_5967);
and U6495 (N_6495,N_5671,N_5745);
nor U6496 (N_6496,N_5748,N_5700);
nor U6497 (N_6497,N_5721,N_5904);
and U6498 (N_6498,N_5687,N_5600);
nand U6499 (N_6499,N_5763,N_5802);
and U6500 (N_6500,N_6148,N_6477);
or U6501 (N_6501,N_6163,N_6198);
or U6502 (N_6502,N_6373,N_6174);
or U6503 (N_6503,N_6172,N_6106);
nor U6504 (N_6504,N_6103,N_6001);
nor U6505 (N_6505,N_6279,N_6259);
and U6506 (N_6506,N_6293,N_6067);
nor U6507 (N_6507,N_6117,N_6335);
and U6508 (N_6508,N_6239,N_6384);
or U6509 (N_6509,N_6202,N_6395);
nor U6510 (N_6510,N_6421,N_6402);
or U6511 (N_6511,N_6015,N_6314);
or U6512 (N_6512,N_6256,N_6466);
and U6513 (N_6513,N_6344,N_6127);
nor U6514 (N_6514,N_6330,N_6320);
nor U6515 (N_6515,N_6418,N_6084);
nand U6516 (N_6516,N_6371,N_6283);
and U6517 (N_6517,N_6407,N_6058);
nand U6518 (N_6518,N_6463,N_6444);
xnor U6519 (N_6519,N_6438,N_6302);
and U6520 (N_6520,N_6312,N_6240);
and U6521 (N_6521,N_6383,N_6009);
nand U6522 (N_6522,N_6059,N_6204);
and U6523 (N_6523,N_6190,N_6471);
and U6524 (N_6524,N_6265,N_6455);
nor U6525 (N_6525,N_6218,N_6213);
nand U6526 (N_6526,N_6237,N_6439);
or U6527 (N_6527,N_6269,N_6416);
nor U6528 (N_6528,N_6028,N_6219);
or U6529 (N_6529,N_6031,N_6456);
nand U6530 (N_6530,N_6257,N_6496);
or U6531 (N_6531,N_6020,N_6398);
nand U6532 (N_6532,N_6199,N_6183);
nand U6533 (N_6533,N_6404,N_6113);
or U6534 (N_6534,N_6227,N_6484);
and U6535 (N_6535,N_6173,N_6436);
nand U6536 (N_6536,N_6136,N_6372);
and U6537 (N_6537,N_6331,N_6222);
nor U6538 (N_6538,N_6369,N_6073);
or U6539 (N_6539,N_6038,N_6128);
nor U6540 (N_6540,N_6425,N_6268);
nand U6541 (N_6541,N_6286,N_6003);
nand U6542 (N_6542,N_6005,N_6196);
and U6543 (N_6543,N_6068,N_6147);
and U6544 (N_6544,N_6332,N_6493);
nand U6545 (N_6545,N_6182,N_6276);
nand U6546 (N_6546,N_6132,N_6441);
nor U6547 (N_6547,N_6055,N_6270);
nor U6548 (N_6548,N_6299,N_6318);
nor U6549 (N_6549,N_6004,N_6029);
and U6550 (N_6550,N_6111,N_6470);
or U6551 (N_6551,N_6390,N_6062);
or U6552 (N_6552,N_6216,N_6448);
or U6553 (N_6553,N_6426,N_6053);
or U6554 (N_6554,N_6467,N_6008);
nand U6555 (N_6555,N_6277,N_6090);
and U6556 (N_6556,N_6074,N_6359);
nand U6557 (N_6557,N_6356,N_6255);
nor U6558 (N_6558,N_6485,N_6487);
nor U6559 (N_6559,N_6480,N_6377);
or U6560 (N_6560,N_6307,N_6306);
nor U6561 (N_6561,N_6245,N_6066);
or U6562 (N_6562,N_6475,N_6429);
or U6563 (N_6563,N_6305,N_6350);
nand U6564 (N_6564,N_6134,N_6251);
nand U6565 (N_6565,N_6181,N_6243);
and U6566 (N_6566,N_6322,N_6178);
xor U6567 (N_6567,N_6288,N_6011);
or U6568 (N_6568,N_6358,N_6378);
nor U6569 (N_6569,N_6042,N_6459);
or U6570 (N_6570,N_6370,N_6201);
nor U6571 (N_6571,N_6121,N_6401);
and U6572 (N_6572,N_6451,N_6267);
or U6573 (N_6573,N_6380,N_6458);
nand U6574 (N_6574,N_6413,N_6221);
and U6575 (N_6575,N_6294,N_6379);
or U6576 (N_6576,N_6056,N_6083);
nor U6577 (N_6577,N_6206,N_6290);
or U6578 (N_6578,N_6076,N_6272);
nor U6579 (N_6579,N_6144,N_6474);
and U6580 (N_6580,N_6108,N_6386);
xor U6581 (N_6581,N_6040,N_6476);
nor U6582 (N_6582,N_6140,N_6046);
or U6583 (N_6583,N_6328,N_6399);
nor U6584 (N_6584,N_6215,N_6497);
or U6585 (N_6585,N_6102,N_6149);
or U6586 (N_6586,N_6273,N_6498);
nor U6587 (N_6587,N_6481,N_6192);
or U6588 (N_6588,N_6397,N_6469);
or U6589 (N_6589,N_6247,N_6316);
or U6590 (N_6590,N_6478,N_6043);
nand U6591 (N_6591,N_6453,N_6394);
nand U6592 (N_6592,N_6156,N_6197);
and U6593 (N_6593,N_6050,N_6080);
xnor U6594 (N_6594,N_6354,N_6006);
nor U6595 (N_6595,N_6142,N_6262);
or U6596 (N_6596,N_6100,N_6440);
nor U6597 (N_6597,N_6443,N_6464);
nor U6598 (N_6598,N_6032,N_6069);
nand U6599 (N_6599,N_6097,N_6363);
and U6600 (N_6600,N_6093,N_6139);
or U6601 (N_6601,N_6408,N_6391);
nor U6602 (N_6602,N_6002,N_6264);
nand U6603 (N_6603,N_6352,N_6234);
or U6604 (N_6604,N_6492,N_6452);
and U6605 (N_6605,N_6168,N_6368);
and U6606 (N_6606,N_6327,N_6057);
or U6607 (N_6607,N_6019,N_6157);
or U6608 (N_6608,N_6315,N_6289);
nor U6609 (N_6609,N_6082,N_6026);
nand U6610 (N_6610,N_6253,N_6249);
or U6611 (N_6611,N_6014,N_6392);
nand U6612 (N_6612,N_6280,N_6292);
nor U6613 (N_6613,N_6472,N_6226);
and U6614 (N_6614,N_6336,N_6349);
nand U6615 (N_6615,N_6342,N_6343);
and U6616 (N_6616,N_6339,N_6027);
nor U6617 (N_6617,N_6217,N_6169);
and U6618 (N_6618,N_6200,N_6152);
nor U6619 (N_6619,N_6462,N_6012);
nand U6620 (N_6620,N_6319,N_6232);
or U6621 (N_6621,N_6039,N_6186);
and U6622 (N_6622,N_6116,N_6007);
nand U6623 (N_6623,N_6329,N_6065);
nand U6624 (N_6624,N_6308,N_6301);
or U6625 (N_6625,N_6271,N_6258);
or U6626 (N_6626,N_6374,N_6044);
or U6627 (N_6627,N_6048,N_6410);
nor U6628 (N_6628,N_6141,N_6387);
or U6629 (N_6629,N_6220,N_6284);
and U6630 (N_6630,N_6291,N_6365);
or U6631 (N_6631,N_6021,N_6094);
or U6632 (N_6632,N_6414,N_6486);
or U6633 (N_6633,N_6023,N_6449);
and U6634 (N_6634,N_6081,N_6252);
nand U6635 (N_6635,N_6110,N_6208);
or U6636 (N_6636,N_6045,N_6236);
xnor U6637 (N_6637,N_6261,N_6010);
or U6638 (N_6638,N_6468,N_6096);
nor U6639 (N_6639,N_6223,N_6211);
or U6640 (N_6640,N_6295,N_6022);
nand U6641 (N_6641,N_6406,N_6346);
nor U6642 (N_6642,N_6278,N_6483);
nor U6643 (N_6643,N_6422,N_6184);
and U6644 (N_6644,N_6311,N_6494);
nand U6645 (N_6645,N_6489,N_6203);
or U6646 (N_6646,N_6437,N_6465);
nand U6647 (N_6647,N_6125,N_6145);
and U6648 (N_6648,N_6423,N_6340);
nor U6649 (N_6649,N_6432,N_6310);
or U6650 (N_6650,N_6088,N_6431);
or U6651 (N_6651,N_6034,N_6054);
nor U6652 (N_6652,N_6499,N_6357);
or U6653 (N_6653,N_6445,N_6018);
nand U6654 (N_6654,N_6360,N_6348);
or U6655 (N_6655,N_6275,N_6176);
and U6656 (N_6656,N_6415,N_6450);
or U6657 (N_6657,N_6341,N_6167);
nor U6658 (N_6658,N_6266,N_6427);
nor U6659 (N_6659,N_6159,N_6160);
and U6660 (N_6660,N_6228,N_6177);
or U6661 (N_6661,N_6274,N_6171);
or U6662 (N_6662,N_6424,N_6325);
nand U6663 (N_6663,N_6114,N_6188);
or U6664 (N_6664,N_6130,N_6324);
or U6665 (N_6665,N_6353,N_6104);
nor U6666 (N_6666,N_6309,N_6131);
or U6667 (N_6667,N_6085,N_6442);
nand U6668 (N_6668,N_6433,N_6495);
and U6669 (N_6669,N_6382,N_6334);
nand U6670 (N_6670,N_6351,N_6000);
and U6671 (N_6671,N_6072,N_6013);
or U6672 (N_6672,N_6036,N_6389);
nor U6673 (N_6673,N_6405,N_6151);
nand U6674 (N_6674,N_6304,N_6297);
nor U6675 (N_6675,N_6347,N_6385);
xor U6676 (N_6676,N_6154,N_6242);
or U6677 (N_6677,N_6099,N_6393);
or U6678 (N_6678,N_6367,N_6428);
and U6679 (N_6679,N_6194,N_6229);
nand U6680 (N_6680,N_6143,N_6138);
nand U6681 (N_6681,N_6230,N_6321);
nand U6682 (N_6682,N_6193,N_6488);
nand U6683 (N_6683,N_6017,N_6079);
and U6684 (N_6684,N_6187,N_6260);
or U6685 (N_6685,N_6482,N_6086);
or U6686 (N_6686,N_6119,N_6430);
nand U6687 (N_6687,N_6388,N_6233);
nor U6688 (N_6688,N_6313,N_6095);
or U6689 (N_6689,N_6375,N_6403);
or U6690 (N_6690,N_6135,N_6175);
nand U6691 (N_6691,N_6191,N_6189);
xnor U6692 (N_6692,N_6241,N_6420);
or U6693 (N_6693,N_6460,N_6248);
or U6694 (N_6694,N_6060,N_6091);
or U6695 (N_6695,N_6089,N_6366);
or U6696 (N_6696,N_6063,N_6323);
or U6697 (N_6697,N_6250,N_6207);
and U6698 (N_6698,N_6212,N_6195);
or U6699 (N_6699,N_6030,N_6118);
and U6700 (N_6700,N_6150,N_6419);
nand U6701 (N_6701,N_6112,N_6285);
nor U6702 (N_6702,N_6109,N_6170);
nand U6703 (N_6703,N_6361,N_6161);
nand U6704 (N_6704,N_6244,N_6123);
nor U6705 (N_6705,N_6396,N_6166);
nand U6706 (N_6706,N_6337,N_6025);
and U6707 (N_6707,N_6446,N_6333);
and U6708 (N_6708,N_6078,N_6298);
or U6709 (N_6709,N_6120,N_6129);
nand U6710 (N_6710,N_6345,N_6461);
and U6711 (N_6711,N_6362,N_6473);
and U6712 (N_6712,N_6179,N_6303);
and U6713 (N_6713,N_6326,N_6035);
and U6714 (N_6714,N_6263,N_6282);
or U6715 (N_6715,N_6454,N_6209);
nand U6716 (N_6716,N_6479,N_6254);
nor U6717 (N_6717,N_6124,N_6409);
or U6718 (N_6718,N_6158,N_6047);
nor U6719 (N_6719,N_6355,N_6051);
and U6720 (N_6720,N_6235,N_6077);
nor U6721 (N_6721,N_6153,N_6435);
nor U6722 (N_6722,N_6064,N_6447);
and U6723 (N_6723,N_6126,N_6364);
or U6724 (N_6724,N_6434,N_6457);
and U6725 (N_6725,N_6155,N_6033);
and U6726 (N_6726,N_6107,N_6338);
nand U6727 (N_6727,N_6164,N_6101);
xnor U6728 (N_6728,N_6412,N_6185);
and U6729 (N_6729,N_6376,N_6317);
nand U6730 (N_6730,N_6417,N_6041);
and U6731 (N_6731,N_6214,N_6092);
nor U6732 (N_6732,N_6281,N_6087);
and U6733 (N_6733,N_6052,N_6071);
and U6734 (N_6734,N_6224,N_6238);
nand U6735 (N_6735,N_6205,N_6381);
nand U6736 (N_6736,N_6490,N_6162);
nand U6737 (N_6737,N_6122,N_6210);
nand U6738 (N_6738,N_6300,N_6146);
or U6739 (N_6739,N_6024,N_6180);
nand U6740 (N_6740,N_6049,N_6115);
nand U6741 (N_6741,N_6061,N_6491);
nor U6742 (N_6742,N_6225,N_6105);
and U6743 (N_6743,N_6400,N_6133);
or U6744 (N_6744,N_6165,N_6075);
nor U6745 (N_6745,N_6287,N_6016);
and U6746 (N_6746,N_6411,N_6137);
nor U6747 (N_6747,N_6231,N_6246);
or U6748 (N_6748,N_6098,N_6296);
nor U6749 (N_6749,N_6037,N_6070);
and U6750 (N_6750,N_6374,N_6311);
or U6751 (N_6751,N_6069,N_6209);
and U6752 (N_6752,N_6198,N_6318);
or U6753 (N_6753,N_6123,N_6397);
nor U6754 (N_6754,N_6375,N_6088);
and U6755 (N_6755,N_6302,N_6399);
nand U6756 (N_6756,N_6363,N_6269);
nor U6757 (N_6757,N_6235,N_6382);
nor U6758 (N_6758,N_6066,N_6076);
nor U6759 (N_6759,N_6268,N_6301);
nand U6760 (N_6760,N_6010,N_6067);
and U6761 (N_6761,N_6413,N_6460);
nor U6762 (N_6762,N_6135,N_6431);
nor U6763 (N_6763,N_6199,N_6493);
nand U6764 (N_6764,N_6185,N_6284);
nor U6765 (N_6765,N_6065,N_6002);
nor U6766 (N_6766,N_6211,N_6485);
nand U6767 (N_6767,N_6011,N_6002);
or U6768 (N_6768,N_6322,N_6350);
or U6769 (N_6769,N_6334,N_6144);
nand U6770 (N_6770,N_6162,N_6190);
nor U6771 (N_6771,N_6151,N_6187);
nor U6772 (N_6772,N_6494,N_6084);
nor U6773 (N_6773,N_6188,N_6241);
nand U6774 (N_6774,N_6215,N_6430);
or U6775 (N_6775,N_6062,N_6495);
nand U6776 (N_6776,N_6441,N_6403);
nor U6777 (N_6777,N_6337,N_6497);
and U6778 (N_6778,N_6089,N_6093);
nor U6779 (N_6779,N_6163,N_6055);
and U6780 (N_6780,N_6222,N_6474);
and U6781 (N_6781,N_6139,N_6176);
nand U6782 (N_6782,N_6316,N_6074);
or U6783 (N_6783,N_6100,N_6168);
nor U6784 (N_6784,N_6487,N_6355);
or U6785 (N_6785,N_6494,N_6195);
nor U6786 (N_6786,N_6030,N_6414);
and U6787 (N_6787,N_6395,N_6315);
nand U6788 (N_6788,N_6290,N_6357);
and U6789 (N_6789,N_6314,N_6495);
nand U6790 (N_6790,N_6485,N_6494);
nand U6791 (N_6791,N_6432,N_6449);
nor U6792 (N_6792,N_6395,N_6080);
nand U6793 (N_6793,N_6449,N_6333);
and U6794 (N_6794,N_6294,N_6040);
and U6795 (N_6795,N_6088,N_6090);
or U6796 (N_6796,N_6123,N_6005);
and U6797 (N_6797,N_6390,N_6055);
nor U6798 (N_6798,N_6168,N_6432);
nor U6799 (N_6799,N_6246,N_6108);
xnor U6800 (N_6800,N_6182,N_6077);
nor U6801 (N_6801,N_6309,N_6283);
nand U6802 (N_6802,N_6354,N_6124);
xnor U6803 (N_6803,N_6392,N_6278);
nand U6804 (N_6804,N_6105,N_6475);
and U6805 (N_6805,N_6317,N_6454);
nor U6806 (N_6806,N_6030,N_6069);
or U6807 (N_6807,N_6316,N_6288);
nor U6808 (N_6808,N_6491,N_6236);
nand U6809 (N_6809,N_6396,N_6395);
or U6810 (N_6810,N_6065,N_6045);
and U6811 (N_6811,N_6329,N_6080);
xor U6812 (N_6812,N_6066,N_6253);
and U6813 (N_6813,N_6271,N_6054);
nand U6814 (N_6814,N_6189,N_6219);
nor U6815 (N_6815,N_6221,N_6401);
nand U6816 (N_6816,N_6072,N_6032);
nor U6817 (N_6817,N_6221,N_6364);
nor U6818 (N_6818,N_6343,N_6252);
or U6819 (N_6819,N_6136,N_6227);
nand U6820 (N_6820,N_6366,N_6495);
or U6821 (N_6821,N_6318,N_6125);
nand U6822 (N_6822,N_6132,N_6224);
nand U6823 (N_6823,N_6016,N_6235);
nand U6824 (N_6824,N_6242,N_6356);
nor U6825 (N_6825,N_6227,N_6157);
and U6826 (N_6826,N_6398,N_6488);
and U6827 (N_6827,N_6134,N_6456);
or U6828 (N_6828,N_6392,N_6317);
or U6829 (N_6829,N_6458,N_6040);
or U6830 (N_6830,N_6429,N_6014);
or U6831 (N_6831,N_6263,N_6209);
nand U6832 (N_6832,N_6458,N_6027);
or U6833 (N_6833,N_6342,N_6007);
nand U6834 (N_6834,N_6231,N_6238);
or U6835 (N_6835,N_6032,N_6473);
nor U6836 (N_6836,N_6409,N_6184);
nor U6837 (N_6837,N_6126,N_6395);
and U6838 (N_6838,N_6146,N_6268);
nand U6839 (N_6839,N_6366,N_6418);
nor U6840 (N_6840,N_6045,N_6113);
nand U6841 (N_6841,N_6450,N_6192);
nor U6842 (N_6842,N_6028,N_6152);
or U6843 (N_6843,N_6421,N_6186);
nor U6844 (N_6844,N_6084,N_6451);
and U6845 (N_6845,N_6361,N_6096);
nand U6846 (N_6846,N_6067,N_6352);
nor U6847 (N_6847,N_6137,N_6127);
nor U6848 (N_6848,N_6177,N_6183);
nor U6849 (N_6849,N_6039,N_6237);
xor U6850 (N_6850,N_6490,N_6487);
and U6851 (N_6851,N_6472,N_6289);
nor U6852 (N_6852,N_6438,N_6474);
and U6853 (N_6853,N_6140,N_6250);
or U6854 (N_6854,N_6295,N_6174);
nand U6855 (N_6855,N_6352,N_6197);
and U6856 (N_6856,N_6278,N_6062);
or U6857 (N_6857,N_6071,N_6105);
or U6858 (N_6858,N_6231,N_6338);
nand U6859 (N_6859,N_6347,N_6251);
and U6860 (N_6860,N_6493,N_6204);
nand U6861 (N_6861,N_6311,N_6267);
xnor U6862 (N_6862,N_6350,N_6436);
nor U6863 (N_6863,N_6298,N_6256);
or U6864 (N_6864,N_6027,N_6424);
or U6865 (N_6865,N_6411,N_6339);
or U6866 (N_6866,N_6111,N_6055);
nor U6867 (N_6867,N_6075,N_6333);
nor U6868 (N_6868,N_6183,N_6314);
or U6869 (N_6869,N_6448,N_6096);
nor U6870 (N_6870,N_6232,N_6322);
nor U6871 (N_6871,N_6474,N_6013);
and U6872 (N_6872,N_6451,N_6335);
and U6873 (N_6873,N_6056,N_6372);
and U6874 (N_6874,N_6410,N_6420);
nand U6875 (N_6875,N_6420,N_6271);
and U6876 (N_6876,N_6222,N_6370);
nor U6877 (N_6877,N_6209,N_6022);
nor U6878 (N_6878,N_6363,N_6354);
and U6879 (N_6879,N_6068,N_6111);
or U6880 (N_6880,N_6146,N_6071);
nor U6881 (N_6881,N_6325,N_6297);
or U6882 (N_6882,N_6213,N_6212);
or U6883 (N_6883,N_6422,N_6061);
or U6884 (N_6884,N_6464,N_6024);
and U6885 (N_6885,N_6261,N_6062);
nor U6886 (N_6886,N_6211,N_6416);
nor U6887 (N_6887,N_6417,N_6341);
nor U6888 (N_6888,N_6285,N_6456);
nor U6889 (N_6889,N_6069,N_6161);
nand U6890 (N_6890,N_6117,N_6166);
nor U6891 (N_6891,N_6395,N_6240);
or U6892 (N_6892,N_6466,N_6088);
and U6893 (N_6893,N_6077,N_6031);
and U6894 (N_6894,N_6291,N_6061);
or U6895 (N_6895,N_6486,N_6381);
nand U6896 (N_6896,N_6164,N_6096);
nand U6897 (N_6897,N_6418,N_6411);
and U6898 (N_6898,N_6027,N_6279);
or U6899 (N_6899,N_6236,N_6292);
nor U6900 (N_6900,N_6011,N_6067);
and U6901 (N_6901,N_6310,N_6269);
and U6902 (N_6902,N_6048,N_6112);
nor U6903 (N_6903,N_6415,N_6337);
and U6904 (N_6904,N_6076,N_6373);
and U6905 (N_6905,N_6327,N_6126);
nor U6906 (N_6906,N_6300,N_6095);
or U6907 (N_6907,N_6424,N_6328);
and U6908 (N_6908,N_6412,N_6465);
xor U6909 (N_6909,N_6023,N_6146);
nand U6910 (N_6910,N_6486,N_6434);
or U6911 (N_6911,N_6091,N_6234);
nand U6912 (N_6912,N_6379,N_6086);
nand U6913 (N_6913,N_6466,N_6355);
and U6914 (N_6914,N_6112,N_6354);
and U6915 (N_6915,N_6085,N_6026);
or U6916 (N_6916,N_6063,N_6228);
nor U6917 (N_6917,N_6270,N_6118);
nand U6918 (N_6918,N_6183,N_6407);
nor U6919 (N_6919,N_6380,N_6182);
nand U6920 (N_6920,N_6263,N_6403);
nor U6921 (N_6921,N_6090,N_6353);
or U6922 (N_6922,N_6297,N_6403);
and U6923 (N_6923,N_6113,N_6479);
nand U6924 (N_6924,N_6423,N_6050);
nand U6925 (N_6925,N_6214,N_6429);
nor U6926 (N_6926,N_6285,N_6152);
nor U6927 (N_6927,N_6099,N_6142);
nor U6928 (N_6928,N_6222,N_6046);
or U6929 (N_6929,N_6078,N_6034);
and U6930 (N_6930,N_6373,N_6254);
nand U6931 (N_6931,N_6239,N_6144);
nand U6932 (N_6932,N_6147,N_6215);
nand U6933 (N_6933,N_6411,N_6275);
nor U6934 (N_6934,N_6225,N_6029);
and U6935 (N_6935,N_6344,N_6272);
nand U6936 (N_6936,N_6074,N_6188);
nor U6937 (N_6937,N_6272,N_6395);
and U6938 (N_6938,N_6362,N_6246);
nand U6939 (N_6939,N_6343,N_6063);
or U6940 (N_6940,N_6382,N_6440);
or U6941 (N_6941,N_6262,N_6086);
xnor U6942 (N_6942,N_6044,N_6160);
nor U6943 (N_6943,N_6253,N_6275);
and U6944 (N_6944,N_6347,N_6265);
nor U6945 (N_6945,N_6097,N_6147);
nand U6946 (N_6946,N_6010,N_6172);
nand U6947 (N_6947,N_6325,N_6334);
or U6948 (N_6948,N_6270,N_6212);
or U6949 (N_6949,N_6012,N_6380);
nand U6950 (N_6950,N_6243,N_6452);
nor U6951 (N_6951,N_6463,N_6206);
nor U6952 (N_6952,N_6470,N_6230);
and U6953 (N_6953,N_6025,N_6323);
nand U6954 (N_6954,N_6126,N_6259);
and U6955 (N_6955,N_6100,N_6234);
or U6956 (N_6956,N_6285,N_6031);
or U6957 (N_6957,N_6139,N_6277);
nor U6958 (N_6958,N_6396,N_6434);
nor U6959 (N_6959,N_6314,N_6249);
or U6960 (N_6960,N_6313,N_6418);
nand U6961 (N_6961,N_6375,N_6165);
and U6962 (N_6962,N_6145,N_6159);
or U6963 (N_6963,N_6424,N_6163);
or U6964 (N_6964,N_6494,N_6303);
or U6965 (N_6965,N_6103,N_6146);
or U6966 (N_6966,N_6070,N_6385);
xnor U6967 (N_6967,N_6351,N_6320);
nor U6968 (N_6968,N_6300,N_6431);
nand U6969 (N_6969,N_6286,N_6321);
nor U6970 (N_6970,N_6464,N_6397);
and U6971 (N_6971,N_6439,N_6117);
nand U6972 (N_6972,N_6217,N_6347);
xnor U6973 (N_6973,N_6458,N_6148);
or U6974 (N_6974,N_6146,N_6282);
or U6975 (N_6975,N_6014,N_6082);
nor U6976 (N_6976,N_6270,N_6159);
and U6977 (N_6977,N_6055,N_6117);
nor U6978 (N_6978,N_6286,N_6189);
or U6979 (N_6979,N_6039,N_6225);
xor U6980 (N_6980,N_6448,N_6061);
nor U6981 (N_6981,N_6329,N_6395);
or U6982 (N_6982,N_6015,N_6089);
nand U6983 (N_6983,N_6083,N_6100);
and U6984 (N_6984,N_6460,N_6024);
and U6985 (N_6985,N_6137,N_6264);
and U6986 (N_6986,N_6289,N_6123);
and U6987 (N_6987,N_6001,N_6215);
and U6988 (N_6988,N_6366,N_6035);
or U6989 (N_6989,N_6097,N_6177);
nor U6990 (N_6990,N_6092,N_6271);
nand U6991 (N_6991,N_6040,N_6488);
or U6992 (N_6992,N_6029,N_6000);
or U6993 (N_6993,N_6320,N_6453);
and U6994 (N_6994,N_6065,N_6217);
and U6995 (N_6995,N_6261,N_6204);
and U6996 (N_6996,N_6052,N_6098);
and U6997 (N_6997,N_6045,N_6287);
or U6998 (N_6998,N_6253,N_6025);
nand U6999 (N_6999,N_6115,N_6362);
or U7000 (N_7000,N_6814,N_6801);
nand U7001 (N_7001,N_6768,N_6882);
nand U7002 (N_7002,N_6777,N_6592);
nand U7003 (N_7003,N_6857,N_6707);
and U7004 (N_7004,N_6754,N_6574);
or U7005 (N_7005,N_6719,N_6678);
nand U7006 (N_7006,N_6842,N_6909);
nor U7007 (N_7007,N_6552,N_6543);
and U7008 (N_7008,N_6674,N_6876);
nand U7009 (N_7009,N_6737,N_6630);
nor U7010 (N_7010,N_6721,N_6911);
or U7011 (N_7011,N_6900,N_6528);
nor U7012 (N_7012,N_6818,N_6583);
nand U7013 (N_7013,N_6783,N_6736);
or U7014 (N_7014,N_6729,N_6647);
and U7015 (N_7015,N_6710,N_6692);
and U7016 (N_7016,N_6699,N_6503);
or U7017 (N_7017,N_6603,N_6550);
and U7018 (N_7018,N_6709,N_6978);
nor U7019 (N_7019,N_6995,N_6970);
or U7020 (N_7020,N_6878,N_6686);
nand U7021 (N_7021,N_6659,N_6837);
nand U7022 (N_7022,N_6834,N_6501);
and U7023 (N_7023,N_6648,N_6936);
or U7024 (N_7024,N_6875,N_6943);
and U7025 (N_7025,N_6865,N_6852);
nand U7026 (N_7026,N_6607,N_6920);
nand U7027 (N_7027,N_6618,N_6750);
nor U7028 (N_7028,N_6535,N_6919);
nand U7029 (N_7029,N_6657,N_6964);
nand U7030 (N_7030,N_6652,N_6741);
nor U7031 (N_7031,N_6606,N_6530);
nor U7032 (N_7032,N_6944,N_6985);
or U7033 (N_7033,N_6661,N_6811);
or U7034 (N_7034,N_6585,N_6604);
nor U7035 (N_7035,N_6646,N_6788);
or U7036 (N_7036,N_6664,N_6724);
nor U7037 (N_7037,N_6689,N_6907);
or U7038 (N_7038,N_6713,N_6778);
and U7039 (N_7039,N_6605,N_6714);
nand U7040 (N_7040,N_6701,N_6525);
or U7041 (N_7041,N_6864,N_6720);
nor U7042 (N_7042,N_6725,N_6663);
nor U7043 (N_7043,N_6708,N_6620);
or U7044 (N_7044,N_6961,N_6690);
or U7045 (N_7045,N_6682,N_6787);
or U7046 (N_7046,N_6895,N_6655);
or U7047 (N_7047,N_6718,N_6639);
or U7048 (N_7048,N_6817,N_6803);
or U7049 (N_7049,N_6636,N_6982);
and U7050 (N_7050,N_6634,N_6960);
nor U7051 (N_7051,N_6749,N_6967);
nor U7052 (N_7052,N_6973,N_6739);
nand U7053 (N_7053,N_6835,N_6742);
nand U7054 (N_7054,N_6877,N_6623);
and U7055 (N_7055,N_6993,N_6669);
nand U7056 (N_7056,N_6587,N_6923);
and U7057 (N_7057,N_6770,N_6573);
nor U7058 (N_7058,N_6931,N_6560);
or U7059 (N_7059,N_6809,N_6601);
nand U7060 (N_7060,N_6904,N_6554);
nor U7061 (N_7061,N_6555,N_6633);
or U7062 (N_7062,N_6883,N_6522);
nand U7063 (N_7063,N_6846,N_6934);
and U7064 (N_7064,N_6597,N_6539);
nor U7065 (N_7065,N_6752,N_6916);
or U7066 (N_7066,N_6516,N_6793);
nor U7067 (N_7067,N_6640,N_6631);
and U7068 (N_7068,N_6772,N_6807);
and U7069 (N_7069,N_6975,N_6628);
and U7070 (N_7070,N_6764,N_6802);
or U7071 (N_7071,N_6565,N_6829);
nand U7072 (N_7072,N_6621,N_6513);
or U7073 (N_7073,N_6782,N_6612);
or U7074 (N_7074,N_6712,N_6775);
or U7075 (N_7075,N_6624,N_6509);
or U7076 (N_7076,N_6862,N_6962);
nand U7077 (N_7077,N_6722,N_6518);
nand U7078 (N_7078,N_6765,N_6951);
nor U7079 (N_7079,N_6937,N_6950);
nand U7080 (N_7080,N_6644,N_6885);
nand U7081 (N_7081,N_6515,N_6563);
nor U7082 (N_7082,N_6537,N_6558);
nand U7083 (N_7083,N_6897,N_6728);
nor U7084 (N_7084,N_6711,N_6918);
nor U7085 (N_7085,N_6589,N_6963);
or U7086 (N_7086,N_6523,N_6653);
nand U7087 (N_7087,N_6965,N_6823);
and U7088 (N_7088,N_6697,N_6533);
and U7089 (N_7089,N_6939,N_6832);
and U7090 (N_7090,N_6602,N_6824);
and U7091 (N_7091,N_6941,N_6654);
and U7092 (N_7092,N_6766,N_6517);
nor U7093 (N_7093,N_6688,N_6781);
nand U7094 (N_7094,N_6898,N_6969);
nand U7095 (N_7095,N_6820,N_6671);
nand U7096 (N_7096,N_6785,N_6507);
nor U7097 (N_7097,N_6726,N_6798);
or U7098 (N_7098,N_6512,N_6828);
and U7099 (N_7099,N_6784,N_6683);
nand U7100 (N_7100,N_6984,N_6886);
xor U7101 (N_7101,N_6700,N_6567);
and U7102 (N_7102,N_6616,N_6795);
and U7103 (N_7103,N_6760,N_6696);
nand U7104 (N_7104,N_6847,N_6800);
nor U7105 (N_7105,N_6608,N_6979);
or U7106 (N_7106,N_6974,N_6925);
and U7107 (N_7107,N_6761,N_6703);
or U7108 (N_7108,N_6933,N_6727);
nand U7109 (N_7109,N_6773,N_6839);
or U7110 (N_7110,N_6954,N_6921);
nor U7111 (N_7111,N_6945,N_6680);
nor U7112 (N_7112,N_6861,N_6556);
nor U7113 (N_7113,N_6792,N_6698);
or U7114 (N_7114,N_6559,N_6850);
or U7115 (N_7115,N_6745,N_6526);
and U7116 (N_7116,N_6805,N_6968);
nor U7117 (N_7117,N_6893,N_6600);
nor U7118 (N_7118,N_6856,N_6996);
nand U7119 (N_7119,N_6681,N_6940);
and U7120 (N_7120,N_6626,N_6586);
or U7121 (N_7121,N_6966,N_6716);
and U7122 (N_7122,N_6870,N_6922);
or U7123 (N_7123,N_6582,N_6638);
nor U7124 (N_7124,N_6929,N_6987);
nand U7125 (N_7125,N_6956,N_6695);
nor U7126 (N_7126,N_6740,N_6858);
and U7127 (N_7127,N_6524,N_6572);
or U7128 (N_7128,N_6908,N_6905);
or U7129 (N_7129,N_6685,N_6562);
nand U7130 (N_7130,N_6953,N_6992);
or U7131 (N_7131,N_6930,N_6958);
nor U7132 (N_7132,N_6632,N_6771);
and U7133 (N_7133,N_6570,N_6762);
and U7134 (N_7134,N_6527,N_6851);
and U7135 (N_7135,N_6677,N_6825);
nand U7136 (N_7136,N_6545,N_6627);
or U7137 (N_7137,N_6853,N_6510);
nor U7138 (N_7138,N_6806,N_6650);
nand U7139 (N_7139,N_6948,N_6926);
and U7140 (N_7140,N_6816,N_6836);
or U7141 (N_7141,N_6549,N_6693);
and U7142 (N_7142,N_6860,N_6917);
or U7143 (N_7143,N_6981,N_6881);
xor U7144 (N_7144,N_6880,N_6548);
or U7145 (N_7145,N_6849,N_6946);
or U7146 (N_7146,N_6643,N_6578);
nand U7147 (N_7147,N_6957,N_6879);
nor U7148 (N_7148,N_6769,N_6924);
or U7149 (N_7149,N_6577,N_6841);
or U7150 (N_7150,N_6889,N_6675);
nand U7151 (N_7151,N_6821,N_6542);
nand U7152 (N_7152,N_6774,N_6547);
nor U7153 (N_7153,N_6635,N_6932);
or U7154 (N_7154,N_6611,N_6983);
or U7155 (N_7155,N_6734,N_6999);
xnor U7156 (N_7156,N_6658,N_6896);
or U7157 (N_7157,N_6927,N_6872);
nand U7158 (N_7158,N_6759,N_6668);
nor U7159 (N_7159,N_6593,N_6833);
or U7160 (N_7160,N_6913,N_6912);
or U7161 (N_7161,N_6986,N_6753);
nand U7162 (N_7162,N_6947,N_6591);
nor U7163 (N_7163,N_6822,N_6609);
and U7164 (N_7164,N_6763,N_6799);
and U7165 (N_7165,N_6590,N_6551);
nor U7166 (N_7166,N_6901,N_6534);
and U7167 (N_7167,N_6990,N_6952);
and U7168 (N_7168,N_6536,N_6519);
nand U7169 (N_7169,N_6502,N_6564);
nand U7170 (N_7170,N_6887,N_6830);
or U7171 (N_7171,N_6579,N_6935);
nor U7172 (N_7172,N_6684,N_6972);
nand U7173 (N_7173,N_6906,N_6662);
and U7174 (N_7174,N_6815,N_6756);
or U7175 (N_7175,N_6672,N_6959);
and U7176 (N_7176,N_6910,N_6827);
nor U7177 (N_7177,N_6642,N_6637);
nand U7178 (N_7178,N_6831,N_6546);
nor U7179 (N_7179,N_6665,N_6767);
nand U7180 (N_7180,N_6744,N_6641);
and U7181 (N_7181,N_6949,N_6667);
or U7182 (N_7182,N_6531,N_6691);
nand U7183 (N_7183,N_6505,N_6666);
or U7184 (N_7184,N_6557,N_6625);
xnor U7185 (N_7185,N_6575,N_6670);
nand U7186 (N_7186,N_6796,N_6994);
or U7187 (N_7187,N_6676,N_6649);
nor U7188 (N_7188,N_6679,N_6888);
nand U7189 (N_7189,N_6514,N_6617);
or U7190 (N_7190,N_6894,N_6694);
or U7191 (N_7191,N_6645,N_6706);
nor U7192 (N_7192,N_6808,N_6873);
nor U7193 (N_7193,N_6891,N_6629);
or U7194 (N_7194,N_6704,N_6614);
nand U7195 (N_7195,N_6500,N_6673);
nor U7196 (N_7196,N_6863,N_6702);
nor U7197 (N_7197,N_6855,N_6902);
nor U7198 (N_7198,N_6687,N_6890);
or U7199 (N_7199,N_6568,N_6791);
xnor U7200 (N_7200,N_6871,N_6884);
and U7201 (N_7201,N_6529,N_6892);
or U7202 (N_7202,N_6776,N_6596);
nor U7203 (N_7203,N_6731,N_6779);
and U7204 (N_7204,N_6656,N_6976);
nand U7205 (N_7205,N_6854,N_6651);
or U7206 (N_7206,N_6595,N_6997);
or U7207 (N_7207,N_6928,N_6748);
and U7208 (N_7208,N_6598,N_6758);
xor U7209 (N_7209,N_6733,N_6743);
nand U7210 (N_7210,N_6723,N_6610);
or U7211 (N_7211,N_6843,N_6566);
nand U7212 (N_7212,N_6615,N_6903);
or U7213 (N_7213,N_6715,N_6826);
and U7214 (N_7214,N_6511,N_6867);
nor U7215 (N_7215,N_6732,N_6599);
and U7216 (N_7216,N_6506,N_6738);
nor U7217 (N_7217,N_6751,N_6594);
and U7218 (N_7218,N_6735,N_6804);
and U7219 (N_7219,N_6810,N_6532);
or U7220 (N_7220,N_6991,N_6540);
nor U7221 (N_7221,N_6859,N_6866);
nand U7222 (N_7222,N_6838,N_6914);
and U7223 (N_7223,N_6840,N_6869);
nor U7224 (N_7224,N_6786,N_6613);
nor U7225 (N_7225,N_6622,N_6553);
nor U7226 (N_7226,N_6746,N_6520);
nand U7227 (N_7227,N_6569,N_6789);
and U7228 (N_7228,N_6580,N_6584);
nand U7229 (N_7229,N_6757,N_6561);
and U7230 (N_7230,N_6571,N_6989);
nand U7231 (N_7231,N_6915,N_6508);
nor U7232 (N_7232,N_6730,N_6521);
or U7233 (N_7233,N_6942,N_6797);
nor U7234 (N_7234,N_6938,N_6504);
or U7235 (N_7235,N_6977,N_6790);
or U7236 (N_7236,N_6844,N_6980);
nand U7237 (N_7237,N_6588,N_6812);
nor U7238 (N_7238,N_6541,N_6619);
nand U7239 (N_7239,N_6899,N_6538);
or U7240 (N_7240,N_6813,N_6780);
nand U7241 (N_7241,N_6998,N_6660);
and U7242 (N_7242,N_6581,N_6845);
and U7243 (N_7243,N_6988,N_6747);
and U7244 (N_7244,N_6717,N_6848);
or U7245 (N_7245,N_6874,N_6794);
nand U7246 (N_7246,N_6971,N_6576);
nand U7247 (N_7247,N_6544,N_6705);
or U7248 (N_7248,N_6868,N_6819);
or U7249 (N_7249,N_6955,N_6755);
nand U7250 (N_7250,N_6895,N_6731);
or U7251 (N_7251,N_6763,N_6533);
nor U7252 (N_7252,N_6684,N_6822);
nor U7253 (N_7253,N_6710,N_6711);
nand U7254 (N_7254,N_6956,N_6570);
and U7255 (N_7255,N_6567,N_6841);
nor U7256 (N_7256,N_6564,N_6621);
nor U7257 (N_7257,N_6548,N_6806);
or U7258 (N_7258,N_6978,N_6727);
nor U7259 (N_7259,N_6530,N_6677);
nor U7260 (N_7260,N_6572,N_6819);
and U7261 (N_7261,N_6719,N_6868);
and U7262 (N_7262,N_6777,N_6675);
and U7263 (N_7263,N_6991,N_6627);
or U7264 (N_7264,N_6713,N_6901);
and U7265 (N_7265,N_6976,N_6731);
nand U7266 (N_7266,N_6903,N_6587);
nor U7267 (N_7267,N_6603,N_6548);
nor U7268 (N_7268,N_6945,N_6872);
nor U7269 (N_7269,N_6661,N_6707);
or U7270 (N_7270,N_6940,N_6628);
and U7271 (N_7271,N_6961,N_6919);
nor U7272 (N_7272,N_6764,N_6693);
nor U7273 (N_7273,N_6978,N_6746);
nor U7274 (N_7274,N_6671,N_6573);
and U7275 (N_7275,N_6890,N_6999);
nor U7276 (N_7276,N_6827,N_6580);
or U7277 (N_7277,N_6592,N_6622);
nand U7278 (N_7278,N_6984,N_6824);
or U7279 (N_7279,N_6628,N_6989);
or U7280 (N_7280,N_6520,N_6961);
xnor U7281 (N_7281,N_6675,N_6697);
nand U7282 (N_7282,N_6577,N_6811);
nor U7283 (N_7283,N_6723,N_6546);
or U7284 (N_7284,N_6635,N_6961);
nor U7285 (N_7285,N_6718,N_6873);
nor U7286 (N_7286,N_6732,N_6881);
nor U7287 (N_7287,N_6836,N_6541);
and U7288 (N_7288,N_6814,N_6758);
nor U7289 (N_7289,N_6928,N_6877);
nor U7290 (N_7290,N_6513,N_6724);
xnor U7291 (N_7291,N_6552,N_6853);
nand U7292 (N_7292,N_6759,N_6604);
nor U7293 (N_7293,N_6791,N_6973);
or U7294 (N_7294,N_6620,N_6658);
nor U7295 (N_7295,N_6793,N_6970);
and U7296 (N_7296,N_6524,N_6762);
and U7297 (N_7297,N_6848,N_6823);
and U7298 (N_7298,N_6708,N_6883);
nor U7299 (N_7299,N_6514,N_6903);
or U7300 (N_7300,N_6763,N_6735);
nand U7301 (N_7301,N_6817,N_6642);
nand U7302 (N_7302,N_6809,N_6659);
or U7303 (N_7303,N_6619,N_6646);
or U7304 (N_7304,N_6754,N_6705);
nand U7305 (N_7305,N_6816,N_6987);
nor U7306 (N_7306,N_6855,N_6979);
nand U7307 (N_7307,N_6586,N_6754);
nand U7308 (N_7308,N_6920,N_6979);
nand U7309 (N_7309,N_6926,N_6947);
nor U7310 (N_7310,N_6783,N_6905);
and U7311 (N_7311,N_6503,N_6632);
xnor U7312 (N_7312,N_6989,N_6738);
and U7313 (N_7313,N_6849,N_6745);
and U7314 (N_7314,N_6657,N_6578);
nand U7315 (N_7315,N_6580,N_6751);
or U7316 (N_7316,N_6664,N_6739);
or U7317 (N_7317,N_6511,N_6844);
or U7318 (N_7318,N_6848,N_6960);
xor U7319 (N_7319,N_6545,N_6509);
nand U7320 (N_7320,N_6712,N_6527);
xor U7321 (N_7321,N_6975,N_6734);
nor U7322 (N_7322,N_6697,N_6643);
or U7323 (N_7323,N_6985,N_6901);
nor U7324 (N_7324,N_6793,N_6929);
nand U7325 (N_7325,N_6668,N_6981);
nor U7326 (N_7326,N_6685,N_6544);
nand U7327 (N_7327,N_6540,N_6677);
or U7328 (N_7328,N_6662,N_6690);
and U7329 (N_7329,N_6837,N_6858);
or U7330 (N_7330,N_6863,N_6864);
nor U7331 (N_7331,N_6810,N_6948);
nand U7332 (N_7332,N_6663,N_6677);
nand U7333 (N_7333,N_6988,N_6942);
and U7334 (N_7334,N_6788,N_6715);
and U7335 (N_7335,N_6854,N_6540);
nor U7336 (N_7336,N_6839,N_6997);
and U7337 (N_7337,N_6774,N_6627);
or U7338 (N_7338,N_6983,N_6947);
nand U7339 (N_7339,N_6899,N_6548);
nand U7340 (N_7340,N_6588,N_6852);
or U7341 (N_7341,N_6638,N_6674);
or U7342 (N_7342,N_6624,N_6913);
or U7343 (N_7343,N_6723,N_6701);
nor U7344 (N_7344,N_6616,N_6510);
and U7345 (N_7345,N_6575,N_6910);
nor U7346 (N_7346,N_6754,N_6693);
and U7347 (N_7347,N_6602,N_6801);
nor U7348 (N_7348,N_6981,N_6987);
nor U7349 (N_7349,N_6562,N_6869);
or U7350 (N_7350,N_6890,N_6725);
or U7351 (N_7351,N_6855,N_6878);
nand U7352 (N_7352,N_6540,N_6707);
nand U7353 (N_7353,N_6607,N_6523);
or U7354 (N_7354,N_6622,N_6880);
and U7355 (N_7355,N_6966,N_6928);
nand U7356 (N_7356,N_6835,N_6645);
nand U7357 (N_7357,N_6696,N_6826);
or U7358 (N_7358,N_6769,N_6667);
or U7359 (N_7359,N_6764,N_6699);
and U7360 (N_7360,N_6846,N_6542);
or U7361 (N_7361,N_6700,N_6828);
and U7362 (N_7362,N_6937,N_6905);
nor U7363 (N_7363,N_6699,N_6981);
nor U7364 (N_7364,N_6565,N_6535);
nand U7365 (N_7365,N_6845,N_6811);
and U7366 (N_7366,N_6550,N_6791);
or U7367 (N_7367,N_6985,N_6896);
or U7368 (N_7368,N_6902,N_6950);
or U7369 (N_7369,N_6870,N_6599);
and U7370 (N_7370,N_6712,N_6949);
nand U7371 (N_7371,N_6840,N_6929);
nor U7372 (N_7372,N_6769,N_6750);
or U7373 (N_7373,N_6790,N_6993);
nand U7374 (N_7374,N_6895,N_6624);
or U7375 (N_7375,N_6580,N_6811);
xnor U7376 (N_7376,N_6709,N_6879);
nand U7377 (N_7377,N_6695,N_6705);
nor U7378 (N_7378,N_6669,N_6931);
or U7379 (N_7379,N_6515,N_6603);
nor U7380 (N_7380,N_6623,N_6727);
or U7381 (N_7381,N_6718,N_6517);
nand U7382 (N_7382,N_6528,N_6821);
xor U7383 (N_7383,N_6848,N_6838);
or U7384 (N_7384,N_6604,N_6620);
nor U7385 (N_7385,N_6536,N_6793);
or U7386 (N_7386,N_6738,N_6833);
or U7387 (N_7387,N_6834,N_6763);
nor U7388 (N_7388,N_6885,N_6563);
nor U7389 (N_7389,N_6937,N_6731);
nand U7390 (N_7390,N_6790,N_6659);
nand U7391 (N_7391,N_6531,N_6778);
xor U7392 (N_7392,N_6920,N_6853);
or U7393 (N_7393,N_6714,N_6501);
or U7394 (N_7394,N_6650,N_6879);
or U7395 (N_7395,N_6837,N_6937);
xor U7396 (N_7396,N_6916,N_6982);
or U7397 (N_7397,N_6896,N_6510);
and U7398 (N_7398,N_6761,N_6975);
and U7399 (N_7399,N_6970,N_6786);
xor U7400 (N_7400,N_6634,N_6542);
and U7401 (N_7401,N_6890,N_6921);
xnor U7402 (N_7402,N_6640,N_6626);
and U7403 (N_7403,N_6815,N_6754);
nor U7404 (N_7404,N_6964,N_6690);
or U7405 (N_7405,N_6908,N_6577);
or U7406 (N_7406,N_6636,N_6705);
or U7407 (N_7407,N_6815,N_6504);
nor U7408 (N_7408,N_6942,N_6695);
nor U7409 (N_7409,N_6950,N_6525);
nor U7410 (N_7410,N_6747,N_6813);
nor U7411 (N_7411,N_6535,N_6668);
nand U7412 (N_7412,N_6973,N_6622);
nand U7413 (N_7413,N_6960,N_6833);
nand U7414 (N_7414,N_6913,N_6657);
nand U7415 (N_7415,N_6673,N_6695);
or U7416 (N_7416,N_6630,N_6957);
or U7417 (N_7417,N_6777,N_6557);
or U7418 (N_7418,N_6886,N_6897);
or U7419 (N_7419,N_6681,N_6744);
nor U7420 (N_7420,N_6896,N_6748);
nor U7421 (N_7421,N_6901,N_6604);
and U7422 (N_7422,N_6733,N_6669);
or U7423 (N_7423,N_6539,N_6789);
nand U7424 (N_7424,N_6929,N_6994);
or U7425 (N_7425,N_6948,N_6943);
nand U7426 (N_7426,N_6791,N_6740);
xor U7427 (N_7427,N_6999,N_6529);
nand U7428 (N_7428,N_6744,N_6833);
and U7429 (N_7429,N_6528,N_6983);
or U7430 (N_7430,N_6916,N_6883);
nand U7431 (N_7431,N_6724,N_6786);
or U7432 (N_7432,N_6699,N_6589);
nand U7433 (N_7433,N_6589,N_6733);
nand U7434 (N_7434,N_6927,N_6610);
or U7435 (N_7435,N_6725,N_6685);
nand U7436 (N_7436,N_6608,N_6840);
nand U7437 (N_7437,N_6951,N_6586);
nor U7438 (N_7438,N_6693,N_6932);
nand U7439 (N_7439,N_6545,N_6658);
and U7440 (N_7440,N_6607,N_6956);
and U7441 (N_7441,N_6548,N_6656);
or U7442 (N_7442,N_6768,N_6930);
nor U7443 (N_7443,N_6668,N_6661);
nand U7444 (N_7444,N_6709,N_6873);
nor U7445 (N_7445,N_6811,N_6558);
and U7446 (N_7446,N_6681,N_6844);
nor U7447 (N_7447,N_6973,N_6679);
nor U7448 (N_7448,N_6576,N_6718);
nand U7449 (N_7449,N_6810,N_6572);
and U7450 (N_7450,N_6975,N_6657);
or U7451 (N_7451,N_6507,N_6829);
xor U7452 (N_7452,N_6928,N_6638);
and U7453 (N_7453,N_6831,N_6734);
and U7454 (N_7454,N_6573,N_6814);
nor U7455 (N_7455,N_6926,N_6542);
nand U7456 (N_7456,N_6895,N_6973);
nor U7457 (N_7457,N_6875,N_6916);
nor U7458 (N_7458,N_6671,N_6775);
nor U7459 (N_7459,N_6641,N_6839);
and U7460 (N_7460,N_6882,N_6994);
nand U7461 (N_7461,N_6713,N_6772);
nand U7462 (N_7462,N_6884,N_6683);
nor U7463 (N_7463,N_6739,N_6659);
nor U7464 (N_7464,N_6865,N_6656);
nor U7465 (N_7465,N_6757,N_6784);
nand U7466 (N_7466,N_6799,N_6891);
or U7467 (N_7467,N_6947,N_6795);
xnor U7468 (N_7468,N_6947,N_6869);
and U7469 (N_7469,N_6782,N_6739);
and U7470 (N_7470,N_6667,N_6755);
nand U7471 (N_7471,N_6834,N_6596);
nor U7472 (N_7472,N_6637,N_6817);
nand U7473 (N_7473,N_6856,N_6900);
nand U7474 (N_7474,N_6913,N_6835);
nor U7475 (N_7475,N_6669,N_6920);
or U7476 (N_7476,N_6537,N_6944);
and U7477 (N_7477,N_6591,N_6716);
nor U7478 (N_7478,N_6944,N_6615);
nand U7479 (N_7479,N_6930,N_6642);
or U7480 (N_7480,N_6856,N_6994);
and U7481 (N_7481,N_6828,N_6881);
nand U7482 (N_7482,N_6930,N_6723);
or U7483 (N_7483,N_6725,N_6965);
and U7484 (N_7484,N_6583,N_6761);
or U7485 (N_7485,N_6668,N_6909);
nor U7486 (N_7486,N_6602,N_6654);
nor U7487 (N_7487,N_6867,N_6576);
or U7488 (N_7488,N_6775,N_6861);
nand U7489 (N_7489,N_6689,N_6811);
and U7490 (N_7490,N_6800,N_6676);
and U7491 (N_7491,N_6754,N_6666);
or U7492 (N_7492,N_6767,N_6960);
xnor U7493 (N_7493,N_6611,N_6942);
nor U7494 (N_7494,N_6571,N_6713);
or U7495 (N_7495,N_6589,N_6606);
nand U7496 (N_7496,N_6844,N_6778);
nand U7497 (N_7497,N_6954,N_6555);
and U7498 (N_7498,N_6614,N_6609);
nor U7499 (N_7499,N_6599,N_6942);
xnor U7500 (N_7500,N_7130,N_7225);
nand U7501 (N_7501,N_7230,N_7101);
nand U7502 (N_7502,N_7194,N_7308);
and U7503 (N_7503,N_7413,N_7298);
and U7504 (N_7504,N_7009,N_7155);
or U7505 (N_7505,N_7336,N_7113);
xor U7506 (N_7506,N_7364,N_7421);
or U7507 (N_7507,N_7258,N_7076);
xor U7508 (N_7508,N_7482,N_7006);
nand U7509 (N_7509,N_7081,N_7313);
nor U7510 (N_7510,N_7071,N_7349);
nand U7511 (N_7511,N_7247,N_7165);
nor U7512 (N_7512,N_7468,N_7399);
nor U7513 (N_7513,N_7223,N_7379);
nor U7514 (N_7514,N_7167,N_7255);
nand U7515 (N_7515,N_7237,N_7064);
nand U7516 (N_7516,N_7418,N_7034);
nand U7517 (N_7517,N_7220,N_7050);
or U7518 (N_7518,N_7493,N_7361);
and U7519 (N_7519,N_7036,N_7047);
nand U7520 (N_7520,N_7376,N_7024);
or U7521 (N_7521,N_7330,N_7262);
or U7522 (N_7522,N_7461,N_7254);
nor U7523 (N_7523,N_7185,N_7429);
or U7524 (N_7524,N_7248,N_7492);
nor U7525 (N_7525,N_7335,N_7256);
or U7526 (N_7526,N_7234,N_7285);
and U7527 (N_7527,N_7021,N_7069);
or U7528 (N_7528,N_7326,N_7344);
nand U7529 (N_7529,N_7297,N_7372);
nor U7530 (N_7530,N_7388,N_7156);
nand U7531 (N_7531,N_7083,N_7133);
nor U7532 (N_7532,N_7019,N_7191);
or U7533 (N_7533,N_7368,N_7187);
nor U7534 (N_7534,N_7434,N_7206);
and U7535 (N_7535,N_7480,N_7366);
and U7536 (N_7536,N_7450,N_7169);
or U7537 (N_7537,N_7268,N_7014);
xor U7538 (N_7538,N_7420,N_7168);
and U7539 (N_7539,N_7246,N_7102);
and U7540 (N_7540,N_7271,N_7467);
nand U7541 (N_7541,N_7057,N_7031);
nand U7542 (N_7542,N_7337,N_7222);
nand U7543 (N_7543,N_7438,N_7445);
nor U7544 (N_7544,N_7452,N_7079);
nand U7545 (N_7545,N_7091,N_7098);
and U7546 (N_7546,N_7407,N_7403);
nand U7547 (N_7547,N_7389,N_7043);
and U7548 (N_7548,N_7498,N_7320);
or U7549 (N_7549,N_7177,N_7158);
nor U7550 (N_7550,N_7245,N_7317);
nor U7551 (N_7551,N_7454,N_7477);
and U7552 (N_7552,N_7040,N_7475);
nor U7553 (N_7553,N_7373,N_7088);
nor U7554 (N_7554,N_7182,N_7189);
nor U7555 (N_7555,N_7375,N_7201);
nand U7556 (N_7556,N_7427,N_7473);
nor U7557 (N_7557,N_7260,N_7026);
and U7558 (N_7558,N_7382,N_7179);
nand U7559 (N_7559,N_7353,N_7145);
or U7560 (N_7560,N_7488,N_7431);
nand U7561 (N_7561,N_7294,N_7061);
and U7562 (N_7562,N_7097,N_7152);
nand U7563 (N_7563,N_7491,N_7453);
nand U7564 (N_7564,N_7345,N_7018);
nand U7565 (N_7565,N_7395,N_7065);
nor U7566 (N_7566,N_7045,N_7470);
or U7567 (N_7567,N_7111,N_7448);
or U7568 (N_7568,N_7282,N_7086);
nor U7569 (N_7569,N_7243,N_7471);
and U7570 (N_7570,N_7135,N_7154);
nor U7571 (N_7571,N_7261,N_7134);
and U7572 (N_7572,N_7304,N_7020);
nand U7573 (N_7573,N_7137,N_7440);
nand U7574 (N_7574,N_7417,N_7249);
and U7575 (N_7575,N_7439,N_7163);
nor U7576 (N_7576,N_7153,N_7046);
nor U7577 (N_7577,N_7310,N_7324);
nor U7578 (N_7578,N_7385,N_7339);
or U7579 (N_7579,N_7178,N_7289);
nand U7580 (N_7580,N_7224,N_7227);
or U7581 (N_7581,N_7303,N_7028);
nand U7582 (N_7582,N_7105,N_7210);
or U7583 (N_7583,N_7402,N_7193);
nor U7584 (N_7584,N_7184,N_7327);
xor U7585 (N_7585,N_7404,N_7212);
and U7586 (N_7586,N_7497,N_7307);
nand U7587 (N_7587,N_7240,N_7226);
nand U7588 (N_7588,N_7002,N_7486);
nor U7589 (N_7589,N_7038,N_7484);
or U7590 (N_7590,N_7096,N_7430);
nor U7591 (N_7591,N_7350,N_7048);
and U7592 (N_7592,N_7348,N_7338);
nand U7593 (N_7593,N_7116,N_7296);
or U7594 (N_7594,N_7235,N_7478);
nand U7595 (N_7595,N_7406,N_7494);
nand U7596 (N_7596,N_7358,N_7013);
or U7597 (N_7597,N_7216,N_7322);
or U7598 (N_7598,N_7263,N_7284);
or U7599 (N_7599,N_7272,N_7059);
or U7600 (N_7600,N_7029,N_7401);
nand U7601 (N_7601,N_7392,N_7144);
and U7602 (N_7602,N_7011,N_7411);
or U7603 (N_7603,N_7356,N_7054);
and U7604 (N_7604,N_7360,N_7170);
or U7605 (N_7605,N_7472,N_7332);
xor U7606 (N_7606,N_7090,N_7044);
xor U7607 (N_7607,N_7299,N_7215);
or U7608 (N_7608,N_7208,N_7328);
nor U7609 (N_7609,N_7100,N_7426);
and U7610 (N_7610,N_7200,N_7396);
and U7611 (N_7611,N_7490,N_7140);
or U7612 (N_7612,N_7008,N_7139);
and U7613 (N_7613,N_7123,N_7037);
or U7614 (N_7614,N_7085,N_7242);
or U7615 (N_7615,N_7386,N_7387);
and U7616 (N_7616,N_7481,N_7425);
nand U7617 (N_7617,N_7384,N_7073);
nor U7618 (N_7618,N_7005,N_7093);
and U7619 (N_7619,N_7355,N_7039);
nor U7620 (N_7620,N_7213,N_7455);
nor U7621 (N_7621,N_7391,N_7127);
or U7622 (N_7622,N_7241,N_7365);
nor U7623 (N_7623,N_7084,N_7280);
or U7624 (N_7624,N_7124,N_7414);
and U7625 (N_7625,N_7067,N_7423);
nand U7626 (N_7626,N_7264,N_7007);
nor U7627 (N_7627,N_7499,N_7003);
nor U7628 (N_7628,N_7197,N_7346);
or U7629 (N_7629,N_7070,N_7056);
nand U7630 (N_7630,N_7228,N_7080);
nand U7631 (N_7631,N_7314,N_7078);
nor U7632 (N_7632,N_7265,N_7267);
or U7633 (N_7633,N_7437,N_7283);
nor U7634 (N_7634,N_7231,N_7292);
and U7635 (N_7635,N_7412,N_7341);
and U7636 (N_7636,N_7012,N_7068);
or U7637 (N_7637,N_7305,N_7433);
or U7638 (N_7638,N_7394,N_7128);
and U7639 (N_7639,N_7117,N_7221);
nand U7640 (N_7640,N_7251,N_7118);
and U7641 (N_7641,N_7319,N_7175);
and U7642 (N_7642,N_7143,N_7072);
nand U7643 (N_7643,N_7259,N_7469);
nor U7644 (N_7644,N_7334,N_7362);
nand U7645 (N_7645,N_7172,N_7351);
nor U7646 (N_7646,N_7257,N_7016);
nor U7647 (N_7647,N_7035,N_7199);
or U7648 (N_7648,N_7390,N_7103);
nand U7649 (N_7649,N_7410,N_7383);
nand U7650 (N_7650,N_7015,N_7207);
nand U7651 (N_7651,N_7340,N_7219);
or U7652 (N_7652,N_7354,N_7457);
nor U7653 (N_7653,N_7465,N_7196);
nand U7654 (N_7654,N_7449,N_7075);
and U7655 (N_7655,N_7150,N_7082);
nor U7656 (N_7656,N_7087,N_7162);
nor U7657 (N_7657,N_7107,N_7363);
nand U7658 (N_7658,N_7458,N_7211);
and U7659 (N_7659,N_7001,N_7108);
nand U7660 (N_7660,N_7273,N_7301);
and U7661 (N_7661,N_7321,N_7278);
or U7662 (N_7662,N_7487,N_7424);
nor U7663 (N_7663,N_7146,N_7266);
or U7664 (N_7664,N_7325,N_7333);
nor U7665 (N_7665,N_7004,N_7342);
nor U7666 (N_7666,N_7371,N_7309);
or U7667 (N_7667,N_7432,N_7062);
nand U7668 (N_7668,N_7329,N_7112);
and U7669 (N_7669,N_7074,N_7126);
and U7670 (N_7670,N_7495,N_7459);
nor U7671 (N_7671,N_7466,N_7323);
nand U7672 (N_7672,N_7052,N_7122);
nor U7673 (N_7673,N_7214,N_7159);
and U7674 (N_7674,N_7239,N_7094);
nor U7675 (N_7675,N_7233,N_7274);
nand U7676 (N_7676,N_7496,N_7232);
nor U7677 (N_7677,N_7171,N_7218);
nor U7678 (N_7678,N_7288,N_7176);
nor U7679 (N_7679,N_7311,N_7446);
nor U7680 (N_7680,N_7370,N_7106);
nand U7681 (N_7681,N_7295,N_7483);
xor U7682 (N_7682,N_7109,N_7476);
or U7683 (N_7683,N_7205,N_7397);
nor U7684 (N_7684,N_7291,N_7447);
and U7685 (N_7685,N_7316,N_7464);
nand U7686 (N_7686,N_7136,N_7367);
nand U7687 (N_7687,N_7204,N_7023);
nand U7688 (N_7688,N_7164,N_7149);
xor U7689 (N_7689,N_7281,N_7151);
nand U7690 (N_7690,N_7489,N_7027);
nand U7691 (N_7691,N_7060,N_7374);
nand U7692 (N_7692,N_7422,N_7030);
or U7693 (N_7693,N_7236,N_7441);
xnor U7694 (N_7694,N_7408,N_7442);
or U7695 (N_7695,N_7017,N_7393);
and U7696 (N_7696,N_7238,N_7209);
xor U7697 (N_7697,N_7252,N_7275);
xnor U7698 (N_7698,N_7250,N_7066);
nand U7699 (N_7699,N_7217,N_7053);
nand U7700 (N_7700,N_7435,N_7331);
nand U7701 (N_7701,N_7095,N_7244);
nor U7702 (N_7702,N_7198,N_7049);
nor U7703 (N_7703,N_7293,N_7474);
or U7704 (N_7704,N_7192,N_7022);
nor U7705 (N_7705,N_7451,N_7110);
or U7706 (N_7706,N_7147,N_7033);
or U7707 (N_7707,N_7443,N_7479);
nand U7708 (N_7708,N_7099,N_7378);
nor U7709 (N_7709,N_7318,N_7058);
nand U7710 (N_7710,N_7312,N_7286);
and U7711 (N_7711,N_7114,N_7188);
and U7712 (N_7712,N_7398,N_7180);
or U7713 (N_7713,N_7302,N_7063);
or U7714 (N_7714,N_7269,N_7202);
xnor U7715 (N_7715,N_7148,N_7357);
and U7716 (N_7716,N_7462,N_7173);
nand U7717 (N_7717,N_7183,N_7306);
nor U7718 (N_7718,N_7120,N_7055);
or U7719 (N_7719,N_7300,N_7463);
nand U7720 (N_7720,N_7186,N_7077);
nand U7721 (N_7721,N_7419,N_7129);
or U7722 (N_7722,N_7025,N_7377);
and U7723 (N_7723,N_7119,N_7181);
and U7724 (N_7724,N_7138,N_7276);
nand U7725 (N_7725,N_7160,N_7253);
nand U7726 (N_7726,N_7436,N_7157);
or U7727 (N_7727,N_7460,N_7400);
or U7728 (N_7728,N_7428,N_7041);
or U7729 (N_7729,N_7190,N_7161);
nor U7730 (N_7730,N_7115,N_7277);
nor U7731 (N_7731,N_7010,N_7166);
and U7732 (N_7732,N_7174,N_7092);
nand U7733 (N_7733,N_7287,N_7444);
or U7734 (N_7734,N_7089,N_7290);
nand U7735 (N_7735,N_7195,N_7132);
nand U7736 (N_7736,N_7416,N_7369);
nor U7737 (N_7737,N_7104,N_7032);
and U7738 (N_7738,N_7359,N_7131);
or U7739 (N_7739,N_7456,N_7142);
nand U7740 (N_7740,N_7000,N_7279);
and U7741 (N_7741,N_7409,N_7315);
and U7742 (N_7742,N_7229,N_7343);
and U7743 (N_7743,N_7380,N_7121);
nand U7744 (N_7744,N_7381,N_7141);
or U7745 (N_7745,N_7347,N_7051);
nor U7746 (N_7746,N_7415,N_7042);
nand U7747 (N_7747,N_7203,N_7270);
nor U7748 (N_7748,N_7485,N_7352);
nand U7749 (N_7749,N_7125,N_7405);
nor U7750 (N_7750,N_7409,N_7435);
or U7751 (N_7751,N_7278,N_7009);
or U7752 (N_7752,N_7307,N_7470);
and U7753 (N_7753,N_7023,N_7047);
or U7754 (N_7754,N_7325,N_7291);
nand U7755 (N_7755,N_7040,N_7147);
and U7756 (N_7756,N_7060,N_7311);
or U7757 (N_7757,N_7137,N_7277);
nor U7758 (N_7758,N_7136,N_7346);
nand U7759 (N_7759,N_7332,N_7221);
nor U7760 (N_7760,N_7114,N_7135);
or U7761 (N_7761,N_7492,N_7001);
nor U7762 (N_7762,N_7031,N_7271);
and U7763 (N_7763,N_7109,N_7009);
nand U7764 (N_7764,N_7274,N_7131);
nand U7765 (N_7765,N_7202,N_7467);
or U7766 (N_7766,N_7404,N_7124);
xor U7767 (N_7767,N_7003,N_7151);
and U7768 (N_7768,N_7342,N_7306);
nor U7769 (N_7769,N_7080,N_7483);
nor U7770 (N_7770,N_7333,N_7301);
nand U7771 (N_7771,N_7045,N_7495);
nor U7772 (N_7772,N_7259,N_7376);
and U7773 (N_7773,N_7045,N_7336);
and U7774 (N_7774,N_7215,N_7472);
nand U7775 (N_7775,N_7482,N_7215);
nor U7776 (N_7776,N_7138,N_7091);
or U7777 (N_7777,N_7398,N_7478);
or U7778 (N_7778,N_7481,N_7276);
and U7779 (N_7779,N_7361,N_7487);
nor U7780 (N_7780,N_7065,N_7346);
nand U7781 (N_7781,N_7243,N_7311);
and U7782 (N_7782,N_7244,N_7021);
and U7783 (N_7783,N_7357,N_7365);
or U7784 (N_7784,N_7128,N_7355);
nand U7785 (N_7785,N_7376,N_7436);
nand U7786 (N_7786,N_7291,N_7056);
nor U7787 (N_7787,N_7084,N_7336);
nor U7788 (N_7788,N_7178,N_7347);
or U7789 (N_7789,N_7218,N_7483);
and U7790 (N_7790,N_7032,N_7246);
and U7791 (N_7791,N_7462,N_7499);
or U7792 (N_7792,N_7281,N_7089);
or U7793 (N_7793,N_7100,N_7026);
nor U7794 (N_7794,N_7488,N_7172);
nand U7795 (N_7795,N_7304,N_7478);
or U7796 (N_7796,N_7410,N_7152);
and U7797 (N_7797,N_7429,N_7225);
or U7798 (N_7798,N_7391,N_7196);
or U7799 (N_7799,N_7372,N_7200);
nor U7800 (N_7800,N_7468,N_7273);
and U7801 (N_7801,N_7389,N_7049);
nand U7802 (N_7802,N_7430,N_7137);
or U7803 (N_7803,N_7278,N_7065);
or U7804 (N_7804,N_7169,N_7017);
or U7805 (N_7805,N_7461,N_7089);
and U7806 (N_7806,N_7366,N_7410);
nor U7807 (N_7807,N_7393,N_7090);
and U7808 (N_7808,N_7377,N_7449);
and U7809 (N_7809,N_7247,N_7203);
nor U7810 (N_7810,N_7140,N_7161);
and U7811 (N_7811,N_7006,N_7353);
nor U7812 (N_7812,N_7118,N_7321);
nor U7813 (N_7813,N_7245,N_7063);
and U7814 (N_7814,N_7157,N_7042);
and U7815 (N_7815,N_7450,N_7191);
or U7816 (N_7816,N_7464,N_7298);
and U7817 (N_7817,N_7293,N_7114);
nand U7818 (N_7818,N_7104,N_7417);
or U7819 (N_7819,N_7471,N_7036);
nor U7820 (N_7820,N_7383,N_7266);
nor U7821 (N_7821,N_7260,N_7003);
nand U7822 (N_7822,N_7419,N_7060);
nand U7823 (N_7823,N_7008,N_7410);
or U7824 (N_7824,N_7220,N_7047);
nand U7825 (N_7825,N_7495,N_7348);
nor U7826 (N_7826,N_7140,N_7305);
nand U7827 (N_7827,N_7135,N_7190);
nand U7828 (N_7828,N_7269,N_7244);
nor U7829 (N_7829,N_7070,N_7281);
and U7830 (N_7830,N_7303,N_7087);
or U7831 (N_7831,N_7008,N_7144);
nor U7832 (N_7832,N_7180,N_7342);
and U7833 (N_7833,N_7459,N_7133);
and U7834 (N_7834,N_7116,N_7009);
nand U7835 (N_7835,N_7250,N_7436);
nor U7836 (N_7836,N_7018,N_7281);
xnor U7837 (N_7837,N_7224,N_7111);
and U7838 (N_7838,N_7232,N_7115);
and U7839 (N_7839,N_7131,N_7000);
nand U7840 (N_7840,N_7216,N_7180);
and U7841 (N_7841,N_7319,N_7273);
nand U7842 (N_7842,N_7009,N_7072);
nor U7843 (N_7843,N_7499,N_7038);
and U7844 (N_7844,N_7482,N_7446);
nor U7845 (N_7845,N_7096,N_7205);
and U7846 (N_7846,N_7396,N_7490);
or U7847 (N_7847,N_7183,N_7081);
or U7848 (N_7848,N_7301,N_7250);
nand U7849 (N_7849,N_7123,N_7249);
and U7850 (N_7850,N_7128,N_7180);
or U7851 (N_7851,N_7318,N_7056);
and U7852 (N_7852,N_7018,N_7088);
and U7853 (N_7853,N_7140,N_7495);
or U7854 (N_7854,N_7388,N_7115);
and U7855 (N_7855,N_7192,N_7129);
and U7856 (N_7856,N_7086,N_7109);
and U7857 (N_7857,N_7147,N_7298);
or U7858 (N_7858,N_7094,N_7284);
and U7859 (N_7859,N_7320,N_7315);
and U7860 (N_7860,N_7213,N_7472);
nor U7861 (N_7861,N_7310,N_7192);
nand U7862 (N_7862,N_7081,N_7291);
and U7863 (N_7863,N_7434,N_7481);
and U7864 (N_7864,N_7249,N_7491);
nand U7865 (N_7865,N_7017,N_7079);
or U7866 (N_7866,N_7195,N_7121);
nand U7867 (N_7867,N_7377,N_7320);
nand U7868 (N_7868,N_7295,N_7489);
or U7869 (N_7869,N_7473,N_7132);
or U7870 (N_7870,N_7100,N_7422);
or U7871 (N_7871,N_7112,N_7364);
or U7872 (N_7872,N_7017,N_7199);
xnor U7873 (N_7873,N_7401,N_7027);
or U7874 (N_7874,N_7174,N_7272);
nand U7875 (N_7875,N_7313,N_7102);
nand U7876 (N_7876,N_7235,N_7414);
and U7877 (N_7877,N_7020,N_7394);
and U7878 (N_7878,N_7059,N_7057);
nand U7879 (N_7879,N_7381,N_7256);
or U7880 (N_7880,N_7322,N_7457);
nor U7881 (N_7881,N_7239,N_7373);
or U7882 (N_7882,N_7356,N_7021);
and U7883 (N_7883,N_7406,N_7274);
nand U7884 (N_7884,N_7404,N_7221);
or U7885 (N_7885,N_7011,N_7032);
or U7886 (N_7886,N_7409,N_7305);
and U7887 (N_7887,N_7134,N_7254);
nand U7888 (N_7888,N_7206,N_7122);
nor U7889 (N_7889,N_7209,N_7229);
nor U7890 (N_7890,N_7015,N_7239);
nor U7891 (N_7891,N_7381,N_7124);
nand U7892 (N_7892,N_7403,N_7446);
nand U7893 (N_7893,N_7274,N_7186);
or U7894 (N_7894,N_7208,N_7350);
or U7895 (N_7895,N_7168,N_7326);
nor U7896 (N_7896,N_7283,N_7185);
and U7897 (N_7897,N_7207,N_7089);
or U7898 (N_7898,N_7322,N_7353);
and U7899 (N_7899,N_7439,N_7303);
and U7900 (N_7900,N_7186,N_7469);
and U7901 (N_7901,N_7383,N_7130);
nor U7902 (N_7902,N_7060,N_7112);
nor U7903 (N_7903,N_7301,N_7089);
or U7904 (N_7904,N_7472,N_7048);
and U7905 (N_7905,N_7196,N_7488);
or U7906 (N_7906,N_7486,N_7219);
nand U7907 (N_7907,N_7404,N_7494);
or U7908 (N_7908,N_7399,N_7350);
or U7909 (N_7909,N_7392,N_7297);
and U7910 (N_7910,N_7470,N_7419);
nand U7911 (N_7911,N_7084,N_7362);
nand U7912 (N_7912,N_7021,N_7314);
nor U7913 (N_7913,N_7408,N_7325);
and U7914 (N_7914,N_7321,N_7348);
or U7915 (N_7915,N_7429,N_7489);
nor U7916 (N_7916,N_7150,N_7291);
nor U7917 (N_7917,N_7130,N_7177);
or U7918 (N_7918,N_7202,N_7213);
nor U7919 (N_7919,N_7475,N_7141);
xor U7920 (N_7920,N_7346,N_7418);
nor U7921 (N_7921,N_7161,N_7254);
nor U7922 (N_7922,N_7156,N_7427);
and U7923 (N_7923,N_7092,N_7094);
nor U7924 (N_7924,N_7133,N_7422);
nor U7925 (N_7925,N_7417,N_7451);
nor U7926 (N_7926,N_7007,N_7144);
and U7927 (N_7927,N_7093,N_7236);
nor U7928 (N_7928,N_7372,N_7253);
nor U7929 (N_7929,N_7286,N_7413);
or U7930 (N_7930,N_7029,N_7343);
nand U7931 (N_7931,N_7126,N_7227);
and U7932 (N_7932,N_7120,N_7492);
or U7933 (N_7933,N_7055,N_7069);
nor U7934 (N_7934,N_7355,N_7410);
nand U7935 (N_7935,N_7091,N_7420);
nor U7936 (N_7936,N_7201,N_7193);
nand U7937 (N_7937,N_7091,N_7426);
or U7938 (N_7938,N_7170,N_7064);
and U7939 (N_7939,N_7195,N_7126);
xnor U7940 (N_7940,N_7430,N_7390);
nand U7941 (N_7941,N_7277,N_7075);
or U7942 (N_7942,N_7101,N_7458);
and U7943 (N_7943,N_7257,N_7276);
nand U7944 (N_7944,N_7008,N_7204);
and U7945 (N_7945,N_7122,N_7425);
nor U7946 (N_7946,N_7126,N_7326);
and U7947 (N_7947,N_7271,N_7382);
nand U7948 (N_7948,N_7300,N_7146);
nor U7949 (N_7949,N_7281,N_7175);
or U7950 (N_7950,N_7139,N_7078);
nor U7951 (N_7951,N_7065,N_7397);
nor U7952 (N_7952,N_7411,N_7178);
nor U7953 (N_7953,N_7187,N_7119);
or U7954 (N_7954,N_7046,N_7377);
nor U7955 (N_7955,N_7088,N_7238);
nand U7956 (N_7956,N_7303,N_7066);
xor U7957 (N_7957,N_7152,N_7322);
nand U7958 (N_7958,N_7032,N_7436);
nor U7959 (N_7959,N_7278,N_7453);
and U7960 (N_7960,N_7138,N_7158);
and U7961 (N_7961,N_7403,N_7202);
or U7962 (N_7962,N_7425,N_7044);
nand U7963 (N_7963,N_7421,N_7096);
or U7964 (N_7964,N_7470,N_7463);
nand U7965 (N_7965,N_7279,N_7184);
nor U7966 (N_7966,N_7464,N_7072);
nor U7967 (N_7967,N_7390,N_7494);
nand U7968 (N_7968,N_7430,N_7066);
and U7969 (N_7969,N_7393,N_7315);
or U7970 (N_7970,N_7263,N_7377);
and U7971 (N_7971,N_7389,N_7295);
nor U7972 (N_7972,N_7071,N_7140);
nor U7973 (N_7973,N_7452,N_7340);
nor U7974 (N_7974,N_7080,N_7286);
and U7975 (N_7975,N_7086,N_7022);
nor U7976 (N_7976,N_7449,N_7366);
and U7977 (N_7977,N_7157,N_7333);
nand U7978 (N_7978,N_7012,N_7223);
or U7979 (N_7979,N_7137,N_7158);
or U7980 (N_7980,N_7022,N_7085);
nor U7981 (N_7981,N_7157,N_7358);
and U7982 (N_7982,N_7415,N_7144);
and U7983 (N_7983,N_7247,N_7310);
nor U7984 (N_7984,N_7467,N_7486);
nand U7985 (N_7985,N_7093,N_7131);
nand U7986 (N_7986,N_7430,N_7068);
nor U7987 (N_7987,N_7186,N_7288);
and U7988 (N_7988,N_7266,N_7304);
nor U7989 (N_7989,N_7426,N_7101);
or U7990 (N_7990,N_7090,N_7269);
nand U7991 (N_7991,N_7198,N_7071);
nand U7992 (N_7992,N_7477,N_7104);
and U7993 (N_7993,N_7457,N_7386);
nand U7994 (N_7994,N_7448,N_7363);
or U7995 (N_7995,N_7075,N_7133);
or U7996 (N_7996,N_7320,N_7405);
xnor U7997 (N_7997,N_7043,N_7481);
or U7998 (N_7998,N_7178,N_7362);
nand U7999 (N_7999,N_7086,N_7285);
nor U8000 (N_8000,N_7642,N_7675);
or U8001 (N_8001,N_7985,N_7669);
xor U8002 (N_8002,N_7668,N_7592);
nand U8003 (N_8003,N_7628,N_7830);
and U8004 (N_8004,N_7562,N_7992);
and U8005 (N_8005,N_7800,N_7920);
nor U8006 (N_8006,N_7597,N_7833);
nor U8007 (N_8007,N_7853,N_7858);
nor U8008 (N_8008,N_7590,N_7620);
or U8009 (N_8009,N_7684,N_7703);
nand U8010 (N_8010,N_7740,N_7772);
nand U8011 (N_8011,N_7728,N_7661);
and U8012 (N_8012,N_7542,N_7673);
nor U8013 (N_8013,N_7569,N_7945);
nor U8014 (N_8014,N_7984,N_7877);
nand U8015 (N_8015,N_7901,N_7835);
xnor U8016 (N_8016,N_7730,N_7818);
and U8017 (N_8017,N_7852,N_7868);
nor U8018 (N_8018,N_7894,N_7911);
nor U8019 (N_8019,N_7618,N_7545);
or U8020 (N_8020,N_7790,N_7714);
and U8021 (N_8021,N_7507,N_7718);
or U8022 (N_8022,N_7954,N_7505);
or U8023 (N_8023,N_7902,N_7660);
nor U8024 (N_8024,N_7764,N_7948);
or U8025 (N_8025,N_7706,N_7797);
nor U8026 (N_8026,N_7587,N_7938);
or U8027 (N_8027,N_7515,N_7971);
xnor U8028 (N_8028,N_7688,N_7544);
nor U8029 (N_8029,N_7546,N_7994);
nor U8030 (N_8030,N_7957,N_7978);
nor U8031 (N_8031,N_7799,N_7863);
or U8032 (N_8032,N_7804,N_7605);
or U8033 (N_8033,N_7603,N_7834);
nor U8034 (N_8034,N_7696,N_7500);
xnor U8035 (N_8035,N_7904,N_7773);
nand U8036 (N_8036,N_7807,N_7870);
nor U8037 (N_8037,N_7925,N_7942);
nand U8038 (N_8038,N_7778,N_7591);
and U8039 (N_8039,N_7671,N_7980);
nor U8040 (N_8040,N_7792,N_7513);
nand U8041 (N_8041,N_7878,N_7855);
or U8042 (N_8042,N_7599,N_7916);
nor U8043 (N_8043,N_7653,N_7887);
nor U8044 (N_8044,N_7953,N_7727);
nand U8045 (N_8045,N_7708,N_7608);
xnor U8046 (N_8046,N_7848,N_7707);
nand U8047 (N_8047,N_7538,N_7930);
and U8048 (N_8048,N_7729,N_7625);
nor U8049 (N_8049,N_7556,N_7525);
nor U8050 (N_8050,N_7826,N_7865);
or U8051 (N_8051,N_7864,N_7931);
and U8052 (N_8052,N_7510,N_7548);
nand U8053 (N_8053,N_7717,N_7781);
nand U8054 (N_8054,N_7828,N_7667);
nor U8055 (N_8055,N_7988,N_7615);
nand U8056 (N_8056,N_7937,N_7838);
nand U8057 (N_8057,N_7851,N_7643);
nor U8058 (N_8058,N_7919,N_7960);
nand U8059 (N_8059,N_7511,N_7568);
or U8060 (N_8060,N_7629,N_7927);
nand U8061 (N_8061,N_7641,N_7640);
nor U8062 (N_8062,N_7777,N_7757);
and U8063 (N_8063,N_7572,N_7837);
or U8064 (N_8064,N_7898,N_7841);
nor U8065 (N_8065,N_7793,N_7810);
and U8066 (N_8066,N_7861,N_7540);
nand U8067 (N_8067,N_7829,N_7873);
nand U8068 (N_8068,N_7915,N_7979);
and U8069 (N_8069,N_7682,N_7533);
or U8070 (N_8070,N_7549,N_7600);
nor U8071 (N_8071,N_7914,N_7903);
nor U8072 (N_8072,N_7921,N_7748);
nor U8073 (N_8073,N_7593,N_7766);
nand U8074 (N_8074,N_7630,N_7683);
nand U8075 (N_8075,N_7687,N_7739);
nor U8076 (N_8076,N_7563,N_7601);
or U8077 (N_8077,N_7951,N_7967);
nand U8078 (N_8078,N_7633,N_7842);
nand U8079 (N_8079,N_7503,N_7553);
nand U8080 (N_8080,N_7731,N_7836);
and U8081 (N_8081,N_7832,N_7849);
nor U8082 (N_8082,N_7856,N_7987);
nand U8083 (N_8083,N_7716,N_7632);
nor U8084 (N_8084,N_7813,N_7536);
and U8085 (N_8085,N_7753,N_7885);
or U8086 (N_8086,N_7997,N_7962);
nand U8087 (N_8087,N_7588,N_7875);
and U8088 (N_8088,N_7963,N_7516);
and U8089 (N_8089,N_7932,N_7543);
xnor U8090 (N_8090,N_7528,N_7535);
nor U8091 (N_8091,N_7741,N_7690);
or U8092 (N_8092,N_7803,N_7644);
or U8093 (N_8093,N_7570,N_7974);
nor U8094 (N_8094,N_7524,N_7784);
and U8095 (N_8095,N_7762,N_7656);
nand U8096 (N_8096,N_7821,N_7843);
nand U8097 (N_8097,N_7733,N_7783);
and U8098 (N_8098,N_7808,N_7596);
nor U8099 (N_8099,N_7602,N_7941);
and U8100 (N_8100,N_7831,N_7977);
or U8101 (N_8101,N_7509,N_7635);
or U8102 (N_8102,N_7996,N_7647);
nor U8103 (N_8103,N_7558,N_7795);
or U8104 (N_8104,N_7820,N_7884);
nor U8105 (N_8105,N_7972,N_7964);
or U8106 (N_8106,N_7541,N_7787);
or U8107 (N_8107,N_7697,N_7754);
and U8108 (N_8108,N_7634,N_7889);
and U8109 (N_8109,N_7906,N_7521);
or U8110 (N_8110,N_7617,N_7585);
or U8111 (N_8111,N_7681,N_7664);
or U8112 (N_8112,N_7770,N_7504);
nand U8113 (N_8113,N_7622,N_7532);
nand U8114 (N_8114,N_7619,N_7639);
nand U8115 (N_8115,N_7665,N_7699);
or U8116 (N_8116,N_7638,N_7819);
or U8117 (N_8117,N_7710,N_7610);
or U8118 (N_8118,N_7575,N_7794);
nor U8119 (N_8119,N_7655,N_7659);
nor U8120 (N_8120,N_7825,N_7695);
and U8121 (N_8121,N_7958,N_7771);
and U8122 (N_8122,N_7709,N_7751);
nor U8123 (N_8123,N_7760,N_7614);
nand U8124 (N_8124,N_7947,N_7574);
and U8125 (N_8125,N_7900,N_7782);
and U8126 (N_8126,N_7726,N_7850);
or U8127 (N_8127,N_7908,N_7822);
and U8128 (N_8128,N_7583,N_7989);
nor U8129 (N_8129,N_7577,N_7943);
or U8130 (N_8130,N_7999,N_7518);
nor U8131 (N_8131,N_7779,N_7724);
nor U8132 (N_8132,N_7711,N_7694);
nand U8133 (N_8133,N_7567,N_7743);
nor U8134 (N_8134,N_7955,N_7926);
nand U8135 (N_8135,N_7522,N_7611);
nand U8136 (N_8136,N_7715,N_7859);
nor U8137 (N_8137,N_7721,N_7952);
nor U8138 (N_8138,N_7654,N_7559);
nand U8139 (N_8139,N_7879,N_7554);
and U8140 (N_8140,N_7775,N_7537);
nand U8141 (N_8141,N_7805,N_7720);
or U8142 (N_8142,N_7909,N_7589);
and U8143 (N_8143,N_7899,N_7531);
nor U8144 (N_8144,N_7670,N_7944);
nand U8145 (N_8145,N_7949,N_7514);
and U8146 (N_8146,N_7789,N_7975);
and U8147 (N_8147,N_7750,N_7674);
nand U8148 (N_8148,N_7680,N_7982);
and U8149 (N_8149,N_7689,N_7811);
nand U8150 (N_8150,N_7649,N_7840);
and U8151 (N_8151,N_7744,N_7986);
and U8152 (N_8152,N_7594,N_7888);
nand U8153 (N_8153,N_7929,N_7704);
and U8154 (N_8154,N_7939,N_7565);
nor U8155 (N_8155,N_7882,N_7579);
nand U8156 (N_8156,N_7785,N_7780);
nand U8157 (N_8157,N_7817,N_7891);
nand U8158 (N_8158,N_7876,N_7517);
nor U8159 (N_8159,N_7746,N_7648);
nor U8160 (N_8160,N_7658,N_7786);
nor U8161 (N_8161,N_7561,N_7923);
nor U8162 (N_8162,N_7626,N_7768);
and U8163 (N_8163,N_7998,N_7895);
nand U8164 (N_8164,N_7956,N_7530);
and U8165 (N_8165,N_7763,N_7935);
nand U8166 (N_8166,N_7607,N_7712);
nor U8167 (N_8167,N_7586,N_7892);
nor U8168 (N_8168,N_7886,N_7755);
or U8169 (N_8169,N_7823,N_7815);
and U8170 (N_8170,N_7961,N_7523);
nand U8171 (N_8171,N_7995,N_7651);
and U8172 (N_8172,N_7910,N_7736);
or U8173 (N_8173,N_7526,N_7950);
nand U8174 (N_8174,N_7646,N_7924);
or U8175 (N_8175,N_7564,N_7512);
nor U8176 (N_8176,N_7581,N_7765);
and U8177 (N_8177,N_7502,N_7501);
xnor U8178 (N_8178,N_7896,N_7839);
or U8179 (N_8179,N_7874,N_7918);
or U8180 (N_8180,N_7802,N_7552);
and U8181 (N_8181,N_7737,N_7759);
or U8182 (N_8182,N_7508,N_7806);
or U8183 (N_8183,N_7539,N_7970);
nand U8184 (N_8184,N_7613,N_7857);
or U8185 (N_8185,N_7637,N_7652);
nand U8186 (N_8186,N_7735,N_7860);
or U8187 (N_8187,N_7529,N_7907);
or U8188 (N_8188,N_7940,N_7871);
nor U8189 (N_8189,N_7854,N_7756);
nand U8190 (N_8190,N_7571,N_7598);
or U8191 (N_8191,N_7686,N_7881);
and U8192 (N_8192,N_7550,N_7913);
nor U8193 (N_8193,N_7844,N_7893);
nand U8194 (N_8194,N_7679,N_7560);
nand U8195 (N_8195,N_7936,N_7547);
or U8196 (N_8196,N_7692,N_7606);
nor U8197 (N_8197,N_7557,N_7616);
or U8198 (N_8198,N_7890,N_7912);
or U8199 (N_8199,N_7922,N_7595);
nor U8200 (N_8200,N_7973,N_7934);
nor U8201 (N_8201,N_7928,N_7872);
or U8202 (N_8202,N_7693,N_7788);
nor U8203 (N_8203,N_7812,N_7933);
nand U8204 (N_8204,N_7993,N_7666);
or U8205 (N_8205,N_7621,N_7678);
and U8206 (N_8206,N_7981,N_7676);
or U8207 (N_8207,N_7767,N_7732);
nor U8208 (N_8208,N_7677,N_7747);
nand U8209 (N_8209,N_7774,N_7758);
nor U8210 (N_8210,N_7827,N_7866);
nand U8211 (N_8211,N_7698,N_7609);
and U8212 (N_8212,N_7965,N_7761);
and U8213 (N_8213,N_7796,N_7551);
or U8214 (N_8214,N_7719,N_7749);
or U8215 (N_8215,N_7816,N_7520);
nor U8216 (N_8216,N_7969,N_7672);
nand U8217 (N_8217,N_7578,N_7990);
xor U8218 (N_8218,N_7612,N_7662);
and U8219 (N_8219,N_7705,N_7734);
nand U8220 (N_8220,N_7959,N_7691);
nand U8221 (N_8221,N_7745,N_7582);
or U8222 (N_8222,N_7555,N_7685);
nor U8223 (N_8223,N_7752,N_7519);
nand U8224 (N_8224,N_7645,N_7738);
and U8225 (N_8225,N_7701,N_7534);
and U8226 (N_8226,N_7847,N_7657);
nand U8227 (N_8227,N_7814,N_7723);
or U8228 (N_8228,N_7702,N_7636);
nor U8229 (N_8229,N_7862,N_7976);
nor U8230 (N_8230,N_7580,N_7623);
or U8231 (N_8231,N_7573,N_7700);
xor U8232 (N_8232,N_7769,N_7627);
nand U8233 (N_8233,N_7576,N_7801);
and U8234 (N_8234,N_7725,N_7968);
and U8235 (N_8235,N_7722,N_7604);
or U8236 (N_8236,N_7776,N_7880);
and U8237 (N_8237,N_7663,N_7824);
or U8238 (N_8238,N_7846,N_7845);
nand U8239 (N_8239,N_7798,N_7584);
or U8240 (N_8240,N_7869,N_7917);
or U8241 (N_8241,N_7742,N_7527);
or U8242 (N_8242,N_7991,N_7946);
and U8243 (N_8243,N_7809,N_7966);
nor U8244 (N_8244,N_7506,N_7883);
nand U8245 (N_8245,N_7791,N_7624);
nand U8246 (N_8246,N_7983,N_7867);
nand U8247 (N_8247,N_7566,N_7631);
and U8248 (N_8248,N_7897,N_7650);
nor U8249 (N_8249,N_7905,N_7713);
or U8250 (N_8250,N_7884,N_7770);
nand U8251 (N_8251,N_7819,N_7803);
nand U8252 (N_8252,N_7598,N_7565);
or U8253 (N_8253,N_7674,N_7684);
and U8254 (N_8254,N_7859,N_7993);
and U8255 (N_8255,N_7741,N_7636);
nand U8256 (N_8256,N_7598,N_7765);
and U8257 (N_8257,N_7782,N_7981);
or U8258 (N_8258,N_7579,N_7775);
nor U8259 (N_8259,N_7913,N_7750);
and U8260 (N_8260,N_7707,N_7964);
nand U8261 (N_8261,N_7682,N_7695);
nand U8262 (N_8262,N_7975,N_7571);
and U8263 (N_8263,N_7518,N_7535);
nand U8264 (N_8264,N_7972,N_7575);
or U8265 (N_8265,N_7831,N_7566);
nor U8266 (N_8266,N_7714,N_7947);
and U8267 (N_8267,N_7734,N_7691);
nand U8268 (N_8268,N_7849,N_7759);
nand U8269 (N_8269,N_7625,N_7525);
nand U8270 (N_8270,N_7992,N_7958);
and U8271 (N_8271,N_7870,N_7928);
or U8272 (N_8272,N_7841,N_7697);
and U8273 (N_8273,N_7636,N_7813);
nand U8274 (N_8274,N_7973,N_7910);
or U8275 (N_8275,N_7651,N_7754);
nand U8276 (N_8276,N_7904,N_7518);
nand U8277 (N_8277,N_7897,N_7970);
or U8278 (N_8278,N_7557,N_7784);
or U8279 (N_8279,N_7602,N_7912);
nand U8280 (N_8280,N_7633,N_7662);
nor U8281 (N_8281,N_7537,N_7809);
or U8282 (N_8282,N_7999,N_7730);
or U8283 (N_8283,N_7926,N_7709);
or U8284 (N_8284,N_7588,N_7816);
nor U8285 (N_8285,N_7709,N_7953);
nand U8286 (N_8286,N_7844,N_7586);
and U8287 (N_8287,N_7991,N_7533);
and U8288 (N_8288,N_7890,N_7923);
nor U8289 (N_8289,N_7834,N_7840);
nand U8290 (N_8290,N_7540,N_7945);
or U8291 (N_8291,N_7883,N_7620);
xor U8292 (N_8292,N_7596,N_7669);
and U8293 (N_8293,N_7738,N_7664);
nand U8294 (N_8294,N_7903,N_7589);
nor U8295 (N_8295,N_7644,N_7818);
nand U8296 (N_8296,N_7681,N_7809);
nor U8297 (N_8297,N_7626,N_7779);
nor U8298 (N_8298,N_7854,N_7959);
or U8299 (N_8299,N_7857,N_7764);
nand U8300 (N_8300,N_7773,N_7897);
and U8301 (N_8301,N_7799,N_7823);
nor U8302 (N_8302,N_7920,N_7834);
xnor U8303 (N_8303,N_7889,N_7582);
or U8304 (N_8304,N_7712,N_7921);
and U8305 (N_8305,N_7708,N_7624);
or U8306 (N_8306,N_7897,N_7569);
or U8307 (N_8307,N_7952,N_7920);
nand U8308 (N_8308,N_7631,N_7571);
or U8309 (N_8309,N_7553,N_7855);
and U8310 (N_8310,N_7907,N_7718);
nor U8311 (N_8311,N_7822,N_7813);
and U8312 (N_8312,N_7790,N_7961);
nor U8313 (N_8313,N_7976,N_7655);
xnor U8314 (N_8314,N_7660,N_7840);
nand U8315 (N_8315,N_7939,N_7778);
xor U8316 (N_8316,N_7711,N_7579);
nand U8317 (N_8317,N_7554,N_7567);
nand U8318 (N_8318,N_7869,N_7804);
and U8319 (N_8319,N_7673,N_7954);
and U8320 (N_8320,N_7661,N_7816);
nor U8321 (N_8321,N_7808,N_7594);
nand U8322 (N_8322,N_7549,N_7986);
nand U8323 (N_8323,N_7680,N_7963);
and U8324 (N_8324,N_7655,N_7536);
nor U8325 (N_8325,N_7985,N_7832);
nand U8326 (N_8326,N_7542,N_7997);
and U8327 (N_8327,N_7854,N_7806);
nand U8328 (N_8328,N_7861,N_7788);
nor U8329 (N_8329,N_7767,N_7868);
nor U8330 (N_8330,N_7941,N_7739);
nor U8331 (N_8331,N_7642,N_7898);
or U8332 (N_8332,N_7767,N_7942);
nand U8333 (N_8333,N_7822,N_7749);
or U8334 (N_8334,N_7970,N_7572);
nand U8335 (N_8335,N_7546,N_7760);
nand U8336 (N_8336,N_7522,N_7526);
xor U8337 (N_8337,N_7561,N_7534);
nand U8338 (N_8338,N_7873,N_7848);
and U8339 (N_8339,N_7501,N_7848);
and U8340 (N_8340,N_7825,N_7902);
nand U8341 (N_8341,N_7750,N_7697);
or U8342 (N_8342,N_7501,N_7822);
nor U8343 (N_8343,N_7973,N_7538);
and U8344 (N_8344,N_7675,N_7792);
nor U8345 (N_8345,N_7761,N_7674);
nor U8346 (N_8346,N_7820,N_7977);
or U8347 (N_8347,N_7920,N_7957);
or U8348 (N_8348,N_7509,N_7792);
and U8349 (N_8349,N_7708,N_7735);
nor U8350 (N_8350,N_7702,N_7950);
nand U8351 (N_8351,N_7849,N_7613);
and U8352 (N_8352,N_7546,N_7865);
or U8353 (N_8353,N_7825,N_7879);
nor U8354 (N_8354,N_7529,N_7640);
nand U8355 (N_8355,N_7954,N_7616);
or U8356 (N_8356,N_7814,N_7726);
or U8357 (N_8357,N_7873,N_7628);
nor U8358 (N_8358,N_7700,N_7762);
nor U8359 (N_8359,N_7716,N_7746);
nand U8360 (N_8360,N_7624,N_7561);
or U8361 (N_8361,N_7766,N_7590);
or U8362 (N_8362,N_7953,N_7819);
nor U8363 (N_8363,N_7713,N_7817);
and U8364 (N_8364,N_7836,N_7595);
nor U8365 (N_8365,N_7669,N_7620);
or U8366 (N_8366,N_7901,N_7937);
or U8367 (N_8367,N_7723,N_7922);
or U8368 (N_8368,N_7873,N_7768);
nor U8369 (N_8369,N_7831,N_7515);
nand U8370 (N_8370,N_7552,N_7909);
or U8371 (N_8371,N_7559,N_7971);
and U8372 (N_8372,N_7533,N_7677);
nand U8373 (N_8373,N_7530,N_7840);
nor U8374 (N_8374,N_7559,N_7902);
and U8375 (N_8375,N_7585,N_7588);
nand U8376 (N_8376,N_7709,N_7592);
or U8377 (N_8377,N_7676,N_7590);
xor U8378 (N_8378,N_7633,N_7674);
or U8379 (N_8379,N_7706,N_7821);
or U8380 (N_8380,N_7734,N_7779);
or U8381 (N_8381,N_7547,N_7576);
nor U8382 (N_8382,N_7538,N_7901);
and U8383 (N_8383,N_7756,N_7611);
or U8384 (N_8384,N_7623,N_7964);
nor U8385 (N_8385,N_7511,N_7520);
or U8386 (N_8386,N_7868,N_7896);
nand U8387 (N_8387,N_7671,N_7889);
nor U8388 (N_8388,N_7700,N_7945);
nand U8389 (N_8389,N_7759,N_7887);
nand U8390 (N_8390,N_7781,N_7791);
and U8391 (N_8391,N_7588,N_7958);
or U8392 (N_8392,N_7672,N_7744);
nand U8393 (N_8393,N_7914,N_7904);
or U8394 (N_8394,N_7770,N_7904);
or U8395 (N_8395,N_7715,N_7541);
or U8396 (N_8396,N_7838,N_7791);
and U8397 (N_8397,N_7543,N_7698);
or U8398 (N_8398,N_7654,N_7893);
and U8399 (N_8399,N_7508,N_7834);
and U8400 (N_8400,N_7943,N_7848);
or U8401 (N_8401,N_7883,N_7572);
or U8402 (N_8402,N_7924,N_7645);
or U8403 (N_8403,N_7910,N_7520);
nor U8404 (N_8404,N_7917,N_7700);
or U8405 (N_8405,N_7980,N_7988);
and U8406 (N_8406,N_7652,N_7509);
nor U8407 (N_8407,N_7739,N_7894);
or U8408 (N_8408,N_7729,N_7832);
nand U8409 (N_8409,N_7517,N_7987);
xnor U8410 (N_8410,N_7557,N_7542);
and U8411 (N_8411,N_7609,N_7838);
nand U8412 (N_8412,N_7738,N_7584);
nor U8413 (N_8413,N_7878,N_7951);
or U8414 (N_8414,N_7806,N_7567);
nor U8415 (N_8415,N_7556,N_7651);
nor U8416 (N_8416,N_7692,N_7540);
or U8417 (N_8417,N_7633,N_7553);
and U8418 (N_8418,N_7929,N_7825);
nand U8419 (N_8419,N_7883,N_7862);
nor U8420 (N_8420,N_7912,N_7915);
nor U8421 (N_8421,N_7884,N_7945);
nor U8422 (N_8422,N_7972,N_7908);
nor U8423 (N_8423,N_7602,N_7571);
and U8424 (N_8424,N_7972,N_7898);
nand U8425 (N_8425,N_7814,N_7947);
or U8426 (N_8426,N_7541,N_7878);
or U8427 (N_8427,N_7951,N_7809);
and U8428 (N_8428,N_7988,N_7783);
nand U8429 (N_8429,N_7566,N_7967);
nor U8430 (N_8430,N_7821,N_7971);
and U8431 (N_8431,N_7896,N_7667);
or U8432 (N_8432,N_7997,N_7886);
or U8433 (N_8433,N_7873,N_7540);
or U8434 (N_8434,N_7646,N_7966);
nand U8435 (N_8435,N_7565,N_7647);
nand U8436 (N_8436,N_7893,N_7629);
nor U8437 (N_8437,N_7898,N_7872);
and U8438 (N_8438,N_7643,N_7995);
or U8439 (N_8439,N_7891,N_7711);
and U8440 (N_8440,N_7785,N_7682);
or U8441 (N_8441,N_7700,N_7531);
and U8442 (N_8442,N_7851,N_7883);
or U8443 (N_8443,N_7937,N_7589);
and U8444 (N_8444,N_7514,N_7868);
nor U8445 (N_8445,N_7658,N_7903);
and U8446 (N_8446,N_7687,N_7657);
or U8447 (N_8447,N_7931,N_7556);
or U8448 (N_8448,N_7923,N_7627);
nand U8449 (N_8449,N_7730,N_7963);
xor U8450 (N_8450,N_7867,N_7744);
nor U8451 (N_8451,N_7570,N_7996);
and U8452 (N_8452,N_7678,N_7694);
or U8453 (N_8453,N_7901,N_7753);
xor U8454 (N_8454,N_7861,N_7996);
or U8455 (N_8455,N_7829,N_7644);
and U8456 (N_8456,N_7550,N_7788);
nor U8457 (N_8457,N_7768,N_7539);
nand U8458 (N_8458,N_7575,N_7736);
nor U8459 (N_8459,N_7609,N_7847);
nor U8460 (N_8460,N_7851,N_7700);
nor U8461 (N_8461,N_7764,N_7546);
nor U8462 (N_8462,N_7631,N_7715);
and U8463 (N_8463,N_7773,N_7785);
nand U8464 (N_8464,N_7801,N_7949);
nor U8465 (N_8465,N_7811,N_7846);
nor U8466 (N_8466,N_7831,N_7769);
xor U8467 (N_8467,N_7967,N_7700);
nand U8468 (N_8468,N_7899,N_7728);
and U8469 (N_8469,N_7825,N_7654);
nand U8470 (N_8470,N_7713,N_7681);
nor U8471 (N_8471,N_7807,N_7606);
nand U8472 (N_8472,N_7805,N_7924);
and U8473 (N_8473,N_7905,N_7853);
and U8474 (N_8474,N_7731,N_7590);
and U8475 (N_8475,N_7912,N_7944);
or U8476 (N_8476,N_7846,N_7572);
and U8477 (N_8477,N_7710,N_7795);
or U8478 (N_8478,N_7940,N_7950);
and U8479 (N_8479,N_7521,N_7555);
and U8480 (N_8480,N_7504,N_7637);
or U8481 (N_8481,N_7895,N_7879);
nor U8482 (N_8482,N_7617,N_7572);
or U8483 (N_8483,N_7812,N_7860);
xor U8484 (N_8484,N_7724,N_7817);
xnor U8485 (N_8485,N_7529,N_7795);
and U8486 (N_8486,N_7556,N_7697);
nand U8487 (N_8487,N_7750,N_7903);
or U8488 (N_8488,N_7861,N_7685);
nand U8489 (N_8489,N_7795,N_7984);
and U8490 (N_8490,N_7709,N_7560);
or U8491 (N_8491,N_7735,N_7788);
nand U8492 (N_8492,N_7628,N_7994);
and U8493 (N_8493,N_7646,N_7681);
nand U8494 (N_8494,N_7678,N_7535);
nand U8495 (N_8495,N_7747,N_7661);
nor U8496 (N_8496,N_7694,N_7813);
nand U8497 (N_8497,N_7735,N_7701);
nand U8498 (N_8498,N_7762,N_7579);
nand U8499 (N_8499,N_7957,N_7926);
nand U8500 (N_8500,N_8158,N_8032);
and U8501 (N_8501,N_8022,N_8451);
nor U8502 (N_8502,N_8450,N_8034);
or U8503 (N_8503,N_8388,N_8029);
nor U8504 (N_8504,N_8030,N_8351);
nor U8505 (N_8505,N_8169,N_8366);
nor U8506 (N_8506,N_8201,N_8418);
nand U8507 (N_8507,N_8268,N_8224);
or U8508 (N_8508,N_8109,N_8210);
nor U8509 (N_8509,N_8216,N_8409);
and U8510 (N_8510,N_8484,N_8118);
or U8511 (N_8511,N_8402,N_8037);
nand U8512 (N_8512,N_8083,N_8187);
nor U8513 (N_8513,N_8394,N_8139);
or U8514 (N_8514,N_8302,N_8249);
and U8515 (N_8515,N_8411,N_8434);
or U8516 (N_8516,N_8204,N_8212);
nor U8517 (N_8517,N_8255,N_8496);
or U8518 (N_8518,N_8129,N_8321);
xnor U8519 (N_8519,N_8382,N_8058);
nand U8520 (N_8520,N_8307,N_8476);
and U8521 (N_8521,N_8208,N_8150);
or U8522 (N_8522,N_8246,N_8011);
nand U8523 (N_8523,N_8261,N_8236);
nor U8524 (N_8524,N_8159,N_8452);
nor U8525 (N_8525,N_8341,N_8317);
nand U8526 (N_8526,N_8119,N_8316);
or U8527 (N_8527,N_8262,N_8256);
or U8528 (N_8528,N_8071,N_8379);
xnor U8529 (N_8529,N_8168,N_8333);
and U8530 (N_8530,N_8436,N_8435);
nand U8531 (N_8531,N_8339,N_8219);
nand U8532 (N_8532,N_8326,N_8322);
nand U8533 (N_8533,N_8313,N_8360);
nor U8534 (N_8534,N_8188,N_8397);
nand U8535 (N_8535,N_8495,N_8059);
nor U8536 (N_8536,N_8039,N_8403);
nand U8537 (N_8537,N_8220,N_8384);
or U8538 (N_8538,N_8026,N_8231);
nand U8539 (N_8539,N_8444,N_8069);
nand U8540 (N_8540,N_8370,N_8343);
and U8541 (N_8541,N_8222,N_8260);
or U8542 (N_8542,N_8153,N_8065);
and U8543 (N_8543,N_8448,N_8148);
or U8544 (N_8544,N_8284,N_8016);
or U8545 (N_8545,N_8116,N_8209);
and U8546 (N_8546,N_8463,N_8214);
or U8547 (N_8547,N_8354,N_8486);
nor U8548 (N_8548,N_8293,N_8286);
nor U8549 (N_8549,N_8334,N_8130);
nor U8550 (N_8550,N_8373,N_8458);
and U8551 (N_8551,N_8193,N_8346);
nor U8552 (N_8552,N_8376,N_8283);
nand U8553 (N_8553,N_8425,N_8154);
or U8554 (N_8554,N_8036,N_8252);
or U8555 (N_8555,N_8429,N_8191);
and U8556 (N_8556,N_8126,N_8002);
nor U8557 (N_8557,N_8266,N_8421);
nor U8558 (N_8558,N_8498,N_8361);
nor U8559 (N_8559,N_8371,N_8438);
and U8560 (N_8560,N_8004,N_8456);
or U8561 (N_8561,N_8289,N_8142);
nor U8562 (N_8562,N_8094,N_8424);
nor U8563 (N_8563,N_8028,N_8157);
or U8564 (N_8564,N_8018,N_8355);
nand U8565 (N_8565,N_8386,N_8096);
nor U8566 (N_8566,N_8362,N_8211);
and U8567 (N_8567,N_8171,N_8430);
nand U8568 (N_8568,N_8184,N_8198);
nor U8569 (N_8569,N_8189,N_8137);
nor U8570 (N_8570,N_8033,N_8367);
or U8571 (N_8571,N_8047,N_8152);
and U8572 (N_8572,N_8233,N_8296);
nor U8573 (N_8573,N_8015,N_8335);
nor U8574 (N_8574,N_8396,N_8064);
or U8575 (N_8575,N_8471,N_8112);
or U8576 (N_8576,N_8115,N_8248);
and U8577 (N_8577,N_8461,N_8259);
nand U8578 (N_8578,N_8074,N_8177);
or U8579 (N_8579,N_8257,N_8348);
and U8580 (N_8580,N_8320,N_8263);
or U8581 (N_8581,N_8055,N_8372);
nand U8582 (N_8582,N_8217,N_8197);
nor U8583 (N_8583,N_8353,N_8491);
nand U8584 (N_8584,N_8025,N_8291);
nand U8585 (N_8585,N_8270,N_8297);
or U8586 (N_8586,N_8108,N_8049);
nand U8587 (N_8587,N_8027,N_8063);
nor U8588 (N_8588,N_8133,N_8123);
or U8589 (N_8589,N_8079,N_8493);
and U8590 (N_8590,N_8420,N_8410);
nand U8591 (N_8591,N_8325,N_8227);
nand U8592 (N_8592,N_8172,N_8019);
nor U8593 (N_8593,N_8113,N_8488);
and U8594 (N_8594,N_8331,N_8277);
and U8595 (N_8595,N_8138,N_8087);
nor U8596 (N_8596,N_8295,N_8462);
or U8597 (N_8597,N_8243,N_8303);
or U8598 (N_8598,N_8253,N_8431);
nor U8599 (N_8599,N_8147,N_8164);
or U8600 (N_8600,N_8401,N_8440);
nand U8601 (N_8601,N_8267,N_8009);
and U8602 (N_8602,N_8368,N_8010);
nand U8603 (N_8603,N_8280,N_8186);
nand U8604 (N_8604,N_8090,N_8489);
nor U8605 (N_8605,N_8427,N_8377);
or U8606 (N_8606,N_8443,N_8180);
nand U8607 (N_8607,N_8413,N_8294);
and U8608 (N_8608,N_8332,N_8151);
or U8609 (N_8609,N_8281,N_8099);
or U8610 (N_8610,N_8043,N_8292);
and U8611 (N_8611,N_8194,N_8230);
nand U8612 (N_8612,N_8162,N_8419);
and U8613 (N_8613,N_8245,N_8469);
or U8614 (N_8614,N_8499,N_8389);
and U8615 (N_8615,N_8490,N_8311);
nand U8616 (N_8616,N_8363,N_8338);
and U8617 (N_8617,N_8156,N_8086);
nand U8618 (N_8618,N_8051,N_8244);
and U8619 (N_8619,N_8358,N_8121);
or U8620 (N_8620,N_8170,N_8276);
nor U8621 (N_8621,N_8480,N_8020);
and U8622 (N_8622,N_8299,N_8092);
nor U8623 (N_8623,N_8306,N_8237);
nor U8624 (N_8624,N_8218,N_8250);
nand U8625 (N_8625,N_8017,N_8160);
or U8626 (N_8626,N_8298,N_8046);
and U8627 (N_8627,N_8433,N_8356);
or U8628 (N_8628,N_8050,N_8124);
nand U8629 (N_8629,N_8076,N_8042);
nand U8630 (N_8630,N_8439,N_8125);
nand U8631 (N_8631,N_8131,N_8352);
nand U8632 (N_8632,N_8272,N_8182);
nand U8633 (N_8633,N_8405,N_8487);
nand U8634 (N_8634,N_8441,N_8102);
or U8635 (N_8635,N_8329,N_8144);
nor U8636 (N_8636,N_8207,N_8460);
or U8637 (N_8637,N_8008,N_8347);
or U8638 (N_8638,N_8196,N_8475);
or U8639 (N_8639,N_8225,N_8199);
or U8640 (N_8640,N_8279,N_8408);
or U8641 (N_8641,N_8359,N_8464);
nor U8642 (N_8642,N_8140,N_8416);
nand U8643 (N_8643,N_8229,N_8345);
nor U8644 (N_8644,N_8481,N_8497);
nor U8645 (N_8645,N_8141,N_8449);
nand U8646 (N_8646,N_8155,N_8457);
or U8647 (N_8647,N_8364,N_8024);
and U8648 (N_8648,N_8414,N_8235);
or U8649 (N_8649,N_8274,N_8479);
nand U8650 (N_8650,N_8422,N_8003);
or U8651 (N_8651,N_8387,N_8062);
xnor U8652 (N_8652,N_8412,N_8078);
nand U8653 (N_8653,N_8374,N_8455);
or U8654 (N_8654,N_8149,N_8007);
xor U8655 (N_8655,N_8472,N_8091);
or U8656 (N_8656,N_8205,N_8380);
or U8657 (N_8657,N_8470,N_8175);
nor U8658 (N_8658,N_8098,N_8073);
nor U8659 (N_8659,N_8107,N_8179);
nand U8660 (N_8660,N_8369,N_8127);
and U8661 (N_8661,N_8221,N_8089);
nor U8662 (N_8662,N_8340,N_8285);
nor U8663 (N_8663,N_8327,N_8135);
or U8664 (N_8664,N_8012,N_8392);
nor U8665 (N_8665,N_8206,N_8190);
nand U8666 (N_8666,N_8328,N_8305);
nor U8667 (N_8667,N_8195,N_8223);
nor U8668 (N_8668,N_8185,N_8163);
nor U8669 (N_8669,N_8324,N_8391);
and U8670 (N_8670,N_8104,N_8066);
nand U8671 (N_8671,N_8383,N_8466);
or U8672 (N_8672,N_8085,N_8428);
or U8673 (N_8673,N_8181,N_8084);
nor U8674 (N_8674,N_8178,N_8473);
nand U8675 (N_8675,N_8375,N_8278);
nor U8676 (N_8676,N_8453,N_8241);
nor U8677 (N_8677,N_8271,N_8075);
or U8678 (N_8678,N_8056,N_8040);
or U8679 (N_8679,N_8308,N_8093);
nand U8680 (N_8680,N_8398,N_8167);
or U8681 (N_8681,N_8390,N_8399);
or U8682 (N_8682,N_8264,N_8045);
nand U8683 (N_8683,N_8106,N_8315);
or U8684 (N_8684,N_8437,N_8323);
nand U8685 (N_8685,N_8415,N_8146);
nor U8686 (N_8686,N_8483,N_8395);
xnor U8687 (N_8687,N_8053,N_8203);
or U8688 (N_8688,N_8060,N_8110);
and U8689 (N_8689,N_8145,N_8021);
and U8690 (N_8690,N_8122,N_8068);
nand U8691 (N_8691,N_8136,N_8406);
or U8692 (N_8692,N_8454,N_8035);
or U8693 (N_8693,N_8215,N_8247);
and U8694 (N_8694,N_8290,N_8273);
and U8695 (N_8695,N_8006,N_8265);
nand U8696 (N_8696,N_8304,N_8057);
nand U8697 (N_8697,N_8173,N_8143);
xor U8698 (N_8698,N_8300,N_8070);
and U8699 (N_8699,N_8357,N_8097);
nor U8700 (N_8700,N_8105,N_8319);
and U8701 (N_8701,N_8350,N_8226);
nand U8702 (N_8702,N_8213,N_8120);
nor U8703 (N_8703,N_8330,N_8166);
nand U8704 (N_8704,N_8013,N_8282);
nor U8705 (N_8705,N_8128,N_8041);
or U8706 (N_8706,N_8318,N_8478);
nor U8707 (N_8707,N_8442,N_8165);
or U8708 (N_8708,N_8407,N_8474);
nand U8709 (N_8709,N_8254,N_8426);
nand U8710 (N_8710,N_8349,N_8459);
and U8711 (N_8711,N_8385,N_8067);
nor U8712 (N_8712,N_8038,N_8031);
nor U8713 (N_8713,N_8005,N_8465);
nor U8714 (N_8714,N_8000,N_8228);
nor U8715 (N_8715,N_8423,N_8072);
and U8716 (N_8716,N_8301,N_8052);
and U8717 (N_8717,N_8365,N_8378);
nor U8718 (N_8718,N_8192,N_8001);
xnor U8719 (N_8719,N_8393,N_8061);
and U8720 (N_8720,N_8269,N_8309);
and U8721 (N_8721,N_8232,N_8400);
nor U8722 (N_8722,N_8111,N_8044);
or U8723 (N_8723,N_8081,N_8023);
nand U8724 (N_8724,N_8312,N_8485);
nand U8725 (N_8725,N_8100,N_8103);
or U8726 (N_8726,N_8134,N_8239);
nand U8727 (N_8727,N_8258,N_8468);
and U8728 (N_8728,N_8494,N_8132);
nand U8729 (N_8729,N_8467,N_8251);
nand U8730 (N_8730,N_8161,N_8336);
xnor U8731 (N_8731,N_8242,N_8095);
nand U8732 (N_8732,N_8240,N_8417);
nand U8733 (N_8733,N_8200,N_8176);
or U8734 (N_8734,N_8287,N_8174);
and U8735 (N_8735,N_8447,N_8238);
and U8736 (N_8736,N_8492,N_8101);
nor U8737 (N_8737,N_8082,N_8014);
and U8738 (N_8738,N_8314,N_8275);
nor U8739 (N_8739,N_8183,N_8117);
or U8740 (N_8740,N_8404,N_8310);
and U8741 (N_8741,N_8088,N_8344);
and U8742 (N_8742,N_8381,N_8077);
and U8743 (N_8743,N_8048,N_8054);
nor U8744 (N_8744,N_8482,N_8445);
nand U8745 (N_8745,N_8234,N_8114);
or U8746 (N_8746,N_8432,N_8080);
xnor U8747 (N_8747,N_8477,N_8446);
nand U8748 (N_8748,N_8202,N_8337);
and U8749 (N_8749,N_8288,N_8342);
and U8750 (N_8750,N_8158,N_8253);
xor U8751 (N_8751,N_8052,N_8456);
or U8752 (N_8752,N_8183,N_8263);
nor U8753 (N_8753,N_8047,N_8173);
nand U8754 (N_8754,N_8466,N_8180);
or U8755 (N_8755,N_8496,N_8324);
nand U8756 (N_8756,N_8268,N_8255);
and U8757 (N_8757,N_8299,N_8290);
and U8758 (N_8758,N_8297,N_8439);
and U8759 (N_8759,N_8459,N_8042);
xor U8760 (N_8760,N_8375,N_8460);
nor U8761 (N_8761,N_8461,N_8398);
nor U8762 (N_8762,N_8144,N_8333);
nor U8763 (N_8763,N_8215,N_8001);
or U8764 (N_8764,N_8465,N_8076);
and U8765 (N_8765,N_8079,N_8215);
or U8766 (N_8766,N_8248,N_8496);
or U8767 (N_8767,N_8466,N_8305);
or U8768 (N_8768,N_8312,N_8194);
or U8769 (N_8769,N_8016,N_8162);
nand U8770 (N_8770,N_8223,N_8108);
nor U8771 (N_8771,N_8265,N_8377);
and U8772 (N_8772,N_8078,N_8344);
xor U8773 (N_8773,N_8495,N_8165);
or U8774 (N_8774,N_8211,N_8489);
nand U8775 (N_8775,N_8224,N_8210);
nand U8776 (N_8776,N_8359,N_8380);
nand U8777 (N_8777,N_8316,N_8325);
or U8778 (N_8778,N_8373,N_8198);
or U8779 (N_8779,N_8025,N_8201);
or U8780 (N_8780,N_8010,N_8086);
nand U8781 (N_8781,N_8407,N_8154);
and U8782 (N_8782,N_8018,N_8243);
nor U8783 (N_8783,N_8072,N_8036);
or U8784 (N_8784,N_8054,N_8011);
nand U8785 (N_8785,N_8435,N_8416);
nor U8786 (N_8786,N_8210,N_8239);
and U8787 (N_8787,N_8455,N_8158);
and U8788 (N_8788,N_8183,N_8428);
and U8789 (N_8789,N_8269,N_8254);
nor U8790 (N_8790,N_8011,N_8498);
nand U8791 (N_8791,N_8314,N_8068);
nand U8792 (N_8792,N_8333,N_8097);
nand U8793 (N_8793,N_8494,N_8204);
nor U8794 (N_8794,N_8359,N_8450);
and U8795 (N_8795,N_8261,N_8414);
nor U8796 (N_8796,N_8424,N_8457);
and U8797 (N_8797,N_8389,N_8313);
nor U8798 (N_8798,N_8342,N_8361);
or U8799 (N_8799,N_8212,N_8225);
and U8800 (N_8800,N_8072,N_8102);
and U8801 (N_8801,N_8452,N_8262);
nand U8802 (N_8802,N_8373,N_8302);
or U8803 (N_8803,N_8082,N_8022);
or U8804 (N_8804,N_8392,N_8411);
or U8805 (N_8805,N_8272,N_8279);
and U8806 (N_8806,N_8239,N_8238);
nor U8807 (N_8807,N_8418,N_8156);
and U8808 (N_8808,N_8460,N_8301);
or U8809 (N_8809,N_8239,N_8151);
or U8810 (N_8810,N_8282,N_8074);
nor U8811 (N_8811,N_8298,N_8135);
nand U8812 (N_8812,N_8040,N_8210);
or U8813 (N_8813,N_8432,N_8232);
and U8814 (N_8814,N_8464,N_8051);
nor U8815 (N_8815,N_8229,N_8401);
or U8816 (N_8816,N_8396,N_8158);
nand U8817 (N_8817,N_8133,N_8210);
or U8818 (N_8818,N_8230,N_8183);
and U8819 (N_8819,N_8272,N_8292);
or U8820 (N_8820,N_8219,N_8443);
nor U8821 (N_8821,N_8032,N_8222);
xnor U8822 (N_8822,N_8259,N_8454);
nor U8823 (N_8823,N_8244,N_8041);
nand U8824 (N_8824,N_8341,N_8171);
or U8825 (N_8825,N_8418,N_8132);
or U8826 (N_8826,N_8102,N_8050);
or U8827 (N_8827,N_8092,N_8421);
xnor U8828 (N_8828,N_8194,N_8255);
and U8829 (N_8829,N_8269,N_8317);
nand U8830 (N_8830,N_8484,N_8240);
or U8831 (N_8831,N_8465,N_8009);
and U8832 (N_8832,N_8053,N_8419);
nor U8833 (N_8833,N_8242,N_8161);
xor U8834 (N_8834,N_8245,N_8242);
or U8835 (N_8835,N_8172,N_8116);
nor U8836 (N_8836,N_8445,N_8248);
or U8837 (N_8837,N_8285,N_8342);
nand U8838 (N_8838,N_8440,N_8454);
nand U8839 (N_8839,N_8063,N_8254);
or U8840 (N_8840,N_8117,N_8149);
and U8841 (N_8841,N_8142,N_8420);
and U8842 (N_8842,N_8463,N_8180);
nand U8843 (N_8843,N_8082,N_8313);
and U8844 (N_8844,N_8421,N_8343);
nor U8845 (N_8845,N_8182,N_8333);
nand U8846 (N_8846,N_8298,N_8249);
nand U8847 (N_8847,N_8114,N_8101);
or U8848 (N_8848,N_8404,N_8321);
and U8849 (N_8849,N_8122,N_8087);
or U8850 (N_8850,N_8334,N_8482);
or U8851 (N_8851,N_8442,N_8356);
nor U8852 (N_8852,N_8205,N_8069);
or U8853 (N_8853,N_8164,N_8075);
nand U8854 (N_8854,N_8282,N_8125);
nor U8855 (N_8855,N_8243,N_8317);
nand U8856 (N_8856,N_8368,N_8088);
nand U8857 (N_8857,N_8304,N_8105);
and U8858 (N_8858,N_8141,N_8442);
and U8859 (N_8859,N_8255,N_8282);
nor U8860 (N_8860,N_8125,N_8297);
or U8861 (N_8861,N_8067,N_8371);
nor U8862 (N_8862,N_8472,N_8111);
nand U8863 (N_8863,N_8035,N_8462);
nor U8864 (N_8864,N_8090,N_8385);
nor U8865 (N_8865,N_8357,N_8072);
nor U8866 (N_8866,N_8336,N_8335);
xor U8867 (N_8867,N_8488,N_8015);
nand U8868 (N_8868,N_8084,N_8222);
nor U8869 (N_8869,N_8297,N_8192);
nand U8870 (N_8870,N_8229,N_8247);
xnor U8871 (N_8871,N_8343,N_8233);
or U8872 (N_8872,N_8242,N_8224);
nor U8873 (N_8873,N_8401,N_8134);
and U8874 (N_8874,N_8112,N_8025);
or U8875 (N_8875,N_8171,N_8301);
nand U8876 (N_8876,N_8006,N_8360);
nand U8877 (N_8877,N_8157,N_8000);
and U8878 (N_8878,N_8224,N_8002);
nand U8879 (N_8879,N_8468,N_8486);
nand U8880 (N_8880,N_8026,N_8201);
and U8881 (N_8881,N_8262,N_8145);
nand U8882 (N_8882,N_8449,N_8122);
or U8883 (N_8883,N_8094,N_8142);
nor U8884 (N_8884,N_8484,N_8238);
or U8885 (N_8885,N_8083,N_8284);
nor U8886 (N_8886,N_8461,N_8480);
nor U8887 (N_8887,N_8191,N_8033);
nand U8888 (N_8888,N_8053,N_8238);
nor U8889 (N_8889,N_8345,N_8361);
nand U8890 (N_8890,N_8362,N_8289);
nor U8891 (N_8891,N_8494,N_8035);
nand U8892 (N_8892,N_8123,N_8291);
nand U8893 (N_8893,N_8166,N_8418);
nand U8894 (N_8894,N_8454,N_8215);
and U8895 (N_8895,N_8432,N_8158);
or U8896 (N_8896,N_8078,N_8375);
or U8897 (N_8897,N_8181,N_8346);
or U8898 (N_8898,N_8489,N_8481);
or U8899 (N_8899,N_8466,N_8222);
or U8900 (N_8900,N_8056,N_8191);
nand U8901 (N_8901,N_8237,N_8234);
and U8902 (N_8902,N_8057,N_8034);
and U8903 (N_8903,N_8372,N_8123);
xnor U8904 (N_8904,N_8477,N_8431);
or U8905 (N_8905,N_8337,N_8429);
and U8906 (N_8906,N_8409,N_8404);
or U8907 (N_8907,N_8236,N_8223);
or U8908 (N_8908,N_8223,N_8384);
or U8909 (N_8909,N_8454,N_8368);
nand U8910 (N_8910,N_8415,N_8283);
xor U8911 (N_8911,N_8005,N_8333);
nand U8912 (N_8912,N_8250,N_8300);
or U8913 (N_8913,N_8101,N_8242);
xor U8914 (N_8914,N_8146,N_8360);
nor U8915 (N_8915,N_8310,N_8247);
nand U8916 (N_8916,N_8198,N_8476);
nor U8917 (N_8917,N_8166,N_8125);
and U8918 (N_8918,N_8454,N_8136);
or U8919 (N_8919,N_8210,N_8362);
nor U8920 (N_8920,N_8475,N_8118);
nand U8921 (N_8921,N_8461,N_8123);
nand U8922 (N_8922,N_8191,N_8480);
and U8923 (N_8923,N_8366,N_8458);
nand U8924 (N_8924,N_8458,N_8060);
nor U8925 (N_8925,N_8331,N_8452);
nor U8926 (N_8926,N_8036,N_8114);
nand U8927 (N_8927,N_8263,N_8438);
or U8928 (N_8928,N_8137,N_8093);
nand U8929 (N_8929,N_8395,N_8273);
and U8930 (N_8930,N_8480,N_8315);
nor U8931 (N_8931,N_8323,N_8339);
nor U8932 (N_8932,N_8216,N_8439);
and U8933 (N_8933,N_8223,N_8040);
nand U8934 (N_8934,N_8355,N_8303);
and U8935 (N_8935,N_8370,N_8435);
nand U8936 (N_8936,N_8426,N_8483);
or U8937 (N_8937,N_8394,N_8364);
or U8938 (N_8938,N_8224,N_8260);
nor U8939 (N_8939,N_8144,N_8478);
and U8940 (N_8940,N_8024,N_8348);
nor U8941 (N_8941,N_8047,N_8297);
and U8942 (N_8942,N_8381,N_8467);
nor U8943 (N_8943,N_8000,N_8025);
nand U8944 (N_8944,N_8455,N_8356);
or U8945 (N_8945,N_8445,N_8375);
or U8946 (N_8946,N_8199,N_8240);
nor U8947 (N_8947,N_8213,N_8453);
and U8948 (N_8948,N_8453,N_8421);
nand U8949 (N_8949,N_8201,N_8360);
or U8950 (N_8950,N_8377,N_8171);
nor U8951 (N_8951,N_8463,N_8128);
or U8952 (N_8952,N_8307,N_8336);
nor U8953 (N_8953,N_8345,N_8386);
or U8954 (N_8954,N_8389,N_8375);
and U8955 (N_8955,N_8149,N_8289);
nor U8956 (N_8956,N_8064,N_8429);
nor U8957 (N_8957,N_8283,N_8279);
nand U8958 (N_8958,N_8365,N_8472);
nand U8959 (N_8959,N_8366,N_8010);
nand U8960 (N_8960,N_8466,N_8039);
nand U8961 (N_8961,N_8121,N_8234);
and U8962 (N_8962,N_8486,N_8374);
nor U8963 (N_8963,N_8139,N_8089);
or U8964 (N_8964,N_8371,N_8365);
nand U8965 (N_8965,N_8011,N_8424);
nor U8966 (N_8966,N_8108,N_8129);
nand U8967 (N_8967,N_8309,N_8481);
or U8968 (N_8968,N_8131,N_8394);
and U8969 (N_8969,N_8042,N_8092);
nand U8970 (N_8970,N_8334,N_8234);
or U8971 (N_8971,N_8207,N_8095);
nor U8972 (N_8972,N_8314,N_8488);
nor U8973 (N_8973,N_8228,N_8314);
nor U8974 (N_8974,N_8455,N_8025);
or U8975 (N_8975,N_8283,N_8244);
nor U8976 (N_8976,N_8253,N_8401);
and U8977 (N_8977,N_8298,N_8139);
nor U8978 (N_8978,N_8400,N_8377);
or U8979 (N_8979,N_8303,N_8161);
nor U8980 (N_8980,N_8334,N_8369);
nand U8981 (N_8981,N_8442,N_8090);
nand U8982 (N_8982,N_8322,N_8486);
and U8983 (N_8983,N_8168,N_8476);
nor U8984 (N_8984,N_8497,N_8224);
nor U8985 (N_8985,N_8031,N_8304);
nor U8986 (N_8986,N_8334,N_8242);
or U8987 (N_8987,N_8253,N_8124);
or U8988 (N_8988,N_8307,N_8406);
and U8989 (N_8989,N_8055,N_8345);
nor U8990 (N_8990,N_8065,N_8433);
or U8991 (N_8991,N_8459,N_8455);
nand U8992 (N_8992,N_8374,N_8040);
and U8993 (N_8993,N_8010,N_8491);
xor U8994 (N_8994,N_8284,N_8495);
or U8995 (N_8995,N_8256,N_8223);
nor U8996 (N_8996,N_8257,N_8045);
nand U8997 (N_8997,N_8292,N_8047);
or U8998 (N_8998,N_8461,N_8053);
nand U8999 (N_8999,N_8199,N_8078);
or U9000 (N_9000,N_8968,N_8787);
nor U9001 (N_9001,N_8526,N_8752);
or U9002 (N_9002,N_8726,N_8953);
nor U9003 (N_9003,N_8841,N_8917);
nor U9004 (N_9004,N_8609,N_8505);
nor U9005 (N_9005,N_8608,N_8734);
and U9006 (N_9006,N_8569,N_8692);
and U9007 (N_9007,N_8924,N_8804);
nand U9008 (N_9008,N_8696,N_8993);
or U9009 (N_9009,N_8894,N_8768);
or U9010 (N_9010,N_8670,N_8691);
nand U9011 (N_9011,N_8688,N_8948);
and U9012 (N_9012,N_8888,N_8982);
and U9013 (N_9013,N_8748,N_8703);
and U9014 (N_9014,N_8746,N_8519);
or U9015 (N_9015,N_8643,N_8880);
and U9016 (N_9016,N_8862,N_8818);
or U9017 (N_9017,N_8977,N_8925);
and U9018 (N_9018,N_8795,N_8758);
and U9019 (N_9019,N_8771,N_8646);
and U9020 (N_9020,N_8914,N_8549);
nor U9021 (N_9021,N_8855,N_8567);
and U9022 (N_9022,N_8834,N_8551);
or U9023 (N_9023,N_8920,N_8513);
and U9024 (N_9024,N_8521,N_8750);
or U9025 (N_9025,N_8582,N_8839);
nor U9026 (N_9026,N_8742,N_8681);
xor U9027 (N_9027,N_8859,N_8927);
nand U9028 (N_9028,N_8808,N_8861);
nor U9029 (N_9029,N_8868,N_8659);
nand U9030 (N_9030,N_8676,N_8538);
or U9031 (N_9031,N_8805,N_8835);
or U9032 (N_9032,N_8731,N_8934);
or U9033 (N_9033,N_8810,N_8829);
nor U9034 (N_9034,N_8864,N_8600);
nor U9035 (N_9035,N_8830,N_8735);
or U9036 (N_9036,N_8556,N_8890);
and U9037 (N_9037,N_8933,N_8824);
nand U9038 (N_9038,N_8509,N_8929);
or U9039 (N_9039,N_8913,N_8852);
and U9040 (N_9040,N_8812,N_8882);
nand U9041 (N_9041,N_8940,N_8561);
nand U9042 (N_9042,N_8784,N_8789);
nor U9043 (N_9043,N_8632,N_8751);
and U9044 (N_9044,N_8557,N_8571);
and U9045 (N_9045,N_8649,N_8544);
or U9046 (N_9046,N_8781,N_8870);
nand U9047 (N_9047,N_8564,N_8858);
nand U9048 (N_9048,N_8941,N_8554);
nor U9049 (N_9049,N_8798,N_8959);
nand U9050 (N_9050,N_8840,N_8767);
xnor U9051 (N_9051,N_8598,N_8972);
nand U9052 (N_9052,N_8764,N_8645);
nand U9053 (N_9053,N_8685,N_8727);
and U9054 (N_9054,N_8639,N_8740);
or U9055 (N_9055,N_8694,N_8893);
xnor U9056 (N_9056,N_8618,N_8744);
and U9057 (N_9057,N_8823,N_8826);
and U9058 (N_9058,N_8991,N_8833);
nor U9059 (N_9059,N_8821,N_8850);
nand U9060 (N_9060,N_8867,N_8715);
xor U9061 (N_9061,N_8552,N_8563);
nand U9062 (N_9062,N_8875,N_8510);
xor U9063 (N_9063,N_8966,N_8816);
or U9064 (N_9064,N_8626,N_8535);
xnor U9065 (N_9065,N_8760,N_8678);
nor U9066 (N_9066,N_8709,N_8625);
or U9067 (N_9067,N_8668,N_8539);
and U9068 (N_9068,N_8857,N_8895);
and U9069 (N_9069,N_8911,N_8842);
and U9070 (N_9070,N_8517,N_8838);
nor U9071 (N_9071,N_8931,N_8613);
or U9072 (N_9072,N_8910,N_8997);
nor U9073 (N_9073,N_8956,N_8873);
nor U9074 (N_9074,N_8515,N_8932);
nand U9075 (N_9075,N_8674,N_8516);
or U9076 (N_9076,N_8642,N_8507);
and U9077 (N_9077,N_8522,N_8963);
nor U9078 (N_9078,N_8733,N_8908);
or U9079 (N_9079,N_8905,N_8624);
and U9080 (N_9080,N_8992,N_8780);
nor U9081 (N_9081,N_8954,N_8779);
nand U9082 (N_9082,N_8669,N_8884);
or U9083 (N_9083,N_8774,N_8930);
nor U9084 (N_9084,N_8573,N_8949);
nor U9085 (N_9085,N_8813,N_8874);
and U9086 (N_9086,N_8541,N_8753);
and U9087 (N_9087,N_8595,N_8897);
nor U9088 (N_9088,N_8602,N_8596);
nand U9089 (N_9089,N_8979,N_8553);
or U9090 (N_9090,N_8887,N_8629);
nor U9091 (N_9091,N_8854,N_8711);
nand U9092 (N_9092,N_8778,N_8540);
nor U9093 (N_9093,N_8807,N_8757);
or U9094 (N_9094,N_8714,N_8971);
and U9095 (N_9095,N_8577,N_8891);
or U9096 (N_9096,N_8630,N_8654);
nor U9097 (N_9097,N_8756,N_8743);
nor U9098 (N_9098,N_8721,N_8947);
or U9099 (N_9099,N_8885,N_8531);
nand U9100 (N_9100,N_8975,N_8783);
or U9101 (N_9101,N_8699,N_8621);
and U9102 (N_9102,N_8590,N_8586);
nand U9103 (N_9103,N_8550,N_8759);
or U9104 (N_9104,N_8723,N_8653);
or U9105 (N_9105,N_8533,N_8926);
nor U9106 (N_9106,N_8631,N_8928);
nor U9107 (N_9107,N_8876,N_8652);
and U9108 (N_9108,N_8606,N_8555);
and U9109 (N_9109,N_8747,N_8901);
nand U9110 (N_9110,N_8846,N_8523);
and U9111 (N_9111,N_8529,N_8601);
nand U9112 (N_9112,N_8922,N_8945);
nor U9113 (N_9113,N_8660,N_8524);
nand U9114 (N_9114,N_8782,N_8607);
or U9115 (N_9115,N_8961,N_8650);
nor U9116 (N_9116,N_8615,N_8981);
and U9117 (N_9117,N_8984,N_8628);
nand U9118 (N_9118,N_8623,N_8988);
or U9119 (N_9119,N_8937,N_8728);
nand U9120 (N_9120,N_8872,N_8849);
nand U9121 (N_9121,N_8869,N_8587);
nor U9122 (N_9122,N_8525,N_8677);
nand U9123 (N_9123,N_8800,N_8558);
nand U9124 (N_9124,N_8773,N_8597);
xnor U9125 (N_9125,N_8796,N_8527);
and U9126 (N_9126,N_8866,N_8634);
nand U9127 (N_9127,N_8762,N_8579);
or U9128 (N_9128,N_8766,N_8665);
and U9129 (N_9129,N_8970,N_8548);
nor U9130 (N_9130,N_8967,N_8831);
or U9131 (N_9131,N_8794,N_8916);
and U9132 (N_9132,N_8611,N_8679);
or U9133 (N_9133,N_8730,N_8955);
nand U9134 (N_9134,N_8655,N_8819);
nand U9135 (N_9135,N_8612,N_8543);
and U9136 (N_9136,N_8680,N_8969);
nor U9137 (N_9137,N_8616,N_8575);
nor U9138 (N_9138,N_8705,N_8990);
nand U9139 (N_9139,N_8675,N_8536);
xnor U9140 (N_9140,N_8799,N_8713);
or U9141 (N_9141,N_8589,N_8903);
or U9142 (N_9142,N_8724,N_8614);
or U9143 (N_9143,N_8985,N_8879);
nand U9144 (N_9144,N_8749,N_8820);
or U9145 (N_9145,N_8907,N_8702);
or U9146 (N_9146,N_8761,N_8664);
or U9147 (N_9147,N_8738,N_8877);
nand U9148 (N_9148,N_8998,N_8801);
or U9149 (N_9149,N_8637,N_8690);
nand U9150 (N_9150,N_8958,N_8619);
or U9151 (N_9151,N_8562,N_8851);
or U9152 (N_9152,N_8732,N_8938);
nand U9153 (N_9153,N_8964,N_8661);
or U9154 (N_9154,N_8772,N_8693);
and U9155 (N_9155,N_8904,N_8547);
nand U9156 (N_9156,N_8936,N_8909);
or U9157 (N_9157,N_8776,N_8765);
nand U9158 (N_9158,N_8594,N_8974);
or U9159 (N_9159,N_8737,N_8710);
nor U9160 (N_9160,N_8500,N_8528);
nor U9161 (N_9161,N_8912,N_8657);
nor U9162 (N_9162,N_8817,N_8576);
and U9163 (N_9163,N_8745,N_8865);
or U9164 (N_9164,N_8504,N_8574);
or U9165 (N_9165,N_8610,N_8683);
and U9166 (N_9166,N_8844,N_8514);
nor U9167 (N_9167,N_8542,N_8792);
and U9168 (N_9168,N_8572,N_8845);
nor U9169 (N_9169,N_8718,N_8532);
nor U9170 (N_9170,N_8518,N_8899);
or U9171 (N_9171,N_8682,N_8648);
or U9172 (N_9172,N_8565,N_8863);
nand U9173 (N_9173,N_8503,N_8950);
nor U9174 (N_9174,N_8622,N_8803);
or U9175 (N_9175,N_8987,N_8739);
nand U9176 (N_9176,N_8906,N_8627);
nor U9177 (N_9177,N_8814,N_8822);
xnor U9178 (N_9178,N_8825,N_8667);
nand U9179 (N_9179,N_8508,N_8791);
nand U9180 (N_9180,N_8722,N_8832);
and U9181 (N_9181,N_8843,N_8881);
xnor U9182 (N_9182,N_8944,N_8570);
and U9183 (N_9183,N_8725,N_8896);
and U9184 (N_9184,N_8797,N_8883);
or U9185 (N_9185,N_8530,N_8915);
and U9186 (N_9186,N_8889,N_8785);
nand U9187 (N_9187,N_8546,N_8697);
nand U9188 (N_9188,N_8684,N_8999);
or U9189 (N_9189,N_8886,N_8566);
nor U9190 (N_9190,N_8698,N_8689);
or U9191 (N_9191,N_8658,N_8617);
nand U9192 (N_9192,N_8581,N_8996);
nand U9193 (N_9193,N_8712,N_8716);
nand U9194 (N_9194,N_8636,N_8847);
nand U9195 (N_9195,N_8770,N_8662);
nor U9196 (N_9196,N_8520,N_8793);
or U9197 (N_9197,N_8786,N_8837);
nand U9198 (N_9198,N_8788,N_8647);
nand U9199 (N_9199,N_8918,N_8695);
nor U9200 (N_9200,N_8871,N_8989);
and U9201 (N_9201,N_8605,N_8860);
nand U9202 (N_9202,N_8651,N_8700);
and U9203 (N_9203,N_8736,N_8878);
nand U9204 (N_9204,N_8960,N_8671);
nor U9205 (N_9205,N_8923,N_8717);
or U9206 (N_9206,N_8638,N_8635);
nand U9207 (N_9207,N_8811,N_8719);
nand U9208 (N_9208,N_8640,N_8603);
or U9209 (N_9209,N_8560,N_8707);
nand U9210 (N_9210,N_8973,N_8686);
nor U9211 (N_9211,N_8900,N_8806);
or U9212 (N_9212,N_8815,N_8720);
and U9213 (N_9213,N_8836,N_8965);
and U9214 (N_9214,N_8763,N_8980);
nand U9215 (N_9215,N_8978,N_8583);
nor U9216 (N_9216,N_8501,N_8604);
and U9217 (N_9217,N_8592,N_8706);
nor U9218 (N_9218,N_8943,N_8939);
and U9219 (N_9219,N_8942,N_8741);
or U9220 (N_9220,N_8957,N_8620);
and U9221 (N_9221,N_8673,N_8827);
or U9222 (N_9222,N_8599,N_8666);
nor U9223 (N_9223,N_8809,N_8769);
or U9224 (N_9224,N_8585,N_8946);
and U9225 (N_9225,N_8580,N_8790);
nor U9226 (N_9226,N_8672,N_8545);
and U9227 (N_9227,N_8952,N_8593);
or U9228 (N_9228,N_8512,N_8578);
or U9229 (N_9229,N_8708,N_8898);
nor U9230 (N_9230,N_8633,N_8919);
nor U9231 (N_9231,N_8962,N_8754);
or U9232 (N_9232,N_8951,N_8892);
or U9233 (N_9233,N_8986,N_8511);
nor U9234 (N_9234,N_8502,N_8644);
and U9235 (N_9235,N_8663,N_8687);
nand U9236 (N_9236,N_8534,N_8995);
or U9237 (N_9237,N_8588,N_8976);
or U9238 (N_9238,N_8902,N_8537);
nor U9239 (N_9239,N_8559,N_8568);
xor U9240 (N_9240,N_8729,N_8921);
nand U9241 (N_9241,N_8994,N_8584);
or U9242 (N_9242,N_8591,N_8755);
or U9243 (N_9243,N_8802,N_8641);
nor U9244 (N_9244,N_8656,N_8848);
nand U9245 (N_9245,N_8853,N_8828);
or U9246 (N_9246,N_8506,N_8704);
nor U9247 (N_9247,N_8777,N_8856);
nor U9248 (N_9248,N_8701,N_8983);
nand U9249 (N_9249,N_8935,N_8775);
nand U9250 (N_9250,N_8741,N_8685);
or U9251 (N_9251,N_8927,N_8686);
nor U9252 (N_9252,N_8898,N_8692);
nand U9253 (N_9253,N_8961,N_8820);
or U9254 (N_9254,N_8806,N_8701);
nor U9255 (N_9255,N_8877,N_8663);
nor U9256 (N_9256,N_8940,N_8590);
or U9257 (N_9257,N_8909,N_8852);
nand U9258 (N_9258,N_8784,N_8739);
nand U9259 (N_9259,N_8558,N_8713);
nor U9260 (N_9260,N_8536,N_8812);
and U9261 (N_9261,N_8935,N_8653);
nand U9262 (N_9262,N_8560,N_8523);
nand U9263 (N_9263,N_8969,N_8950);
or U9264 (N_9264,N_8551,N_8920);
and U9265 (N_9265,N_8651,N_8883);
nand U9266 (N_9266,N_8559,N_8746);
or U9267 (N_9267,N_8683,N_8767);
and U9268 (N_9268,N_8572,N_8522);
nand U9269 (N_9269,N_8773,N_8762);
nor U9270 (N_9270,N_8553,N_8551);
nand U9271 (N_9271,N_8607,N_8685);
nand U9272 (N_9272,N_8908,N_8634);
and U9273 (N_9273,N_8817,N_8704);
nor U9274 (N_9274,N_8979,N_8622);
nor U9275 (N_9275,N_8507,N_8708);
nand U9276 (N_9276,N_8563,N_8638);
nor U9277 (N_9277,N_8920,N_8884);
or U9278 (N_9278,N_8529,N_8903);
or U9279 (N_9279,N_8627,N_8790);
and U9280 (N_9280,N_8841,N_8591);
nand U9281 (N_9281,N_8928,N_8728);
nor U9282 (N_9282,N_8590,N_8577);
and U9283 (N_9283,N_8931,N_8989);
nand U9284 (N_9284,N_8738,N_8623);
nor U9285 (N_9285,N_8966,N_8832);
nand U9286 (N_9286,N_8790,N_8702);
nand U9287 (N_9287,N_8656,N_8799);
or U9288 (N_9288,N_8540,N_8828);
nor U9289 (N_9289,N_8579,N_8694);
and U9290 (N_9290,N_8522,N_8752);
nor U9291 (N_9291,N_8527,N_8898);
and U9292 (N_9292,N_8709,N_8507);
and U9293 (N_9293,N_8829,N_8989);
or U9294 (N_9294,N_8555,N_8982);
and U9295 (N_9295,N_8512,N_8624);
nand U9296 (N_9296,N_8715,N_8811);
nor U9297 (N_9297,N_8980,N_8516);
nor U9298 (N_9298,N_8771,N_8592);
or U9299 (N_9299,N_8550,N_8713);
xor U9300 (N_9300,N_8679,N_8542);
nor U9301 (N_9301,N_8517,N_8625);
nand U9302 (N_9302,N_8645,N_8692);
or U9303 (N_9303,N_8959,N_8517);
nand U9304 (N_9304,N_8694,N_8516);
nand U9305 (N_9305,N_8580,N_8599);
and U9306 (N_9306,N_8626,N_8856);
and U9307 (N_9307,N_8859,N_8772);
nor U9308 (N_9308,N_8950,N_8979);
and U9309 (N_9309,N_8817,N_8889);
nand U9310 (N_9310,N_8956,N_8558);
nor U9311 (N_9311,N_8967,N_8648);
nor U9312 (N_9312,N_8575,N_8742);
or U9313 (N_9313,N_8820,N_8805);
nor U9314 (N_9314,N_8904,N_8655);
or U9315 (N_9315,N_8678,N_8568);
nand U9316 (N_9316,N_8563,N_8537);
or U9317 (N_9317,N_8920,N_8742);
or U9318 (N_9318,N_8988,N_8554);
or U9319 (N_9319,N_8641,N_8574);
or U9320 (N_9320,N_8646,N_8688);
or U9321 (N_9321,N_8813,N_8732);
or U9322 (N_9322,N_8614,N_8839);
and U9323 (N_9323,N_8963,N_8670);
nand U9324 (N_9324,N_8766,N_8947);
nor U9325 (N_9325,N_8555,N_8560);
and U9326 (N_9326,N_8632,N_8611);
nor U9327 (N_9327,N_8767,N_8596);
and U9328 (N_9328,N_8536,N_8725);
nand U9329 (N_9329,N_8542,N_8893);
and U9330 (N_9330,N_8549,N_8974);
nand U9331 (N_9331,N_8849,N_8946);
nand U9332 (N_9332,N_8806,N_8983);
nor U9333 (N_9333,N_8912,N_8969);
nand U9334 (N_9334,N_8569,N_8675);
or U9335 (N_9335,N_8529,N_8620);
and U9336 (N_9336,N_8934,N_8521);
or U9337 (N_9337,N_8653,N_8567);
nor U9338 (N_9338,N_8994,N_8975);
nor U9339 (N_9339,N_8735,N_8574);
and U9340 (N_9340,N_8714,N_8602);
nand U9341 (N_9341,N_8582,N_8615);
nand U9342 (N_9342,N_8872,N_8560);
nand U9343 (N_9343,N_8719,N_8895);
or U9344 (N_9344,N_8709,N_8510);
or U9345 (N_9345,N_8988,N_8933);
and U9346 (N_9346,N_8996,N_8641);
or U9347 (N_9347,N_8691,N_8846);
and U9348 (N_9348,N_8854,N_8930);
and U9349 (N_9349,N_8815,N_8524);
nand U9350 (N_9350,N_8815,N_8772);
nand U9351 (N_9351,N_8725,N_8780);
nor U9352 (N_9352,N_8914,N_8964);
xnor U9353 (N_9353,N_8549,N_8515);
or U9354 (N_9354,N_8747,N_8552);
and U9355 (N_9355,N_8706,N_8854);
and U9356 (N_9356,N_8664,N_8876);
nor U9357 (N_9357,N_8845,N_8502);
or U9358 (N_9358,N_8517,N_8579);
and U9359 (N_9359,N_8747,N_8870);
nor U9360 (N_9360,N_8789,N_8737);
or U9361 (N_9361,N_8788,N_8797);
and U9362 (N_9362,N_8912,N_8862);
nand U9363 (N_9363,N_8696,N_8569);
nand U9364 (N_9364,N_8915,N_8933);
or U9365 (N_9365,N_8675,N_8897);
nand U9366 (N_9366,N_8650,N_8670);
nand U9367 (N_9367,N_8611,N_8633);
nor U9368 (N_9368,N_8812,N_8803);
or U9369 (N_9369,N_8735,N_8904);
nand U9370 (N_9370,N_8974,N_8747);
xor U9371 (N_9371,N_8894,N_8694);
nor U9372 (N_9372,N_8918,N_8814);
or U9373 (N_9373,N_8894,N_8555);
and U9374 (N_9374,N_8976,N_8863);
and U9375 (N_9375,N_8864,N_8646);
or U9376 (N_9376,N_8611,N_8523);
and U9377 (N_9377,N_8905,N_8973);
and U9378 (N_9378,N_8620,N_8521);
nor U9379 (N_9379,N_8713,N_8528);
or U9380 (N_9380,N_8545,N_8613);
and U9381 (N_9381,N_8599,N_8989);
nand U9382 (N_9382,N_8514,N_8649);
or U9383 (N_9383,N_8674,N_8520);
nor U9384 (N_9384,N_8998,N_8938);
nor U9385 (N_9385,N_8860,N_8571);
nor U9386 (N_9386,N_8550,N_8564);
nand U9387 (N_9387,N_8514,N_8577);
and U9388 (N_9388,N_8908,N_8570);
nand U9389 (N_9389,N_8918,N_8938);
nor U9390 (N_9390,N_8613,N_8723);
nor U9391 (N_9391,N_8898,N_8978);
or U9392 (N_9392,N_8760,N_8554);
and U9393 (N_9393,N_8674,N_8765);
or U9394 (N_9394,N_8641,N_8842);
nor U9395 (N_9395,N_8573,N_8602);
nand U9396 (N_9396,N_8549,N_8925);
or U9397 (N_9397,N_8953,N_8893);
nand U9398 (N_9398,N_8639,N_8977);
or U9399 (N_9399,N_8746,N_8741);
nand U9400 (N_9400,N_8711,N_8945);
nand U9401 (N_9401,N_8914,N_8627);
nand U9402 (N_9402,N_8524,N_8980);
or U9403 (N_9403,N_8724,N_8519);
nand U9404 (N_9404,N_8672,N_8687);
or U9405 (N_9405,N_8823,N_8710);
nand U9406 (N_9406,N_8742,N_8504);
and U9407 (N_9407,N_8838,N_8679);
and U9408 (N_9408,N_8992,N_8713);
and U9409 (N_9409,N_8652,N_8547);
and U9410 (N_9410,N_8770,N_8772);
and U9411 (N_9411,N_8890,N_8657);
nand U9412 (N_9412,N_8801,N_8645);
xor U9413 (N_9413,N_8831,N_8731);
or U9414 (N_9414,N_8584,N_8877);
nand U9415 (N_9415,N_8971,N_8628);
nor U9416 (N_9416,N_8606,N_8633);
nor U9417 (N_9417,N_8763,N_8800);
or U9418 (N_9418,N_8710,N_8578);
xor U9419 (N_9419,N_8868,N_8803);
and U9420 (N_9420,N_8760,N_8884);
and U9421 (N_9421,N_8668,N_8721);
nand U9422 (N_9422,N_8795,N_8905);
nor U9423 (N_9423,N_8682,N_8608);
nor U9424 (N_9424,N_8653,N_8608);
nor U9425 (N_9425,N_8500,N_8744);
nor U9426 (N_9426,N_8826,N_8780);
and U9427 (N_9427,N_8610,N_8552);
and U9428 (N_9428,N_8538,N_8847);
or U9429 (N_9429,N_8755,N_8598);
nand U9430 (N_9430,N_8800,N_8660);
nand U9431 (N_9431,N_8578,N_8972);
nor U9432 (N_9432,N_8905,N_8955);
or U9433 (N_9433,N_8514,N_8973);
nor U9434 (N_9434,N_8682,N_8892);
nand U9435 (N_9435,N_8976,N_8566);
or U9436 (N_9436,N_8678,N_8507);
nor U9437 (N_9437,N_8650,N_8560);
nand U9438 (N_9438,N_8978,N_8837);
or U9439 (N_9439,N_8746,N_8542);
nor U9440 (N_9440,N_8878,N_8851);
or U9441 (N_9441,N_8895,N_8835);
or U9442 (N_9442,N_8660,N_8619);
or U9443 (N_9443,N_8836,N_8719);
nand U9444 (N_9444,N_8649,N_8989);
nor U9445 (N_9445,N_8547,N_8775);
or U9446 (N_9446,N_8672,N_8962);
or U9447 (N_9447,N_8674,N_8638);
and U9448 (N_9448,N_8522,N_8684);
nor U9449 (N_9449,N_8641,N_8541);
nor U9450 (N_9450,N_8610,N_8910);
or U9451 (N_9451,N_8576,N_8505);
or U9452 (N_9452,N_8630,N_8638);
nand U9453 (N_9453,N_8673,N_8894);
nor U9454 (N_9454,N_8990,N_8587);
or U9455 (N_9455,N_8692,N_8771);
and U9456 (N_9456,N_8562,N_8998);
nor U9457 (N_9457,N_8716,N_8688);
xor U9458 (N_9458,N_8729,N_8747);
xnor U9459 (N_9459,N_8960,N_8891);
nor U9460 (N_9460,N_8586,N_8894);
nand U9461 (N_9461,N_8634,N_8631);
nor U9462 (N_9462,N_8526,N_8598);
or U9463 (N_9463,N_8853,N_8987);
and U9464 (N_9464,N_8517,N_8704);
or U9465 (N_9465,N_8595,N_8652);
nor U9466 (N_9466,N_8755,N_8722);
and U9467 (N_9467,N_8618,N_8907);
or U9468 (N_9468,N_8772,N_8624);
and U9469 (N_9469,N_8600,N_8885);
or U9470 (N_9470,N_8627,N_8666);
or U9471 (N_9471,N_8532,N_8939);
nand U9472 (N_9472,N_8598,N_8663);
nand U9473 (N_9473,N_8854,N_8747);
or U9474 (N_9474,N_8564,N_8915);
nor U9475 (N_9475,N_8561,N_8801);
and U9476 (N_9476,N_8500,N_8752);
or U9477 (N_9477,N_8772,N_8670);
nor U9478 (N_9478,N_8809,N_8552);
xnor U9479 (N_9479,N_8915,N_8678);
and U9480 (N_9480,N_8695,N_8689);
or U9481 (N_9481,N_8588,N_8543);
nand U9482 (N_9482,N_8988,N_8981);
nor U9483 (N_9483,N_8925,N_8778);
nor U9484 (N_9484,N_8789,N_8779);
nor U9485 (N_9485,N_8786,N_8618);
or U9486 (N_9486,N_8605,N_8625);
nor U9487 (N_9487,N_8546,N_8553);
nor U9488 (N_9488,N_8600,N_8856);
nand U9489 (N_9489,N_8817,N_8811);
nor U9490 (N_9490,N_8677,N_8522);
nor U9491 (N_9491,N_8714,N_8736);
or U9492 (N_9492,N_8952,N_8655);
and U9493 (N_9493,N_8606,N_8567);
nand U9494 (N_9494,N_8721,N_8823);
and U9495 (N_9495,N_8911,N_8713);
and U9496 (N_9496,N_8984,N_8867);
nor U9497 (N_9497,N_8526,N_8844);
nor U9498 (N_9498,N_8839,N_8829);
nand U9499 (N_9499,N_8749,N_8623);
nand U9500 (N_9500,N_9105,N_9466);
nand U9501 (N_9501,N_9184,N_9320);
or U9502 (N_9502,N_9279,N_9432);
or U9503 (N_9503,N_9021,N_9433);
or U9504 (N_9504,N_9296,N_9383);
nor U9505 (N_9505,N_9339,N_9423);
or U9506 (N_9506,N_9262,N_9335);
nand U9507 (N_9507,N_9273,N_9196);
and U9508 (N_9508,N_9133,N_9067);
or U9509 (N_9509,N_9134,N_9309);
and U9510 (N_9510,N_9243,N_9303);
nand U9511 (N_9511,N_9030,N_9493);
or U9512 (N_9512,N_9097,N_9409);
or U9513 (N_9513,N_9122,N_9393);
nor U9514 (N_9514,N_9033,N_9077);
nor U9515 (N_9515,N_9421,N_9463);
or U9516 (N_9516,N_9132,N_9026);
nand U9517 (N_9517,N_9338,N_9149);
nor U9518 (N_9518,N_9252,N_9036);
and U9519 (N_9519,N_9025,N_9424);
nand U9520 (N_9520,N_9152,N_9169);
nand U9521 (N_9521,N_9498,N_9297);
nor U9522 (N_9522,N_9141,N_9478);
nand U9523 (N_9523,N_9354,N_9238);
and U9524 (N_9524,N_9011,N_9101);
nor U9525 (N_9525,N_9391,N_9356);
nand U9526 (N_9526,N_9480,N_9221);
and U9527 (N_9527,N_9427,N_9364);
nor U9528 (N_9528,N_9130,N_9476);
nand U9529 (N_9529,N_9250,N_9107);
nand U9530 (N_9530,N_9345,N_9247);
nand U9531 (N_9531,N_9485,N_9127);
nor U9532 (N_9532,N_9254,N_9298);
nor U9533 (N_9533,N_9363,N_9275);
and U9534 (N_9534,N_9484,N_9435);
and U9535 (N_9535,N_9190,N_9106);
or U9536 (N_9536,N_9379,N_9355);
nand U9537 (N_9537,N_9426,N_9131);
or U9538 (N_9538,N_9136,N_9139);
or U9539 (N_9539,N_9145,N_9199);
and U9540 (N_9540,N_9397,N_9018);
nand U9541 (N_9541,N_9035,N_9471);
nand U9542 (N_9542,N_9209,N_9447);
nor U9543 (N_9543,N_9094,N_9366);
and U9544 (N_9544,N_9392,N_9388);
and U9545 (N_9545,N_9082,N_9038);
and U9546 (N_9546,N_9405,N_9037);
or U9547 (N_9547,N_9472,N_9245);
or U9548 (N_9548,N_9013,N_9231);
nor U9549 (N_9549,N_9182,N_9284);
or U9550 (N_9550,N_9114,N_9009);
nor U9551 (N_9551,N_9088,N_9176);
nor U9552 (N_9552,N_9193,N_9055);
nand U9553 (N_9553,N_9420,N_9099);
nand U9554 (N_9554,N_9234,N_9064);
nand U9555 (N_9555,N_9043,N_9163);
nor U9556 (N_9556,N_9085,N_9179);
nor U9557 (N_9557,N_9161,N_9491);
or U9558 (N_9558,N_9063,N_9201);
or U9559 (N_9559,N_9357,N_9416);
or U9560 (N_9560,N_9398,N_9007);
and U9561 (N_9561,N_9189,N_9028);
or U9562 (N_9562,N_9352,N_9168);
and U9563 (N_9563,N_9039,N_9041);
nand U9564 (N_9564,N_9171,N_9386);
nor U9565 (N_9565,N_9422,N_9124);
nand U9566 (N_9566,N_9080,N_9151);
or U9567 (N_9567,N_9429,N_9205);
or U9568 (N_9568,N_9256,N_9289);
or U9569 (N_9569,N_9265,N_9206);
or U9570 (N_9570,N_9116,N_9058);
xor U9571 (N_9571,N_9321,N_9396);
nor U9572 (N_9572,N_9075,N_9344);
or U9573 (N_9573,N_9170,N_9316);
xor U9574 (N_9574,N_9081,N_9479);
nor U9575 (N_9575,N_9291,N_9071);
nor U9576 (N_9576,N_9327,N_9411);
nor U9577 (N_9577,N_9306,N_9470);
or U9578 (N_9578,N_9283,N_9331);
nand U9579 (N_9579,N_9192,N_9436);
and U9580 (N_9580,N_9312,N_9109);
or U9581 (N_9581,N_9126,N_9008);
and U9582 (N_9582,N_9380,N_9328);
and U9583 (N_9583,N_9230,N_9207);
or U9584 (N_9584,N_9223,N_9147);
nand U9585 (N_9585,N_9314,N_9117);
or U9586 (N_9586,N_9015,N_9334);
and U9587 (N_9587,N_9438,N_9072);
and U9588 (N_9588,N_9084,N_9437);
and U9589 (N_9589,N_9271,N_9294);
and U9590 (N_9590,N_9371,N_9146);
nand U9591 (N_9591,N_9195,N_9227);
and U9592 (N_9592,N_9244,N_9374);
or U9593 (N_9593,N_9459,N_9128);
nor U9594 (N_9594,N_9369,N_9166);
and U9595 (N_9595,N_9157,N_9496);
and U9596 (N_9596,N_9029,N_9135);
nand U9597 (N_9597,N_9104,N_9083);
or U9598 (N_9598,N_9290,N_9341);
nor U9599 (N_9599,N_9482,N_9158);
or U9600 (N_9600,N_9382,N_9465);
nor U9601 (N_9601,N_9185,N_9242);
and U9602 (N_9602,N_9113,N_9311);
or U9603 (N_9603,N_9346,N_9300);
nand U9604 (N_9604,N_9457,N_9213);
and U9605 (N_9605,N_9248,N_9458);
or U9606 (N_9606,N_9415,N_9110);
and U9607 (N_9607,N_9065,N_9093);
nor U9608 (N_9608,N_9045,N_9073);
nor U9609 (N_9609,N_9180,N_9211);
nor U9610 (N_9610,N_9164,N_9014);
or U9611 (N_9611,N_9467,N_9302);
nand U9612 (N_9612,N_9020,N_9385);
nand U9613 (N_9613,N_9389,N_9486);
or U9614 (N_9614,N_9129,N_9317);
nor U9615 (N_9615,N_9236,N_9270);
nor U9616 (N_9616,N_9160,N_9413);
nor U9617 (N_9617,N_9016,N_9068);
and U9618 (N_9618,N_9006,N_9191);
nand U9619 (N_9619,N_9024,N_9431);
and U9620 (N_9620,N_9325,N_9174);
nand U9621 (N_9621,N_9451,N_9017);
nor U9622 (N_9622,N_9367,N_9208);
nand U9623 (N_9623,N_9225,N_9483);
and U9624 (N_9624,N_9142,N_9153);
or U9625 (N_9625,N_9333,N_9137);
and U9626 (N_9626,N_9468,N_9313);
nor U9627 (N_9627,N_9140,N_9258);
nand U9628 (N_9628,N_9469,N_9443);
or U9629 (N_9629,N_9010,N_9378);
or U9630 (N_9630,N_9299,N_9100);
and U9631 (N_9631,N_9375,N_9488);
nand U9632 (N_9632,N_9319,N_9220);
and U9633 (N_9633,N_9454,N_9102);
or U9634 (N_9634,N_9342,N_9499);
nor U9635 (N_9635,N_9418,N_9237);
or U9636 (N_9636,N_9439,N_9349);
or U9637 (N_9637,N_9069,N_9044);
and U9638 (N_9638,N_9387,N_9059);
nor U9639 (N_9639,N_9376,N_9054);
or U9640 (N_9640,N_9188,N_9074);
nor U9641 (N_9641,N_9359,N_9241);
nand U9642 (N_9642,N_9475,N_9172);
nor U9643 (N_9643,N_9155,N_9125);
and U9644 (N_9644,N_9060,N_9365);
nor U9645 (N_9645,N_9259,N_9143);
nor U9646 (N_9646,N_9086,N_9138);
nor U9647 (N_9647,N_9453,N_9204);
or U9648 (N_9648,N_9358,N_9285);
nand U9649 (N_9649,N_9308,N_9473);
nor U9650 (N_9650,N_9148,N_9490);
nor U9651 (N_9651,N_9032,N_9156);
nor U9652 (N_9652,N_9048,N_9034);
nor U9653 (N_9653,N_9202,N_9090);
nor U9654 (N_9654,N_9047,N_9162);
nand U9655 (N_9655,N_9005,N_9348);
nand U9656 (N_9656,N_9360,N_9425);
nor U9657 (N_9657,N_9448,N_9159);
nand U9658 (N_9658,N_9061,N_9347);
nand U9659 (N_9659,N_9350,N_9450);
and U9660 (N_9660,N_9003,N_9278);
or U9661 (N_9661,N_9261,N_9257);
and U9662 (N_9662,N_9052,N_9251);
and U9663 (N_9663,N_9144,N_9089);
or U9664 (N_9664,N_9178,N_9362);
or U9665 (N_9665,N_9304,N_9353);
or U9666 (N_9666,N_9210,N_9440);
or U9667 (N_9667,N_9315,N_9264);
or U9668 (N_9668,N_9194,N_9004);
xnor U9669 (N_9669,N_9268,N_9217);
nand U9670 (N_9670,N_9407,N_9332);
or U9671 (N_9671,N_9049,N_9070);
nand U9672 (N_9672,N_9098,N_9076);
or U9673 (N_9673,N_9377,N_9461);
nand U9674 (N_9674,N_9286,N_9400);
nand U9675 (N_9675,N_9489,N_9287);
or U9676 (N_9676,N_9492,N_9428);
and U9677 (N_9677,N_9119,N_9233);
or U9678 (N_9678,N_9305,N_9408);
nor U9679 (N_9679,N_9118,N_9295);
or U9680 (N_9680,N_9023,N_9318);
or U9681 (N_9681,N_9343,N_9430);
nand U9682 (N_9682,N_9307,N_9121);
nand U9683 (N_9683,N_9460,N_9051);
xor U9684 (N_9684,N_9456,N_9095);
or U9685 (N_9685,N_9120,N_9477);
nand U9686 (N_9686,N_9449,N_9226);
and U9687 (N_9687,N_9372,N_9246);
nand U9688 (N_9688,N_9370,N_9404);
nand U9689 (N_9689,N_9173,N_9310);
nor U9690 (N_9690,N_9249,N_9288);
and U9691 (N_9691,N_9228,N_9481);
nor U9692 (N_9692,N_9495,N_9103);
or U9693 (N_9693,N_9002,N_9464);
or U9694 (N_9694,N_9012,N_9445);
and U9695 (N_9695,N_9027,N_9175);
nor U9696 (N_9696,N_9000,N_9019);
or U9697 (N_9697,N_9001,N_9402);
nor U9698 (N_9698,N_9212,N_9022);
or U9699 (N_9699,N_9293,N_9269);
nor U9700 (N_9700,N_9232,N_9455);
nor U9701 (N_9701,N_9292,N_9337);
nor U9702 (N_9702,N_9394,N_9263);
nor U9703 (N_9703,N_9446,N_9487);
nand U9704 (N_9704,N_9336,N_9066);
and U9705 (N_9705,N_9253,N_9218);
nor U9706 (N_9706,N_9274,N_9260);
nor U9707 (N_9707,N_9096,N_9167);
nand U9708 (N_9708,N_9462,N_9046);
or U9709 (N_9709,N_9200,N_9277);
xor U9710 (N_9710,N_9031,N_9497);
or U9711 (N_9711,N_9414,N_9267);
nand U9712 (N_9712,N_9150,N_9324);
or U9713 (N_9713,N_9123,N_9239);
nor U9714 (N_9714,N_9087,N_9474);
or U9715 (N_9715,N_9406,N_9078);
or U9716 (N_9716,N_9272,N_9111);
and U9717 (N_9717,N_9494,N_9419);
nor U9718 (N_9718,N_9390,N_9255);
nand U9719 (N_9719,N_9444,N_9057);
and U9720 (N_9720,N_9216,N_9042);
xnor U9721 (N_9721,N_9224,N_9301);
or U9722 (N_9722,N_9115,N_9053);
nor U9723 (N_9723,N_9410,N_9229);
and U9724 (N_9724,N_9340,N_9197);
and U9725 (N_9725,N_9282,N_9280);
nor U9726 (N_9726,N_9154,N_9351);
or U9727 (N_9727,N_9403,N_9203);
or U9728 (N_9728,N_9441,N_9091);
and U9729 (N_9729,N_9399,N_9381);
nor U9730 (N_9730,N_9395,N_9281);
nor U9731 (N_9731,N_9417,N_9215);
and U9732 (N_9732,N_9442,N_9276);
or U9733 (N_9733,N_9326,N_9183);
nor U9734 (N_9734,N_9177,N_9368);
nor U9735 (N_9735,N_9112,N_9434);
nor U9736 (N_9736,N_9401,N_9050);
and U9737 (N_9737,N_9187,N_9373);
or U9738 (N_9738,N_9452,N_9219);
nand U9739 (N_9739,N_9240,N_9079);
and U9740 (N_9740,N_9108,N_9222);
nand U9741 (N_9741,N_9092,N_9181);
xor U9742 (N_9742,N_9361,N_9040);
and U9743 (N_9743,N_9198,N_9323);
nor U9744 (N_9744,N_9165,N_9266);
and U9745 (N_9745,N_9329,N_9214);
nand U9746 (N_9746,N_9322,N_9056);
and U9747 (N_9747,N_9384,N_9235);
nor U9748 (N_9748,N_9062,N_9186);
nor U9749 (N_9749,N_9412,N_9330);
or U9750 (N_9750,N_9063,N_9116);
nand U9751 (N_9751,N_9042,N_9093);
nor U9752 (N_9752,N_9400,N_9461);
or U9753 (N_9753,N_9463,N_9032);
and U9754 (N_9754,N_9439,N_9025);
and U9755 (N_9755,N_9345,N_9369);
or U9756 (N_9756,N_9186,N_9033);
and U9757 (N_9757,N_9475,N_9278);
nor U9758 (N_9758,N_9089,N_9341);
or U9759 (N_9759,N_9004,N_9099);
and U9760 (N_9760,N_9053,N_9255);
or U9761 (N_9761,N_9089,N_9215);
nor U9762 (N_9762,N_9292,N_9133);
nand U9763 (N_9763,N_9482,N_9201);
and U9764 (N_9764,N_9386,N_9076);
and U9765 (N_9765,N_9327,N_9276);
or U9766 (N_9766,N_9430,N_9038);
or U9767 (N_9767,N_9123,N_9268);
nand U9768 (N_9768,N_9074,N_9195);
nand U9769 (N_9769,N_9226,N_9317);
and U9770 (N_9770,N_9317,N_9334);
and U9771 (N_9771,N_9040,N_9157);
nand U9772 (N_9772,N_9126,N_9000);
or U9773 (N_9773,N_9139,N_9070);
and U9774 (N_9774,N_9182,N_9392);
nand U9775 (N_9775,N_9252,N_9492);
nor U9776 (N_9776,N_9049,N_9190);
nor U9777 (N_9777,N_9158,N_9163);
nand U9778 (N_9778,N_9399,N_9364);
or U9779 (N_9779,N_9487,N_9294);
nor U9780 (N_9780,N_9310,N_9359);
xnor U9781 (N_9781,N_9402,N_9306);
nor U9782 (N_9782,N_9120,N_9085);
and U9783 (N_9783,N_9180,N_9143);
nor U9784 (N_9784,N_9283,N_9494);
and U9785 (N_9785,N_9199,N_9429);
xor U9786 (N_9786,N_9190,N_9091);
nand U9787 (N_9787,N_9164,N_9089);
and U9788 (N_9788,N_9071,N_9321);
nor U9789 (N_9789,N_9356,N_9411);
or U9790 (N_9790,N_9054,N_9152);
nor U9791 (N_9791,N_9396,N_9101);
nor U9792 (N_9792,N_9151,N_9272);
nor U9793 (N_9793,N_9144,N_9072);
or U9794 (N_9794,N_9011,N_9137);
and U9795 (N_9795,N_9203,N_9126);
nor U9796 (N_9796,N_9211,N_9226);
nand U9797 (N_9797,N_9065,N_9154);
nand U9798 (N_9798,N_9157,N_9472);
or U9799 (N_9799,N_9212,N_9450);
or U9800 (N_9800,N_9133,N_9267);
and U9801 (N_9801,N_9087,N_9111);
or U9802 (N_9802,N_9001,N_9369);
nand U9803 (N_9803,N_9365,N_9064);
and U9804 (N_9804,N_9022,N_9065);
and U9805 (N_9805,N_9093,N_9116);
and U9806 (N_9806,N_9181,N_9013);
and U9807 (N_9807,N_9256,N_9358);
nand U9808 (N_9808,N_9296,N_9326);
nor U9809 (N_9809,N_9395,N_9116);
nor U9810 (N_9810,N_9283,N_9244);
nand U9811 (N_9811,N_9236,N_9419);
xor U9812 (N_9812,N_9032,N_9038);
or U9813 (N_9813,N_9080,N_9037);
nor U9814 (N_9814,N_9317,N_9131);
or U9815 (N_9815,N_9468,N_9205);
and U9816 (N_9816,N_9101,N_9224);
nand U9817 (N_9817,N_9002,N_9490);
nor U9818 (N_9818,N_9349,N_9084);
nor U9819 (N_9819,N_9146,N_9261);
and U9820 (N_9820,N_9207,N_9105);
or U9821 (N_9821,N_9008,N_9317);
nand U9822 (N_9822,N_9365,N_9261);
nand U9823 (N_9823,N_9102,N_9142);
or U9824 (N_9824,N_9171,N_9491);
nand U9825 (N_9825,N_9016,N_9354);
nand U9826 (N_9826,N_9318,N_9195);
nand U9827 (N_9827,N_9299,N_9312);
nor U9828 (N_9828,N_9155,N_9499);
and U9829 (N_9829,N_9462,N_9225);
nand U9830 (N_9830,N_9481,N_9157);
and U9831 (N_9831,N_9252,N_9084);
nand U9832 (N_9832,N_9073,N_9118);
nand U9833 (N_9833,N_9339,N_9182);
and U9834 (N_9834,N_9434,N_9208);
nor U9835 (N_9835,N_9345,N_9254);
nand U9836 (N_9836,N_9051,N_9124);
and U9837 (N_9837,N_9287,N_9152);
nor U9838 (N_9838,N_9444,N_9278);
or U9839 (N_9839,N_9245,N_9478);
nor U9840 (N_9840,N_9040,N_9462);
nand U9841 (N_9841,N_9121,N_9368);
nand U9842 (N_9842,N_9318,N_9055);
and U9843 (N_9843,N_9460,N_9255);
and U9844 (N_9844,N_9377,N_9366);
nand U9845 (N_9845,N_9219,N_9111);
nand U9846 (N_9846,N_9478,N_9265);
and U9847 (N_9847,N_9143,N_9484);
xnor U9848 (N_9848,N_9024,N_9038);
nand U9849 (N_9849,N_9444,N_9355);
and U9850 (N_9850,N_9386,N_9292);
nor U9851 (N_9851,N_9092,N_9192);
nor U9852 (N_9852,N_9426,N_9477);
nand U9853 (N_9853,N_9169,N_9168);
and U9854 (N_9854,N_9176,N_9463);
nand U9855 (N_9855,N_9272,N_9226);
or U9856 (N_9856,N_9447,N_9286);
nor U9857 (N_9857,N_9353,N_9293);
or U9858 (N_9858,N_9381,N_9004);
nand U9859 (N_9859,N_9283,N_9326);
or U9860 (N_9860,N_9481,N_9065);
or U9861 (N_9861,N_9474,N_9279);
nand U9862 (N_9862,N_9352,N_9235);
nand U9863 (N_9863,N_9004,N_9009);
and U9864 (N_9864,N_9324,N_9018);
and U9865 (N_9865,N_9067,N_9369);
or U9866 (N_9866,N_9104,N_9034);
xor U9867 (N_9867,N_9433,N_9256);
nand U9868 (N_9868,N_9437,N_9480);
nand U9869 (N_9869,N_9194,N_9134);
and U9870 (N_9870,N_9499,N_9470);
nor U9871 (N_9871,N_9463,N_9002);
nor U9872 (N_9872,N_9171,N_9066);
nand U9873 (N_9873,N_9341,N_9426);
and U9874 (N_9874,N_9009,N_9310);
or U9875 (N_9875,N_9155,N_9337);
nor U9876 (N_9876,N_9327,N_9144);
nand U9877 (N_9877,N_9298,N_9269);
nand U9878 (N_9878,N_9370,N_9273);
and U9879 (N_9879,N_9019,N_9203);
nor U9880 (N_9880,N_9209,N_9456);
nor U9881 (N_9881,N_9498,N_9484);
nor U9882 (N_9882,N_9381,N_9451);
or U9883 (N_9883,N_9367,N_9194);
nor U9884 (N_9884,N_9176,N_9468);
nand U9885 (N_9885,N_9027,N_9455);
or U9886 (N_9886,N_9202,N_9441);
nor U9887 (N_9887,N_9484,N_9042);
nor U9888 (N_9888,N_9186,N_9240);
and U9889 (N_9889,N_9037,N_9038);
or U9890 (N_9890,N_9216,N_9118);
nor U9891 (N_9891,N_9468,N_9082);
nor U9892 (N_9892,N_9172,N_9294);
and U9893 (N_9893,N_9448,N_9128);
or U9894 (N_9894,N_9131,N_9412);
or U9895 (N_9895,N_9166,N_9167);
nand U9896 (N_9896,N_9094,N_9175);
and U9897 (N_9897,N_9102,N_9339);
and U9898 (N_9898,N_9177,N_9324);
nor U9899 (N_9899,N_9095,N_9357);
nor U9900 (N_9900,N_9183,N_9221);
nor U9901 (N_9901,N_9129,N_9078);
nand U9902 (N_9902,N_9400,N_9303);
or U9903 (N_9903,N_9136,N_9455);
nand U9904 (N_9904,N_9315,N_9229);
nor U9905 (N_9905,N_9152,N_9319);
and U9906 (N_9906,N_9175,N_9111);
nand U9907 (N_9907,N_9269,N_9494);
nand U9908 (N_9908,N_9387,N_9414);
and U9909 (N_9909,N_9009,N_9100);
and U9910 (N_9910,N_9111,N_9156);
nand U9911 (N_9911,N_9306,N_9395);
nand U9912 (N_9912,N_9264,N_9035);
and U9913 (N_9913,N_9482,N_9043);
xor U9914 (N_9914,N_9124,N_9228);
nand U9915 (N_9915,N_9391,N_9197);
or U9916 (N_9916,N_9264,N_9236);
or U9917 (N_9917,N_9126,N_9048);
or U9918 (N_9918,N_9474,N_9053);
or U9919 (N_9919,N_9186,N_9200);
nand U9920 (N_9920,N_9279,N_9186);
and U9921 (N_9921,N_9219,N_9107);
and U9922 (N_9922,N_9486,N_9236);
or U9923 (N_9923,N_9306,N_9062);
or U9924 (N_9924,N_9352,N_9111);
nor U9925 (N_9925,N_9143,N_9415);
nand U9926 (N_9926,N_9310,N_9484);
nand U9927 (N_9927,N_9417,N_9030);
and U9928 (N_9928,N_9069,N_9201);
and U9929 (N_9929,N_9328,N_9133);
and U9930 (N_9930,N_9386,N_9159);
or U9931 (N_9931,N_9027,N_9379);
nand U9932 (N_9932,N_9249,N_9278);
nand U9933 (N_9933,N_9400,N_9448);
and U9934 (N_9934,N_9360,N_9064);
or U9935 (N_9935,N_9280,N_9391);
and U9936 (N_9936,N_9110,N_9210);
nand U9937 (N_9937,N_9136,N_9080);
nand U9938 (N_9938,N_9286,N_9022);
or U9939 (N_9939,N_9150,N_9249);
nor U9940 (N_9940,N_9268,N_9260);
or U9941 (N_9941,N_9211,N_9354);
xnor U9942 (N_9942,N_9221,N_9283);
xor U9943 (N_9943,N_9358,N_9400);
or U9944 (N_9944,N_9398,N_9045);
and U9945 (N_9945,N_9293,N_9208);
nor U9946 (N_9946,N_9309,N_9443);
and U9947 (N_9947,N_9019,N_9274);
nand U9948 (N_9948,N_9386,N_9194);
or U9949 (N_9949,N_9182,N_9145);
nor U9950 (N_9950,N_9431,N_9067);
nor U9951 (N_9951,N_9228,N_9445);
nor U9952 (N_9952,N_9405,N_9220);
nand U9953 (N_9953,N_9120,N_9142);
and U9954 (N_9954,N_9194,N_9411);
xnor U9955 (N_9955,N_9365,N_9233);
xor U9956 (N_9956,N_9003,N_9127);
or U9957 (N_9957,N_9460,N_9116);
or U9958 (N_9958,N_9479,N_9390);
and U9959 (N_9959,N_9078,N_9442);
and U9960 (N_9960,N_9249,N_9049);
and U9961 (N_9961,N_9404,N_9186);
or U9962 (N_9962,N_9318,N_9096);
and U9963 (N_9963,N_9125,N_9476);
and U9964 (N_9964,N_9174,N_9008);
nor U9965 (N_9965,N_9204,N_9282);
and U9966 (N_9966,N_9453,N_9111);
nor U9967 (N_9967,N_9124,N_9497);
or U9968 (N_9968,N_9295,N_9187);
or U9969 (N_9969,N_9307,N_9048);
nand U9970 (N_9970,N_9400,N_9447);
nor U9971 (N_9971,N_9373,N_9169);
and U9972 (N_9972,N_9163,N_9272);
nand U9973 (N_9973,N_9482,N_9016);
nand U9974 (N_9974,N_9177,N_9064);
nand U9975 (N_9975,N_9081,N_9238);
nor U9976 (N_9976,N_9283,N_9185);
or U9977 (N_9977,N_9199,N_9329);
nor U9978 (N_9978,N_9075,N_9009);
and U9979 (N_9979,N_9116,N_9440);
and U9980 (N_9980,N_9171,N_9387);
or U9981 (N_9981,N_9072,N_9123);
or U9982 (N_9982,N_9292,N_9150);
and U9983 (N_9983,N_9298,N_9425);
nor U9984 (N_9984,N_9323,N_9054);
nand U9985 (N_9985,N_9087,N_9414);
or U9986 (N_9986,N_9044,N_9445);
or U9987 (N_9987,N_9344,N_9331);
nand U9988 (N_9988,N_9315,N_9452);
nor U9989 (N_9989,N_9426,N_9421);
nor U9990 (N_9990,N_9321,N_9108);
and U9991 (N_9991,N_9341,N_9449);
or U9992 (N_9992,N_9356,N_9461);
or U9993 (N_9993,N_9341,N_9313);
or U9994 (N_9994,N_9154,N_9410);
or U9995 (N_9995,N_9076,N_9475);
and U9996 (N_9996,N_9243,N_9335);
and U9997 (N_9997,N_9350,N_9188);
nor U9998 (N_9998,N_9100,N_9094);
nor U9999 (N_9999,N_9255,N_9413);
nand U10000 (N_10000,N_9718,N_9608);
nor U10001 (N_10001,N_9980,N_9559);
nor U10002 (N_10002,N_9902,N_9536);
nor U10003 (N_10003,N_9794,N_9522);
and U10004 (N_10004,N_9564,N_9929);
or U10005 (N_10005,N_9835,N_9747);
and U10006 (N_10006,N_9948,N_9978);
nor U10007 (N_10007,N_9821,N_9971);
nor U10008 (N_10008,N_9828,N_9659);
and U10009 (N_10009,N_9903,N_9745);
and U10010 (N_10010,N_9735,N_9531);
and U10011 (N_10011,N_9734,N_9969);
or U10012 (N_10012,N_9778,N_9644);
or U10013 (N_10013,N_9693,N_9962);
nor U10014 (N_10014,N_9733,N_9934);
nand U10015 (N_10015,N_9710,N_9918);
or U10016 (N_10016,N_9993,N_9761);
nor U10017 (N_10017,N_9753,N_9612);
and U10018 (N_10018,N_9864,N_9613);
and U10019 (N_10019,N_9807,N_9770);
nand U10020 (N_10020,N_9860,N_9744);
nor U10021 (N_10021,N_9558,N_9580);
nand U10022 (N_10022,N_9957,N_9758);
nor U10023 (N_10023,N_9703,N_9822);
or U10024 (N_10024,N_9781,N_9690);
xnor U10025 (N_10025,N_9931,N_9808);
nand U10026 (N_10026,N_9731,N_9856);
nor U10027 (N_10027,N_9803,N_9512);
nor U10028 (N_10028,N_9910,N_9595);
nand U10029 (N_10029,N_9721,N_9867);
or U10030 (N_10030,N_9941,N_9937);
and U10031 (N_10031,N_9886,N_9581);
or U10032 (N_10032,N_9709,N_9795);
nor U10033 (N_10033,N_9513,N_9707);
nor U10034 (N_10034,N_9945,N_9812);
nand U10035 (N_10035,N_9774,N_9639);
and U10036 (N_10036,N_9650,N_9930);
and U10037 (N_10037,N_9911,N_9848);
or U10038 (N_10038,N_9515,N_9858);
and U10039 (N_10039,N_9798,N_9928);
and U10040 (N_10040,N_9590,N_9868);
nor U10041 (N_10041,N_9925,N_9916);
nand U10042 (N_10042,N_9763,N_9742);
and U10043 (N_10043,N_9722,N_9637);
and U10044 (N_10044,N_9765,N_9533);
and U10045 (N_10045,N_9702,N_9626);
or U10046 (N_10046,N_9643,N_9524);
nor U10047 (N_10047,N_9965,N_9769);
nand U10048 (N_10048,N_9802,N_9907);
nor U10049 (N_10049,N_9668,N_9529);
nand U10050 (N_10050,N_9509,N_9849);
or U10051 (N_10051,N_9615,N_9727);
or U10052 (N_10052,N_9566,N_9815);
nand U10053 (N_10053,N_9764,N_9783);
nand U10054 (N_10054,N_9501,N_9576);
and U10055 (N_10055,N_9839,N_9726);
and U10056 (N_10056,N_9625,N_9920);
and U10057 (N_10057,N_9573,N_9751);
nor U10058 (N_10058,N_9572,N_9938);
nand U10059 (N_10059,N_9593,N_9646);
nand U10060 (N_10060,N_9972,N_9953);
nand U10061 (N_10061,N_9997,N_9888);
and U10062 (N_10062,N_9989,N_9852);
or U10063 (N_10063,N_9670,N_9956);
and U10064 (N_10064,N_9843,N_9904);
nand U10065 (N_10065,N_9627,N_9649);
and U10066 (N_10066,N_9561,N_9960);
and U10067 (N_10067,N_9876,N_9741);
nand U10068 (N_10068,N_9568,N_9699);
nand U10069 (N_10069,N_9725,N_9569);
and U10070 (N_10070,N_9716,N_9708);
or U10071 (N_10071,N_9618,N_9805);
and U10072 (N_10072,N_9688,N_9660);
nor U10073 (N_10073,N_9811,N_9676);
and U10074 (N_10074,N_9819,N_9933);
nor U10075 (N_10075,N_9617,N_9674);
nor U10076 (N_10076,N_9678,N_9793);
xor U10077 (N_10077,N_9611,N_9991);
and U10078 (N_10078,N_9782,N_9662);
nand U10079 (N_10079,N_9840,N_9584);
nand U10080 (N_10080,N_9954,N_9825);
nand U10081 (N_10081,N_9691,N_9963);
nor U10082 (N_10082,N_9766,N_9588);
nor U10083 (N_10083,N_9817,N_9653);
and U10084 (N_10084,N_9983,N_9975);
nor U10085 (N_10085,N_9877,N_9999);
or U10086 (N_10086,N_9966,N_9899);
or U10087 (N_10087,N_9586,N_9942);
and U10088 (N_10088,N_9525,N_9939);
nor U10089 (N_10089,N_9974,N_9909);
and U10090 (N_10090,N_9689,N_9979);
nor U10091 (N_10091,N_9892,N_9647);
nand U10092 (N_10092,N_9996,N_9535);
nand U10093 (N_10093,N_9671,N_9679);
and U10094 (N_10094,N_9698,N_9508);
and U10095 (N_10095,N_9829,N_9986);
nand U10096 (N_10096,N_9816,N_9771);
or U10097 (N_10097,N_9833,N_9597);
nand U10098 (N_10098,N_9885,N_9516);
and U10099 (N_10099,N_9832,N_9838);
or U10100 (N_10100,N_9567,N_9896);
nor U10101 (N_10101,N_9655,N_9984);
nor U10102 (N_10102,N_9820,N_9701);
nor U10103 (N_10103,N_9505,N_9680);
nand U10104 (N_10104,N_9717,N_9589);
nor U10105 (N_10105,N_9830,N_9579);
nor U10106 (N_10106,N_9882,N_9756);
or U10107 (N_10107,N_9517,N_9792);
nand U10108 (N_10108,N_9503,N_9967);
nand U10109 (N_10109,N_9622,N_9988);
and U10110 (N_10110,N_9661,N_9874);
nor U10111 (N_10111,N_9720,N_9504);
nand U10112 (N_10112,N_9634,N_9827);
nor U10113 (N_10113,N_9872,N_9906);
and U10114 (N_10114,N_9800,N_9801);
or U10115 (N_10115,N_9601,N_9797);
nor U10116 (N_10116,N_9638,N_9880);
nor U10117 (N_10117,N_9528,N_9694);
nand U10118 (N_10118,N_9842,N_9631);
nor U10119 (N_10119,N_9736,N_9648);
or U10120 (N_10120,N_9636,N_9729);
xor U10121 (N_10121,N_9895,N_9606);
xnor U10122 (N_10122,N_9544,N_9550);
or U10123 (N_10123,N_9549,N_9824);
and U10124 (N_10124,N_9784,N_9511);
nor U10125 (N_10125,N_9871,N_9844);
or U10126 (N_10126,N_9554,N_9813);
or U10127 (N_10127,N_9705,N_9681);
and U10128 (N_10128,N_9624,N_9776);
nor U10129 (N_10129,N_9878,N_9796);
and U10130 (N_10130,N_9905,N_9632);
or U10131 (N_10131,N_9697,N_9869);
and U10132 (N_10132,N_9754,N_9917);
or U10133 (N_10133,N_9919,N_9587);
and U10134 (N_10134,N_9667,N_9913);
nor U10135 (N_10135,N_9946,N_9943);
or U10136 (N_10136,N_9675,N_9894);
nand U10137 (N_10137,N_9599,N_9514);
and U10138 (N_10138,N_9686,N_9542);
or U10139 (N_10139,N_9773,N_9540);
nor U10140 (N_10140,N_9510,N_9865);
nand U10141 (N_10141,N_9951,N_9621);
nand U10142 (N_10142,N_9949,N_9940);
nor U10143 (N_10143,N_9633,N_9994);
and U10144 (N_10144,N_9565,N_9804);
and U10145 (N_10145,N_9610,N_9932);
or U10146 (N_10146,N_9926,N_9788);
or U10147 (N_10147,N_9651,N_9787);
and U10148 (N_10148,N_9523,N_9563);
and U10149 (N_10149,N_9887,N_9982);
nand U10150 (N_10150,N_9538,N_9604);
nor U10151 (N_10151,N_9924,N_9746);
or U10152 (N_10152,N_9921,N_9959);
nor U10153 (N_10153,N_9645,N_9507);
nand U10154 (N_10154,N_9737,N_9657);
and U10155 (N_10155,N_9623,N_9981);
nand U10156 (N_10156,N_9866,N_9518);
nand U10157 (N_10157,N_9749,N_9711);
nand U10158 (N_10158,N_9723,N_9958);
nor U10159 (N_10159,N_9809,N_9799);
or U10160 (N_10160,N_9665,N_9692);
nand U10161 (N_10161,N_9552,N_9609);
and U10162 (N_10162,N_9810,N_9775);
and U10163 (N_10163,N_9786,N_9873);
or U10164 (N_10164,N_9891,N_9944);
xor U10165 (N_10165,N_9952,N_9673);
and U10166 (N_10166,N_9582,N_9598);
and U10167 (N_10167,N_9641,N_9664);
nor U10168 (N_10168,N_9682,N_9927);
nand U10169 (N_10169,N_9998,N_9577);
nand U10170 (N_10170,N_9669,N_9592);
nand U10171 (N_10171,N_9846,N_9575);
nand U10172 (N_10172,N_9527,N_9826);
and U10173 (N_10173,N_9719,N_9700);
nor U10174 (N_10174,N_9837,N_9672);
nand U10175 (N_10175,N_9539,N_9687);
and U10176 (N_10176,N_9976,N_9897);
nand U10177 (N_10177,N_9912,N_9574);
and U10178 (N_10178,N_9831,N_9578);
nand U10179 (N_10179,N_9857,N_9502);
or U10180 (N_10180,N_9875,N_9859);
or U10181 (N_10181,N_9603,N_9922);
nor U10182 (N_10182,N_9521,N_9654);
and U10183 (N_10183,N_9964,N_9543);
nor U10184 (N_10184,N_9847,N_9546);
nor U10185 (N_10185,N_9755,N_9740);
and U10186 (N_10186,N_9914,N_9743);
nand U10187 (N_10187,N_9530,N_9936);
nand U10188 (N_10188,N_9684,N_9884);
nand U10189 (N_10189,N_9855,N_9663);
nor U10190 (N_10190,N_9898,N_9834);
and U10191 (N_10191,N_9750,N_9630);
nand U10192 (N_10192,N_9712,N_9893);
and U10193 (N_10193,N_9519,N_9570);
nor U10194 (N_10194,N_9652,N_9724);
and U10195 (N_10195,N_9841,N_9500);
nand U10196 (N_10196,N_9973,N_9616);
nor U10197 (N_10197,N_9987,N_9704);
or U10198 (N_10198,N_9985,N_9977);
and U10199 (N_10199,N_9950,N_9814);
nor U10200 (N_10200,N_9594,N_9789);
and U10201 (N_10201,N_9555,N_9551);
nand U10202 (N_10202,N_9541,N_9779);
and U10203 (N_10203,N_9583,N_9714);
and U10204 (N_10204,N_9683,N_9970);
nand U10205 (N_10205,N_9547,N_9995);
nand U10206 (N_10206,N_9879,N_9619);
nor U10207 (N_10207,N_9772,N_9602);
and U10208 (N_10208,N_9635,N_9889);
nor U10209 (N_10209,N_9767,N_9526);
nor U10210 (N_10210,N_9900,N_9656);
or U10211 (N_10211,N_9908,N_9629);
and U10212 (N_10212,N_9915,N_9628);
nor U10213 (N_10213,N_9677,N_9780);
and U10214 (N_10214,N_9706,N_9861);
or U10215 (N_10215,N_9658,N_9968);
nor U10216 (N_10216,N_9640,N_9738);
nor U10217 (N_10217,N_9537,N_9881);
nor U10218 (N_10218,N_9560,N_9666);
nand U10219 (N_10219,N_9520,N_9768);
or U10220 (N_10220,N_9863,N_9728);
and U10221 (N_10221,N_9935,N_9961);
and U10222 (N_10222,N_9823,N_9556);
nand U10223 (N_10223,N_9748,N_9854);
or U10224 (N_10224,N_9752,N_9732);
nor U10225 (N_10225,N_9553,N_9818);
nor U10226 (N_10226,N_9990,N_9992);
nor U10227 (N_10227,N_9545,N_9685);
xor U10228 (N_10228,N_9600,N_9790);
nand U10229 (N_10229,N_9695,N_9901);
nand U10230 (N_10230,N_9923,N_9713);
nand U10231 (N_10231,N_9883,N_9620);
nor U10232 (N_10232,N_9850,N_9506);
nor U10233 (N_10233,N_9947,N_9605);
or U10234 (N_10234,N_9596,N_9532);
or U10235 (N_10235,N_9762,N_9851);
nand U10236 (N_10236,N_9862,N_9548);
and U10237 (N_10237,N_9557,N_9845);
or U10238 (N_10238,N_9785,N_9870);
nand U10239 (N_10239,N_9571,N_9614);
nor U10240 (N_10240,N_9757,N_9760);
or U10241 (N_10241,N_9715,N_9534);
nor U10242 (N_10242,N_9890,N_9777);
or U10243 (N_10243,N_9955,N_9836);
or U10244 (N_10244,N_9696,N_9730);
and U10245 (N_10245,N_9759,N_9585);
xnor U10246 (N_10246,N_9642,N_9591);
nand U10247 (N_10247,N_9562,N_9607);
nor U10248 (N_10248,N_9806,N_9791);
and U10249 (N_10249,N_9853,N_9739);
nor U10250 (N_10250,N_9731,N_9930);
nand U10251 (N_10251,N_9984,N_9891);
or U10252 (N_10252,N_9770,N_9797);
or U10253 (N_10253,N_9736,N_9832);
nand U10254 (N_10254,N_9538,N_9686);
and U10255 (N_10255,N_9679,N_9654);
or U10256 (N_10256,N_9740,N_9936);
and U10257 (N_10257,N_9711,N_9913);
nand U10258 (N_10258,N_9952,N_9594);
and U10259 (N_10259,N_9850,N_9575);
xnor U10260 (N_10260,N_9587,N_9529);
and U10261 (N_10261,N_9795,N_9712);
nor U10262 (N_10262,N_9824,N_9570);
or U10263 (N_10263,N_9841,N_9921);
nor U10264 (N_10264,N_9500,N_9816);
and U10265 (N_10265,N_9925,N_9966);
or U10266 (N_10266,N_9828,N_9634);
or U10267 (N_10267,N_9930,N_9831);
nor U10268 (N_10268,N_9594,N_9571);
nor U10269 (N_10269,N_9548,N_9988);
or U10270 (N_10270,N_9983,N_9592);
xnor U10271 (N_10271,N_9840,N_9695);
nand U10272 (N_10272,N_9741,N_9543);
nor U10273 (N_10273,N_9967,N_9943);
and U10274 (N_10274,N_9588,N_9584);
nor U10275 (N_10275,N_9558,N_9648);
xor U10276 (N_10276,N_9935,N_9972);
nor U10277 (N_10277,N_9946,N_9835);
nand U10278 (N_10278,N_9756,N_9822);
and U10279 (N_10279,N_9939,N_9756);
or U10280 (N_10280,N_9834,N_9756);
nand U10281 (N_10281,N_9759,N_9817);
or U10282 (N_10282,N_9551,N_9536);
nand U10283 (N_10283,N_9928,N_9922);
nand U10284 (N_10284,N_9967,N_9898);
nor U10285 (N_10285,N_9573,N_9618);
nor U10286 (N_10286,N_9789,N_9523);
and U10287 (N_10287,N_9530,N_9675);
and U10288 (N_10288,N_9973,N_9865);
or U10289 (N_10289,N_9627,N_9643);
nand U10290 (N_10290,N_9827,N_9907);
nor U10291 (N_10291,N_9828,N_9539);
and U10292 (N_10292,N_9955,N_9931);
and U10293 (N_10293,N_9539,N_9564);
or U10294 (N_10294,N_9811,N_9520);
or U10295 (N_10295,N_9858,N_9694);
and U10296 (N_10296,N_9714,N_9767);
and U10297 (N_10297,N_9686,N_9535);
and U10298 (N_10298,N_9692,N_9775);
nand U10299 (N_10299,N_9755,N_9507);
nand U10300 (N_10300,N_9789,N_9942);
nand U10301 (N_10301,N_9666,N_9927);
nor U10302 (N_10302,N_9543,N_9695);
and U10303 (N_10303,N_9683,N_9553);
nor U10304 (N_10304,N_9707,N_9822);
nand U10305 (N_10305,N_9654,N_9582);
nor U10306 (N_10306,N_9529,N_9598);
and U10307 (N_10307,N_9893,N_9854);
or U10308 (N_10308,N_9775,N_9717);
nor U10309 (N_10309,N_9950,N_9579);
nor U10310 (N_10310,N_9637,N_9847);
nand U10311 (N_10311,N_9802,N_9869);
nor U10312 (N_10312,N_9691,N_9545);
nand U10313 (N_10313,N_9668,N_9616);
or U10314 (N_10314,N_9807,N_9742);
nor U10315 (N_10315,N_9940,N_9711);
nand U10316 (N_10316,N_9507,N_9523);
and U10317 (N_10317,N_9787,N_9844);
and U10318 (N_10318,N_9782,N_9824);
nand U10319 (N_10319,N_9809,N_9606);
nand U10320 (N_10320,N_9546,N_9525);
or U10321 (N_10321,N_9731,N_9944);
and U10322 (N_10322,N_9790,N_9516);
nand U10323 (N_10323,N_9590,N_9677);
nor U10324 (N_10324,N_9899,N_9693);
nand U10325 (N_10325,N_9611,N_9738);
or U10326 (N_10326,N_9928,N_9942);
or U10327 (N_10327,N_9597,N_9937);
or U10328 (N_10328,N_9614,N_9556);
nor U10329 (N_10329,N_9745,N_9622);
nand U10330 (N_10330,N_9722,N_9980);
nor U10331 (N_10331,N_9915,N_9913);
and U10332 (N_10332,N_9663,N_9962);
and U10333 (N_10333,N_9656,N_9778);
nand U10334 (N_10334,N_9602,N_9839);
or U10335 (N_10335,N_9862,N_9858);
or U10336 (N_10336,N_9779,N_9772);
nand U10337 (N_10337,N_9551,N_9876);
nand U10338 (N_10338,N_9763,N_9985);
and U10339 (N_10339,N_9790,N_9523);
nor U10340 (N_10340,N_9633,N_9783);
nor U10341 (N_10341,N_9840,N_9619);
and U10342 (N_10342,N_9762,N_9811);
nand U10343 (N_10343,N_9761,N_9515);
nor U10344 (N_10344,N_9690,N_9709);
nand U10345 (N_10345,N_9691,N_9939);
or U10346 (N_10346,N_9695,N_9512);
or U10347 (N_10347,N_9865,N_9970);
nor U10348 (N_10348,N_9843,N_9988);
or U10349 (N_10349,N_9615,N_9629);
or U10350 (N_10350,N_9943,N_9783);
nand U10351 (N_10351,N_9950,N_9668);
and U10352 (N_10352,N_9902,N_9544);
and U10353 (N_10353,N_9865,N_9669);
and U10354 (N_10354,N_9751,N_9818);
nor U10355 (N_10355,N_9646,N_9869);
and U10356 (N_10356,N_9831,N_9508);
or U10357 (N_10357,N_9965,N_9738);
xnor U10358 (N_10358,N_9570,N_9555);
or U10359 (N_10359,N_9538,N_9806);
nand U10360 (N_10360,N_9963,N_9855);
nor U10361 (N_10361,N_9794,N_9916);
or U10362 (N_10362,N_9538,N_9803);
nand U10363 (N_10363,N_9959,N_9882);
and U10364 (N_10364,N_9542,N_9921);
nor U10365 (N_10365,N_9830,N_9957);
or U10366 (N_10366,N_9518,N_9746);
or U10367 (N_10367,N_9727,N_9958);
or U10368 (N_10368,N_9650,N_9640);
or U10369 (N_10369,N_9878,N_9772);
and U10370 (N_10370,N_9566,N_9965);
nor U10371 (N_10371,N_9869,N_9786);
nor U10372 (N_10372,N_9794,N_9586);
nand U10373 (N_10373,N_9861,N_9641);
or U10374 (N_10374,N_9872,N_9506);
nand U10375 (N_10375,N_9663,N_9896);
and U10376 (N_10376,N_9592,N_9644);
nor U10377 (N_10377,N_9607,N_9744);
xor U10378 (N_10378,N_9882,N_9593);
and U10379 (N_10379,N_9899,N_9760);
and U10380 (N_10380,N_9817,N_9515);
nand U10381 (N_10381,N_9524,N_9717);
or U10382 (N_10382,N_9607,N_9881);
nand U10383 (N_10383,N_9793,N_9943);
nand U10384 (N_10384,N_9782,N_9761);
or U10385 (N_10385,N_9950,N_9844);
nand U10386 (N_10386,N_9792,N_9938);
nor U10387 (N_10387,N_9875,N_9738);
nor U10388 (N_10388,N_9664,N_9917);
nor U10389 (N_10389,N_9867,N_9716);
and U10390 (N_10390,N_9846,N_9948);
nor U10391 (N_10391,N_9992,N_9871);
nor U10392 (N_10392,N_9857,N_9676);
and U10393 (N_10393,N_9528,N_9956);
or U10394 (N_10394,N_9866,N_9690);
nor U10395 (N_10395,N_9617,N_9972);
or U10396 (N_10396,N_9954,N_9594);
nor U10397 (N_10397,N_9567,N_9572);
nor U10398 (N_10398,N_9863,N_9628);
or U10399 (N_10399,N_9517,N_9902);
xnor U10400 (N_10400,N_9804,N_9574);
nor U10401 (N_10401,N_9678,N_9523);
and U10402 (N_10402,N_9536,N_9955);
nand U10403 (N_10403,N_9624,N_9926);
or U10404 (N_10404,N_9540,N_9953);
or U10405 (N_10405,N_9571,N_9878);
and U10406 (N_10406,N_9950,N_9649);
nor U10407 (N_10407,N_9743,N_9758);
and U10408 (N_10408,N_9869,N_9616);
or U10409 (N_10409,N_9625,N_9733);
nor U10410 (N_10410,N_9834,N_9538);
or U10411 (N_10411,N_9815,N_9662);
or U10412 (N_10412,N_9856,N_9634);
or U10413 (N_10413,N_9887,N_9631);
nor U10414 (N_10414,N_9898,N_9680);
nor U10415 (N_10415,N_9842,N_9561);
or U10416 (N_10416,N_9915,N_9844);
nor U10417 (N_10417,N_9689,N_9710);
nand U10418 (N_10418,N_9596,N_9594);
nand U10419 (N_10419,N_9901,N_9989);
nand U10420 (N_10420,N_9618,N_9728);
xnor U10421 (N_10421,N_9610,N_9521);
nand U10422 (N_10422,N_9504,N_9881);
and U10423 (N_10423,N_9817,N_9544);
or U10424 (N_10424,N_9710,N_9913);
nand U10425 (N_10425,N_9588,N_9837);
nor U10426 (N_10426,N_9971,N_9551);
nor U10427 (N_10427,N_9875,N_9669);
nor U10428 (N_10428,N_9917,N_9700);
nand U10429 (N_10429,N_9544,N_9849);
nor U10430 (N_10430,N_9500,N_9713);
or U10431 (N_10431,N_9577,N_9576);
nand U10432 (N_10432,N_9724,N_9936);
or U10433 (N_10433,N_9607,N_9904);
and U10434 (N_10434,N_9930,N_9506);
nand U10435 (N_10435,N_9726,N_9871);
nand U10436 (N_10436,N_9615,N_9826);
nor U10437 (N_10437,N_9731,N_9849);
nor U10438 (N_10438,N_9708,N_9695);
nand U10439 (N_10439,N_9867,N_9887);
and U10440 (N_10440,N_9896,N_9616);
nand U10441 (N_10441,N_9635,N_9801);
xor U10442 (N_10442,N_9766,N_9652);
nor U10443 (N_10443,N_9901,N_9835);
nand U10444 (N_10444,N_9505,N_9847);
or U10445 (N_10445,N_9730,N_9578);
nor U10446 (N_10446,N_9799,N_9616);
or U10447 (N_10447,N_9585,N_9543);
nand U10448 (N_10448,N_9698,N_9620);
and U10449 (N_10449,N_9916,N_9718);
nor U10450 (N_10450,N_9991,N_9608);
and U10451 (N_10451,N_9926,N_9952);
and U10452 (N_10452,N_9852,N_9648);
nor U10453 (N_10453,N_9571,N_9529);
or U10454 (N_10454,N_9548,N_9677);
and U10455 (N_10455,N_9888,N_9625);
and U10456 (N_10456,N_9864,N_9629);
nand U10457 (N_10457,N_9610,N_9898);
nor U10458 (N_10458,N_9775,N_9988);
and U10459 (N_10459,N_9510,N_9506);
or U10460 (N_10460,N_9815,N_9676);
and U10461 (N_10461,N_9796,N_9895);
or U10462 (N_10462,N_9875,N_9946);
or U10463 (N_10463,N_9857,N_9793);
xor U10464 (N_10464,N_9651,N_9539);
and U10465 (N_10465,N_9774,N_9934);
and U10466 (N_10466,N_9632,N_9777);
or U10467 (N_10467,N_9938,N_9548);
nor U10468 (N_10468,N_9602,N_9551);
nand U10469 (N_10469,N_9693,N_9989);
nor U10470 (N_10470,N_9524,N_9798);
and U10471 (N_10471,N_9816,N_9840);
nand U10472 (N_10472,N_9847,N_9868);
nor U10473 (N_10473,N_9781,N_9693);
nor U10474 (N_10474,N_9768,N_9800);
or U10475 (N_10475,N_9971,N_9545);
or U10476 (N_10476,N_9890,N_9631);
nand U10477 (N_10477,N_9955,N_9737);
and U10478 (N_10478,N_9801,N_9979);
nand U10479 (N_10479,N_9744,N_9826);
and U10480 (N_10480,N_9515,N_9548);
nor U10481 (N_10481,N_9551,N_9568);
or U10482 (N_10482,N_9721,N_9652);
or U10483 (N_10483,N_9685,N_9618);
and U10484 (N_10484,N_9999,N_9545);
nand U10485 (N_10485,N_9500,N_9852);
and U10486 (N_10486,N_9920,N_9597);
nand U10487 (N_10487,N_9947,N_9825);
nor U10488 (N_10488,N_9784,N_9917);
or U10489 (N_10489,N_9894,N_9677);
nor U10490 (N_10490,N_9831,N_9639);
and U10491 (N_10491,N_9949,N_9698);
and U10492 (N_10492,N_9572,N_9987);
nand U10493 (N_10493,N_9751,N_9886);
nor U10494 (N_10494,N_9589,N_9634);
nor U10495 (N_10495,N_9518,N_9824);
and U10496 (N_10496,N_9977,N_9759);
nor U10497 (N_10497,N_9993,N_9570);
and U10498 (N_10498,N_9505,N_9573);
or U10499 (N_10499,N_9841,N_9887);
nor U10500 (N_10500,N_10250,N_10113);
and U10501 (N_10501,N_10323,N_10498);
xnor U10502 (N_10502,N_10349,N_10386);
or U10503 (N_10503,N_10181,N_10270);
and U10504 (N_10504,N_10001,N_10253);
nand U10505 (N_10505,N_10082,N_10173);
nand U10506 (N_10506,N_10102,N_10475);
and U10507 (N_10507,N_10421,N_10021);
or U10508 (N_10508,N_10306,N_10132);
nor U10509 (N_10509,N_10031,N_10047);
or U10510 (N_10510,N_10368,N_10107);
or U10511 (N_10511,N_10317,N_10260);
xor U10512 (N_10512,N_10159,N_10118);
or U10513 (N_10513,N_10030,N_10259);
or U10514 (N_10514,N_10456,N_10397);
nor U10515 (N_10515,N_10169,N_10350);
nand U10516 (N_10516,N_10455,N_10236);
xnor U10517 (N_10517,N_10227,N_10239);
or U10518 (N_10518,N_10088,N_10376);
and U10519 (N_10519,N_10049,N_10203);
nor U10520 (N_10520,N_10366,N_10197);
and U10521 (N_10521,N_10426,N_10002);
and U10522 (N_10522,N_10210,N_10122);
nand U10523 (N_10523,N_10328,N_10193);
nor U10524 (N_10524,N_10037,N_10019);
nor U10525 (N_10525,N_10178,N_10420);
nor U10526 (N_10526,N_10053,N_10111);
nand U10527 (N_10527,N_10060,N_10123);
nand U10528 (N_10528,N_10240,N_10115);
nor U10529 (N_10529,N_10235,N_10453);
or U10530 (N_10530,N_10369,N_10084);
or U10531 (N_10531,N_10375,N_10352);
nand U10532 (N_10532,N_10042,N_10414);
nor U10533 (N_10533,N_10175,N_10283);
nand U10534 (N_10534,N_10033,N_10373);
and U10535 (N_10535,N_10055,N_10472);
or U10536 (N_10536,N_10075,N_10480);
nand U10537 (N_10537,N_10061,N_10231);
nor U10538 (N_10538,N_10171,N_10223);
and U10539 (N_10539,N_10464,N_10158);
nor U10540 (N_10540,N_10219,N_10412);
or U10541 (N_10541,N_10092,N_10285);
nand U10542 (N_10542,N_10150,N_10196);
and U10543 (N_10543,N_10449,N_10457);
nor U10544 (N_10544,N_10229,N_10416);
and U10545 (N_10545,N_10380,N_10089);
xor U10546 (N_10546,N_10172,N_10331);
nand U10547 (N_10547,N_10012,N_10090);
nand U10548 (N_10548,N_10126,N_10351);
nor U10549 (N_10549,N_10269,N_10013);
nor U10550 (N_10550,N_10070,N_10446);
nor U10551 (N_10551,N_10432,N_10281);
or U10552 (N_10552,N_10043,N_10182);
xor U10553 (N_10553,N_10304,N_10409);
or U10554 (N_10554,N_10322,N_10309);
or U10555 (N_10555,N_10356,N_10408);
and U10556 (N_10556,N_10257,N_10488);
or U10557 (N_10557,N_10363,N_10041);
nor U10558 (N_10558,N_10057,N_10212);
nor U10559 (N_10559,N_10010,N_10301);
or U10560 (N_10560,N_10339,N_10124);
and U10561 (N_10561,N_10401,N_10162);
nand U10562 (N_10562,N_10395,N_10467);
nor U10563 (N_10563,N_10147,N_10136);
nand U10564 (N_10564,N_10161,N_10149);
nand U10565 (N_10565,N_10438,N_10016);
or U10566 (N_10566,N_10462,N_10135);
nand U10567 (N_10567,N_10489,N_10388);
nor U10568 (N_10568,N_10121,N_10288);
nor U10569 (N_10569,N_10476,N_10479);
and U10570 (N_10570,N_10248,N_10407);
or U10571 (N_10571,N_10244,N_10371);
nor U10572 (N_10572,N_10068,N_10080);
nor U10573 (N_10573,N_10417,N_10059);
and U10574 (N_10574,N_10286,N_10374);
nand U10575 (N_10575,N_10278,N_10028);
nor U10576 (N_10576,N_10390,N_10074);
or U10577 (N_10577,N_10251,N_10141);
or U10578 (N_10578,N_10246,N_10180);
nor U10579 (N_10579,N_10461,N_10392);
nand U10580 (N_10580,N_10105,N_10473);
nand U10581 (N_10581,N_10382,N_10142);
or U10582 (N_10582,N_10297,N_10367);
or U10583 (N_10583,N_10311,N_10497);
xnor U10584 (N_10584,N_10496,N_10011);
nor U10585 (N_10585,N_10035,N_10213);
or U10586 (N_10586,N_10291,N_10134);
and U10587 (N_10587,N_10381,N_10211);
nor U10588 (N_10588,N_10316,N_10282);
nor U10589 (N_10589,N_10048,N_10441);
or U10590 (N_10590,N_10184,N_10129);
or U10591 (N_10591,N_10450,N_10263);
and U10592 (N_10592,N_10003,N_10085);
or U10593 (N_10593,N_10146,N_10287);
nand U10594 (N_10594,N_10387,N_10333);
or U10595 (N_10595,N_10303,N_10199);
and U10596 (N_10596,N_10233,N_10261);
nor U10597 (N_10597,N_10471,N_10298);
or U10598 (N_10598,N_10360,N_10133);
and U10599 (N_10599,N_10299,N_10204);
nand U10600 (N_10600,N_10018,N_10344);
xnor U10601 (N_10601,N_10396,N_10022);
nor U10602 (N_10602,N_10237,N_10329);
or U10603 (N_10603,N_10069,N_10034);
and U10604 (N_10604,N_10170,N_10198);
or U10605 (N_10605,N_10241,N_10209);
nor U10606 (N_10606,N_10341,N_10137);
nand U10607 (N_10607,N_10347,N_10429);
nor U10608 (N_10608,N_10091,N_10385);
xor U10609 (N_10609,N_10076,N_10358);
nor U10610 (N_10610,N_10109,N_10004);
nor U10611 (N_10611,N_10495,N_10086);
nand U10612 (N_10612,N_10087,N_10112);
and U10613 (N_10613,N_10362,N_10389);
or U10614 (N_10614,N_10359,N_10006);
nor U10615 (N_10615,N_10063,N_10202);
nand U10616 (N_10616,N_10007,N_10312);
and U10617 (N_10617,N_10348,N_10065);
or U10618 (N_10618,N_10214,N_10313);
and U10619 (N_10619,N_10459,N_10024);
nand U10620 (N_10620,N_10415,N_10258);
xnor U10621 (N_10621,N_10234,N_10200);
nor U10622 (N_10622,N_10195,N_10393);
nor U10623 (N_10623,N_10208,N_10096);
and U10624 (N_10624,N_10160,N_10145);
and U10625 (N_10625,N_10230,N_10155);
nor U10626 (N_10626,N_10454,N_10337);
and U10627 (N_10627,N_10399,N_10081);
nand U10628 (N_10628,N_10310,N_10130);
nand U10629 (N_10629,N_10361,N_10465);
and U10630 (N_10630,N_10190,N_10383);
or U10631 (N_10631,N_10384,N_10357);
and U10632 (N_10632,N_10242,N_10424);
and U10633 (N_10633,N_10120,N_10015);
nor U10634 (N_10634,N_10413,N_10174);
and U10635 (N_10635,N_10143,N_10046);
or U10636 (N_10636,N_10486,N_10494);
and U10637 (N_10637,N_10425,N_10493);
and U10638 (N_10638,N_10218,N_10404);
and U10639 (N_10639,N_10305,N_10423);
nand U10640 (N_10640,N_10083,N_10192);
nor U10641 (N_10641,N_10452,N_10247);
or U10642 (N_10642,N_10179,N_10378);
xor U10643 (N_10643,N_10443,N_10419);
or U10644 (N_10644,N_10290,N_10463);
or U10645 (N_10645,N_10164,N_10428);
or U10646 (N_10646,N_10029,N_10444);
nand U10647 (N_10647,N_10405,N_10418);
or U10648 (N_10648,N_10117,N_10077);
or U10649 (N_10649,N_10294,N_10321);
nor U10650 (N_10650,N_10326,N_10436);
or U10651 (N_10651,N_10252,N_10153);
and U10652 (N_10652,N_10140,N_10460);
and U10653 (N_10653,N_10435,N_10110);
nand U10654 (N_10654,N_10266,N_10220);
nand U10655 (N_10655,N_10157,N_10325);
or U10656 (N_10656,N_10481,N_10265);
nor U10657 (N_10657,N_10009,N_10051);
xnor U10658 (N_10658,N_10127,N_10335);
nor U10659 (N_10659,N_10165,N_10400);
or U10660 (N_10660,N_10119,N_10274);
nor U10661 (N_10661,N_10295,N_10207);
or U10662 (N_10662,N_10152,N_10045);
and U10663 (N_10663,N_10292,N_10072);
and U10664 (N_10664,N_10078,N_10353);
and U10665 (N_10665,N_10094,N_10040);
and U10666 (N_10666,N_10098,N_10492);
and U10667 (N_10667,N_10267,N_10448);
and U10668 (N_10668,N_10330,N_10319);
nor U10669 (N_10669,N_10422,N_10314);
and U10670 (N_10670,N_10289,N_10279);
or U10671 (N_10671,N_10485,N_10437);
or U10672 (N_10672,N_10372,N_10017);
nor U10673 (N_10673,N_10228,N_10044);
and U10674 (N_10674,N_10243,N_10280);
or U10675 (N_10675,N_10490,N_10308);
nor U10676 (N_10676,N_10249,N_10014);
or U10677 (N_10677,N_10073,N_10458);
and U10678 (N_10678,N_10032,N_10410);
nand U10679 (N_10679,N_10254,N_10217);
and U10680 (N_10680,N_10340,N_10271);
nand U10681 (N_10681,N_10020,N_10238);
nor U10682 (N_10682,N_10370,N_10054);
nand U10683 (N_10683,N_10148,N_10005);
nand U10684 (N_10684,N_10483,N_10255);
and U10685 (N_10685,N_10008,N_10262);
nand U10686 (N_10686,N_10038,N_10245);
nand U10687 (N_10687,N_10000,N_10491);
and U10688 (N_10688,N_10232,N_10320);
or U10689 (N_10689,N_10183,N_10264);
and U10690 (N_10690,N_10050,N_10433);
or U10691 (N_10691,N_10469,N_10151);
and U10692 (N_10692,N_10205,N_10499);
nand U10693 (N_10693,N_10191,N_10027);
nor U10694 (N_10694,N_10166,N_10125);
nand U10695 (N_10695,N_10036,N_10188);
nor U10696 (N_10696,N_10206,N_10201);
or U10697 (N_10697,N_10163,N_10277);
and U10698 (N_10698,N_10300,N_10144);
nor U10699 (N_10699,N_10345,N_10466);
or U10700 (N_10700,N_10156,N_10355);
and U10701 (N_10701,N_10186,N_10104);
nor U10702 (N_10702,N_10365,N_10324);
and U10703 (N_10703,N_10484,N_10114);
and U10704 (N_10704,N_10430,N_10411);
and U10705 (N_10705,N_10403,N_10058);
nor U10706 (N_10706,N_10442,N_10071);
and U10707 (N_10707,N_10406,N_10256);
nand U10708 (N_10708,N_10176,N_10434);
nand U10709 (N_10709,N_10336,N_10154);
nand U10710 (N_10710,N_10346,N_10477);
nor U10711 (N_10711,N_10099,N_10215);
xnor U10712 (N_10712,N_10440,N_10116);
and U10713 (N_10713,N_10026,N_10445);
nand U10714 (N_10714,N_10189,N_10097);
and U10715 (N_10715,N_10474,N_10284);
and U10716 (N_10716,N_10108,N_10342);
or U10717 (N_10717,N_10025,N_10296);
or U10718 (N_10718,N_10398,N_10222);
nor U10719 (N_10719,N_10302,N_10293);
nand U10720 (N_10720,N_10128,N_10221);
and U10721 (N_10721,N_10167,N_10106);
or U10722 (N_10722,N_10187,N_10185);
and U10723 (N_10723,N_10138,N_10427);
or U10724 (N_10724,N_10327,N_10268);
or U10725 (N_10725,N_10354,N_10470);
nand U10726 (N_10726,N_10343,N_10067);
and U10727 (N_10727,N_10225,N_10039);
and U10728 (N_10728,N_10095,N_10194);
or U10729 (N_10729,N_10377,N_10272);
and U10730 (N_10730,N_10103,N_10131);
nor U10731 (N_10731,N_10139,N_10402);
or U10732 (N_10732,N_10468,N_10066);
and U10733 (N_10733,N_10275,N_10334);
or U10734 (N_10734,N_10226,N_10273);
xnor U10735 (N_10735,N_10079,N_10447);
xor U10736 (N_10736,N_10332,N_10224);
nand U10737 (N_10737,N_10431,N_10487);
nand U10738 (N_10738,N_10216,N_10338);
or U10739 (N_10739,N_10100,N_10478);
nor U10740 (N_10740,N_10062,N_10093);
or U10741 (N_10741,N_10379,N_10168);
and U10742 (N_10742,N_10177,N_10023);
nand U10743 (N_10743,N_10315,N_10101);
nand U10744 (N_10744,N_10394,N_10052);
or U10745 (N_10745,N_10482,N_10056);
nor U10746 (N_10746,N_10318,N_10307);
nand U10747 (N_10747,N_10364,N_10391);
and U10748 (N_10748,N_10064,N_10451);
nand U10749 (N_10749,N_10276,N_10439);
or U10750 (N_10750,N_10396,N_10051);
nand U10751 (N_10751,N_10300,N_10054);
xnor U10752 (N_10752,N_10250,N_10045);
and U10753 (N_10753,N_10492,N_10398);
nand U10754 (N_10754,N_10260,N_10062);
and U10755 (N_10755,N_10120,N_10212);
or U10756 (N_10756,N_10286,N_10382);
nor U10757 (N_10757,N_10063,N_10346);
or U10758 (N_10758,N_10094,N_10090);
or U10759 (N_10759,N_10339,N_10197);
nand U10760 (N_10760,N_10212,N_10308);
and U10761 (N_10761,N_10043,N_10039);
or U10762 (N_10762,N_10048,N_10288);
or U10763 (N_10763,N_10015,N_10072);
nor U10764 (N_10764,N_10060,N_10052);
nor U10765 (N_10765,N_10056,N_10185);
nor U10766 (N_10766,N_10478,N_10381);
nor U10767 (N_10767,N_10479,N_10369);
xor U10768 (N_10768,N_10434,N_10047);
and U10769 (N_10769,N_10008,N_10272);
and U10770 (N_10770,N_10440,N_10443);
and U10771 (N_10771,N_10170,N_10187);
nor U10772 (N_10772,N_10311,N_10023);
or U10773 (N_10773,N_10119,N_10458);
nor U10774 (N_10774,N_10483,N_10061);
and U10775 (N_10775,N_10432,N_10167);
nor U10776 (N_10776,N_10115,N_10283);
or U10777 (N_10777,N_10209,N_10004);
nand U10778 (N_10778,N_10028,N_10309);
nand U10779 (N_10779,N_10011,N_10424);
or U10780 (N_10780,N_10355,N_10001);
nor U10781 (N_10781,N_10426,N_10402);
nor U10782 (N_10782,N_10437,N_10039);
nor U10783 (N_10783,N_10412,N_10116);
nand U10784 (N_10784,N_10103,N_10355);
nand U10785 (N_10785,N_10019,N_10175);
nand U10786 (N_10786,N_10196,N_10099);
nor U10787 (N_10787,N_10422,N_10460);
or U10788 (N_10788,N_10324,N_10371);
xnor U10789 (N_10789,N_10346,N_10466);
and U10790 (N_10790,N_10195,N_10063);
nor U10791 (N_10791,N_10088,N_10136);
and U10792 (N_10792,N_10360,N_10484);
nor U10793 (N_10793,N_10342,N_10223);
nor U10794 (N_10794,N_10011,N_10262);
or U10795 (N_10795,N_10327,N_10008);
or U10796 (N_10796,N_10194,N_10209);
and U10797 (N_10797,N_10057,N_10409);
or U10798 (N_10798,N_10304,N_10324);
or U10799 (N_10799,N_10061,N_10069);
nor U10800 (N_10800,N_10455,N_10469);
and U10801 (N_10801,N_10128,N_10089);
nor U10802 (N_10802,N_10436,N_10189);
nor U10803 (N_10803,N_10267,N_10391);
nand U10804 (N_10804,N_10054,N_10434);
or U10805 (N_10805,N_10426,N_10291);
and U10806 (N_10806,N_10227,N_10361);
nand U10807 (N_10807,N_10059,N_10309);
xor U10808 (N_10808,N_10305,N_10309);
nor U10809 (N_10809,N_10366,N_10114);
nand U10810 (N_10810,N_10375,N_10343);
nor U10811 (N_10811,N_10262,N_10268);
and U10812 (N_10812,N_10143,N_10206);
xor U10813 (N_10813,N_10328,N_10368);
and U10814 (N_10814,N_10423,N_10252);
nor U10815 (N_10815,N_10182,N_10380);
nor U10816 (N_10816,N_10131,N_10319);
and U10817 (N_10817,N_10282,N_10019);
nor U10818 (N_10818,N_10207,N_10072);
and U10819 (N_10819,N_10374,N_10234);
and U10820 (N_10820,N_10041,N_10111);
nand U10821 (N_10821,N_10037,N_10206);
nor U10822 (N_10822,N_10031,N_10349);
and U10823 (N_10823,N_10146,N_10159);
and U10824 (N_10824,N_10314,N_10016);
nand U10825 (N_10825,N_10080,N_10023);
nor U10826 (N_10826,N_10285,N_10106);
and U10827 (N_10827,N_10405,N_10157);
nand U10828 (N_10828,N_10118,N_10339);
xnor U10829 (N_10829,N_10308,N_10085);
nand U10830 (N_10830,N_10061,N_10004);
nand U10831 (N_10831,N_10075,N_10210);
nand U10832 (N_10832,N_10160,N_10006);
or U10833 (N_10833,N_10080,N_10345);
nand U10834 (N_10834,N_10278,N_10208);
nor U10835 (N_10835,N_10252,N_10295);
and U10836 (N_10836,N_10407,N_10234);
or U10837 (N_10837,N_10430,N_10406);
nor U10838 (N_10838,N_10074,N_10019);
nor U10839 (N_10839,N_10433,N_10065);
nand U10840 (N_10840,N_10128,N_10312);
nand U10841 (N_10841,N_10099,N_10481);
or U10842 (N_10842,N_10121,N_10369);
nor U10843 (N_10843,N_10226,N_10394);
or U10844 (N_10844,N_10094,N_10296);
nor U10845 (N_10845,N_10269,N_10137);
or U10846 (N_10846,N_10338,N_10445);
or U10847 (N_10847,N_10293,N_10059);
or U10848 (N_10848,N_10474,N_10445);
or U10849 (N_10849,N_10303,N_10020);
and U10850 (N_10850,N_10350,N_10151);
nand U10851 (N_10851,N_10341,N_10322);
nand U10852 (N_10852,N_10236,N_10255);
or U10853 (N_10853,N_10215,N_10425);
and U10854 (N_10854,N_10425,N_10481);
nand U10855 (N_10855,N_10343,N_10089);
nor U10856 (N_10856,N_10132,N_10104);
xor U10857 (N_10857,N_10085,N_10474);
or U10858 (N_10858,N_10251,N_10488);
nand U10859 (N_10859,N_10064,N_10118);
and U10860 (N_10860,N_10139,N_10114);
or U10861 (N_10861,N_10240,N_10316);
and U10862 (N_10862,N_10091,N_10074);
nor U10863 (N_10863,N_10302,N_10474);
and U10864 (N_10864,N_10463,N_10473);
nand U10865 (N_10865,N_10107,N_10442);
nor U10866 (N_10866,N_10442,N_10000);
nand U10867 (N_10867,N_10083,N_10011);
or U10868 (N_10868,N_10429,N_10448);
or U10869 (N_10869,N_10089,N_10236);
or U10870 (N_10870,N_10201,N_10004);
nand U10871 (N_10871,N_10476,N_10410);
nor U10872 (N_10872,N_10415,N_10366);
nor U10873 (N_10873,N_10101,N_10442);
nor U10874 (N_10874,N_10255,N_10045);
and U10875 (N_10875,N_10112,N_10327);
nor U10876 (N_10876,N_10337,N_10231);
and U10877 (N_10877,N_10004,N_10334);
and U10878 (N_10878,N_10148,N_10292);
nor U10879 (N_10879,N_10180,N_10253);
or U10880 (N_10880,N_10476,N_10150);
xor U10881 (N_10881,N_10072,N_10181);
or U10882 (N_10882,N_10247,N_10204);
nand U10883 (N_10883,N_10368,N_10267);
nand U10884 (N_10884,N_10404,N_10360);
nand U10885 (N_10885,N_10337,N_10388);
or U10886 (N_10886,N_10017,N_10307);
nand U10887 (N_10887,N_10462,N_10421);
or U10888 (N_10888,N_10211,N_10241);
or U10889 (N_10889,N_10312,N_10155);
or U10890 (N_10890,N_10024,N_10424);
nor U10891 (N_10891,N_10490,N_10407);
and U10892 (N_10892,N_10020,N_10315);
or U10893 (N_10893,N_10265,N_10331);
nor U10894 (N_10894,N_10007,N_10001);
nor U10895 (N_10895,N_10078,N_10251);
and U10896 (N_10896,N_10198,N_10027);
nor U10897 (N_10897,N_10459,N_10346);
nand U10898 (N_10898,N_10302,N_10001);
nor U10899 (N_10899,N_10016,N_10367);
or U10900 (N_10900,N_10241,N_10445);
nor U10901 (N_10901,N_10362,N_10413);
and U10902 (N_10902,N_10356,N_10047);
nor U10903 (N_10903,N_10390,N_10397);
nor U10904 (N_10904,N_10316,N_10024);
nand U10905 (N_10905,N_10345,N_10203);
xor U10906 (N_10906,N_10052,N_10458);
and U10907 (N_10907,N_10098,N_10154);
nor U10908 (N_10908,N_10271,N_10026);
nand U10909 (N_10909,N_10077,N_10044);
nand U10910 (N_10910,N_10120,N_10251);
or U10911 (N_10911,N_10320,N_10304);
nor U10912 (N_10912,N_10113,N_10005);
nor U10913 (N_10913,N_10064,N_10423);
nor U10914 (N_10914,N_10492,N_10461);
nand U10915 (N_10915,N_10006,N_10117);
nor U10916 (N_10916,N_10479,N_10277);
nor U10917 (N_10917,N_10281,N_10360);
or U10918 (N_10918,N_10033,N_10219);
nand U10919 (N_10919,N_10231,N_10382);
and U10920 (N_10920,N_10101,N_10019);
nor U10921 (N_10921,N_10285,N_10429);
nand U10922 (N_10922,N_10421,N_10280);
nor U10923 (N_10923,N_10430,N_10296);
nand U10924 (N_10924,N_10135,N_10028);
and U10925 (N_10925,N_10088,N_10153);
and U10926 (N_10926,N_10137,N_10319);
nor U10927 (N_10927,N_10496,N_10089);
nor U10928 (N_10928,N_10129,N_10323);
nor U10929 (N_10929,N_10237,N_10038);
nor U10930 (N_10930,N_10119,N_10324);
and U10931 (N_10931,N_10489,N_10161);
or U10932 (N_10932,N_10093,N_10243);
nand U10933 (N_10933,N_10187,N_10427);
and U10934 (N_10934,N_10324,N_10461);
nor U10935 (N_10935,N_10091,N_10097);
nand U10936 (N_10936,N_10293,N_10252);
nand U10937 (N_10937,N_10329,N_10307);
and U10938 (N_10938,N_10147,N_10351);
nand U10939 (N_10939,N_10469,N_10186);
nand U10940 (N_10940,N_10470,N_10035);
and U10941 (N_10941,N_10317,N_10320);
or U10942 (N_10942,N_10208,N_10197);
nor U10943 (N_10943,N_10033,N_10027);
nor U10944 (N_10944,N_10487,N_10213);
and U10945 (N_10945,N_10309,N_10063);
and U10946 (N_10946,N_10090,N_10064);
nand U10947 (N_10947,N_10106,N_10401);
or U10948 (N_10948,N_10315,N_10054);
nor U10949 (N_10949,N_10237,N_10158);
nor U10950 (N_10950,N_10049,N_10196);
nand U10951 (N_10951,N_10466,N_10090);
nand U10952 (N_10952,N_10170,N_10255);
or U10953 (N_10953,N_10082,N_10060);
or U10954 (N_10954,N_10124,N_10359);
nand U10955 (N_10955,N_10144,N_10418);
nor U10956 (N_10956,N_10102,N_10438);
and U10957 (N_10957,N_10068,N_10429);
nand U10958 (N_10958,N_10333,N_10090);
nor U10959 (N_10959,N_10269,N_10057);
nand U10960 (N_10960,N_10223,N_10287);
and U10961 (N_10961,N_10237,N_10318);
and U10962 (N_10962,N_10002,N_10385);
or U10963 (N_10963,N_10497,N_10084);
xor U10964 (N_10964,N_10090,N_10365);
nor U10965 (N_10965,N_10151,N_10012);
nand U10966 (N_10966,N_10159,N_10014);
or U10967 (N_10967,N_10285,N_10355);
or U10968 (N_10968,N_10477,N_10440);
nor U10969 (N_10969,N_10048,N_10123);
or U10970 (N_10970,N_10312,N_10149);
nand U10971 (N_10971,N_10052,N_10325);
or U10972 (N_10972,N_10147,N_10409);
and U10973 (N_10973,N_10461,N_10346);
or U10974 (N_10974,N_10471,N_10096);
nand U10975 (N_10975,N_10284,N_10405);
and U10976 (N_10976,N_10446,N_10107);
nor U10977 (N_10977,N_10316,N_10280);
or U10978 (N_10978,N_10022,N_10473);
or U10979 (N_10979,N_10131,N_10022);
and U10980 (N_10980,N_10326,N_10002);
and U10981 (N_10981,N_10097,N_10295);
or U10982 (N_10982,N_10355,N_10483);
or U10983 (N_10983,N_10080,N_10467);
xor U10984 (N_10984,N_10058,N_10217);
nand U10985 (N_10985,N_10267,N_10293);
or U10986 (N_10986,N_10398,N_10115);
nand U10987 (N_10987,N_10308,N_10422);
or U10988 (N_10988,N_10288,N_10123);
and U10989 (N_10989,N_10047,N_10438);
nand U10990 (N_10990,N_10495,N_10397);
nand U10991 (N_10991,N_10371,N_10436);
or U10992 (N_10992,N_10290,N_10360);
and U10993 (N_10993,N_10094,N_10113);
or U10994 (N_10994,N_10012,N_10219);
xor U10995 (N_10995,N_10228,N_10059);
and U10996 (N_10996,N_10110,N_10234);
and U10997 (N_10997,N_10179,N_10046);
nand U10998 (N_10998,N_10114,N_10175);
and U10999 (N_10999,N_10014,N_10023);
and U11000 (N_11000,N_10523,N_10916);
xor U11001 (N_11001,N_10884,N_10737);
and U11002 (N_11002,N_10664,N_10872);
or U11003 (N_11003,N_10663,N_10711);
and U11004 (N_11004,N_10649,N_10639);
nand U11005 (N_11005,N_10821,N_10651);
or U11006 (N_11006,N_10689,N_10814);
nor U11007 (N_11007,N_10927,N_10815);
or U11008 (N_11008,N_10577,N_10706);
nor U11009 (N_11009,N_10501,N_10589);
nor U11010 (N_11010,N_10882,N_10991);
or U11011 (N_11011,N_10963,N_10655);
nand U11012 (N_11012,N_10946,N_10970);
nor U11013 (N_11013,N_10835,N_10820);
nand U11014 (N_11014,N_10583,N_10903);
nor U11015 (N_11015,N_10531,N_10964);
nor U11016 (N_11016,N_10770,N_10848);
or U11017 (N_11017,N_10829,N_10900);
or U11018 (N_11018,N_10701,N_10819);
and U11019 (N_11019,N_10792,N_10873);
nand U11020 (N_11020,N_10541,N_10671);
nor U11021 (N_11021,N_10551,N_10666);
or U11022 (N_11022,N_10597,N_10846);
nor U11023 (N_11023,N_10885,N_10746);
nor U11024 (N_11024,N_10606,N_10847);
nand U11025 (N_11025,N_10795,N_10668);
and U11026 (N_11026,N_10537,N_10911);
nor U11027 (N_11027,N_10810,N_10894);
nor U11028 (N_11028,N_10607,N_10506);
and U11029 (N_11029,N_10683,N_10625);
or U11030 (N_11030,N_10773,N_10776);
or U11031 (N_11031,N_10553,N_10744);
or U11032 (N_11032,N_10966,N_10850);
and U11033 (N_11033,N_10640,N_10648);
and U11034 (N_11034,N_10700,N_10581);
or U11035 (N_11035,N_10834,N_10529);
or U11036 (N_11036,N_10520,N_10984);
nor U11037 (N_11037,N_10684,N_10713);
xnor U11038 (N_11038,N_10590,N_10538);
and U11039 (N_11039,N_10856,N_10533);
nor U11040 (N_11040,N_10790,N_10886);
nor U11041 (N_11041,N_10967,N_10564);
and U11042 (N_11042,N_10867,N_10877);
or U11043 (N_11043,N_10956,N_10679);
and U11044 (N_11044,N_10839,N_10576);
xor U11045 (N_11045,N_10628,N_10986);
or U11046 (N_11046,N_10889,N_10527);
or U11047 (N_11047,N_10643,N_10945);
nand U11048 (N_11048,N_10854,N_10552);
and U11049 (N_11049,N_10980,N_10785);
or U11050 (N_11050,N_10682,N_10557);
and U11051 (N_11051,N_10898,N_10563);
nand U11052 (N_11052,N_10755,N_10862);
and U11053 (N_11053,N_10811,N_10917);
nor U11054 (N_11054,N_10543,N_10601);
or U11055 (N_11055,N_10592,N_10787);
nor U11056 (N_11056,N_10715,N_10705);
nor U11057 (N_11057,N_10824,N_10925);
nor U11058 (N_11058,N_10570,N_10922);
nand U11059 (N_11059,N_10812,N_10940);
and U11060 (N_11060,N_10871,N_10818);
nand U11061 (N_11061,N_10636,N_10968);
or U11062 (N_11062,N_10864,N_10539);
and U11063 (N_11063,N_10909,N_10626);
nor U11064 (N_11064,N_10727,N_10765);
nor U11065 (N_11065,N_10514,N_10961);
or U11066 (N_11066,N_10841,N_10883);
nand U11067 (N_11067,N_10604,N_10960);
nor U11068 (N_11068,N_10645,N_10914);
or U11069 (N_11069,N_10575,N_10594);
and U11070 (N_11070,N_10730,N_10751);
nor U11071 (N_11071,N_10504,N_10611);
nor U11072 (N_11072,N_10673,N_10972);
xor U11073 (N_11073,N_10653,N_10709);
and U11074 (N_11074,N_10941,N_10723);
nand U11075 (N_11075,N_10919,N_10708);
or U11076 (N_11076,N_10974,N_10778);
nand U11077 (N_11077,N_10769,N_10665);
or U11078 (N_11078,N_10609,N_10851);
nand U11079 (N_11079,N_10912,N_10513);
and U11080 (N_11080,N_10863,N_10540);
nor U11081 (N_11081,N_10585,N_10977);
nor U11082 (N_11082,N_10996,N_10608);
nand U11083 (N_11083,N_10624,N_10870);
or U11084 (N_11084,N_10627,N_10943);
nor U11085 (N_11085,N_10750,N_10722);
nor U11086 (N_11086,N_10754,N_10830);
nor U11087 (N_11087,N_10717,N_10779);
nor U11088 (N_11088,N_10837,N_10800);
nor U11089 (N_11089,N_10955,N_10733);
or U11090 (N_11090,N_10740,N_10735);
and U11091 (N_11091,N_10780,N_10893);
nand U11092 (N_11092,N_10749,N_10803);
or U11093 (N_11093,N_10549,N_10562);
nand U11094 (N_11094,N_10822,N_10808);
nor U11095 (N_11095,N_10516,N_10798);
and U11096 (N_11096,N_10794,N_10888);
nor U11097 (N_11097,N_10556,N_10638);
and U11098 (N_11098,N_10853,N_10857);
nand U11099 (N_11099,N_10633,N_10817);
nand U11100 (N_11100,N_10695,N_10542);
nand U11101 (N_11101,N_10567,N_10505);
or U11102 (N_11102,N_10997,N_10752);
nor U11103 (N_11103,N_10712,N_10586);
nand U11104 (N_11104,N_10936,N_10660);
nor U11105 (N_11105,N_10572,N_10860);
nor U11106 (N_11106,N_10699,N_10659);
nor U11107 (N_11107,N_10587,N_10518);
or U11108 (N_11108,N_10844,N_10908);
nor U11109 (N_11109,N_10758,N_10521);
or U11110 (N_11110,N_10995,N_10732);
nor U11111 (N_11111,N_10990,N_10958);
nor U11112 (N_11112,N_10681,N_10729);
and U11113 (N_11113,N_10550,N_10804);
nor U11114 (N_11114,N_10767,N_10985);
or U11115 (N_11115,N_10670,N_10704);
or U11116 (N_11116,N_10612,N_10509);
and U11117 (N_11117,N_10630,N_10992);
or U11118 (N_11118,N_10788,N_10632);
or U11119 (N_11119,N_10545,N_10957);
nand U11120 (N_11120,N_10634,N_10703);
nand U11121 (N_11121,N_10881,N_10535);
and U11122 (N_11122,N_10629,N_10823);
nor U11123 (N_11123,N_10502,N_10865);
and U11124 (N_11124,N_10775,N_10813);
or U11125 (N_11125,N_10678,N_10993);
and U11126 (N_11126,N_10906,N_10616);
or U11127 (N_11127,N_10652,N_10667);
or U11128 (N_11128,N_10661,N_10532);
or U11129 (N_11129,N_10641,N_10613);
nor U11130 (N_11130,N_10631,N_10987);
or U11131 (N_11131,N_10547,N_10675);
nand U11132 (N_11132,N_10680,N_10897);
and U11133 (N_11133,N_10763,N_10947);
nor U11134 (N_11134,N_10603,N_10544);
or U11135 (N_11135,N_10726,N_10582);
or U11136 (N_11136,N_10852,N_10528);
nor U11137 (N_11137,N_10784,N_10588);
nor U11138 (N_11138,N_10696,N_10646);
and U11139 (N_11139,N_10685,N_10791);
or U11140 (N_11140,N_10650,N_10716);
and U11141 (N_11141,N_10904,N_10560);
and U11142 (N_11142,N_10962,N_10831);
nand U11143 (N_11143,N_10500,N_10915);
nand U11144 (N_11144,N_10690,N_10969);
and U11145 (N_11145,N_10738,N_10524);
nor U11146 (N_11146,N_10918,N_10789);
nand U11147 (N_11147,N_10954,N_10921);
or U11148 (N_11148,N_10939,N_10694);
or U11149 (N_11149,N_10658,N_10714);
or U11150 (N_11150,N_10797,N_10507);
and U11151 (N_11151,N_10774,N_10756);
and U11152 (N_11152,N_10933,N_10981);
xnor U11153 (N_11153,N_10760,N_10907);
or U11154 (N_11154,N_10623,N_10517);
or U11155 (N_11155,N_10994,N_10747);
and U11156 (N_11156,N_10595,N_10574);
nand U11157 (N_11157,N_10619,N_10771);
nand U11158 (N_11158,N_10686,N_10832);
nand U11159 (N_11159,N_10736,N_10620);
or U11160 (N_11160,N_10905,N_10944);
and U11161 (N_11161,N_10875,N_10555);
nand U11162 (N_11162,N_10827,N_10838);
nand U11163 (N_11163,N_10739,N_10573);
nand U11164 (N_11164,N_10635,N_10859);
or U11165 (N_11165,N_10975,N_10759);
or U11166 (N_11166,N_10833,N_10828);
nor U11167 (N_11167,N_10669,N_10610);
and U11168 (N_11168,N_10536,N_10546);
and U11169 (N_11169,N_10932,N_10742);
nor U11170 (N_11170,N_10887,N_10615);
nand U11171 (N_11171,N_10973,N_10558);
or U11172 (N_11172,N_10692,N_10777);
nor U11173 (N_11173,N_10948,N_10725);
nor U11174 (N_11174,N_10796,N_10766);
nor U11175 (N_11175,N_10805,N_10728);
nand U11176 (N_11176,N_10724,N_10757);
and U11177 (N_11177,N_10861,N_10534);
or U11178 (N_11178,N_10976,N_10935);
or U11179 (N_11179,N_10734,N_10998);
nand U11180 (N_11180,N_10866,N_10772);
nor U11181 (N_11181,N_10710,N_10930);
nor U11182 (N_11182,N_10929,N_10858);
nor U11183 (N_11183,N_10720,N_10598);
nand U11184 (N_11184,N_10674,N_10868);
and U11185 (N_11185,N_10702,N_10559);
nor U11186 (N_11186,N_10693,N_10845);
or U11187 (N_11187,N_10983,N_10842);
nor U11188 (N_11188,N_10978,N_10515);
nand U11189 (N_11189,N_10526,N_10876);
or U11190 (N_11190,N_10783,N_10719);
nand U11191 (N_11191,N_10878,N_10647);
and U11192 (N_11192,N_10949,N_10618);
nand U11193 (N_11193,N_10745,N_10806);
and U11194 (N_11194,N_10512,N_10591);
nor U11195 (N_11195,N_10913,N_10923);
nand U11196 (N_11196,N_10764,N_10741);
nand U11197 (N_11197,N_10743,N_10687);
or U11198 (N_11198,N_10895,N_10579);
and U11199 (N_11199,N_10952,N_10731);
nor U11200 (N_11200,N_10892,N_10879);
or U11201 (N_11201,N_10644,N_10698);
or U11202 (N_11202,N_10677,N_10799);
nand U11203 (N_11203,N_10931,N_10571);
or U11204 (N_11204,N_10561,N_10816);
nand U11205 (N_11205,N_10707,N_10938);
nor U11206 (N_11206,N_10530,N_10762);
and U11207 (N_11207,N_10662,N_10718);
nand U11208 (N_11208,N_10924,N_10672);
or U11209 (N_11209,N_10926,N_10599);
nand U11210 (N_11210,N_10578,N_10999);
and U11211 (N_11211,N_10901,N_10843);
or U11212 (N_11212,N_10593,N_10637);
and U11213 (N_11213,N_10951,N_10910);
or U11214 (N_11214,N_10617,N_10782);
nor U11215 (N_11215,N_10836,N_10809);
xnor U11216 (N_11216,N_10807,N_10874);
xor U11217 (N_11217,N_10982,N_10826);
or U11218 (N_11218,N_10781,N_10849);
nand U11219 (N_11219,N_10596,N_10891);
and U11220 (N_11220,N_10569,N_10965);
nand U11221 (N_11221,N_10519,N_10642);
nor U11222 (N_11222,N_10676,N_10934);
nand U11223 (N_11223,N_10953,N_10880);
and U11224 (N_11224,N_10602,N_10657);
and U11225 (N_11225,N_10768,N_10656);
nand U11226 (N_11226,N_10748,N_10614);
and U11227 (N_11227,N_10793,N_10688);
or U11228 (N_11228,N_10840,N_10950);
and U11229 (N_11229,N_10959,N_10855);
nor U11230 (N_11230,N_10761,N_10525);
nand U11231 (N_11231,N_10511,N_10786);
nand U11232 (N_11232,N_10896,N_10825);
or U11233 (N_11233,N_10802,N_10565);
nand U11234 (N_11234,N_10584,N_10621);
or U11235 (N_11235,N_10697,N_10890);
and U11236 (N_11236,N_10753,N_10979);
nand U11237 (N_11237,N_10920,N_10928);
or U11238 (N_11238,N_10622,N_10605);
nand U11239 (N_11239,N_10503,N_10522);
and U11240 (N_11240,N_10510,N_10508);
and U11241 (N_11241,N_10554,N_10801);
and U11242 (N_11242,N_10902,N_10566);
and U11243 (N_11243,N_10580,N_10691);
nand U11244 (N_11244,N_10869,N_10942);
nor U11245 (N_11245,N_10721,N_10548);
nand U11246 (N_11246,N_10899,N_10988);
nand U11247 (N_11247,N_10989,N_10600);
or U11248 (N_11248,N_10971,N_10654);
nor U11249 (N_11249,N_10568,N_10937);
or U11250 (N_11250,N_10793,N_10672);
and U11251 (N_11251,N_10747,N_10590);
and U11252 (N_11252,N_10751,N_10613);
or U11253 (N_11253,N_10675,N_10632);
and U11254 (N_11254,N_10589,N_10957);
nor U11255 (N_11255,N_10783,N_10935);
nor U11256 (N_11256,N_10828,N_10577);
and U11257 (N_11257,N_10589,N_10795);
or U11258 (N_11258,N_10833,N_10794);
or U11259 (N_11259,N_10532,N_10557);
nor U11260 (N_11260,N_10700,N_10994);
and U11261 (N_11261,N_10583,N_10936);
and U11262 (N_11262,N_10517,N_10797);
or U11263 (N_11263,N_10831,N_10749);
nand U11264 (N_11264,N_10905,N_10647);
or U11265 (N_11265,N_10537,N_10912);
nand U11266 (N_11266,N_10572,N_10942);
or U11267 (N_11267,N_10693,N_10995);
and U11268 (N_11268,N_10883,N_10609);
and U11269 (N_11269,N_10647,N_10529);
xor U11270 (N_11270,N_10879,N_10860);
nor U11271 (N_11271,N_10610,N_10609);
nor U11272 (N_11272,N_10549,N_10786);
nand U11273 (N_11273,N_10772,N_10903);
nor U11274 (N_11274,N_10935,N_10763);
nor U11275 (N_11275,N_10662,N_10558);
and U11276 (N_11276,N_10998,N_10672);
nand U11277 (N_11277,N_10795,N_10663);
nor U11278 (N_11278,N_10620,N_10712);
nand U11279 (N_11279,N_10979,N_10988);
and U11280 (N_11280,N_10649,N_10988);
and U11281 (N_11281,N_10805,N_10612);
nor U11282 (N_11282,N_10774,N_10753);
or U11283 (N_11283,N_10889,N_10505);
or U11284 (N_11284,N_10580,N_10649);
nand U11285 (N_11285,N_10727,N_10591);
and U11286 (N_11286,N_10552,N_10906);
and U11287 (N_11287,N_10701,N_10590);
or U11288 (N_11288,N_10668,N_10685);
and U11289 (N_11289,N_10937,N_10929);
or U11290 (N_11290,N_10694,N_10770);
nand U11291 (N_11291,N_10758,N_10990);
and U11292 (N_11292,N_10576,N_10979);
xor U11293 (N_11293,N_10523,N_10551);
or U11294 (N_11294,N_10838,N_10941);
and U11295 (N_11295,N_10511,N_10813);
nor U11296 (N_11296,N_10726,N_10616);
and U11297 (N_11297,N_10992,N_10602);
or U11298 (N_11298,N_10684,N_10886);
nor U11299 (N_11299,N_10657,N_10967);
nand U11300 (N_11300,N_10682,N_10878);
xnor U11301 (N_11301,N_10545,N_10868);
or U11302 (N_11302,N_10662,N_10669);
nand U11303 (N_11303,N_10898,N_10543);
or U11304 (N_11304,N_10549,N_10963);
nor U11305 (N_11305,N_10839,N_10780);
nor U11306 (N_11306,N_10681,N_10532);
and U11307 (N_11307,N_10846,N_10836);
nand U11308 (N_11308,N_10849,N_10862);
and U11309 (N_11309,N_10587,N_10615);
nor U11310 (N_11310,N_10564,N_10629);
nand U11311 (N_11311,N_10705,N_10703);
nor U11312 (N_11312,N_10963,N_10594);
nand U11313 (N_11313,N_10504,N_10591);
nand U11314 (N_11314,N_10500,N_10749);
nand U11315 (N_11315,N_10876,N_10755);
and U11316 (N_11316,N_10525,N_10537);
and U11317 (N_11317,N_10699,N_10683);
and U11318 (N_11318,N_10945,N_10998);
xnor U11319 (N_11319,N_10774,N_10995);
or U11320 (N_11320,N_10694,N_10522);
nand U11321 (N_11321,N_10726,N_10986);
and U11322 (N_11322,N_10620,N_10708);
or U11323 (N_11323,N_10626,N_10775);
nand U11324 (N_11324,N_10648,N_10779);
and U11325 (N_11325,N_10782,N_10835);
or U11326 (N_11326,N_10933,N_10998);
nand U11327 (N_11327,N_10788,N_10515);
and U11328 (N_11328,N_10660,N_10649);
nor U11329 (N_11329,N_10618,N_10955);
or U11330 (N_11330,N_10710,N_10983);
or U11331 (N_11331,N_10731,N_10968);
or U11332 (N_11332,N_10766,N_10642);
nor U11333 (N_11333,N_10702,N_10615);
nor U11334 (N_11334,N_10613,N_10975);
nor U11335 (N_11335,N_10897,N_10972);
nor U11336 (N_11336,N_10657,N_10821);
or U11337 (N_11337,N_10761,N_10895);
or U11338 (N_11338,N_10864,N_10948);
nand U11339 (N_11339,N_10816,N_10804);
and U11340 (N_11340,N_10855,N_10975);
nor U11341 (N_11341,N_10569,N_10534);
nand U11342 (N_11342,N_10903,N_10804);
and U11343 (N_11343,N_10544,N_10516);
and U11344 (N_11344,N_10533,N_10808);
nand U11345 (N_11345,N_10997,N_10980);
nor U11346 (N_11346,N_10553,N_10578);
or U11347 (N_11347,N_10787,N_10926);
or U11348 (N_11348,N_10905,N_10885);
or U11349 (N_11349,N_10953,N_10797);
nor U11350 (N_11350,N_10643,N_10528);
and U11351 (N_11351,N_10860,N_10795);
nand U11352 (N_11352,N_10849,N_10949);
nand U11353 (N_11353,N_10555,N_10753);
xnor U11354 (N_11354,N_10719,N_10790);
nand U11355 (N_11355,N_10608,N_10712);
and U11356 (N_11356,N_10526,N_10628);
xnor U11357 (N_11357,N_10708,N_10678);
nor U11358 (N_11358,N_10780,N_10919);
or U11359 (N_11359,N_10770,N_10506);
nor U11360 (N_11360,N_10868,N_10846);
or U11361 (N_11361,N_10693,N_10563);
nand U11362 (N_11362,N_10975,N_10653);
and U11363 (N_11363,N_10993,N_10930);
nand U11364 (N_11364,N_10935,N_10637);
and U11365 (N_11365,N_10658,N_10574);
and U11366 (N_11366,N_10891,N_10555);
or U11367 (N_11367,N_10957,N_10682);
and U11368 (N_11368,N_10503,N_10950);
and U11369 (N_11369,N_10560,N_10836);
nor U11370 (N_11370,N_10899,N_10553);
or U11371 (N_11371,N_10894,N_10758);
nand U11372 (N_11372,N_10629,N_10646);
nand U11373 (N_11373,N_10903,N_10952);
and U11374 (N_11374,N_10994,N_10557);
nand U11375 (N_11375,N_10536,N_10713);
nand U11376 (N_11376,N_10932,N_10983);
or U11377 (N_11377,N_10841,N_10676);
nor U11378 (N_11378,N_10504,N_10533);
or U11379 (N_11379,N_10775,N_10835);
and U11380 (N_11380,N_10927,N_10866);
and U11381 (N_11381,N_10612,N_10522);
nor U11382 (N_11382,N_10524,N_10600);
or U11383 (N_11383,N_10527,N_10601);
nor U11384 (N_11384,N_10837,N_10529);
nand U11385 (N_11385,N_10672,N_10881);
or U11386 (N_11386,N_10639,N_10553);
or U11387 (N_11387,N_10815,N_10634);
and U11388 (N_11388,N_10774,N_10690);
or U11389 (N_11389,N_10768,N_10841);
nor U11390 (N_11390,N_10661,N_10620);
or U11391 (N_11391,N_10613,N_10807);
or U11392 (N_11392,N_10746,N_10902);
or U11393 (N_11393,N_10801,N_10570);
nor U11394 (N_11394,N_10774,N_10607);
nand U11395 (N_11395,N_10661,N_10791);
nand U11396 (N_11396,N_10509,N_10704);
nand U11397 (N_11397,N_10937,N_10932);
or U11398 (N_11398,N_10978,N_10998);
nand U11399 (N_11399,N_10615,N_10590);
nor U11400 (N_11400,N_10781,N_10719);
nor U11401 (N_11401,N_10661,N_10517);
nor U11402 (N_11402,N_10662,N_10990);
and U11403 (N_11403,N_10580,N_10508);
nor U11404 (N_11404,N_10524,N_10633);
and U11405 (N_11405,N_10564,N_10804);
nand U11406 (N_11406,N_10698,N_10517);
and U11407 (N_11407,N_10857,N_10774);
and U11408 (N_11408,N_10905,N_10728);
and U11409 (N_11409,N_10818,N_10992);
or U11410 (N_11410,N_10866,N_10512);
nor U11411 (N_11411,N_10881,N_10836);
nand U11412 (N_11412,N_10851,N_10764);
nand U11413 (N_11413,N_10757,N_10732);
nand U11414 (N_11414,N_10984,N_10906);
and U11415 (N_11415,N_10634,N_10560);
nor U11416 (N_11416,N_10874,N_10800);
nand U11417 (N_11417,N_10809,N_10729);
and U11418 (N_11418,N_10731,N_10524);
or U11419 (N_11419,N_10642,N_10989);
nand U11420 (N_11420,N_10975,N_10543);
nand U11421 (N_11421,N_10853,N_10682);
and U11422 (N_11422,N_10584,N_10840);
nor U11423 (N_11423,N_10655,N_10562);
nand U11424 (N_11424,N_10986,N_10906);
or U11425 (N_11425,N_10573,N_10671);
nor U11426 (N_11426,N_10733,N_10693);
or U11427 (N_11427,N_10529,N_10915);
xor U11428 (N_11428,N_10792,N_10504);
nor U11429 (N_11429,N_10850,N_10533);
and U11430 (N_11430,N_10622,N_10722);
and U11431 (N_11431,N_10979,N_10578);
or U11432 (N_11432,N_10916,N_10609);
and U11433 (N_11433,N_10689,N_10726);
nor U11434 (N_11434,N_10723,N_10908);
nor U11435 (N_11435,N_10861,N_10514);
nand U11436 (N_11436,N_10713,N_10967);
nor U11437 (N_11437,N_10856,N_10520);
and U11438 (N_11438,N_10647,N_10994);
nor U11439 (N_11439,N_10896,N_10561);
nor U11440 (N_11440,N_10919,N_10640);
or U11441 (N_11441,N_10958,N_10560);
or U11442 (N_11442,N_10739,N_10965);
nand U11443 (N_11443,N_10606,N_10531);
nand U11444 (N_11444,N_10715,N_10682);
xnor U11445 (N_11445,N_10940,N_10725);
nor U11446 (N_11446,N_10650,N_10742);
nand U11447 (N_11447,N_10750,N_10763);
nand U11448 (N_11448,N_10516,N_10682);
nor U11449 (N_11449,N_10944,N_10900);
nand U11450 (N_11450,N_10913,N_10718);
nor U11451 (N_11451,N_10561,N_10962);
and U11452 (N_11452,N_10557,N_10702);
and U11453 (N_11453,N_10871,N_10717);
nand U11454 (N_11454,N_10943,N_10826);
nand U11455 (N_11455,N_10786,N_10815);
or U11456 (N_11456,N_10938,N_10831);
nor U11457 (N_11457,N_10927,N_10678);
nor U11458 (N_11458,N_10565,N_10591);
and U11459 (N_11459,N_10611,N_10853);
xnor U11460 (N_11460,N_10769,N_10744);
nor U11461 (N_11461,N_10768,N_10531);
or U11462 (N_11462,N_10910,N_10673);
and U11463 (N_11463,N_10795,N_10878);
and U11464 (N_11464,N_10754,N_10636);
nand U11465 (N_11465,N_10802,N_10879);
nand U11466 (N_11466,N_10720,N_10608);
nand U11467 (N_11467,N_10770,N_10683);
nand U11468 (N_11468,N_10947,N_10837);
nand U11469 (N_11469,N_10934,N_10822);
and U11470 (N_11470,N_10721,N_10569);
nand U11471 (N_11471,N_10819,N_10728);
nand U11472 (N_11472,N_10686,N_10622);
or U11473 (N_11473,N_10633,N_10962);
nor U11474 (N_11474,N_10754,N_10941);
or U11475 (N_11475,N_10783,N_10893);
or U11476 (N_11476,N_10539,N_10972);
nor U11477 (N_11477,N_10702,N_10736);
nand U11478 (N_11478,N_10689,N_10900);
or U11479 (N_11479,N_10716,N_10806);
xnor U11480 (N_11480,N_10553,N_10927);
or U11481 (N_11481,N_10882,N_10589);
nor U11482 (N_11482,N_10540,N_10962);
nand U11483 (N_11483,N_10938,N_10797);
nor U11484 (N_11484,N_10737,N_10967);
xnor U11485 (N_11485,N_10611,N_10793);
nor U11486 (N_11486,N_10931,N_10867);
nor U11487 (N_11487,N_10544,N_10826);
nor U11488 (N_11488,N_10758,N_10535);
and U11489 (N_11489,N_10637,N_10598);
and U11490 (N_11490,N_10959,N_10514);
nor U11491 (N_11491,N_10860,N_10577);
nor U11492 (N_11492,N_10929,N_10928);
or U11493 (N_11493,N_10878,N_10891);
nor U11494 (N_11494,N_10954,N_10985);
nor U11495 (N_11495,N_10650,N_10692);
nor U11496 (N_11496,N_10662,N_10861);
nor U11497 (N_11497,N_10855,N_10609);
xor U11498 (N_11498,N_10577,N_10939);
and U11499 (N_11499,N_10965,N_10718);
and U11500 (N_11500,N_11487,N_11334);
or U11501 (N_11501,N_11303,N_11025);
nand U11502 (N_11502,N_11309,N_11445);
nor U11503 (N_11503,N_11053,N_11114);
xor U11504 (N_11504,N_11351,N_11472);
or U11505 (N_11505,N_11086,N_11227);
or U11506 (N_11506,N_11450,N_11352);
nor U11507 (N_11507,N_11387,N_11207);
and U11508 (N_11508,N_11278,N_11170);
nor U11509 (N_11509,N_11435,N_11331);
nand U11510 (N_11510,N_11413,N_11267);
and U11511 (N_11511,N_11168,N_11266);
and U11512 (N_11512,N_11046,N_11084);
nor U11513 (N_11513,N_11483,N_11393);
nor U11514 (N_11514,N_11213,N_11332);
and U11515 (N_11515,N_11191,N_11252);
nor U11516 (N_11516,N_11100,N_11087);
nor U11517 (N_11517,N_11109,N_11263);
or U11518 (N_11518,N_11117,N_11382);
nor U11519 (N_11519,N_11036,N_11482);
nor U11520 (N_11520,N_11014,N_11449);
or U11521 (N_11521,N_11237,N_11074);
or U11522 (N_11522,N_11369,N_11041);
or U11523 (N_11523,N_11268,N_11405);
or U11524 (N_11524,N_11419,N_11121);
or U11525 (N_11525,N_11307,N_11188);
nand U11526 (N_11526,N_11443,N_11200);
nand U11527 (N_11527,N_11427,N_11283);
nand U11528 (N_11528,N_11002,N_11302);
xnor U11529 (N_11529,N_11239,N_11498);
nand U11530 (N_11530,N_11226,N_11313);
nand U11531 (N_11531,N_11253,N_11490);
and U11532 (N_11532,N_11311,N_11330);
and U11533 (N_11533,N_11447,N_11143);
xnor U11534 (N_11534,N_11156,N_11485);
nand U11535 (N_11535,N_11315,N_11214);
and U11536 (N_11536,N_11107,N_11178);
nor U11537 (N_11537,N_11030,N_11415);
nand U11538 (N_11538,N_11059,N_11383);
or U11539 (N_11539,N_11098,N_11069);
nor U11540 (N_11540,N_11115,N_11306);
nand U11541 (N_11541,N_11495,N_11029);
nor U11542 (N_11542,N_11328,N_11094);
nand U11543 (N_11543,N_11265,N_11397);
xor U11544 (N_11544,N_11368,N_11391);
nor U11545 (N_11545,N_11080,N_11233);
xnor U11546 (N_11546,N_11050,N_11219);
nand U11547 (N_11547,N_11335,N_11235);
nand U11548 (N_11548,N_11297,N_11499);
or U11549 (N_11549,N_11139,N_11051);
and U11550 (N_11550,N_11476,N_11055);
nor U11551 (N_11551,N_11011,N_11097);
or U11552 (N_11552,N_11392,N_11079);
or U11553 (N_11553,N_11039,N_11007);
nor U11554 (N_11554,N_11018,N_11385);
nand U11555 (N_11555,N_11316,N_11367);
and U11556 (N_11556,N_11292,N_11095);
nand U11557 (N_11557,N_11416,N_11257);
nor U11558 (N_11558,N_11293,N_11269);
or U11559 (N_11559,N_11323,N_11158);
nand U11560 (N_11560,N_11091,N_11048);
nand U11561 (N_11561,N_11439,N_11128);
or U11562 (N_11562,N_11338,N_11388);
nand U11563 (N_11563,N_11221,N_11040);
nor U11564 (N_11564,N_11333,N_11364);
nor U11565 (N_11565,N_11035,N_11058);
nor U11566 (N_11566,N_11061,N_11147);
or U11567 (N_11567,N_11277,N_11026);
and U11568 (N_11568,N_11358,N_11197);
or U11569 (N_11569,N_11099,N_11248);
nand U11570 (N_11570,N_11123,N_11144);
or U11571 (N_11571,N_11111,N_11344);
and U11572 (N_11572,N_11361,N_11125);
nor U11573 (N_11573,N_11324,N_11149);
and U11574 (N_11574,N_11337,N_11258);
and U11575 (N_11575,N_11142,N_11438);
nand U11576 (N_11576,N_11282,N_11470);
nor U11577 (N_11577,N_11310,N_11436);
and U11578 (N_11578,N_11196,N_11118);
and U11579 (N_11579,N_11464,N_11017);
and U11580 (N_11580,N_11373,N_11187);
or U11581 (N_11581,N_11384,N_11246);
nor U11582 (N_11582,N_11215,N_11120);
nand U11583 (N_11583,N_11360,N_11295);
nand U11584 (N_11584,N_11045,N_11174);
or U11585 (N_11585,N_11318,N_11232);
and U11586 (N_11586,N_11060,N_11243);
and U11587 (N_11587,N_11262,N_11294);
and U11588 (N_11588,N_11299,N_11418);
nand U11589 (N_11589,N_11380,N_11096);
nor U11590 (N_11590,N_11083,N_11461);
and U11591 (N_11591,N_11440,N_11212);
nand U11592 (N_11592,N_11127,N_11350);
or U11593 (N_11593,N_11071,N_11027);
nand U11594 (N_11594,N_11455,N_11157);
nor U11595 (N_11595,N_11231,N_11122);
nor U11596 (N_11596,N_11280,N_11329);
and U11597 (N_11597,N_11028,N_11112);
nor U11598 (N_11598,N_11291,N_11210);
or U11599 (N_11599,N_11494,N_11363);
or U11600 (N_11600,N_11167,N_11463);
and U11601 (N_11601,N_11459,N_11377);
or U11602 (N_11602,N_11275,N_11371);
nand U11603 (N_11603,N_11468,N_11421);
and U11604 (N_11604,N_11005,N_11024);
or U11605 (N_11605,N_11285,N_11209);
nor U11606 (N_11606,N_11240,N_11396);
nand U11607 (N_11607,N_11153,N_11003);
nor U11608 (N_11608,N_11346,N_11223);
or U11609 (N_11609,N_11204,N_11001);
nand U11610 (N_11610,N_11013,N_11211);
or U11611 (N_11611,N_11406,N_11010);
nand U11612 (N_11612,N_11376,N_11130);
nand U11613 (N_11613,N_11177,N_11065);
nor U11614 (N_11614,N_11261,N_11032);
nand U11615 (N_11615,N_11473,N_11217);
or U11616 (N_11616,N_11417,N_11356);
and U11617 (N_11617,N_11260,N_11366);
xor U11618 (N_11618,N_11184,N_11116);
nand U11619 (N_11619,N_11251,N_11090);
or U11620 (N_11620,N_11195,N_11172);
or U11621 (N_11621,N_11180,N_11199);
nor U11622 (N_11622,N_11414,N_11326);
nand U11623 (N_11623,N_11192,N_11437);
xor U11624 (N_11624,N_11386,N_11428);
nand U11625 (N_11625,N_11300,N_11342);
or U11626 (N_11626,N_11401,N_11343);
xnor U11627 (N_11627,N_11327,N_11247);
or U11628 (N_11628,N_11425,N_11359);
or U11629 (N_11629,N_11379,N_11113);
nor U11630 (N_11630,N_11161,N_11457);
nor U11631 (N_11631,N_11370,N_11137);
nor U11632 (N_11632,N_11155,N_11190);
nor U11633 (N_11633,N_11082,N_11365);
nor U11634 (N_11634,N_11408,N_11076);
nor U11635 (N_11635,N_11471,N_11341);
and U11636 (N_11636,N_11133,N_11110);
and U11637 (N_11637,N_11474,N_11467);
or U11638 (N_11638,N_11272,N_11395);
nand U11639 (N_11639,N_11104,N_11288);
and U11640 (N_11640,N_11466,N_11321);
or U11641 (N_11641,N_11006,N_11453);
and U11642 (N_11642,N_11208,N_11189);
or U11643 (N_11643,N_11353,N_11420);
or U11644 (N_11644,N_11254,N_11194);
nand U11645 (N_11645,N_11159,N_11398);
nor U11646 (N_11646,N_11012,N_11234);
or U11647 (N_11647,N_11102,N_11236);
or U11648 (N_11648,N_11312,N_11179);
nand U11649 (N_11649,N_11052,N_11340);
nor U11650 (N_11650,N_11484,N_11290);
nor U11651 (N_11651,N_11070,N_11108);
nor U11652 (N_11652,N_11452,N_11429);
nand U11653 (N_11653,N_11164,N_11374);
nand U11654 (N_11654,N_11412,N_11442);
nor U11655 (N_11655,N_11270,N_11322);
xor U11656 (N_11656,N_11238,N_11357);
or U11657 (N_11657,N_11230,N_11255);
and U11658 (N_11658,N_11296,N_11066);
and U11659 (N_11659,N_11347,N_11441);
and U11660 (N_11660,N_11206,N_11446);
nand U11661 (N_11661,N_11222,N_11336);
or U11662 (N_11662,N_11286,N_11033);
and U11663 (N_11663,N_11201,N_11148);
nor U11664 (N_11664,N_11444,N_11354);
nor U11665 (N_11665,N_11456,N_11085);
nor U11666 (N_11666,N_11081,N_11182);
and U11667 (N_11667,N_11093,N_11454);
and U11668 (N_11668,N_11362,N_11228);
and U11669 (N_11669,N_11281,N_11349);
nand U11670 (N_11670,N_11478,N_11432);
or U11671 (N_11671,N_11043,N_11403);
nor U11672 (N_11672,N_11038,N_11193);
and U11673 (N_11673,N_11119,N_11103);
xnor U11674 (N_11674,N_11105,N_11497);
or U11675 (N_11675,N_11244,N_11134);
nor U11676 (N_11676,N_11430,N_11245);
nand U11677 (N_11677,N_11078,N_11220);
nor U11678 (N_11678,N_11410,N_11073);
nor U11679 (N_11679,N_11250,N_11274);
nand U11680 (N_11680,N_11462,N_11169);
or U11681 (N_11681,N_11020,N_11150);
nor U11682 (N_11682,N_11422,N_11241);
and U11683 (N_11683,N_11037,N_11314);
nand U11684 (N_11684,N_11229,N_11000);
nor U11685 (N_11685,N_11031,N_11493);
or U11686 (N_11686,N_11325,N_11047);
nor U11687 (N_11687,N_11273,N_11101);
nand U11688 (N_11688,N_11400,N_11279);
nor U11689 (N_11689,N_11381,N_11138);
or U11690 (N_11690,N_11092,N_11259);
or U11691 (N_11691,N_11448,N_11481);
nand U11692 (N_11692,N_11173,N_11126);
nor U11693 (N_11693,N_11488,N_11489);
or U11694 (N_11694,N_11433,N_11140);
or U11695 (N_11695,N_11339,N_11106);
nor U11696 (N_11696,N_11480,N_11034);
or U11697 (N_11697,N_11152,N_11141);
or U11698 (N_11698,N_11064,N_11469);
or U11699 (N_11699,N_11008,N_11271);
or U11700 (N_11700,N_11077,N_11063);
nor U11701 (N_11701,N_11399,N_11287);
nand U11702 (N_11702,N_11072,N_11264);
nor U11703 (N_11703,N_11320,N_11019);
and U11704 (N_11704,N_11372,N_11319);
nor U11705 (N_11705,N_11056,N_11460);
or U11706 (N_11706,N_11062,N_11289);
and U11707 (N_11707,N_11205,N_11394);
and U11708 (N_11708,N_11426,N_11375);
nor U11709 (N_11709,N_11402,N_11160);
or U11710 (N_11710,N_11203,N_11424);
and U11711 (N_11711,N_11411,N_11166);
nand U11712 (N_11712,N_11404,N_11496);
or U11713 (N_11713,N_11256,N_11458);
nor U11714 (N_11714,N_11049,N_11162);
or U11715 (N_11715,N_11491,N_11124);
nand U11716 (N_11716,N_11042,N_11216);
nor U11717 (N_11717,N_11089,N_11015);
or U11718 (N_11718,N_11298,N_11431);
and U11719 (N_11719,N_11304,N_11378);
and U11720 (N_11720,N_11345,N_11183);
nor U11721 (N_11721,N_11423,N_11317);
or U11722 (N_11722,N_11475,N_11186);
and U11723 (N_11723,N_11218,N_11154);
and U11724 (N_11724,N_11301,N_11175);
and U11725 (N_11725,N_11171,N_11390);
or U11726 (N_11726,N_11198,N_11486);
and U11727 (N_11727,N_11242,N_11044);
or U11728 (N_11728,N_11129,N_11492);
nand U11729 (N_11729,N_11135,N_11068);
xnor U11730 (N_11730,N_11407,N_11145);
and U11731 (N_11731,N_11249,N_11004);
or U11732 (N_11732,N_11308,N_11477);
nand U11733 (N_11733,N_11284,N_11409);
and U11734 (N_11734,N_11131,N_11057);
and U11735 (N_11735,N_11355,N_11009);
or U11736 (N_11736,N_11348,N_11151);
nand U11737 (N_11737,N_11016,N_11132);
nand U11738 (N_11738,N_11022,N_11479);
nor U11739 (N_11739,N_11075,N_11451);
nand U11740 (N_11740,N_11225,N_11181);
nor U11741 (N_11741,N_11165,N_11146);
and U11742 (N_11742,N_11163,N_11023);
nor U11743 (N_11743,N_11176,N_11276);
nor U11744 (N_11744,N_11054,N_11088);
nand U11745 (N_11745,N_11434,N_11202);
or U11746 (N_11746,N_11136,N_11465);
nand U11747 (N_11747,N_11185,N_11389);
xnor U11748 (N_11748,N_11067,N_11021);
and U11749 (N_11749,N_11224,N_11305);
nand U11750 (N_11750,N_11069,N_11493);
nand U11751 (N_11751,N_11331,N_11203);
or U11752 (N_11752,N_11166,N_11464);
xor U11753 (N_11753,N_11363,N_11423);
or U11754 (N_11754,N_11265,N_11083);
nor U11755 (N_11755,N_11303,N_11351);
and U11756 (N_11756,N_11466,N_11056);
or U11757 (N_11757,N_11039,N_11095);
nand U11758 (N_11758,N_11327,N_11097);
nand U11759 (N_11759,N_11362,N_11322);
or U11760 (N_11760,N_11476,N_11463);
and U11761 (N_11761,N_11239,N_11449);
nand U11762 (N_11762,N_11075,N_11019);
nand U11763 (N_11763,N_11340,N_11401);
and U11764 (N_11764,N_11273,N_11429);
or U11765 (N_11765,N_11368,N_11218);
and U11766 (N_11766,N_11037,N_11332);
nand U11767 (N_11767,N_11403,N_11267);
or U11768 (N_11768,N_11049,N_11002);
nand U11769 (N_11769,N_11450,N_11039);
nor U11770 (N_11770,N_11035,N_11228);
or U11771 (N_11771,N_11054,N_11493);
or U11772 (N_11772,N_11418,N_11045);
nand U11773 (N_11773,N_11329,N_11373);
nand U11774 (N_11774,N_11367,N_11433);
nand U11775 (N_11775,N_11042,N_11444);
nor U11776 (N_11776,N_11181,N_11315);
or U11777 (N_11777,N_11466,N_11129);
or U11778 (N_11778,N_11453,N_11331);
nor U11779 (N_11779,N_11434,N_11269);
and U11780 (N_11780,N_11363,N_11145);
or U11781 (N_11781,N_11040,N_11212);
nand U11782 (N_11782,N_11392,N_11373);
nand U11783 (N_11783,N_11158,N_11438);
nor U11784 (N_11784,N_11172,N_11454);
nand U11785 (N_11785,N_11265,N_11341);
nor U11786 (N_11786,N_11279,N_11495);
or U11787 (N_11787,N_11360,N_11073);
and U11788 (N_11788,N_11221,N_11458);
nand U11789 (N_11789,N_11199,N_11124);
nor U11790 (N_11790,N_11186,N_11448);
nand U11791 (N_11791,N_11274,N_11409);
nor U11792 (N_11792,N_11109,N_11491);
nor U11793 (N_11793,N_11254,N_11170);
or U11794 (N_11794,N_11391,N_11177);
and U11795 (N_11795,N_11134,N_11304);
nor U11796 (N_11796,N_11365,N_11334);
or U11797 (N_11797,N_11180,N_11050);
or U11798 (N_11798,N_11334,N_11235);
nand U11799 (N_11799,N_11417,N_11031);
nor U11800 (N_11800,N_11422,N_11381);
or U11801 (N_11801,N_11128,N_11231);
and U11802 (N_11802,N_11305,N_11454);
or U11803 (N_11803,N_11151,N_11204);
nor U11804 (N_11804,N_11128,N_11336);
or U11805 (N_11805,N_11112,N_11050);
or U11806 (N_11806,N_11231,N_11486);
or U11807 (N_11807,N_11010,N_11438);
xnor U11808 (N_11808,N_11185,N_11448);
nand U11809 (N_11809,N_11362,N_11278);
and U11810 (N_11810,N_11389,N_11382);
nor U11811 (N_11811,N_11152,N_11179);
and U11812 (N_11812,N_11208,N_11096);
nand U11813 (N_11813,N_11034,N_11152);
and U11814 (N_11814,N_11404,N_11330);
or U11815 (N_11815,N_11286,N_11067);
or U11816 (N_11816,N_11115,N_11104);
nand U11817 (N_11817,N_11122,N_11246);
nand U11818 (N_11818,N_11255,N_11102);
or U11819 (N_11819,N_11443,N_11238);
or U11820 (N_11820,N_11204,N_11033);
nor U11821 (N_11821,N_11239,N_11304);
nand U11822 (N_11822,N_11076,N_11424);
or U11823 (N_11823,N_11302,N_11138);
or U11824 (N_11824,N_11151,N_11072);
or U11825 (N_11825,N_11149,N_11125);
nor U11826 (N_11826,N_11439,N_11321);
and U11827 (N_11827,N_11241,N_11230);
or U11828 (N_11828,N_11244,N_11461);
nor U11829 (N_11829,N_11260,N_11236);
and U11830 (N_11830,N_11470,N_11401);
and U11831 (N_11831,N_11311,N_11342);
nand U11832 (N_11832,N_11489,N_11353);
nor U11833 (N_11833,N_11441,N_11481);
nor U11834 (N_11834,N_11321,N_11079);
and U11835 (N_11835,N_11324,N_11018);
nor U11836 (N_11836,N_11114,N_11042);
and U11837 (N_11837,N_11383,N_11250);
and U11838 (N_11838,N_11106,N_11460);
and U11839 (N_11839,N_11237,N_11104);
nor U11840 (N_11840,N_11224,N_11339);
nand U11841 (N_11841,N_11448,N_11445);
or U11842 (N_11842,N_11465,N_11491);
nor U11843 (N_11843,N_11337,N_11266);
nand U11844 (N_11844,N_11006,N_11092);
and U11845 (N_11845,N_11163,N_11168);
nand U11846 (N_11846,N_11440,N_11041);
nand U11847 (N_11847,N_11208,N_11120);
nor U11848 (N_11848,N_11028,N_11036);
nor U11849 (N_11849,N_11290,N_11226);
or U11850 (N_11850,N_11387,N_11148);
and U11851 (N_11851,N_11494,N_11250);
nand U11852 (N_11852,N_11134,N_11210);
and U11853 (N_11853,N_11245,N_11127);
or U11854 (N_11854,N_11060,N_11438);
nand U11855 (N_11855,N_11193,N_11334);
nand U11856 (N_11856,N_11016,N_11332);
nand U11857 (N_11857,N_11451,N_11429);
and U11858 (N_11858,N_11295,N_11299);
and U11859 (N_11859,N_11140,N_11082);
nor U11860 (N_11860,N_11175,N_11152);
nand U11861 (N_11861,N_11319,N_11248);
and U11862 (N_11862,N_11440,N_11468);
nor U11863 (N_11863,N_11118,N_11462);
nand U11864 (N_11864,N_11140,N_11262);
nor U11865 (N_11865,N_11383,N_11116);
nand U11866 (N_11866,N_11067,N_11150);
nor U11867 (N_11867,N_11336,N_11226);
xnor U11868 (N_11868,N_11023,N_11377);
nand U11869 (N_11869,N_11061,N_11451);
and U11870 (N_11870,N_11344,N_11490);
nand U11871 (N_11871,N_11151,N_11404);
nand U11872 (N_11872,N_11019,N_11454);
and U11873 (N_11873,N_11309,N_11466);
or U11874 (N_11874,N_11151,N_11225);
nor U11875 (N_11875,N_11199,N_11186);
or U11876 (N_11876,N_11465,N_11101);
or U11877 (N_11877,N_11270,N_11014);
nor U11878 (N_11878,N_11311,N_11450);
nand U11879 (N_11879,N_11372,N_11472);
nand U11880 (N_11880,N_11390,N_11214);
nor U11881 (N_11881,N_11038,N_11412);
nand U11882 (N_11882,N_11464,N_11201);
nand U11883 (N_11883,N_11045,N_11462);
and U11884 (N_11884,N_11397,N_11148);
nand U11885 (N_11885,N_11042,N_11105);
and U11886 (N_11886,N_11335,N_11432);
and U11887 (N_11887,N_11180,N_11257);
nand U11888 (N_11888,N_11196,N_11267);
nor U11889 (N_11889,N_11458,N_11379);
nor U11890 (N_11890,N_11493,N_11180);
nor U11891 (N_11891,N_11210,N_11393);
or U11892 (N_11892,N_11188,N_11422);
nor U11893 (N_11893,N_11144,N_11063);
xor U11894 (N_11894,N_11023,N_11489);
nor U11895 (N_11895,N_11127,N_11133);
or U11896 (N_11896,N_11203,N_11276);
or U11897 (N_11897,N_11299,N_11372);
and U11898 (N_11898,N_11089,N_11436);
xnor U11899 (N_11899,N_11068,N_11014);
or U11900 (N_11900,N_11132,N_11010);
or U11901 (N_11901,N_11376,N_11439);
and U11902 (N_11902,N_11075,N_11461);
and U11903 (N_11903,N_11061,N_11414);
nand U11904 (N_11904,N_11255,N_11005);
or U11905 (N_11905,N_11268,N_11338);
nor U11906 (N_11906,N_11463,N_11394);
nand U11907 (N_11907,N_11392,N_11465);
nand U11908 (N_11908,N_11061,N_11257);
or U11909 (N_11909,N_11123,N_11430);
and U11910 (N_11910,N_11221,N_11486);
nor U11911 (N_11911,N_11076,N_11361);
nor U11912 (N_11912,N_11404,N_11278);
or U11913 (N_11913,N_11367,N_11306);
and U11914 (N_11914,N_11481,N_11215);
nor U11915 (N_11915,N_11181,N_11342);
nor U11916 (N_11916,N_11108,N_11163);
nor U11917 (N_11917,N_11365,N_11235);
or U11918 (N_11918,N_11421,N_11279);
nor U11919 (N_11919,N_11154,N_11287);
or U11920 (N_11920,N_11099,N_11447);
xor U11921 (N_11921,N_11276,N_11092);
and U11922 (N_11922,N_11252,N_11293);
and U11923 (N_11923,N_11132,N_11200);
or U11924 (N_11924,N_11329,N_11174);
nand U11925 (N_11925,N_11474,N_11126);
nand U11926 (N_11926,N_11077,N_11078);
nor U11927 (N_11927,N_11452,N_11425);
nor U11928 (N_11928,N_11349,N_11134);
nor U11929 (N_11929,N_11231,N_11394);
nand U11930 (N_11930,N_11303,N_11092);
and U11931 (N_11931,N_11444,N_11231);
nand U11932 (N_11932,N_11163,N_11127);
nor U11933 (N_11933,N_11458,N_11124);
nand U11934 (N_11934,N_11299,N_11075);
or U11935 (N_11935,N_11342,N_11341);
or U11936 (N_11936,N_11431,N_11263);
and U11937 (N_11937,N_11181,N_11089);
nor U11938 (N_11938,N_11472,N_11416);
or U11939 (N_11939,N_11413,N_11117);
or U11940 (N_11940,N_11321,N_11415);
and U11941 (N_11941,N_11328,N_11472);
and U11942 (N_11942,N_11308,N_11258);
nand U11943 (N_11943,N_11271,N_11255);
and U11944 (N_11944,N_11378,N_11272);
nor U11945 (N_11945,N_11030,N_11318);
nand U11946 (N_11946,N_11057,N_11025);
nor U11947 (N_11947,N_11251,N_11275);
nand U11948 (N_11948,N_11357,N_11381);
and U11949 (N_11949,N_11113,N_11376);
and U11950 (N_11950,N_11222,N_11335);
and U11951 (N_11951,N_11108,N_11176);
nand U11952 (N_11952,N_11466,N_11114);
and U11953 (N_11953,N_11276,N_11090);
nand U11954 (N_11954,N_11319,N_11370);
and U11955 (N_11955,N_11202,N_11352);
nor U11956 (N_11956,N_11114,N_11420);
and U11957 (N_11957,N_11481,N_11443);
and U11958 (N_11958,N_11442,N_11446);
nand U11959 (N_11959,N_11322,N_11292);
or U11960 (N_11960,N_11082,N_11354);
nor U11961 (N_11961,N_11417,N_11471);
nor U11962 (N_11962,N_11477,N_11079);
or U11963 (N_11963,N_11049,N_11404);
nand U11964 (N_11964,N_11349,N_11381);
nor U11965 (N_11965,N_11183,N_11181);
or U11966 (N_11966,N_11282,N_11034);
nor U11967 (N_11967,N_11242,N_11201);
nand U11968 (N_11968,N_11132,N_11245);
nand U11969 (N_11969,N_11380,N_11382);
or U11970 (N_11970,N_11128,N_11196);
or U11971 (N_11971,N_11016,N_11125);
and U11972 (N_11972,N_11338,N_11110);
and U11973 (N_11973,N_11072,N_11083);
nor U11974 (N_11974,N_11039,N_11306);
nand U11975 (N_11975,N_11472,N_11122);
or U11976 (N_11976,N_11270,N_11150);
nor U11977 (N_11977,N_11350,N_11384);
nor U11978 (N_11978,N_11383,N_11446);
or U11979 (N_11979,N_11015,N_11442);
xor U11980 (N_11980,N_11142,N_11317);
nand U11981 (N_11981,N_11203,N_11248);
nand U11982 (N_11982,N_11483,N_11459);
or U11983 (N_11983,N_11185,N_11375);
nor U11984 (N_11984,N_11120,N_11080);
or U11985 (N_11985,N_11366,N_11294);
or U11986 (N_11986,N_11210,N_11381);
nor U11987 (N_11987,N_11087,N_11416);
and U11988 (N_11988,N_11327,N_11348);
and U11989 (N_11989,N_11013,N_11334);
or U11990 (N_11990,N_11110,N_11382);
or U11991 (N_11991,N_11163,N_11352);
nor U11992 (N_11992,N_11380,N_11456);
or U11993 (N_11993,N_11097,N_11111);
or U11994 (N_11994,N_11068,N_11202);
nand U11995 (N_11995,N_11211,N_11295);
and U11996 (N_11996,N_11105,N_11347);
nand U11997 (N_11997,N_11304,N_11455);
and U11998 (N_11998,N_11135,N_11157);
or U11999 (N_11999,N_11368,N_11144);
or U12000 (N_12000,N_11817,N_11930);
and U12001 (N_12001,N_11613,N_11949);
and U12002 (N_12002,N_11976,N_11687);
or U12003 (N_12003,N_11628,N_11725);
nand U12004 (N_12004,N_11850,N_11945);
xnor U12005 (N_12005,N_11540,N_11656);
nor U12006 (N_12006,N_11999,N_11708);
nand U12007 (N_12007,N_11788,N_11853);
or U12008 (N_12008,N_11884,N_11589);
nand U12009 (N_12009,N_11948,N_11849);
or U12010 (N_12010,N_11966,N_11610);
and U12011 (N_12011,N_11916,N_11583);
or U12012 (N_12012,N_11691,N_11739);
nor U12013 (N_12013,N_11991,N_11764);
nor U12014 (N_12014,N_11501,N_11649);
nor U12015 (N_12015,N_11676,N_11517);
nand U12016 (N_12016,N_11506,N_11942);
or U12017 (N_12017,N_11634,N_11967);
or U12018 (N_12018,N_11908,N_11975);
nor U12019 (N_12019,N_11572,N_11742);
nor U12020 (N_12020,N_11507,N_11671);
or U12021 (N_12021,N_11757,N_11547);
nand U12022 (N_12022,N_11789,N_11630);
or U12023 (N_12023,N_11543,N_11515);
nor U12024 (N_12024,N_11877,N_11792);
and U12025 (N_12025,N_11796,N_11524);
and U12026 (N_12026,N_11844,N_11898);
nor U12027 (N_12027,N_11805,N_11683);
nor U12028 (N_12028,N_11845,N_11903);
and U12029 (N_12029,N_11637,N_11670);
nand U12030 (N_12030,N_11565,N_11837);
or U12031 (N_12031,N_11654,N_11762);
or U12032 (N_12032,N_11773,N_11765);
nor U12033 (N_12033,N_11582,N_11960);
and U12034 (N_12034,N_11887,N_11592);
nand U12035 (N_12035,N_11816,N_11994);
nand U12036 (N_12036,N_11801,N_11738);
and U12037 (N_12037,N_11617,N_11910);
nor U12038 (N_12038,N_11591,N_11595);
nor U12039 (N_12039,N_11866,N_11744);
nor U12040 (N_12040,N_11748,N_11705);
or U12041 (N_12041,N_11558,N_11797);
nand U12042 (N_12042,N_11891,N_11888);
or U12043 (N_12043,N_11746,N_11855);
nand U12044 (N_12044,N_11938,N_11596);
nor U12045 (N_12045,N_11892,N_11560);
nor U12046 (N_12046,N_11751,N_11710);
or U12047 (N_12047,N_11927,N_11714);
or U12048 (N_12048,N_11585,N_11526);
or U12049 (N_12049,N_11950,N_11562);
and U12050 (N_12050,N_11568,N_11566);
or U12051 (N_12051,N_11874,N_11689);
nand U12052 (N_12052,N_11749,N_11939);
and U12053 (N_12053,N_11747,N_11814);
and U12054 (N_12054,N_11545,N_11509);
nor U12055 (N_12055,N_11889,N_11707);
and U12056 (N_12056,N_11775,N_11620);
and U12057 (N_12057,N_11902,N_11922);
and U12058 (N_12058,N_11546,N_11754);
nand U12059 (N_12059,N_11542,N_11651);
nand U12060 (N_12060,N_11755,N_11859);
nand U12061 (N_12061,N_11586,N_11752);
nand U12062 (N_12062,N_11815,N_11590);
nor U12063 (N_12063,N_11989,N_11614);
xor U12064 (N_12064,N_11988,N_11522);
nand U12065 (N_12065,N_11606,N_11777);
nor U12066 (N_12066,N_11909,N_11786);
nor U12067 (N_12067,N_11694,N_11635);
nand U12068 (N_12068,N_11735,N_11642);
or U12069 (N_12069,N_11803,N_11520);
nor U12070 (N_12070,N_11525,N_11569);
nor U12071 (N_12071,N_11799,N_11693);
nor U12072 (N_12072,N_11829,N_11530);
or U12073 (N_12073,N_11821,N_11669);
or U12074 (N_12074,N_11605,N_11963);
nand U12075 (N_12075,N_11657,N_11624);
nor U12076 (N_12076,N_11798,N_11718);
and U12077 (N_12077,N_11984,N_11518);
and U12078 (N_12078,N_11808,N_11852);
nand U12079 (N_12079,N_11774,N_11760);
and U12080 (N_12080,N_11643,N_11502);
or U12081 (N_12081,N_11848,N_11954);
or U12082 (N_12082,N_11871,N_11740);
or U12083 (N_12083,N_11512,N_11882);
or U12084 (N_12084,N_11548,N_11987);
nand U12085 (N_12085,N_11629,N_11559);
xnor U12086 (N_12086,N_11841,N_11990);
and U12087 (N_12087,N_11860,N_11609);
nor U12088 (N_12088,N_11593,N_11872);
nand U12089 (N_12089,N_11573,N_11958);
and U12090 (N_12090,N_11771,N_11625);
nor U12091 (N_12091,N_11701,N_11696);
and U12092 (N_12092,N_11897,N_11679);
or U12093 (N_12093,N_11835,N_11787);
nand U12094 (N_12094,N_11791,N_11597);
and U12095 (N_12095,N_11535,N_11552);
or U12096 (N_12096,N_11985,N_11648);
nor U12097 (N_12097,N_11794,N_11682);
or U12098 (N_12098,N_11615,N_11660);
nand U12099 (N_12099,N_11719,N_11951);
and U12100 (N_12100,N_11536,N_11932);
and U12101 (N_12101,N_11946,N_11686);
xnor U12102 (N_12102,N_11825,N_11864);
nand U12103 (N_12103,N_11832,N_11539);
nand U12104 (N_12104,N_11564,N_11971);
and U12105 (N_12105,N_11551,N_11905);
nor U12106 (N_12106,N_11956,N_11544);
and U12107 (N_12107,N_11918,N_11639);
nand U12108 (N_12108,N_11587,N_11827);
and U12109 (N_12109,N_11528,N_11661);
or U12110 (N_12110,N_11576,N_11875);
or U12111 (N_12111,N_11955,N_11684);
nor U12112 (N_12112,N_11914,N_11830);
nor U12113 (N_12113,N_11846,N_11965);
or U12114 (N_12114,N_11869,N_11741);
or U12115 (N_12115,N_11726,N_11695);
and U12116 (N_12116,N_11729,N_11745);
and U12117 (N_12117,N_11953,N_11778);
nand U12118 (N_12118,N_11861,N_11769);
nor U12119 (N_12119,N_11813,N_11868);
nand U12120 (N_12120,N_11961,N_11776);
nor U12121 (N_12121,N_11603,N_11608);
or U12122 (N_12122,N_11828,N_11503);
nor U12123 (N_12123,N_11921,N_11867);
and U12124 (N_12124,N_11998,N_11857);
or U12125 (N_12125,N_11979,N_11833);
and U12126 (N_12126,N_11940,N_11863);
nand U12127 (N_12127,N_11824,N_11978);
nor U12128 (N_12128,N_11681,N_11982);
nand U12129 (N_12129,N_11728,N_11598);
and U12130 (N_12130,N_11934,N_11619);
nand U12131 (N_12131,N_11578,N_11736);
or U12132 (N_12132,N_11655,N_11793);
nor U12133 (N_12133,N_11785,N_11980);
and U12134 (N_12134,N_11928,N_11699);
nor U12135 (N_12135,N_11756,N_11510);
or U12136 (N_12136,N_11663,N_11981);
or U12137 (N_12137,N_11668,N_11915);
or U12138 (N_12138,N_11843,N_11581);
nor U12139 (N_12139,N_11553,N_11790);
or U12140 (N_12140,N_11621,N_11783);
or U12141 (N_12141,N_11917,N_11622);
nand U12142 (N_12142,N_11865,N_11862);
and U12143 (N_12143,N_11674,N_11957);
or U12144 (N_12144,N_11632,N_11645);
nand U12145 (N_12145,N_11733,N_11926);
or U12146 (N_12146,N_11895,N_11724);
nand U12147 (N_12147,N_11839,N_11952);
nor U12148 (N_12148,N_11537,N_11716);
or U12149 (N_12149,N_11924,N_11662);
nor U12150 (N_12150,N_11667,N_11672);
or U12151 (N_12151,N_11594,N_11720);
or U12152 (N_12152,N_11907,N_11549);
nand U12153 (N_12153,N_11680,N_11819);
and U12154 (N_12154,N_11723,N_11604);
xor U12155 (N_12155,N_11623,N_11513);
and U12156 (N_12156,N_11870,N_11713);
or U12157 (N_12157,N_11931,N_11880);
xor U12158 (N_12158,N_11504,N_11678);
and U12159 (N_12159,N_11636,N_11626);
nand U12160 (N_12160,N_11904,N_11890);
nand U12161 (N_12161,N_11750,N_11781);
nand U12162 (N_12162,N_11554,N_11533);
and U12163 (N_12163,N_11986,N_11532);
and U12164 (N_12164,N_11732,N_11563);
or U12165 (N_12165,N_11944,N_11556);
nand U12166 (N_12166,N_11858,N_11800);
or U12167 (N_12167,N_11700,N_11806);
nand U12168 (N_12168,N_11767,N_11936);
or U12169 (N_12169,N_11659,N_11579);
nand U12170 (N_12170,N_11712,N_11727);
nor U12171 (N_12171,N_11584,N_11650);
nor U12172 (N_12172,N_11500,N_11838);
xnor U12173 (N_12173,N_11962,N_11709);
and U12174 (N_12174,N_11664,N_11570);
and U12175 (N_12175,N_11514,N_11531);
nand U12176 (N_12176,N_11899,N_11935);
nand U12177 (N_12177,N_11658,N_11571);
or U12178 (N_12178,N_11826,N_11995);
nor U12179 (N_12179,N_11809,N_11652);
nand U12180 (N_12180,N_11703,N_11780);
and U12181 (N_12181,N_11779,N_11666);
or U12182 (N_12182,N_11929,N_11900);
nor U12183 (N_12183,N_11600,N_11618);
and U12184 (N_12184,N_11947,N_11722);
nand U12185 (N_12185,N_11685,N_11675);
and U12186 (N_12186,N_11879,N_11627);
or U12187 (N_12187,N_11697,N_11937);
nor U12188 (N_12188,N_11529,N_11577);
and U12189 (N_12189,N_11519,N_11784);
nor U12190 (N_12190,N_11943,N_11856);
nor U12191 (N_12191,N_11920,N_11973);
nor U12192 (N_12192,N_11969,N_11766);
xor U12193 (N_12193,N_11541,N_11840);
or U12194 (N_12194,N_11612,N_11919);
nor U12195 (N_12195,N_11823,N_11883);
and U12196 (N_12196,N_11818,N_11616);
or U12197 (N_12197,N_11893,N_11761);
nand U12198 (N_12198,N_11802,N_11561);
nand U12199 (N_12199,N_11873,N_11601);
nand U12200 (N_12200,N_11959,N_11731);
and U12201 (N_12201,N_11804,N_11550);
and U12202 (N_12202,N_11511,N_11811);
or U12203 (N_12203,N_11768,N_11925);
nor U12204 (N_12204,N_11996,N_11702);
nand U12205 (N_12205,N_11646,N_11836);
or U12206 (N_12206,N_11633,N_11631);
or U12207 (N_12207,N_11647,N_11574);
nand U12208 (N_12208,N_11782,N_11923);
nand U12209 (N_12209,N_11698,N_11812);
nor U12210 (N_12210,N_11894,N_11810);
xnor U12211 (N_12211,N_11567,N_11557);
or U12212 (N_12212,N_11820,N_11602);
or U12213 (N_12213,N_11822,N_11993);
nor U12214 (N_12214,N_11977,N_11854);
and U12215 (N_12215,N_11737,N_11770);
nand U12216 (N_12216,N_11521,N_11527);
and U12217 (N_12217,N_11906,N_11665);
or U12218 (N_12218,N_11607,N_11831);
nor U12219 (N_12219,N_11638,N_11640);
and U12220 (N_12220,N_11878,N_11653);
nor U12221 (N_12221,N_11641,N_11972);
nor U12222 (N_12222,N_11516,N_11588);
nand U12223 (N_12223,N_11968,N_11688);
xnor U12224 (N_12224,N_11992,N_11711);
or U12225 (N_12225,N_11912,N_11847);
nor U12226 (N_12226,N_11795,N_11734);
nand U12227 (N_12227,N_11580,N_11523);
nand U12228 (N_12228,N_11772,N_11886);
or U12229 (N_12229,N_11970,N_11913);
or U12230 (N_12230,N_11538,N_11851);
or U12231 (N_12231,N_11941,N_11964);
or U12232 (N_12232,N_11885,N_11730);
and U12233 (N_12233,N_11911,N_11717);
or U12234 (N_12234,N_11673,N_11555);
nand U12235 (N_12235,N_11834,N_11706);
and U12236 (N_12236,N_11508,N_11997);
nor U12237 (N_12237,N_11575,N_11715);
or U12238 (N_12238,N_11896,N_11611);
nor U12239 (N_12239,N_11974,N_11759);
nor U12240 (N_12240,N_11758,N_11599);
or U12241 (N_12241,N_11763,N_11690);
and U12242 (N_12242,N_11876,N_11807);
nand U12243 (N_12243,N_11704,N_11842);
nand U12244 (N_12244,N_11743,N_11933);
and U12245 (N_12245,N_11753,N_11721);
nand U12246 (N_12246,N_11901,N_11505);
nor U12247 (N_12247,N_11644,N_11881);
nor U12248 (N_12248,N_11534,N_11983);
and U12249 (N_12249,N_11677,N_11692);
xnor U12250 (N_12250,N_11706,N_11943);
and U12251 (N_12251,N_11833,N_11956);
nand U12252 (N_12252,N_11992,N_11681);
nor U12253 (N_12253,N_11554,N_11633);
nor U12254 (N_12254,N_11823,N_11843);
nand U12255 (N_12255,N_11738,N_11927);
nor U12256 (N_12256,N_11644,N_11638);
and U12257 (N_12257,N_11800,N_11686);
and U12258 (N_12258,N_11816,N_11503);
and U12259 (N_12259,N_11939,N_11785);
nand U12260 (N_12260,N_11877,N_11546);
and U12261 (N_12261,N_11707,N_11579);
and U12262 (N_12262,N_11715,N_11591);
or U12263 (N_12263,N_11525,N_11762);
and U12264 (N_12264,N_11890,N_11966);
and U12265 (N_12265,N_11943,N_11765);
or U12266 (N_12266,N_11678,N_11783);
or U12267 (N_12267,N_11631,N_11990);
nor U12268 (N_12268,N_11583,N_11646);
or U12269 (N_12269,N_11918,N_11969);
and U12270 (N_12270,N_11859,N_11714);
nand U12271 (N_12271,N_11729,N_11670);
and U12272 (N_12272,N_11664,N_11735);
nor U12273 (N_12273,N_11702,N_11870);
and U12274 (N_12274,N_11929,N_11735);
and U12275 (N_12275,N_11662,N_11676);
and U12276 (N_12276,N_11511,N_11614);
nor U12277 (N_12277,N_11737,N_11560);
and U12278 (N_12278,N_11769,N_11587);
and U12279 (N_12279,N_11693,N_11696);
or U12280 (N_12280,N_11812,N_11866);
or U12281 (N_12281,N_11608,N_11841);
nand U12282 (N_12282,N_11548,N_11869);
nand U12283 (N_12283,N_11637,N_11924);
nand U12284 (N_12284,N_11840,N_11692);
nor U12285 (N_12285,N_11715,N_11922);
nand U12286 (N_12286,N_11959,N_11597);
nor U12287 (N_12287,N_11932,N_11513);
or U12288 (N_12288,N_11888,N_11989);
and U12289 (N_12289,N_11528,N_11943);
nor U12290 (N_12290,N_11984,N_11752);
nand U12291 (N_12291,N_11633,N_11897);
nor U12292 (N_12292,N_11989,N_11532);
and U12293 (N_12293,N_11701,N_11600);
or U12294 (N_12294,N_11532,N_11898);
nor U12295 (N_12295,N_11913,N_11978);
and U12296 (N_12296,N_11692,N_11809);
nor U12297 (N_12297,N_11952,N_11942);
or U12298 (N_12298,N_11850,N_11527);
and U12299 (N_12299,N_11993,N_11899);
nor U12300 (N_12300,N_11824,N_11986);
nand U12301 (N_12301,N_11558,N_11886);
xor U12302 (N_12302,N_11911,N_11764);
nand U12303 (N_12303,N_11572,N_11870);
or U12304 (N_12304,N_11516,N_11594);
nand U12305 (N_12305,N_11518,N_11555);
and U12306 (N_12306,N_11563,N_11753);
and U12307 (N_12307,N_11833,N_11547);
nand U12308 (N_12308,N_11738,N_11890);
or U12309 (N_12309,N_11951,N_11928);
xnor U12310 (N_12310,N_11587,N_11584);
and U12311 (N_12311,N_11782,N_11810);
nor U12312 (N_12312,N_11551,N_11776);
nor U12313 (N_12313,N_11713,N_11985);
nand U12314 (N_12314,N_11909,N_11990);
nor U12315 (N_12315,N_11712,N_11956);
nand U12316 (N_12316,N_11677,N_11857);
nor U12317 (N_12317,N_11512,N_11861);
nand U12318 (N_12318,N_11748,N_11729);
and U12319 (N_12319,N_11865,N_11718);
nand U12320 (N_12320,N_11681,N_11608);
nand U12321 (N_12321,N_11888,N_11955);
nor U12322 (N_12322,N_11798,N_11566);
and U12323 (N_12323,N_11947,N_11793);
or U12324 (N_12324,N_11695,N_11798);
nor U12325 (N_12325,N_11874,N_11815);
nand U12326 (N_12326,N_11850,N_11641);
or U12327 (N_12327,N_11745,N_11759);
and U12328 (N_12328,N_11609,N_11735);
and U12329 (N_12329,N_11652,N_11946);
nand U12330 (N_12330,N_11937,N_11651);
nor U12331 (N_12331,N_11873,N_11665);
nand U12332 (N_12332,N_11563,N_11871);
and U12333 (N_12333,N_11727,N_11759);
and U12334 (N_12334,N_11673,N_11667);
nand U12335 (N_12335,N_11946,N_11829);
nor U12336 (N_12336,N_11542,N_11525);
nor U12337 (N_12337,N_11931,N_11687);
or U12338 (N_12338,N_11712,N_11945);
or U12339 (N_12339,N_11949,N_11595);
or U12340 (N_12340,N_11997,N_11679);
nand U12341 (N_12341,N_11979,N_11622);
and U12342 (N_12342,N_11998,N_11785);
nor U12343 (N_12343,N_11562,N_11641);
or U12344 (N_12344,N_11657,N_11965);
nand U12345 (N_12345,N_11929,N_11992);
nand U12346 (N_12346,N_11564,N_11648);
or U12347 (N_12347,N_11592,N_11566);
and U12348 (N_12348,N_11988,N_11947);
nand U12349 (N_12349,N_11561,N_11770);
nor U12350 (N_12350,N_11633,N_11548);
or U12351 (N_12351,N_11815,N_11779);
or U12352 (N_12352,N_11514,N_11723);
nor U12353 (N_12353,N_11667,N_11873);
nor U12354 (N_12354,N_11982,N_11773);
or U12355 (N_12355,N_11746,N_11989);
nand U12356 (N_12356,N_11774,N_11786);
nand U12357 (N_12357,N_11862,N_11720);
nand U12358 (N_12358,N_11560,N_11943);
nor U12359 (N_12359,N_11699,N_11677);
nand U12360 (N_12360,N_11965,N_11645);
and U12361 (N_12361,N_11848,N_11811);
nor U12362 (N_12362,N_11882,N_11916);
nor U12363 (N_12363,N_11797,N_11687);
nor U12364 (N_12364,N_11655,N_11857);
and U12365 (N_12365,N_11568,N_11774);
or U12366 (N_12366,N_11974,N_11545);
and U12367 (N_12367,N_11555,N_11785);
or U12368 (N_12368,N_11912,N_11715);
or U12369 (N_12369,N_11845,N_11503);
nor U12370 (N_12370,N_11691,N_11936);
or U12371 (N_12371,N_11544,N_11507);
nand U12372 (N_12372,N_11606,N_11610);
and U12373 (N_12373,N_11505,N_11700);
and U12374 (N_12374,N_11689,N_11685);
nor U12375 (N_12375,N_11869,N_11803);
and U12376 (N_12376,N_11656,N_11776);
nand U12377 (N_12377,N_11677,N_11536);
nor U12378 (N_12378,N_11793,N_11533);
or U12379 (N_12379,N_11976,N_11754);
or U12380 (N_12380,N_11531,N_11861);
or U12381 (N_12381,N_11736,N_11768);
nor U12382 (N_12382,N_11560,N_11918);
and U12383 (N_12383,N_11764,N_11829);
nor U12384 (N_12384,N_11677,N_11621);
nor U12385 (N_12385,N_11981,N_11820);
nor U12386 (N_12386,N_11539,N_11777);
and U12387 (N_12387,N_11934,N_11944);
nor U12388 (N_12388,N_11838,N_11860);
or U12389 (N_12389,N_11825,N_11955);
nor U12390 (N_12390,N_11797,N_11802);
or U12391 (N_12391,N_11761,N_11632);
nor U12392 (N_12392,N_11575,N_11889);
or U12393 (N_12393,N_11665,N_11742);
nand U12394 (N_12394,N_11831,N_11937);
and U12395 (N_12395,N_11849,N_11901);
nor U12396 (N_12396,N_11987,N_11544);
and U12397 (N_12397,N_11502,N_11825);
nand U12398 (N_12398,N_11795,N_11923);
or U12399 (N_12399,N_11614,N_11508);
nand U12400 (N_12400,N_11623,N_11778);
nand U12401 (N_12401,N_11885,N_11579);
or U12402 (N_12402,N_11988,N_11787);
and U12403 (N_12403,N_11878,N_11860);
or U12404 (N_12404,N_11888,N_11806);
nand U12405 (N_12405,N_11512,N_11581);
and U12406 (N_12406,N_11859,N_11851);
and U12407 (N_12407,N_11757,N_11770);
or U12408 (N_12408,N_11981,N_11848);
and U12409 (N_12409,N_11807,N_11562);
xor U12410 (N_12410,N_11972,N_11967);
or U12411 (N_12411,N_11781,N_11770);
or U12412 (N_12412,N_11500,N_11794);
or U12413 (N_12413,N_11661,N_11824);
or U12414 (N_12414,N_11689,N_11832);
or U12415 (N_12415,N_11802,N_11695);
nand U12416 (N_12416,N_11753,N_11889);
and U12417 (N_12417,N_11859,N_11637);
or U12418 (N_12418,N_11898,N_11820);
and U12419 (N_12419,N_11549,N_11887);
or U12420 (N_12420,N_11764,N_11522);
nor U12421 (N_12421,N_11764,N_11682);
nor U12422 (N_12422,N_11819,N_11681);
or U12423 (N_12423,N_11705,N_11951);
or U12424 (N_12424,N_11877,N_11517);
nor U12425 (N_12425,N_11763,N_11950);
nand U12426 (N_12426,N_11850,N_11786);
nand U12427 (N_12427,N_11994,N_11723);
or U12428 (N_12428,N_11544,N_11678);
nor U12429 (N_12429,N_11930,N_11966);
and U12430 (N_12430,N_11559,N_11582);
and U12431 (N_12431,N_11526,N_11642);
nand U12432 (N_12432,N_11816,N_11615);
xor U12433 (N_12433,N_11850,N_11615);
nand U12434 (N_12434,N_11938,N_11662);
or U12435 (N_12435,N_11598,N_11994);
nand U12436 (N_12436,N_11954,N_11917);
nor U12437 (N_12437,N_11507,N_11873);
nor U12438 (N_12438,N_11939,N_11853);
nor U12439 (N_12439,N_11766,N_11702);
and U12440 (N_12440,N_11950,N_11597);
or U12441 (N_12441,N_11532,N_11862);
and U12442 (N_12442,N_11852,N_11594);
nor U12443 (N_12443,N_11755,N_11599);
nor U12444 (N_12444,N_11569,N_11584);
and U12445 (N_12445,N_11799,N_11663);
nand U12446 (N_12446,N_11843,N_11671);
and U12447 (N_12447,N_11735,N_11996);
or U12448 (N_12448,N_11521,N_11955);
nand U12449 (N_12449,N_11649,N_11891);
and U12450 (N_12450,N_11857,N_11587);
nand U12451 (N_12451,N_11796,N_11570);
or U12452 (N_12452,N_11702,N_11713);
nand U12453 (N_12453,N_11660,N_11913);
nand U12454 (N_12454,N_11973,N_11617);
nor U12455 (N_12455,N_11901,N_11779);
or U12456 (N_12456,N_11761,N_11780);
or U12457 (N_12457,N_11934,N_11741);
and U12458 (N_12458,N_11889,N_11537);
nand U12459 (N_12459,N_11954,N_11541);
nor U12460 (N_12460,N_11863,N_11992);
and U12461 (N_12461,N_11764,N_11509);
or U12462 (N_12462,N_11978,N_11770);
and U12463 (N_12463,N_11610,N_11571);
and U12464 (N_12464,N_11797,N_11703);
and U12465 (N_12465,N_11776,N_11815);
and U12466 (N_12466,N_11981,N_11588);
nor U12467 (N_12467,N_11751,N_11623);
and U12468 (N_12468,N_11533,N_11596);
nor U12469 (N_12469,N_11575,N_11779);
and U12470 (N_12470,N_11590,N_11825);
nor U12471 (N_12471,N_11800,N_11691);
nand U12472 (N_12472,N_11699,N_11762);
nand U12473 (N_12473,N_11758,N_11591);
or U12474 (N_12474,N_11663,N_11590);
nor U12475 (N_12475,N_11988,N_11922);
nand U12476 (N_12476,N_11975,N_11939);
nand U12477 (N_12477,N_11762,N_11808);
or U12478 (N_12478,N_11624,N_11605);
and U12479 (N_12479,N_11546,N_11934);
nand U12480 (N_12480,N_11976,N_11674);
nand U12481 (N_12481,N_11804,N_11803);
and U12482 (N_12482,N_11724,N_11685);
nand U12483 (N_12483,N_11783,N_11874);
nor U12484 (N_12484,N_11661,N_11529);
nand U12485 (N_12485,N_11574,N_11679);
or U12486 (N_12486,N_11857,N_11816);
nand U12487 (N_12487,N_11555,N_11533);
nor U12488 (N_12488,N_11641,N_11901);
nand U12489 (N_12489,N_11751,N_11862);
and U12490 (N_12490,N_11744,N_11660);
nor U12491 (N_12491,N_11527,N_11896);
nand U12492 (N_12492,N_11553,N_11513);
or U12493 (N_12493,N_11841,N_11785);
and U12494 (N_12494,N_11821,N_11591);
nor U12495 (N_12495,N_11523,N_11818);
and U12496 (N_12496,N_11515,N_11622);
nor U12497 (N_12497,N_11521,N_11755);
or U12498 (N_12498,N_11923,N_11798);
nor U12499 (N_12499,N_11935,N_11883);
or U12500 (N_12500,N_12272,N_12154);
nand U12501 (N_12501,N_12381,N_12443);
nand U12502 (N_12502,N_12486,N_12495);
or U12503 (N_12503,N_12025,N_12431);
nor U12504 (N_12504,N_12153,N_12198);
nand U12505 (N_12505,N_12117,N_12467);
xnor U12506 (N_12506,N_12440,N_12020);
and U12507 (N_12507,N_12307,N_12365);
nand U12508 (N_12508,N_12261,N_12089);
and U12509 (N_12509,N_12048,N_12230);
or U12510 (N_12510,N_12418,N_12062);
and U12511 (N_12511,N_12296,N_12489);
and U12512 (N_12512,N_12090,N_12411);
nand U12513 (N_12513,N_12094,N_12445);
and U12514 (N_12514,N_12339,N_12394);
or U12515 (N_12515,N_12400,N_12469);
and U12516 (N_12516,N_12192,N_12060);
and U12517 (N_12517,N_12099,N_12268);
nor U12518 (N_12518,N_12386,N_12485);
nor U12519 (N_12519,N_12208,N_12321);
nor U12520 (N_12520,N_12404,N_12237);
nand U12521 (N_12521,N_12005,N_12465);
or U12522 (N_12522,N_12328,N_12408);
and U12523 (N_12523,N_12317,N_12419);
xnor U12524 (N_12524,N_12430,N_12122);
or U12525 (N_12525,N_12481,N_12401);
nor U12526 (N_12526,N_12361,N_12068);
nand U12527 (N_12527,N_12113,N_12206);
and U12528 (N_12528,N_12392,N_12450);
or U12529 (N_12529,N_12039,N_12422);
or U12530 (N_12530,N_12405,N_12340);
nand U12531 (N_12531,N_12045,N_12463);
nor U12532 (N_12532,N_12058,N_12146);
xor U12533 (N_12533,N_12003,N_12133);
or U12534 (N_12534,N_12499,N_12442);
nand U12535 (N_12535,N_12051,N_12216);
nand U12536 (N_12536,N_12454,N_12246);
nand U12537 (N_12537,N_12102,N_12239);
and U12538 (N_12538,N_12140,N_12397);
nor U12539 (N_12539,N_12007,N_12281);
and U12540 (N_12540,N_12047,N_12364);
nor U12541 (N_12541,N_12081,N_12278);
and U12542 (N_12542,N_12209,N_12118);
or U12543 (N_12543,N_12366,N_12053);
nor U12544 (N_12544,N_12085,N_12238);
nand U12545 (N_12545,N_12114,N_12242);
xnor U12546 (N_12546,N_12232,N_12357);
or U12547 (N_12547,N_12087,N_12257);
or U12548 (N_12548,N_12160,N_12464);
and U12549 (N_12549,N_12233,N_12001);
or U12550 (N_12550,N_12120,N_12217);
or U12551 (N_12551,N_12398,N_12327);
nand U12552 (N_12552,N_12303,N_12016);
xor U12553 (N_12553,N_12011,N_12482);
nor U12554 (N_12554,N_12144,N_12338);
or U12555 (N_12555,N_12346,N_12282);
nor U12556 (N_12556,N_12182,N_12207);
nor U12557 (N_12557,N_12258,N_12323);
or U12558 (N_12558,N_12121,N_12457);
nand U12559 (N_12559,N_12247,N_12292);
nor U12560 (N_12560,N_12287,N_12377);
and U12561 (N_12561,N_12075,N_12002);
and U12562 (N_12562,N_12289,N_12336);
or U12563 (N_12563,N_12096,N_12195);
nand U12564 (N_12564,N_12064,N_12213);
and U12565 (N_12565,N_12362,N_12265);
or U12566 (N_12566,N_12460,N_12395);
or U12567 (N_12567,N_12479,N_12201);
nor U12568 (N_12568,N_12355,N_12474);
and U12569 (N_12569,N_12125,N_12290);
or U12570 (N_12570,N_12131,N_12251);
nand U12571 (N_12571,N_12214,N_12260);
or U12572 (N_12572,N_12342,N_12147);
and U12573 (N_12573,N_12167,N_12384);
or U12574 (N_12574,N_12176,N_12368);
xnor U12575 (N_12575,N_12017,N_12145);
or U12576 (N_12576,N_12471,N_12014);
nor U12577 (N_12577,N_12097,N_12177);
nor U12578 (N_12578,N_12286,N_12351);
and U12579 (N_12579,N_12028,N_12337);
and U12580 (N_12580,N_12032,N_12390);
and U12581 (N_12581,N_12441,N_12234);
nand U12582 (N_12582,N_12226,N_12139);
nand U12583 (N_12583,N_12447,N_12250);
nand U12584 (N_12584,N_12124,N_12403);
and U12585 (N_12585,N_12370,N_12313);
nand U12586 (N_12586,N_12197,N_12104);
nand U12587 (N_12587,N_12106,N_12136);
and U12588 (N_12588,N_12449,N_12150);
or U12589 (N_12589,N_12222,N_12379);
or U12590 (N_12590,N_12107,N_12249);
nand U12591 (N_12591,N_12253,N_12335);
or U12592 (N_12592,N_12036,N_12175);
nor U12593 (N_12593,N_12241,N_12204);
and U12594 (N_12594,N_12166,N_12484);
or U12595 (N_12595,N_12185,N_12179);
nand U12596 (N_12596,N_12428,N_12000);
and U12597 (N_12597,N_12318,N_12172);
and U12598 (N_12598,N_12314,N_12149);
nand U12599 (N_12599,N_12389,N_12297);
or U12600 (N_12600,N_12043,N_12284);
or U12601 (N_12601,N_12425,N_12376);
nor U12602 (N_12602,N_12240,N_12426);
nand U12603 (N_12603,N_12203,N_12162);
nand U12604 (N_12604,N_12347,N_12356);
nor U12605 (N_12605,N_12191,N_12302);
or U12606 (N_12606,N_12061,N_12385);
nand U12607 (N_12607,N_12415,N_12212);
xnor U12608 (N_12608,N_12410,N_12046);
and U12609 (N_12609,N_12012,N_12300);
nor U12610 (N_12610,N_12076,N_12088);
or U12611 (N_12611,N_12072,N_12071);
nand U12612 (N_12612,N_12274,N_12128);
nand U12613 (N_12613,N_12433,N_12034);
nor U12614 (N_12614,N_12372,N_12013);
nor U12615 (N_12615,N_12049,N_12159);
or U12616 (N_12616,N_12151,N_12438);
nor U12617 (N_12617,N_12252,N_12388);
and U12618 (N_12618,N_12082,N_12171);
and U12619 (N_12619,N_12473,N_12205);
and U12620 (N_12620,N_12331,N_12414);
xnor U12621 (N_12621,N_12359,N_12084);
nor U12622 (N_12622,N_12135,N_12353);
nor U12623 (N_12623,N_12446,N_12164);
nand U12624 (N_12624,N_12295,N_12273);
and U12625 (N_12625,N_12026,N_12320);
or U12626 (N_12626,N_12210,N_12468);
nor U12627 (N_12627,N_12306,N_12037);
nor U12628 (N_12628,N_12283,N_12218);
or U12629 (N_12629,N_12006,N_12236);
or U12630 (N_12630,N_12453,N_12050);
nand U12631 (N_12631,N_12275,N_12267);
and U12632 (N_12632,N_12288,N_12009);
or U12633 (N_12633,N_12285,N_12312);
or U12634 (N_12634,N_12475,N_12180);
and U12635 (N_12635,N_12349,N_12190);
nand U12636 (N_12636,N_12183,N_12341);
nor U12637 (N_12637,N_12493,N_12200);
and U12638 (N_12638,N_12077,N_12225);
nor U12639 (N_12639,N_12030,N_12137);
or U12640 (N_12640,N_12054,N_12245);
and U12641 (N_12641,N_12399,N_12086);
and U12642 (N_12642,N_12008,N_12031);
nor U12643 (N_12643,N_12483,N_12276);
nand U12644 (N_12644,N_12148,N_12427);
and U12645 (N_12645,N_12256,N_12324);
or U12646 (N_12646,N_12116,N_12193);
nor U12647 (N_12647,N_12004,N_12315);
nand U12648 (N_12648,N_12266,N_12138);
nand U12649 (N_12649,N_12027,N_12134);
nand U12650 (N_12650,N_12413,N_12262);
or U12651 (N_12651,N_12477,N_12199);
and U12652 (N_12652,N_12322,N_12263);
or U12653 (N_12653,N_12022,N_12057);
or U12654 (N_12654,N_12174,N_12316);
nor U12655 (N_12655,N_12196,N_12420);
or U12656 (N_12656,N_12458,N_12396);
nor U12657 (N_12657,N_12310,N_12163);
and U12658 (N_12658,N_12480,N_12123);
and U12659 (N_12659,N_12059,N_12040);
nand U12660 (N_12660,N_12109,N_12070);
nor U12661 (N_12661,N_12434,N_12126);
nand U12662 (N_12662,N_12055,N_12065);
xor U12663 (N_12663,N_12079,N_12024);
nor U12664 (N_12664,N_12211,N_12156);
nor U12665 (N_12665,N_12492,N_12462);
nor U12666 (N_12666,N_12091,N_12093);
or U12667 (N_12667,N_12033,N_12228);
nand U12668 (N_12668,N_12439,N_12170);
nand U12669 (N_12669,N_12215,N_12035);
or U12670 (N_12670,N_12360,N_12452);
and U12671 (N_12671,N_12301,N_12044);
nor U12672 (N_12672,N_12298,N_12299);
or U12673 (N_12673,N_12019,N_12023);
or U12674 (N_12674,N_12456,N_12455);
nand U12675 (N_12675,N_12132,N_12038);
and U12676 (N_12676,N_12248,N_12374);
nand U12677 (N_12677,N_12141,N_12496);
nor U12678 (N_12678,N_12178,N_12305);
and U12679 (N_12679,N_12119,N_12169);
and U12680 (N_12680,N_12373,N_12291);
and U12681 (N_12681,N_12461,N_12383);
nor U12682 (N_12682,N_12319,N_12115);
and U12683 (N_12683,N_12378,N_12103);
nor U12684 (N_12684,N_12476,N_12459);
and U12685 (N_12685,N_12010,N_12437);
or U12686 (N_12686,N_12421,N_12412);
nor U12687 (N_12687,N_12158,N_12490);
nor U12688 (N_12688,N_12333,N_12189);
nor U12689 (N_12689,N_12095,N_12498);
nand U12690 (N_12690,N_12041,N_12407);
nor U12691 (N_12691,N_12435,N_12098);
and U12692 (N_12692,N_12371,N_12108);
or U12693 (N_12693,N_12063,N_12345);
and U12694 (N_12694,N_12387,N_12105);
nor U12695 (N_12695,N_12352,N_12083);
or U12696 (N_12696,N_12402,N_12129);
nand U12697 (N_12697,N_12270,N_12161);
or U12698 (N_12698,N_12491,N_12066);
nor U12699 (N_12699,N_12309,N_12423);
nor U12700 (N_12700,N_12255,N_12326);
nand U12701 (N_12701,N_12254,N_12015);
or U12702 (N_12702,N_12332,N_12073);
or U12703 (N_12703,N_12354,N_12194);
nand U12704 (N_12704,N_12494,N_12101);
or U12705 (N_12705,N_12111,N_12184);
and U12706 (N_12706,N_12311,N_12466);
or U12707 (N_12707,N_12181,N_12021);
nor U12708 (N_12708,N_12369,N_12220);
nand U12709 (N_12709,N_12069,N_12173);
and U12710 (N_12710,N_12269,N_12152);
and U12711 (N_12711,N_12100,N_12470);
and U12712 (N_12712,N_12451,N_12074);
and U12713 (N_12713,N_12358,N_12110);
or U12714 (N_12714,N_12367,N_12280);
nor U12715 (N_12715,N_12127,N_12293);
xor U12716 (N_12716,N_12334,N_12130);
and U12717 (N_12717,N_12056,N_12157);
nor U12718 (N_12718,N_12329,N_12279);
nor U12719 (N_12719,N_12330,N_12078);
nand U12720 (N_12720,N_12488,N_12229);
nor U12721 (N_12721,N_12363,N_12243);
or U12722 (N_12722,N_12406,N_12052);
and U12723 (N_12723,N_12187,N_12429);
or U12724 (N_12724,N_12231,N_12472);
nand U12725 (N_12725,N_12325,N_12497);
nand U12726 (N_12726,N_12417,N_12080);
and U12727 (N_12727,N_12344,N_12067);
nand U12728 (N_12728,N_12350,N_12432);
and U12729 (N_12729,N_12223,N_12142);
and U12730 (N_12730,N_12294,N_12478);
nand U12731 (N_12731,N_12343,N_12487);
xnor U12732 (N_12732,N_12380,N_12304);
xor U12733 (N_12733,N_12277,N_12029);
or U12734 (N_12734,N_12221,N_12018);
nor U12735 (N_12735,N_12348,N_12202);
and U12736 (N_12736,N_12219,N_12244);
nand U12737 (N_12737,N_12424,N_12375);
or U12738 (N_12738,N_12448,N_12042);
nand U12739 (N_12739,N_12168,N_12264);
xor U12740 (N_12740,N_12259,N_12155);
nand U12741 (N_12741,N_12186,N_12227);
and U12742 (N_12742,N_12235,N_12112);
nand U12743 (N_12743,N_12165,N_12143);
nor U12744 (N_12744,N_12271,N_12409);
nand U12745 (N_12745,N_12308,N_12391);
and U12746 (N_12746,N_12382,N_12436);
nor U12747 (N_12747,N_12444,N_12416);
and U12748 (N_12748,N_12188,N_12224);
nor U12749 (N_12749,N_12393,N_12092);
or U12750 (N_12750,N_12189,N_12427);
nand U12751 (N_12751,N_12407,N_12487);
xor U12752 (N_12752,N_12007,N_12474);
and U12753 (N_12753,N_12064,N_12425);
and U12754 (N_12754,N_12451,N_12106);
or U12755 (N_12755,N_12228,N_12472);
nand U12756 (N_12756,N_12396,N_12024);
and U12757 (N_12757,N_12250,N_12323);
nand U12758 (N_12758,N_12016,N_12362);
and U12759 (N_12759,N_12032,N_12189);
and U12760 (N_12760,N_12492,N_12126);
or U12761 (N_12761,N_12488,N_12336);
nor U12762 (N_12762,N_12485,N_12210);
nand U12763 (N_12763,N_12279,N_12154);
nor U12764 (N_12764,N_12337,N_12133);
nand U12765 (N_12765,N_12258,N_12488);
and U12766 (N_12766,N_12041,N_12299);
nand U12767 (N_12767,N_12075,N_12194);
nand U12768 (N_12768,N_12405,N_12469);
nand U12769 (N_12769,N_12308,N_12052);
and U12770 (N_12770,N_12495,N_12470);
nor U12771 (N_12771,N_12459,N_12170);
and U12772 (N_12772,N_12286,N_12419);
nor U12773 (N_12773,N_12483,N_12028);
nor U12774 (N_12774,N_12246,N_12107);
nand U12775 (N_12775,N_12465,N_12073);
nor U12776 (N_12776,N_12482,N_12165);
nor U12777 (N_12777,N_12225,N_12288);
and U12778 (N_12778,N_12084,N_12138);
xor U12779 (N_12779,N_12463,N_12111);
or U12780 (N_12780,N_12412,N_12232);
and U12781 (N_12781,N_12344,N_12096);
or U12782 (N_12782,N_12230,N_12249);
and U12783 (N_12783,N_12289,N_12003);
or U12784 (N_12784,N_12057,N_12040);
and U12785 (N_12785,N_12007,N_12095);
nor U12786 (N_12786,N_12042,N_12437);
nand U12787 (N_12787,N_12066,N_12302);
and U12788 (N_12788,N_12259,N_12186);
nand U12789 (N_12789,N_12456,N_12142);
xor U12790 (N_12790,N_12418,N_12101);
nor U12791 (N_12791,N_12260,N_12342);
or U12792 (N_12792,N_12144,N_12016);
and U12793 (N_12793,N_12273,N_12455);
or U12794 (N_12794,N_12053,N_12376);
nand U12795 (N_12795,N_12212,N_12454);
nand U12796 (N_12796,N_12207,N_12086);
nand U12797 (N_12797,N_12440,N_12047);
nand U12798 (N_12798,N_12407,N_12079);
nand U12799 (N_12799,N_12216,N_12416);
nand U12800 (N_12800,N_12222,N_12463);
nor U12801 (N_12801,N_12481,N_12477);
nor U12802 (N_12802,N_12262,N_12088);
nand U12803 (N_12803,N_12362,N_12004);
nand U12804 (N_12804,N_12224,N_12405);
or U12805 (N_12805,N_12481,N_12154);
nand U12806 (N_12806,N_12457,N_12294);
nor U12807 (N_12807,N_12375,N_12216);
nand U12808 (N_12808,N_12326,N_12025);
or U12809 (N_12809,N_12193,N_12181);
or U12810 (N_12810,N_12084,N_12303);
nand U12811 (N_12811,N_12259,N_12316);
nor U12812 (N_12812,N_12141,N_12222);
and U12813 (N_12813,N_12335,N_12491);
and U12814 (N_12814,N_12347,N_12137);
nand U12815 (N_12815,N_12047,N_12025);
or U12816 (N_12816,N_12166,N_12103);
nor U12817 (N_12817,N_12101,N_12455);
nand U12818 (N_12818,N_12002,N_12266);
nor U12819 (N_12819,N_12470,N_12197);
nand U12820 (N_12820,N_12106,N_12006);
nor U12821 (N_12821,N_12161,N_12104);
and U12822 (N_12822,N_12164,N_12053);
nor U12823 (N_12823,N_12107,N_12157);
nand U12824 (N_12824,N_12147,N_12008);
or U12825 (N_12825,N_12165,N_12357);
nor U12826 (N_12826,N_12445,N_12037);
nor U12827 (N_12827,N_12200,N_12416);
nor U12828 (N_12828,N_12434,N_12116);
or U12829 (N_12829,N_12209,N_12438);
and U12830 (N_12830,N_12477,N_12349);
nor U12831 (N_12831,N_12095,N_12188);
nor U12832 (N_12832,N_12212,N_12479);
and U12833 (N_12833,N_12096,N_12016);
or U12834 (N_12834,N_12189,N_12450);
nor U12835 (N_12835,N_12291,N_12446);
or U12836 (N_12836,N_12213,N_12342);
nand U12837 (N_12837,N_12165,N_12449);
or U12838 (N_12838,N_12010,N_12327);
or U12839 (N_12839,N_12164,N_12317);
and U12840 (N_12840,N_12088,N_12273);
nor U12841 (N_12841,N_12116,N_12015);
nor U12842 (N_12842,N_12351,N_12301);
xor U12843 (N_12843,N_12496,N_12225);
or U12844 (N_12844,N_12116,N_12198);
and U12845 (N_12845,N_12034,N_12444);
and U12846 (N_12846,N_12171,N_12326);
and U12847 (N_12847,N_12329,N_12266);
nand U12848 (N_12848,N_12065,N_12425);
nor U12849 (N_12849,N_12296,N_12268);
nand U12850 (N_12850,N_12349,N_12479);
nor U12851 (N_12851,N_12035,N_12417);
nor U12852 (N_12852,N_12343,N_12403);
xnor U12853 (N_12853,N_12119,N_12483);
or U12854 (N_12854,N_12398,N_12229);
or U12855 (N_12855,N_12102,N_12117);
nor U12856 (N_12856,N_12451,N_12264);
nand U12857 (N_12857,N_12169,N_12030);
or U12858 (N_12858,N_12358,N_12398);
nand U12859 (N_12859,N_12076,N_12414);
and U12860 (N_12860,N_12053,N_12049);
nor U12861 (N_12861,N_12159,N_12190);
or U12862 (N_12862,N_12371,N_12101);
nor U12863 (N_12863,N_12013,N_12323);
or U12864 (N_12864,N_12433,N_12074);
nand U12865 (N_12865,N_12323,N_12114);
nand U12866 (N_12866,N_12097,N_12447);
and U12867 (N_12867,N_12306,N_12036);
nand U12868 (N_12868,N_12149,N_12394);
nor U12869 (N_12869,N_12397,N_12087);
nand U12870 (N_12870,N_12113,N_12441);
nor U12871 (N_12871,N_12443,N_12023);
nor U12872 (N_12872,N_12158,N_12232);
nand U12873 (N_12873,N_12329,N_12104);
or U12874 (N_12874,N_12485,N_12135);
and U12875 (N_12875,N_12164,N_12402);
nor U12876 (N_12876,N_12083,N_12364);
and U12877 (N_12877,N_12366,N_12497);
nor U12878 (N_12878,N_12283,N_12036);
nand U12879 (N_12879,N_12279,N_12082);
nand U12880 (N_12880,N_12374,N_12122);
nor U12881 (N_12881,N_12046,N_12290);
or U12882 (N_12882,N_12379,N_12391);
or U12883 (N_12883,N_12396,N_12191);
or U12884 (N_12884,N_12020,N_12146);
and U12885 (N_12885,N_12477,N_12402);
nand U12886 (N_12886,N_12077,N_12364);
nand U12887 (N_12887,N_12363,N_12460);
nor U12888 (N_12888,N_12404,N_12215);
nand U12889 (N_12889,N_12345,N_12210);
or U12890 (N_12890,N_12336,N_12394);
nand U12891 (N_12891,N_12110,N_12160);
nor U12892 (N_12892,N_12262,N_12352);
nor U12893 (N_12893,N_12092,N_12083);
and U12894 (N_12894,N_12180,N_12339);
nand U12895 (N_12895,N_12289,N_12460);
nand U12896 (N_12896,N_12025,N_12280);
or U12897 (N_12897,N_12437,N_12363);
xnor U12898 (N_12898,N_12222,N_12147);
nor U12899 (N_12899,N_12058,N_12007);
nand U12900 (N_12900,N_12361,N_12431);
nor U12901 (N_12901,N_12315,N_12066);
and U12902 (N_12902,N_12235,N_12106);
and U12903 (N_12903,N_12117,N_12336);
or U12904 (N_12904,N_12337,N_12079);
nor U12905 (N_12905,N_12299,N_12117);
nor U12906 (N_12906,N_12198,N_12233);
nor U12907 (N_12907,N_12238,N_12168);
nor U12908 (N_12908,N_12188,N_12176);
nor U12909 (N_12909,N_12367,N_12238);
and U12910 (N_12910,N_12206,N_12387);
and U12911 (N_12911,N_12136,N_12151);
nor U12912 (N_12912,N_12015,N_12324);
or U12913 (N_12913,N_12166,N_12235);
or U12914 (N_12914,N_12188,N_12498);
nor U12915 (N_12915,N_12473,N_12176);
or U12916 (N_12916,N_12291,N_12077);
and U12917 (N_12917,N_12090,N_12418);
nor U12918 (N_12918,N_12087,N_12207);
or U12919 (N_12919,N_12011,N_12213);
nand U12920 (N_12920,N_12208,N_12035);
nand U12921 (N_12921,N_12047,N_12299);
or U12922 (N_12922,N_12329,N_12458);
xor U12923 (N_12923,N_12274,N_12436);
nor U12924 (N_12924,N_12307,N_12187);
nor U12925 (N_12925,N_12344,N_12281);
nor U12926 (N_12926,N_12375,N_12364);
or U12927 (N_12927,N_12098,N_12071);
nand U12928 (N_12928,N_12259,N_12042);
or U12929 (N_12929,N_12467,N_12248);
and U12930 (N_12930,N_12265,N_12214);
or U12931 (N_12931,N_12048,N_12008);
or U12932 (N_12932,N_12421,N_12346);
nand U12933 (N_12933,N_12145,N_12295);
or U12934 (N_12934,N_12272,N_12009);
xor U12935 (N_12935,N_12069,N_12368);
or U12936 (N_12936,N_12177,N_12448);
and U12937 (N_12937,N_12379,N_12182);
and U12938 (N_12938,N_12256,N_12249);
nand U12939 (N_12939,N_12264,N_12038);
or U12940 (N_12940,N_12186,N_12485);
or U12941 (N_12941,N_12295,N_12323);
and U12942 (N_12942,N_12326,N_12201);
and U12943 (N_12943,N_12451,N_12483);
nand U12944 (N_12944,N_12228,N_12218);
nand U12945 (N_12945,N_12229,N_12091);
nand U12946 (N_12946,N_12060,N_12387);
nor U12947 (N_12947,N_12088,N_12103);
and U12948 (N_12948,N_12305,N_12187);
and U12949 (N_12949,N_12125,N_12311);
nor U12950 (N_12950,N_12399,N_12029);
and U12951 (N_12951,N_12181,N_12145);
or U12952 (N_12952,N_12412,N_12229);
nand U12953 (N_12953,N_12405,N_12382);
nand U12954 (N_12954,N_12000,N_12107);
or U12955 (N_12955,N_12015,N_12420);
or U12956 (N_12956,N_12449,N_12348);
nand U12957 (N_12957,N_12215,N_12255);
nor U12958 (N_12958,N_12103,N_12343);
nor U12959 (N_12959,N_12393,N_12000);
xor U12960 (N_12960,N_12300,N_12124);
nor U12961 (N_12961,N_12014,N_12165);
and U12962 (N_12962,N_12068,N_12120);
and U12963 (N_12963,N_12041,N_12282);
and U12964 (N_12964,N_12459,N_12343);
nand U12965 (N_12965,N_12166,N_12205);
and U12966 (N_12966,N_12384,N_12190);
nor U12967 (N_12967,N_12483,N_12190);
or U12968 (N_12968,N_12394,N_12052);
xor U12969 (N_12969,N_12414,N_12086);
or U12970 (N_12970,N_12317,N_12274);
and U12971 (N_12971,N_12459,N_12257);
nand U12972 (N_12972,N_12255,N_12252);
or U12973 (N_12973,N_12306,N_12066);
nand U12974 (N_12974,N_12345,N_12467);
or U12975 (N_12975,N_12024,N_12255);
and U12976 (N_12976,N_12280,N_12213);
or U12977 (N_12977,N_12474,N_12025);
nor U12978 (N_12978,N_12193,N_12481);
and U12979 (N_12979,N_12364,N_12314);
nor U12980 (N_12980,N_12019,N_12480);
and U12981 (N_12981,N_12007,N_12268);
and U12982 (N_12982,N_12374,N_12322);
nand U12983 (N_12983,N_12078,N_12120);
and U12984 (N_12984,N_12299,N_12434);
nor U12985 (N_12985,N_12076,N_12359);
nand U12986 (N_12986,N_12341,N_12297);
and U12987 (N_12987,N_12051,N_12401);
or U12988 (N_12988,N_12279,N_12141);
nand U12989 (N_12989,N_12048,N_12356);
nand U12990 (N_12990,N_12186,N_12376);
nor U12991 (N_12991,N_12264,N_12233);
and U12992 (N_12992,N_12262,N_12417);
or U12993 (N_12993,N_12309,N_12364);
nor U12994 (N_12994,N_12172,N_12203);
nor U12995 (N_12995,N_12092,N_12455);
nand U12996 (N_12996,N_12091,N_12470);
and U12997 (N_12997,N_12277,N_12300);
and U12998 (N_12998,N_12222,N_12172);
nand U12999 (N_12999,N_12376,N_12359);
nor U13000 (N_13000,N_12562,N_12929);
xnor U13001 (N_13001,N_12776,N_12937);
nand U13002 (N_13002,N_12629,N_12561);
nand U13003 (N_13003,N_12762,N_12731);
or U13004 (N_13004,N_12799,N_12963);
and U13005 (N_13005,N_12950,N_12990);
and U13006 (N_13006,N_12861,N_12645);
nand U13007 (N_13007,N_12701,N_12864);
or U13008 (N_13008,N_12570,N_12623);
or U13009 (N_13009,N_12761,N_12828);
or U13010 (N_13010,N_12932,N_12572);
nor U13011 (N_13011,N_12696,N_12555);
or U13012 (N_13012,N_12594,N_12979);
or U13013 (N_13013,N_12604,N_12906);
nand U13014 (N_13014,N_12569,N_12903);
or U13015 (N_13015,N_12796,N_12521);
xor U13016 (N_13016,N_12620,N_12916);
xnor U13017 (N_13017,N_12954,N_12636);
nand U13018 (N_13018,N_12786,N_12563);
nor U13019 (N_13019,N_12969,N_12850);
nor U13020 (N_13020,N_12613,N_12726);
or U13021 (N_13021,N_12592,N_12751);
nand U13022 (N_13022,N_12525,N_12920);
and U13023 (N_13023,N_12879,N_12797);
and U13024 (N_13024,N_12893,N_12805);
or U13025 (N_13025,N_12809,N_12512);
or U13026 (N_13026,N_12885,N_12977);
or U13027 (N_13027,N_12652,N_12812);
nand U13028 (N_13028,N_12576,N_12754);
xor U13029 (N_13029,N_12635,N_12985);
nor U13030 (N_13030,N_12948,N_12806);
or U13031 (N_13031,N_12826,N_12608);
nor U13032 (N_13032,N_12825,N_12559);
nor U13033 (N_13033,N_12778,N_12574);
nand U13034 (N_13034,N_12624,N_12681);
and U13035 (N_13035,N_12891,N_12831);
nor U13036 (N_13036,N_12853,N_12838);
or U13037 (N_13037,N_12863,N_12504);
and U13038 (N_13038,N_12527,N_12852);
and U13039 (N_13039,N_12578,N_12600);
nor U13040 (N_13040,N_12571,N_12999);
nor U13041 (N_13041,N_12974,N_12707);
or U13042 (N_13042,N_12859,N_12738);
or U13043 (N_13043,N_12533,N_12649);
and U13044 (N_13044,N_12709,N_12936);
or U13045 (N_13045,N_12908,N_12529);
and U13046 (N_13046,N_12736,N_12952);
nor U13047 (N_13047,N_12711,N_12914);
or U13048 (N_13048,N_12585,N_12710);
or U13049 (N_13049,N_12595,N_12591);
and U13050 (N_13050,N_12759,N_12794);
nand U13051 (N_13051,N_12811,N_12921);
and U13052 (N_13052,N_12982,N_12993);
nor U13053 (N_13053,N_12820,N_12757);
nor U13054 (N_13054,N_12808,N_12606);
nor U13055 (N_13055,N_12832,N_12933);
nor U13056 (N_13056,N_12669,N_12745);
xnor U13057 (N_13057,N_12617,N_12763);
xor U13058 (N_13058,N_12945,N_12889);
nor U13059 (N_13059,N_12520,N_12780);
and U13060 (N_13060,N_12637,N_12934);
and U13061 (N_13061,N_12741,N_12522);
and U13062 (N_13062,N_12719,N_12654);
nor U13063 (N_13063,N_12566,N_12717);
nand U13064 (N_13064,N_12560,N_12940);
nor U13065 (N_13065,N_12946,N_12735);
nor U13066 (N_13066,N_12573,N_12845);
nor U13067 (N_13067,N_12925,N_12777);
or U13068 (N_13068,N_12800,N_12765);
or U13069 (N_13069,N_12750,N_12854);
or U13070 (N_13070,N_12856,N_12550);
nor U13071 (N_13071,N_12840,N_12848);
nand U13072 (N_13072,N_12650,N_12989);
and U13073 (N_13073,N_12674,N_12515);
nand U13074 (N_13074,N_12638,N_12737);
and U13075 (N_13075,N_12643,N_12807);
nand U13076 (N_13076,N_12683,N_12770);
nor U13077 (N_13077,N_12822,N_12657);
and U13078 (N_13078,N_12723,N_12911);
or U13079 (N_13079,N_12729,N_12835);
nand U13080 (N_13080,N_12813,N_12603);
and U13081 (N_13081,N_12827,N_12746);
or U13082 (N_13082,N_12703,N_12714);
and U13083 (N_13083,N_12919,N_12695);
nand U13084 (N_13084,N_12855,N_12689);
nor U13085 (N_13085,N_12915,N_12802);
nand U13086 (N_13086,N_12791,N_12542);
and U13087 (N_13087,N_12733,N_12615);
and U13088 (N_13088,N_12716,N_12953);
or U13089 (N_13089,N_12679,N_12756);
nand U13090 (N_13090,N_12534,N_12642);
nor U13091 (N_13091,N_12720,N_12888);
nor U13092 (N_13092,N_12740,N_12590);
nor U13093 (N_13093,N_12935,N_12506);
nor U13094 (N_13094,N_12616,N_12607);
xor U13095 (N_13095,N_12941,N_12535);
nor U13096 (N_13096,N_12837,N_12959);
nand U13097 (N_13097,N_12579,N_12818);
and U13098 (N_13098,N_12849,N_12668);
nor U13099 (N_13099,N_12902,N_12787);
nand U13100 (N_13100,N_12869,N_12687);
or U13101 (N_13101,N_12973,N_12829);
or U13102 (N_13102,N_12552,N_12942);
and U13103 (N_13103,N_12532,N_12988);
and U13104 (N_13104,N_12773,N_12632);
nor U13105 (N_13105,N_12898,N_12841);
and U13106 (N_13106,N_12670,N_12510);
and U13107 (N_13107,N_12602,N_12793);
and U13108 (N_13108,N_12847,N_12685);
nor U13109 (N_13109,N_12697,N_12749);
or U13110 (N_13110,N_12732,N_12634);
or U13111 (N_13111,N_12890,N_12927);
or U13112 (N_13112,N_12747,N_12951);
nor U13113 (N_13113,N_12851,N_12580);
or U13114 (N_13114,N_12865,N_12713);
and U13115 (N_13115,N_12795,N_12609);
or U13116 (N_13116,N_12972,N_12782);
nand U13117 (N_13117,N_12955,N_12748);
nor U13118 (N_13118,N_12528,N_12682);
nor U13119 (N_13119,N_12882,N_12753);
xnor U13120 (N_13120,N_12507,N_12577);
nor U13121 (N_13121,N_12768,N_12673);
nor U13122 (N_13122,N_12675,N_12834);
nor U13123 (N_13123,N_12666,N_12862);
or U13124 (N_13124,N_12548,N_12901);
and U13125 (N_13125,N_12596,N_12992);
nand U13126 (N_13126,N_12539,N_12551);
or U13127 (N_13127,N_12910,N_12790);
and U13128 (N_13128,N_12651,N_12949);
or U13129 (N_13129,N_12783,N_12547);
and U13130 (N_13130,N_12785,N_12663);
and U13131 (N_13131,N_12544,N_12692);
nand U13132 (N_13132,N_12870,N_12630);
nand U13133 (N_13133,N_12897,N_12508);
and U13134 (N_13134,N_12715,N_12625);
nand U13135 (N_13135,N_12612,N_12691);
nor U13136 (N_13136,N_12967,N_12830);
and U13137 (N_13137,N_12819,N_12994);
nand U13138 (N_13138,N_12976,N_12775);
nand U13139 (N_13139,N_12917,N_12628);
or U13140 (N_13140,N_12839,N_12621);
or U13141 (N_13141,N_12907,N_12611);
nand U13142 (N_13142,N_12878,N_12699);
xor U13143 (N_13143,N_12743,N_12928);
nor U13144 (N_13144,N_12700,N_12727);
nor U13145 (N_13145,N_12526,N_12693);
nand U13146 (N_13146,N_12918,N_12694);
nor U13147 (N_13147,N_12833,N_12789);
nor U13148 (N_13148,N_12704,N_12997);
nand U13149 (N_13149,N_12788,N_12771);
and U13150 (N_13150,N_12686,N_12958);
or U13151 (N_13151,N_12960,N_12734);
and U13152 (N_13152,N_12905,N_12721);
nand U13153 (N_13153,N_12647,N_12610);
nor U13154 (N_13154,N_12639,N_12947);
and U13155 (N_13155,N_12658,N_12678);
or U13156 (N_13156,N_12671,N_12892);
or U13157 (N_13157,N_12633,N_12540);
or U13158 (N_13158,N_12648,N_12755);
or U13159 (N_13159,N_12883,N_12896);
nand U13160 (N_13160,N_12660,N_12900);
nor U13161 (N_13161,N_12922,N_12659);
nand U13162 (N_13162,N_12913,N_12517);
nand U13163 (N_13163,N_12509,N_12501);
or U13164 (N_13164,N_12981,N_12646);
xnor U13165 (N_13165,N_12655,N_12823);
nand U13166 (N_13166,N_12582,N_12871);
nor U13167 (N_13167,N_12939,N_12866);
nor U13168 (N_13168,N_12868,N_12965);
or U13169 (N_13169,N_12876,N_12505);
and U13170 (N_13170,N_12998,N_12676);
and U13171 (N_13171,N_12764,N_12886);
nand U13172 (N_13172,N_12986,N_12564);
nor U13173 (N_13173,N_12565,N_12618);
or U13174 (N_13174,N_12518,N_12516);
and U13175 (N_13175,N_12567,N_12817);
and U13176 (N_13176,N_12792,N_12556);
nor U13177 (N_13177,N_12500,N_12537);
or U13178 (N_13178,N_12712,N_12698);
nor U13179 (N_13179,N_12545,N_12758);
and U13180 (N_13180,N_12543,N_12597);
and U13181 (N_13181,N_12943,N_12502);
and U13182 (N_13182,N_12656,N_12684);
nand U13183 (N_13183,N_12867,N_12996);
and U13184 (N_13184,N_12593,N_12706);
xnor U13185 (N_13185,N_12575,N_12798);
or U13186 (N_13186,N_12702,N_12641);
nand U13187 (N_13187,N_12843,N_12962);
nand U13188 (N_13188,N_12944,N_12583);
nand U13189 (N_13189,N_12983,N_12991);
nand U13190 (N_13190,N_12664,N_12554);
and U13191 (N_13191,N_12665,N_12752);
xnor U13192 (N_13192,N_12588,N_12690);
nand U13193 (N_13193,N_12586,N_12730);
nor U13194 (N_13194,N_12672,N_12601);
and U13195 (N_13195,N_12987,N_12514);
nand U13196 (N_13196,N_12966,N_12667);
or U13197 (N_13197,N_12557,N_12688);
nor U13198 (N_13198,N_12880,N_12513);
or U13199 (N_13199,N_12899,N_12875);
and U13200 (N_13200,N_12774,N_12558);
and U13201 (N_13201,N_12661,N_12677);
nand U13202 (N_13202,N_12810,N_12769);
and U13203 (N_13203,N_12541,N_12549);
nor U13204 (N_13204,N_12626,N_12779);
nor U13205 (N_13205,N_12857,N_12873);
nor U13206 (N_13206,N_12728,N_12894);
nor U13207 (N_13207,N_12722,N_12538);
nor U13208 (N_13208,N_12824,N_12524);
nand U13209 (N_13209,N_12815,N_12877);
nand U13210 (N_13210,N_12725,N_12530);
or U13211 (N_13211,N_12971,N_12909);
or U13212 (N_13212,N_12961,N_12804);
or U13213 (N_13213,N_12975,N_12846);
nand U13214 (N_13214,N_12904,N_12619);
nand U13215 (N_13215,N_12640,N_12842);
nor U13216 (N_13216,N_12772,N_12803);
nand U13217 (N_13217,N_12860,N_12598);
and U13218 (N_13218,N_12938,N_12984);
or U13219 (N_13219,N_12568,N_12821);
nand U13220 (N_13220,N_12653,N_12964);
and U13221 (N_13221,N_12995,N_12519);
or U13222 (N_13222,N_12887,N_12881);
and U13223 (N_13223,N_12644,N_12605);
and U13224 (N_13224,N_12872,N_12926);
or U13225 (N_13225,N_12784,N_12708);
nor U13226 (N_13226,N_12724,N_12622);
nand U13227 (N_13227,N_12742,N_12718);
nand U13228 (N_13228,N_12924,N_12912);
and U13229 (N_13229,N_12614,N_12662);
or U13230 (N_13230,N_12631,N_12523);
nor U13231 (N_13231,N_12739,N_12980);
or U13232 (N_13232,N_12744,N_12766);
nor U13233 (N_13233,N_12705,N_12531);
or U13234 (N_13234,N_12781,N_12767);
nand U13235 (N_13235,N_12801,N_12923);
nor U13236 (N_13236,N_12581,N_12931);
and U13237 (N_13237,N_12844,N_12930);
nor U13238 (N_13238,N_12956,N_12874);
or U13239 (N_13239,N_12584,N_12836);
nor U13240 (N_13240,N_12536,N_12858);
or U13241 (N_13241,N_12895,N_12760);
nand U13242 (N_13242,N_12814,N_12627);
nand U13243 (N_13243,N_12884,N_12599);
xnor U13244 (N_13244,N_12816,N_12957);
and U13245 (N_13245,N_12680,N_12978);
and U13246 (N_13246,N_12970,N_12546);
or U13247 (N_13247,N_12968,N_12553);
or U13248 (N_13248,N_12589,N_12587);
nor U13249 (N_13249,N_12511,N_12503);
nand U13250 (N_13250,N_12814,N_12698);
nand U13251 (N_13251,N_12678,N_12734);
or U13252 (N_13252,N_12607,N_12997);
nor U13253 (N_13253,N_12994,N_12850);
and U13254 (N_13254,N_12768,N_12565);
and U13255 (N_13255,N_12752,N_12613);
and U13256 (N_13256,N_12650,N_12737);
or U13257 (N_13257,N_12656,N_12519);
or U13258 (N_13258,N_12574,N_12702);
nor U13259 (N_13259,N_12595,N_12691);
nor U13260 (N_13260,N_12934,N_12697);
nand U13261 (N_13261,N_12984,N_12507);
nand U13262 (N_13262,N_12616,N_12565);
nor U13263 (N_13263,N_12799,N_12905);
nor U13264 (N_13264,N_12818,N_12864);
nor U13265 (N_13265,N_12559,N_12566);
and U13266 (N_13266,N_12926,N_12910);
nand U13267 (N_13267,N_12631,N_12992);
and U13268 (N_13268,N_12801,N_12955);
nand U13269 (N_13269,N_12774,N_12661);
nand U13270 (N_13270,N_12503,N_12607);
nor U13271 (N_13271,N_12918,N_12987);
or U13272 (N_13272,N_12843,N_12715);
nor U13273 (N_13273,N_12511,N_12516);
and U13274 (N_13274,N_12878,N_12605);
nand U13275 (N_13275,N_12935,N_12699);
nand U13276 (N_13276,N_12801,N_12757);
and U13277 (N_13277,N_12618,N_12891);
or U13278 (N_13278,N_12649,N_12993);
and U13279 (N_13279,N_12511,N_12755);
xnor U13280 (N_13280,N_12919,N_12614);
and U13281 (N_13281,N_12707,N_12787);
nand U13282 (N_13282,N_12678,N_12919);
nand U13283 (N_13283,N_12522,N_12798);
nand U13284 (N_13284,N_12908,N_12584);
or U13285 (N_13285,N_12934,N_12679);
or U13286 (N_13286,N_12642,N_12660);
or U13287 (N_13287,N_12627,N_12604);
nor U13288 (N_13288,N_12942,N_12544);
or U13289 (N_13289,N_12637,N_12710);
nor U13290 (N_13290,N_12855,N_12995);
or U13291 (N_13291,N_12980,N_12517);
nand U13292 (N_13292,N_12889,N_12878);
nor U13293 (N_13293,N_12556,N_12904);
and U13294 (N_13294,N_12821,N_12656);
nor U13295 (N_13295,N_12544,N_12879);
nor U13296 (N_13296,N_12630,N_12606);
nor U13297 (N_13297,N_12635,N_12871);
nor U13298 (N_13298,N_12511,N_12502);
nor U13299 (N_13299,N_12571,N_12904);
xnor U13300 (N_13300,N_12679,N_12901);
nand U13301 (N_13301,N_12530,N_12999);
nor U13302 (N_13302,N_12951,N_12786);
or U13303 (N_13303,N_12822,N_12925);
and U13304 (N_13304,N_12760,N_12979);
nor U13305 (N_13305,N_12779,N_12735);
nor U13306 (N_13306,N_12687,N_12871);
xnor U13307 (N_13307,N_12502,N_12968);
and U13308 (N_13308,N_12763,N_12598);
and U13309 (N_13309,N_12679,N_12604);
nand U13310 (N_13310,N_12988,N_12848);
and U13311 (N_13311,N_12520,N_12979);
nor U13312 (N_13312,N_12614,N_12834);
nand U13313 (N_13313,N_12783,N_12842);
and U13314 (N_13314,N_12779,N_12792);
nor U13315 (N_13315,N_12813,N_12691);
nand U13316 (N_13316,N_12858,N_12577);
nor U13317 (N_13317,N_12788,N_12765);
nand U13318 (N_13318,N_12636,N_12899);
nand U13319 (N_13319,N_12831,N_12569);
nand U13320 (N_13320,N_12864,N_12516);
and U13321 (N_13321,N_12847,N_12662);
or U13322 (N_13322,N_12765,N_12576);
nor U13323 (N_13323,N_12637,N_12739);
and U13324 (N_13324,N_12677,N_12519);
nand U13325 (N_13325,N_12635,N_12804);
and U13326 (N_13326,N_12586,N_12947);
nor U13327 (N_13327,N_12985,N_12887);
nor U13328 (N_13328,N_12737,N_12532);
or U13329 (N_13329,N_12584,N_12878);
and U13330 (N_13330,N_12776,N_12749);
nor U13331 (N_13331,N_12839,N_12611);
xnor U13332 (N_13332,N_12608,N_12554);
or U13333 (N_13333,N_12833,N_12971);
nor U13334 (N_13334,N_12784,N_12845);
or U13335 (N_13335,N_12783,N_12993);
nand U13336 (N_13336,N_12918,N_12506);
nor U13337 (N_13337,N_12865,N_12841);
nand U13338 (N_13338,N_12831,N_12821);
or U13339 (N_13339,N_12692,N_12695);
or U13340 (N_13340,N_12874,N_12757);
and U13341 (N_13341,N_12876,N_12979);
nand U13342 (N_13342,N_12777,N_12780);
nand U13343 (N_13343,N_12685,N_12898);
nor U13344 (N_13344,N_12803,N_12841);
and U13345 (N_13345,N_12842,N_12672);
nand U13346 (N_13346,N_12983,N_12885);
nor U13347 (N_13347,N_12622,N_12753);
or U13348 (N_13348,N_12961,N_12855);
nor U13349 (N_13349,N_12542,N_12599);
or U13350 (N_13350,N_12900,N_12608);
and U13351 (N_13351,N_12624,N_12502);
and U13352 (N_13352,N_12506,N_12986);
and U13353 (N_13353,N_12843,N_12800);
and U13354 (N_13354,N_12879,N_12883);
nor U13355 (N_13355,N_12766,N_12507);
nor U13356 (N_13356,N_12657,N_12500);
nand U13357 (N_13357,N_12522,N_12500);
nand U13358 (N_13358,N_12589,N_12566);
nor U13359 (N_13359,N_12815,N_12548);
nand U13360 (N_13360,N_12600,N_12937);
nor U13361 (N_13361,N_12843,N_12727);
and U13362 (N_13362,N_12613,N_12994);
nor U13363 (N_13363,N_12676,N_12988);
nor U13364 (N_13364,N_12673,N_12986);
and U13365 (N_13365,N_12736,N_12770);
and U13366 (N_13366,N_12824,N_12567);
or U13367 (N_13367,N_12799,N_12866);
or U13368 (N_13368,N_12727,N_12525);
and U13369 (N_13369,N_12549,N_12724);
nand U13370 (N_13370,N_12619,N_12858);
and U13371 (N_13371,N_12740,N_12748);
xor U13372 (N_13372,N_12796,N_12509);
nand U13373 (N_13373,N_12523,N_12961);
and U13374 (N_13374,N_12970,N_12611);
xnor U13375 (N_13375,N_12656,N_12693);
or U13376 (N_13376,N_12780,N_12819);
and U13377 (N_13377,N_12702,N_12733);
nand U13378 (N_13378,N_12715,N_12604);
nor U13379 (N_13379,N_12905,N_12611);
and U13380 (N_13380,N_12552,N_12882);
and U13381 (N_13381,N_12928,N_12519);
nor U13382 (N_13382,N_12931,N_12545);
and U13383 (N_13383,N_12924,N_12694);
or U13384 (N_13384,N_12673,N_12753);
nand U13385 (N_13385,N_12530,N_12501);
and U13386 (N_13386,N_12588,N_12740);
and U13387 (N_13387,N_12676,N_12928);
or U13388 (N_13388,N_12699,N_12681);
and U13389 (N_13389,N_12888,N_12516);
nor U13390 (N_13390,N_12960,N_12841);
and U13391 (N_13391,N_12825,N_12619);
and U13392 (N_13392,N_12562,N_12661);
and U13393 (N_13393,N_12868,N_12937);
xnor U13394 (N_13394,N_12979,N_12574);
nand U13395 (N_13395,N_12644,N_12529);
or U13396 (N_13396,N_12908,N_12725);
and U13397 (N_13397,N_12822,N_12744);
and U13398 (N_13398,N_12659,N_12522);
nand U13399 (N_13399,N_12956,N_12693);
nand U13400 (N_13400,N_12850,N_12539);
nand U13401 (N_13401,N_12573,N_12593);
nor U13402 (N_13402,N_12647,N_12885);
nor U13403 (N_13403,N_12911,N_12756);
or U13404 (N_13404,N_12899,N_12694);
nor U13405 (N_13405,N_12725,N_12880);
or U13406 (N_13406,N_12747,N_12577);
nor U13407 (N_13407,N_12904,N_12966);
and U13408 (N_13408,N_12727,N_12699);
nor U13409 (N_13409,N_12614,N_12811);
or U13410 (N_13410,N_12661,N_12992);
nand U13411 (N_13411,N_12744,N_12866);
nand U13412 (N_13412,N_12639,N_12764);
and U13413 (N_13413,N_12564,N_12683);
nor U13414 (N_13414,N_12613,N_12688);
nor U13415 (N_13415,N_12539,N_12979);
nor U13416 (N_13416,N_12513,N_12949);
or U13417 (N_13417,N_12834,N_12646);
and U13418 (N_13418,N_12702,N_12667);
and U13419 (N_13419,N_12853,N_12956);
nand U13420 (N_13420,N_12706,N_12995);
nor U13421 (N_13421,N_12756,N_12519);
nor U13422 (N_13422,N_12720,N_12906);
and U13423 (N_13423,N_12789,N_12602);
and U13424 (N_13424,N_12873,N_12983);
nand U13425 (N_13425,N_12534,N_12914);
or U13426 (N_13426,N_12713,N_12980);
or U13427 (N_13427,N_12525,N_12880);
or U13428 (N_13428,N_12612,N_12989);
or U13429 (N_13429,N_12911,N_12628);
nor U13430 (N_13430,N_12932,N_12900);
or U13431 (N_13431,N_12978,N_12522);
nand U13432 (N_13432,N_12907,N_12616);
xnor U13433 (N_13433,N_12747,N_12798);
nand U13434 (N_13434,N_12544,N_12924);
and U13435 (N_13435,N_12861,N_12844);
nand U13436 (N_13436,N_12653,N_12630);
nor U13437 (N_13437,N_12708,N_12871);
or U13438 (N_13438,N_12905,N_12933);
and U13439 (N_13439,N_12870,N_12633);
xor U13440 (N_13440,N_12958,N_12973);
nor U13441 (N_13441,N_12840,N_12639);
and U13442 (N_13442,N_12705,N_12923);
xor U13443 (N_13443,N_12849,N_12635);
and U13444 (N_13444,N_12569,N_12660);
and U13445 (N_13445,N_12896,N_12952);
nand U13446 (N_13446,N_12944,N_12998);
nor U13447 (N_13447,N_12789,N_12794);
nor U13448 (N_13448,N_12592,N_12728);
and U13449 (N_13449,N_12898,N_12699);
or U13450 (N_13450,N_12781,N_12680);
or U13451 (N_13451,N_12626,N_12698);
nor U13452 (N_13452,N_12892,N_12874);
nand U13453 (N_13453,N_12735,N_12665);
or U13454 (N_13454,N_12623,N_12979);
and U13455 (N_13455,N_12695,N_12862);
or U13456 (N_13456,N_12657,N_12928);
or U13457 (N_13457,N_12655,N_12815);
and U13458 (N_13458,N_12650,N_12534);
or U13459 (N_13459,N_12915,N_12748);
or U13460 (N_13460,N_12681,N_12568);
nand U13461 (N_13461,N_12981,N_12596);
or U13462 (N_13462,N_12736,N_12777);
nor U13463 (N_13463,N_12958,N_12730);
or U13464 (N_13464,N_12582,N_12524);
or U13465 (N_13465,N_12754,N_12567);
nor U13466 (N_13466,N_12842,N_12643);
or U13467 (N_13467,N_12935,N_12736);
and U13468 (N_13468,N_12998,N_12788);
nor U13469 (N_13469,N_12515,N_12636);
nand U13470 (N_13470,N_12852,N_12501);
and U13471 (N_13471,N_12763,N_12960);
and U13472 (N_13472,N_12547,N_12773);
nand U13473 (N_13473,N_12929,N_12526);
or U13474 (N_13474,N_12733,N_12889);
nor U13475 (N_13475,N_12598,N_12972);
and U13476 (N_13476,N_12968,N_12910);
nor U13477 (N_13477,N_12709,N_12825);
nor U13478 (N_13478,N_12688,N_12569);
nor U13479 (N_13479,N_12836,N_12880);
nand U13480 (N_13480,N_12864,N_12837);
and U13481 (N_13481,N_12757,N_12569);
or U13482 (N_13482,N_12638,N_12506);
nor U13483 (N_13483,N_12945,N_12999);
and U13484 (N_13484,N_12939,N_12677);
nand U13485 (N_13485,N_12698,N_12612);
nand U13486 (N_13486,N_12840,N_12752);
nor U13487 (N_13487,N_12843,N_12936);
and U13488 (N_13488,N_12749,N_12522);
nor U13489 (N_13489,N_12697,N_12815);
or U13490 (N_13490,N_12747,N_12566);
nor U13491 (N_13491,N_12576,N_12866);
nor U13492 (N_13492,N_12782,N_12850);
nor U13493 (N_13493,N_12978,N_12717);
or U13494 (N_13494,N_12841,N_12555);
or U13495 (N_13495,N_12836,N_12825);
or U13496 (N_13496,N_12807,N_12871);
nand U13497 (N_13497,N_12558,N_12967);
and U13498 (N_13498,N_12894,N_12746);
nand U13499 (N_13499,N_12596,N_12926);
or U13500 (N_13500,N_13244,N_13214);
or U13501 (N_13501,N_13484,N_13075);
or U13502 (N_13502,N_13094,N_13285);
nor U13503 (N_13503,N_13167,N_13002);
or U13504 (N_13504,N_13202,N_13170);
or U13505 (N_13505,N_13052,N_13207);
or U13506 (N_13506,N_13031,N_13462);
nand U13507 (N_13507,N_13158,N_13287);
or U13508 (N_13508,N_13335,N_13100);
and U13509 (N_13509,N_13069,N_13422);
nor U13510 (N_13510,N_13453,N_13276);
or U13511 (N_13511,N_13470,N_13406);
nor U13512 (N_13512,N_13416,N_13062);
nand U13513 (N_13513,N_13138,N_13349);
nand U13514 (N_13514,N_13384,N_13454);
and U13515 (N_13515,N_13277,N_13171);
xor U13516 (N_13516,N_13284,N_13354);
or U13517 (N_13517,N_13457,N_13319);
nor U13518 (N_13518,N_13491,N_13231);
or U13519 (N_13519,N_13212,N_13123);
and U13520 (N_13520,N_13303,N_13118);
and U13521 (N_13521,N_13221,N_13488);
and U13522 (N_13522,N_13217,N_13059);
nand U13523 (N_13523,N_13371,N_13172);
and U13524 (N_13524,N_13005,N_13022);
and U13525 (N_13525,N_13072,N_13429);
and U13526 (N_13526,N_13139,N_13197);
nand U13527 (N_13527,N_13015,N_13314);
nand U13528 (N_13528,N_13196,N_13086);
nor U13529 (N_13529,N_13003,N_13134);
nand U13530 (N_13530,N_13074,N_13001);
or U13531 (N_13531,N_13033,N_13154);
or U13532 (N_13532,N_13157,N_13340);
and U13533 (N_13533,N_13203,N_13364);
nand U13534 (N_13534,N_13498,N_13255);
nand U13535 (N_13535,N_13328,N_13449);
nand U13536 (N_13536,N_13324,N_13159);
nand U13537 (N_13537,N_13288,N_13427);
or U13538 (N_13538,N_13050,N_13205);
and U13539 (N_13539,N_13258,N_13093);
xor U13540 (N_13540,N_13473,N_13497);
nand U13541 (N_13541,N_13073,N_13325);
nand U13542 (N_13542,N_13351,N_13252);
or U13543 (N_13543,N_13249,N_13192);
nand U13544 (N_13544,N_13432,N_13496);
nor U13545 (N_13545,N_13297,N_13299);
nand U13546 (N_13546,N_13327,N_13257);
nor U13547 (N_13547,N_13101,N_13129);
nor U13548 (N_13548,N_13256,N_13004);
nand U13549 (N_13549,N_13108,N_13467);
nor U13550 (N_13550,N_13119,N_13136);
and U13551 (N_13551,N_13346,N_13048);
nand U13552 (N_13552,N_13060,N_13085);
and U13553 (N_13553,N_13260,N_13239);
nor U13554 (N_13554,N_13487,N_13087);
nand U13555 (N_13555,N_13341,N_13020);
nand U13556 (N_13556,N_13238,N_13195);
or U13557 (N_13557,N_13402,N_13440);
or U13558 (N_13558,N_13306,N_13153);
nor U13559 (N_13559,N_13392,N_13263);
or U13560 (N_13560,N_13317,N_13178);
nand U13561 (N_13561,N_13420,N_13266);
or U13562 (N_13562,N_13103,N_13366);
nand U13563 (N_13563,N_13273,N_13436);
and U13564 (N_13564,N_13039,N_13415);
nand U13565 (N_13565,N_13320,N_13289);
or U13566 (N_13566,N_13458,N_13146);
or U13567 (N_13567,N_13193,N_13318);
nor U13568 (N_13568,N_13477,N_13378);
nand U13569 (N_13569,N_13216,N_13127);
or U13570 (N_13570,N_13471,N_13408);
nor U13571 (N_13571,N_13247,N_13077);
nor U13572 (N_13572,N_13067,N_13267);
nand U13573 (N_13573,N_13053,N_13082);
and U13574 (N_13574,N_13381,N_13226);
nor U13575 (N_13575,N_13095,N_13390);
and U13576 (N_13576,N_13499,N_13271);
or U13577 (N_13577,N_13316,N_13301);
or U13578 (N_13578,N_13021,N_13110);
nand U13579 (N_13579,N_13128,N_13208);
nor U13580 (N_13580,N_13389,N_13142);
and U13581 (N_13581,N_13494,N_13469);
nor U13582 (N_13582,N_13163,N_13315);
nor U13583 (N_13583,N_13274,N_13054);
nor U13584 (N_13584,N_13220,N_13042);
nand U13585 (N_13585,N_13492,N_13359);
or U13586 (N_13586,N_13369,N_13357);
nand U13587 (N_13587,N_13362,N_13292);
nor U13588 (N_13588,N_13379,N_13293);
and U13589 (N_13589,N_13233,N_13188);
nor U13590 (N_13590,N_13330,N_13385);
nand U13591 (N_13591,N_13468,N_13122);
and U13592 (N_13592,N_13310,N_13076);
and U13593 (N_13593,N_13291,N_13463);
or U13594 (N_13594,N_13223,N_13311);
or U13595 (N_13595,N_13116,N_13112);
nand U13596 (N_13596,N_13438,N_13140);
and U13597 (N_13597,N_13115,N_13162);
nand U13598 (N_13598,N_13040,N_13456);
nand U13599 (N_13599,N_13344,N_13012);
nand U13600 (N_13600,N_13080,N_13133);
nand U13601 (N_13601,N_13368,N_13485);
and U13602 (N_13602,N_13345,N_13332);
nand U13603 (N_13603,N_13298,N_13281);
nand U13604 (N_13604,N_13236,N_13472);
nand U13605 (N_13605,N_13017,N_13044);
or U13606 (N_13606,N_13437,N_13355);
nand U13607 (N_13607,N_13079,N_13227);
nor U13608 (N_13608,N_13176,N_13296);
or U13609 (N_13609,N_13398,N_13204);
and U13610 (N_13610,N_13387,N_13229);
or U13611 (N_13611,N_13113,N_13377);
nor U13612 (N_13612,N_13024,N_13117);
xnor U13613 (N_13613,N_13006,N_13419);
and U13614 (N_13614,N_13361,N_13265);
or U13615 (N_13615,N_13184,N_13414);
nor U13616 (N_13616,N_13036,N_13027);
or U13617 (N_13617,N_13312,N_13465);
nand U13618 (N_13618,N_13401,N_13160);
nor U13619 (N_13619,N_13211,N_13342);
nor U13620 (N_13620,N_13025,N_13261);
nor U13621 (N_13621,N_13026,N_13206);
and U13622 (N_13622,N_13373,N_13121);
nand U13623 (N_13623,N_13007,N_13089);
nor U13624 (N_13624,N_13348,N_13283);
or U13625 (N_13625,N_13337,N_13386);
or U13626 (N_13626,N_13186,N_13441);
nor U13627 (N_13627,N_13105,N_13466);
or U13628 (N_13628,N_13034,N_13019);
nor U13629 (N_13629,N_13347,N_13264);
nor U13630 (N_13630,N_13008,N_13329);
and U13631 (N_13631,N_13222,N_13032);
or U13632 (N_13632,N_13097,N_13495);
nand U13633 (N_13633,N_13307,N_13225);
nor U13634 (N_13634,N_13442,N_13413);
or U13635 (N_13635,N_13391,N_13464);
nor U13636 (N_13636,N_13251,N_13125);
nor U13637 (N_13637,N_13295,N_13322);
or U13638 (N_13638,N_13434,N_13201);
nand U13639 (N_13639,N_13275,N_13164);
nor U13640 (N_13640,N_13189,N_13180);
nand U13641 (N_13641,N_13124,N_13417);
or U13642 (N_13642,N_13070,N_13200);
nor U13643 (N_13643,N_13057,N_13240);
nor U13644 (N_13644,N_13383,N_13372);
nand U13645 (N_13645,N_13209,N_13043);
nand U13646 (N_13646,N_13111,N_13451);
nor U13647 (N_13647,N_13421,N_13083);
nand U13648 (N_13648,N_13148,N_13305);
and U13649 (N_13649,N_13166,N_13445);
nor U13650 (N_13650,N_13308,N_13068);
or U13651 (N_13651,N_13182,N_13107);
or U13652 (N_13652,N_13165,N_13365);
xor U13653 (N_13653,N_13219,N_13334);
nand U13654 (N_13654,N_13055,N_13278);
and U13655 (N_13655,N_13374,N_13397);
nand U13656 (N_13656,N_13047,N_13137);
and U13657 (N_13657,N_13155,N_13412);
or U13658 (N_13658,N_13000,N_13168);
nor U13659 (N_13659,N_13323,N_13131);
or U13660 (N_13660,N_13143,N_13038);
or U13661 (N_13661,N_13248,N_13407);
nand U13662 (N_13662,N_13404,N_13064);
nor U13663 (N_13663,N_13161,N_13302);
and U13664 (N_13664,N_13078,N_13237);
nor U13665 (N_13665,N_13213,N_13290);
and U13666 (N_13666,N_13423,N_13049);
xor U13667 (N_13667,N_13030,N_13411);
nand U13668 (N_13668,N_13210,N_13280);
nand U13669 (N_13669,N_13246,N_13375);
or U13670 (N_13670,N_13241,N_13056);
nor U13671 (N_13671,N_13191,N_13099);
or U13672 (N_13672,N_13058,N_13370);
xnor U13673 (N_13673,N_13151,N_13224);
or U13674 (N_13674,N_13363,N_13272);
nand U13675 (N_13675,N_13106,N_13424);
and U13676 (N_13676,N_13190,N_13091);
nand U13677 (N_13677,N_13144,N_13018);
nand U13678 (N_13678,N_13230,N_13382);
nand U13679 (N_13679,N_13388,N_13259);
nor U13680 (N_13680,N_13326,N_13313);
and U13681 (N_13681,N_13482,N_13141);
nor U13682 (N_13682,N_13145,N_13051);
xor U13683 (N_13683,N_13336,N_13367);
or U13684 (N_13684,N_13029,N_13393);
nor U13685 (N_13685,N_13218,N_13120);
xnor U13686 (N_13686,N_13490,N_13028);
nand U13687 (N_13687,N_13198,N_13450);
or U13688 (N_13688,N_13061,N_13135);
nand U13689 (N_13689,N_13199,N_13035);
nand U13690 (N_13690,N_13126,N_13480);
nand U13691 (N_13691,N_13268,N_13479);
nand U13692 (N_13692,N_13353,N_13046);
nor U13693 (N_13693,N_13262,N_13460);
nor U13694 (N_13694,N_13183,N_13179);
and U13695 (N_13695,N_13010,N_13399);
nor U13696 (N_13696,N_13333,N_13114);
and U13697 (N_13697,N_13081,N_13147);
and U13698 (N_13698,N_13452,N_13152);
nor U13699 (N_13699,N_13489,N_13169);
xor U13700 (N_13700,N_13483,N_13394);
nor U13701 (N_13701,N_13090,N_13185);
nand U13702 (N_13702,N_13228,N_13352);
nor U13703 (N_13703,N_13254,N_13011);
nor U13704 (N_13704,N_13242,N_13215);
nand U13705 (N_13705,N_13433,N_13279);
nor U13706 (N_13706,N_13459,N_13013);
or U13707 (N_13707,N_13426,N_13016);
and U13708 (N_13708,N_13096,N_13448);
and U13709 (N_13709,N_13177,N_13187);
nor U13710 (N_13710,N_13132,N_13425);
xnor U13711 (N_13711,N_13338,N_13009);
nand U13712 (N_13712,N_13023,N_13234);
nand U13713 (N_13713,N_13173,N_13321);
nor U13714 (N_13714,N_13376,N_13065);
or U13715 (N_13715,N_13109,N_13300);
and U13716 (N_13716,N_13396,N_13294);
nor U13717 (N_13717,N_13245,N_13088);
or U13718 (N_13718,N_13235,N_13475);
and U13719 (N_13719,N_13447,N_13250);
nor U13720 (N_13720,N_13474,N_13418);
nand U13721 (N_13721,N_13098,N_13084);
or U13722 (N_13722,N_13493,N_13356);
and U13723 (N_13723,N_13243,N_13410);
or U13724 (N_13724,N_13149,N_13104);
nor U13725 (N_13725,N_13286,N_13405);
nand U13726 (N_13726,N_13102,N_13150);
or U13727 (N_13727,N_13430,N_13063);
and U13728 (N_13728,N_13269,N_13071);
nor U13729 (N_13729,N_13270,N_13041);
nor U13730 (N_13730,N_13092,N_13309);
and U13731 (N_13731,N_13350,N_13400);
and U13732 (N_13732,N_13486,N_13409);
or U13733 (N_13733,N_13045,N_13443);
nor U13734 (N_13734,N_13282,N_13476);
and U13735 (N_13735,N_13435,N_13194);
xnor U13736 (N_13736,N_13343,N_13478);
nand U13737 (N_13737,N_13439,N_13395);
and U13738 (N_13738,N_13253,N_13175);
nand U13739 (N_13739,N_13431,N_13232);
nor U13740 (N_13740,N_13174,N_13428);
and U13741 (N_13741,N_13066,N_13331);
xor U13742 (N_13742,N_13181,N_13358);
nand U13743 (N_13743,N_13037,N_13339);
or U13744 (N_13744,N_13461,N_13130);
nand U13745 (N_13745,N_13403,N_13014);
and U13746 (N_13746,N_13360,N_13481);
or U13747 (N_13747,N_13380,N_13156);
nand U13748 (N_13748,N_13446,N_13455);
nand U13749 (N_13749,N_13444,N_13304);
nand U13750 (N_13750,N_13379,N_13316);
nor U13751 (N_13751,N_13156,N_13247);
nor U13752 (N_13752,N_13240,N_13445);
nand U13753 (N_13753,N_13242,N_13327);
and U13754 (N_13754,N_13157,N_13332);
and U13755 (N_13755,N_13140,N_13011);
nand U13756 (N_13756,N_13198,N_13346);
nor U13757 (N_13757,N_13277,N_13402);
or U13758 (N_13758,N_13135,N_13447);
nand U13759 (N_13759,N_13243,N_13010);
nand U13760 (N_13760,N_13476,N_13011);
nand U13761 (N_13761,N_13217,N_13345);
nor U13762 (N_13762,N_13328,N_13351);
or U13763 (N_13763,N_13454,N_13330);
nor U13764 (N_13764,N_13289,N_13167);
nand U13765 (N_13765,N_13048,N_13375);
nand U13766 (N_13766,N_13229,N_13035);
nand U13767 (N_13767,N_13390,N_13180);
xor U13768 (N_13768,N_13090,N_13451);
or U13769 (N_13769,N_13048,N_13104);
nand U13770 (N_13770,N_13387,N_13149);
nand U13771 (N_13771,N_13282,N_13276);
nor U13772 (N_13772,N_13238,N_13014);
and U13773 (N_13773,N_13436,N_13367);
and U13774 (N_13774,N_13230,N_13341);
nand U13775 (N_13775,N_13005,N_13076);
nand U13776 (N_13776,N_13464,N_13090);
or U13777 (N_13777,N_13097,N_13489);
and U13778 (N_13778,N_13415,N_13431);
nand U13779 (N_13779,N_13292,N_13279);
or U13780 (N_13780,N_13299,N_13317);
and U13781 (N_13781,N_13140,N_13055);
and U13782 (N_13782,N_13144,N_13272);
nand U13783 (N_13783,N_13492,N_13255);
and U13784 (N_13784,N_13442,N_13099);
nor U13785 (N_13785,N_13400,N_13118);
nor U13786 (N_13786,N_13234,N_13221);
and U13787 (N_13787,N_13178,N_13166);
nand U13788 (N_13788,N_13331,N_13349);
nand U13789 (N_13789,N_13468,N_13301);
nand U13790 (N_13790,N_13154,N_13034);
nand U13791 (N_13791,N_13195,N_13115);
or U13792 (N_13792,N_13193,N_13449);
nor U13793 (N_13793,N_13177,N_13314);
nor U13794 (N_13794,N_13400,N_13454);
nand U13795 (N_13795,N_13494,N_13228);
and U13796 (N_13796,N_13397,N_13054);
or U13797 (N_13797,N_13120,N_13301);
xnor U13798 (N_13798,N_13013,N_13442);
or U13799 (N_13799,N_13304,N_13277);
nand U13800 (N_13800,N_13033,N_13399);
or U13801 (N_13801,N_13407,N_13039);
or U13802 (N_13802,N_13251,N_13456);
nor U13803 (N_13803,N_13047,N_13177);
or U13804 (N_13804,N_13342,N_13465);
or U13805 (N_13805,N_13323,N_13425);
nor U13806 (N_13806,N_13485,N_13087);
and U13807 (N_13807,N_13109,N_13224);
or U13808 (N_13808,N_13090,N_13326);
or U13809 (N_13809,N_13458,N_13103);
xor U13810 (N_13810,N_13133,N_13103);
nor U13811 (N_13811,N_13312,N_13077);
nand U13812 (N_13812,N_13151,N_13118);
or U13813 (N_13813,N_13240,N_13466);
and U13814 (N_13814,N_13055,N_13479);
nand U13815 (N_13815,N_13089,N_13201);
and U13816 (N_13816,N_13437,N_13124);
nand U13817 (N_13817,N_13444,N_13264);
or U13818 (N_13818,N_13053,N_13491);
and U13819 (N_13819,N_13384,N_13399);
and U13820 (N_13820,N_13323,N_13455);
nor U13821 (N_13821,N_13325,N_13479);
nand U13822 (N_13822,N_13384,N_13463);
or U13823 (N_13823,N_13270,N_13056);
and U13824 (N_13824,N_13279,N_13076);
or U13825 (N_13825,N_13326,N_13485);
nand U13826 (N_13826,N_13443,N_13478);
or U13827 (N_13827,N_13408,N_13063);
and U13828 (N_13828,N_13210,N_13403);
nand U13829 (N_13829,N_13136,N_13155);
or U13830 (N_13830,N_13325,N_13458);
or U13831 (N_13831,N_13221,N_13216);
nand U13832 (N_13832,N_13089,N_13457);
nand U13833 (N_13833,N_13363,N_13469);
and U13834 (N_13834,N_13257,N_13399);
nand U13835 (N_13835,N_13472,N_13160);
and U13836 (N_13836,N_13100,N_13449);
and U13837 (N_13837,N_13125,N_13020);
nor U13838 (N_13838,N_13134,N_13169);
and U13839 (N_13839,N_13187,N_13358);
nand U13840 (N_13840,N_13204,N_13293);
nor U13841 (N_13841,N_13023,N_13384);
nand U13842 (N_13842,N_13287,N_13155);
nand U13843 (N_13843,N_13006,N_13061);
nor U13844 (N_13844,N_13283,N_13207);
or U13845 (N_13845,N_13407,N_13073);
and U13846 (N_13846,N_13121,N_13402);
xnor U13847 (N_13847,N_13350,N_13113);
or U13848 (N_13848,N_13282,N_13447);
nor U13849 (N_13849,N_13189,N_13288);
nor U13850 (N_13850,N_13376,N_13445);
xor U13851 (N_13851,N_13101,N_13337);
and U13852 (N_13852,N_13110,N_13218);
and U13853 (N_13853,N_13449,N_13401);
nand U13854 (N_13854,N_13053,N_13213);
nand U13855 (N_13855,N_13272,N_13156);
nor U13856 (N_13856,N_13027,N_13070);
nand U13857 (N_13857,N_13429,N_13430);
nand U13858 (N_13858,N_13466,N_13297);
nor U13859 (N_13859,N_13370,N_13353);
or U13860 (N_13860,N_13249,N_13166);
nor U13861 (N_13861,N_13089,N_13042);
or U13862 (N_13862,N_13132,N_13160);
or U13863 (N_13863,N_13329,N_13471);
xor U13864 (N_13864,N_13072,N_13183);
and U13865 (N_13865,N_13151,N_13006);
xnor U13866 (N_13866,N_13343,N_13120);
or U13867 (N_13867,N_13473,N_13068);
nand U13868 (N_13868,N_13126,N_13205);
and U13869 (N_13869,N_13042,N_13353);
nor U13870 (N_13870,N_13042,N_13202);
or U13871 (N_13871,N_13125,N_13079);
nand U13872 (N_13872,N_13433,N_13449);
nand U13873 (N_13873,N_13028,N_13108);
and U13874 (N_13874,N_13090,N_13490);
nor U13875 (N_13875,N_13302,N_13220);
and U13876 (N_13876,N_13217,N_13236);
or U13877 (N_13877,N_13358,N_13390);
and U13878 (N_13878,N_13038,N_13416);
and U13879 (N_13879,N_13048,N_13252);
and U13880 (N_13880,N_13468,N_13094);
and U13881 (N_13881,N_13407,N_13453);
xor U13882 (N_13882,N_13024,N_13428);
or U13883 (N_13883,N_13083,N_13187);
nand U13884 (N_13884,N_13203,N_13411);
and U13885 (N_13885,N_13321,N_13048);
and U13886 (N_13886,N_13452,N_13080);
nand U13887 (N_13887,N_13242,N_13046);
or U13888 (N_13888,N_13359,N_13386);
or U13889 (N_13889,N_13315,N_13380);
xor U13890 (N_13890,N_13014,N_13336);
nand U13891 (N_13891,N_13428,N_13209);
and U13892 (N_13892,N_13095,N_13250);
nand U13893 (N_13893,N_13015,N_13264);
nand U13894 (N_13894,N_13352,N_13305);
or U13895 (N_13895,N_13194,N_13011);
or U13896 (N_13896,N_13112,N_13167);
nor U13897 (N_13897,N_13376,N_13051);
and U13898 (N_13898,N_13492,N_13213);
nor U13899 (N_13899,N_13469,N_13129);
and U13900 (N_13900,N_13184,N_13231);
or U13901 (N_13901,N_13427,N_13214);
nand U13902 (N_13902,N_13371,N_13492);
and U13903 (N_13903,N_13498,N_13152);
and U13904 (N_13904,N_13400,N_13163);
xnor U13905 (N_13905,N_13210,N_13135);
and U13906 (N_13906,N_13054,N_13431);
nor U13907 (N_13907,N_13349,N_13313);
nor U13908 (N_13908,N_13131,N_13242);
nand U13909 (N_13909,N_13016,N_13443);
and U13910 (N_13910,N_13019,N_13027);
or U13911 (N_13911,N_13358,N_13174);
or U13912 (N_13912,N_13309,N_13454);
or U13913 (N_13913,N_13296,N_13116);
and U13914 (N_13914,N_13259,N_13102);
nor U13915 (N_13915,N_13308,N_13449);
nor U13916 (N_13916,N_13180,N_13335);
nand U13917 (N_13917,N_13444,N_13075);
and U13918 (N_13918,N_13153,N_13023);
or U13919 (N_13919,N_13069,N_13415);
nor U13920 (N_13920,N_13285,N_13249);
and U13921 (N_13921,N_13072,N_13017);
and U13922 (N_13922,N_13348,N_13208);
nand U13923 (N_13923,N_13109,N_13465);
or U13924 (N_13924,N_13097,N_13210);
nand U13925 (N_13925,N_13373,N_13382);
nand U13926 (N_13926,N_13471,N_13005);
nand U13927 (N_13927,N_13390,N_13437);
nand U13928 (N_13928,N_13054,N_13281);
nand U13929 (N_13929,N_13297,N_13493);
or U13930 (N_13930,N_13175,N_13084);
nor U13931 (N_13931,N_13260,N_13094);
nand U13932 (N_13932,N_13223,N_13337);
nand U13933 (N_13933,N_13427,N_13221);
nor U13934 (N_13934,N_13327,N_13207);
or U13935 (N_13935,N_13021,N_13027);
and U13936 (N_13936,N_13335,N_13388);
nand U13937 (N_13937,N_13343,N_13370);
or U13938 (N_13938,N_13494,N_13108);
and U13939 (N_13939,N_13244,N_13175);
xor U13940 (N_13940,N_13050,N_13014);
or U13941 (N_13941,N_13242,N_13043);
or U13942 (N_13942,N_13235,N_13467);
nor U13943 (N_13943,N_13338,N_13060);
nand U13944 (N_13944,N_13435,N_13481);
nand U13945 (N_13945,N_13005,N_13045);
and U13946 (N_13946,N_13211,N_13418);
or U13947 (N_13947,N_13252,N_13123);
nor U13948 (N_13948,N_13120,N_13201);
or U13949 (N_13949,N_13013,N_13237);
and U13950 (N_13950,N_13244,N_13109);
or U13951 (N_13951,N_13267,N_13240);
nand U13952 (N_13952,N_13059,N_13238);
and U13953 (N_13953,N_13138,N_13474);
nor U13954 (N_13954,N_13378,N_13273);
nand U13955 (N_13955,N_13039,N_13362);
xor U13956 (N_13956,N_13182,N_13196);
nor U13957 (N_13957,N_13085,N_13095);
and U13958 (N_13958,N_13161,N_13435);
nand U13959 (N_13959,N_13305,N_13398);
nand U13960 (N_13960,N_13064,N_13385);
nor U13961 (N_13961,N_13059,N_13400);
or U13962 (N_13962,N_13486,N_13118);
nand U13963 (N_13963,N_13042,N_13100);
nand U13964 (N_13964,N_13478,N_13273);
nand U13965 (N_13965,N_13214,N_13300);
nor U13966 (N_13966,N_13056,N_13457);
and U13967 (N_13967,N_13214,N_13091);
nand U13968 (N_13968,N_13368,N_13461);
nand U13969 (N_13969,N_13481,N_13059);
or U13970 (N_13970,N_13026,N_13270);
nand U13971 (N_13971,N_13282,N_13456);
or U13972 (N_13972,N_13009,N_13476);
nor U13973 (N_13973,N_13370,N_13225);
or U13974 (N_13974,N_13391,N_13081);
nand U13975 (N_13975,N_13464,N_13275);
nand U13976 (N_13976,N_13167,N_13411);
or U13977 (N_13977,N_13193,N_13334);
nor U13978 (N_13978,N_13260,N_13227);
nand U13979 (N_13979,N_13317,N_13479);
or U13980 (N_13980,N_13033,N_13283);
nand U13981 (N_13981,N_13173,N_13457);
nor U13982 (N_13982,N_13379,N_13389);
or U13983 (N_13983,N_13470,N_13044);
nand U13984 (N_13984,N_13047,N_13438);
or U13985 (N_13985,N_13228,N_13356);
nand U13986 (N_13986,N_13323,N_13128);
xnor U13987 (N_13987,N_13394,N_13025);
and U13988 (N_13988,N_13390,N_13233);
and U13989 (N_13989,N_13336,N_13129);
nand U13990 (N_13990,N_13292,N_13101);
and U13991 (N_13991,N_13497,N_13396);
nand U13992 (N_13992,N_13090,N_13486);
and U13993 (N_13993,N_13258,N_13170);
and U13994 (N_13994,N_13415,N_13279);
and U13995 (N_13995,N_13080,N_13139);
or U13996 (N_13996,N_13406,N_13036);
or U13997 (N_13997,N_13311,N_13119);
nand U13998 (N_13998,N_13363,N_13425);
and U13999 (N_13999,N_13168,N_13461);
or U14000 (N_14000,N_13682,N_13514);
nand U14001 (N_14001,N_13804,N_13852);
and U14002 (N_14002,N_13912,N_13923);
or U14003 (N_14003,N_13958,N_13547);
or U14004 (N_14004,N_13582,N_13945);
nand U14005 (N_14005,N_13932,N_13810);
nor U14006 (N_14006,N_13877,N_13548);
and U14007 (N_14007,N_13893,N_13839);
nor U14008 (N_14008,N_13806,N_13896);
nor U14009 (N_14009,N_13568,N_13573);
nand U14010 (N_14010,N_13976,N_13751);
or U14011 (N_14011,N_13972,N_13508);
nand U14012 (N_14012,N_13605,N_13812);
nor U14013 (N_14013,N_13661,N_13516);
nand U14014 (N_14014,N_13635,N_13634);
or U14015 (N_14015,N_13591,N_13814);
nor U14016 (N_14016,N_13665,N_13894);
and U14017 (N_14017,N_13915,N_13562);
or U14018 (N_14018,N_13553,N_13895);
nand U14019 (N_14019,N_13968,N_13808);
or U14020 (N_14020,N_13578,N_13986);
nand U14021 (N_14021,N_13965,N_13775);
or U14022 (N_14022,N_13997,N_13747);
nand U14023 (N_14023,N_13966,N_13837);
and U14024 (N_14024,N_13755,N_13580);
or U14025 (N_14025,N_13779,N_13761);
nor U14026 (N_14026,N_13821,N_13974);
and U14027 (N_14027,N_13726,N_13550);
nor U14028 (N_14028,N_13956,N_13969);
nand U14029 (N_14029,N_13543,N_13612);
and U14030 (N_14030,N_13787,N_13936);
nand U14031 (N_14031,N_13544,N_13630);
nor U14032 (N_14032,N_13691,N_13638);
nand U14033 (N_14033,N_13700,N_13595);
nand U14034 (N_14034,N_13650,N_13699);
nand U14035 (N_14035,N_13872,N_13698);
or U14036 (N_14036,N_13921,N_13739);
nor U14037 (N_14037,N_13614,N_13913);
or U14038 (N_14038,N_13811,N_13758);
nand U14039 (N_14039,N_13598,N_13704);
or U14040 (N_14040,N_13827,N_13566);
nand U14041 (N_14041,N_13909,N_13782);
nand U14042 (N_14042,N_13863,N_13599);
xor U14043 (N_14043,N_13799,N_13813);
or U14044 (N_14044,N_13924,N_13937);
or U14045 (N_14045,N_13719,N_13693);
nand U14046 (N_14046,N_13639,N_13750);
or U14047 (N_14047,N_13823,N_13664);
and U14048 (N_14048,N_13979,N_13831);
nand U14049 (N_14049,N_13585,N_13886);
and U14050 (N_14050,N_13994,N_13525);
and U14051 (N_14051,N_13529,N_13535);
and U14052 (N_14052,N_13637,N_13753);
and U14053 (N_14053,N_13767,N_13606);
nor U14054 (N_14054,N_13703,N_13982);
nand U14055 (N_14055,N_13731,N_13795);
or U14056 (N_14056,N_13933,N_13926);
nand U14057 (N_14057,N_13871,N_13939);
nor U14058 (N_14058,N_13970,N_13816);
or U14059 (N_14059,N_13769,N_13803);
and U14060 (N_14060,N_13626,N_13928);
or U14061 (N_14061,N_13555,N_13672);
or U14062 (N_14062,N_13511,N_13674);
nand U14063 (N_14063,N_13618,N_13569);
nor U14064 (N_14064,N_13929,N_13844);
nor U14065 (N_14065,N_13991,N_13961);
and U14066 (N_14066,N_13935,N_13727);
or U14067 (N_14067,N_13917,N_13594);
or U14068 (N_14068,N_13696,N_13631);
or U14069 (N_14069,N_13644,N_13820);
nor U14070 (N_14070,N_13841,N_13518);
nor U14071 (N_14071,N_13981,N_13660);
xnor U14072 (N_14072,N_13579,N_13946);
nor U14073 (N_14073,N_13534,N_13581);
and U14074 (N_14074,N_13680,N_13642);
nor U14075 (N_14075,N_13818,N_13616);
and U14076 (N_14076,N_13504,N_13717);
nand U14077 (N_14077,N_13975,N_13987);
and U14078 (N_14078,N_13780,N_13980);
or U14079 (N_14079,N_13705,N_13744);
nor U14080 (N_14080,N_13558,N_13609);
nand U14081 (N_14081,N_13984,N_13902);
nor U14082 (N_14082,N_13584,N_13603);
and U14083 (N_14083,N_13601,N_13523);
nor U14084 (N_14084,N_13608,N_13819);
and U14085 (N_14085,N_13517,N_13918);
and U14086 (N_14086,N_13802,N_13941);
nor U14087 (N_14087,N_13824,N_13919);
nand U14088 (N_14088,N_13718,N_13985);
and U14089 (N_14089,N_13536,N_13645);
or U14090 (N_14090,N_13791,N_13990);
nand U14091 (N_14091,N_13515,N_13989);
or U14092 (N_14092,N_13654,N_13675);
nor U14093 (N_14093,N_13653,N_13526);
and U14094 (N_14094,N_13537,N_13890);
or U14095 (N_14095,N_13754,N_13860);
nand U14096 (N_14096,N_13792,N_13623);
or U14097 (N_14097,N_13746,N_13914);
and U14098 (N_14098,N_13858,N_13549);
nand U14099 (N_14099,N_13659,N_13565);
nor U14100 (N_14100,N_13859,N_13545);
nor U14101 (N_14101,N_13853,N_13829);
or U14102 (N_14102,N_13764,N_13898);
and U14103 (N_14103,N_13776,N_13686);
nor U14104 (N_14104,N_13993,N_13842);
nor U14105 (N_14105,N_13593,N_13540);
nor U14106 (N_14106,N_13762,N_13855);
and U14107 (N_14107,N_13783,N_13790);
nand U14108 (N_14108,N_13607,N_13587);
nand U14109 (N_14109,N_13907,N_13728);
nor U14110 (N_14110,N_13788,N_13501);
or U14111 (N_14111,N_13633,N_13867);
and U14112 (N_14112,N_13528,N_13538);
nor U14113 (N_14113,N_13882,N_13978);
and U14114 (N_14114,N_13772,N_13571);
or U14115 (N_14115,N_13648,N_13800);
nand U14116 (N_14116,N_13815,N_13621);
nand U14117 (N_14117,N_13873,N_13866);
and U14118 (N_14118,N_13657,N_13955);
nand U14119 (N_14119,N_13570,N_13862);
or U14120 (N_14120,N_13702,N_13556);
nor U14121 (N_14121,N_13797,N_13711);
nand U14122 (N_14122,N_13690,N_13967);
nand U14123 (N_14123,N_13785,N_13574);
or U14124 (N_14124,N_13628,N_13983);
nand U14125 (N_14125,N_13602,N_13760);
nor U14126 (N_14126,N_13520,N_13663);
or U14127 (N_14127,N_13998,N_13927);
and U14128 (N_14128,N_13830,N_13851);
nand U14129 (N_14129,N_13888,N_13940);
and U14130 (N_14130,N_13625,N_13695);
and U14131 (N_14131,N_13743,N_13825);
nor U14132 (N_14132,N_13590,N_13950);
and U14133 (N_14133,N_13706,N_13658);
nor U14134 (N_14134,N_13656,N_13794);
nand U14135 (N_14135,N_13713,N_13600);
nand U14136 (N_14136,N_13733,N_13554);
and U14137 (N_14137,N_13885,N_13883);
nand U14138 (N_14138,N_13916,N_13817);
or U14139 (N_14139,N_13732,N_13577);
and U14140 (N_14140,N_13527,N_13583);
nor U14141 (N_14141,N_13905,N_13901);
nor U14142 (N_14142,N_13938,N_13843);
nand U14143 (N_14143,N_13533,N_13521);
or U14144 (N_14144,N_13532,N_13673);
and U14145 (N_14145,N_13708,N_13736);
nor U14146 (N_14146,N_13530,N_13738);
nor U14147 (N_14147,N_13793,N_13567);
nor U14148 (N_14148,N_13992,N_13509);
and U14149 (N_14149,N_13962,N_13756);
nor U14150 (N_14150,N_13949,N_13519);
or U14151 (N_14151,N_13925,N_13506);
or U14152 (N_14152,N_13689,N_13712);
or U14153 (N_14153,N_13889,N_13845);
or U14154 (N_14154,N_13957,N_13522);
nand U14155 (N_14155,N_13944,N_13765);
and U14156 (N_14156,N_13903,N_13908);
xor U14157 (N_14157,N_13768,N_13922);
and U14158 (N_14158,N_13920,N_13900);
and U14159 (N_14159,N_13838,N_13692);
and U14160 (N_14160,N_13597,N_13617);
nand U14161 (N_14161,N_13715,N_13833);
nand U14162 (N_14162,N_13655,N_13671);
xnor U14163 (N_14163,N_13500,N_13615);
nand U14164 (N_14164,N_13687,N_13724);
and U14165 (N_14165,N_13763,N_13505);
nor U14166 (N_14166,N_13546,N_13561);
and U14167 (N_14167,N_13757,N_13971);
nor U14168 (N_14168,N_13931,N_13835);
nand U14169 (N_14169,N_13773,N_13539);
xor U14170 (N_14170,N_13670,N_13541);
and U14171 (N_14171,N_13951,N_13876);
nand U14172 (N_14172,N_13683,N_13759);
and U14173 (N_14173,N_13619,N_13503);
nand U14174 (N_14174,N_13847,N_13942);
nand U14175 (N_14175,N_13973,N_13934);
nand U14176 (N_14176,N_13778,N_13828);
nand U14177 (N_14177,N_13822,N_13510);
or U14178 (N_14178,N_13575,N_13777);
and U14179 (N_14179,N_13770,N_13807);
and U14180 (N_14180,N_13564,N_13688);
or U14181 (N_14181,N_13875,N_13604);
nand U14182 (N_14182,N_13666,N_13507);
and U14183 (N_14183,N_13846,N_13848);
nand U14184 (N_14184,N_13589,N_13960);
or U14185 (N_14185,N_13781,N_13721);
nand U14186 (N_14186,N_13911,N_13801);
and U14187 (N_14187,N_13906,N_13943);
or U14188 (N_14188,N_13643,N_13869);
nor U14189 (N_14189,N_13742,N_13892);
nand U14190 (N_14190,N_13999,N_13735);
nand U14191 (N_14191,N_13796,N_13857);
nor U14192 (N_14192,N_13722,N_13502);
nand U14193 (N_14193,N_13752,N_13627);
or U14194 (N_14194,N_13662,N_13679);
nor U14195 (N_14195,N_13745,N_13694);
or U14196 (N_14196,N_13865,N_13588);
or U14197 (N_14197,N_13899,N_13647);
and U14198 (N_14198,N_13512,N_13576);
and U14199 (N_14199,N_13551,N_13709);
nand U14200 (N_14200,N_13880,N_13707);
and U14201 (N_14201,N_13884,N_13572);
or U14202 (N_14202,N_13881,N_13749);
and U14203 (N_14203,N_13771,N_13636);
nor U14204 (N_14204,N_13849,N_13878);
nor U14205 (N_14205,N_13861,N_13887);
nor U14206 (N_14206,N_13542,N_13676);
nand U14207 (N_14207,N_13870,N_13952);
or U14208 (N_14208,N_13641,N_13836);
nor U14209 (N_14209,N_13826,N_13684);
nor U14210 (N_14210,N_13667,N_13766);
and U14211 (N_14211,N_13620,N_13629);
nand U14212 (N_14212,N_13954,N_13910);
nor U14213 (N_14213,N_13646,N_13685);
and U14214 (N_14214,N_13798,N_13904);
nand U14215 (N_14215,N_13681,N_13964);
nor U14216 (N_14216,N_13741,N_13834);
or U14217 (N_14217,N_13805,N_13897);
nand U14218 (N_14218,N_13531,N_13963);
nor U14219 (N_14219,N_13716,N_13977);
nand U14220 (N_14220,N_13840,N_13586);
or U14221 (N_14221,N_13557,N_13891);
nand U14222 (N_14222,N_13610,N_13652);
nand U14223 (N_14223,N_13809,N_13559);
and U14224 (N_14224,N_13864,N_13701);
or U14225 (N_14225,N_13774,N_13714);
and U14226 (N_14226,N_13953,N_13611);
and U14227 (N_14227,N_13710,N_13832);
nand U14228 (N_14228,N_13730,N_13868);
nor U14229 (N_14229,N_13668,N_13789);
nand U14230 (N_14230,N_13988,N_13640);
nor U14231 (N_14231,N_13552,N_13729);
nand U14232 (N_14232,N_13856,N_13596);
and U14233 (N_14233,N_13737,N_13720);
nand U14234 (N_14234,N_13930,N_13996);
xor U14235 (N_14235,N_13879,N_13854);
nand U14236 (N_14236,N_13677,N_13784);
nor U14237 (N_14237,N_13850,N_13513);
nand U14238 (N_14238,N_13697,N_13632);
nand U14239 (N_14239,N_13734,N_13947);
or U14240 (N_14240,N_13613,N_13669);
or U14241 (N_14241,N_13723,N_13748);
and U14242 (N_14242,N_13649,N_13560);
and U14243 (N_14243,N_13524,N_13624);
or U14244 (N_14244,N_13874,N_13651);
or U14245 (N_14245,N_13740,N_13592);
nor U14246 (N_14246,N_13959,N_13678);
and U14247 (N_14247,N_13622,N_13563);
and U14248 (N_14248,N_13725,N_13995);
nor U14249 (N_14249,N_13948,N_13786);
or U14250 (N_14250,N_13621,N_13824);
nand U14251 (N_14251,N_13829,N_13886);
or U14252 (N_14252,N_13984,N_13560);
nor U14253 (N_14253,N_13723,N_13655);
and U14254 (N_14254,N_13527,N_13629);
nor U14255 (N_14255,N_13550,N_13830);
xnor U14256 (N_14256,N_13840,N_13863);
nor U14257 (N_14257,N_13817,N_13981);
nor U14258 (N_14258,N_13927,N_13530);
nand U14259 (N_14259,N_13919,N_13904);
and U14260 (N_14260,N_13673,N_13993);
nand U14261 (N_14261,N_13561,N_13586);
or U14262 (N_14262,N_13744,N_13940);
or U14263 (N_14263,N_13568,N_13648);
nand U14264 (N_14264,N_13581,N_13567);
nor U14265 (N_14265,N_13596,N_13960);
nand U14266 (N_14266,N_13997,N_13791);
or U14267 (N_14267,N_13556,N_13586);
nand U14268 (N_14268,N_13520,N_13535);
or U14269 (N_14269,N_13695,N_13899);
or U14270 (N_14270,N_13642,N_13511);
and U14271 (N_14271,N_13832,N_13538);
nand U14272 (N_14272,N_13753,N_13980);
nor U14273 (N_14273,N_13974,N_13890);
and U14274 (N_14274,N_13752,N_13743);
or U14275 (N_14275,N_13754,N_13808);
nand U14276 (N_14276,N_13705,N_13752);
nor U14277 (N_14277,N_13938,N_13944);
nor U14278 (N_14278,N_13578,N_13987);
and U14279 (N_14279,N_13754,N_13669);
and U14280 (N_14280,N_13617,N_13622);
nand U14281 (N_14281,N_13805,N_13723);
or U14282 (N_14282,N_13629,N_13521);
nor U14283 (N_14283,N_13647,N_13910);
nor U14284 (N_14284,N_13521,N_13728);
nand U14285 (N_14285,N_13856,N_13901);
nand U14286 (N_14286,N_13836,N_13959);
or U14287 (N_14287,N_13957,N_13899);
and U14288 (N_14288,N_13798,N_13825);
nand U14289 (N_14289,N_13701,N_13783);
or U14290 (N_14290,N_13514,N_13829);
nor U14291 (N_14291,N_13908,N_13798);
and U14292 (N_14292,N_13737,N_13924);
and U14293 (N_14293,N_13634,N_13552);
xnor U14294 (N_14294,N_13626,N_13688);
or U14295 (N_14295,N_13740,N_13579);
nand U14296 (N_14296,N_13590,N_13893);
and U14297 (N_14297,N_13760,N_13929);
nor U14298 (N_14298,N_13511,N_13925);
xnor U14299 (N_14299,N_13697,N_13624);
nand U14300 (N_14300,N_13806,N_13606);
nand U14301 (N_14301,N_13578,N_13915);
and U14302 (N_14302,N_13938,N_13799);
xnor U14303 (N_14303,N_13688,N_13544);
and U14304 (N_14304,N_13601,N_13504);
nand U14305 (N_14305,N_13973,N_13754);
or U14306 (N_14306,N_13750,N_13505);
nand U14307 (N_14307,N_13714,N_13708);
nand U14308 (N_14308,N_13959,N_13506);
or U14309 (N_14309,N_13671,N_13776);
and U14310 (N_14310,N_13781,N_13505);
and U14311 (N_14311,N_13880,N_13979);
nand U14312 (N_14312,N_13514,N_13533);
nor U14313 (N_14313,N_13642,N_13750);
or U14314 (N_14314,N_13894,N_13549);
or U14315 (N_14315,N_13939,N_13910);
nand U14316 (N_14316,N_13963,N_13949);
nand U14317 (N_14317,N_13960,N_13674);
or U14318 (N_14318,N_13639,N_13790);
or U14319 (N_14319,N_13995,N_13518);
nand U14320 (N_14320,N_13902,N_13649);
or U14321 (N_14321,N_13650,N_13505);
and U14322 (N_14322,N_13900,N_13513);
nand U14323 (N_14323,N_13708,N_13664);
and U14324 (N_14324,N_13766,N_13999);
nor U14325 (N_14325,N_13753,N_13942);
nand U14326 (N_14326,N_13588,N_13525);
and U14327 (N_14327,N_13513,N_13954);
nand U14328 (N_14328,N_13710,N_13949);
nor U14329 (N_14329,N_13903,N_13832);
or U14330 (N_14330,N_13726,N_13819);
or U14331 (N_14331,N_13964,N_13662);
nor U14332 (N_14332,N_13814,N_13932);
nor U14333 (N_14333,N_13653,N_13962);
or U14334 (N_14334,N_13534,N_13637);
or U14335 (N_14335,N_13905,N_13532);
nor U14336 (N_14336,N_13783,N_13534);
nor U14337 (N_14337,N_13801,N_13821);
nor U14338 (N_14338,N_13655,N_13908);
or U14339 (N_14339,N_13717,N_13678);
and U14340 (N_14340,N_13505,N_13601);
nor U14341 (N_14341,N_13895,N_13557);
and U14342 (N_14342,N_13902,N_13623);
and U14343 (N_14343,N_13832,N_13631);
or U14344 (N_14344,N_13518,N_13986);
nor U14345 (N_14345,N_13943,N_13734);
or U14346 (N_14346,N_13815,N_13817);
nor U14347 (N_14347,N_13937,N_13675);
nor U14348 (N_14348,N_13921,N_13555);
nor U14349 (N_14349,N_13927,N_13942);
nor U14350 (N_14350,N_13794,N_13787);
nor U14351 (N_14351,N_13894,N_13677);
nor U14352 (N_14352,N_13654,N_13940);
and U14353 (N_14353,N_13924,N_13668);
or U14354 (N_14354,N_13591,N_13934);
nor U14355 (N_14355,N_13503,N_13778);
or U14356 (N_14356,N_13756,N_13989);
nor U14357 (N_14357,N_13576,N_13661);
and U14358 (N_14358,N_13772,N_13646);
or U14359 (N_14359,N_13736,N_13992);
or U14360 (N_14360,N_13996,N_13717);
and U14361 (N_14361,N_13917,N_13696);
xor U14362 (N_14362,N_13945,N_13913);
or U14363 (N_14363,N_13628,N_13805);
and U14364 (N_14364,N_13558,N_13852);
and U14365 (N_14365,N_13826,N_13853);
xor U14366 (N_14366,N_13912,N_13527);
nand U14367 (N_14367,N_13568,N_13954);
and U14368 (N_14368,N_13611,N_13654);
nor U14369 (N_14369,N_13959,N_13881);
and U14370 (N_14370,N_13850,N_13565);
nor U14371 (N_14371,N_13685,N_13502);
or U14372 (N_14372,N_13629,N_13692);
nand U14373 (N_14373,N_13945,N_13992);
nand U14374 (N_14374,N_13752,N_13779);
nand U14375 (N_14375,N_13701,N_13703);
nor U14376 (N_14376,N_13683,N_13805);
nor U14377 (N_14377,N_13850,N_13598);
or U14378 (N_14378,N_13578,N_13622);
nor U14379 (N_14379,N_13793,N_13502);
nand U14380 (N_14380,N_13652,N_13675);
or U14381 (N_14381,N_13516,N_13575);
nor U14382 (N_14382,N_13501,N_13554);
nand U14383 (N_14383,N_13741,N_13931);
or U14384 (N_14384,N_13800,N_13666);
and U14385 (N_14385,N_13640,N_13752);
or U14386 (N_14386,N_13754,N_13847);
or U14387 (N_14387,N_13684,N_13883);
nand U14388 (N_14388,N_13936,N_13729);
or U14389 (N_14389,N_13770,N_13590);
nor U14390 (N_14390,N_13640,N_13585);
and U14391 (N_14391,N_13957,N_13552);
and U14392 (N_14392,N_13926,N_13961);
or U14393 (N_14393,N_13806,N_13944);
or U14394 (N_14394,N_13701,N_13821);
nand U14395 (N_14395,N_13637,N_13732);
nor U14396 (N_14396,N_13649,N_13816);
nor U14397 (N_14397,N_13769,N_13923);
or U14398 (N_14398,N_13682,N_13844);
or U14399 (N_14399,N_13932,N_13878);
nand U14400 (N_14400,N_13845,N_13983);
xor U14401 (N_14401,N_13663,N_13730);
nand U14402 (N_14402,N_13903,N_13708);
or U14403 (N_14403,N_13711,N_13503);
nor U14404 (N_14404,N_13669,N_13721);
nand U14405 (N_14405,N_13809,N_13591);
nand U14406 (N_14406,N_13600,N_13861);
and U14407 (N_14407,N_13502,N_13557);
nor U14408 (N_14408,N_13984,N_13597);
or U14409 (N_14409,N_13898,N_13706);
nand U14410 (N_14410,N_13617,N_13671);
and U14411 (N_14411,N_13967,N_13767);
nor U14412 (N_14412,N_13875,N_13560);
nor U14413 (N_14413,N_13914,N_13871);
nand U14414 (N_14414,N_13756,N_13894);
nor U14415 (N_14415,N_13750,N_13609);
and U14416 (N_14416,N_13712,N_13750);
or U14417 (N_14417,N_13977,N_13700);
or U14418 (N_14418,N_13829,N_13772);
nor U14419 (N_14419,N_13740,N_13696);
and U14420 (N_14420,N_13558,N_13633);
nand U14421 (N_14421,N_13733,N_13696);
and U14422 (N_14422,N_13845,N_13574);
or U14423 (N_14423,N_13727,N_13575);
nand U14424 (N_14424,N_13766,N_13555);
or U14425 (N_14425,N_13671,N_13772);
or U14426 (N_14426,N_13978,N_13751);
nand U14427 (N_14427,N_13977,N_13837);
nor U14428 (N_14428,N_13585,N_13735);
and U14429 (N_14429,N_13791,N_13686);
or U14430 (N_14430,N_13668,N_13736);
xor U14431 (N_14431,N_13911,N_13902);
xnor U14432 (N_14432,N_13747,N_13629);
nor U14433 (N_14433,N_13983,N_13546);
and U14434 (N_14434,N_13611,N_13736);
or U14435 (N_14435,N_13929,N_13997);
and U14436 (N_14436,N_13841,N_13571);
and U14437 (N_14437,N_13966,N_13660);
and U14438 (N_14438,N_13836,N_13941);
or U14439 (N_14439,N_13609,N_13625);
or U14440 (N_14440,N_13610,N_13518);
nand U14441 (N_14441,N_13575,N_13663);
nor U14442 (N_14442,N_13971,N_13681);
nor U14443 (N_14443,N_13898,N_13907);
nand U14444 (N_14444,N_13786,N_13936);
xnor U14445 (N_14445,N_13710,N_13517);
nor U14446 (N_14446,N_13807,N_13574);
nand U14447 (N_14447,N_13676,N_13582);
or U14448 (N_14448,N_13715,N_13653);
and U14449 (N_14449,N_13742,N_13816);
or U14450 (N_14450,N_13808,N_13568);
and U14451 (N_14451,N_13508,N_13546);
and U14452 (N_14452,N_13820,N_13921);
and U14453 (N_14453,N_13565,N_13687);
or U14454 (N_14454,N_13837,N_13662);
and U14455 (N_14455,N_13662,N_13628);
and U14456 (N_14456,N_13723,N_13686);
or U14457 (N_14457,N_13605,N_13761);
and U14458 (N_14458,N_13608,N_13693);
or U14459 (N_14459,N_13664,N_13957);
or U14460 (N_14460,N_13693,N_13959);
or U14461 (N_14461,N_13608,N_13541);
nor U14462 (N_14462,N_13706,N_13809);
nand U14463 (N_14463,N_13812,N_13521);
nor U14464 (N_14464,N_13893,N_13848);
nor U14465 (N_14465,N_13566,N_13768);
or U14466 (N_14466,N_13717,N_13831);
or U14467 (N_14467,N_13647,N_13831);
nand U14468 (N_14468,N_13896,N_13944);
nor U14469 (N_14469,N_13522,N_13671);
nand U14470 (N_14470,N_13971,N_13987);
nand U14471 (N_14471,N_13848,N_13795);
and U14472 (N_14472,N_13573,N_13528);
nor U14473 (N_14473,N_13791,N_13900);
nand U14474 (N_14474,N_13710,N_13962);
and U14475 (N_14475,N_13861,N_13694);
nand U14476 (N_14476,N_13533,N_13973);
and U14477 (N_14477,N_13814,N_13997);
and U14478 (N_14478,N_13811,N_13807);
nor U14479 (N_14479,N_13612,N_13998);
nor U14480 (N_14480,N_13791,N_13925);
nor U14481 (N_14481,N_13675,N_13579);
or U14482 (N_14482,N_13667,N_13585);
nand U14483 (N_14483,N_13907,N_13708);
and U14484 (N_14484,N_13868,N_13553);
nand U14485 (N_14485,N_13787,N_13997);
nor U14486 (N_14486,N_13710,N_13564);
and U14487 (N_14487,N_13815,N_13889);
and U14488 (N_14488,N_13520,N_13991);
nor U14489 (N_14489,N_13632,N_13561);
and U14490 (N_14490,N_13868,N_13820);
or U14491 (N_14491,N_13636,N_13966);
and U14492 (N_14492,N_13835,N_13825);
and U14493 (N_14493,N_13990,N_13549);
nor U14494 (N_14494,N_13906,N_13864);
or U14495 (N_14495,N_13792,N_13788);
nor U14496 (N_14496,N_13768,N_13735);
nor U14497 (N_14497,N_13533,N_13541);
nor U14498 (N_14498,N_13792,N_13959);
or U14499 (N_14499,N_13908,N_13532);
nand U14500 (N_14500,N_14278,N_14232);
nor U14501 (N_14501,N_14431,N_14148);
nand U14502 (N_14502,N_14184,N_14300);
nor U14503 (N_14503,N_14306,N_14233);
and U14504 (N_14504,N_14066,N_14017);
nand U14505 (N_14505,N_14238,N_14458);
nand U14506 (N_14506,N_14234,N_14104);
and U14507 (N_14507,N_14413,N_14373);
or U14508 (N_14508,N_14029,N_14489);
or U14509 (N_14509,N_14124,N_14016);
nor U14510 (N_14510,N_14209,N_14085);
nand U14511 (N_14511,N_14275,N_14246);
nand U14512 (N_14512,N_14331,N_14376);
nand U14513 (N_14513,N_14102,N_14341);
or U14514 (N_14514,N_14022,N_14248);
or U14515 (N_14515,N_14342,N_14173);
xnor U14516 (N_14516,N_14031,N_14440);
nand U14517 (N_14517,N_14150,N_14055);
nand U14518 (N_14518,N_14486,N_14210);
and U14519 (N_14519,N_14129,N_14044);
nor U14520 (N_14520,N_14059,N_14038);
or U14521 (N_14521,N_14241,N_14294);
nor U14522 (N_14522,N_14033,N_14012);
nand U14523 (N_14523,N_14023,N_14324);
or U14524 (N_14524,N_14349,N_14409);
or U14525 (N_14525,N_14302,N_14109);
and U14526 (N_14526,N_14323,N_14135);
and U14527 (N_14527,N_14309,N_14107);
or U14528 (N_14528,N_14236,N_14161);
nand U14529 (N_14529,N_14137,N_14158);
nor U14530 (N_14530,N_14179,N_14384);
nor U14531 (N_14531,N_14126,N_14213);
and U14532 (N_14532,N_14277,N_14292);
and U14533 (N_14533,N_14403,N_14163);
nor U14534 (N_14534,N_14100,N_14344);
and U14535 (N_14535,N_14400,N_14370);
or U14536 (N_14536,N_14166,N_14103);
nor U14537 (N_14537,N_14174,N_14045);
or U14538 (N_14538,N_14139,N_14439);
and U14539 (N_14539,N_14426,N_14216);
and U14540 (N_14540,N_14473,N_14145);
or U14541 (N_14541,N_14401,N_14206);
nor U14542 (N_14542,N_14030,N_14243);
or U14543 (N_14543,N_14437,N_14357);
and U14544 (N_14544,N_14498,N_14024);
or U14545 (N_14545,N_14385,N_14254);
nand U14546 (N_14546,N_14147,N_14361);
and U14547 (N_14547,N_14408,N_14308);
nand U14548 (N_14548,N_14272,N_14194);
nand U14549 (N_14549,N_14001,N_14436);
and U14550 (N_14550,N_14168,N_14366);
nor U14551 (N_14551,N_14050,N_14032);
and U14552 (N_14552,N_14339,N_14482);
and U14553 (N_14553,N_14425,N_14072);
nand U14554 (N_14554,N_14322,N_14328);
or U14555 (N_14555,N_14281,N_14468);
xnor U14556 (N_14556,N_14470,N_14442);
nand U14557 (N_14557,N_14493,N_14132);
or U14558 (N_14558,N_14424,N_14247);
or U14559 (N_14559,N_14364,N_14067);
nand U14560 (N_14560,N_14221,N_14289);
and U14561 (N_14561,N_14064,N_14201);
or U14562 (N_14562,N_14305,N_14368);
and U14563 (N_14563,N_14013,N_14242);
and U14564 (N_14564,N_14097,N_14367);
nand U14565 (N_14565,N_14006,N_14393);
and U14566 (N_14566,N_14450,N_14093);
nand U14567 (N_14567,N_14405,N_14452);
and U14568 (N_14568,N_14231,N_14467);
or U14569 (N_14569,N_14003,N_14229);
nor U14570 (N_14570,N_14418,N_14407);
nand U14571 (N_14571,N_14215,N_14313);
or U14572 (N_14572,N_14297,N_14079);
or U14573 (N_14573,N_14378,N_14274);
or U14574 (N_14574,N_14360,N_14390);
and U14575 (N_14575,N_14268,N_14088);
and U14576 (N_14576,N_14453,N_14181);
and U14577 (N_14577,N_14200,N_14058);
nor U14578 (N_14578,N_14451,N_14435);
nand U14579 (N_14579,N_14220,N_14375);
nor U14580 (N_14580,N_14081,N_14295);
and U14581 (N_14581,N_14414,N_14134);
and U14582 (N_14582,N_14253,N_14034);
and U14583 (N_14583,N_14164,N_14138);
nor U14584 (N_14584,N_14252,N_14388);
nand U14585 (N_14585,N_14293,N_14131);
nand U14586 (N_14586,N_14040,N_14185);
and U14587 (N_14587,N_14290,N_14165);
and U14588 (N_14588,N_14217,N_14020);
nor U14589 (N_14589,N_14307,N_14061);
and U14590 (N_14590,N_14052,N_14264);
nand U14591 (N_14591,N_14039,N_14410);
and U14592 (N_14592,N_14394,N_14494);
nand U14593 (N_14593,N_14351,N_14392);
xor U14594 (N_14594,N_14154,N_14094);
nand U14595 (N_14595,N_14149,N_14311);
nor U14596 (N_14596,N_14089,N_14495);
and U14597 (N_14597,N_14069,N_14472);
nor U14598 (N_14598,N_14249,N_14283);
and U14599 (N_14599,N_14214,N_14075);
nand U14600 (N_14600,N_14071,N_14212);
nor U14601 (N_14601,N_14086,N_14343);
or U14602 (N_14602,N_14228,N_14002);
and U14603 (N_14603,N_14488,N_14317);
nand U14604 (N_14604,N_14255,N_14333);
or U14605 (N_14605,N_14389,N_14224);
or U14606 (N_14606,N_14207,N_14019);
and U14607 (N_14607,N_14225,N_14186);
or U14608 (N_14608,N_14411,N_14227);
nor U14609 (N_14609,N_14329,N_14198);
and U14610 (N_14610,N_14448,N_14485);
or U14611 (N_14611,N_14118,N_14026);
nand U14612 (N_14612,N_14122,N_14304);
nor U14613 (N_14613,N_14128,N_14320);
and U14614 (N_14614,N_14011,N_14053);
nor U14615 (N_14615,N_14037,N_14007);
and U14616 (N_14616,N_14258,N_14415);
or U14617 (N_14617,N_14018,N_14171);
and U14618 (N_14618,N_14116,N_14204);
nand U14619 (N_14619,N_14459,N_14065);
nor U14620 (N_14620,N_14298,N_14434);
and U14621 (N_14621,N_14355,N_14062);
nor U14622 (N_14622,N_14159,N_14133);
and U14623 (N_14623,N_14162,N_14091);
nor U14624 (N_14624,N_14199,N_14365);
nor U14625 (N_14625,N_14345,N_14005);
or U14626 (N_14626,N_14074,N_14047);
nand U14627 (N_14627,N_14348,N_14314);
nor U14628 (N_14628,N_14422,N_14196);
or U14629 (N_14629,N_14175,N_14178);
or U14630 (N_14630,N_14021,N_14136);
or U14631 (N_14631,N_14101,N_14108);
xor U14632 (N_14632,N_14155,N_14025);
nand U14633 (N_14633,N_14014,N_14077);
and U14634 (N_14634,N_14337,N_14379);
and U14635 (N_14635,N_14326,N_14219);
nor U14636 (N_14636,N_14280,N_14099);
nor U14637 (N_14637,N_14444,N_14261);
nor U14638 (N_14638,N_14446,N_14015);
and U14639 (N_14639,N_14478,N_14499);
or U14640 (N_14640,N_14096,N_14152);
and U14641 (N_14641,N_14237,N_14433);
nand U14642 (N_14642,N_14338,N_14170);
nor U14643 (N_14643,N_14296,N_14256);
or U14644 (N_14644,N_14250,N_14358);
or U14645 (N_14645,N_14299,N_14176);
nand U14646 (N_14646,N_14190,N_14105);
and U14647 (N_14647,N_14265,N_14336);
and U14648 (N_14648,N_14363,N_14078);
and U14649 (N_14649,N_14208,N_14113);
and U14650 (N_14650,N_14117,N_14353);
and U14651 (N_14651,N_14193,N_14288);
and U14652 (N_14652,N_14406,N_14454);
or U14653 (N_14653,N_14449,N_14027);
nand U14654 (N_14654,N_14203,N_14028);
and U14655 (N_14655,N_14443,N_14460);
and U14656 (N_14656,N_14354,N_14497);
and U14657 (N_14657,N_14279,N_14447);
or U14658 (N_14658,N_14475,N_14235);
xor U14659 (N_14659,N_14192,N_14477);
and U14660 (N_14660,N_14483,N_14245);
and U14661 (N_14661,N_14466,N_14240);
nor U14662 (N_14662,N_14257,N_14464);
and U14663 (N_14663,N_14462,N_14391);
nor U14664 (N_14664,N_14319,N_14315);
or U14665 (N_14665,N_14041,N_14419);
nor U14666 (N_14666,N_14262,N_14141);
nor U14667 (N_14667,N_14153,N_14119);
nor U14668 (N_14668,N_14356,N_14087);
and U14669 (N_14669,N_14092,N_14432);
and U14670 (N_14670,N_14143,N_14423);
and U14671 (N_14671,N_14350,N_14396);
nor U14672 (N_14672,N_14082,N_14120);
and U14673 (N_14673,N_14397,N_14282);
nand U14674 (N_14674,N_14455,N_14416);
nor U14675 (N_14675,N_14172,N_14438);
and U14676 (N_14676,N_14112,N_14043);
nor U14677 (N_14677,N_14267,N_14189);
and U14678 (N_14678,N_14270,N_14010);
or U14679 (N_14679,N_14068,N_14266);
nand U14680 (N_14680,N_14481,N_14377);
nor U14681 (N_14681,N_14076,N_14312);
nor U14682 (N_14682,N_14110,N_14427);
nor U14683 (N_14683,N_14404,N_14146);
nor U14684 (N_14684,N_14310,N_14445);
nor U14685 (N_14685,N_14430,N_14054);
nand U14686 (N_14686,N_14476,N_14321);
nor U14687 (N_14687,N_14084,N_14035);
nor U14688 (N_14688,N_14125,N_14276);
and U14689 (N_14689,N_14048,N_14441);
xor U14690 (N_14690,N_14420,N_14380);
or U14691 (N_14691,N_14332,N_14183);
and U14692 (N_14692,N_14083,N_14273);
and U14693 (N_14693,N_14340,N_14382);
nor U14694 (N_14694,N_14421,N_14070);
xnor U14695 (N_14695,N_14359,N_14008);
and U14696 (N_14696,N_14490,N_14057);
and U14697 (N_14697,N_14301,N_14098);
or U14698 (N_14698,N_14090,N_14325);
xor U14699 (N_14699,N_14195,N_14417);
and U14700 (N_14700,N_14398,N_14352);
nand U14701 (N_14701,N_14095,N_14334);
and U14702 (N_14702,N_14484,N_14480);
nand U14703 (N_14703,N_14156,N_14457);
nand U14704 (N_14704,N_14197,N_14374);
nor U14705 (N_14705,N_14479,N_14036);
or U14706 (N_14706,N_14042,N_14412);
nor U14707 (N_14707,N_14263,N_14182);
nor U14708 (N_14708,N_14169,N_14335);
or U14709 (N_14709,N_14383,N_14063);
nor U14710 (N_14710,N_14271,N_14461);
nand U14711 (N_14711,N_14303,N_14318);
nand U14712 (N_14712,N_14151,N_14130);
and U14713 (N_14713,N_14144,N_14188);
nand U14714 (N_14714,N_14429,N_14046);
and U14715 (N_14715,N_14140,N_14239);
and U14716 (N_14716,N_14284,N_14160);
nor U14717 (N_14717,N_14123,N_14114);
nor U14718 (N_14718,N_14226,N_14330);
nor U14719 (N_14719,N_14106,N_14286);
and U14720 (N_14720,N_14491,N_14463);
and U14721 (N_14721,N_14496,N_14080);
or U14722 (N_14722,N_14381,N_14191);
nand U14723 (N_14723,N_14287,N_14218);
nand U14724 (N_14724,N_14399,N_14060);
nand U14725 (N_14725,N_14492,N_14291);
nor U14726 (N_14726,N_14259,N_14115);
or U14727 (N_14727,N_14372,N_14230);
and U14728 (N_14728,N_14073,N_14369);
and U14729 (N_14729,N_14049,N_14387);
and U14730 (N_14730,N_14395,N_14000);
nand U14731 (N_14731,N_14428,N_14142);
nand U14732 (N_14732,N_14269,N_14051);
nand U14733 (N_14733,N_14222,N_14202);
nand U14734 (N_14734,N_14180,N_14402);
xnor U14735 (N_14735,N_14223,N_14471);
and U14736 (N_14736,N_14009,N_14244);
and U14737 (N_14737,N_14167,N_14371);
and U14738 (N_14738,N_14346,N_14316);
nand U14739 (N_14739,N_14474,N_14111);
and U14740 (N_14740,N_14004,N_14487);
and U14741 (N_14741,N_14362,N_14465);
and U14742 (N_14742,N_14469,N_14205);
or U14743 (N_14743,N_14456,N_14347);
nor U14744 (N_14744,N_14285,N_14327);
and U14745 (N_14745,N_14157,N_14211);
nor U14746 (N_14746,N_14121,N_14177);
and U14747 (N_14747,N_14056,N_14251);
nand U14748 (N_14748,N_14127,N_14187);
or U14749 (N_14749,N_14386,N_14260);
or U14750 (N_14750,N_14306,N_14373);
nor U14751 (N_14751,N_14269,N_14395);
nand U14752 (N_14752,N_14170,N_14232);
nor U14753 (N_14753,N_14134,N_14061);
nand U14754 (N_14754,N_14080,N_14387);
or U14755 (N_14755,N_14111,N_14345);
nand U14756 (N_14756,N_14428,N_14326);
nand U14757 (N_14757,N_14369,N_14474);
nor U14758 (N_14758,N_14379,N_14033);
and U14759 (N_14759,N_14442,N_14490);
and U14760 (N_14760,N_14165,N_14492);
nor U14761 (N_14761,N_14459,N_14271);
and U14762 (N_14762,N_14320,N_14498);
or U14763 (N_14763,N_14383,N_14288);
and U14764 (N_14764,N_14420,N_14229);
nand U14765 (N_14765,N_14492,N_14219);
and U14766 (N_14766,N_14410,N_14219);
and U14767 (N_14767,N_14143,N_14296);
and U14768 (N_14768,N_14449,N_14136);
or U14769 (N_14769,N_14278,N_14260);
or U14770 (N_14770,N_14199,N_14260);
and U14771 (N_14771,N_14166,N_14455);
and U14772 (N_14772,N_14282,N_14491);
nor U14773 (N_14773,N_14363,N_14011);
xnor U14774 (N_14774,N_14231,N_14244);
or U14775 (N_14775,N_14106,N_14198);
and U14776 (N_14776,N_14300,N_14176);
and U14777 (N_14777,N_14301,N_14305);
and U14778 (N_14778,N_14007,N_14018);
nand U14779 (N_14779,N_14192,N_14422);
nand U14780 (N_14780,N_14135,N_14370);
or U14781 (N_14781,N_14021,N_14429);
nand U14782 (N_14782,N_14266,N_14140);
or U14783 (N_14783,N_14212,N_14261);
nor U14784 (N_14784,N_14046,N_14031);
nand U14785 (N_14785,N_14085,N_14064);
or U14786 (N_14786,N_14287,N_14173);
nand U14787 (N_14787,N_14299,N_14381);
nand U14788 (N_14788,N_14227,N_14285);
and U14789 (N_14789,N_14200,N_14344);
nand U14790 (N_14790,N_14169,N_14224);
nand U14791 (N_14791,N_14187,N_14120);
and U14792 (N_14792,N_14155,N_14286);
and U14793 (N_14793,N_14333,N_14177);
or U14794 (N_14794,N_14427,N_14384);
or U14795 (N_14795,N_14419,N_14165);
nor U14796 (N_14796,N_14445,N_14400);
nand U14797 (N_14797,N_14024,N_14344);
nor U14798 (N_14798,N_14015,N_14069);
nor U14799 (N_14799,N_14492,N_14245);
nor U14800 (N_14800,N_14056,N_14152);
nor U14801 (N_14801,N_14310,N_14154);
or U14802 (N_14802,N_14149,N_14102);
and U14803 (N_14803,N_14027,N_14023);
nor U14804 (N_14804,N_14144,N_14466);
and U14805 (N_14805,N_14422,N_14355);
nand U14806 (N_14806,N_14090,N_14069);
or U14807 (N_14807,N_14357,N_14352);
nand U14808 (N_14808,N_14458,N_14090);
or U14809 (N_14809,N_14018,N_14464);
nor U14810 (N_14810,N_14208,N_14321);
or U14811 (N_14811,N_14195,N_14019);
or U14812 (N_14812,N_14497,N_14337);
or U14813 (N_14813,N_14209,N_14314);
and U14814 (N_14814,N_14155,N_14049);
nand U14815 (N_14815,N_14167,N_14428);
nand U14816 (N_14816,N_14282,N_14128);
nor U14817 (N_14817,N_14219,N_14120);
nor U14818 (N_14818,N_14431,N_14320);
nand U14819 (N_14819,N_14440,N_14088);
and U14820 (N_14820,N_14024,N_14430);
nand U14821 (N_14821,N_14151,N_14308);
nand U14822 (N_14822,N_14056,N_14403);
and U14823 (N_14823,N_14194,N_14047);
and U14824 (N_14824,N_14328,N_14374);
nand U14825 (N_14825,N_14372,N_14442);
and U14826 (N_14826,N_14290,N_14429);
nor U14827 (N_14827,N_14406,N_14379);
or U14828 (N_14828,N_14282,N_14205);
nor U14829 (N_14829,N_14035,N_14498);
and U14830 (N_14830,N_14400,N_14379);
xor U14831 (N_14831,N_14051,N_14215);
nor U14832 (N_14832,N_14313,N_14129);
and U14833 (N_14833,N_14113,N_14314);
and U14834 (N_14834,N_14309,N_14145);
nor U14835 (N_14835,N_14215,N_14070);
nand U14836 (N_14836,N_14220,N_14112);
nand U14837 (N_14837,N_14020,N_14210);
nand U14838 (N_14838,N_14493,N_14091);
and U14839 (N_14839,N_14491,N_14306);
or U14840 (N_14840,N_14070,N_14023);
nor U14841 (N_14841,N_14395,N_14484);
or U14842 (N_14842,N_14409,N_14396);
and U14843 (N_14843,N_14172,N_14125);
nand U14844 (N_14844,N_14133,N_14033);
nand U14845 (N_14845,N_14013,N_14403);
xnor U14846 (N_14846,N_14052,N_14046);
or U14847 (N_14847,N_14042,N_14136);
nor U14848 (N_14848,N_14473,N_14007);
nand U14849 (N_14849,N_14022,N_14411);
and U14850 (N_14850,N_14299,N_14251);
and U14851 (N_14851,N_14314,N_14464);
nand U14852 (N_14852,N_14104,N_14398);
nand U14853 (N_14853,N_14431,N_14032);
nor U14854 (N_14854,N_14059,N_14203);
nand U14855 (N_14855,N_14417,N_14297);
or U14856 (N_14856,N_14194,N_14331);
or U14857 (N_14857,N_14424,N_14273);
nand U14858 (N_14858,N_14263,N_14466);
or U14859 (N_14859,N_14222,N_14474);
nand U14860 (N_14860,N_14251,N_14103);
or U14861 (N_14861,N_14383,N_14179);
nand U14862 (N_14862,N_14109,N_14338);
nor U14863 (N_14863,N_14015,N_14205);
and U14864 (N_14864,N_14498,N_14039);
nor U14865 (N_14865,N_14114,N_14112);
and U14866 (N_14866,N_14211,N_14163);
or U14867 (N_14867,N_14326,N_14442);
and U14868 (N_14868,N_14177,N_14151);
nor U14869 (N_14869,N_14308,N_14000);
and U14870 (N_14870,N_14092,N_14067);
xor U14871 (N_14871,N_14345,N_14225);
and U14872 (N_14872,N_14114,N_14210);
nand U14873 (N_14873,N_14343,N_14435);
and U14874 (N_14874,N_14116,N_14141);
or U14875 (N_14875,N_14160,N_14342);
or U14876 (N_14876,N_14210,N_14141);
nand U14877 (N_14877,N_14377,N_14269);
and U14878 (N_14878,N_14066,N_14020);
nand U14879 (N_14879,N_14024,N_14393);
nand U14880 (N_14880,N_14438,N_14208);
nor U14881 (N_14881,N_14232,N_14153);
nand U14882 (N_14882,N_14428,N_14137);
and U14883 (N_14883,N_14361,N_14036);
nand U14884 (N_14884,N_14125,N_14242);
nand U14885 (N_14885,N_14272,N_14322);
nor U14886 (N_14886,N_14071,N_14213);
and U14887 (N_14887,N_14072,N_14070);
or U14888 (N_14888,N_14111,N_14236);
or U14889 (N_14889,N_14065,N_14299);
or U14890 (N_14890,N_14337,N_14267);
nor U14891 (N_14891,N_14051,N_14406);
nor U14892 (N_14892,N_14290,N_14173);
nand U14893 (N_14893,N_14298,N_14107);
nor U14894 (N_14894,N_14364,N_14446);
xor U14895 (N_14895,N_14151,N_14236);
or U14896 (N_14896,N_14115,N_14026);
nand U14897 (N_14897,N_14455,N_14490);
and U14898 (N_14898,N_14446,N_14215);
nor U14899 (N_14899,N_14005,N_14230);
and U14900 (N_14900,N_14198,N_14352);
or U14901 (N_14901,N_14434,N_14075);
nand U14902 (N_14902,N_14015,N_14499);
or U14903 (N_14903,N_14392,N_14357);
or U14904 (N_14904,N_14430,N_14418);
or U14905 (N_14905,N_14097,N_14297);
nor U14906 (N_14906,N_14257,N_14481);
and U14907 (N_14907,N_14162,N_14137);
nand U14908 (N_14908,N_14481,N_14217);
xnor U14909 (N_14909,N_14306,N_14462);
and U14910 (N_14910,N_14359,N_14297);
xor U14911 (N_14911,N_14380,N_14218);
xnor U14912 (N_14912,N_14152,N_14199);
nand U14913 (N_14913,N_14143,N_14056);
or U14914 (N_14914,N_14139,N_14383);
nand U14915 (N_14915,N_14472,N_14419);
nand U14916 (N_14916,N_14025,N_14290);
and U14917 (N_14917,N_14040,N_14210);
or U14918 (N_14918,N_14460,N_14001);
or U14919 (N_14919,N_14162,N_14314);
nor U14920 (N_14920,N_14303,N_14092);
or U14921 (N_14921,N_14139,N_14137);
and U14922 (N_14922,N_14491,N_14214);
or U14923 (N_14923,N_14061,N_14443);
nand U14924 (N_14924,N_14064,N_14171);
nor U14925 (N_14925,N_14213,N_14324);
or U14926 (N_14926,N_14087,N_14220);
or U14927 (N_14927,N_14172,N_14275);
nand U14928 (N_14928,N_14416,N_14423);
nor U14929 (N_14929,N_14368,N_14472);
and U14930 (N_14930,N_14250,N_14177);
or U14931 (N_14931,N_14338,N_14379);
nand U14932 (N_14932,N_14339,N_14465);
and U14933 (N_14933,N_14233,N_14091);
nand U14934 (N_14934,N_14063,N_14456);
or U14935 (N_14935,N_14485,N_14204);
nor U14936 (N_14936,N_14301,N_14304);
xnor U14937 (N_14937,N_14445,N_14094);
and U14938 (N_14938,N_14141,N_14341);
nor U14939 (N_14939,N_14405,N_14209);
and U14940 (N_14940,N_14230,N_14229);
nand U14941 (N_14941,N_14409,N_14433);
or U14942 (N_14942,N_14230,N_14326);
or U14943 (N_14943,N_14107,N_14399);
nor U14944 (N_14944,N_14097,N_14182);
or U14945 (N_14945,N_14237,N_14496);
nand U14946 (N_14946,N_14028,N_14337);
nand U14947 (N_14947,N_14255,N_14486);
or U14948 (N_14948,N_14288,N_14301);
nand U14949 (N_14949,N_14192,N_14268);
nand U14950 (N_14950,N_14360,N_14210);
and U14951 (N_14951,N_14491,N_14111);
nor U14952 (N_14952,N_14271,N_14279);
nand U14953 (N_14953,N_14379,N_14386);
or U14954 (N_14954,N_14456,N_14377);
nand U14955 (N_14955,N_14386,N_14133);
and U14956 (N_14956,N_14375,N_14385);
nor U14957 (N_14957,N_14034,N_14172);
nand U14958 (N_14958,N_14070,N_14286);
nand U14959 (N_14959,N_14037,N_14246);
nor U14960 (N_14960,N_14146,N_14336);
nor U14961 (N_14961,N_14048,N_14420);
and U14962 (N_14962,N_14149,N_14144);
nor U14963 (N_14963,N_14375,N_14459);
and U14964 (N_14964,N_14309,N_14448);
and U14965 (N_14965,N_14187,N_14136);
nand U14966 (N_14966,N_14287,N_14350);
and U14967 (N_14967,N_14356,N_14178);
nand U14968 (N_14968,N_14228,N_14044);
or U14969 (N_14969,N_14148,N_14156);
nor U14970 (N_14970,N_14224,N_14417);
nor U14971 (N_14971,N_14450,N_14493);
xnor U14972 (N_14972,N_14127,N_14465);
or U14973 (N_14973,N_14308,N_14186);
nor U14974 (N_14974,N_14318,N_14221);
or U14975 (N_14975,N_14459,N_14022);
and U14976 (N_14976,N_14190,N_14246);
and U14977 (N_14977,N_14078,N_14018);
and U14978 (N_14978,N_14278,N_14264);
and U14979 (N_14979,N_14153,N_14337);
and U14980 (N_14980,N_14218,N_14018);
or U14981 (N_14981,N_14122,N_14492);
and U14982 (N_14982,N_14035,N_14447);
or U14983 (N_14983,N_14052,N_14406);
nor U14984 (N_14984,N_14367,N_14249);
and U14985 (N_14985,N_14140,N_14339);
nor U14986 (N_14986,N_14377,N_14385);
or U14987 (N_14987,N_14446,N_14466);
nor U14988 (N_14988,N_14367,N_14268);
nor U14989 (N_14989,N_14133,N_14210);
nand U14990 (N_14990,N_14411,N_14038);
and U14991 (N_14991,N_14194,N_14410);
nand U14992 (N_14992,N_14297,N_14189);
nor U14993 (N_14993,N_14029,N_14057);
nand U14994 (N_14994,N_14208,N_14201);
nand U14995 (N_14995,N_14382,N_14114);
or U14996 (N_14996,N_14328,N_14292);
nor U14997 (N_14997,N_14113,N_14382);
and U14998 (N_14998,N_14448,N_14282);
nand U14999 (N_14999,N_14423,N_14259);
nor U15000 (N_15000,N_14791,N_14811);
nor U15001 (N_15001,N_14943,N_14795);
or U15002 (N_15002,N_14886,N_14860);
and U15003 (N_15003,N_14808,N_14897);
nand U15004 (N_15004,N_14855,N_14707);
nor U15005 (N_15005,N_14734,N_14869);
or U15006 (N_15006,N_14597,N_14879);
and U15007 (N_15007,N_14701,N_14698);
or U15008 (N_15008,N_14523,N_14673);
and U15009 (N_15009,N_14745,N_14772);
nand U15010 (N_15010,N_14946,N_14834);
and U15011 (N_15011,N_14802,N_14573);
and U15012 (N_15012,N_14562,N_14694);
nand U15013 (N_15013,N_14598,N_14748);
or U15014 (N_15014,N_14865,N_14963);
or U15015 (N_15015,N_14732,N_14526);
or U15016 (N_15016,N_14516,N_14567);
and U15017 (N_15017,N_14851,N_14611);
and U15018 (N_15018,N_14984,N_14884);
nor U15019 (N_15019,N_14789,N_14690);
or U15020 (N_15020,N_14689,N_14818);
and U15021 (N_15021,N_14557,N_14828);
nor U15022 (N_15022,N_14650,N_14661);
xnor U15023 (N_15023,N_14827,N_14665);
or U15024 (N_15024,N_14922,N_14520);
nor U15025 (N_15025,N_14569,N_14982);
nand U15026 (N_15026,N_14647,N_14655);
or U15027 (N_15027,N_14594,N_14524);
nand U15028 (N_15028,N_14646,N_14682);
and U15029 (N_15029,N_14662,N_14907);
and U15030 (N_15030,N_14841,N_14553);
xor U15031 (N_15031,N_14925,N_14586);
and U15032 (N_15032,N_14874,N_14950);
nor U15033 (N_15033,N_14730,N_14699);
and U15034 (N_15034,N_14546,N_14541);
nor U15035 (N_15035,N_14686,N_14697);
nor U15036 (N_15036,N_14550,N_14876);
nor U15037 (N_15037,N_14551,N_14660);
and U15038 (N_15038,N_14738,N_14769);
and U15039 (N_15039,N_14838,N_14857);
nor U15040 (N_15040,N_14853,N_14831);
nor U15041 (N_15041,N_14538,N_14792);
nand U15042 (N_15042,N_14637,N_14521);
and U15043 (N_15043,N_14989,N_14644);
or U15044 (N_15044,N_14608,N_14940);
or U15045 (N_15045,N_14938,N_14900);
nor U15046 (N_15046,N_14930,N_14901);
nand U15047 (N_15047,N_14672,N_14914);
or U15048 (N_15048,N_14799,N_14656);
nand U15049 (N_15049,N_14547,N_14727);
nand U15050 (N_15050,N_14592,N_14728);
nand U15051 (N_15051,N_14577,N_14558);
nand U15052 (N_15052,N_14658,N_14702);
and U15053 (N_15053,N_14926,N_14713);
or U15054 (N_15054,N_14905,N_14561);
nand U15055 (N_15055,N_14895,N_14625);
or U15056 (N_15056,N_14513,N_14812);
nand U15057 (N_15057,N_14842,N_14966);
nor U15058 (N_15058,N_14778,N_14677);
and U15059 (N_15059,N_14892,N_14962);
nor U15060 (N_15060,N_14596,N_14885);
nand U15061 (N_15061,N_14953,N_14581);
or U15062 (N_15062,N_14643,N_14934);
or U15063 (N_15063,N_14539,N_14579);
nand U15064 (N_15064,N_14839,N_14503);
and U15065 (N_15065,N_14898,N_14850);
nor U15066 (N_15066,N_14896,N_14858);
nand U15067 (N_15067,N_14584,N_14847);
nand U15068 (N_15068,N_14856,N_14729);
and U15069 (N_15069,N_14867,N_14645);
nor U15070 (N_15070,N_14525,N_14915);
and U15071 (N_15071,N_14555,N_14893);
nand U15072 (N_15072,N_14717,N_14622);
nand U15073 (N_15073,N_14969,N_14648);
or U15074 (N_15074,N_14623,N_14691);
and U15075 (N_15075,N_14754,N_14714);
or U15076 (N_15076,N_14911,N_14903);
nor U15077 (N_15077,N_14890,N_14632);
or U15078 (N_15078,N_14642,N_14935);
nor U15079 (N_15079,N_14941,N_14663);
or U15080 (N_15080,N_14837,N_14944);
or U15081 (N_15081,N_14532,N_14878);
nor U15082 (N_15082,N_14985,N_14747);
or U15083 (N_15083,N_14651,N_14704);
and U15084 (N_15084,N_14527,N_14721);
nor U15085 (N_15085,N_14640,N_14657);
nor U15086 (N_15086,N_14518,N_14751);
or U15087 (N_15087,N_14961,N_14733);
nor U15088 (N_15088,N_14829,N_14716);
nand U15089 (N_15089,N_14502,N_14774);
or U15090 (N_15090,N_14676,N_14675);
nor U15091 (N_15091,N_14861,N_14987);
and U15092 (N_15092,N_14515,N_14737);
nor U15093 (N_15093,N_14565,N_14529);
and U15094 (N_15094,N_14883,N_14544);
or U15095 (N_15095,N_14760,N_14619);
and U15096 (N_15096,N_14980,N_14788);
or U15097 (N_15097,N_14606,N_14548);
xnor U15098 (N_15098,N_14726,N_14805);
and U15099 (N_15099,N_14617,N_14820);
or U15100 (N_15100,N_14859,N_14923);
nand U15101 (N_15101,N_14904,N_14889);
or U15102 (N_15102,N_14782,N_14685);
or U15103 (N_15103,N_14758,N_14936);
and U15104 (N_15104,N_14948,N_14679);
and U15105 (N_15105,N_14986,N_14771);
or U15106 (N_15106,N_14563,N_14703);
nor U15107 (N_15107,N_14832,N_14687);
and U15108 (N_15108,N_14618,N_14591);
xor U15109 (N_15109,N_14945,N_14528);
or U15110 (N_15110,N_14695,N_14863);
nand U15111 (N_15111,N_14995,N_14742);
nor U15112 (N_15112,N_14710,N_14583);
nor U15113 (N_15113,N_14512,N_14678);
nor U15114 (N_15114,N_14786,N_14568);
and U15115 (N_15115,N_14531,N_14504);
nor U15116 (N_15116,N_14556,N_14759);
nor U15117 (N_15117,N_14997,N_14667);
nand U15118 (N_15118,N_14830,N_14652);
and U15119 (N_15119,N_14870,N_14564);
and U15120 (N_15120,N_14975,N_14956);
or U15121 (N_15121,N_14959,N_14803);
nor U15122 (N_15122,N_14605,N_14981);
or U15123 (N_15123,N_14743,N_14501);
nand U15124 (N_15124,N_14913,N_14955);
or U15125 (N_15125,N_14607,N_14821);
nand U15126 (N_15126,N_14852,N_14965);
and U15127 (N_15127,N_14712,N_14779);
and U15128 (N_15128,N_14825,N_14773);
nand U15129 (N_15129,N_14988,N_14537);
nand U15130 (N_15130,N_14845,N_14917);
nand U15131 (N_15131,N_14627,N_14735);
or U15132 (N_15132,N_14641,N_14517);
and U15133 (N_15133,N_14921,N_14931);
or U15134 (N_15134,N_14724,N_14543);
nor U15135 (N_15135,N_14559,N_14777);
nor U15136 (N_15136,N_14991,N_14817);
and U15137 (N_15137,N_14800,N_14887);
or U15138 (N_15138,N_14587,N_14653);
nand U15139 (N_15139,N_14620,N_14849);
and U15140 (N_15140,N_14998,N_14628);
and U15141 (N_15141,N_14508,N_14888);
or U15142 (N_15142,N_14813,N_14616);
nor U15143 (N_15143,N_14809,N_14633);
nor U15144 (N_15144,N_14947,N_14666);
or U15145 (N_15145,N_14739,N_14576);
or U15146 (N_15146,N_14971,N_14670);
or U15147 (N_15147,N_14862,N_14854);
and U15148 (N_15148,N_14951,N_14680);
or U15149 (N_15149,N_14804,N_14990);
or U15150 (N_15150,N_14582,N_14920);
and U15151 (N_15151,N_14770,N_14600);
nand U15152 (N_15152,N_14933,N_14500);
and U15153 (N_15153,N_14744,N_14542);
nor U15154 (N_15154,N_14725,N_14970);
nor U15155 (N_15155,N_14785,N_14902);
nand U15156 (N_15156,N_14967,N_14624);
nand U15157 (N_15157,N_14614,N_14794);
nand U15158 (N_15158,N_14899,N_14880);
and U15159 (N_15159,N_14848,N_14602);
and U15160 (N_15160,N_14932,N_14688);
xor U15161 (N_15161,N_14601,N_14768);
or U15162 (N_15162,N_14752,N_14696);
nor U15163 (N_15163,N_14806,N_14976);
or U15164 (N_15164,N_14736,N_14864);
and U15165 (N_15165,N_14615,N_14630);
nand U15166 (N_15166,N_14882,N_14575);
or U15167 (N_15167,N_14979,N_14798);
and U15168 (N_15168,N_14534,N_14761);
nand U15169 (N_15169,N_14571,N_14983);
nor U15170 (N_15170,N_14909,N_14612);
or U15171 (N_15171,N_14871,N_14636);
nor U15172 (N_15172,N_14664,N_14588);
nor U15173 (N_15173,N_14545,N_14767);
or U15174 (N_15174,N_14919,N_14881);
nor U15175 (N_15175,N_14572,N_14578);
and U15176 (N_15176,N_14836,N_14843);
and U15177 (N_15177,N_14824,N_14719);
nand U15178 (N_15178,N_14877,N_14891);
nor U15179 (N_15179,N_14639,N_14756);
nand U15180 (N_15180,N_14807,N_14720);
and U15181 (N_15181,N_14912,N_14604);
nor U15182 (N_15182,N_14992,N_14942);
nand U15183 (N_15183,N_14610,N_14634);
and U15184 (N_15184,N_14974,N_14775);
nand U15185 (N_15185,N_14613,N_14635);
and U15186 (N_15186,N_14715,N_14741);
nand U15187 (N_15187,N_14753,N_14505);
xnor U15188 (N_15188,N_14784,N_14603);
and U15189 (N_15189,N_14928,N_14693);
or U15190 (N_15190,N_14766,N_14629);
nand U15191 (N_15191,N_14790,N_14875);
nand U15192 (N_15192,N_14535,N_14823);
nand U15193 (N_15193,N_14908,N_14801);
or U15194 (N_15194,N_14780,N_14519);
and U15195 (N_15195,N_14993,N_14684);
or U15196 (N_15196,N_14958,N_14894);
or U15197 (N_15197,N_14781,N_14833);
nand U15198 (N_15198,N_14787,N_14755);
nor U15199 (N_15199,N_14826,N_14810);
or U15200 (N_15200,N_14654,N_14723);
and U15201 (N_15201,N_14700,N_14814);
and U15202 (N_15202,N_14595,N_14949);
nor U15203 (N_15203,N_14509,N_14960);
nor U15204 (N_15204,N_14554,N_14731);
and U15205 (N_15205,N_14996,N_14840);
or U15206 (N_15206,N_14764,N_14822);
and U15207 (N_15207,N_14906,N_14815);
or U15208 (N_15208,N_14570,N_14507);
or U15209 (N_15209,N_14846,N_14793);
or U15210 (N_15210,N_14918,N_14552);
nor U15211 (N_15211,N_14589,N_14939);
or U15212 (N_15212,N_14540,N_14954);
nand U15213 (N_15213,N_14566,N_14964);
nand U15214 (N_15214,N_14593,N_14506);
nand U15215 (N_15215,N_14763,N_14749);
or U15216 (N_15216,N_14511,N_14626);
nor U15217 (N_15217,N_14708,N_14977);
nand U15218 (N_15218,N_14580,N_14796);
nor U15219 (N_15219,N_14994,N_14621);
and U15220 (N_15220,N_14927,N_14972);
nor U15221 (N_15221,N_14683,N_14746);
nand U15222 (N_15222,N_14631,N_14514);
and U15223 (N_15223,N_14978,N_14674);
xnor U15224 (N_15224,N_14757,N_14668);
nor U15225 (N_15225,N_14522,N_14722);
and U15226 (N_15226,N_14762,N_14718);
nor U15227 (N_15227,N_14929,N_14816);
or U15228 (N_15228,N_14649,N_14916);
nor U15229 (N_15229,N_14590,N_14910);
nor U15230 (N_15230,N_14560,N_14669);
nor U15231 (N_15231,N_14671,N_14868);
nor U15232 (N_15232,N_14819,N_14973);
nor U15233 (N_15233,N_14952,N_14705);
and U15234 (N_15234,N_14536,N_14765);
nand U15235 (N_15235,N_14968,N_14585);
nand U15236 (N_15236,N_14937,N_14638);
and U15237 (N_15237,N_14957,N_14530);
nor U15238 (N_15238,N_14681,N_14999);
nand U15239 (N_15239,N_14692,N_14609);
nor U15240 (N_15240,N_14866,N_14574);
or U15241 (N_15241,N_14776,N_14797);
or U15242 (N_15242,N_14835,N_14711);
or U15243 (N_15243,N_14750,N_14873);
and U15244 (N_15244,N_14924,N_14599);
nor U15245 (N_15245,N_14510,N_14740);
nor U15246 (N_15246,N_14659,N_14844);
nand U15247 (N_15247,N_14709,N_14706);
nor U15248 (N_15248,N_14549,N_14533);
nand U15249 (N_15249,N_14783,N_14872);
xnor U15250 (N_15250,N_14876,N_14871);
or U15251 (N_15251,N_14574,N_14885);
or U15252 (N_15252,N_14552,N_14662);
or U15253 (N_15253,N_14776,N_14661);
nand U15254 (N_15254,N_14870,N_14733);
and U15255 (N_15255,N_14881,N_14543);
nor U15256 (N_15256,N_14552,N_14933);
nor U15257 (N_15257,N_14972,N_14622);
and U15258 (N_15258,N_14946,N_14597);
and U15259 (N_15259,N_14901,N_14991);
and U15260 (N_15260,N_14737,N_14708);
nand U15261 (N_15261,N_14627,N_14861);
or U15262 (N_15262,N_14786,N_14793);
nand U15263 (N_15263,N_14669,N_14951);
nor U15264 (N_15264,N_14741,N_14717);
and U15265 (N_15265,N_14836,N_14519);
and U15266 (N_15266,N_14585,N_14609);
nand U15267 (N_15267,N_14716,N_14507);
or U15268 (N_15268,N_14790,N_14739);
nor U15269 (N_15269,N_14952,N_14551);
nand U15270 (N_15270,N_14642,N_14976);
nor U15271 (N_15271,N_14500,N_14628);
nand U15272 (N_15272,N_14672,N_14578);
and U15273 (N_15273,N_14722,N_14832);
nand U15274 (N_15274,N_14779,N_14657);
and U15275 (N_15275,N_14576,N_14787);
and U15276 (N_15276,N_14636,N_14556);
nor U15277 (N_15277,N_14795,N_14658);
and U15278 (N_15278,N_14941,N_14513);
nand U15279 (N_15279,N_14689,N_14595);
nand U15280 (N_15280,N_14814,N_14627);
or U15281 (N_15281,N_14811,N_14539);
nand U15282 (N_15282,N_14808,N_14629);
or U15283 (N_15283,N_14802,N_14832);
or U15284 (N_15284,N_14790,N_14873);
nand U15285 (N_15285,N_14686,N_14769);
and U15286 (N_15286,N_14846,N_14892);
or U15287 (N_15287,N_14895,N_14968);
and U15288 (N_15288,N_14592,N_14856);
or U15289 (N_15289,N_14750,N_14638);
or U15290 (N_15290,N_14927,N_14568);
and U15291 (N_15291,N_14920,N_14880);
and U15292 (N_15292,N_14876,N_14822);
or U15293 (N_15293,N_14987,N_14792);
nor U15294 (N_15294,N_14685,N_14681);
nor U15295 (N_15295,N_14939,N_14744);
and U15296 (N_15296,N_14861,N_14872);
and U15297 (N_15297,N_14612,N_14986);
nor U15298 (N_15298,N_14877,N_14523);
and U15299 (N_15299,N_14796,N_14998);
nand U15300 (N_15300,N_14761,N_14986);
nand U15301 (N_15301,N_14596,N_14993);
nor U15302 (N_15302,N_14963,N_14914);
or U15303 (N_15303,N_14594,N_14686);
and U15304 (N_15304,N_14551,N_14702);
and U15305 (N_15305,N_14828,N_14834);
nor U15306 (N_15306,N_14949,N_14600);
nor U15307 (N_15307,N_14978,N_14639);
and U15308 (N_15308,N_14651,N_14894);
or U15309 (N_15309,N_14568,N_14645);
and U15310 (N_15310,N_14608,N_14615);
nand U15311 (N_15311,N_14604,N_14986);
or U15312 (N_15312,N_14965,N_14627);
nor U15313 (N_15313,N_14509,N_14693);
nand U15314 (N_15314,N_14521,N_14639);
nand U15315 (N_15315,N_14727,N_14875);
nand U15316 (N_15316,N_14956,N_14938);
nor U15317 (N_15317,N_14521,N_14598);
nor U15318 (N_15318,N_14515,N_14863);
or U15319 (N_15319,N_14962,N_14639);
nand U15320 (N_15320,N_14751,N_14774);
nor U15321 (N_15321,N_14546,N_14962);
or U15322 (N_15322,N_14829,N_14783);
and U15323 (N_15323,N_14732,N_14606);
nand U15324 (N_15324,N_14587,N_14632);
or U15325 (N_15325,N_14668,N_14901);
or U15326 (N_15326,N_14511,N_14706);
and U15327 (N_15327,N_14672,N_14658);
or U15328 (N_15328,N_14787,N_14901);
nand U15329 (N_15329,N_14916,N_14904);
nor U15330 (N_15330,N_14556,N_14659);
or U15331 (N_15331,N_14701,N_14980);
nand U15332 (N_15332,N_14687,N_14673);
or U15333 (N_15333,N_14718,N_14629);
nor U15334 (N_15334,N_14963,N_14918);
nand U15335 (N_15335,N_14940,N_14801);
or U15336 (N_15336,N_14846,N_14624);
nor U15337 (N_15337,N_14806,N_14801);
or U15338 (N_15338,N_14899,N_14547);
and U15339 (N_15339,N_14622,N_14891);
or U15340 (N_15340,N_14637,N_14935);
nand U15341 (N_15341,N_14706,N_14605);
nor U15342 (N_15342,N_14785,N_14582);
or U15343 (N_15343,N_14848,N_14716);
xor U15344 (N_15344,N_14581,N_14573);
or U15345 (N_15345,N_14717,N_14645);
nor U15346 (N_15346,N_14518,N_14913);
and U15347 (N_15347,N_14695,N_14813);
and U15348 (N_15348,N_14996,N_14506);
nor U15349 (N_15349,N_14723,N_14823);
and U15350 (N_15350,N_14711,N_14912);
or U15351 (N_15351,N_14545,N_14601);
nand U15352 (N_15352,N_14596,N_14527);
nand U15353 (N_15353,N_14568,N_14854);
nor U15354 (N_15354,N_14862,N_14896);
xor U15355 (N_15355,N_14752,N_14600);
and U15356 (N_15356,N_14520,N_14521);
nand U15357 (N_15357,N_14662,N_14847);
nand U15358 (N_15358,N_14876,N_14712);
xor U15359 (N_15359,N_14710,N_14998);
or U15360 (N_15360,N_14592,N_14576);
and U15361 (N_15361,N_14993,N_14869);
nor U15362 (N_15362,N_14536,N_14757);
nor U15363 (N_15363,N_14575,N_14557);
nor U15364 (N_15364,N_14706,N_14769);
nor U15365 (N_15365,N_14800,N_14990);
and U15366 (N_15366,N_14982,N_14636);
nor U15367 (N_15367,N_14685,N_14717);
and U15368 (N_15368,N_14916,N_14671);
and U15369 (N_15369,N_14671,N_14835);
nand U15370 (N_15370,N_14987,N_14964);
nand U15371 (N_15371,N_14955,N_14603);
and U15372 (N_15372,N_14730,N_14862);
or U15373 (N_15373,N_14974,N_14982);
nor U15374 (N_15374,N_14525,N_14940);
nand U15375 (N_15375,N_14738,N_14833);
or U15376 (N_15376,N_14702,N_14757);
nand U15377 (N_15377,N_14978,N_14810);
or U15378 (N_15378,N_14987,N_14531);
or U15379 (N_15379,N_14754,N_14925);
nor U15380 (N_15380,N_14674,N_14501);
or U15381 (N_15381,N_14690,N_14897);
or U15382 (N_15382,N_14513,N_14989);
or U15383 (N_15383,N_14634,N_14975);
and U15384 (N_15384,N_14785,N_14587);
and U15385 (N_15385,N_14862,N_14938);
nor U15386 (N_15386,N_14969,N_14856);
and U15387 (N_15387,N_14880,N_14538);
or U15388 (N_15388,N_14965,N_14666);
or U15389 (N_15389,N_14656,N_14585);
or U15390 (N_15390,N_14946,N_14716);
nor U15391 (N_15391,N_14718,N_14907);
nor U15392 (N_15392,N_14974,N_14598);
and U15393 (N_15393,N_14657,N_14887);
nand U15394 (N_15394,N_14793,N_14767);
nand U15395 (N_15395,N_14663,N_14835);
nand U15396 (N_15396,N_14856,N_14842);
and U15397 (N_15397,N_14788,N_14731);
xor U15398 (N_15398,N_14851,N_14854);
nand U15399 (N_15399,N_14692,N_14620);
nand U15400 (N_15400,N_14996,N_14782);
or U15401 (N_15401,N_14583,N_14715);
and U15402 (N_15402,N_14781,N_14622);
nor U15403 (N_15403,N_14717,N_14727);
nand U15404 (N_15404,N_14745,N_14685);
or U15405 (N_15405,N_14920,N_14777);
and U15406 (N_15406,N_14605,N_14546);
nand U15407 (N_15407,N_14860,N_14833);
and U15408 (N_15408,N_14805,N_14969);
nand U15409 (N_15409,N_14516,N_14751);
nand U15410 (N_15410,N_14790,N_14709);
and U15411 (N_15411,N_14980,N_14782);
nand U15412 (N_15412,N_14989,N_14583);
and U15413 (N_15413,N_14581,N_14961);
or U15414 (N_15414,N_14769,N_14791);
nand U15415 (N_15415,N_14769,N_14799);
or U15416 (N_15416,N_14882,N_14650);
nor U15417 (N_15417,N_14701,N_14916);
and U15418 (N_15418,N_14885,N_14962);
and U15419 (N_15419,N_14595,N_14713);
or U15420 (N_15420,N_14665,N_14553);
or U15421 (N_15421,N_14646,N_14803);
nor U15422 (N_15422,N_14948,N_14655);
nand U15423 (N_15423,N_14698,N_14734);
and U15424 (N_15424,N_14545,N_14636);
or U15425 (N_15425,N_14643,N_14505);
nand U15426 (N_15426,N_14780,N_14745);
nor U15427 (N_15427,N_14701,N_14542);
and U15428 (N_15428,N_14651,N_14897);
nor U15429 (N_15429,N_14559,N_14731);
or U15430 (N_15430,N_14585,N_14710);
or U15431 (N_15431,N_14727,N_14858);
nor U15432 (N_15432,N_14567,N_14620);
nand U15433 (N_15433,N_14811,N_14739);
nor U15434 (N_15434,N_14805,N_14900);
or U15435 (N_15435,N_14923,N_14738);
and U15436 (N_15436,N_14619,N_14921);
and U15437 (N_15437,N_14837,N_14680);
and U15438 (N_15438,N_14525,N_14762);
xnor U15439 (N_15439,N_14825,N_14859);
nand U15440 (N_15440,N_14840,N_14843);
nor U15441 (N_15441,N_14645,N_14779);
nand U15442 (N_15442,N_14871,N_14544);
nand U15443 (N_15443,N_14590,N_14759);
or U15444 (N_15444,N_14871,N_14951);
nor U15445 (N_15445,N_14692,N_14954);
or U15446 (N_15446,N_14537,N_14663);
or U15447 (N_15447,N_14549,N_14532);
and U15448 (N_15448,N_14660,N_14863);
xor U15449 (N_15449,N_14727,N_14767);
nor U15450 (N_15450,N_14944,N_14870);
or U15451 (N_15451,N_14784,N_14808);
nand U15452 (N_15452,N_14666,N_14773);
nand U15453 (N_15453,N_14852,N_14502);
and U15454 (N_15454,N_14693,N_14862);
nand U15455 (N_15455,N_14730,N_14671);
nor U15456 (N_15456,N_14917,N_14557);
or U15457 (N_15457,N_14543,N_14621);
or U15458 (N_15458,N_14599,N_14764);
or U15459 (N_15459,N_14956,N_14691);
nor U15460 (N_15460,N_14791,N_14708);
and U15461 (N_15461,N_14904,N_14841);
or U15462 (N_15462,N_14715,N_14835);
nand U15463 (N_15463,N_14857,N_14676);
nand U15464 (N_15464,N_14771,N_14963);
or U15465 (N_15465,N_14795,N_14922);
nand U15466 (N_15466,N_14697,N_14651);
nor U15467 (N_15467,N_14772,N_14633);
and U15468 (N_15468,N_14902,N_14876);
or U15469 (N_15469,N_14510,N_14831);
and U15470 (N_15470,N_14522,N_14854);
or U15471 (N_15471,N_14683,N_14756);
or U15472 (N_15472,N_14733,N_14512);
and U15473 (N_15473,N_14952,N_14997);
nand U15474 (N_15474,N_14751,N_14841);
nor U15475 (N_15475,N_14934,N_14757);
nand U15476 (N_15476,N_14987,N_14881);
and U15477 (N_15477,N_14594,N_14654);
nor U15478 (N_15478,N_14794,N_14870);
nor U15479 (N_15479,N_14978,N_14969);
nand U15480 (N_15480,N_14575,N_14598);
or U15481 (N_15481,N_14986,N_14773);
nor U15482 (N_15482,N_14594,N_14897);
xnor U15483 (N_15483,N_14995,N_14577);
or U15484 (N_15484,N_14672,N_14789);
xnor U15485 (N_15485,N_14544,N_14810);
and U15486 (N_15486,N_14615,N_14809);
xor U15487 (N_15487,N_14682,N_14749);
or U15488 (N_15488,N_14890,N_14766);
nor U15489 (N_15489,N_14517,N_14870);
nand U15490 (N_15490,N_14689,N_14708);
and U15491 (N_15491,N_14781,N_14948);
and U15492 (N_15492,N_14514,N_14726);
and U15493 (N_15493,N_14827,N_14906);
nand U15494 (N_15494,N_14563,N_14859);
and U15495 (N_15495,N_14928,N_14545);
or U15496 (N_15496,N_14642,N_14921);
and U15497 (N_15497,N_14939,N_14737);
xnor U15498 (N_15498,N_14615,N_14861);
and U15499 (N_15499,N_14594,N_14889);
and U15500 (N_15500,N_15484,N_15225);
nand U15501 (N_15501,N_15442,N_15354);
nand U15502 (N_15502,N_15104,N_15251);
nor U15503 (N_15503,N_15388,N_15202);
and U15504 (N_15504,N_15499,N_15065);
and U15505 (N_15505,N_15491,N_15019);
xnor U15506 (N_15506,N_15493,N_15322);
nor U15507 (N_15507,N_15003,N_15471);
or U15508 (N_15508,N_15261,N_15037);
nand U15509 (N_15509,N_15283,N_15011);
nor U15510 (N_15510,N_15004,N_15394);
or U15511 (N_15511,N_15460,N_15205);
nand U15512 (N_15512,N_15178,N_15403);
or U15513 (N_15513,N_15463,N_15103);
nor U15514 (N_15514,N_15142,N_15120);
nor U15515 (N_15515,N_15296,N_15404);
and U15516 (N_15516,N_15305,N_15468);
and U15517 (N_15517,N_15073,N_15113);
xor U15518 (N_15518,N_15370,N_15076);
nand U15519 (N_15519,N_15380,N_15030);
nand U15520 (N_15520,N_15222,N_15413);
nor U15521 (N_15521,N_15208,N_15436);
nor U15522 (N_15522,N_15349,N_15236);
nand U15523 (N_15523,N_15284,N_15034);
nor U15524 (N_15524,N_15280,N_15395);
or U15525 (N_15525,N_15494,N_15143);
or U15526 (N_15526,N_15425,N_15459);
nor U15527 (N_15527,N_15376,N_15072);
and U15528 (N_15528,N_15458,N_15195);
xor U15529 (N_15529,N_15124,N_15247);
nor U15530 (N_15530,N_15488,N_15125);
xnor U15531 (N_15531,N_15316,N_15387);
nor U15532 (N_15532,N_15415,N_15430);
nand U15533 (N_15533,N_15188,N_15258);
and U15534 (N_15534,N_15437,N_15221);
nor U15535 (N_15535,N_15432,N_15393);
or U15536 (N_15536,N_15276,N_15181);
and U15537 (N_15537,N_15097,N_15472);
and U15538 (N_15538,N_15228,N_15277);
nand U15539 (N_15539,N_15074,N_15197);
or U15540 (N_15540,N_15264,N_15287);
or U15541 (N_15541,N_15153,N_15420);
nor U15542 (N_15542,N_15151,N_15235);
nand U15543 (N_15543,N_15344,N_15162);
and U15544 (N_15544,N_15043,N_15330);
and U15545 (N_15545,N_15165,N_15269);
or U15546 (N_15546,N_15428,N_15058);
nand U15547 (N_15547,N_15050,N_15313);
nand U15548 (N_15548,N_15026,N_15010);
or U15549 (N_15549,N_15231,N_15408);
nand U15550 (N_15550,N_15136,N_15441);
xnor U15551 (N_15551,N_15377,N_15273);
nor U15552 (N_15552,N_15489,N_15244);
and U15553 (N_15553,N_15379,N_15454);
nor U15554 (N_15554,N_15137,N_15149);
nor U15555 (N_15555,N_15014,N_15071);
or U15556 (N_15556,N_15315,N_15041);
xor U15557 (N_15557,N_15170,N_15200);
and U15558 (N_15558,N_15084,N_15046);
nand U15559 (N_15559,N_15443,N_15422);
or U15560 (N_15560,N_15374,N_15333);
nand U15561 (N_15561,N_15444,N_15232);
or U15562 (N_15562,N_15497,N_15135);
nand U15563 (N_15563,N_15433,N_15411);
and U15564 (N_15564,N_15020,N_15075);
or U15565 (N_15565,N_15006,N_15007);
or U15566 (N_15566,N_15255,N_15173);
or U15567 (N_15567,N_15320,N_15217);
xor U15568 (N_15568,N_15310,N_15329);
nor U15569 (N_15569,N_15187,N_15111);
nand U15570 (N_15570,N_15319,N_15015);
and U15571 (N_15571,N_15029,N_15048);
nor U15572 (N_15572,N_15201,N_15271);
nand U15573 (N_15573,N_15345,N_15331);
or U15574 (N_15574,N_15378,N_15101);
nand U15575 (N_15575,N_15138,N_15160);
or U15576 (N_15576,N_15241,N_15355);
nand U15577 (N_15577,N_15382,N_15177);
nor U15578 (N_15578,N_15438,N_15230);
or U15579 (N_15579,N_15154,N_15148);
nor U15580 (N_15580,N_15086,N_15397);
nor U15581 (N_15581,N_15309,N_15409);
and U15582 (N_15582,N_15040,N_15326);
nor U15583 (N_15583,N_15146,N_15233);
or U15584 (N_15584,N_15418,N_15018);
or U15585 (N_15585,N_15121,N_15439);
nand U15586 (N_15586,N_15293,N_15013);
or U15587 (N_15587,N_15301,N_15461);
nor U15588 (N_15588,N_15448,N_15304);
or U15589 (N_15589,N_15297,N_15130);
or U15590 (N_15590,N_15424,N_15412);
and U15591 (N_15591,N_15134,N_15179);
nor U15592 (N_15592,N_15279,N_15226);
or U15593 (N_15593,N_15328,N_15381);
nand U15594 (N_15594,N_15465,N_15352);
and U15595 (N_15595,N_15335,N_15294);
and U15596 (N_15596,N_15431,N_15435);
nand U15597 (N_15597,N_15174,N_15254);
nand U15598 (N_15598,N_15051,N_15194);
nand U15599 (N_15599,N_15350,N_15105);
and U15600 (N_15600,N_15373,N_15429);
nor U15601 (N_15601,N_15317,N_15008);
or U15602 (N_15602,N_15166,N_15371);
nand U15603 (N_15603,N_15383,N_15392);
and U15604 (N_15604,N_15060,N_15203);
nand U15605 (N_15605,N_15385,N_15238);
or U15606 (N_15606,N_15475,N_15325);
and U15607 (N_15607,N_15139,N_15152);
and U15608 (N_15608,N_15110,N_15298);
nor U15609 (N_15609,N_15286,N_15089);
and U15610 (N_15610,N_15260,N_15155);
or U15611 (N_15611,N_15082,N_15033);
nor U15612 (N_15612,N_15240,N_15314);
or U15613 (N_15613,N_15126,N_15064);
and U15614 (N_15614,N_15311,N_15038);
nor U15615 (N_15615,N_15398,N_15306);
or U15616 (N_15616,N_15281,N_15133);
and U15617 (N_15617,N_15342,N_15009);
and U15618 (N_15618,N_15036,N_15172);
or U15619 (N_15619,N_15481,N_15114);
nor U15620 (N_15620,N_15396,N_15066);
or U15621 (N_15621,N_15140,N_15289);
or U15622 (N_15622,N_15272,N_15318);
or U15623 (N_15623,N_15375,N_15427);
or U15624 (N_15624,N_15183,N_15091);
xnor U15625 (N_15625,N_15312,N_15469);
and U15626 (N_15626,N_15421,N_15423);
and U15627 (N_15627,N_15122,N_15163);
nand U15628 (N_15628,N_15372,N_15031);
nor U15629 (N_15629,N_15452,N_15078);
or U15630 (N_15630,N_15099,N_15270);
and U15631 (N_15631,N_15478,N_15157);
and U15632 (N_15632,N_15016,N_15213);
nand U15633 (N_15633,N_15303,N_15467);
xnor U15634 (N_15634,N_15250,N_15159);
nor U15635 (N_15635,N_15035,N_15485);
nand U15636 (N_15636,N_15132,N_15257);
or U15637 (N_15637,N_15189,N_15062);
nor U15638 (N_15638,N_15324,N_15219);
and U15639 (N_15639,N_15131,N_15307);
nor U15640 (N_15640,N_15256,N_15025);
xnor U15641 (N_15641,N_15285,N_15184);
and U15642 (N_15642,N_15449,N_15211);
nor U15643 (N_15643,N_15477,N_15480);
nand U15644 (N_15644,N_15268,N_15321);
and U15645 (N_15645,N_15115,N_15399);
and U15646 (N_15646,N_15087,N_15360);
or U15647 (N_15647,N_15106,N_15447);
nand U15648 (N_15648,N_15128,N_15168);
and U15649 (N_15649,N_15190,N_15340);
or U15650 (N_15650,N_15061,N_15021);
nand U15651 (N_15651,N_15186,N_15220);
or U15652 (N_15652,N_15407,N_15118);
nand U15653 (N_15653,N_15196,N_15248);
nand U15654 (N_15654,N_15470,N_15414);
nor U15655 (N_15655,N_15042,N_15039);
and U15656 (N_15656,N_15457,N_15098);
nor U15657 (N_15657,N_15391,N_15364);
nand U15658 (N_15658,N_15056,N_15492);
nor U15659 (N_15659,N_15332,N_15292);
nor U15660 (N_15660,N_15299,N_15486);
and U15661 (N_15661,N_15339,N_15107);
and U15662 (N_15662,N_15147,N_15027);
or U15663 (N_15663,N_15327,N_15450);
or U15664 (N_15664,N_15367,N_15145);
nor U15665 (N_15665,N_15265,N_15227);
nand U15666 (N_15666,N_15047,N_15001);
nand U15667 (N_15667,N_15094,N_15192);
and U15668 (N_15668,N_15384,N_15090);
or U15669 (N_15669,N_15479,N_15077);
or U15670 (N_15670,N_15070,N_15063);
and U15671 (N_15671,N_15356,N_15055);
nor U15672 (N_15672,N_15237,N_15456);
nor U15673 (N_15673,N_15109,N_15229);
or U15674 (N_15674,N_15095,N_15363);
and U15675 (N_15675,N_15338,N_15275);
or U15676 (N_15676,N_15290,N_15167);
or U15677 (N_15677,N_15405,N_15182);
and U15678 (N_15678,N_15215,N_15218);
and U15679 (N_15679,N_15081,N_15127);
and U15680 (N_15680,N_15348,N_15359);
nor U15681 (N_15681,N_15417,N_15259);
nand U15682 (N_15682,N_15053,N_15185);
nor U15683 (N_15683,N_15093,N_15453);
xor U15684 (N_15684,N_15473,N_15161);
nand U15685 (N_15685,N_15171,N_15028);
or U15686 (N_15686,N_15052,N_15193);
and U15687 (N_15687,N_15141,N_15401);
or U15688 (N_15688,N_15012,N_15206);
nor U15689 (N_15689,N_15302,N_15362);
nor U15690 (N_15690,N_15239,N_15024);
nand U15691 (N_15691,N_15390,N_15117);
nand U15692 (N_15692,N_15234,N_15365);
nand U15693 (N_15693,N_15446,N_15323);
and U15694 (N_15694,N_15180,N_15005);
nand U15695 (N_15695,N_15358,N_15069);
nor U15696 (N_15696,N_15341,N_15156);
and U15697 (N_15697,N_15088,N_15266);
nand U15698 (N_15698,N_15245,N_15368);
nand U15699 (N_15699,N_15123,N_15083);
xor U15700 (N_15700,N_15002,N_15386);
and U15701 (N_15701,N_15022,N_15000);
nand U15702 (N_15702,N_15402,N_15487);
or U15703 (N_15703,N_15267,N_15476);
nand U15704 (N_15704,N_15426,N_15212);
nand U15705 (N_15705,N_15464,N_15278);
nand U15706 (N_15706,N_15490,N_15274);
or U15707 (N_15707,N_15351,N_15210);
nor U15708 (N_15708,N_15334,N_15249);
and U15709 (N_15709,N_15346,N_15445);
nand U15710 (N_15710,N_15482,N_15455);
nand U15711 (N_15711,N_15389,N_15410);
or U15712 (N_15712,N_15353,N_15288);
and U15713 (N_15713,N_15451,N_15300);
nand U15714 (N_15714,N_15116,N_15291);
nand U15715 (N_15715,N_15295,N_15357);
nor U15716 (N_15716,N_15252,N_15242);
nand U15717 (N_15717,N_15045,N_15400);
nand U15718 (N_15718,N_15336,N_15308);
or U15719 (N_15719,N_15096,N_15102);
nand U15720 (N_15720,N_15158,N_15495);
nor U15721 (N_15721,N_15017,N_15207);
nand U15722 (N_15722,N_15059,N_15496);
nor U15723 (N_15723,N_15092,N_15068);
nand U15724 (N_15724,N_15150,N_15049);
and U15725 (N_15725,N_15243,N_15204);
nor U15726 (N_15726,N_15085,N_15246);
or U15727 (N_15727,N_15366,N_15369);
nor U15728 (N_15728,N_15209,N_15112);
nand U15729 (N_15729,N_15044,N_15067);
and U15730 (N_15730,N_15483,N_15253);
nor U15731 (N_15731,N_15199,N_15080);
and U15732 (N_15732,N_15119,N_15169);
nand U15733 (N_15733,N_15224,N_15100);
or U15734 (N_15734,N_15191,N_15032);
and U15735 (N_15735,N_15108,N_15198);
and U15736 (N_15736,N_15223,N_15347);
nor U15737 (N_15737,N_15023,N_15343);
nand U15738 (N_15738,N_15434,N_15263);
nor U15739 (N_15739,N_15164,N_15419);
xnor U15740 (N_15740,N_15498,N_15214);
nand U15741 (N_15741,N_15262,N_15361);
and U15742 (N_15742,N_15175,N_15406);
and U15743 (N_15743,N_15176,N_15054);
nor U15744 (N_15744,N_15474,N_15466);
nor U15745 (N_15745,N_15057,N_15144);
or U15746 (N_15746,N_15337,N_15216);
nor U15747 (N_15747,N_15079,N_15462);
and U15748 (N_15748,N_15440,N_15129);
and U15749 (N_15749,N_15282,N_15416);
or U15750 (N_15750,N_15474,N_15457);
or U15751 (N_15751,N_15166,N_15016);
nand U15752 (N_15752,N_15158,N_15303);
nor U15753 (N_15753,N_15218,N_15291);
or U15754 (N_15754,N_15333,N_15034);
nor U15755 (N_15755,N_15089,N_15013);
and U15756 (N_15756,N_15212,N_15086);
and U15757 (N_15757,N_15410,N_15328);
or U15758 (N_15758,N_15083,N_15480);
nand U15759 (N_15759,N_15359,N_15284);
and U15760 (N_15760,N_15125,N_15222);
and U15761 (N_15761,N_15451,N_15058);
nand U15762 (N_15762,N_15468,N_15050);
and U15763 (N_15763,N_15096,N_15024);
or U15764 (N_15764,N_15432,N_15451);
nand U15765 (N_15765,N_15481,N_15259);
nor U15766 (N_15766,N_15376,N_15409);
or U15767 (N_15767,N_15283,N_15431);
nor U15768 (N_15768,N_15194,N_15416);
or U15769 (N_15769,N_15310,N_15403);
or U15770 (N_15770,N_15267,N_15135);
and U15771 (N_15771,N_15249,N_15188);
nand U15772 (N_15772,N_15388,N_15411);
nor U15773 (N_15773,N_15438,N_15492);
nor U15774 (N_15774,N_15319,N_15048);
nor U15775 (N_15775,N_15440,N_15127);
or U15776 (N_15776,N_15301,N_15494);
nand U15777 (N_15777,N_15262,N_15339);
and U15778 (N_15778,N_15342,N_15169);
or U15779 (N_15779,N_15424,N_15346);
and U15780 (N_15780,N_15477,N_15474);
nor U15781 (N_15781,N_15022,N_15194);
or U15782 (N_15782,N_15269,N_15169);
or U15783 (N_15783,N_15283,N_15416);
and U15784 (N_15784,N_15417,N_15297);
or U15785 (N_15785,N_15373,N_15327);
nand U15786 (N_15786,N_15459,N_15305);
and U15787 (N_15787,N_15452,N_15107);
nand U15788 (N_15788,N_15056,N_15489);
nand U15789 (N_15789,N_15333,N_15384);
and U15790 (N_15790,N_15182,N_15378);
nor U15791 (N_15791,N_15322,N_15240);
nand U15792 (N_15792,N_15205,N_15307);
nor U15793 (N_15793,N_15268,N_15428);
or U15794 (N_15794,N_15063,N_15173);
nor U15795 (N_15795,N_15068,N_15365);
or U15796 (N_15796,N_15452,N_15317);
or U15797 (N_15797,N_15138,N_15016);
and U15798 (N_15798,N_15063,N_15119);
nand U15799 (N_15799,N_15274,N_15115);
or U15800 (N_15800,N_15131,N_15366);
nand U15801 (N_15801,N_15454,N_15120);
and U15802 (N_15802,N_15303,N_15094);
or U15803 (N_15803,N_15383,N_15265);
nand U15804 (N_15804,N_15031,N_15352);
and U15805 (N_15805,N_15271,N_15146);
nor U15806 (N_15806,N_15054,N_15470);
and U15807 (N_15807,N_15029,N_15471);
nand U15808 (N_15808,N_15132,N_15110);
nor U15809 (N_15809,N_15046,N_15391);
or U15810 (N_15810,N_15416,N_15392);
or U15811 (N_15811,N_15039,N_15453);
nand U15812 (N_15812,N_15218,N_15010);
nor U15813 (N_15813,N_15401,N_15244);
and U15814 (N_15814,N_15163,N_15154);
or U15815 (N_15815,N_15141,N_15402);
or U15816 (N_15816,N_15424,N_15454);
nand U15817 (N_15817,N_15163,N_15260);
nor U15818 (N_15818,N_15026,N_15054);
xnor U15819 (N_15819,N_15200,N_15378);
nand U15820 (N_15820,N_15116,N_15412);
or U15821 (N_15821,N_15047,N_15164);
or U15822 (N_15822,N_15195,N_15381);
nand U15823 (N_15823,N_15130,N_15306);
or U15824 (N_15824,N_15025,N_15337);
and U15825 (N_15825,N_15313,N_15448);
nor U15826 (N_15826,N_15299,N_15414);
nand U15827 (N_15827,N_15033,N_15158);
nand U15828 (N_15828,N_15149,N_15153);
or U15829 (N_15829,N_15101,N_15480);
or U15830 (N_15830,N_15037,N_15336);
nand U15831 (N_15831,N_15199,N_15064);
nand U15832 (N_15832,N_15483,N_15426);
nand U15833 (N_15833,N_15477,N_15347);
nor U15834 (N_15834,N_15332,N_15019);
or U15835 (N_15835,N_15093,N_15413);
or U15836 (N_15836,N_15454,N_15014);
or U15837 (N_15837,N_15476,N_15208);
xnor U15838 (N_15838,N_15025,N_15052);
or U15839 (N_15839,N_15003,N_15342);
xnor U15840 (N_15840,N_15427,N_15048);
and U15841 (N_15841,N_15376,N_15135);
or U15842 (N_15842,N_15205,N_15399);
nand U15843 (N_15843,N_15455,N_15302);
or U15844 (N_15844,N_15441,N_15182);
and U15845 (N_15845,N_15097,N_15117);
or U15846 (N_15846,N_15109,N_15035);
nor U15847 (N_15847,N_15054,N_15286);
nand U15848 (N_15848,N_15480,N_15461);
and U15849 (N_15849,N_15079,N_15235);
nand U15850 (N_15850,N_15063,N_15107);
xor U15851 (N_15851,N_15411,N_15410);
and U15852 (N_15852,N_15369,N_15359);
nor U15853 (N_15853,N_15074,N_15105);
nor U15854 (N_15854,N_15359,N_15102);
nor U15855 (N_15855,N_15434,N_15224);
nand U15856 (N_15856,N_15066,N_15432);
nor U15857 (N_15857,N_15301,N_15264);
nor U15858 (N_15858,N_15360,N_15081);
or U15859 (N_15859,N_15448,N_15339);
and U15860 (N_15860,N_15442,N_15240);
nand U15861 (N_15861,N_15184,N_15176);
or U15862 (N_15862,N_15187,N_15247);
or U15863 (N_15863,N_15327,N_15046);
or U15864 (N_15864,N_15444,N_15144);
or U15865 (N_15865,N_15276,N_15258);
or U15866 (N_15866,N_15027,N_15105);
or U15867 (N_15867,N_15107,N_15054);
or U15868 (N_15868,N_15108,N_15178);
or U15869 (N_15869,N_15493,N_15407);
and U15870 (N_15870,N_15024,N_15165);
and U15871 (N_15871,N_15120,N_15395);
nand U15872 (N_15872,N_15206,N_15020);
nand U15873 (N_15873,N_15137,N_15160);
nor U15874 (N_15874,N_15153,N_15209);
nor U15875 (N_15875,N_15104,N_15387);
and U15876 (N_15876,N_15044,N_15297);
and U15877 (N_15877,N_15282,N_15345);
and U15878 (N_15878,N_15208,N_15487);
or U15879 (N_15879,N_15290,N_15346);
nand U15880 (N_15880,N_15008,N_15197);
and U15881 (N_15881,N_15150,N_15151);
nor U15882 (N_15882,N_15429,N_15194);
or U15883 (N_15883,N_15342,N_15263);
and U15884 (N_15884,N_15317,N_15208);
nor U15885 (N_15885,N_15457,N_15200);
or U15886 (N_15886,N_15149,N_15476);
nand U15887 (N_15887,N_15034,N_15110);
or U15888 (N_15888,N_15221,N_15083);
nand U15889 (N_15889,N_15205,N_15365);
or U15890 (N_15890,N_15415,N_15309);
and U15891 (N_15891,N_15174,N_15173);
and U15892 (N_15892,N_15101,N_15177);
nand U15893 (N_15893,N_15417,N_15263);
or U15894 (N_15894,N_15488,N_15183);
or U15895 (N_15895,N_15041,N_15425);
or U15896 (N_15896,N_15176,N_15470);
nor U15897 (N_15897,N_15177,N_15453);
nand U15898 (N_15898,N_15370,N_15309);
and U15899 (N_15899,N_15336,N_15278);
nand U15900 (N_15900,N_15191,N_15178);
nand U15901 (N_15901,N_15183,N_15346);
nand U15902 (N_15902,N_15075,N_15190);
nand U15903 (N_15903,N_15102,N_15339);
or U15904 (N_15904,N_15411,N_15114);
and U15905 (N_15905,N_15222,N_15096);
and U15906 (N_15906,N_15292,N_15477);
or U15907 (N_15907,N_15451,N_15346);
nor U15908 (N_15908,N_15034,N_15328);
and U15909 (N_15909,N_15046,N_15086);
or U15910 (N_15910,N_15438,N_15327);
and U15911 (N_15911,N_15431,N_15109);
nand U15912 (N_15912,N_15139,N_15484);
xor U15913 (N_15913,N_15331,N_15073);
and U15914 (N_15914,N_15382,N_15227);
or U15915 (N_15915,N_15336,N_15161);
and U15916 (N_15916,N_15228,N_15410);
nor U15917 (N_15917,N_15010,N_15496);
nand U15918 (N_15918,N_15044,N_15390);
and U15919 (N_15919,N_15212,N_15120);
or U15920 (N_15920,N_15066,N_15000);
nor U15921 (N_15921,N_15041,N_15038);
nand U15922 (N_15922,N_15425,N_15345);
and U15923 (N_15923,N_15027,N_15349);
or U15924 (N_15924,N_15407,N_15497);
nand U15925 (N_15925,N_15236,N_15068);
nand U15926 (N_15926,N_15109,N_15070);
or U15927 (N_15927,N_15011,N_15114);
nor U15928 (N_15928,N_15384,N_15211);
and U15929 (N_15929,N_15090,N_15428);
or U15930 (N_15930,N_15154,N_15174);
nor U15931 (N_15931,N_15385,N_15156);
xnor U15932 (N_15932,N_15251,N_15336);
nor U15933 (N_15933,N_15331,N_15342);
or U15934 (N_15934,N_15170,N_15291);
and U15935 (N_15935,N_15112,N_15407);
and U15936 (N_15936,N_15354,N_15286);
and U15937 (N_15937,N_15089,N_15301);
nor U15938 (N_15938,N_15262,N_15234);
nor U15939 (N_15939,N_15266,N_15015);
nand U15940 (N_15940,N_15161,N_15067);
and U15941 (N_15941,N_15467,N_15022);
nand U15942 (N_15942,N_15248,N_15359);
and U15943 (N_15943,N_15048,N_15106);
nand U15944 (N_15944,N_15303,N_15401);
nand U15945 (N_15945,N_15381,N_15145);
xnor U15946 (N_15946,N_15031,N_15435);
nor U15947 (N_15947,N_15036,N_15063);
nand U15948 (N_15948,N_15136,N_15283);
nand U15949 (N_15949,N_15322,N_15049);
nor U15950 (N_15950,N_15048,N_15450);
nand U15951 (N_15951,N_15430,N_15088);
or U15952 (N_15952,N_15146,N_15336);
or U15953 (N_15953,N_15240,N_15470);
nor U15954 (N_15954,N_15422,N_15404);
and U15955 (N_15955,N_15380,N_15070);
nand U15956 (N_15956,N_15242,N_15400);
nand U15957 (N_15957,N_15483,N_15131);
xnor U15958 (N_15958,N_15474,N_15482);
and U15959 (N_15959,N_15382,N_15461);
nor U15960 (N_15960,N_15158,N_15227);
or U15961 (N_15961,N_15298,N_15369);
nor U15962 (N_15962,N_15054,N_15042);
nor U15963 (N_15963,N_15118,N_15347);
nor U15964 (N_15964,N_15021,N_15189);
or U15965 (N_15965,N_15294,N_15263);
or U15966 (N_15966,N_15497,N_15386);
and U15967 (N_15967,N_15155,N_15420);
nand U15968 (N_15968,N_15486,N_15370);
or U15969 (N_15969,N_15335,N_15291);
xor U15970 (N_15970,N_15116,N_15462);
or U15971 (N_15971,N_15223,N_15496);
or U15972 (N_15972,N_15089,N_15297);
nor U15973 (N_15973,N_15478,N_15206);
or U15974 (N_15974,N_15298,N_15201);
nand U15975 (N_15975,N_15086,N_15090);
nand U15976 (N_15976,N_15349,N_15400);
nand U15977 (N_15977,N_15037,N_15194);
and U15978 (N_15978,N_15103,N_15294);
xnor U15979 (N_15979,N_15064,N_15194);
nand U15980 (N_15980,N_15429,N_15360);
nor U15981 (N_15981,N_15454,N_15022);
or U15982 (N_15982,N_15142,N_15257);
or U15983 (N_15983,N_15288,N_15253);
nand U15984 (N_15984,N_15414,N_15237);
nor U15985 (N_15985,N_15283,N_15060);
and U15986 (N_15986,N_15315,N_15158);
and U15987 (N_15987,N_15463,N_15423);
or U15988 (N_15988,N_15289,N_15171);
xnor U15989 (N_15989,N_15240,N_15134);
and U15990 (N_15990,N_15045,N_15021);
nor U15991 (N_15991,N_15167,N_15085);
and U15992 (N_15992,N_15418,N_15428);
or U15993 (N_15993,N_15142,N_15352);
nand U15994 (N_15994,N_15364,N_15221);
nor U15995 (N_15995,N_15163,N_15441);
and U15996 (N_15996,N_15152,N_15051);
and U15997 (N_15997,N_15382,N_15386);
or U15998 (N_15998,N_15302,N_15238);
nand U15999 (N_15999,N_15255,N_15156);
nor U16000 (N_16000,N_15933,N_15915);
nand U16001 (N_16001,N_15779,N_15921);
or U16002 (N_16002,N_15524,N_15908);
nor U16003 (N_16003,N_15606,N_15842);
or U16004 (N_16004,N_15574,N_15830);
nand U16005 (N_16005,N_15537,N_15515);
or U16006 (N_16006,N_15698,N_15520);
or U16007 (N_16007,N_15901,N_15594);
and U16008 (N_16008,N_15807,N_15794);
or U16009 (N_16009,N_15723,N_15964);
nor U16010 (N_16010,N_15751,N_15957);
or U16011 (N_16011,N_15589,N_15963);
nor U16012 (N_16012,N_15668,N_15682);
nand U16013 (N_16013,N_15982,N_15743);
and U16014 (N_16014,N_15930,N_15732);
nor U16015 (N_16015,N_15678,N_15927);
nand U16016 (N_16016,N_15812,N_15755);
nand U16017 (N_16017,N_15644,N_15893);
nand U16018 (N_16018,N_15632,N_15689);
xnor U16019 (N_16019,N_15825,N_15772);
nand U16020 (N_16020,N_15838,N_15836);
and U16021 (N_16021,N_15934,N_15938);
nor U16022 (N_16022,N_15502,N_15602);
nand U16023 (N_16023,N_15786,N_15558);
or U16024 (N_16024,N_15652,N_15551);
nand U16025 (N_16025,N_15722,N_15912);
or U16026 (N_16026,N_15840,N_15747);
or U16027 (N_16027,N_15849,N_15834);
nor U16028 (N_16028,N_15960,N_15603);
nor U16029 (N_16029,N_15846,N_15641);
and U16030 (N_16030,N_15752,N_15782);
xnor U16031 (N_16031,N_15775,N_15870);
nand U16032 (N_16032,N_15529,N_15648);
and U16033 (N_16033,N_15561,N_15700);
and U16034 (N_16034,N_15598,N_15985);
and U16035 (N_16035,N_15793,N_15923);
xor U16036 (N_16036,N_15549,N_15882);
nand U16037 (N_16037,N_15528,N_15599);
or U16038 (N_16038,N_15504,N_15925);
or U16039 (N_16039,N_15991,N_15725);
or U16040 (N_16040,N_15523,N_15926);
and U16041 (N_16041,N_15658,N_15684);
nor U16042 (N_16042,N_15685,N_15919);
and U16043 (N_16043,N_15745,N_15571);
nor U16044 (N_16044,N_15810,N_15997);
and U16045 (N_16045,N_15992,N_15680);
nor U16046 (N_16046,N_15897,N_15541);
nor U16047 (N_16047,N_15800,N_15760);
or U16048 (N_16048,N_15629,N_15735);
nand U16049 (N_16049,N_15969,N_15970);
nor U16050 (N_16050,N_15601,N_15519);
nor U16051 (N_16051,N_15681,N_15729);
nor U16052 (N_16052,N_15777,N_15567);
nand U16053 (N_16053,N_15819,N_15778);
xor U16054 (N_16054,N_15693,N_15539);
nor U16055 (N_16055,N_15889,N_15742);
nor U16056 (N_16056,N_15851,N_15974);
nor U16057 (N_16057,N_15749,N_15733);
nor U16058 (N_16058,N_15983,N_15814);
and U16059 (N_16059,N_15904,N_15978);
nor U16060 (N_16060,N_15844,N_15922);
or U16061 (N_16061,N_15590,N_15998);
or U16062 (N_16062,N_15894,N_15500);
and U16063 (N_16063,N_15587,N_15959);
nor U16064 (N_16064,N_15667,N_15746);
nor U16065 (N_16065,N_15664,N_15562);
nand U16066 (N_16066,N_15815,N_15554);
or U16067 (N_16067,N_15649,N_15993);
nor U16068 (N_16068,N_15877,N_15967);
and U16069 (N_16069,N_15999,N_15710);
xor U16070 (N_16070,N_15903,N_15826);
nand U16071 (N_16071,N_15508,N_15679);
xor U16072 (N_16072,N_15550,N_15699);
or U16073 (N_16073,N_15538,N_15696);
nor U16074 (N_16074,N_15885,N_15773);
and U16075 (N_16075,N_15808,N_15929);
nand U16076 (N_16076,N_15707,N_15705);
nor U16077 (N_16077,N_15791,N_15886);
and U16078 (N_16078,N_15940,N_15756);
or U16079 (N_16079,N_15787,N_15823);
or U16080 (N_16080,N_15931,N_15556);
or U16081 (N_16081,N_15637,N_15996);
nand U16082 (N_16082,N_15918,N_15780);
nor U16083 (N_16083,N_15509,N_15513);
nand U16084 (N_16084,N_15741,N_15888);
nand U16085 (N_16085,N_15720,N_15616);
nor U16086 (N_16086,N_15661,N_15552);
or U16087 (N_16087,N_15712,N_15716);
nand U16088 (N_16088,N_15608,N_15687);
and U16089 (N_16089,N_15892,N_15605);
or U16090 (N_16090,N_15543,N_15572);
and U16091 (N_16091,N_15578,N_15953);
or U16092 (N_16092,N_15654,N_15977);
nand U16093 (N_16093,N_15622,N_15692);
or U16094 (N_16094,N_15837,N_15790);
nand U16095 (N_16095,N_15717,N_15560);
nor U16096 (N_16096,N_15765,N_15956);
or U16097 (N_16097,N_15548,N_15845);
and U16098 (N_16098,N_15936,N_15868);
nand U16099 (N_16099,N_15738,N_15950);
and U16100 (N_16100,N_15788,N_15626);
or U16101 (N_16101,N_15517,N_15688);
nor U16102 (N_16102,N_15740,N_15961);
nand U16103 (N_16103,N_15914,N_15505);
nor U16104 (N_16104,N_15564,N_15588);
or U16105 (N_16105,N_15905,N_15766);
nor U16106 (N_16106,N_15816,N_15631);
nand U16107 (N_16107,N_15653,N_15620);
and U16108 (N_16108,N_15609,N_15909);
nor U16109 (N_16109,N_15853,N_15824);
and U16110 (N_16110,N_15623,N_15597);
and U16111 (N_16111,N_15945,N_15569);
nand U16112 (N_16112,N_15625,N_15805);
and U16113 (N_16113,N_15511,N_15833);
nand U16114 (N_16114,N_15878,N_15916);
nand U16115 (N_16115,N_15635,N_15595);
and U16116 (N_16116,N_15636,N_15943);
nor U16117 (N_16117,N_15863,N_15579);
nand U16118 (N_16118,N_15619,N_15618);
and U16119 (N_16119,N_15976,N_15911);
or U16120 (N_16120,N_15984,N_15646);
nor U16121 (N_16121,N_15660,N_15835);
and U16122 (N_16122,N_15932,N_15874);
nor U16123 (N_16123,N_15757,N_15891);
nor U16124 (N_16124,N_15872,N_15762);
xnor U16125 (N_16125,N_15503,N_15890);
nand U16126 (N_16126,N_15785,N_15607);
or U16127 (N_16127,N_15727,N_15758);
nor U16128 (N_16128,N_15827,N_15792);
nand U16129 (N_16129,N_15898,N_15736);
and U16130 (N_16130,N_15718,N_15873);
or U16131 (N_16131,N_15828,N_15686);
and U16132 (N_16132,N_15563,N_15802);
or U16133 (N_16133,N_15713,N_15676);
or U16134 (N_16134,N_15640,N_15638);
and U16135 (N_16135,N_15989,N_15847);
nand U16136 (N_16136,N_15724,N_15744);
nor U16137 (N_16137,N_15737,N_15797);
and U16138 (N_16138,N_15612,N_15952);
and U16139 (N_16139,N_15944,N_15981);
nor U16140 (N_16140,N_15701,N_15973);
nand U16141 (N_16141,N_15941,N_15647);
and U16142 (N_16142,N_15670,N_15665);
or U16143 (N_16143,N_15753,N_15948);
or U16144 (N_16144,N_15799,N_15867);
nand U16145 (N_16145,N_15582,N_15994);
or U16146 (N_16146,N_15795,N_15839);
or U16147 (N_16147,N_15801,N_15798);
and U16148 (N_16148,N_15856,N_15610);
nor U16149 (N_16149,N_15821,N_15883);
nand U16150 (N_16150,N_15881,N_15568);
or U16151 (N_16151,N_15781,N_15734);
nor U16152 (N_16152,N_15591,N_15553);
nor U16153 (N_16153,N_15857,N_15559);
and U16154 (N_16154,N_15596,N_15709);
nand U16155 (N_16155,N_15906,N_15971);
and U16156 (N_16156,N_15672,N_15506);
nand U16157 (N_16157,N_15869,N_15990);
nand U16158 (N_16158,N_15955,N_15593);
nand U16159 (N_16159,N_15613,N_15771);
nand U16160 (N_16160,N_15750,N_15655);
and U16161 (N_16161,N_15659,N_15864);
and U16162 (N_16162,N_15774,N_15817);
and U16163 (N_16163,N_15575,N_15674);
nor U16164 (N_16164,N_15630,N_15580);
nor U16165 (N_16165,N_15565,N_15951);
nor U16166 (N_16166,N_15592,N_15900);
nor U16167 (N_16167,N_15866,N_15545);
nor U16168 (N_16168,N_15577,N_15604);
nand U16169 (N_16169,N_15706,N_15617);
or U16170 (N_16170,N_15980,N_15697);
nor U16171 (N_16171,N_15715,N_15547);
nand U16172 (N_16172,N_15995,N_15731);
and U16173 (N_16173,N_15666,N_15576);
or U16174 (N_16174,N_15586,N_15555);
and U16175 (N_16175,N_15536,N_15895);
nor U16176 (N_16176,N_15841,N_15962);
or U16177 (N_16177,N_15848,N_15739);
or U16178 (N_16178,N_15714,N_15673);
nor U16179 (N_16179,N_15645,N_15763);
or U16180 (N_16180,N_15761,N_15913);
nand U16181 (N_16181,N_15704,N_15861);
nor U16182 (N_16182,N_15979,N_15776);
nor U16183 (N_16183,N_15811,N_15708);
and U16184 (N_16184,N_15691,N_15946);
nand U16185 (N_16185,N_15643,N_15860);
nand U16186 (N_16186,N_15822,N_15510);
and U16187 (N_16187,N_15784,N_15726);
nor U16188 (N_16188,N_15767,N_15690);
nand U16189 (N_16189,N_15942,N_15975);
nand U16190 (N_16190,N_15862,N_15768);
or U16191 (N_16191,N_15702,N_15884);
nor U16192 (N_16192,N_15854,N_15907);
and U16193 (N_16193,N_15879,N_15829);
xor U16194 (N_16194,N_15624,N_15831);
nor U16195 (N_16195,N_15677,N_15516);
nand U16196 (N_16196,N_15642,N_15535);
nor U16197 (N_16197,N_15512,N_15695);
and U16198 (N_16198,N_15533,N_15614);
nand U16199 (N_16199,N_15628,N_15651);
and U16200 (N_16200,N_15947,N_15669);
nor U16201 (N_16201,N_15966,N_15570);
and U16202 (N_16202,N_15526,N_15859);
and U16203 (N_16203,N_15711,N_15852);
and U16204 (N_16204,N_15887,N_15540);
and U16205 (N_16205,N_15656,N_15759);
nand U16206 (N_16206,N_15809,N_15764);
nand U16207 (N_16207,N_15968,N_15939);
xor U16208 (N_16208,N_15583,N_15719);
or U16209 (N_16209,N_15899,N_15518);
or U16210 (N_16210,N_15544,N_15585);
nand U16211 (N_16211,N_15843,N_15965);
or U16212 (N_16212,N_15910,N_15858);
and U16213 (N_16213,N_15611,N_15527);
nand U16214 (N_16214,N_15820,N_15972);
nand U16215 (N_16215,N_15657,N_15662);
or U16216 (N_16216,N_15789,N_15871);
or U16217 (N_16217,N_15850,N_15748);
nand U16218 (N_16218,N_15522,N_15986);
xnor U16219 (N_16219,N_15675,N_15530);
nand U16220 (N_16220,N_15573,N_15896);
or U16221 (N_16221,N_15615,N_15639);
nor U16222 (N_16222,N_15514,N_15832);
nor U16223 (N_16223,N_15683,N_15525);
or U16224 (N_16224,N_15803,N_15581);
or U16225 (N_16225,N_15621,N_15855);
or U16226 (N_16226,N_15521,N_15730);
nand U16227 (N_16227,N_15880,N_15671);
or U16228 (N_16228,N_15917,N_15532);
nand U16229 (N_16229,N_15876,N_15958);
and U16230 (N_16230,N_15806,N_15627);
nand U16231 (N_16231,N_15988,N_15935);
nor U16232 (N_16232,N_15531,N_15542);
nor U16233 (N_16233,N_15703,N_15928);
nor U16234 (N_16234,N_15813,N_15920);
nor U16235 (N_16235,N_15600,N_15584);
nand U16236 (N_16236,N_15783,N_15796);
and U16237 (N_16237,N_15875,N_15566);
and U16238 (N_16238,N_15770,N_15987);
or U16239 (N_16239,N_15804,N_15507);
xor U16240 (N_16240,N_15721,N_15865);
or U16241 (N_16241,N_15949,N_15902);
nor U16242 (N_16242,N_15557,N_15769);
nand U16243 (N_16243,N_15924,N_15663);
or U16244 (N_16244,N_15501,N_15534);
and U16245 (N_16245,N_15633,N_15546);
and U16246 (N_16246,N_15728,N_15650);
or U16247 (N_16247,N_15754,N_15954);
or U16248 (N_16248,N_15694,N_15634);
and U16249 (N_16249,N_15818,N_15937);
nand U16250 (N_16250,N_15833,N_15990);
nor U16251 (N_16251,N_15545,N_15574);
and U16252 (N_16252,N_15780,N_15509);
nor U16253 (N_16253,N_15516,N_15518);
and U16254 (N_16254,N_15619,N_15871);
or U16255 (N_16255,N_15659,N_15777);
nor U16256 (N_16256,N_15700,N_15782);
nand U16257 (N_16257,N_15823,N_15707);
nor U16258 (N_16258,N_15908,N_15858);
and U16259 (N_16259,N_15932,N_15992);
nor U16260 (N_16260,N_15545,N_15597);
or U16261 (N_16261,N_15662,N_15520);
and U16262 (N_16262,N_15637,N_15728);
and U16263 (N_16263,N_15709,N_15881);
nor U16264 (N_16264,N_15767,N_15709);
or U16265 (N_16265,N_15786,N_15808);
nand U16266 (N_16266,N_15653,N_15740);
or U16267 (N_16267,N_15814,N_15770);
or U16268 (N_16268,N_15759,N_15635);
nand U16269 (N_16269,N_15999,N_15963);
and U16270 (N_16270,N_15966,N_15738);
and U16271 (N_16271,N_15730,N_15749);
and U16272 (N_16272,N_15845,N_15526);
and U16273 (N_16273,N_15534,N_15662);
xnor U16274 (N_16274,N_15644,N_15546);
and U16275 (N_16275,N_15524,N_15876);
xor U16276 (N_16276,N_15689,N_15995);
and U16277 (N_16277,N_15743,N_15585);
nor U16278 (N_16278,N_15683,N_15916);
nand U16279 (N_16279,N_15889,N_15874);
nand U16280 (N_16280,N_15816,N_15857);
or U16281 (N_16281,N_15596,N_15560);
nor U16282 (N_16282,N_15809,N_15674);
or U16283 (N_16283,N_15584,N_15597);
nand U16284 (N_16284,N_15755,N_15945);
and U16285 (N_16285,N_15749,N_15598);
nand U16286 (N_16286,N_15577,N_15995);
nor U16287 (N_16287,N_15720,N_15936);
nand U16288 (N_16288,N_15535,N_15669);
nor U16289 (N_16289,N_15894,N_15584);
nor U16290 (N_16290,N_15786,N_15615);
xor U16291 (N_16291,N_15852,N_15721);
nor U16292 (N_16292,N_15724,N_15890);
nand U16293 (N_16293,N_15908,N_15646);
nand U16294 (N_16294,N_15788,N_15793);
and U16295 (N_16295,N_15791,N_15955);
nor U16296 (N_16296,N_15959,N_15564);
and U16297 (N_16297,N_15879,N_15838);
nand U16298 (N_16298,N_15961,N_15814);
nor U16299 (N_16299,N_15869,N_15772);
or U16300 (N_16300,N_15649,N_15798);
nor U16301 (N_16301,N_15931,N_15713);
nand U16302 (N_16302,N_15668,N_15844);
or U16303 (N_16303,N_15953,N_15966);
and U16304 (N_16304,N_15992,N_15591);
nor U16305 (N_16305,N_15892,N_15662);
or U16306 (N_16306,N_15938,N_15723);
nor U16307 (N_16307,N_15676,N_15929);
or U16308 (N_16308,N_15776,N_15849);
and U16309 (N_16309,N_15670,N_15685);
nand U16310 (N_16310,N_15950,N_15505);
nor U16311 (N_16311,N_15794,N_15732);
nand U16312 (N_16312,N_15825,N_15774);
nand U16313 (N_16313,N_15857,N_15582);
or U16314 (N_16314,N_15703,N_15919);
xor U16315 (N_16315,N_15861,N_15600);
and U16316 (N_16316,N_15872,N_15695);
nor U16317 (N_16317,N_15993,N_15629);
nor U16318 (N_16318,N_15837,N_15607);
nand U16319 (N_16319,N_15677,N_15901);
or U16320 (N_16320,N_15656,N_15711);
and U16321 (N_16321,N_15847,N_15888);
and U16322 (N_16322,N_15929,N_15666);
nor U16323 (N_16323,N_15798,N_15819);
or U16324 (N_16324,N_15720,N_15609);
nor U16325 (N_16325,N_15998,N_15501);
nor U16326 (N_16326,N_15870,N_15603);
xnor U16327 (N_16327,N_15663,N_15662);
nor U16328 (N_16328,N_15957,N_15885);
or U16329 (N_16329,N_15623,N_15667);
and U16330 (N_16330,N_15751,N_15856);
nor U16331 (N_16331,N_15910,N_15816);
or U16332 (N_16332,N_15727,N_15916);
nor U16333 (N_16333,N_15965,N_15678);
nand U16334 (N_16334,N_15796,N_15651);
or U16335 (N_16335,N_15689,N_15733);
or U16336 (N_16336,N_15814,N_15889);
xor U16337 (N_16337,N_15624,N_15658);
and U16338 (N_16338,N_15548,N_15791);
nor U16339 (N_16339,N_15668,N_15981);
or U16340 (N_16340,N_15812,N_15900);
or U16341 (N_16341,N_15862,N_15662);
nand U16342 (N_16342,N_15853,N_15735);
or U16343 (N_16343,N_15660,N_15685);
and U16344 (N_16344,N_15899,N_15670);
nor U16345 (N_16345,N_15840,N_15689);
and U16346 (N_16346,N_15540,N_15566);
nor U16347 (N_16347,N_15590,N_15752);
nor U16348 (N_16348,N_15912,N_15581);
or U16349 (N_16349,N_15803,N_15876);
and U16350 (N_16350,N_15727,N_15786);
nor U16351 (N_16351,N_15924,N_15614);
nor U16352 (N_16352,N_15711,N_15846);
or U16353 (N_16353,N_15867,N_15910);
nor U16354 (N_16354,N_15836,N_15941);
nor U16355 (N_16355,N_15910,N_15979);
and U16356 (N_16356,N_15753,N_15800);
and U16357 (N_16357,N_15674,N_15658);
nor U16358 (N_16358,N_15740,N_15707);
nor U16359 (N_16359,N_15503,N_15707);
or U16360 (N_16360,N_15806,N_15964);
and U16361 (N_16361,N_15993,N_15949);
nand U16362 (N_16362,N_15873,N_15840);
or U16363 (N_16363,N_15845,N_15738);
xor U16364 (N_16364,N_15765,N_15822);
or U16365 (N_16365,N_15872,N_15626);
nand U16366 (N_16366,N_15969,N_15745);
nor U16367 (N_16367,N_15633,N_15845);
xnor U16368 (N_16368,N_15663,N_15695);
and U16369 (N_16369,N_15631,N_15797);
or U16370 (N_16370,N_15692,N_15965);
nor U16371 (N_16371,N_15509,N_15994);
nor U16372 (N_16372,N_15860,N_15846);
nor U16373 (N_16373,N_15845,N_15663);
nor U16374 (N_16374,N_15533,N_15570);
nor U16375 (N_16375,N_15772,N_15936);
or U16376 (N_16376,N_15774,N_15585);
and U16377 (N_16377,N_15581,N_15731);
nand U16378 (N_16378,N_15766,N_15589);
nor U16379 (N_16379,N_15558,N_15987);
nor U16380 (N_16380,N_15952,N_15833);
nand U16381 (N_16381,N_15570,N_15783);
and U16382 (N_16382,N_15539,N_15662);
or U16383 (N_16383,N_15687,N_15658);
nand U16384 (N_16384,N_15565,N_15506);
and U16385 (N_16385,N_15534,N_15847);
nand U16386 (N_16386,N_15864,N_15603);
nand U16387 (N_16387,N_15582,N_15828);
nor U16388 (N_16388,N_15875,N_15780);
and U16389 (N_16389,N_15854,N_15600);
nand U16390 (N_16390,N_15857,N_15712);
and U16391 (N_16391,N_15866,N_15953);
nand U16392 (N_16392,N_15695,N_15696);
and U16393 (N_16393,N_15994,N_15876);
or U16394 (N_16394,N_15874,N_15777);
and U16395 (N_16395,N_15849,N_15931);
nor U16396 (N_16396,N_15845,N_15524);
nor U16397 (N_16397,N_15577,N_15501);
xnor U16398 (N_16398,N_15902,N_15619);
and U16399 (N_16399,N_15692,N_15826);
nor U16400 (N_16400,N_15912,N_15982);
or U16401 (N_16401,N_15753,N_15761);
or U16402 (N_16402,N_15733,N_15685);
nand U16403 (N_16403,N_15969,N_15640);
nor U16404 (N_16404,N_15747,N_15906);
nor U16405 (N_16405,N_15626,N_15967);
nand U16406 (N_16406,N_15814,N_15581);
nand U16407 (N_16407,N_15853,N_15899);
nor U16408 (N_16408,N_15580,N_15894);
nand U16409 (N_16409,N_15686,N_15977);
nand U16410 (N_16410,N_15972,N_15509);
nor U16411 (N_16411,N_15556,N_15676);
and U16412 (N_16412,N_15943,N_15628);
and U16413 (N_16413,N_15763,N_15556);
nand U16414 (N_16414,N_15769,N_15512);
and U16415 (N_16415,N_15554,N_15929);
nand U16416 (N_16416,N_15863,N_15509);
and U16417 (N_16417,N_15851,N_15824);
or U16418 (N_16418,N_15571,N_15539);
nand U16419 (N_16419,N_15883,N_15852);
and U16420 (N_16420,N_15736,N_15800);
or U16421 (N_16421,N_15885,N_15534);
nand U16422 (N_16422,N_15698,N_15742);
and U16423 (N_16423,N_15898,N_15658);
nand U16424 (N_16424,N_15515,N_15610);
nor U16425 (N_16425,N_15983,N_15963);
nand U16426 (N_16426,N_15822,N_15600);
nor U16427 (N_16427,N_15724,N_15987);
or U16428 (N_16428,N_15706,N_15624);
or U16429 (N_16429,N_15834,N_15855);
nand U16430 (N_16430,N_15999,N_15638);
nand U16431 (N_16431,N_15963,N_15954);
and U16432 (N_16432,N_15683,N_15684);
nand U16433 (N_16433,N_15622,N_15696);
nor U16434 (N_16434,N_15721,N_15609);
and U16435 (N_16435,N_15754,N_15580);
and U16436 (N_16436,N_15923,N_15879);
and U16437 (N_16437,N_15513,N_15832);
nand U16438 (N_16438,N_15523,N_15974);
and U16439 (N_16439,N_15629,N_15972);
and U16440 (N_16440,N_15915,N_15906);
and U16441 (N_16441,N_15760,N_15588);
nand U16442 (N_16442,N_15990,N_15538);
nand U16443 (N_16443,N_15681,N_15644);
nand U16444 (N_16444,N_15828,N_15517);
or U16445 (N_16445,N_15615,N_15698);
xor U16446 (N_16446,N_15506,N_15623);
or U16447 (N_16447,N_15866,N_15757);
nor U16448 (N_16448,N_15689,N_15774);
and U16449 (N_16449,N_15567,N_15822);
nand U16450 (N_16450,N_15834,N_15726);
nor U16451 (N_16451,N_15648,N_15832);
nor U16452 (N_16452,N_15732,N_15954);
or U16453 (N_16453,N_15792,N_15812);
nor U16454 (N_16454,N_15874,N_15583);
and U16455 (N_16455,N_15601,N_15755);
nor U16456 (N_16456,N_15937,N_15971);
nor U16457 (N_16457,N_15945,N_15808);
and U16458 (N_16458,N_15837,N_15516);
and U16459 (N_16459,N_15795,N_15863);
nor U16460 (N_16460,N_15808,N_15871);
nor U16461 (N_16461,N_15694,N_15972);
nor U16462 (N_16462,N_15572,N_15986);
or U16463 (N_16463,N_15849,N_15786);
nand U16464 (N_16464,N_15710,N_15955);
nor U16465 (N_16465,N_15588,N_15678);
nand U16466 (N_16466,N_15621,N_15859);
nor U16467 (N_16467,N_15679,N_15631);
or U16468 (N_16468,N_15866,N_15723);
or U16469 (N_16469,N_15717,N_15854);
nor U16470 (N_16470,N_15638,N_15674);
or U16471 (N_16471,N_15981,N_15861);
nor U16472 (N_16472,N_15852,N_15734);
nand U16473 (N_16473,N_15889,N_15611);
nand U16474 (N_16474,N_15867,N_15797);
nand U16475 (N_16475,N_15506,N_15799);
and U16476 (N_16476,N_15626,N_15759);
or U16477 (N_16477,N_15828,N_15545);
or U16478 (N_16478,N_15753,N_15591);
nand U16479 (N_16479,N_15990,N_15672);
nand U16480 (N_16480,N_15585,N_15812);
nor U16481 (N_16481,N_15886,N_15665);
or U16482 (N_16482,N_15563,N_15575);
nand U16483 (N_16483,N_15650,N_15667);
nor U16484 (N_16484,N_15520,N_15743);
nand U16485 (N_16485,N_15757,N_15570);
and U16486 (N_16486,N_15541,N_15932);
nor U16487 (N_16487,N_15746,N_15972);
nor U16488 (N_16488,N_15503,N_15795);
nand U16489 (N_16489,N_15944,N_15516);
xor U16490 (N_16490,N_15881,N_15656);
nand U16491 (N_16491,N_15764,N_15556);
and U16492 (N_16492,N_15679,N_15855);
xnor U16493 (N_16493,N_15852,N_15779);
or U16494 (N_16494,N_15520,N_15970);
xnor U16495 (N_16495,N_15550,N_15504);
nand U16496 (N_16496,N_15912,N_15511);
nand U16497 (N_16497,N_15820,N_15531);
nor U16498 (N_16498,N_15954,N_15678);
nand U16499 (N_16499,N_15759,N_15838);
and U16500 (N_16500,N_16435,N_16417);
nor U16501 (N_16501,N_16133,N_16480);
xor U16502 (N_16502,N_16363,N_16042);
nand U16503 (N_16503,N_16051,N_16348);
and U16504 (N_16504,N_16370,N_16441);
and U16505 (N_16505,N_16488,N_16162);
and U16506 (N_16506,N_16379,N_16131);
or U16507 (N_16507,N_16030,N_16038);
nand U16508 (N_16508,N_16144,N_16227);
nand U16509 (N_16509,N_16338,N_16235);
nand U16510 (N_16510,N_16310,N_16397);
nand U16511 (N_16511,N_16386,N_16306);
or U16512 (N_16512,N_16195,N_16389);
or U16513 (N_16513,N_16199,N_16164);
or U16514 (N_16514,N_16076,N_16058);
nand U16515 (N_16515,N_16097,N_16203);
and U16516 (N_16516,N_16433,N_16439);
nor U16517 (N_16517,N_16110,N_16192);
and U16518 (N_16518,N_16005,N_16047);
and U16519 (N_16519,N_16443,N_16425);
nor U16520 (N_16520,N_16326,N_16213);
nand U16521 (N_16521,N_16266,N_16264);
or U16522 (N_16522,N_16428,N_16265);
and U16523 (N_16523,N_16314,N_16095);
or U16524 (N_16524,N_16469,N_16361);
nor U16525 (N_16525,N_16218,N_16115);
xnor U16526 (N_16526,N_16378,N_16109);
or U16527 (N_16527,N_16478,N_16082);
nand U16528 (N_16528,N_16270,N_16028);
nand U16529 (N_16529,N_16394,N_16299);
nor U16530 (N_16530,N_16219,N_16209);
and U16531 (N_16531,N_16268,N_16188);
nand U16532 (N_16532,N_16059,N_16016);
nor U16533 (N_16533,N_16167,N_16273);
nand U16534 (N_16534,N_16071,N_16367);
nand U16535 (N_16535,N_16026,N_16241);
xor U16536 (N_16536,N_16248,N_16420);
or U16537 (N_16537,N_16201,N_16399);
or U16538 (N_16538,N_16422,N_16407);
and U16539 (N_16539,N_16410,N_16369);
or U16540 (N_16540,N_16359,N_16258);
or U16541 (N_16541,N_16357,N_16458);
xor U16542 (N_16542,N_16223,N_16060);
nand U16543 (N_16543,N_16096,N_16020);
and U16544 (N_16544,N_16288,N_16175);
xor U16545 (N_16545,N_16041,N_16050);
xnor U16546 (N_16546,N_16197,N_16090);
nand U16547 (N_16547,N_16143,N_16491);
and U16548 (N_16548,N_16252,N_16474);
nand U16549 (N_16549,N_16345,N_16204);
nor U16550 (N_16550,N_16151,N_16230);
nor U16551 (N_16551,N_16382,N_16154);
nor U16552 (N_16552,N_16206,N_16298);
xor U16553 (N_16553,N_16043,N_16499);
nand U16554 (N_16554,N_16086,N_16044);
or U16555 (N_16555,N_16452,N_16275);
and U16556 (N_16556,N_16457,N_16472);
and U16557 (N_16557,N_16125,N_16145);
and U16558 (N_16558,N_16036,N_16494);
nand U16559 (N_16559,N_16496,N_16261);
nand U16560 (N_16560,N_16277,N_16205);
nor U16561 (N_16561,N_16099,N_16000);
nand U16562 (N_16562,N_16210,N_16001);
nand U16563 (N_16563,N_16136,N_16490);
or U16564 (N_16564,N_16214,N_16272);
nand U16565 (N_16565,N_16291,N_16098);
and U16566 (N_16566,N_16347,N_16448);
nor U16567 (N_16567,N_16054,N_16108);
and U16568 (N_16568,N_16321,N_16148);
nor U16569 (N_16569,N_16146,N_16202);
or U16570 (N_16570,N_16160,N_16333);
or U16571 (N_16571,N_16405,N_16374);
nor U16572 (N_16572,N_16328,N_16150);
nor U16573 (N_16573,N_16411,N_16116);
nor U16574 (N_16574,N_16222,N_16142);
nand U16575 (N_16575,N_16445,N_16487);
nand U16576 (N_16576,N_16147,N_16119);
xnor U16577 (N_16577,N_16062,N_16406);
and U16578 (N_16578,N_16346,N_16126);
or U16579 (N_16579,N_16093,N_16106);
or U16580 (N_16580,N_16416,N_16052);
nor U16581 (N_16581,N_16372,N_16412);
nor U16582 (N_16582,N_16069,N_16470);
and U16583 (N_16583,N_16007,N_16293);
nand U16584 (N_16584,N_16233,N_16077);
nor U16585 (N_16585,N_16262,N_16200);
or U16586 (N_16586,N_16246,N_16174);
and U16587 (N_16587,N_16396,N_16239);
or U16588 (N_16588,N_16232,N_16418);
nor U16589 (N_16589,N_16249,N_16476);
nand U16590 (N_16590,N_16074,N_16274);
or U16591 (N_16591,N_16295,N_16193);
nor U16592 (N_16592,N_16353,N_16294);
or U16593 (N_16593,N_16449,N_16065);
and U16594 (N_16594,N_16240,N_16319);
or U16595 (N_16595,N_16178,N_16256);
and U16596 (N_16596,N_16434,N_16247);
and U16597 (N_16597,N_16339,N_16023);
nor U16598 (N_16598,N_16008,N_16032);
and U16599 (N_16599,N_16413,N_16436);
nand U16600 (N_16600,N_16152,N_16226);
and U16601 (N_16601,N_16373,N_16066);
nor U16602 (N_16602,N_16254,N_16037);
nand U16603 (N_16603,N_16045,N_16191);
and U16604 (N_16604,N_16013,N_16228);
and U16605 (N_16605,N_16376,N_16313);
and U16606 (N_16606,N_16278,N_16383);
or U16607 (N_16607,N_16215,N_16401);
xor U16608 (N_16608,N_16207,N_16498);
and U16609 (N_16609,N_16300,N_16068);
nor U16610 (N_16610,N_16092,N_16094);
nand U16611 (N_16611,N_16010,N_16465);
or U16612 (N_16612,N_16385,N_16332);
or U16613 (N_16613,N_16260,N_16061);
nor U16614 (N_16614,N_16320,N_16113);
or U16615 (N_16615,N_16212,N_16006);
and U16616 (N_16616,N_16466,N_16134);
or U16617 (N_16617,N_16170,N_16414);
or U16618 (N_16618,N_16075,N_16089);
and U16619 (N_16619,N_16473,N_16390);
nor U16620 (N_16620,N_16444,N_16477);
nand U16621 (N_16621,N_16194,N_16381);
nand U16622 (N_16622,N_16427,N_16137);
or U16623 (N_16623,N_16269,N_16351);
nor U16624 (N_16624,N_16423,N_16451);
nor U16625 (N_16625,N_16067,N_16308);
nor U16626 (N_16626,N_16124,N_16190);
and U16627 (N_16627,N_16362,N_16341);
nor U16628 (N_16628,N_16208,N_16325);
and U16629 (N_16629,N_16336,N_16029);
and U16630 (N_16630,N_16460,N_16140);
nand U16631 (N_16631,N_16404,N_16039);
nor U16632 (N_16632,N_16078,N_16118);
or U16633 (N_16633,N_16450,N_16127);
or U16634 (N_16634,N_16354,N_16327);
xor U16635 (N_16635,N_16112,N_16081);
nand U16636 (N_16636,N_16316,N_16022);
and U16637 (N_16637,N_16305,N_16189);
nor U16638 (N_16638,N_16440,N_16350);
or U16639 (N_16639,N_16244,N_16056);
and U16640 (N_16640,N_16107,N_16177);
nor U16641 (N_16641,N_16419,N_16392);
and U16642 (N_16642,N_16117,N_16253);
xor U16643 (N_16643,N_16138,N_16358);
nand U16644 (N_16644,N_16464,N_16055);
nand U16645 (N_16645,N_16122,N_16403);
nand U16646 (N_16646,N_16322,N_16475);
xnor U16647 (N_16647,N_16159,N_16085);
and U16648 (N_16648,N_16461,N_16371);
and U16649 (N_16649,N_16290,N_16395);
or U16650 (N_16650,N_16432,N_16187);
nand U16651 (N_16651,N_16317,N_16088);
nor U16652 (N_16652,N_16287,N_16297);
or U16653 (N_16653,N_16083,N_16179);
and U16654 (N_16654,N_16468,N_16072);
nor U16655 (N_16655,N_16015,N_16103);
and U16656 (N_16656,N_16387,N_16285);
nand U16657 (N_16657,N_16349,N_16046);
and U16658 (N_16658,N_16485,N_16454);
nand U16659 (N_16659,N_16211,N_16400);
nand U16660 (N_16660,N_16289,N_16421);
and U16661 (N_16661,N_16302,N_16459);
and U16662 (N_16662,N_16084,N_16132);
and U16663 (N_16663,N_16257,N_16493);
or U16664 (N_16664,N_16331,N_16365);
nand U16665 (N_16665,N_16196,N_16180);
nor U16666 (N_16666,N_16442,N_16337);
nand U16667 (N_16667,N_16017,N_16087);
nand U16668 (N_16668,N_16157,N_16121);
and U16669 (N_16669,N_16323,N_16217);
or U16670 (N_16670,N_16255,N_16415);
nor U16671 (N_16671,N_16155,N_16161);
or U16672 (N_16672,N_16221,N_16169);
nor U16673 (N_16673,N_16250,N_16281);
and U16674 (N_16674,N_16156,N_16114);
and U16675 (N_16675,N_16398,N_16158);
or U16676 (N_16676,N_16426,N_16334);
and U16677 (N_16677,N_16111,N_16120);
nand U16678 (N_16678,N_16479,N_16129);
nor U16679 (N_16679,N_16024,N_16329);
or U16680 (N_16680,N_16003,N_16021);
nand U16681 (N_16681,N_16267,N_16002);
nor U16682 (N_16682,N_16163,N_16139);
nor U16683 (N_16683,N_16079,N_16318);
nor U16684 (N_16684,N_16027,N_16409);
xor U16685 (N_16685,N_16276,N_16324);
nand U16686 (N_16686,N_16463,N_16360);
or U16687 (N_16687,N_16183,N_16040);
xnor U16688 (N_16688,N_16186,N_16467);
and U16689 (N_16689,N_16063,N_16438);
nand U16690 (N_16690,N_16057,N_16185);
nor U16691 (N_16691,N_16446,N_16198);
xnor U16692 (N_16692,N_16303,N_16296);
nor U16693 (N_16693,N_16408,N_16166);
and U16694 (N_16694,N_16286,N_16242);
and U16695 (N_16695,N_16388,N_16168);
nor U16696 (N_16696,N_16355,N_16455);
nand U16697 (N_16697,N_16173,N_16482);
nor U16698 (N_16698,N_16238,N_16128);
and U16699 (N_16699,N_16181,N_16031);
and U16700 (N_16700,N_16123,N_16453);
nor U16701 (N_16701,N_16053,N_16149);
nor U16702 (N_16702,N_16271,N_16391);
nand U16703 (N_16703,N_16251,N_16343);
nor U16704 (N_16704,N_16033,N_16165);
or U16705 (N_16705,N_16495,N_16224);
nor U16706 (N_16706,N_16497,N_16301);
nor U16707 (N_16707,N_16462,N_16234);
nor U16708 (N_16708,N_16034,N_16153);
and U16709 (N_16709,N_16014,N_16486);
or U16710 (N_16710,N_16080,N_16259);
and U16711 (N_16711,N_16292,N_16375);
nand U16712 (N_16712,N_16431,N_16130);
nand U16713 (N_16713,N_16100,N_16216);
and U16714 (N_16714,N_16492,N_16048);
and U16715 (N_16715,N_16073,N_16012);
nand U16716 (N_16716,N_16340,N_16035);
and U16717 (N_16717,N_16245,N_16447);
nand U16718 (N_16718,N_16064,N_16309);
xnor U16719 (N_16719,N_16311,N_16330);
or U16720 (N_16720,N_16380,N_16489);
and U16721 (N_16721,N_16049,N_16011);
nand U16722 (N_16722,N_16220,N_16229);
nor U16723 (N_16723,N_16101,N_16104);
or U16724 (N_16724,N_16171,N_16018);
nand U16725 (N_16725,N_16364,N_16025);
nor U16726 (N_16726,N_16283,N_16182);
nor U16727 (N_16727,N_16172,N_16236);
nand U16728 (N_16728,N_16377,N_16004);
nand U16729 (N_16729,N_16263,N_16437);
nor U16730 (N_16730,N_16019,N_16481);
nor U16731 (N_16731,N_16237,N_16231);
or U16732 (N_16732,N_16282,N_16105);
and U16733 (N_16733,N_16091,N_16483);
nand U16734 (N_16734,N_16456,N_16307);
or U16735 (N_16735,N_16070,N_16315);
or U16736 (N_16736,N_16280,N_16368);
and U16737 (N_16737,N_16312,N_16366);
and U16738 (N_16738,N_16335,N_16184);
nand U16739 (N_16739,N_16102,N_16342);
nor U16740 (N_16740,N_16384,N_16430);
or U16741 (N_16741,N_16352,N_16393);
nor U16742 (N_16742,N_16429,N_16225);
and U16743 (N_16743,N_16484,N_16141);
nor U16744 (N_16744,N_16284,N_16243);
or U16745 (N_16745,N_16471,N_16135);
nand U16746 (N_16746,N_16304,N_16424);
nand U16747 (N_16747,N_16402,N_16356);
nand U16748 (N_16748,N_16344,N_16009);
or U16749 (N_16749,N_16176,N_16279);
nor U16750 (N_16750,N_16080,N_16245);
nor U16751 (N_16751,N_16214,N_16094);
nor U16752 (N_16752,N_16032,N_16005);
or U16753 (N_16753,N_16283,N_16161);
nand U16754 (N_16754,N_16103,N_16457);
nand U16755 (N_16755,N_16163,N_16122);
or U16756 (N_16756,N_16320,N_16479);
nor U16757 (N_16757,N_16277,N_16330);
nor U16758 (N_16758,N_16043,N_16479);
or U16759 (N_16759,N_16081,N_16226);
or U16760 (N_16760,N_16090,N_16055);
and U16761 (N_16761,N_16107,N_16081);
nor U16762 (N_16762,N_16018,N_16465);
or U16763 (N_16763,N_16472,N_16284);
nand U16764 (N_16764,N_16256,N_16289);
nor U16765 (N_16765,N_16098,N_16256);
and U16766 (N_16766,N_16188,N_16489);
xnor U16767 (N_16767,N_16266,N_16339);
and U16768 (N_16768,N_16361,N_16221);
nand U16769 (N_16769,N_16304,N_16473);
or U16770 (N_16770,N_16102,N_16013);
and U16771 (N_16771,N_16412,N_16084);
nand U16772 (N_16772,N_16359,N_16366);
and U16773 (N_16773,N_16260,N_16213);
nor U16774 (N_16774,N_16330,N_16005);
nand U16775 (N_16775,N_16404,N_16498);
and U16776 (N_16776,N_16112,N_16007);
nand U16777 (N_16777,N_16018,N_16054);
nor U16778 (N_16778,N_16439,N_16494);
or U16779 (N_16779,N_16406,N_16337);
and U16780 (N_16780,N_16197,N_16116);
nor U16781 (N_16781,N_16385,N_16151);
nand U16782 (N_16782,N_16401,N_16253);
nor U16783 (N_16783,N_16291,N_16312);
or U16784 (N_16784,N_16243,N_16324);
and U16785 (N_16785,N_16302,N_16309);
and U16786 (N_16786,N_16484,N_16071);
nand U16787 (N_16787,N_16445,N_16184);
and U16788 (N_16788,N_16392,N_16231);
or U16789 (N_16789,N_16201,N_16403);
nor U16790 (N_16790,N_16437,N_16488);
nand U16791 (N_16791,N_16481,N_16012);
or U16792 (N_16792,N_16106,N_16114);
nor U16793 (N_16793,N_16356,N_16020);
nor U16794 (N_16794,N_16090,N_16315);
and U16795 (N_16795,N_16035,N_16341);
or U16796 (N_16796,N_16453,N_16203);
nand U16797 (N_16797,N_16193,N_16409);
or U16798 (N_16798,N_16044,N_16377);
nor U16799 (N_16799,N_16437,N_16313);
or U16800 (N_16800,N_16299,N_16013);
and U16801 (N_16801,N_16111,N_16287);
and U16802 (N_16802,N_16277,N_16292);
or U16803 (N_16803,N_16237,N_16049);
nor U16804 (N_16804,N_16328,N_16496);
nor U16805 (N_16805,N_16004,N_16345);
nor U16806 (N_16806,N_16437,N_16325);
nor U16807 (N_16807,N_16180,N_16232);
nand U16808 (N_16808,N_16176,N_16433);
or U16809 (N_16809,N_16034,N_16170);
nor U16810 (N_16810,N_16207,N_16490);
and U16811 (N_16811,N_16417,N_16323);
or U16812 (N_16812,N_16038,N_16237);
nor U16813 (N_16813,N_16455,N_16196);
nand U16814 (N_16814,N_16031,N_16377);
and U16815 (N_16815,N_16096,N_16245);
or U16816 (N_16816,N_16389,N_16202);
or U16817 (N_16817,N_16074,N_16340);
nand U16818 (N_16818,N_16098,N_16406);
nand U16819 (N_16819,N_16267,N_16461);
and U16820 (N_16820,N_16371,N_16468);
or U16821 (N_16821,N_16171,N_16499);
or U16822 (N_16822,N_16071,N_16405);
nand U16823 (N_16823,N_16369,N_16067);
or U16824 (N_16824,N_16448,N_16008);
or U16825 (N_16825,N_16212,N_16050);
nor U16826 (N_16826,N_16294,N_16239);
and U16827 (N_16827,N_16262,N_16221);
nand U16828 (N_16828,N_16233,N_16305);
and U16829 (N_16829,N_16378,N_16408);
nand U16830 (N_16830,N_16047,N_16361);
and U16831 (N_16831,N_16314,N_16226);
nand U16832 (N_16832,N_16051,N_16037);
and U16833 (N_16833,N_16349,N_16391);
and U16834 (N_16834,N_16079,N_16217);
nor U16835 (N_16835,N_16446,N_16141);
nand U16836 (N_16836,N_16127,N_16227);
or U16837 (N_16837,N_16269,N_16108);
nor U16838 (N_16838,N_16281,N_16478);
xnor U16839 (N_16839,N_16408,N_16177);
nor U16840 (N_16840,N_16069,N_16011);
or U16841 (N_16841,N_16162,N_16464);
nand U16842 (N_16842,N_16005,N_16056);
nor U16843 (N_16843,N_16283,N_16372);
and U16844 (N_16844,N_16258,N_16158);
and U16845 (N_16845,N_16080,N_16188);
nor U16846 (N_16846,N_16074,N_16299);
or U16847 (N_16847,N_16167,N_16368);
nand U16848 (N_16848,N_16466,N_16232);
nor U16849 (N_16849,N_16327,N_16028);
and U16850 (N_16850,N_16270,N_16172);
or U16851 (N_16851,N_16163,N_16476);
and U16852 (N_16852,N_16122,N_16259);
nand U16853 (N_16853,N_16213,N_16078);
nand U16854 (N_16854,N_16371,N_16072);
or U16855 (N_16855,N_16274,N_16490);
or U16856 (N_16856,N_16089,N_16204);
nand U16857 (N_16857,N_16308,N_16463);
nand U16858 (N_16858,N_16227,N_16330);
nand U16859 (N_16859,N_16317,N_16030);
nor U16860 (N_16860,N_16032,N_16073);
nand U16861 (N_16861,N_16281,N_16056);
nor U16862 (N_16862,N_16302,N_16294);
and U16863 (N_16863,N_16161,N_16046);
xor U16864 (N_16864,N_16074,N_16008);
nand U16865 (N_16865,N_16147,N_16139);
nor U16866 (N_16866,N_16002,N_16088);
and U16867 (N_16867,N_16313,N_16347);
or U16868 (N_16868,N_16008,N_16346);
nand U16869 (N_16869,N_16136,N_16446);
or U16870 (N_16870,N_16365,N_16230);
nor U16871 (N_16871,N_16468,N_16237);
and U16872 (N_16872,N_16440,N_16001);
or U16873 (N_16873,N_16400,N_16334);
nand U16874 (N_16874,N_16048,N_16167);
or U16875 (N_16875,N_16350,N_16013);
nand U16876 (N_16876,N_16369,N_16052);
and U16877 (N_16877,N_16446,N_16168);
or U16878 (N_16878,N_16465,N_16474);
nand U16879 (N_16879,N_16205,N_16080);
nand U16880 (N_16880,N_16368,N_16292);
nand U16881 (N_16881,N_16226,N_16353);
nor U16882 (N_16882,N_16394,N_16196);
or U16883 (N_16883,N_16200,N_16494);
xnor U16884 (N_16884,N_16363,N_16164);
and U16885 (N_16885,N_16296,N_16321);
and U16886 (N_16886,N_16324,N_16001);
or U16887 (N_16887,N_16010,N_16107);
nor U16888 (N_16888,N_16059,N_16004);
nand U16889 (N_16889,N_16015,N_16283);
and U16890 (N_16890,N_16490,N_16171);
nand U16891 (N_16891,N_16134,N_16275);
or U16892 (N_16892,N_16275,N_16477);
and U16893 (N_16893,N_16212,N_16039);
nand U16894 (N_16894,N_16407,N_16354);
xor U16895 (N_16895,N_16111,N_16202);
and U16896 (N_16896,N_16301,N_16084);
nand U16897 (N_16897,N_16082,N_16156);
nor U16898 (N_16898,N_16303,N_16146);
nand U16899 (N_16899,N_16293,N_16042);
or U16900 (N_16900,N_16326,N_16324);
nand U16901 (N_16901,N_16214,N_16382);
or U16902 (N_16902,N_16383,N_16498);
nor U16903 (N_16903,N_16070,N_16012);
or U16904 (N_16904,N_16217,N_16305);
and U16905 (N_16905,N_16185,N_16427);
nand U16906 (N_16906,N_16209,N_16247);
nand U16907 (N_16907,N_16320,N_16196);
or U16908 (N_16908,N_16379,N_16470);
nor U16909 (N_16909,N_16485,N_16199);
nor U16910 (N_16910,N_16390,N_16357);
nor U16911 (N_16911,N_16487,N_16189);
nor U16912 (N_16912,N_16021,N_16296);
and U16913 (N_16913,N_16489,N_16105);
and U16914 (N_16914,N_16223,N_16032);
nor U16915 (N_16915,N_16002,N_16021);
nor U16916 (N_16916,N_16317,N_16444);
nor U16917 (N_16917,N_16046,N_16093);
or U16918 (N_16918,N_16453,N_16356);
and U16919 (N_16919,N_16426,N_16154);
nor U16920 (N_16920,N_16319,N_16436);
or U16921 (N_16921,N_16000,N_16265);
nand U16922 (N_16922,N_16053,N_16301);
or U16923 (N_16923,N_16173,N_16365);
nor U16924 (N_16924,N_16187,N_16169);
nor U16925 (N_16925,N_16316,N_16093);
or U16926 (N_16926,N_16214,N_16375);
and U16927 (N_16927,N_16382,N_16035);
or U16928 (N_16928,N_16385,N_16335);
nand U16929 (N_16929,N_16007,N_16354);
nor U16930 (N_16930,N_16004,N_16172);
nor U16931 (N_16931,N_16037,N_16364);
xor U16932 (N_16932,N_16333,N_16499);
or U16933 (N_16933,N_16259,N_16076);
or U16934 (N_16934,N_16179,N_16191);
or U16935 (N_16935,N_16287,N_16235);
nor U16936 (N_16936,N_16419,N_16312);
nand U16937 (N_16937,N_16162,N_16104);
and U16938 (N_16938,N_16197,N_16203);
or U16939 (N_16939,N_16326,N_16342);
nor U16940 (N_16940,N_16372,N_16109);
and U16941 (N_16941,N_16070,N_16428);
or U16942 (N_16942,N_16441,N_16422);
and U16943 (N_16943,N_16028,N_16073);
nand U16944 (N_16944,N_16059,N_16322);
nand U16945 (N_16945,N_16178,N_16149);
and U16946 (N_16946,N_16482,N_16142);
nand U16947 (N_16947,N_16060,N_16320);
nor U16948 (N_16948,N_16324,N_16122);
nand U16949 (N_16949,N_16035,N_16147);
or U16950 (N_16950,N_16396,N_16274);
nand U16951 (N_16951,N_16298,N_16100);
nand U16952 (N_16952,N_16324,N_16394);
and U16953 (N_16953,N_16191,N_16426);
nor U16954 (N_16954,N_16144,N_16134);
or U16955 (N_16955,N_16435,N_16265);
nor U16956 (N_16956,N_16363,N_16394);
nor U16957 (N_16957,N_16102,N_16115);
and U16958 (N_16958,N_16144,N_16101);
nand U16959 (N_16959,N_16170,N_16129);
or U16960 (N_16960,N_16442,N_16087);
and U16961 (N_16961,N_16364,N_16341);
nand U16962 (N_16962,N_16041,N_16419);
and U16963 (N_16963,N_16090,N_16037);
nand U16964 (N_16964,N_16046,N_16120);
or U16965 (N_16965,N_16033,N_16106);
nor U16966 (N_16966,N_16092,N_16122);
or U16967 (N_16967,N_16133,N_16432);
and U16968 (N_16968,N_16173,N_16318);
and U16969 (N_16969,N_16255,N_16264);
or U16970 (N_16970,N_16343,N_16346);
nor U16971 (N_16971,N_16176,N_16056);
nor U16972 (N_16972,N_16159,N_16331);
and U16973 (N_16973,N_16397,N_16039);
nand U16974 (N_16974,N_16426,N_16410);
xnor U16975 (N_16975,N_16320,N_16084);
or U16976 (N_16976,N_16439,N_16319);
nor U16977 (N_16977,N_16165,N_16422);
or U16978 (N_16978,N_16347,N_16400);
nand U16979 (N_16979,N_16103,N_16059);
nand U16980 (N_16980,N_16282,N_16323);
nand U16981 (N_16981,N_16481,N_16321);
and U16982 (N_16982,N_16021,N_16095);
or U16983 (N_16983,N_16119,N_16084);
or U16984 (N_16984,N_16223,N_16121);
nor U16985 (N_16985,N_16044,N_16034);
nand U16986 (N_16986,N_16291,N_16270);
and U16987 (N_16987,N_16009,N_16099);
or U16988 (N_16988,N_16157,N_16202);
and U16989 (N_16989,N_16030,N_16310);
or U16990 (N_16990,N_16006,N_16351);
or U16991 (N_16991,N_16023,N_16081);
nand U16992 (N_16992,N_16422,N_16175);
and U16993 (N_16993,N_16406,N_16443);
nor U16994 (N_16994,N_16204,N_16066);
nand U16995 (N_16995,N_16384,N_16171);
or U16996 (N_16996,N_16095,N_16213);
and U16997 (N_16997,N_16141,N_16483);
or U16998 (N_16998,N_16384,N_16449);
nand U16999 (N_16999,N_16135,N_16074);
nand U17000 (N_17000,N_16511,N_16751);
nand U17001 (N_17001,N_16505,N_16647);
nand U17002 (N_17002,N_16825,N_16772);
nand U17003 (N_17003,N_16895,N_16946);
nor U17004 (N_17004,N_16595,N_16676);
nand U17005 (N_17005,N_16904,N_16761);
or U17006 (N_17006,N_16737,N_16528);
or U17007 (N_17007,N_16576,N_16951);
nor U17008 (N_17008,N_16715,N_16679);
nor U17009 (N_17009,N_16801,N_16985);
or U17010 (N_17010,N_16845,N_16780);
or U17011 (N_17011,N_16953,N_16609);
nor U17012 (N_17012,N_16673,N_16902);
and U17013 (N_17013,N_16981,N_16894);
nor U17014 (N_17014,N_16945,N_16515);
and U17015 (N_17015,N_16674,N_16596);
nor U17016 (N_17016,N_16608,N_16557);
nand U17017 (N_17017,N_16814,N_16849);
nor U17018 (N_17018,N_16886,N_16513);
nor U17019 (N_17019,N_16549,N_16732);
and U17020 (N_17020,N_16962,N_16618);
nand U17021 (N_17021,N_16575,N_16767);
nor U17022 (N_17022,N_16977,N_16854);
or U17023 (N_17023,N_16968,N_16571);
and U17024 (N_17024,N_16824,N_16719);
nand U17025 (N_17025,N_16606,N_16592);
and U17026 (N_17026,N_16859,N_16873);
or U17027 (N_17027,N_16941,N_16760);
and U17028 (N_17028,N_16918,N_16632);
nor U17029 (N_17029,N_16857,N_16762);
xor U17030 (N_17030,N_16917,N_16909);
nor U17031 (N_17031,N_16774,N_16957);
and U17032 (N_17032,N_16795,N_16562);
and U17033 (N_17033,N_16791,N_16856);
nor U17034 (N_17034,N_16623,N_16921);
nand U17035 (N_17035,N_16517,N_16599);
xnor U17036 (N_17036,N_16806,N_16874);
nand U17037 (N_17037,N_16919,N_16826);
nand U17038 (N_17038,N_16996,N_16912);
and U17039 (N_17039,N_16982,N_16882);
and U17040 (N_17040,N_16759,N_16703);
nand U17041 (N_17041,N_16850,N_16649);
and U17042 (N_17042,N_16847,N_16682);
and U17043 (N_17043,N_16510,N_16799);
nand U17044 (N_17044,N_16709,N_16600);
nor U17045 (N_17045,N_16666,N_16998);
or U17046 (N_17046,N_16949,N_16591);
or U17047 (N_17047,N_16524,N_16535);
and U17048 (N_17048,N_16546,N_16516);
or U17049 (N_17049,N_16586,N_16842);
nor U17050 (N_17050,N_16727,N_16852);
nor U17051 (N_17051,N_16626,N_16819);
nand U17052 (N_17052,N_16785,N_16580);
nor U17053 (N_17053,N_16537,N_16602);
or U17054 (N_17054,N_16613,N_16698);
nand U17055 (N_17055,N_16790,N_16956);
nand U17056 (N_17056,N_16520,N_16988);
nor U17057 (N_17057,N_16925,N_16574);
and U17058 (N_17058,N_16955,N_16533);
and U17059 (N_17059,N_16696,N_16853);
nand U17060 (N_17060,N_16697,N_16783);
nand U17061 (N_17061,N_16634,N_16743);
nand U17062 (N_17062,N_16648,N_16621);
nor U17063 (N_17063,N_16619,N_16633);
nand U17064 (N_17064,N_16514,N_16866);
and U17065 (N_17065,N_16663,N_16542);
or U17066 (N_17066,N_16989,N_16833);
nor U17067 (N_17067,N_16758,N_16942);
nand U17068 (N_17068,N_16802,N_16637);
and U17069 (N_17069,N_16792,N_16526);
and U17070 (N_17070,N_16813,N_16865);
and U17071 (N_17071,N_16552,N_16640);
or U17072 (N_17072,N_16950,N_16808);
nand U17073 (N_17073,N_16993,N_16502);
nor U17074 (N_17074,N_16876,N_16501);
nor U17075 (N_17075,N_16610,N_16999);
nand U17076 (N_17076,N_16724,N_16539);
nand U17077 (N_17077,N_16601,N_16954);
nand U17078 (N_17078,N_16581,N_16922);
or U17079 (N_17079,N_16641,N_16923);
nand U17080 (N_17080,N_16573,N_16887);
nor U17081 (N_17081,N_16689,N_16839);
nor U17082 (N_17082,N_16965,N_16797);
or U17083 (N_17083,N_16820,N_16810);
or U17084 (N_17084,N_16629,N_16734);
nor U17085 (N_17085,N_16771,N_16594);
nand U17086 (N_17086,N_16855,N_16749);
nor U17087 (N_17087,N_16607,N_16907);
and U17088 (N_17088,N_16544,N_16911);
nor U17089 (N_17089,N_16702,N_16821);
and U17090 (N_17090,N_16567,N_16714);
and U17091 (N_17091,N_16670,N_16585);
or U17092 (N_17092,N_16937,N_16652);
and U17093 (N_17093,N_16731,N_16775);
or U17094 (N_17094,N_16536,N_16800);
nand U17095 (N_17095,N_16718,N_16527);
nor U17096 (N_17096,N_16916,N_16947);
and U17097 (N_17097,N_16784,N_16672);
nor U17098 (N_17098,N_16915,N_16890);
and U17099 (N_17099,N_16952,N_16938);
or U17100 (N_17100,N_16617,N_16582);
and U17101 (N_17101,N_16995,N_16897);
or U17102 (N_17102,N_16973,N_16794);
nand U17103 (N_17103,N_16867,N_16862);
nor U17104 (N_17104,N_16570,N_16830);
nor U17105 (N_17105,N_16750,N_16803);
and U17106 (N_17106,N_16615,N_16929);
and U17107 (N_17107,N_16782,N_16644);
or U17108 (N_17108,N_16645,N_16503);
nand U17109 (N_17109,N_16778,N_16540);
nand U17110 (N_17110,N_16829,N_16638);
and U17111 (N_17111,N_16765,N_16597);
or U17112 (N_17112,N_16646,N_16881);
and U17113 (N_17113,N_16753,N_16693);
or U17114 (N_17114,N_16587,N_16675);
nand U17115 (N_17115,N_16726,N_16984);
nand U17116 (N_17116,N_16614,N_16875);
nand U17117 (N_17117,N_16566,N_16843);
or U17118 (N_17118,N_16690,N_16880);
and U17119 (N_17119,N_16891,N_16589);
or U17120 (N_17120,N_16500,N_16838);
nand U17121 (N_17121,N_16986,N_16688);
nand U17122 (N_17122,N_16553,N_16818);
nand U17123 (N_17123,N_16888,N_16969);
nand U17124 (N_17124,N_16654,N_16970);
and U17125 (N_17125,N_16521,N_16756);
and U17126 (N_17126,N_16620,N_16773);
nor U17127 (N_17127,N_16972,N_16992);
and U17128 (N_17128,N_16612,N_16844);
or U17129 (N_17129,N_16745,N_16899);
nor U17130 (N_17130,N_16705,N_16848);
or U17131 (N_17131,N_16694,N_16630);
and U17132 (N_17132,N_16691,N_16708);
nor U17133 (N_17133,N_16658,N_16669);
or U17134 (N_17134,N_16932,N_16828);
and U17135 (N_17135,N_16677,N_16757);
nand U17136 (N_17136,N_16752,N_16870);
and U17137 (N_17137,N_16523,N_16940);
nand U17138 (N_17138,N_16729,N_16628);
nand U17139 (N_17139,N_16643,N_16681);
or U17140 (N_17140,N_16754,N_16991);
or U17141 (N_17141,N_16701,N_16883);
nor U17142 (N_17142,N_16837,N_16590);
nand U17143 (N_17143,N_16508,N_16739);
and U17144 (N_17144,N_16685,N_16742);
or U17145 (N_17145,N_16851,N_16639);
and U17146 (N_17146,N_16979,N_16625);
and U17147 (N_17147,N_16990,N_16519);
nor U17148 (N_17148,N_16860,N_16559);
or U17149 (N_17149,N_16561,N_16678);
xor U17150 (N_17150,N_16730,N_16635);
or U17151 (N_17151,N_16588,N_16906);
xnor U17152 (N_17152,N_16766,N_16611);
and U17153 (N_17153,N_16958,N_16622);
nand U17154 (N_17154,N_16807,N_16728);
nor U17155 (N_17155,N_16636,N_16948);
nor U17156 (N_17156,N_16631,N_16547);
nand U17157 (N_17157,N_16717,N_16763);
nor U17158 (N_17158,N_16563,N_16746);
nor U17159 (N_17159,N_16869,N_16840);
and U17160 (N_17160,N_16683,N_16811);
or U17161 (N_17161,N_16748,N_16805);
nor U17162 (N_17162,N_16668,N_16740);
nand U17163 (N_17163,N_16931,N_16769);
or U17164 (N_17164,N_16879,N_16531);
nor U17165 (N_17165,N_16710,N_16905);
nand U17166 (N_17166,N_16841,N_16930);
or U17167 (N_17167,N_16723,N_16551);
nand U17168 (N_17168,N_16939,N_16827);
nand U17169 (N_17169,N_16720,N_16555);
or U17170 (N_17170,N_16661,N_16812);
and U17171 (N_17171,N_16779,N_16568);
nor U17172 (N_17172,N_16863,N_16987);
and U17173 (N_17173,N_16706,N_16983);
or U17174 (N_17174,N_16593,N_16506);
or U17175 (N_17175,N_16936,N_16616);
nand U17176 (N_17176,N_16660,N_16560);
nor U17177 (N_17177,N_16997,N_16796);
and U17178 (N_17178,N_16736,N_16770);
and U17179 (N_17179,N_16924,N_16603);
and U17180 (N_17180,N_16910,N_16572);
and U17181 (N_17181,N_16822,N_16789);
nor U17182 (N_17182,N_16781,N_16671);
nand U17183 (N_17183,N_16889,N_16550);
and U17184 (N_17184,N_16933,N_16605);
nor U17185 (N_17185,N_16898,N_16583);
or U17186 (N_17186,N_16878,N_16966);
or U17187 (N_17187,N_16926,N_16548);
nand U17188 (N_17188,N_16747,N_16712);
and U17189 (N_17189,N_16518,N_16959);
and U17190 (N_17190,N_16964,N_16655);
or U17191 (N_17191,N_16901,N_16836);
nand U17192 (N_17192,N_16656,N_16816);
and U17193 (N_17193,N_16725,N_16764);
or U17194 (N_17194,N_16787,N_16651);
nand U17195 (N_17195,N_16864,N_16687);
or U17196 (N_17196,N_16963,N_16809);
nor U17197 (N_17197,N_16961,N_16529);
nor U17198 (N_17198,N_16556,N_16768);
nand U17199 (N_17199,N_16699,N_16604);
nor U17200 (N_17200,N_16713,N_16545);
nor U17201 (N_17201,N_16735,N_16662);
or U17202 (N_17202,N_16707,N_16900);
nor U17203 (N_17203,N_16914,N_16716);
or U17204 (N_17204,N_16584,N_16700);
and U17205 (N_17205,N_16744,N_16692);
or U17206 (N_17206,N_16569,N_16884);
nor U17207 (N_17207,N_16832,N_16525);
xor U17208 (N_17208,N_16650,N_16565);
nand U17209 (N_17209,N_16834,N_16913);
nor U17210 (N_17210,N_16776,N_16578);
nand U17211 (N_17211,N_16903,N_16659);
nor U17212 (N_17212,N_16788,N_16579);
and U17213 (N_17213,N_16665,N_16543);
nand U17214 (N_17214,N_16846,N_16927);
nand U17215 (N_17215,N_16512,N_16877);
and U17216 (N_17216,N_16978,N_16893);
nand U17217 (N_17217,N_16695,N_16798);
nor U17218 (N_17218,N_16934,N_16928);
nand U17219 (N_17219,N_16975,N_16653);
nor U17220 (N_17220,N_16738,N_16598);
nor U17221 (N_17221,N_16509,N_16664);
nor U17222 (N_17222,N_16538,N_16667);
nand U17223 (N_17223,N_16704,N_16980);
or U17224 (N_17224,N_16960,N_16755);
or U17225 (N_17225,N_16892,N_16554);
nor U17226 (N_17226,N_16944,N_16534);
nand U17227 (N_17227,N_16680,N_16657);
and U17228 (N_17228,N_16721,N_16943);
and U17229 (N_17229,N_16530,N_16871);
or U17230 (N_17230,N_16967,N_16541);
and U17231 (N_17231,N_16815,N_16974);
nand U17232 (N_17232,N_16935,N_16831);
nor U17233 (N_17233,N_16564,N_16777);
and U17234 (N_17234,N_16722,N_16507);
or U17235 (N_17235,N_16624,N_16976);
or U17236 (N_17236,N_16896,N_16861);
and U17237 (N_17237,N_16741,N_16711);
and U17238 (N_17238,N_16872,N_16642);
or U17239 (N_17239,N_16627,N_16684);
nand U17240 (N_17240,N_16994,N_16804);
and U17241 (N_17241,N_16504,N_16817);
nand U17242 (N_17242,N_16686,N_16885);
nor U17243 (N_17243,N_16858,N_16971);
or U17244 (N_17244,N_16532,N_16793);
nor U17245 (N_17245,N_16868,N_16733);
nand U17246 (N_17246,N_16908,N_16558);
nand U17247 (N_17247,N_16577,N_16522);
and U17248 (N_17248,N_16823,N_16835);
nand U17249 (N_17249,N_16786,N_16920);
or U17250 (N_17250,N_16567,N_16606);
or U17251 (N_17251,N_16844,N_16831);
nand U17252 (N_17252,N_16529,N_16518);
nor U17253 (N_17253,N_16557,N_16520);
nor U17254 (N_17254,N_16897,N_16805);
nand U17255 (N_17255,N_16925,N_16803);
xnor U17256 (N_17256,N_16825,N_16609);
or U17257 (N_17257,N_16720,N_16544);
nand U17258 (N_17258,N_16550,N_16527);
or U17259 (N_17259,N_16694,N_16999);
or U17260 (N_17260,N_16702,N_16863);
or U17261 (N_17261,N_16660,N_16501);
nand U17262 (N_17262,N_16792,N_16936);
and U17263 (N_17263,N_16602,N_16553);
nand U17264 (N_17264,N_16967,N_16670);
nor U17265 (N_17265,N_16977,N_16682);
or U17266 (N_17266,N_16589,N_16652);
and U17267 (N_17267,N_16912,N_16927);
and U17268 (N_17268,N_16620,N_16991);
nor U17269 (N_17269,N_16515,N_16725);
and U17270 (N_17270,N_16532,N_16975);
nor U17271 (N_17271,N_16614,N_16976);
or U17272 (N_17272,N_16591,N_16682);
nor U17273 (N_17273,N_16753,N_16529);
or U17274 (N_17274,N_16597,N_16740);
and U17275 (N_17275,N_16981,N_16611);
nand U17276 (N_17276,N_16716,N_16834);
and U17277 (N_17277,N_16677,N_16903);
xnor U17278 (N_17278,N_16797,N_16932);
nand U17279 (N_17279,N_16790,N_16898);
nand U17280 (N_17280,N_16714,N_16893);
or U17281 (N_17281,N_16673,N_16520);
or U17282 (N_17282,N_16512,N_16933);
and U17283 (N_17283,N_16564,N_16510);
or U17284 (N_17284,N_16940,N_16879);
and U17285 (N_17285,N_16952,N_16633);
or U17286 (N_17286,N_16802,N_16849);
or U17287 (N_17287,N_16678,N_16581);
and U17288 (N_17288,N_16593,N_16842);
or U17289 (N_17289,N_16965,N_16808);
or U17290 (N_17290,N_16779,N_16989);
or U17291 (N_17291,N_16912,N_16668);
nand U17292 (N_17292,N_16908,N_16675);
or U17293 (N_17293,N_16581,N_16782);
xor U17294 (N_17294,N_16772,N_16823);
or U17295 (N_17295,N_16873,N_16590);
and U17296 (N_17296,N_16510,N_16548);
nor U17297 (N_17297,N_16799,N_16578);
nor U17298 (N_17298,N_16814,N_16769);
or U17299 (N_17299,N_16535,N_16843);
xnor U17300 (N_17300,N_16754,N_16713);
or U17301 (N_17301,N_16647,N_16664);
nand U17302 (N_17302,N_16980,N_16755);
nand U17303 (N_17303,N_16758,N_16979);
nor U17304 (N_17304,N_16658,N_16648);
and U17305 (N_17305,N_16994,N_16690);
or U17306 (N_17306,N_16531,N_16791);
and U17307 (N_17307,N_16561,N_16867);
nor U17308 (N_17308,N_16791,N_16544);
nand U17309 (N_17309,N_16771,N_16744);
xor U17310 (N_17310,N_16827,N_16840);
nor U17311 (N_17311,N_16999,N_16820);
or U17312 (N_17312,N_16724,N_16588);
and U17313 (N_17313,N_16648,N_16773);
nand U17314 (N_17314,N_16741,N_16937);
or U17315 (N_17315,N_16819,N_16750);
xor U17316 (N_17316,N_16672,N_16685);
nand U17317 (N_17317,N_16617,N_16686);
or U17318 (N_17318,N_16858,N_16502);
nand U17319 (N_17319,N_16588,N_16543);
nand U17320 (N_17320,N_16819,N_16915);
and U17321 (N_17321,N_16737,N_16927);
and U17322 (N_17322,N_16830,N_16654);
nand U17323 (N_17323,N_16920,N_16602);
or U17324 (N_17324,N_16829,N_16659);
nand U17325 (N_17325,N_16963,N_16724);
nor U17326 (N_17326,N_16513,N_16534);
nand U17327 (N_17327,N_16877,N_16625);
and U17328 (N_17328,N_16682,N_16921);
or U17329 (N_17329,N_16866,N_16533);
nand U17330 (N_17330,N_16758,N_16749);
nor U17331 (N_17331,N_16760,N_16834);
or U17332 (N_17332,N_16647,N_16864);
or U17333 (N_17333,N_16543,N_16605);
nand U17334 (N_17334,N_16728,N_16783);
nor U17335 (N_17335,N_16516,N_16949);
nor U17336 (N_17336,N_16716,N_16768);
or U17337 (N_17337,N_16881,N_16692);
nand U17338 (N_17338,N_16924,N_16578);
nand U17339 (N_17339,N_16855,N_16741);
nand U17340 (N_17340,N_16823,N_16962);
nor U17341 (N_17341,N_16916,N_16543);
or U17342 (N_17342,N_16947,N_16962);
and U17343 (N_17343,N_16536,N_16630);
and U17344 (N_17344,N_16662,N_16960);
nand U17345 (N_17345,N_16645,N_16738);
nor U17346 (N_17346,N_16580,N_16638);
and U17347 (N_17347,N_16661,N_16618);
or U17348 (N_17348,N_16985,N_16606);
and U17349 (N_17349,N_16968,N_16676);
and U17350 (N_17350,N_16596,N_16879);
nor U17351 (N_17351,N_16510,N_16682);
nand U17352 (N_17352,N_16875,N_16550);
nand U17353 (N_17353,N_16825,N_16604);
and U17354 (N_17354,N_16914,N_16861);
xor U17355 (N_17355,N_16759,N_16672);
or U17356 (N_17356,N_16715,N_16786);
nor U17357 (N_17357,N_16883,N_16816);
and U17358 (N_17358,N_16671,N_16582);
nand U17359 (N_17359,N_16814,N_16582);
nand U17360 (N_17360,N_16525,N_16875);
and U17361 (N_17361,N_16815,N_16515);
nor U17362 (N_17362,N_16819,N_16850);
nor U17363 (N_17363,N_16504,N_16532);
nor U17364 (N_17364,N_16606,N_16688);
or U17365 (N_17365,N_16786,N_16775);
and U17366 (N_17366,N_16528,N_16923);
or U17367 (N_17367,N_16923,N_16643);
or U17368 (N_17368,N_16970,N_16782);
or U17369 (N_17369,N_16574,N_16818);
and U17370 (N_17370,N_16983,N_16787);
or U17371 (N_17371,N_16908,N_16789);
or U17372 (N_17372,N_16737,N_16676);
or U17373 (N_17373,N_16809,N_16634);
and U17374 (N_17374,N_16977,N_16730);
nand U17375 (N_17375,N_16792,N_16985);
and U17376 (N_17376,N_16723,N_16648);
and U17377 (N_17377,N_16679,N_16814);
nor U17378 (N_17378,N_16823,N_16707);
and U17379 (N_17379,N_16547,N_16614);
and U17380 (N_17380,N_16805,N_16900);
and U17381 (N_17381,N_16597,N_16854);
nor U17382 (N_17382,N_16621,N_16670);
and U17383 (N_17383,N_16711,N_16873);
nand U17384 (N_17384,N_16753,N_16858);
nand U17385 (N_17385,N_16582,N_16881);
nand U17386 (N_17386,N_16575,N_16938);
nor U17387 (N_17387,N_16904,N_16628);
nand U17388 (N_17388,N_16767,N_16938);
or U17389 (N_17389,N_16704,N_16921);
nor U17390 (N_17390,N_16762,N_16615);
or U17391 (N_17391,N_16864,N_16554);
nand U17392 (N_17392,N_16629,N_16591);
xnor U17393 (N_17393,N_16632,N_16558);
nand U17394 (N_17394,N_16960,N_16979);
nand U17395 (N_17395,N_16651,N_16871);
nor U17396 (N_17396,N_16960,N_16831);
nor U17397 (N_17397,N_16764,N_16601);
and U17398 (N_17398,N_16519,N_16914);
and U17399 (N_17399,N_16711,N_16881);
and U17400 (N_17400,N_16747,N_16670);
or U17401 (N_17401,N_16530,N_16710);
nand U17402 (N_17402,N_16733,N_16831);
nor U17403 (N_17403,N_16512,N_16646);
nand U17404 (N_17404,N_16929,N_16962);
or U17405 (N_17405,N_16716,N_16703);
nor U17406 (N_17406,N_16832,N_16884);
or U17407 (N_17407,N_16859,N_16790);
nand U17408 (N_17408,N_16861,N_16821);
or U17409 (N_17409,N_16709,N_16529);
and U17410 (N_17410,N_16618,N_16969);
or U17411 (N_17411,N_16559,N_16597);
or U17412 (N_17412,N_16571,N_16627);
nor U17413 (N_17413,N_16784,N_16756);
or U17414 (N_17414,N_16568,N_16986);
nand U17415 (N_17415,N_16785,N_16867);
nand U17416 (N_17416,N_16711,N_16545);
nor U17417 (N_17417,N_16601,N_16930);
nand U17418 (N_17418,N_16509,N_16582);
and U17419 (N_17419,N_16505,N_16670);
or U17420 (N_17420,N_16572,N_16700);
nor U17421 (N_17421,N_16527,N_16758);
nor U17422 (N_17422,N_16876,N_16577);
or U17423 (N_17423,N_16823,N_16627);
nor U17424 (N_17424,N_16569,N_16574);
and U17425 (N_17425,N_16687,N_16781);
and U17426 (N_17426,N_16554,N_16511);
nand U17427 (N_17427,N_16742,N_16832);
and U17428 (N_17428,N_16502,N_16524);
nand U17429 (N_17429,N_16701,N_16923);
or U17430 (N_17430,N_16794,N_16525);
or U17431 (N_17431,N_16650,N_16940);
nand U17432 (N_17432,N_16812,N_16904);
nand U17433 (N_17433,N_16826,N_16816);
and U17434 (N_17434,N_16907,N_16944);
or U17435 (N_17435,N_16870,N_16706);
and U17436 (N_17436,N_16783,N_16729);
nand U17437 (N_17437,N_16922,N_16660);
xor U17438 (N_17438,N_16652,N_16565);
and U17439 (N_17439,N_16880,N_16702);
nand U17440 (N_17440,N_16687,N_16701);
and U17441 (N_17441,N_16860,N_16755);
nand U17442 (N_17442,N_16605,N_16844);
nand U17443 (N_17443,N_16648,N_16617);
nand U17444 (N_17444,N_16958,N_16603);
or U17445 (N_17445,N_16801,N_16683);
nand U17446 (N_17446,N_16539,N_16535);
or U17447 (N_17447,N_16756,N_16747);
xnor U17448 (N_17448,N_16668,N_16924);
or U17449 (N_17449,N_16683,N_16505);
and U17450 (N_17450,N_16797,N_16502);
nand U17451 (N_17451,N_16872,N_16944);
or U17452 (N_17452,N_16847,N_16628);
and U17453 (N_17453,N_16944,N_16814);
or U17454 (N_17454,N_16703,N_16556);
and U17455 (N_17455,N_16802,N_16602);
nand U17456 (N_17456,N_16828,N_16833);
or U17457 (N_17457,N_16598,N_16681);
nand U17458 (N_17458,N_16813,N_16636);
nor U17459 (N_17459,N_16778,N_16982);
nor U17460 (N_17460,N_16851,N_16798);
and U17461 (N_17461,N_16681,N_16845);
or U17462 (N_17462,N_16536,N_16549);
nor U17463 (N_17463,N_16964,N_16851);
or U17464 (N_17464,N_16774,N_16768);
nor U17465 (N_17465,N_16891,N_16657);
or U17466 (N_17466,N_16751,N_16545);
and U17467 (N_17467,N_16559,N_16766);
xnor U17468 (N_17468,N_16800,N_16750);
nor U17469 (N_17469,N_16926,N_16730);
nand U17470 (N_17470,N_16554,N_16831);
and U17471 (N_17471,N_16971,N_16610);
nor U17472 (N_17472,N_16771,N_16992);
or U17473 (N_17473,N_16857,N_16540);
nor U17474 (N_17474,N_16631,N_16894);
nand U17475 (N_17475,N_16972,N_16703);
or U17476 (N_17476,N_16905,N_16937);
and U17477 (N_17477,N_16668,N_16544);
nor U17478 (N_17478,N_16813,N_16812);
or U17479 (N_17479,N_16505,N_16964);
or U17480 (N_17480,N_16630,N_16515);
and U17481 (N_17481,N_16926,N_16957);
nand U17482 (N_17482,N_16915,N_16748);
xor U17483 (N_17483,N_16918,N_16662);
or U17484 (N_17484,N_16619,N_16614);
nand U17485 (N_17485,N_16924,N_16927);
and U17486 (N_17486,N_16872,N_16653);
nand U17487 (N_17487,N_16907,N_16515);
nor U17488 (N_17488,N_16793,N_16670);
nor U17489 (N_17489,N_16609,N_16596);
nand U17490 (N_17490,N_16596,N_16959);
nand U17491 (N_17491,N_16826,N_16708);
nand U17492 (N_17492,N_16793,N_16744);
nand U17493 (N_17493,N_16518,N_16687);
or U17494 (N_17494,N_16774,N_16941);
and U17495 (N_17495,N_16692,N_16983);
nor U17496 (N_17496,N_16733,N_16850);
nand U17497 (N_17497,N_16528,N_16537);
or U17498 (N_17498,N_16513,N_16825);
or U17499 (N_17499,N_16548,N_16506);
and U17500 (N_17500,N_17167,N_17083);
nand U17501 (N_17501,N_17307,N_17140);
and U17502 (N_17502,N_17225,N_17036);
or U17503 (N_17503,N_17175,N_17481);
nor U17504 (N_17504,N_17049,N_17238);
and U17505 (N_17505,N_17373,N_17475);
nand U17506 (N_17506,N_17054,N_17398);
and U17507 (N_17507,N_17113,N_17396);
or U17508 (N_17508,N_17151,N_17404);
nor U17509 (N_17509,N_17485,N_17025);
or U17510 (N_17510,N_17335,N_17244);
nand U17511 (N_17511,N_17114,N_17332);
and U17512 (N_17512,N_17435,N_17246);
or U17513 (N_17513,N_17407,N_17183);
nor U17514 (N_17514,N_17078,N_17008);
nor U17515 (N_17515,N_17436,N_17496);
nor U17516 (N_17516,N_17142,N_17339);
or U17517 (N_17517,N_17004,N_17141);
or U17518 (N_17518,N_17185,N_17173);
nand U17519 (N_17519,N_17372,N_17449);
nand U17520 (N_17520,N_17365,N_17383);
nand U17521 (N_17521,N_17128,N_17472);
nand U17522 (N_17522,N_17302,N_17013);
nor U17523 (N_17523,N_17095,N_17170);
and U17524 (N_17524,N_17423,N_17283);
nand U17525 (N_17525,N_17150,N_17099);
nor U17526 (N_17526,N_17438,N_17024);
nand U17527 (N_17527,N_17498,N_17295);
or U17528 (N_17528,N_17259,N_17038);
and U17529 (N_17529,N_17249,N_17409);
and U17530 (N_17530,N_17007,N_17367);
xnor U17531 (N_17531,N_17156,N_17251);
nand U17532 (N_17532,N_17416,N_17002);
and U17533 (N_17533,N_17480,N_17041);
xnor U17534 (N_17534,N_17417,N_17192);
nand U17535 (N_17535,N_17328,N_17021);
nand U17536 (N_17536,N_17040,N_17467);
nand U17537 (N_17537,N_17210,N_17027);
and U17538 (N_17538,N_17430,N_17270);
nand U17539 (N_17539,N_17403,N_17127);
and U17540 (N_17540,N_17331,N_17267);
and U17541 (N_17541,N_17499,N_17233);
or U17542 (N_17542,N_17048,N_17006);
nor U17543 (N_17543,N_17289,N_17291);
nor U17544 (N_17544,N_17317,N_17235);
or U17545 (N_17545,N_17236,N_17305);
and U17546 (N_17546,N_17342,N_17357);
xnor U17547 (N_17547,N_17091,N_17454);
or U17548 (N_17548,N_17477,N_17343);
nor U17549 (N_17549,N_17118,N_17319);
nand U17550 (N_17550,N_17483,N_17418);
nand U17551 (N_17551,N_17205,N_17217);
or U17552 (N_17552,N_17093,N_17152);
nand U17553 (N_17553,N_17463,N_17181);
xor U17554 (N_17554,N_17349,N_17277);
or U17555 (N_17555,N_17077,N_17355);
or U17556 (N_17556,N_17195,N_17257);
nand U17557 (N_17557,N_17088,N_17344);
and U17558 (N_17558,N_17326,N_17161);
nor U17559 (N_17559,N_17374,N_17473);
nand U17560 (N_17560,N_17209,N_17309);
xor U17561 (N_17561,N_17206,N_17442);
or U17562 (N_17562,N_17107,N_17378);
and U17563 (N_17563,N_17452,N_17354);
nor U17564 (N_17564,N_17154,N_17018);
or U17565 (N_17565,N_17338,N_17346);
nand U17566 (N_17566,N_17164,N_17063);
nand U17567 (N_17567,N_17056,N_17102);
or U17568 (N_17568,N_17275,N_17433);
nand U17569 (N_17569,N_17484,N_17062);
nand U17570 (N_17570,N_17379,N_17458);
nor U17571 (N_17571,N_17058,N_17068);
and U17572 (N_17572,N_17368,N_17071);
and U17573 (N_17573,N_17286,N_17239);
nand U17574 (N_17574,N_17492,N_17352);
nor U17575 (N_17575,N_17258,N_17031);
nand U17576 (N_17576,N_17268,N_17123);
nor U17577 (N_17577,N_17131,N_17191);
or U17578 (N_17578,N_17104,N_17139);
and U17579 (N_17579,N_17474,N_17412);
nor U17580 (N_17580,N_17171,N_17026);
nand U17581 (N_17581,N_17124,N_17086);
nor U17582 (N_17582,N_17199,N_17260);
nor U17583 (N_17583,N_17380,N_17432);
or U17584 (N_17584,N_17098,N_17079);
and U17585 (N_17585,N_17136,N_17293);
nand U17586 (N_17586,N_17495,N_17120);
nand U17587 (N_17587,N_17304,N_17299);
and U17588 (N_17588,N_17450,N_17177);
or U17589 (N_17589,N_17096,N_17262);
nor U17590 (N_17590,N_17321,N_17172);
nand U17591 (N_17591,N_17301,N_17497);
or U17592 (N_17592,N_17166,N_17147);
or U17593 (N_17593,N_17457,N_17197);
nor U17594 (N_17594,N_17400,N_17392);
nand U17595 (N_17595,N_17073,N_17381);
or U17596 (N_17596,N_17419,N_17245);
or U17597 (N_17597,N_17255,N_17070);
or U17598 (N_17598,N_17146,N_17320);
nor U17599 (N_17599,N_17316,N_17133);
nand U17600 (N_17600,N_17462,N_17300);
and U17601 (N_17601,N_17471,N_17389);
or U17602 (N_17602,N_17247,N_17461);
nor U17603 (N_17603,N_17313,N_17334);
nor U17604 (N_17604,N_17491,N_17216);
nor U17605 (N_17605,N_17288,N_17388);
nor U17606 (N_17606,N_17405,N_17280);
or U17607 (N_17607,N_17137,N_17263);
nor U17608 (N_17608,N_17399,N_17353);
or U17609 (N_17609,N_17122,N_17310);
nand U17610 (N_17610,N_17090,N_17193);
or U17611 (N_17611,N_17459,N_17108);
and U17612 (N_17612,N_17250,N_17092);
nor U17613 (N_17613,N_17134,N_17384);
or U17614 (N_17614,N_17112,N_17318);
nor U17615 (N_17615,N_17431,N_17001);
or U17616 (N_17616,N_17284,N_17356);
nand U17617 (N_17617,N_17377,N_17067);
nand U17618 (N_17618,N_17162,N_17272);
xnor U17619 (N_17619,N_17012,N_17014);
nor U17620 (N_17620,N_17248,N_17351);
and U17621 (N_17621,N_17408,N_17478);
and U17622 (N_17622,N_17045,N_17149);
nand U17623 (N_17623,N_17411,N_17460);
nor U17624 (N_17624,N_17315,N_17348);
nor U17625 (N_17625,N_17016,N_17111);
and U17626 (N_17626,N_17047,N_17052);
nor U17627 (N_17627,N_17213,N_17240);
xor U17628 (N_17628,N_17469,N_17401);
and U17629 (N_17629,N_17022,N_17386);
xor U17630 (N_17630,N_17228,N_17479);
and U17631 (N_17631,N_17265,N_17311);
nand U17632 (N_17632,N_17116,N_17261);
nand U17633 (N_17633,N_17428,N_17103);
or U17634 (N_17634,N_17312,N_17229);
xor U17635 (N_17635,N_17451,N_17034);
or U17636 (N_17636,N_17153,N_17276);
or U17637 (N_17637,N_17361,N_17358);
nor U17638 (N_17638,N_17144,N_17187);
nor U17639 (N_17639,N_17444,N_17194);
or U17640 (N_17640,N_17069,N_17363);
nor U17641 (N_17641,N_17220,N_17176);
and U17642 (N_17642,N_17287,N_17360);
and U17643 (N_17643,N_17490,N_17097);
nand U17644 (N_17644,N_17044,N_17223);
or U17645 (N_17645,N_17132,N_17129);
and U17646 (N_17646,N_17443,N_17466);
and U17647 (N_17647,N_17105,N_17336);
or U17648 (N_17648,N_17340,N_17028);
or U17649 (N_17649,N_17163,N_17121);
nor U17650 (N_17650,N_17215,N_17350);
and U17651 (N_17651,N_17084,N_17035);
nor U17652 (N_17652,N_17030,N_17230);
and U17653 (N_17653,N_17415,N_17057);
nor U17654 (N_17654,N_17437,N_17135);
nand U17655 (N_17655,N_17019,N_17470);
and U17656 (N_17656,N_17370,N_17003);
and U17657 (N_17657,N_17159,N_17204);
nor U17658 (N_17658,N_17441,N_17157);
nand U17659 (N_17659,N_17371,N_17333);
and U17660 (N_17660,N_17375,N_17202);
or U17661 (N_17661,N_17075,N_17476);
and U17662 (N_17662,N_17385,N_17314);
and U17663 (N_17663,N_17115,N_17242);
nand U17664 (N_17664,N_17222,N_17281);
nor U17665 (N_17665,N_17487,N_17017);
nand U17666 (N_17666,N_17414,N_17413);
nand U17667 (N_17667,N_17279,N_17042);
nor U17668 (N_17668,N_17168,N_17254);
nor U17669 (N_17669,N_17464,N_17190);
and U17670 (N_17670,N_17420,N_17237);
and U17671 (N_17671,N_17196,N_17143);
and U17672 (N_17672,N_17306,N_17180);
nor U17673 (N_17673,N_17234,N_17271);
and U17674 (N_17674,N_17110,N_17297);
or U17675 (N_17675,N_17488,N_17241);
nor U17676 (N_17676,N_17138,N_17422);
or U17677 (N_17677,N_17362,N_17406);
nor U17678 (N_17678,N_17119,N_17020);
nor U17679 (N_17679,N_17065,N_17082);
nand U17680 (N_17680,N_17252,N_17174);
and U17681 (N_17681,N_17325,N_17429);
and U17682 (N_17682,N_17369,N_17274);
xnor U17683 (N_17683,N_17072,N_17155);
nor U17684 (N_17684,N_17169,N_17201);
and U17685 (N_17685,N_17468,N_17125);
and U17686 (N_17686,N_17009,N_17226);
nor U17687 (N_17687,N_17402,N_17264);
or U17688 (N_17688,N_17298,N_17094);
or U17689 (N_17689,N_17043,N_17269);
or U17690 (N_17690,N_17189,N_17033);
nand U17691 (N_17691,N_17290,N_17382);
nand U17692 (N_17692,N_17029,N_17446);
and U17693 (N_17693,N_17482,N_17203);
or U17694 (N_17694,N_17032,N_17303);
xnor U17695 (N_17695,N_17145,N_17066);
or U17696 (N_17696,N_17278,N_17053);
nor U17697 (N_17697,N_17200,N_17076);
nand U17698 (N_17698,N_17158,N_17000);
or U17699 (N_17699,N_17089,N_17359);
or U17700 (N_17700,N_17327,N_17050);
or U17701 (N_17701,N_17051,N_17061);
and U17702 (N_17702,N_17243,N_17322);
nor U17703 (N_17703,N_17010,N_17330);
nand U17704 (N_17704,N_17323,N_17324);
or U17705 (N_17705,N_17465,N_17256);
nor U17706 (N_17706,N_17207,N_17296);
nand U17707 (N_17707,N_17366,N_17046);
nand U17708 (N_17708,N_17117,N_17080);
nand U17709 (N_17709,N_17101,N_17015);
and U17710 (N_17710,N_17221,N_17037);
nand U17711 (N_17711,N_17453,N_17393);
nand U17712 (N_17712,N_17188,N_17055);
nor U17713 (N_17713,N_17179,N_17039);
nor U17714 (N_17714,N_17178,N_17212);
or U17715 (N_17715,N_17160,N_17440);
or U17716 (N_17716,N_17345,N_17165);
or U17717 (N_17717,N_17285,N_17231);
nor U17718 (N_17718,N_17397,N_17266);
nand U17719 (N_17719,N_17456,N_17364);
and U17720 (N_17720,N_17198,N_17448);
or U17721 (N_17721,N_17494,N_17376);
and U17722 (N_17722,N_17074,N_17100);
xnor U17723 (N_17723,N_17391,N_17395);
nor U17724 (N_17724,N_17218,N_17493);
nand U17725 (N_17725,N_17329,N_17060);
or U17726 (N_17726,N_17421,N_17390);
and U17727 (N_17727,N_17253,N_17486);
nor U17728 (N_17728,N_17447,N_17148);
or U17729 (N_17729,N_17232,N_17059);
nand U17730 (N_17730,N_17341,N_17184);
or U17731 (N_17731,N_17219,N_17294);
nand U17732 (N_17732,N_17005,N_17394);
and U17733 (N_17733,N_17489,N_17337);
nand U17734 (N_17734,N_17273,N_17439);
and U17735 (N_17735,N_17011,N_17109);
or U17736 (N_17736,N_17455,N_17427);
and U17737 (N_17737,N_17387,N_17445);
or U17738 (N_17738,N_17410,N_17130);
and U17739 (N_17739,N_17282,N_17085);
or U17740 (N_17740,N_17426,N_17308);
nor U17741 (N_17741,N_17081,N_17434);
nand U17742 (N_17742,N_17208,N_17347);
nor U17743 (N_17743,N_17425,N_17214);
and U17744 (N_17744,N_17211,N_17292);
nor U17745 (N_17745,N_17224,N_17227);
and U17746 (N_17746,N_17106,N_17182);
or U17747 (N_17747,N_17186,N_17087);
xnor U17748 (N_17748,N_17023,N_17126);
nor U17749 (N_17749,N_17424,N_17064);
or U17750 (N_17750,N_17297,N_17244);
nand U17751 (N_17751,N_17322,N_17309);
and U17752 (N_17752,N_17148,N_17495);
or U17753 (N_17753,N_17334,N_17086);
nand U17754 (N_17754,N_17499,N_17282);
nand U17755 (N_17755,N_17167,N_17195);
or U17756 (N_17756,N_17450,N_17307);
or U17757 (N_17757,N_17450,N_17232);
or U17758 (N_17758,N_17066,N_17473);
or U17759 (N_17759,N_17065,N_17463);
or U17760 (N_17760,N_17226,N_17128);
nand U17761 (N_17761,N_17493,N_17313);
nand U17762 (N_17762,N_17304,N_17462);
xor U17763 (N_17763,N_17059,N_17482);
nor U17764 (N_17764,N_17090,N_17311);
nor U17765 (N_17765,N_17004,N_17306);
or U17766 (N_17766,N_17343,N_17286);
nor U17767 (N_17767,N_17370,N_17246);
or U17768 (N_17768,N_17152,N_17100);
nand U17769 (N_17769,N_17346,N_17480);
or U17770 (N_17770,N_17241,N_17360);
and U17771 (N_17771,N_17448,N_17164);
nor U17772 (N_17772,N_17133,N_17079);
nand U17773 (N_17773,N_17414,N_17348);
or U17774 (N_17774,N_17280,N_17162);
nor U17775 (N_17775,N_17120,N_17335);
or U17776 (N_17776,N_17158,N_17188);
or U17777 (N_17777,N_17498,N_17206);
nor U17778 (N_17778,N_17167,N_17175);
or U17779 (N_17779,N_17409,N_17150);
or U17780 (N_17780,N_17053,N_17184);
or U17781 (N_17781,N_17102,N_17224);
or U17782 (N_17782,N_17347,N_17233);
or U17783 (N_17783,N_17191,N_17372);
nor U17784 (N_17784,N_17141,N_17474);
nand U17785 (N_17785,N_17102,N_17407);
nand U17786 (N_17786,N_17348,N_17126);
or U17787 (N_17787,N_17398,N_17238);
nand U17788 (N_17788,N_17104,N_17398);
nand U17789 (N_17789,N_17309,N_17305);
nor U17790 (N_17790,N_17407,N_17453);
nand U17791 (N_17791,N_17128,N_17005);
and U17792 (N_17792,N_17351,N_17176);
and U17793 (N_17793,N_17429,N_17397);
and U17794 (N_17794,N_17382,N_17441);
nand U17795 (N_17795,N_17244,N_17395);
nand U17796 (N_17796,N_17481,N_17215);
or U17797 (N_17797,N_17473,N_17223);
nor U17798 (N_17798,N_17134,N_17195);
and U17799 (N_17799,N_17368,N_17329);
nor U17800 (N_17800,N_17096,N_17012);
nor U17801 (N_17801,N_17153,N_17332);
and U17802 (N_17802,N_17050,N_17104);
or U17803 (N_17803,N_17184,N_17370);
nor U17804 (N_17804,N_17451,N_17271);
xnor U17805 (N_17805,N_17109,N_17376);
nor U17806 (N_17806,N_17158,N_17250);
or U17807 (N_17807,N_17276,N_17101);
nand U17808 (N_17808,N_17158,N_17474);
nor U17809 (N_17809,N_17397,N_17405);
or U17810 (N_17810,N_17458,N_17030);
nand U17811 (N_17811,N_17179,N_17488);
nand U17812 (N_17812,N_17422,N_17143);
or U17813 (N_17813,N_17302,N_17069);
or U17814 (N_17814,N_17372,N_17087);
or U17815 (N_17815,N_17445,N_17006);
and U17816 (N_17816,N_17479,N_17233);
nand U17817 (N_17817,N_17059,N_17475);
and U17818 (N_17818,N_17012,N_17160);
and U17819 (N_17819,N_17092,N_17131);
or U17820 (N_17820,N_17255,N_17413);
or U17821 (N_17821,N_17016,N_17487);
nand U17822 (N_17822,N_17292,N_17145);
or U17823 (N_17823,N_17056,N_17320);
or U17824 (N_17824,N_17366,N_17254);
nand U17825 (N_17825,N_17047,N_17451);
xor U17826 (N_17826,N_17347,N_17061);
or U17827 (N_17827,N_17463,N_17323);
and U17828 (N_17828,N_17119,N_17459);
or U17829 (N_17829,N_17313,N_17224);
nand U17830 (N_17830,N_17280,N_17432);
or U17831 (N_17831,N_17480,N_17263);
nor U17832 (N_17832,N_17401,N_17021);
nor U17833 (N_17833,N_17043,N_17042);
or U17834 (N_17834,N_17112,N_17107);
and U17835 (N_17835,N_17370,N_17373);
nor U17836 (N_17836,N_17383,N_17290);
nand U17837 (N_17837,N_17323,N_17363);
or U17838 (N_17838,N_17364,N_17308);
nand U17839 (N_17839,N_17286,N_17169);
nor U17840 (N_17840,N_17303,N_17409);
and U17841 (N_17841,N_17199,N_17335);
nor U17842 (N_17842,N_17234,N_17214);
and U17843 (N_17843,N_17285,N_17062);
nor U17844 (N_17844,N_17346,N_17395);
nor U17845 (N_17845,N_17488,N_17315);
nor U17846 (N_17846,N_17223,N_17432);
or U17847 (N_17847,N_17452,N_17272);
nor U17848 (N_17848,N_17342,N_17126);
or U17849 (N_17849,N_17204,N_17143);
or U17850 (N_17850,N_17488,N_17189);
nor U17851 (N_17851,N_17221,N_17373);
nand U17852 (N_17852,N_17112,N_17218);
and U17853 (N_17853,N_17111,N_17457);
or U17854 (N_17854,N_17405,N_17191);
nor U17855 (N_17855,N_17329,N_17325);
nand U17856 (N_17856,N_17233,N_17340);
or U17857 (N_17857,N_17356,N_17226);
or U17858 (N_17858,N_17325,N_17307);
nor U17859 (N_17859,N_17098,N_17081);
nor U17860 (N_17860,N_17309,N_17490);
nor U17861 (N_17861,N_17204,N_17141);
nand U17862 (N_17862,N_17222,N_17100);
and U17863 (N_17863,N_17217,N_17279);
or U17864 (N_17864,N_17106,N_17418);
nor U17865 (N_17865,N_17048,N_17148);
nor U17866 (N_17866,N_17071,N_17187);
nand U17867 (N_17867,N_17044,N_17162);
and U17868 (N_17868,N_17130,N_17463);
nor U17869 (N_17869,N_17132,N_17326);
or U17870 (N_17870,N_17285,N_17102);
nor U17871 (N_17871,N_17034,N_17190);
or U17872 (N_17872,N_17043,N_17253);
and U17873 (N_17873,N_17430,N_17414);
or U17874 (N_17874,N_17129,N_17378);
and U17875 (N_17875,N_17397,N_17379);
and U17876 (N_17876,N_17337,N_17371);
and U17877 (N_17877,N_17182,N_17285);
and U17878 (N_17878,N_17226,N_17419);
and U17879 (N_17879,N_17064,N_17040);
and U17880 (N_17880,N_17364,N_17088);
and U17881 (N_17881,N_17282,N_17020);
or U17882 (N_17882,N_17271,N_17099);
nand U17883 (N_17883,N_17426,N_17311);
or U17884 (N_17884,N_17366,N_17275);
nor U17885 (N_17885,N_17272,N_17252);
nand U17886 (N_17886,N_17101,N_17046);
and U17887 (N_17887,N_17490,N_17305);
nand U17888 (N_17888,N_17205,N_17224);
nand U17889 (N_17889,N_17130,N_17269);
and U17890 (N_17890,N_17025,N_17261);
and U17891 (N_17891,N_17020,N_17322);
nor U17892 (N_17892,N_17342,N_17068);
nand U17893 (N_17893,N_17093,N_17192);
and U17894 (N_17894,N_17381,N_17242);
and U17895 (N_17895,N_17186,N_17258);
nand U17896 (N_17896,N_17441,N_17189);
xor U17897 (N_17897,N_17275,N_17249);
or U17898 (N_17898,N_17207,N_17295);
or U17899 (N_17899,N_17473,N_17046);
or U17900 (N_17900,N_17218,N_17262);
or U17901 (N_17901,N_17338,N_17383);
and U17902 (N_17902,N_17424,N_17072);
nand U17903 (N_17903,N_17382,N_17153);
and U17904 (N_17904,N_17370,N_17015);
nor U17905 (N_17905,N_17067,N_17499);
and U17906 (N_17906,N_17070,N_17065);
and U17907 (N_17907,N_17388,N_17033);
nor U17908 (N_17908,N_17202,N_17355);
or U17909 (N_17909,N_17278,N_17113);
and U17910 (N_17910,N_17255,N_17273);
xor U17911 (N_17911,N_17382,N_17363);
xnor U17912 (N_17912,N_17174,N_17220);
nor U17913 (N_17913,N_17320,N_17343);
nand U17914 (N_17914,N_17007,N_17478);
nor U17915 (N_17915,N_17015,N_17035);
and U17916 (N_17916,N_17416,N_17478);
or U17917 (N_17917,N_17219,N_17317);
nand U17918 (N_17918,N_17409,N_17256);
nor U17919 (N_17919,N_17085,N_17136);
and U17920 (N_17920,N_17190,N_17195);
nor U17921 (N_17921,N_17056,N_17259);
nor U17922 (N_17922,N_17390,N_17112);
and U17923 (N_17923,N_17102,N_17359);
or U17924 (N_17924,N_17465,N_17121);
or U17925 (N_17925,N_17390,N_17228);
nor U17926 (N_17926,N_17475,N_17129);
nand U17927 (N_17927,N_17056,N_17453);
or U17928 (N_17928,N_17360,N_17094);
nor U17929 (N_17929,N_17126,N_17015);
or U17930 (N_17930,N_17206,N_17414);
or U17931 (N_17931,N_17284,N_17229);
nor U17932 (N_17932,N_17405,N_17052);
nor U17933 (N_17933,N_17371,N_17087);
nand U17934 (N_17934,N_17277,N_17299);
nand U17935 (N_17935,N_17475,N_17124);
and U17936 (N_17936,N_17198,N_17457);
and U17937 (N_17937,N_17310,N_17037);
and U17938 (N_17938,N_17297,N_17081);
nor U17939 (N_17939,N_17423,N_17178);
nor U17940 (N_17940,N_17449,N_17436);
nor U17941 (N_17941,N_17052,N_17026);
or U17942 (N_17942,N_17087,N_17069);
nor U17943 (N_17943,N_17343,N_17354);
and U17944 (N_17944,N_17040,N_17268);
and U17945 (N_17945,N_17337,N_17017);
or U17946 (N_17946,N_17113,N_17182);
and U17947 (N_17947,N_17017,N_17449);
or U17948 (N_17948,N_17402,N_17406);
nor U17949 (N_17949,N_17393,N_17288);
nor U17950 (N_17950,N_17492,N_17423);
nand U17951 (N_17951,N_17143,N_17002);
or U17952 (N_17952,N_17295,N_17322);
or U17953 (N_17953,N_17265,N_17068);
nand U17954 (N_17954,N_17465,N_17217);
nor U17955 (N_17955,N_17092,N_17231);
and U17956 (N_17956,N_17372,N_17444);
and U17957 (N_17957,N_17123,N_17187);
or U17958 (N_17958,N_17072,N_17430);
nand U17959 (N_17959,N_17394,N_17176);
nand U17960 (N_17960,N_17062,N_17037);
nor U17961 (N_17961,N_17450,N_17166);
nand U17962 (N_17962,N_17479,N_17213);
nor U17963 (N_17963,N_17161,N_17208);
and U17964 (N_17964,N_17309,N_17484);
and U17965 (N_17965,N_17152,N_17321);
or U17966 (N_17966,N_17272,N_17176);
nor U17967 (N_17967,N_17116,N_17013);
nor U17968 (N_17968,N_17320,N_17319);
nand U17969 (N_17969,N_17481,N_17427);
or U17970 (N_17970,N_17392,N_17237);
or U17971 (N_17971,N_17008,N_17225);
or U17972 (N_17972,N_17086,N_17176);
nand U17973 (N_17973,N_17279,N_17340);
or U17974 (N_17974,N_17387,N_17075);
or U17975 (N_17975,N_17403,N_17097);
nand U17976 (N_17976,N_17298,N_17172);
or U17977 (N_17977,N_17364,N_17421);
and U17978 (N_17978,N_17182,N_17313);
nor U17979 (N_17979,N_17351,N_17267);
nand U17980 (N_17980,N_17152,N_17245);
and U17981 (N_17981,N_17420,N_17062);
nand U17982 (N_17982,N_17355,N_17126);
nor U17983 (N_17983,N_17227,N_17125);
nand U17984 (N_17984,N_17498,N_17009);
or U17985 (N_17985,N_17343,N_17402);
nand U17986 (N_17986,N_17398,N_17018);
nor U17987 (N_17987,N_17263,N_17256);
xor U17988 (N_17988,N_17423,N_17124);
or U17989 (N_17989,N_17264,N_17051);
nor U17990 (N_17990,N_17437,N_17196);
nor U17991 (N_17991,N_17253,N_17372);
and U17992 (N_17992,N_17128,N_17320);
nor U17993 (N_17993,N_17130,N_17403);
nand U17994 (N_17994,N_17050,N_17499);
nand U17995 (N_17995,N_17458,N_17115);
or U17996 (N_17996,N_17181,N_17304);
nand U17997 (N_17997,N_17275,N_17331);
nand U17998 (N_17998,N_17392,N_17129);
and U17999 (N_17999,N_17355,N_17132);
or U18000 (N_18000,N_17729,N_17751);
nor U18001 (N_18001,N_17773,N_17667);
and U18002 (N_18002,N_17571,N_17700);
and U18003 (N_18003,N_17770,N_17607);
and U18004 (N_18004,N_17850,N_17831);
nand U18005 (N_18005,N_17643,N_17821);
and U18006 (N_18006,N_17576,N_17845);
nand U18007 (N_18007,N_17923,N_17570);
nor U18008 (N_18008,N_17691,N_17638);
nand U18009 (N_18009,N_17568,N_17893);
nand U18010 (N_18010,N_17901,N_17763);
nand U18011 (N_18011,N_17915,N_17745);
nor U18012 (N_18012,N_17945,N_17617);
nor U18013 (N_18013,N_17952,N_17659);
and U18014 (N_18014,N_17543,N_17723);
or U18015 (N_18015,N_17693,N_17741);
or U18016 (N_18016,N_17550,N_17514);
or U18017 (N_18017,N_17665,N_17602);
nor U18018 (N_18018,N_17728,N_17891);
nand U18019 (N_18019,N_17525,N_17979);
nand U18020 (N_18020,N_17683,N_17623);
nand U18021 (N_18021,N_17881,N_17661);
nor U18022 (N_18022,N_17895,N_17603);
nand U18023 (N_18023,N_17758,N_17557);
and U18024 (N_18024,N_17523,N_17605);
and U18025 (N_18025,N_17775,N_17957);
and U18026 (N_18026,N_17714,N_17584);
nor U18027 (N_18027,N_17960,N_17708);
and U18028 (N_18028,N_17731,N_17580);
and U18029 (N_18029,N_17890,N_17826);
or U18030 (N_18030,N_17833,N_17879);
nor U18031 (N_18031,N_17767,N_17518);
and U18032 (N_18032,N_17882,N_17972);
nand U18033 (N_18033,N_17897,N_17639);
nor U18034 (N_18034,N_17760,N_17990);
xor U18035 (N_18035,N_17809,N_17779);
nand U18036 (N_18036,N_17725,N_17613);
and U18037 (N_18037,N_17694,N_17836);
nand U18038 (N_18038,N_17991,N_17733);
nand U18039 (N_18039,N_17718,N_17766);
nand U18040 (N_18040,N_17963,N_17815);
nor U18041 (N_18041,N_17579,N_17581);
or U18042 (N_18042,N_17712,N_17762);
nor U18043 (N_18043,N_17740,N_17630);
and U18044 (N_18044,N_17716,N_17511);
and U18045 (N_18045,N_17596,N_17983);
nand U18046 (N_18046,N_17540,N_17704);
and U18047 (N_18047,N_17549,N_17526);
or U18048 (N_18048,N_17778,N_17572);
nand U18049 (N_18049,N_17547,N_17995);
nand U18050 (N_18050,N_17675,N_17791);
and U18051 (N_18051,N_17840,N_17843);
nand U18052 (N_18052,N_17590,N_17757);
nand U18053 (N_18053,N_17565,N_17934);
nor U18054 (N_18054,N_17922,N_17832);
xnor U18055 (N_18055,N_17858,N_17848);
or U18056 (N_18056,N_17907,N_17631);
nand U18057 (N_18057,N_17695,N_17561);
nor U18058 (N_18058,N_17905,N_17515);
or U18059 (N_18059,N_17618,N_17956);
and U18060 (N_18060,N_17721,N_17827);
nor U18061 (N_18061,N_17797,N_17994);
nor U18062 (N_18062,N_17755,N_17806);
or U18063 (N_18063,N_17567,N_17984);
xor U18064 (N_18064,N_17982,N_17824);
nor U18065 (N_18065,N_17899,N_17706);
or U18066 (N_18066,N_17955,N_17688);
or U18067 (N_18067,N_17577,N_17864);
nor U18068 (N_18068,N_17900,N_17552);
nor U18069 (N_18069,N_17867,N_17535);
xnor U18070 (N_18070,N_17961,N_17985);
nand U18071 (N_18071,N_17980,N_17774);
nand U18072 (N_18072,N_17847,N_17641);
nor U18073 (N_18073,N_17671,N_17647);
nand U18074 (N_18074,N_17692,N_17871);
and U18075 (N_18075,N_17932,N_17971);
xor U18076 (N_18076,N_17750,N_17844);
nand U18077 (N_18077,N_17697,N_17823);
or U18078 (N_18078,N_17591,N_17841);
nor U18079 (N_18079,N_17888,N_17612);
nor U18080 (N_18080,N_17663,N_17852);
nor U18081 (N_18081,N_17820,N_17886);
nand U18082 (N_18082,N_17735,N_17742);
nand U18083 (N_18083,N_17789,N_17884);
nor U18084 (N_18084,N_17545,N_17551);
nor U18085 (N_18085,N_17539,N_17648);
or U18086 (N_18086,N_17861,N_17673);
and U18087 (N_18087,N_17566,N_17800);
nand U18088 (N_18088,N_17918,N_17593);
nor U18089 (N_18089,N_17805,N_17719);
nand U18090 (N_18090,N_17606,N_17958);
or U18091 (N_18091,N_17794,N_17803);
nor U18092 (N_18092,N_17516,N_17811);
or U18093 (N_18093,N_17658,N_17621);
nor U18094 (N_18094,N_17573,N_17996);
nand U18095 (N_18095,N_17869,N_17894);
nand U18096 (N_18096,N_17676,N_17578);
nand U18097 (N_18097,N_17660,N_17669);
nand U18098 (N_18098,N_17699,N_17720);
and U18099 (N_18099,N_17702,N_17501);
or U18100 (N_18100,N_17634,N_17816);
nor U18101 (N_18101,N_17672,N_17970);
nor U18102 (N_18102,N_17530,N_17834);
and U18103 (N_18103,N_17711,N_17998);
nor U18104 (N_18104,N_17968,N_17622);
or U18105 (N_18105,N_17781,N_17744);
nand U18106 (N_18106,N_17785,N_17737);
or U18107 (N_18107,N_17813,N_17768);
nor U18108 (N_18108,N_17788,N_17657);
and U18109 (N_18109,N_17722,N_17940);
or U18110 (N_18110,N_17862,N_17769);
or U18111 (N_18111,N_17949,N_17527);
nor U18112 (N_18112,N_17628,N_17795);
and U18113 (N_18113,N_17954,N_17609);
or U18114 (N_18114,N_17504,N_17541);
nor U18115 (N_18115,N_17965,N_17889);
nand U18116 (N_18116,N_17611,N_17746);
and U18117 (N_18117,N_17502,N_17610);
xor U18118 (N_18118,N_17765,N_17759);
nor U18119 (N_18119,N_17977,N_17946);
nand U18120 (N_18120,N_17925,N_17974);
or U18121 (N_18121,N_17771,N_17519);
nand U18122 (N_18122,N_17782,N_17804);
and U18123 (N_18123,N_17509,N_17792);
and U18124 (N_18124,N_17796,N_17819);
or U18125 (N_18125,N_17872,N_17687);
nand U18126 (N_18126,N_17927,N_17624);
nand U18127 (N_18127,N_17736,N_17500);
or U18128 (N_18128,N_17589,N_17536);
or U18129 (N_18129,N_17696,N_17558);
nor U18130 (N_18130,N_17625,N_17887);
nand U18131 (N_18131,N_17598,N_17916);
or U18132 (N_18132,N_17875,N_17776);
nand U18133 (N_18133,N_17503,N_17588);
or U18134 (N_18134,N_17967,N_17664);
or U18135 (N_18135,N_17537,N_17701);
nand U18136 (N_18136,N_17912,N_17753);
or U18137 (N_18137,N_17926,N_17600);
or U18138 (N_18138,N_17911,N_17592);
or U18139 (N_18139,N_17531,N_17947);
or U18140 (N_18140,N_17707,N_17583);
or U18141 (N_18141,N_17793,N_17542);
nand U18142 (N_18142,N_17635,N_17724);
and U18143 (N_18143,N_17715,N_17508);
nor U18144 (N_18144,N_17941,N_17962);
or U18145 (N_18145,N_17933,N_17727);
nor U18146 (N_18146,N_17825,N_17987);
or U18147 (N_18147,N_17969,N_17614);
and U18148 (N_18148,N_17920,N_17783);
nor U18149 (N_18149,N_17645,N_17563);
and U18150 (N_18150,N_17559,N_17885);
nand U18151 (N_18151,N_17650,N_17652);
and U18152 (N_18152,N_17685,N_17640);
and U18153 (N_18153,N_17935,N_17555);
nand U18154 (N_18154,N_17880,N_17903);
nand U18155 (N_18155,N_17632,N_17859);
and U18156 (N_18156,N_17822,N_17997);
nand U18157 (N_18157,N_17717,N_17544);
and U18158 (N_18158,N_17554,N_17686);
or U18159 (N_18159,N_17860,N_17680);
and U18160 (N_18160,N_17870,N_17902);
and U18161 (N_18161,N_17520,N_17646);
xnor U18162 (N_18162,N_17857,N_17564);
nand U18163 (N_18163,N_17532,N_17808);
nand U18164 (N_18164,N_17837,N_17863);
and U18165 (N_18165,N_17944,N_17569);
and U18166 (N_18166,N_17575,N_17533);
nand U18167 (N_18167,N_17587,N_17917);
nor U18168 (N_18168,N_17633,N_17684);
xor U18169 (N_18169,N_17528,N_17865);
nor U18170 (N_18170,N_17981,N_17668);
nand U18171 (N_18171,N_17828,N_17642);
nand U18172 (N_18172,N_17914,N_17896);
or U18173 (N_18173,N_17812,N_17942);
and U18174 (N_18174,N_17690,N_17959);
xor U18175 (N_18175,N_17975,N_17976);
nor U18176 (N_18176,N_17839,N_17964);
nor U18177 (N_18177,N_17842,N_17512);
nor U18178 (N_18178,N_17599,N_17999);
nor U18179 (N_18179,N_17931,N_17856);
or U18180 (N_18180,N_17764,N_17883);
or U18181 (N_18181,N_17548,N_17924);
nand U18182 (N_18182,N_17582,N_17978);
nand U18183 (N_18183,N_17802,N_17522);
or U18184 (N_18184,N_17910,N_17689);
or U18185 (N_18185,N_17594,N_17851);
or U18186 (N_18186,N_17798,N_17619);
or U18187 (N_18187,N_17654,N_17772);
or U18188 (N_18188,N_17838,N_17636);
and U18189 (N_18189,N_17898,N_17608);
and U18190 (N_18190,N_17534,N_17989);
or U18191 (N_18191,N_17637,N_17709);
or U18192 (N_18192,N_17597,N_17529);
nor U18193 (N_18193,N_17951,N_17818);
nand U18194 (N_18194,N_17829,N_17574);
nor U18195 (N_18195,N_17877,N_17679);
and U18196 (N_18196,N_17553,N_17681);
nand U18197 (N_18197,N_17556,N_17993);
nand U18198 (N_18198,N_17674,N_17908);
nor U18199 (N_18199,N_17986,N_17601);
nand U18200 (N_18200,N_17817,N_17930);
nand U18201 (N_18201,N_17876,N_17620);
nor U18202 (N_18202,N_17756,N_17849);
and U18203 (N_18203,N_17904,N_17937);
nor U18204 (N_18204,N_17810,N_17929);
and U18205 (N_18205,N_17906,N_17873);
or U18206 (N_18206,N_17615,N_17649);
nor U18207 (N_18207,N_17538,N_17670);
or U18208 (N_18208,N_17586,N_17732);
and U18209 (N_18209,N_17616,N_17505);
nand U18210 (N_18210,N_17513,N_17936);
or U18211 (N_18211,N_17677,N_17604);
and U18212 (N_18212,N_17713,N_17938);
or U18213 (N_18213,N_17913,N_17626);
nor U18214 (N_18214,N_17506,N_17855);
nor U18215 (N_18215,N_17627,N_17546);
nor U18216 (N_18216,N_17510,N_17846);
or U18217 (N_18217,N_17749,N_17966);
and U18218 (N_18218,N_17629,N_17678);
nand U18219 (N_18219,N_17655,N_17743);
xnor U18220 (N_18220,N_17973,N_17754);
nor U18221 (N_18221,N_17507,N_17919);
or U18222 (N_18222,N_17807,N_17909);
nor U18223 (N_18223,N_17786,N_17878);
or U18224 (N_18224,N_17666,N_17730);
nor U18225 (N_18225,N_17854,N_17943);
nor U18226 (N_18226,N_17703,N_17585);
nand U18227 (N_18227,N_17868,N_17662);
nand U18228 (N_18228,N_17950,N_17801);
nand U18229 (N_18229,N_17988,N_17928);
nand U18230 (N_18230,N_17921,N_17866);
and U18231 (N_18231,N_17698,N_17830);
nand U18232 (N_18232,N_17524,N_17682);
or U18233 (N_18233,N_17644,N_17892);
nand U18234 (N_18234,N_17748,N_17939);
or U18235 (N_18235,N_17787,N_17562);
or U18236 (N_18236,N_17761,N_17853);
nor U18237 (N_18237,N_17953,N_17521);
xnor U18238 (N_18238,N_17992,N_17799);
and U18239 (N_18239,N_17835,N_17560);
nand U18240 (N_18240,N_17948,N_17656);
and U18241 (N_18241,N_17752,N_17651);
nand U18242 (N_18242,N_17814,N_17777);
or U18243 (N_18243,N_17710,N_17653);
nor U18244 (N_18244,N_17726,N_17739);
nand U18245 (N_18245,N_17738,N_17595);
nor U18246 (N_18246,N_17790,N_17705);
nor U18247 (N_18247,N_17517,N_17874);
and U18248 (N_18248,N_17747,N_17784);
or U18249 (N_18249,N_17780,N_17734);
or U18250 (N_18250,N_17756,N_17883);
and U18251 (N_18251,N_17819,N_17860);
or U18252 (N_18252,N_17921,N_17687);
or U18253 (N_18253,N_17958,N_17883);
nand U18254 (N_18254,N_17814,N_17849);
or U18255 (N_18255,N_17632,N_17808);
nand U18256 (N_18256,N_17995,N_17724);
nor U18257 (N_18257,N_17601,N_17790);
or U18258 (N_18258,N_17816,N_17505);
or U18259 (N_18259,N_17740,N_17888);
or U18260 (N_18260,N_17583,N_17599);
nor U18261 (N_18261,N_17512,N_17925);
or U18262 (N_18262,N_17926,N_17797);
or U18263 (N_18263,N_17891,N_17963);
nand U18264 (N_18264,N_17940,N_17584);
and U18265 (N_18265,N_17704,N_17682);
nor U18266 (N_18266,N_17949,N_17629);
xor U18267 (N_18267,N_17904,N_17774);
nor U18268 (N_18268,N_17965,N_17909);
or U18269 (N_18269,N_17598,N_17522);
or U18270 (N_18270,N_17669,N_17647);
or U18271 (N_18271,N_17864,N_17785);
nand U18272 (N_18272,N_17566,N_17824);
and U18273 (N_18273,N_17802,N_17855);
and U18274 (N_18274,N_17780,N_17911);
nor U18275 (N_18275,N_17695,N_17534);
nor U18276 (N_18276,N_17973,N_17961);
nand U18277 (N_18277,N_17839,N_17753);
or U18278 (N_18278,N_17606,N_17645);
and U18279 (N_18279,N_17549,N_17559);
or U18280 (N_18280,N_17987,N_17629);
and U18281 (N_18281,N_17748,N_17706);
nand U18282 (N_18282,N_17931,N_17729);
nand U18283 (N_18283,N_17576,N_17816);
and U18284 (N_18284,N_17794,N_17737);
and U18285 (N_18285,N_17946,N_17505);
nand U18286 (N_18286,N_17785,N_17729);
or U18287 (N_18287,N_17890,N_17680);
nor U18288 (N_18288,N_17656,N_17571);
and U18289 (N_18289,N_17652,N_17887);
nor U18290 (N_18290,N_17989,N_17889);
nor U18291 (N_18291,N_17988,N_17723);
nand U18292 (N_18292,N_17811,N_17939);
nand U18293 (N_18293,N_17611,N_17793);
nand U18294 (N_18294,N_17782,N_17502);
and U18295 (N_18295,N_17681,N_17930);
nand U18296 (N_18296,N_17632,N_17624);
and U18297 (N_18297,N_17788,N_17870);
nand U18298 (N_18298,N_17866,N_17677);
or U18299 (N_18299,N_17756,N_17587);
and U18300 (N_18300,N_17945,N_17913);
xnor U18301 (N_18301,N_17817,N_17905);
and U18302 (N_18302,N_17742,N_17986);
nor U18303 (N_18303,N_17555,N_17539);
and U18304 (N_18304,N_17772,N_17704);
nor U18305 (N_18305,N_17565,N_17827);
nor U18306 (N_18306,N_17905,N_17769);
or U18307 (N_18307,N_17861,N_17684);
nor U18308 (N_18308,N_17842,N_17533);
nand U18309 (N_18309,N_17902,N_17951);
or U18310 (N_18310,N_17604,N_17566);
nand U18311 (N_18311,N_17730,N_17629);
nor U18312 (N_18312,N_17695,N_17914);
nor U18313 (N_18313,N_17754,N_17910);
nand U18314 (N_18314,N_17780,N_17768);
nor U18315 (N_18315,N_17619,N_17816);
or U18316 (N_18316,N_17708,N_17730);
and U18317 (N_18317,N_17752,N_17533);
or U18318 (N_18318,N_17778,N_17559);
nor U18319 (N_18319,N_17964,N_17848);
nor U18320 (N_18320,N_17774,N_17748);
and U18321 (N_18321,N_17850,N_17984);
nor U18322 (N_18322,N_17773,N_17573);
nor U18323 (N_18323,N_17792,N_17544);
or U18324 (N_18324,N_17575,N_17674);
nand U18325 (N_18325,N_17578,N_17742);
or U18326 (N_18326,N_17618,N_17913);
or U18327 (N_18327,N_17834,N_17936);
nor U18328 (N_18328,N_17763,N_17589);
nor U18329 (N_18329,N_17527,N_17983);
or U18330 (N_18330,N_17738,N_17629);
or U18331 (N_18331,N_17591,N_17899);
nor U18332 (N_18332,N_17502,N_17565);
and U18333 (N_18333,N_17666,N_17834);
and U18334 (N_18334,N_17953,N_17576);
or U18335 (N_18335,N_17842,N_17850);
and U18336 (N_18336,N_17770,N_17548);
nand U18337 (N_18337,N_17954,N_17697);
nand U18338 (N_18338,N_17682,N_17631);
nand U18339 (N_18339,N_17881,N_17829);
nor U18340 (N_18340,N_17565,N_17869);
nor U18341 (N_18341,N_17800,N_17683);
or U18342 (N_18342,N_17529,N_17535);
nor U18343 (N_18343,N_17569,N_17629);
and U18344 (N_18344,N_17514,N_17883);
or U18345 (N_18345,N_17868,N_17859);
nand U18346 (N_18346,N_17791,N_17666);
or U18347 (N_18347,N_17980,N_17732);
nor U18348 (N_18348,N_17787,N_17829);
or U18349 (N_18349,N_17764,N_17913);
or U18350 (N_18350,N_17695,N_17727);
nor U18351 (N_18351,N_17997,N_17532);
nor U18352 (N_18352,N_17985,N_17554);
nand U18353 (N_18353,N_17959,N_17515);
nor U18354 (N_18354,N_17745,N_17673);
or U18355 (N_18355,N_17657,N_17831);
and U18356 (N_18356,N_17842,N_17540);
or U18357 (N_18357,N_17825,N_17544);
nor U18358 (N_18358,N_17648,N_17997);
or U18359 (N_18359,N_17618,N_17727);
nor U18360 (N_18360,N_17581,N_17727);
nor U18361 (N_18361,N_17670,N_17948);
nand U18362 (N_18362,N_17528,N_17665);
and U18363 (N_18363,N_17774,N_17747);
or U18364 (N_18364,N_17804,N_17718);
or U18365 (N_18365,N_17568,N_17925);
or U18366 (N_18366,N_17718,N_17657);
or U18367 (N_18367,N_17804,N_17727);
and U18368 (N_18368,N_17821,N_17877);
nand U18369 (N_18369,N_17761,N_17518);
nor U18370 (N_18370,N_17707,N_17758);
xor U18371 (N_18371,N_17602,N_17802);
and U18372 (N_18372,N_17760,N_17527);
nor U18373 (N_18373,N_17558,N_17852);
and U18374 (N_18374,N_17841,N_17858);
nand U18375 (N_18375,N_17890,N_17943);
or U18376 (N_18376,N_17729,N_17807);
and U18377 (N_18377,N_17871,N_17879);
and U18378 (N_18378,N_17603,N_17937);
or U18379 (N_18379,N_17981,N_17688);
nand U18380 (N_18380,N_17825,N_17831);
or U18381 (N_18381,N_17578,N_17735);
or U18382 (N_18382,N_17655,N_17757);
or U18383 (N_18383,N_17749,N_17922);
and U18384 (N_18384,N_17620,N_17816);
and U18385 (N_18385,N_17907,N_17744);
and U18386 (N_18386,N_17884,N_17651);
nor U18387 (N_18387,N_17847,N_17640);
and U18388 (N_18388,N_17643,N_17568);
nand U18389 (N_18389,N_17849,N_17948);
nand U18390 (N_18390,N_17561,N_17548);
and U18391 (N_18391,N_17849,N_17623);
nor U18392 (N_18392,N_17691,N_17790);
nor U18393 (N_18393,N_17911,N_17520);
or U18394 (N_18394,N_17841,N_17648);
nor U18395 (N_18395,N_17502,N_17891);
or U18396 (N_18396,N_17593,N_17791);
xnor U18397 (N_18397,N_17705,N_17549);
xor U18398 (N_18398,N_17951,N_17797);
nand U18399 (N_18399,N_17851,N_17563);
nor U18400 (N_18400,N_17621,N_17718);
and U18401 (N_18401,N_17881,N_17684);
xnor U18402 (N_18402,N_17921,N_17542);
or U18403 (N_18403,N_17819,N_17881);
nor U18404 (N_18404,N_17899,N_17857);
nand U18405 (N_18405,N_17926,N_17607);
and U18406 (N_18406,N_17918,N_17573);
nand U18407 (N_18407,N_17549,N_17913);
nor U18408 (N_18408,N_17520,N_17832);
nand U18409 (N_18409,N_17757,N_17776);
or U18410 (N_18410,N_17728,N_17857);
or U18411 (N_18411,N_17540,N_17625);
nand U18412 (N_18412,N_17513,N_17653);
and U18413 (N_18413,N_17997,N_17582);
nor U18414 (N_18414,N_17909,N_17714);
and U18415 (N_18415,N_17976,N_17629);
xor U18416 (N_18416,N_17954,N_17600);
nor U18417 (N_18417,N_17755,N_17641);
or U18418 (N_18418,N_17842,N_17928);
xnor U18419 (N_18419,N_17912,N_17599);
and U18420 (N_18420,N_17749,N_17673);
or U18421 (N_18421,N_17668,N_17813);
nor U18422 (N_18422,N_17543,N_17778);
nor U18423 (N_18423,N_17981,N_17686);
and U18424 (N_18424,N_17950,N_17688);
and U18425 (N_18425,N_17887,N_17796);
or U18426 (N_18426,N_17703,N_17707);
nor U18427 (N_18427,N_17582,N_17871);
nor U18428 (N_18428,N_17854,N_17704);
nor U18429 (N_18429,N_17869,N_17811);
nor U18430 (N_18430,N_17955,N_17721);
nor U18431 (N_18431,N_17914,N_17764);
or U18432 (N_18432,N_17542,N_17947);
and U18433 (N_18433,N_17508,N_17908);
nor U18434 (N_18434,N_17971,N_17593);
nor U18435 (N_18435,N_17592,N_17825);
nor U18436 (N_18436,N_17977,N_17853);
or U18437 (N_18437,N_17509,N_17930);
and U18438 (N_18438,N_17820,N_17510);
and U18439 (N_18439,N_17535,N_17599);
nor U18440 (N_18440,N_17973,N_17676);
nand U18441 (N_18441,N_17717,N_17666);
or U18442 (N_18442,N_17768,N_17965);
nor U18443 (N_18443,N_17599,N_17978);
nand U18444 (N_18444,N_17662,N_17945);
nor U18445 (N_18445,N_17832,N_17556);
nand U18446 (N_18446,N_17904,N_17649);
and U18447 (N_18447,N_17784,N_17652);
or U18448 (N_18448,N_17576,N_17657);
nand U18449 (N_18449,N_17883,N_17704);
nand U18450 (N_18450,N_17719,N_17543);
or U18451 (N_18451,N_17981,N_17750);
nand U18452 (N_18452,N_17619,N_17823);
nor U18453 (N_18453,N_17898,N_17654);
nor U18454 (N_18454,N_17931,N_17559);
and U18455 (N_18455,N_17970,N_17526);
and U18456 (N_18456,N_17841,N_17865);
nand U18457 (N_18457,N_17815,N_17892);
and U18458 (N_18458,N_17908,N_17554);
nor U18459 (N_18459,N_17548,N_17672);
nor U18460 (N_18460,N_17634,N_17923);
nor U18461 (N_18461,N_17850,N_17754);
or U18462 (N_18462,N_17535,N_17826);
nor U18463 (N_18463,N_17943,N_17785);
nand U18464 (N_18464,N_17928,N_17674);
nand U18465 (N_18465,N_17571,N_17825);
nor U18466 (N_18466,N_17746,N_17704);
nand U18467 (N_18467,N_17512,N_17770);
and U18468 (N_18468,N_17671,N_17949);
nor U18469 (N_18469,N_17543,N_17964);
nand U18470 (N_18470,N_17566,N_17964);
or U18471 (N_18471,N_17646,N_17874);
nor U18472 (N_18472,N_17663,N_17518);
or U18473 (N_18473,N_17727,N_17522);
and U18474 (N_18474,N_17660,N_17889);
and U18475 (N_18475,N_17685,N_17555);
nor U18476 (N_18476,N_17640,N_17713);
nand U18477 (N_18477,N_17860,N_17900);
nor U18478 (N_18478,N_17802,N_17632);
nand U18479 (N_18479,N_17644,N_17674);
and U18480 (N_18480,N_17807,N_17919);
and U18481 (N_18481,N_17999,N_17909);
nor U18482 (N_18482,N_17651,N_17594);
nand U18483 (N_18483,N_17549,N_17534);
nor U18484 (N_18484,N_17771,N_17633);
nand U18485 (N_18485,N_17907,N_17652);
and U18486 (N_18486,N_17658,N_17745);
or U18487 (N_18487,N_17706,N_17637);
or U18488 (N_18488,N_17625,N_17870);
nand U18489 (N_18489,N_17607,N_17869);
or U18490 (N_18490,N_17994,N_17847);
or U18491 (N_18491,N_17803,N_17990);
or U18492 (N_18492,N_17789,N_17907);
nand U18493 (N_18493,N_17824,N_17946);
nor U18494 (N_18494,N_17864,N_17882);
nor U18495 (N_18495,N_17790,N_17753);
or U18496 (N_18496,N_17745,N_17773);
and U18497 (N_18497,N_17897,N_17738);
nor U18498 (N_18498,N_17722,N_17908);
nor U18499 (N_18499,N_17553,N_17602);
or U18500 (N_18500,N_18403,N_18078);
nand U18501 (N_18501,N_18192,N_18439);
or U18502 (N_18502,N_18483,N_18111);
nand U18503 (N_18503,N_18297,N_18344);
and U18504 (N_18504,N_18097,N_18148);
nor U18505 (N_18505,N_18212,N_18052);
or U18506 (N_18506,N_18017,N_18405);
nor U18507 (N_18507,N_18061,N_18179);
or U18508 (N_18508,N_18203,N_18376);
and U18509 (N_18509,N_18289,N_18308);
nor U18510 (N_18510,N_18493,N_18230);
or U18511 (N_18511,N_18459,N_18228);
nand U18512 (N_18512,N_18118,N_18051);
and U18513 (N_18513,N_18112,N_18434);
nand U18514 (N_18514,N_18484,N_18214);
nor U18515 (N_18515,N_18425,N_18158);
nor U18516 (N_18516,N_18235,N_18055);
and U18517 (N_18517,N_18360,N_18461);
or U18518 (N_18518,N_18002,N_18342);
or U18519 (N_18519,N_18033,N_18057);
and U18520 (N_18520,N_18077,N_18162);
or U18521 (N_18521,N_18433,N_18045);
nor U18522 (N_18522,N_18027,N_18475);
nand U18523 (N_18523,N_18207,N_18106);
and U18524 (N_18524,N_18307,N_18411);
and U18525 (N_18525,N_18378,N_18181);
or U18526 (N_18526,N_18080,N_18471);
or U18527 (N_18527,N_18088,N_18169);
and U18528 (N_18528,N_18153,N_18117);
and U18529 (N_18529,N_18102,N_18218);
and U18530 (N_18530,N_18401,N_18276);
or U18531 (N_18531,N_18019,N_18053);
nand U18532 (N_18532,N_18274,N_18455);
nor U18533 (N_18533,N_18272,N_18479);
nor U18534 (N_18534,N_18193,N_18238);
or U18535 (N_18535,N_18372,N_18236);
nand U18536 (N_18536,N_18406,N_18195);
and U18537 (N_18537,N_18101,N_18384);
and U18538 (N_18538,N_18056,N_18300);
nand U18539 (N_18539,N_18453,N_18032);
or U18540 (N_18540,N_18438,N_18029);
nand U18541 (N_18541,N_18028,N_18164);
nand U18542 (N_18542,N_18211,N_18256);
nand U18543 (N_18543,N_18059,N_18143);
nand U18544 (N_18544,N_18227,N_18172);
nand U18545 (N_18545,N_18322,N_18496);
or U18546 (N_18546,N_18280,N_18432);
and U18547 (N_18547,N_18240,N_18122);
nor U18548 (N_18548,N_18410,N_18288);
and U18549 (N_18549,N_18377,N_18124);
nand U18550 (N_18550,N_18219,N_18366);
nand U18551 (N_18551,N_18152,N_18160);
or U18552 (N_18552,N_18146,N_18065);
nor U18553 (N_18553,N_18182,N_18351);
and U18554 (N_18554,N_18263,N_18008);
nor U18555 (N_18555,N_18333,N_18290);
and U18556 (N_18556,N_18417,N_18202);
nand U18557 (N_18557,N_18244,N_18408);
nand U18558 (N_18558,N_18311,N_18265);
nand U18559 (N_18559,N_18488,N_18458);
nor U18560 (N_18560,N_18451,N_18119);
or U18561 (N_18561,N_18326,N_18315);
nand U18562 (N_18562,N_18035,N_18069);
nand U18563 (N_18563,N_18220,N_18171);
or U18564 (N_18564,N_18175,N_18463);
nand U18565 (N_18565,N_18382,N_18229);
or U18566 (N_18566,N_18457,N_18015);
nand U18567 (N_18567,N_18054,N_18134);
nor U18568 (N_18568,N_18076,N_18489);
or U18569 (N_18569,N_18103,N_18180);
nor U18570 (N_18570,N_18440,N_18269);
nand U18571 (N_18571,N_18109,N_18167);
nor U18572 (N_18572,N_18003,N_18215);
or U18573 (N_18573,N_18359,N_18329);
nor U18574 (N_18574,N_18092,N_18413);
or U18575 (N_18575,N_18089,N_18096);
nand U18576 (N_18576,N_18173,N_18304);
nor U18577 (N_18577,N_18205,N_18424);
nor U18578 (N_18578,N_18323,N_18198);
or U18579 (N_18579,N_18436,N_18446);
nor U18580 (N_18580,N_18114,N_18213);
or U18581 (N_18581,N_18460,N_18468);
nor U18582 (N_18582,N_18137,N_18121);
nor U18583 (N_18583,N_18155,N_18268);
nor U18584 (N_18584,N_18098,N_18048);
nand U18585 (N_18585,N_18068,N_18264);
nand U18586 (N_18586,N_18324,N_18467);
nor U18587 (N_18587,N_18397,N_18337);
nor U18588 (N_18588,N_18177,N_18282);
or U18589 (N_18589,N_18334,N_18250);
nor U18590 (N_18590,N_18448,N_18099);
and U18591 (N_18591,N_18064,N_18402);
nand U18592 (N_18592,N_18415,N_18414);
and U18593 (N_18593,N_18473,N_18041);
nand U18594 (N_18594,N_18348,N_18336);
or U18595 (N_18595,N_18389,N_18184);
nor U18596 (N_18596,N_18497,N_18233);
or U18597 (N_18597,N_18349,N_18197);
and U18598 (N_18598,N_18150,N_18259);
nand U18599 (N_18599,N_18430,N_18340);
nor U18600 (N_18600,N_18367,N_18454);
or U18601 (N_18601,N_18159,N_18199);
and U18602 (N_18602,N_18094,N_18310);
and U18603 (N_18603,N_18060,N_18083);
or U18604 (N_18604,N_18049,N_18363);
or U18605 (N_18605,N_18115,N_18379);
or U18606 (N_18606,N_18431,N_18185);
and U18607 (N_18607,N_18075,N_18187);
nor U18608 (N_18608,N_18319,N_18277);
nand U18609 (N_18609,N_18317,N_18086);
nor U18610 (N_18610,N_18222,N_18281);
or U18611 (N_18611,N_18084,N_18437);
or U18612 (N_18612,N_18296,N_18302);
nand U18613 (N_18613,N_18252,N_18001);
xor U18614 (N_18614,N_18347,N_18245);
nor U18615 (N_18615,N_18293,N_18320);
nor U18616 (N_18616,N_18313,N_18482);
or U18617 (N_18617,N_18399,N_18144);
xnor U18618 (N_18618,N_18472,N_18125);
nand U18619 (N_18619,N_18224,N_18487);
nand U18620 (N_18620,N_18262,N_18418);
nor U18621 (N_18621,N_18133,N_18168);
and U18622 (N_18622,N_18420,N_18298);
or U18623 (N_18623,N_18025,N_18407);
nor U18624 (N_18624,N_18231,N_18387);
nand U18625 (N_18625,N_18492,N_18191);
or U18626 (N_18626,N_18295,N_18139);
xnor U18627 (N_18627,N_18412,N_18216);
nor U18628 (N_18628,N_18355,N_18243);
xnor U18629 (N_18629,N_18452,N_18450);
or U18630 (N_18630,N_18044,N_18005);
and U18631 (N_18631,N_18163,N_18404);
and U18632 (N_18632,N_18299,N_18200);
or U18633 (N_18633,N_18237,N_18138);
nor U18634 (N_18634,N_18428,N_18157);
nand U18635 (N_18635,N_18232,N_18328);
nor U18636 (N_18636,N_18369,N_18020);
and U18637 (N_18637,N_18022,N_18023);
or U18638 (N_18638,N_18085,N_18046);
or U18639 (N_18639,N_18273,N_18477);
nand U18640 (N_18640,N_18251,N_18206);
nand U18641 (N_18641,N_18338,N_18013);
or U18642 (N_18642,N_18120,N_18267);
nand U18643 (N_18643,N_18325,N_18021);
or U18644 (N_18644,N_18006,N_18257);
xor U18645 (N_18645,N_18043,N_18226);
nor U18646 (N_18646,N_18186,N_18246);
nand U18647 (N_18647,N_18255,N_18287);
nand U18648 (N_18648,N_18066,N_18396);
nor U18649 (N_18649,N_18201,N_18283);
nor U18650 (N_18650,N_18464,N_18070);
or U18651 (N_18651,N_18062,N_18135);
nand U18652 (N_18652,N_18480,N_18161);
and U18653 (N_18653,N_18291,N_18422);
and U18654 (N_18654,N_18266,N_18409);
or U18655 (N_18655,N_18435,N_18470);
and U18656 (N_18656,N_18395,N_18104);
or U18657 (N_18657,N_18332,N_18067);
nand U18658 (N_18658,N_18365,N_18034);
nor U18659 (N_18659,N_18241,N_18016);
nand U18660 (N_18660,N_18474,N_18393);
nor U18661 (N_18661,N_18183,N_18261);
and U18662 (N_18662,N_18305,N_18292);
or U18663 (N_18663,N_18270,N_18113);
and U18664 (N_18664,N_18427,N_18485);
nor U18665 (N_18665,N_18466,N_18381);
or U18666 (N_18666,N_18426,N_18204);
nand U18667 (N_18667,N_18275,N_18284);
nor U18668 (N_18668,N_18358,N_18303);
or U18669 (N_18669,N_18314,N_18419);
nand U18670 (N_18670,N_18140,N_18478);
or U18671 (N_18671,N_18242,N_18239);
nor U18672 (N_18672,N_18354,N_18371);
or U18673 (N_18673,N_18343,N_18040);
and U18674 (N_18674,N_18095,N_18058);
and U18675 (N_18675,N_18105,N_18294);
and U18676 (N_18676,N_18330,N_18312);
and U18677 (N_18677,N_18038,N_18494);
nand U18678 (N_18678,N_18030,N_18126);
and U18679 (N_18679,N_18429,N_18189);
nand U18680 (N_18680,N_18416,N_18026);
or U18681 (N_18681,N_18443,N_18499);
or U18682 (N_18682,N_18301,N_18039);
nor U18683 (N_18683,N_18345,N_18012);
and U18684 (N_18684,N_18190,N_18390);
and U18685 (N_18685,N_18386,N_18210);
and U18686 (N_18686,N_18007,N_18170);
or U18687 (N_18687,N_18271,N_18093);
nor U18688 (N_18688,N_18388,N_18421);
nor U18689 (N_18689,N_18154,N_18130);
or U18690 (N_18690,N_18074,N_18339);
nor U18691 (N_18691,N_18364,N_18221);
nand U18692 (N_18692,N_18374,N_18335);
nand U18693 (N_18693,N_18249,N_18254);
nor U18694 (N_18694,N_18036,N_18341);
and U18695 (N_18695,N_18108,N_18368);
nand U18696 (N_18696,N_18151,N_18072);
or U18697 (N_18697,N_18316,N_18456);
or U18698 (N_18698,N_18286,N_18385);
and U18699 (N_18699,N_18447,N_18209);
nand U18700 (N_18700,N_18361,N_18441);
and U18701 (N_18701,N_18350,N_18423);
or U18702 (N_18702,N_18081,N_18346);
or U18703 (N_18703,N_18178,N_18018);
or U18704 (N_18704,N_18306,N_18498);
or U18705 (N_18705,N_18285,N_18208);
or U18706 (N_18706,N_18165,N_18260);
nand U18707 (N_18707,N_18063,N_18004);
and U18708 (N_18708,N_18073,N_18370);
or U18709 (N_18709,N_18279,N_18142);
nor U18710 (N_18710,N_18194,N_18100);
nand U18711 (N_18711,N_18469,N_18149);
xnor U18712 (N_18712,N_18253,N_18462);
and U18713 (N_18713,N_18107,N_18331);
or U18714 (N_18714,N_18116,N_18373);
nand U18715 (N_18715,N_18491,N_18449);
and U18716 (N_18716,N_18357,N_18147);
nor U18717 (N_18717,N_18188,N_18014);
nor U18718 (N_18718,N_18136,N_18010);
and U18719 (N_18719,N_18129,N_18156);
and U18720 (N_18720,N_18166,N_18087);
nor U18721 (N_18721,N_18380,N_18248);
or U18722 (N_18722,N_18176,N_18217);
nand U18723 (N_18723,N_18037,N_18353);
nor U18724 (N_18724,N_18465,N_18490);
nor U18725 (N_18725,N_18011,N_18000);
nor U18726 (N_18726,N_18225,N_18352);
and U18727 (N_18727,N_18445,N_18082);
nand U18728 (N_18728,N_18174,N_18127);
nor U18729 (N_18729,N_18481,N_18327);
and U18730 (N_18730,N_18258,N_18318);
nand U18731 (N_18731,N_18132,N_18486);
or U18732 (N_18732,N_18383,N_18356);
nand U18733 (N_18733,N_18495,N_18247);
or U18734 (N_18734,N_18050,N_18400);
nand U18735 (N_18735,N_18398,N_18223);
or U18736 (N_18736,N_18476,N_18375);
or U18737 (N_18737,N_18009,N_18128);
xnor U18738 (N_18738,N_18196,N_18047);
nor U18739 (N_18739,N_18234,N_18278);
nor U18740 (N_18740,N_18442,N_18110);
and U18741 (N_18741,N_18091,N_18444);
nand U18742 (N_18742,N_18024,N_18321);
and U18743 (N_18743,N_18391,N_18392);
or U18744 (N_18744,N_18309,N_18131);
and U18745 (N_18745,N_18394,N_18090);
or U18746 (N_18746,N_18042,N_18362);
nand U18747 (N_18747,N_18031,N_18079);
nand U18748 (N_18748,N_18145,N_18123);
or U18749 (N_18749,N_18071,N_18141);
nor U18750 (N_18750,N_18136,N_18083);
nand U18751 (N_18751,N_18199,N_18137);
and U18752 (N_18752,N_18093,N_18372);
or U18753 (N_18753,N_18116,N_18248);
and U18754 (N_18754,N_18126,N_18011);
and U18755 (N_18755,N_18215,N_18441);
and U18756 (N_18756,N_18155,N_18180);
and U18757 (N_18757,N_18198,N_18250);
nor U18758 (N_18758,N_18263,N_18103);
nand U18759 (N_18759,N_18137,N_18187);
xor U18760 (N_18760,N_18220,N_18269);
nand U18761 (N_18761,N_18043,N_18379);
xnor U18762 (N_18762,N_18192,N_18150);
nor U18763 (N_18763,N_18189,N_18276);
or U18764 (N_18764,N_18285,N_18029);
nand U18765 (N_18765,N_18285,N_18202);
nor U18766 (N_18766,N_18235,N_18182);
nand U18767 (N_18767,N_18355,N_18442);
nand U18768 (N_18768,N_18476,N_18139);
nor U18769 (N_18769,N_18104,N_18297);
and U18770 (N_18770,N_18316,N_18247);
and U18771 (N_18771,N_18216,N_18491);
nand U18772 (N_18772,N_18319,N_18459);
or U18773 (N_18773,N_18310,N_18320);
and U18774 (N_18774,N_18312,N_18245);
or U18775 (N_18775,N_18039,N_18292);
nand U18776 (N_18776,N_18302,N_18408);
nand U18777 (N_18777,N_18204,N_18414);
nand U18778 (N_18778,N_18304,N_18371);
or U18779 (N_18779,N_18358,N_18483);
nand U18780 (N_18780,N_18091,N_18328);
and U18781 (N_18781,N_18083,N_18113);
or U18782 (N_18782,N_18189,N_18281);
or U18783 (N_18783,N_18007,N_18332);
and U18784 (N_18784,N_18220,N_18287);
nor U18785 (N_18785,N_18263,N_18117);
and U18786 (N_18786,N_18025,N_18058);
and U18787 (N_18787,N_18069,N_18244);
nor U18788 (N_18788,N_18397,N_18145);
nor U18789 (N_18789,N_18434,N_18012);
nand U18790 (N_18790,N_18078,N_18244);
nor U18791 (N_18791,N_18195,N_18418);
nor U18792 (N_18792,N_18052,N_18149);
or U18793 (N_18793,N_18476,N_18173);
and U18794 (N_18794,N_18394,N_18226);
or U18795 (N_18795,N_18097,N_18395);
nand U18796 (N_18796,N_18082,N_18213);
nor U18797 (N_18797,N_18262,N_18455);
and U18798 (N_18798,N_18261,N_18202);
nand U18799 (N_18799,N_18048,N_18187);
or U18800 (N_18800,N_18363,N_18048);
and U18801 (N_18801,N_18339,N_18118);
or U18802 (N_18802,N_18002,N_18253);
and U18803 (N_18803,N_18406,N_18014);
nor U18804 (N_18804,N_18498,N_18263);
nand U18805 (N_18805,N_18141,N_18155);
nand U18806 (N_18806,N_18254,N_18253);
or U18807 (N_18807,N_18104,N_18009);
and U18808 (N_18808,N_18378,N_18306);
or U18809 (N_18809,N_18340,N_18134);
nor U18810 (N_18810,N_18324,N_18255);
and U18811 (N_18811,N_18132,N_18367);
nand U18812 (N_18812,N_18165,N_18155);
or U18813 (N_18813,N_18453,N_18472);
nor U18814 (N_18814,N_18182,N_18247);
nand U18815 (N_18815,N_18297,N_18402);
nand U18816 (N_18816,N_18471,N_18065);
nand U18817 (N_18817,N_18388,N_18069);
or U18818 (N_18818,N_18013,N_18351);
and U18819 (N_18819,N_18395,N_18166);
xnor U18820 (N_18820,N_18487,N_18061);
and U18821 (N_18821,N_18369,N_18249);
nor U18822 (N_18822,N_18294,N_18239);
or U18823 (N_18823,N_18442,N_18311);
nand U18824 (N_18824,N_18057,N_18291);
or U18825 (N_18825,N_18398,N_18178);
or U18826 (N_18826,N_18273,N_18077);
and U18827 (N_18827,N_18347,N_18420);
nand U18828 (N_18828,N_18201,N_18351);
nor U18829 (N_18829,N_18317,N_18024);
or U18830 (N_18830,N_18289,N_18371);
and U18831 (N_18831,N_18128,N_18358);
and U18832 (N_18832,N_18060,N_18295);
nand U18833 (N_18833,N_18248,N_18013);
and U18834 (N_18834,N_18167,N_18383);
and U18835 (N_18835,N_18490,N_18194);
nor U18836 (N_18836,N_18433,N_18405);
and U18837 (N_18837,N_18213,N_18287);
nor U18838 (N_18838,N_18492,N_18422);
nor U18839 (N_18839,N_18293,N_18311);
nand U18840 (N_18840,N_18279,N_18477);
nand U18841 (N_18841,N_18152,N_18213);
nand U18842 (N_18842,N_18464,N_18452);
and U18843 (N_18843,N_18094,N_18374);
and U18844 (N_18844,N_18450,N_18214);
nor U18845 (N_18845,N_18085,N_18097);
nand U18846 (N_18846,N_18160,N_18433);
and U18847 (N_18847,N_18200,N_18238);
nand U18848 (N_18848,N_18294,N_18055);
or U18849 (N_18849,N_18385,N_18229);
nand U18850 (N_18850,N_18418,N_18347);
or U18851 (N_18851,N_18074,N_18286);
or U18852 (N_18852,N_18190,N_18141);
nand U18853 (N_18853,N_18277,N_18121);
or U18854 (N_18854,N_18133,N_18493);
or U18855 (N_18855,N_18394,N_18066);
and U18856 (N_18856,N_18244,N_18195);
and U18857 (N_18857,N_18186,N_18408);
or U18858 (N_18858,N_18049,N_18424);
and U18859 (N_18859,N_18315,N_18114);
or U18860 (N_18860,N_18494,N_18187);
or U18861 (N_18861,N_18362,N_18240);
and U18862 (N_18862,N_18383,N_18128);
nor U18863 (N_18863,N_18355,N_18118);
or U18864 (N_18864,N_18066,N_18228);
or U18865 (N_18865,N_18249,N_18319);
nand U18866 (N_18866,N_18178,N_18122);
or U18867 (N_18867,N_18318,N_18094);
xor U18868 (N_18868,N_18022,N_18070);
or U18869 (N_18869,N_18199,N_18399);
nor U18870 (N_18870,N_18131,N_18225);
nand U18871 (N_18871,N_18310,N_18156);
nand U18872 (N_18872,N_18126,N_18294);
nor U18873 (N_18873,N_18013,N_18072);
nor U18874 (N_18874,N_18347,N_18110);
nor U18875 (N_18875,N_18355,N_18202);
nor U18876 (N_18876,N_18311,N_18135);
nor U18877 (N_18877,N_18410,N_18253);
or U18878 (N_18878,N_18158,N_18006);
xor U18879 (N_18879,N_18163,N_18006);
nor U18880 (N_18880,N_18375,N_18232);
nor U18881 (N_18881,N_18227,N_18385);
or U18882 (N_18882,N_18372,N_18060);
or U18883 (N_18883,N_18455,N_18167);
nand U18884 (N_18884,N_18008,N_18368);
and U18885 (N_18885,N_18002,N_18029);
nor U18886 (N_18886,N_18464,N_18146);
xor U18887 (N_18887,N_18141,N_18024);
nor U18888 (N_18888,N_18316,N_18335);
nor U18889 (N_18889,N_18315,N_18008);
nor U18890 (N_18890,N_18240,N_18222);
or U18891 (N_18891,N_18307,N_18189);
or U18892 (N_18892,N_18005,N_18381);
nand U18893 (N_18893,N_18301,N_18241);
nand U18894 (N_18894,N_18362,N_18345);
nor U18895 (N_18895,N_18266,N_18385);
and U18896 (N_18896,N_18421,N_18228);
or U18897 (N_18897,N_18463,N_18342);
or U18898 (N_18898,N_18280,N_18313);
or U18899 (N_18899,N_18429,N_18200);
or U18900 (N_18900,N_18491,N_18052);
or U18901 (N_18901,N_18486,N_18125);
nor U18902 (N_18902,N_18204,N_18119);
and U18903 (N_18903,N_18305,N_18153);
nand U18904 (N_18904,N_18456,N_18326);
nor U18905 (N_18905,N_18259,N_18386);
xnor U18906 (N_18906,N_18122,N_18392);
or U18907 (N_18907,N_18185,N_18234);
or U18908 (N_18908,N_18210,N_18428);
and U18909 (N_18909,N_18214,N_18094);
nor U18910 (N_18910,N_18285,N_18324);
nand U18911 (N_18911,N_18250,N_18497);
or U18912 (N_18912,N_18169,N_18403);
nand U18913 (N_18913,N_18012,N_18068);
nand U18914 (N_18914,N_18372,N_18226);
and U18915 (N_18915,N_18476,N_18155);
and U18916 (N_18916,N_18417,N_18251);
nor U18917 (N_18917,N_18411,N_18089);
and U18918 (N_18918,N_18154,N_18236);
nand U18919 (N_18919,N_18090,N_18476);
or U18920 (N_18920,N_18440,N_18057);
nand U18921 (N_18921,N_18441,N_18390);
nor U18922 (N_18922,N_18143,N_18490);
nor U18923 (N_18923,N_18399,N_18204);
nor U18924 (N_18924,N_18105,N_18242);
nand U18925 (N_18925,N_18396,N_18271);
nand U18926 (N_18926,N_18420,N_18243);
nor U18927 (N_18927,N_18030,N_18118);
nand U18928 (N_18928,N_18149,N_18318);
nand U18929 (N_18929,N_18201,N_18006);
and U18930 (N_18930,N_18410,N_18031);
nor U18931 (N_18931,N_18095,N_18112);
or U18932 (N_18932,N_18075,N_18462);
nand U18933 (N_18933,N_18165,N_18133);
nand U18934 (N_18934,N_18162,N_18457);
nand U18935 (N_18935,N_18277,N_18148);
nand U18936 (N_18936,N_18138,N_18408);
and U18937 (N_18937,N_18310,N_18369);
or U18938 (N_18938,N_18349,N_18025);
nor U18939 (N_18939,N_18057,N_18163);
nor U18940 (N_18940,N_18139,N_18369);
nand U18941 (N_18941,N_18485,N_18299);
nor U18942 (N_18942,N_18074,N_18448);
or U18943 (N_18943,N_18374,N_18245);
and U18944 (N_18944,N_18106,N_18047);
nor U18945 (N_18945,N_18310,N_18232);
or U18946 (N_18946,N_18021,N_18320);
and U18947 (N_18947,N_18391,N_18179);
and U18948 (N_18948,N_18112,N_18367);
nand U18949 (N_18949,N_18304,N_18151);
nor U18950 (N_18950,N_18310,N_18143);
and U18951 (N_18951,N_18375,N_18217);
nand U18952 (N_18952,N_18303,N_18109);
and U18953 (N_18953,N_18419,N_18387);
nand U18954 (N_18954,N_18172,N_18020);
nor U18955 (N_18955,N_18078,N_18209);
nor U18956 (N_18956,N_18480,N_18383);
or U18957 (N_18957,N_18096,N_18040);
and U18958 (N_18958,N_18067,N_18372);
and U18959 (N_18959,N_18375,N_18428);
nand U18960 (N_18960,N_18165,N_18427);
nand U18961 (N_18961,N_18498,N_18406);
nand U18962 (N_18962,N_18050,N_18000);
nand U18963 (N_18963,N_18354,N_18321);
or U18964 (N_18964,N_18444,N_18121);
nor U18965 (N_18965,N_18247,N_18075);
nor U18966 (N_18966,N_18097,N_18042);
or U18967 (N_18967,N_18411,N_18257);
or U18968 (N_18968,N_18428,N_18295);
or U18969 (N_18969,N_18412,N_18142);
and U18970 (N_18970,N_18045,N_18342);
and U18971 (N_18971,N_18423,N_18203);
nand U18972 (N_18972,N_18444,N_18083);
nor U18973 (N_18973,N_18433,N_18165);
or U18974 (N_18974,N_18208,N_18089);
nor U18975 (N_18975,N_18181,N_18044);
and U18976 (N_18976,N_18401,N_18268);
and U18977 (N_18977,N_18010,N_18131);
or U18978 (N_18978,N_18013,N_18326);
nand U18979 (N_18979,N_18450,N_18402);
or U18980 (N_18980,N_18486,N_18324);
and U18981 (N_18981,N_18085,N_18399);
nand U18982 (N_18982,N_18150,N_18268);
and U18983 (N_18983,N_18243,N_18421);
and U18984 (N_18984,N_18458,N_18391);
nand U18985 (N_18985,N_18201,N_18147);
nor U18986 (N_18986,N_18060,N_18492);
nor U18987 (N_18987,N_18080,N_18142);
nand U18988 (N_18988,N_18159,N_18216);
nand U18989 (N_18989,N_18345,N_18455);
or U18990 (N_18990,N_18054,N_18196);
or U18991 (N_18991,N_18273,N_18333);
nor U18992 (N_18992,N_18312,N_18453);
nor U18993 (N_18993,N_18116,N_18345);
and U18994 (N_18994,N_18439,N_18197);
or U18995 (N_18995,N_18274,N_18214);
nand U18996 (N_18996,N_18393,N_18295);
and U18997 (N_18997,N_18383,N_18035);
nand U18998 (N_18998,N_18191,N_18142);
and U18999 (N_18999,N_18275,N_18041);
and U19000 (N_19000,N_18759,N_18722);
nand U19001 (N_19001,N_18553,N_18867);
or U19002 (N_19002,N_18510,N_18764);
or U19003 (N_19003,N_18707,N_18820);
and U19004 (N_19004,N_18763,N_18717);
xnor U19005 (N_19005,N_18650,N_18811);
or U19006 (N_19006,N_18581,N_18950);
nand U19007 (N_19007,N_18635,N_18515);
nor U19008 (N_19008,N_18833,N_18830);
and U19009 (N_19009,N_18855,N_18692);
nor U19010 (N_19010,N_18708,N_18980);
and U19011 (N_19011,N_18557,N_18985);
or U19012 (N_19012,N_18518,N_18712);
nor U19013 (N_19013,N_18746,N_18947);
nand U19014 (N_19014,N_18787,N_18979);
or U19015 (N_19015,N_18585,N_18901);
or U19016 (N_19016,N_18528,N_18680);
and U19017 (N_19017,N_18736,N_18517);
xnor U19018 (N_19018,N_18807,N_18597);
and U19019 (N_19019,N_18819,N_18639);
nand U19020 (N_19020,N_18959,N_18823);
and U19021 (N_19021,N_18628,N_18644);
or U19022 (N_19022,N_18610,N_18744);
nor U19023 (N_19023,N_18724,N_18589);
nand U19024 (N_19024,N_18785,N_18932);
and U19025 (N_19025,N_18713,N_18630);
and U19026 (N_19026,N_18852,N_18730);
and U19027 (N_19027,N_18931,N_18691);
and U19028 (N_19028,N_18989,N_18544);
nand U19029 (N_19029,N_18714,N_18667);
and U19030 (N_19030,N_18929,N_18854);
nor U19031 (N_19031,N_18601,N_18758);
nor U19032 (N_19032,N_18834,N_18564);
or U19033 (N_19033,N_18777,N_18728);
nand U19034 (N_19034,N_18827,N_18599);
nor U19035 (N_19035,N_18533,N_18647);
nor U19036 (N_19036,N_18657,N_18732);
or U19037 (N_19037,N_18700,N_18580);
nand U19038 (N_19038,N_18757,N_18706);
or U19039 (N_19039,N_18592,N_18671);
or U19040 (N_19040,N_18864,N_18975);
nor U19041 (N_19041,N_18921,N_18578);
nor U19042 (N_19042,N_18902,N_18905);
nor U19043 (N_19043,N_18966,N_18727);
and U19044 (N_19044,N_18733,N_18535);
nand U19045 (N_19045,N_18917,N_18649);
nand U19046 (N_19046,N_18782,N_18681);
and U19047 (N_19047,N_18600,N_18705);
nor U19048 (N_19048,N_18507,N_18716);
and U19049 (N_19049,N_18735,N_18840);
nor U19050 (N_19050,N_18752,N_18817);
nand U19051 (N_19051,N_18844,N_18933);
and U19052 (N_19052,N_18542,N_18572);
and U19053 (N_19053,N_18586,N_18641);
and U19054 (N_19054,N_18690,N_18894);
and U19055 (N_19055,N_18748,N_18622);
nor U19056 (N_19056,N_18543,N_18783);
and U19057 (N_19057,N_18660,N_18842);
or U19058 (N_19058,N_18829,N_18656);
or U19059 (N_19059,N_18996,N_18743);
nor U19060 (N_19060,N_18973,N_18835);
or U19061 (N_19061,N_18918,N_18673);
nor U19062 (N_19062,N_18879,N_18942);
and U19063 (N_19063,N_18627,N_18825);
nor U19064 (N_19064,N_18792,N_18814);
and U19065 (N_19065,N_18606,N_18974);
nor U19066 (N_19066,N_18780,N_18756);
nor U19067 (N_19067,N_18922,N_18960);
nand U19068 (N_19068,N_18520,N_18948);
or U19069 (N_19069,N_18614,N_18672);
nor U19070 (N_19070,N_18923,N_18915);
or U19071 (N_19071,N_18541,N_18761);
nand U19072 (N_19072,N_18514,N_18984);
nand U19073 (N_19073,N_18935,N_18749);
nor U19074 (N_19074,N_18721,N_18981);
nor U19075 (N_19075,N_18697,N_18593);
nor U19076 (N_19076,N_18781,N_18993);
nor U19077 (N_19077,N_18790,N_18512);
nand U19078 (N_19078,N_18893,N_18669);
or U19079 (N_19079,N_18804,N_18890);
nor U19080 (N_19080,N_18715,N_18693);
nor U19081 (N_19081,N_18686,N_18869);
nor U19082 (N_19082,N_18654,N_18881);
nand U19083 (N_19083,N_18674,N_18958);
or U19084 (N_19084,N_18696,N_18702);
nand U19085 (N_19085,N_18624,N_18768);
and U19086 (N_19086,N_18760,N_18910);
nor U19087 (N_19087,N_18565,N_18784);
and U19088 (N_19088,N_18615,N_18653);
and U19089 (N_19089,N_18848,N_18509);
nor U19090 (N_19090,N_18908,N_18766);
nand U19091 (N_19091,N_18527,N_18583);
nor U19092 (N_19092,N_18786,N_18555);
nor U19093 (N_19093,N_18577,N_18837);
nor U19094 (N_19094,N_18949,N_18658);
nor U19095 (N_19095,N_18661,N_18888);
nor U19096 (N_19096,N_18626,N_18505);
and U19097 (N_19097,N_18591,N_18916);
or U19098 (N_19098,N_18547,N_18988);
nor U19099 (N_19099,N_18548,N_18619);
and U19100 (N_19100,N_18634,N_18638);
nor U19101 (N_19101,N_18519,N_18725);
and U19102 (N_19102,N_18664,N_18957);
nand U19103 (N_19103,N_18865,N_18576);
or U19104 (N_19104,N_18720,N_18675);
nor U19105 (N_19105,N_18907,N_18618);
nor U19106 (N_19106,N_18554,N_18579);
or U19107 (N_19107,N_18801,N_18524);
or U19108 (N_19108,N_18972,N_18739);
and U19109 (N_19109,N_18711,N_18677);
or U19110 (N_19110,N_18682,N_18569);
or U19111 (N_19111,N_18596,N_18952);
nand U19112 (N_19112,N_18631,N_18602);
and U19113 (N_19113,N_18584,N_18611);
and U19114 (N_19114,N_18847,N_18587);
or U19115 (N_19115,N_18856,N_18872);
and U19116 (N_19116,N_18816,N_18843);
and U19117 (N_19117,N_18729,N_18574);
and U19118 (N_19118,N_18617,N_18964);
nand U19119 (N_19119,N_18769,N_18886);
nand U19120 (N_19120,N_18805,N_18689);
and U19121 (N_19121,N_18871,N_18963);
nand U19122 (N_19122,N_18516,N_18562);
nand U19123 (N_19123,N_18740,N_18956);
nor U19124 (N_19124,N_18977,N_18876);
nor U19125 (N_19125,N_18551,N_18803);
xnor U19126 (N_19126,N_18968,N_18919);
and U19127 (N_19127,N_18926,N_18522);
and U19128 (N_19128,N_18889,N_18789);
or U19129 (N_19129,N_18779,N_18534);
nand U19130 (N_19130,N_18699,N_18701);
or U19131 (N_19131,N_18530,N_18986);
nand U19132 (N_19132,N_18796,N_18698);
or U19133 (N_19133,N_18549,N_18637);
nand U19134 (N_19134,N_18550,N_18839);
nand U19135 (N_19135,N_18643,N_18525);
or U19136 (N_19136,N_18772,N_18546);
or U19137 (N_19137,N_18928,N_18815);
nand U19138 (N_19138,N_18531,N_18613);
or U19139 (N_19139,N_18506,N_18845);
nand U19140 (N_19140,N_18883,N_18998);
or U19141 (N_19141,N_18513,N_18994);
or U19142 (N_19142,N_18620,N_18836);
nand U19143 (N_19143,N_18663,N_18911);
and U19144 (N_19144,N_18813,N_18678);
or U19145 (N_19145,N_18665,N_18776);
nand U19146 (N_19146,N_18745,N_18982);
nor U19147 (N_19147,N_18603,N_18967);
nor U19148 (N_19148,N_18906,N_18723);
and U19149 (N_19149,N_18560,N_18539);
nand U19150 (N_19150,N_18751,N_18738);
and U19151 (N_19151,N_18771,N_18762);
nor U19152 (N_19152,N_18969,N_18992);
xor U19153 (N_19153,N_18821,N_18882);
nor U19154 (N_19154,N_18538,N_18508);
nand U19155 (N_19155,N_18863,N_18913);
nand U19156 (N_19156,N_18595,N_18511);
nand U19157 (N_19157,N_18687,N_18795);
nor U19158 (N_19158,N_18559,N_18558);
nand U19159 (N_19159,N_18566,N_18502);
xnor U19160 (N_19160,N_18951,N_18877);
nand U19161 (N_19161,N_18747,N_18642);
or U19162 (N_19162,N_18598,N_18866);
nor U19163 (N_19163,N_18573,N_18978);
nand U19164 (N_19164,N_18582,N_18797);
and U19165 (N_19165,N_18775,N_18874);
nor U19166 (N_19166,N_18588,N_18529);
or U19167 (N_19167,N_18651,N_18523);
or U19168 (N_19168,N_18632,N_18734);
or U19169 (N_19169,N_18897,N_18755);
and U19170 (N_19170,N_18683,N_18640);
nor U19171 (N_19171,N_18636,N_18818);
nand U19172 (N_19172,N_18679,N_18659);
nor U19173 (N_19173,N_18540,N_18793);
and U19174 (N_19174,N_18710,N_18737);
nand U19175 (N_19175,N_18878,N_18885);
nor U19176 (N_19176,N_18545,N_18629);
and U19177 (N_19177,N_18965,N_18718);
nand U19178 (N_19178,N_18612,N_18851);
nor U19179 (N_19179,N_18570,N_18971);
and U19180 (N_19180,N_18767,N_18571);
or U19181 (N_19181,N_18853,N_18970);
xor U19182 (N_19182,N_18501,N_18924);
nor U19183 (N_19183,N_18670,N_18788);
nor U19184 (N_19184,N_18703,N_18940);
or U19185 (N_19185,N_18925,N_18556);
and U19186 (N_19186,N_18791,N_18741);
and U19187 (N_19187,N_18904,N_18857);
nor U19188 (N_19188,N_18754,N_18798);
nor U19189 (N_19189,N_18912,N_18936);
or U19190 (N_19190,N_18704,N_18920);
or U19191 (N_19191,N_18859,N_18983);
nand U19192 (N_19192,N_18770,N_18899);
and U19193 (N_19193,N_18831,N_18891);
or U19194 (N_19194,N_18625,N_18880);
or U19195 (N_19195,N_18567,N_18938);
and U19196 (N_19196,N_18668,N_18731);
or U19197 (N_19197,N_18930,N_18892);
or U19198 (N_19198,N_18896,N_18806);
nand U19199 (N_19199,N_18662,N_18726);
nand U19200 (N_19200,N_18955,N_18563);
or U19201 (N_19201,N_18753,N_18990);
nand U19202 (N_19202,N_18552,N_18694);
and U19203 (N_19203,N_18809,N_18648);
or U19204 (N_19204,N_18646,N_18808);
nor U19205 (N_19205,N_18900,N_18774);
nor U19206 (N_19206,N_18895,N_18939);
nor U19207 (N_19207,N_18794,N_18799);
or U19208 (N_19208,N_18828,N_18575);
nand U19209 (N_19209,N_18991,N_18623);
nand U19210 (N_19210,N_18946,N_18944);
nand U19211 (N_19211,N_18999,N_18750);
and U19212 (N_19212,N_18887,N_18561);
nand U19213 (N_19213,N_18903,N_18800);
nand U19214 (N_19214,N_18868,N_18645);
or U19215 (N_19215,N_18590,N_18607);
nand U19216 (N_19216,N_18873,N_18862);
or U19217 (N_19217,N_18832,N_18841);
and U19218 (N_19218,N_18742,N_18616);
nor U19219 (N_19219,N_18861,N_18500);
nand U19220 (N_19220,N_18909,N_18858);
nand U19221 (N_19221,N_18503,N_18773);
nor U19222 (N_19222,N_18765,N_18568);
or U19223 (N_19223,N_18633,N_18666);
or U19224 (N_19224,N_18521,N_18954);
nor U19225 (N_19225,N_18914,N_18812);
nor U19226 (N_19226,N_18824,N_18526);
nor U19227 (N_19227,N_18962,N_18961);
nor U19228 (N_19228,N_18608,N_18875);
nand U19229 (N_19229,N_18688,N_18719);
and U19230 (N_19230,N_18941,N_18810);
or U19231 (N_19231,N_18532,N_18927);
or U19232 (N_19232,N_18976,N_18953);
nand U19233 (N_19233,N_18860,N_18898);
nor U19234 (N_19234,N_18870,N_18987);
and U19235 (N_19235,N_18822,N_18937);
nand U19236 (N_19236,N_18695,N_18684);
nand U19237 (N_19237,N_18676,N_18537);
nor U19238 (N_19238,N_18778,N_18995);
nand U19239 (N_19239,N_18709,N_18605);
or U19240 (N_19240,N_18838,N_18685);
and U19241 (N_19241,N_18997,N_18536);
nand U19242 (N_19242,N_18849,N_18846);
nand U19243 (N_19243,N_18884,N_18655);
or U19244 (N_19244,N_18934,N_18943);
and U19245 (N_19245,N_18802,N_18609);
nor U19246 (N_19246,N_18604,N_18945);
and U19247 (N_19247,N_18621,N_18826);
or U19248 (N_19248,N_18504,N_18652);
or U19249 (N_19249,N_18850,N_18594);
nand U19250 (N_19250,N_18625,N_18929);
nand U19251 (N_19251,N_18864,N_18535);
or U19252 (N_19252,N_18568,N_18534);
nor U19253 (N_19253,N_18926,N_18931);
and U19254 (N_19254,N_18751,N_18589);
nor U19255 (N_19255,N_18942,N_18779);
and U19256 (N_19256,N_18839,N_18961);
nand U19257 (N_19257,N_18952,N_18515);
or U19258 (N_19258,N_18513,N_18962);
and U19259 (N_19259,N_18877,N_18801);
nor U19260 (N_19260,N_18829,N_18646);
and U19261 (N_19261,N_18984,N_18881);
or U19262 (N_19262,N_18950,N_18615);
nand U19263 (N_19263,N_18622,N_18986);
or U19264 (N_19264,N_18716,N_18929);
or U19265 (N_19265,N_18742,N_18589);
or U19266 (N_19266,N_18743,N_18919);
nand U19267 (N_19267,N_18716,N_18575);
or U19268 (N_19268,N_18683,N_18935);
or U19269 (N_19269,N_18823,N_18747);
nand U19270 (N_19270,N_18738,N_18762);
or U19271 (N_19271,N_18513,N_18986);
nor U19272 (N_19272,N_18506,N_18769);
nand U19273 (N_19273,N_18772,N_18585);
nor U19274 (N_19274,N_18679,N_18526);
or U19275 (N_19275,N_18833,N_18528);
and U19276 (N_19276,N_18743,N_18581);
nor U19277 (N_19277,N_18677,N_18843);
or U19278 (N_19278,N_18910,N_18828);
nand U19279 (N_19279,N_18955,N_18633);
nor U19280 (N_19280,N_18988,N_18607);
or U19281 (N_19281,N_18509,N_18516);
nand U19282 (N_19282,N_18623,N_18827);
nor U19283 (N_19283,N_18975,N_18963);
nor U19284 (N_19284,N_18802,N_18907);
nor U19285 (N_19285,N_18823,N_18768);
nor U19286 (N_19286,N_18771,N_18662);
or U19287 (N_19287,N_18907,N_18741);
or U19288 (N_19288,N_18544,N_18991);
nand U19289 (N_19289,N_18556,N_18901);
or U19290 (N_19290,N_18550,N_18617);
nand U19291 (N_19291,N_18644,N_18974);
or U19292 (N_19292,N_18902,N_18764);
nand U19293 (N_19293,N_18871,N_18969);
nand U19294 (N_19294,N_18959,N_18803);
nor U19295 (N_19295,N_18767,N_18609);
and U19296 (N_19296,N_18975,N_18741);
nand U19297 (N_19297,N_18777,N_18878);
and U19298 (N_19298,N_18784,N_18712);
nor U19299 (N_19299,N_18657,N_18865);
nand U19300 (N_19300,N_18735,N_18640);
and U19301 (N_19301,N_18764,N_18843);
or U19302 (N_19302,N_18981,N_18961);
nor U19303 (N_19303,N_18528,N_18662);
or U19304 (N_19304,N_18612,N_18954);
nor U19305 (N_19305,N_18840,N_18550);
nand U19306 (N_19306,N_18802,N_18807);
or U19307 (N_19307,N_18912,N_18866);
or U19308 (N_19308,N_18519,N_18957);
or U19309 (N_19309,N_18524,N_18729);
nor U19310 (N_19310,N_18530,N_18868);
nor U19311 (N_19311,N_18940,N_18999);
nand U19312 (N_19312,N_18789,N_18893);
nand U19313 (N_19313,N_18679,N_18852);
nor U19314 (N_19314,N_18669,N_18746);
and U19315 (N_19315,N_18925,N_18990);
nor U19316 (N_19316,N_18751,N_18798);
nor U19317 (N_19317,N_18958,N_18814);
and U19318 (N_19318,N_18797,N_18547);
nor U19319 (N_19319,N_18663,N_18609);
nand U19320 (N_19320,N_18846,N_18980);
nor U19321 (N_19321,N_18804,N_18679);
nand U19322 (N_19322,N_18970,N_18589);
nor U19323 (N_19323,N_18989,N_18722);
nor U19324 (N_19324,N_18743,N_18767);
nor U19325 (N_19325,N_18859,N_18610);
nand U19326 (N_19326,N_18518,N_18944);
and U19327 (N_19327,N_18829,N_18737);
and U19328 (N_19328,N_18727,N_18929);
and U19329 (N_19329,N_18638,N_18709);
nand U19330 (N_19330,N_18638,N_18893);
or U19331 (N_19331,N_18744,N_18566);
and U19332 (N_19332,N_18928,N_18989);
and U19333 (N_19333,N_18902,N_18830);
nand U19334 (N_19334,N_18627,N_18820);
and U19335 (N_19335,N_18648,N_18628);
nor U19336 (N_19336,N_18706,N_18882);
and U19337 (N_19337,N_18863,N_18725);
and U19338 (N_19338,N_18745,N_18718);
nand U19339 (N_19339,N_18855,N_18984);
nor U19340 (N_19340,N_18721,N_18593);
nor U19341 (N_19341,N_18871,N_18629);
or U19342 (N_19342,N_18536,N_18869);
nand U19343 (N_19343,N_18629,N_18846);
or U19344 (N_19344,N_18553,N_18932);
nor U19345 (N_19345,N_18573,N_18700);
and U19346 (N_19346,N_18719,N_18817);
xor U19347 (N_19347,N_18888,N_18968);
or U19348 (N_19348,N_18962,N_18949);
or U19349 (N_19349,N_18551,N_18574);
or U19350 (N_19350,N_18823,N_18588);
nor U19351 (N_19351,N_18576,N_18531);
nor U19352 (N_19352,N_18826,N_18961);
nor U19353 (N_19353,N_18620,N_18994);
or U19354 (N_19354,N_18574,N_18926);
and U19355 (N_19355,N_18903,N_18609);
nand U19356 (N_19356,N_18794,N_18969);
nor U19357 (N_19357,N_18901,N_18886);
or U19358 (N_19358,N_18989,N_18655);
or U19359 (N_19359,N_18867,N_18510);
nor U19360 (N_19360,N_18903,N_18912);
or U19361 (N_19361,N_18802,N_18946);
nor U19362 (N_19362,N_18631,N_18706);
nand U19363 (N_19363,N_18518,N_18585);
or U19364 (N_19364,N_18848,N_18757);
xnor U19365 (N_19365,N_18940,N_18590);
nand U19366 (N_19366,N_18843,N_18901);
or U19367 (N_19367,N_18621,N_18875);
nand U19368 (N_19368,N_18745,N_18545);
or U19369 (N_19369,N_18796,N_18644);
and U19370 (N_19370,N_18847,N_18778);
and U19371 (N_19371,N_18713,N_18754);
nor U19372 (N_19372,N_18809,N_18825);
or U19373 (N_19373,N_18697,N_18921);
nand U19374 (N_19374,N_18627,N_18657);
nand U19375 (N_19375,N_18878,N_18958);
nor U19376 (N_19376,N_18838,N_18689);
nand U19377 (N_19377,N_18657,N_18842);
xnor U19378 (N_19378,N_18642,N_18748);
nor U19379 (N_19379,N_18919,N_18730);
nor U19380 (N_19380,N_18507,N_18579);
nand U19381 (N_19381,N_18668,N_18717);
or U19382 (N_19382,N_18723,N_18942);
nand U19383 (N_19383,N_18821,N_18638);
or U19384 (N_19384,N_18863,N_18693);
nand U19385 (N_19385,N_18657,N_18633);
nand U19386 (N_19386,N_18866,N_18790);
or U19387 (N_19387,N_18836,N_18584);
nor U19388 (N_19388,N_18968,N_18596);
nor U19389 (N_19389,N_18921,N_18640);
or U19390 (N_19390,N_18792,N_18526);
and U19391 (N_19391,N_18726,N_18751);
or U19392 (N_19392,N_18602,N_18581);
nor U19393 (N_19393,N_18897,N_18966);
xor U19394 (N_19394,N_18522,N_18815);
nand U19395 (N_19395,N_18807,N_18982);
or U19396 (N_19396,N_18846,N_18732);
nand U19397 (N_19397,N_18563,N_18510);
or U19398 (N_19398,N_18755,N_18890);
nand U19399 (N_19399,N_18950,N_18857);
or U19400 (N_19400,N_18530,N_18901);
nor U19401 (N_19401,N_18828,N_18625);
nor U19402 (N_19402,N_18918,N_18834);
and U19403 (N_19403,N_18506,N_18793);
nor U19404 (N_19404,N_18776,N_18597);
and U19405 (N_19405,N_18592,N_18986);
or U19406 (N_19406,N_18931,N_18865);
and U19407 (N_19407,N_18617,N_18637);
nand U19408 (N_19408,N_18715,N_18654);
nand U19409 (N_19409,N_18991,N_18985);
and U19410 (N_19410,N_18905,N_18617);
and U19411 (N_19411,N_18625,N_18645);
nor U19412 (N_19412,N_18526,N_18897);
and U19413 (N_19413,N_18978,N_18697);
nand U19414 (N_19414,N_18970,N_18686);
and U19415 (N_19415,N_18673,N_18846);
or U19416 (N_19416,N_18527,N_18928);
nand U19417 (N_19417,N_18583,N_18558);
and U19418 (N_19418,N_18781,N_18744);
nand U19419 (N_19419,N_18665,N_18754);
and U19420 (N_19420,N_18775,N_18925);
nand U19421 (N_19421,N_18991,N_18851);
and U19422 (N_19422,N_18648,N_18555);
or U19423 (N_19423,N_18843,N_18742);
nand U19424 (N_19424,N_18807,N_18642);
and U19425 (N_19425,N_18647,N_18923);
and U19426 (N_19426,N_18572,N_18977);
or U19427 (N_19427,N_18618,N_18956);
and U19428 (N_19428,N_18609,N_18777);
nor U19429 (N_19429,N_18766,N_18775);
nor U19430 (N_19430,N_18760,N_18898);
or U19431 (N_19431,N_18871,N_18882);
or U19432 (N_19432,N_18835,N_18768);
xnor U19433 (N_19433,N_18706,N_18568);
xnor U19434 (N_19434,N_18767,N_18834);
nand U19435 (N_19435,N_18947,N_18928);
and U19436 (N_19436,N_18768,N_18672);
nand U19437 (N_19437,N_18803,N_18990);
or U19438 (N_19438,N_18607,N_18866);
xnor U19439 (N_19439,N_18752,N_18779);
nand U19440 (N_19440,N_18733,N_18878);
nand U19441 (N_19441,N_18967,N_18897);
nand U19442 (N_19442,N_18841,N_18574);
and U19443 (N_19443,N_18752,N_18662);
nand U19444 (N_19444,N_18748,N_18680);
and U19445 (N_19445,N_18754,N_18982);
xor U19446 (N_19446,N_18740,N_18798);
xnor U19447 (N_19447,N_18880,N_18799);
nor U19448 (N_19448,N_18503,N_18727);
nand U19449 (N_19449,N_18809,N_18718);
or U19450 (N_19450,N_18506,N_18969);
nor U19451 (N_19451,N_18968,N_18627);
and U19452 (N_19452,N_18932,N_18789);
or U19453 (N_19453,N_18528,N_18742);
and U19454 (N_19454,N_18754,N_18518);
or U19455 (N_19455,N_18569,N_18946);
or U19456 (N_19456,N_18683,N_18673);
nand U19457 (N_19457,N_18850,N_18515);
and U19458 (N_19458,N_18614,N_18546);
or U19459 (N_19459,N_18942,N_18768);
nor U19460 (N_19460,N_18662,N_18532);
and U19461 (N_19461,N_18555,N_18711);
nand U19462 (N_19462,N_18622,N_18803);
nor U19463 (N_19463,N_18823,N_18887);
nand U19464 (N_19464,N_18509,N_18898);
nand U19465 (N_19465,N_18773,N_18677);
nor U19466 (N_19466,N_18559,N_18581);
and U19467 (N_19467,N_18816,N_18576);
and U19468 (N_19468,N_18663,N_18661);
or U19469 (N_19469,N_18775,N_18515);
nor U19470 (N_19470,N_18979,N_18838);
and U19471 (N_19471,N_18619,N_18522);
nor U19472 (N_19472,N_18653,N_18584);
nand U19473 (N_19473,N_18602,N_18617);
nor U19474 (N_19474,N_18886,N_18658);
nand U19475 (N_19475,N_18514,N_18624);
nand U19476 (N_19476,N_18773,N_18750);
or U19477 (N_19477,N_18879,N_18761);
nor U19478 (N_19478,N_18640,N_18527);
nand U19479 (N_19479,N_18700,N_18978);
nor U19480 (N_19480,N_18829,N_18792);
nor U19481 (N_19481,N_18505,N_18898);
and U19482 (N_19482,N_18803,N_18788);
and U19483 (N_19483,N_18630,N_18910);
nand U19484 (N_19484,N_18911,N_18759);
nor U19485 (N_19485,N_18853,N_18851);
or U19486 (N_19486,N_18846,N_18865);
nor U19487 (N_19487,N_18518,N_18928);
or U19488 (N_19488,N_18776,N_18788);
or U19489 (N_19489,N_18930,N_18935);
and U19490 (N_19490,N_18875,N_18563);
and U19491 (N_19491,N_18541,N_18582);
and U19492 (N_19492,N_18747,N_18846);
nand U19493 (N_19493,N_18641,N_18755);
nand U19494 (N_19494,N_18738,N_18995);
nand U19495 (N_19495,N_18698,N_18968);
or U19496 (N_19496,N_18540,N_18908);
nor U19497 (N_19497,N_18930,N_18678);
or U19498 (N_19498,N_18743,N_18869);
nor U19499 (N_19499,N_18590,N_18713);
nor U19500 (N_19500,N_19026,N_19107);
and U19501 (N_19501,N_19486,N_19498);
and U19502 (N_19502,N_19351,N_19074);
nand U19503 (N_19503,N_19173,N_19328);
nand U19504 (N_19504,N_19284,N_19411);
and U19505 (N_19505,N_19196,N_19242);
nor U19506 (N_19506,N_19233,N_19128);
and U19507 (N_19507,N_19169,N_19245);
nand U19508 (N_19508,N_19300,N_19014);
and U19509 (N_19509,N_19135,N_19036);
or U19510 (N_19510,N_19260,N_19216);
and U19511 (N_19511,N_19151,N_19327);
or U19512 (N_19512,N_19046,N_19203);
nor U19513 (N_19513,N_19329,N_19377);
or U19514 (N_19514,N_19413,N_19341);
nand U19515 (N_19515,N_19332,N_19273);
or U19516 (N_19516,N_19405,N_19215);
or U19517 (N_19517,N_19061,N_19314);
and U19518 (N_19518,N_19186,N_19223);
xnor U19519 (N_19519,N_19194,N_19287);
nor U19520 (N_19520,N_19193,N_19356);
nor U19521 (N_19521,N_19491,N_19100);
or U19522 (N_19522,N_19043,N_19362);
nor U19523 (N_19523,N_19392,N_19333);
nand U19524 (N_19524,N_19433,N_19032);
or U19525 (N_19525,N_19040,N_19146);
nor U19526 (N_19526,N_19481,N_19117);
and U19527 (N_19527,N_19134,N_19141);
nor U19528 (N_19528,N_19105,N_19293);
and U19529 (N_19529,N_19072,N_19275);
nand U19530 (N_19530,N_19452,N_19222);
and U19531 (N_19531,N_19276,N_19109);
and U19532 (N_19532,N_19289,N_19115);
or U19533 (N_19533,N_19165,N_19339);
or U19534 (N_19534,N_19160,N_19023);
and U19535 (N_19535,N_19005,N_19375);
or U19536 (N_19536,N_19379,N_19248);
and U19537 (N_19537,N_19201,N_19398);
nand U19538 (N_19538,N_19097,N_19084);
nor U19539 (N_19539,N_19118,N_19095);
and U19540 (N_19540,N_19306,N_19038);
nand U19541 (N_19541,N_19073,N_19258);
and U19542 (N_19542,N_19080,N_19261);
or U19543 (N_19543,N_19060,N_19153);
or U19544 (N_19544,N_19385,N_19085);
nand U19545 (N_19545,N_19003,N_19054);
nor U19546 (N_19546,N_19133,N_19441);
or U19547 (N_19547,N_19378,N_19069);
nor U19548 (N_19548,N_19471,N_19253);
nor U19549 (N_19549,N_19137,N_19006);
nor U19550 (N_19550,N_19156,N_19464);
nor U19551 (N_19551,N_19438,N_19171);
or U19552 (N_19552,N_19182,N_19221);
nand U19553 (N_19553,N_19076,N_19047);
nor U19554 (N_19554,N_19412,N_19466);
and U19555 (N_19555,N_19318,N_19265);
nor U19556 (N_19556,N_19124,N_19359);
nor U19557 (N_19557,N_19334,N_19031);
and U19558 (N_19558,N_19145,N_19219);
nor U19559 (N_19559,N_19150,N_19346);
and U19560 (N_19560,N_19094,N_19390);
or U19561 (N_19561,N_19282,N_19394);
nand U19562 (N_19562,N_19159,N_19475);
nand U19563 (N_19563,N_19051,N_19338);
and U19564 (N_19564,N_19192,N_19088);
nor U19565 (N_19565,N_19168,N_19179);
or U19566 (N_19566,N_19373,N_19343);
and U19567 (N_19567,N_19406,N_19229);
and U19568 (N_19568,N_19497,N_19191);
nand U19569 (N_19569,N_19052,N_19417);
or U19570 (N_19570,N_19075,N_19310);
nor U19571 (N_19571,N_19008,N_19366);
or U19572 (N_19572,N_19017,N_19015);
nor U19573 (N_19573,N_19234,N_19102);
or U19574 (N_19574,N_19232,N_19161);
or U19575 (N_19575,N_19185,N_19446);
and U19576 (N_19576,N_19030,N_19344);
and U19577 (N_19577,N_19345,N_19309);
nand U19578 (N_19578,N_19029,N_19382);
or U19579 (N_19579,N_19132,N_19313);
nor U19580 (N_19580,N_19199,N_19254);
or U19581 (N_19581,N_19138,N_19064);
or U19582 (N_19582,N_19285,N_19025);
nor U19583 (N_19583,N_19077,N_19045);
nor U19584 (N_19584,N_19434,N_19494);
or U19585 (N_19585,N_19093,N_19127);
or U19586 (N_19586,N_19236,N_19478);
nand U19587 (N_19587,N_19206,N_19140);
nand U19588 (N_19588,N_19391,N_19055);
nor U19589 (N_19589,N_19268,N_19407);
and U19590 (N_19590,N_19208,N_19224);
or U19591 (N_19591,N_19263,N_19112);
nand U19592 (N_19592,N_19099,N_19249);
nor U19593 (N_19593,N_19322,N_19239);
and U19594 (N_19594,N_19420,N_19279);
or U19595 (N_19595,N_19469,N_19148);
nand U19596 (N_19596,N_19188,N_19241);
nor U19597 (N_19597,N_19350,N_19483);
nor U19598 (N_19598,N_19057,N_19070);
and U19599 (N_19599,N_19496,N_19335);
or U19600 (N_19600,N_19337,N_19308);
nor U19601 (N_19601,N_19000,N_19012);
and U19602 (N_19602,N_19266,N_19207);
and U19603 (N_19603,N_19035,N_19280);
nand U19604 (N_19604,N_19299,N_19317);
nor U19605 (N_19605,N_19103,N_19376);
and U19606 (N_19606,N_19493,N_19489);
or U19607 (N_19607,N_19319,N_19217);
nand U19608 (N_19608,N_19430,N_19078);
nor U19609 (N_19609,N_19157,N_19324);
and U19610 (N_19610,N_19399,N_19119);
nand U19611 (N_19611,N_19467,N_19068);
nand U19612 (N_19612,N_19360,N_19101);
or U19613 (N_19613,N_19416,N_19455);
or U19614 (N_19614,N_19301,N_19321);
or U19615 (N_19615,N_19062,N_19142);
or U19616 (N_19616,N_19291,N_19041);
nor U19617 (N_19617,N_19357,N_19149);
or U19618 (N_19618,N_19020,N_19154);
and U19619 (N_19619,N_19415,N_19414);
and U19620 (N_19620,N_19401,N_19437);
or U19621 (N_19621,N_19473,N_19247);
nor U19622 (N_19622,N_19108,N_19086);
and U19623 (N_19623,N_19459,N_19380);
or U19624 (N_19624,N_19294,N_19479);
or U19625 (N_19625,N_19250,N_19476);
or U19626 (N_19626,N_19002,N_19226);
or U19627 (N_19627,N_19243,N_19065);
xor U19628 (N_19628,N_19358,N_19238);
or U19629 (N_19629,N_19004,N_19288);
nor U19630 (N_19630,N_19180,N_19364);
or U19631 (N_19631,N_19298,N_19393);
nor U19632 (N_19632,N_19336,N_19458);
nand U19633 (N_19633,N_19384,N_19125);
nand U19634 (N_19634,N_19011,N_19063);
xnor U19635 (N_19635,N_19442,N_19488);
nor U19636 (N_19636,N_19058,N_19400);
and U19637 (N_19637,N_19034,N_19425);
nand U19638 (N_19638,N_19435,N_19286);
nand U19639 (N_19639,N_19059,N_19255);
or U19640 (N_19640,N_19499,N_19089);
or U19641 (N_19641,N_19304,N_19272);
and U19642 (N_19642,N_19492,N_19120);
nand U19643 (N_19643,N_19244,N_19303);
or U19644 (N_19644,N_19262,N_19202);
and U19645 (N_19645,N_19044,N_19079);
or U19646 (N_19646,N_19482,N_19198);
and U19647 (N_19647,N_19422,N_19205);
or U19648 (N_19648,N_19370,N_19418);
nand U19649 (N_19649,N_19451,N_19371);
and U19650 (N_19650,N_19106,N_19315);
nand U19651 (N_19651,N_19450,N_19197);
and U19652 (N_19652,N_19470,N_19374);
or U19653 (N_19653,N_19009,N_19122);
or U19654 (N_19654,N_19028,N_19147);
and U19655 (N_19655,N_19409,N_19001);
or U19656 (N_19656,N_19090,N_19410);
and U19657 (N_19657,N_19311,N_19177);
nand U19658 (N_19658,N_19449,N_19252);
and U19659 (N_19659,N_19155,N_19210);
and U19660 (N_19660,N_19227,N_19269);
nand U19661 (N_19661,N_19386,N_19305);
nor U19662 (N_19662,N_19050,N_19123);
nand U19663 (N_19663,N_19214,N_19428);
nor U19664 (N_19664,N_19440,N_19381);
or U19665 (N_19665,N_19126,N_19307);
nand U19666 (N_19666,N_19421,N_19419);
or U19667 (N_19667,N_19013,N_19111);
nor U19668 (N_19668,N_19424,N_19104);
or U19669 (N_19669,N_19240,N_19457);
nor U19670 (N_19670,N_19181,N_19274);
and U19671 (N_19671,N_19316,N_19408);
and U19672 (N_19672,N_19018,N_19027);
nor U19673 (N_19673,N_19039,N_19448);
or U19674 (N_19674,N_19235,N_19368);
or U19675 (N_19675,N_19264,N_19485);
or U19676 (N_19676,N_19083,N_19130);
nor U19677 (N_19677,N_19016,N_19453);
and U19678 (N_19678,N_19369,N_19228);
or U19679 (N_19679,N_19162,N_19436);
and U19680 (N_19680,N_19049,N_19302);
and U19681 (N_19681,N_19195,N_19152);
nand U19682 (N_19682,N_19454,N_19048);
and U19683 (N_19683,N_19267,N_19220);
and U19684 (N_19684,N_19423,N_19183);
and U19685 (N_19685,N_19121,N_19067);
and U19686 (N_19686,N_19347,N_19429);
and U19687 (N_19687,N_19212,N_19447);
and U19688 (N_19688,N_19456,N_19432);
and U19689 (N_19689,N_19404,N_19353);
nand U19690 (N_19690,N_19087,N_19204);
nand U19691 (N_19691,N_19431,N_19403);
and U19692 (N_19692,N_19445,N_19396);
and U19693 (N_19693,N_19166,N_19022);
nand U19694 (N_19694,N_19184,N_19024);
nand U19695 (N_19695,N_19037,N_19211);
and U19696 (N_19696,N_19129,N_19033);
and U19697 (N_19697,N_19365,N_19395);
or U19698 (N_19698,N_19139,N_19209);
and U19699 (N_19699,N_19271,N_19426);
nand U19700 (N_19700,N_19474,N_19389);
nand U19701 (N_19701,N_19487,N_19320);
and U19702 (N_19702,N_19256,N_19277);
nand U19703 (N_19703,N_19163,N_19091);
or U19704 (N_19704,N_19477,N_19427);
nand U19705 (N_19705,N_19495,N_19355);
and U19706 (N_19706,N_19331,N_19251);
nand U19707 (N_19707,N_19463,N_19113);
and U19708 (N_19708,N_19397,N_19439);
nor U19709 (N_19709,N_19352,N_19213);
or U19710 (N_19710,N_19292,N_19189);
and U19711 (N_19711,N_19326,N_19257);
nand U19712 (N_19712,N_19278,N_19172);
nand U19713 (N_19713,N_19167,N_19174);
or U19714 (N_19714,N_19462,N_19175);
and U19715 (N_19715,N_19114,N_19468);
nand U19716 (N_19716,N_19187,N_19131);
or U19717 (N_19717,N_19281,N_19472);
nor U19718 (N_19718,N_19071,N_19021);
and U19719 (N_19719,N_19231,N_19290);
nor U19720 (N_19720,N_19342,N_19053);
nor U19721 (N_19721,N_19349,N_19270);
or U19722 (N_19722,N_19007,N_19340);
nor U19723 (N_19723,N_19295,N_19312);
and U19724 (N_19724,N_19010,N_19372);
nor U19725 (N_19725,N_19170,N_19297);
or U19726 (N_19726,N_19387,N_19383);
or U19727 (N_19727,N_19283,N_19460);
and U19728 (N_19728,N_19480,N_19096);
and U19729 (N_19729,N_19143,N_19361);
and U19730 (N_19730,N_19081,N_19190);
nor U19731 (N_19731,N_19323,N_19144);
or U19732 (N_19732,N_19230,N_19158);
nor U19733 (N_19733,N_19176,N_19042);
and U19734 (N_19734,N_19237,N_19461);
or U19735 (N_19735,N_19110,N_19225);
or U19736 (N_19736,N_19367,N_19098);
and U19737 (N_19737,N_19465,N_19443);
nor U19738 (N_19738,N_19348,N_19218);
and U19739 (N_19739,N_19363,N_19164);
xor U19740 (N_19740,N_19066,N_19056);
or U19741 (N_19741,N_19200,N_19330);
nor U19742 (N_19742,N_19388,N_19296);
or U19743 (N_19743,N_19116,N_19092);
or U19744 (N_19744,N_19019,N_19246);
nor U19745 (N_19745,N_19325,N_19082);
nor U19746 (N_19746,N_19354,N_19402);
or U19747 (N_19747,N_19178,N_19490);
or U19748 (N_19748,N_19484,N_19259);
nor U19749 (N_19749,N_19136,N_19444);
and U19750 (N_19750,N_19381,N_19027);
nand U19751 (N_19751,N_19321,N_19400);
xnor U19752 (N_19752,N_19265,N_19040);
nand U19753 (N_19753,N_19291,N_19485);
or U19754 (N_19754,N_19366,N_19059);
or U19755 (N_19755,N_19007,N_19301);
and U19756 (N_19756,N_19372,N_19163);
nand U19757 (N_19757,N_19382,N_19033);
nor U19758 (N_19758,N_19233,N_19319);
nor U19759 (N_19759,N_19467,N_19340);
nor U19760 (N_19760,N_19095,N_19479);
or U19761 (N_19761,N_19194,N_19211);
nor U19762 (N_19762,N_19159,N_19424);
and U19763 (N_19763,N_19040,N_19372);
nor U19764 (N_19764,N_19256,N_19250);
nand U19765 (N_19765,N_19414,N_19062);
or U19766 (N_19766,N_19196,N_19234);
and U19767 (N_19767,N_19111,N_19487);
and U19768 (N_19768,N_19025,N_19080);
nor U19769 (N_19769,N_19495,N_19265);
or U19770 (N_19770,N_19141,N_19232);
or U19771 (N_19771,N_19335,N_19304);
nor U19772 (N_19772,N_19496,N_19403);
nor U19773 (N_19773,N_19031,N_19197);
or U19774 (N_19774,N_19093,N_19475);
or U19775 (N_19775,N_19456,N_19194);
or U19776 (N_19776,N_19470,N_19492);
nor U19777 (N_19777,N_19110,N_19209);
nor U19778 (N_19778,N_19457,N_19027);
or U19779 (N_19779,N_19191,N_19030);
nor U19780 (N_19780,N_19194,N_19251);
nand U19781 (N_19781,N_19426,N_19498);
nand U19782 (N_19782,N_19461,N_19378);
nand U19783 (N_19783,N_19445,N_19298);
nor U19784 (N_19784,N_19096,N_19328);
or U19785 (N_19785,N_19051,N_19154);
nor U19786 (N_19786,N_19004,N_19256);
and U19787 (N_19787,N_19344,N_19224);
nand U19788 (N_19788,N_19407,N_19240);
or U19789 (N_19789,N_19310,N_19091);
or U19790 (N_19790,N_19201,N_19226);
and U19791 (N_19791,N_19271,N_19200);
nand U19792 (N_19792,N_19476,N_19377);
or U19793 (N_19793,N_19351,N_19035);
or U19794 (N_19794,N_19000,N_19072);
nor U19795 (N_19795,N_19067,N_19112);
or U19796 (N_19796,N_19132,N_19191);
nand U19797 (N_19797,N_19463,N_19341);
or U19798 (N_19798,N_19195,N_19376);
nor U19799 (N_19799,N_19485,N_19072);
nor U19800 (N_19800,N_19062,N_19214);
or U19801 (N_19801,N_19464,N_19467);
or U19802 (N_19802,N_19353,N_19084);
or U19803 (N_19803,N_19377,N_19078);
and U19804 (N_19804,N_19222,N_19257);
nand U19805 (N_19805,N_19252,N_19255);
nor U19806 (N_19806,N_19079,N_19085);
or U19807 (N_19807,N_19036,N_19010);
and U19808 (N_19808,N_19218,N_19293);
and U19809 (N_19809,N_19268,N_19119);
nand U19810 (N_19810,N_19243,N_19484);
xnor U19811 (N_19811,N_19143,N_19046);
or U19812 (N_19812,N_19000,N_19425);
nor U19813 (N_19813,N_19473,N_19197);
and U19814 (N_19814,N_19196,N_19036);
nor U19815 (N_19815,N_19298,N_19405);
nor U19816 (N_19816,N_19386,N_19070);
and U19817 (N_19817,N_19444,N_19331);
or U19818 (N_19818,N_19326,N_19367);
and U19819 (N_19819,N_19149,N_19496);
nor U19820 (N_19820,N_19139,N_19340);
or U19821 (N_19821,N_19465,N_19131);
nor U19822 (N_19822,N_19319,N_19349);
and U19823 (N_19823,N_19401,N_19099);
and U19824 (N_19824,N_19369,N_19144);
nand U19825 (N_19825,N_19014,N_19192);
nor U19826 (N_19826,N_19138,N_19050);
and U19827 (N_19827,N_19257,N_19418);
or U19828 (N_19828,N_19240,N_19318);
nand U19829 (N_19829,N_19083,N_19305);
nor U19830 (N_19830,N_19420,N_19474);
nand U19831 (N_19831,N_19064,N_19386);
and U19832 (N_19832,N_19253,N_19009);
or U19833 (N_19833,N_19498,N_19334);
nand U19834 (N_19834,N_19171,N_19302);
and U19835 (N_19835,N_19398,N_19354);
or U19836 (N_19836,N_19102,N_19402);
nand U19837 (N_19837,N_19128,N_19167);
or U19838 (N_19838,N_19342,N_19428);
nor U19839 (N_19839,N_19283,N_19035);
and U19840 (N_19840,N_19236,N_19336);
nor U19841 (N_19841,N_19227,N_19140);
or U19842 (N_19842,N_19414,N_19309);
or U19843 (N_19843,N_19242,N_19022);
and U19844 (N_19844,N_19015,N_19069);
nand U19845 (N_19845,N_19421,N_19048);
or U19846 (N_19846,N_19172,N_19332);
nor U19847 (N_19847,N_19458,N_19355);
nand U19848 (N_19848,N_19058,N_19417);
and U19849 (N_19849,N_19202,N_19291);
or U19850 (N_19850,N_19121,N_19430);
or U19851 (N_19851,N_19361,N_19015);
and U19852 (N_19852,N_19110,N_19186);
nand U19853 (N_19853,N_19314,N_19203);
and U19854 (N_19854,N_19254,N_19018);
or U19855 (N_19855,N_19263,N_19059);
and U19856 (N_19856,N_19036,N_19414);
nor U19857 (N_19857,N_19365,N_19116);
nor U19858 (N_19858,N_19437,N_19471);
xnor U19859 (N_19859,N_19043,N_19178);
or U19860 (N_19860,N_19219,N_19263);
nand U19861 (N_19861,N_19366,N_19268);
nand U19862 (N_19862,N_19042,N_19131);
nor U19863 (N_19863,N_19176,N_19415);
nor U19864 (N_19864,N_19242,N_19006);
or U19865 (N_19865,N_19284,N_19312);
nand U19866 (N_19866,N_19208,N_19268);
and U19867 (N_19867,N_19132,N_19404);
and U19868 (N_19868,N_19262,N_19479);
nand U19869 (N_19869,N_19099,N_19012);
nand U19870 (N_19870,N_19204,N_19367);
or U19871 (N_19871,N_19271,N_19014);
nand U19872 (N_19872,N_19123,N_19223);
xor U19873 (N_19873,N_19035,N_19077);
nand U19874 (N_19874,N_19472,N_19312);
nor U19875 (N_19875,N_19429,N_19360);
nor U19876 (N_19876,N_19422,N_19248);
nand U19877 (N_19877,N_19124,N_19498);
nand U19878 (N_19878,N_19075,N_19320);
nor U19879 (N_19879,N_19231,N_19480);
nor U19880 (N_19880,N_19109,N_19070);
nor U19881 (N_19881,N_19283,N_19286);
or U19882 (N_19882,N_19335,N_19431);
and U19883 (N_19883,N_19155,N_19198);
or U19884 (N_19884,N_19477,N_19144);
or U19885 (N_19885,N_19000,N_19097);
or U19886 (N_19886,N_19285,N_19255);
xnor U19887 (N_19887,N_19363,N_19019);
or U19888 (N_19888,N_19231,N_19456);
or U19889 (N_19889,N_19077,N_19036);
nor U19890 (N_19890,N_19154,N_19339);
or U19891 (N_19891,N_19497,N_19408);
or U19892 (N_19892,N_19432,N_19229);
nand U19893 (N_19893,N_19110,N_19413);
or U19894 (N_19894,N_19027,N_19214);
nand U19895 (N_19895,N_19128,N_19312);
nor U19896 (N_19896,N_19298,N_19435);
or U19897 (N_19897,N_19079,N_19312);
or U19898 (N_19898,N_19349,N_19162);
nor U19899 (N_19899,N_19105,N_19412);
nand U19900 (N_19900,N_19214,N_19208);
and U19901 (N_19901,N_19181,N_19295);
nand U19902 (N_19902,N_19460,N_19189);
and U19903 (N_19903,N_19201,N_19165);
xnor U19904 (N_19904,N_19424,N_19288);
nand U19905 (N_19905,N_19304,N_19456);
or U19906 (N_19906,N_19242,N_19350);
nor U19907 (N_19907,N_19322,N_19157);
nand U19908 (N_19908,N_19285,N_19233);
and U19909 (N_19909,N_19307,N_19343);
and U19910 (N_19910,N_19047,N_19451);
nor U19911 (N_19911,N_19257,N_19251);
or U19912 (N_19912,N_19043,N_19380);
or U19913 (N_19913,N_19149,N_19211);
or U19914 (N_19914,N_19498,N_19487);
nand U19915 (N_19915,N_19071,N_19358);
or U19916 (N_19916,N_19184,N_19308);
nor U19917 (N_19917,N_19405,N_19392);
or U19918 (N_19918,N_19035,N_19495);
and U19919 (N_19919,N_19167,N_19057);
or U19920 (N_19920,N_19155,N_19331);
nand U19921 (N_19921,N_19103,N_19004);
or U19922 (N_19922,N_19245,N_19052);
nor U19923 (N_19923,N_19481,N_19351);
and U19924 (N_19924,N_19235,N_19206);
nand U19925 (N_19925,N_19103,N_19020);
nand U19926 (N_19926,N_19209,N_19372);
nor U19927 (N_19927,N_19208,N_19261);
and U19928 (N_19928,N_19341,N_19488);
nor U19929 (N_19929,N_19009,N_19139);
nor U19930 (N_19930,N_19393,N_19386);
nand U19931 (N_19931,N_19368,N_19334);
nand U19932 (N_19932,N_19428,N_19270);
or U19933 (N_19933,N_19350,N_19351);
nor U19934 (N_19934,N_19099,N_19392);
nand U19935 (N_19935,N_19197,N_19278);
or U19936 (N_19936,N_19456,N_19433);
and U19937 (N_19937,N_19415,N_19216);
or U19938 (N_19938,N_19104,N_19224);
or U19939 (N_19939,N_19147,N_19272);
and U19940 (N_19940,N_19458,N_19013);
nor U19941 (N_19941,N_19336,N_19400);
or U19942 (N_19942,N_19456,N_19070);
and U19943 (N_19943,N_19178,N_19242);
or U19944 (N_19944,N_19469,N_19353);
nand U19945 (N_19945,N_19087,N_19430);
or U19946 (N_19946,N_19320,N_19020);
or U19947 (N_19947,N_19236,N_19215);
nor U19948 (N_19948,N_19180,N_19083);
nand U19949 (N_19949,N_19342,N_19196);
and U19950 (N_19950,N_19029,N_19020);
and U19951 (N_19951,N_19225,N_19329);
or U19952 (N_19952,N_19448,N_19172);
or U19953 (N_19953,N_19290,N_19237);
and U19954 (N_19954,N_19227,N_19196);
nor U19955 (N_19955,N_19174,N_19186);
or U19956 (N_19956,N_19327,N_19120);
and U19957 (N_19957,N_19083,N_19404);
nand U19958 (N_19958,N_19287,N_19263);
or U19959 (N_19959,N_19493,N_19472);
nor U19960 (N_19960,N_19346,N_19297);
and U19961 (N_19961,N_19209,N_19320);
or U19962 (N_19962,N_19486,N_19449);
or U19963 (N_19963,N_19097,N_19483);
xnor U19964 (N_19964,N_19143,N_19389);
and U19965 (N_19965,N_19381,N_19213);
nor U19966 (N_19966,N_19123,N_19032);
nor U19967 (N_19967,N_19141,N_19392);
and U19968 (N_19968,N_19487,N_19286);
nand U19969 (N_19969,N_19249,N_19193);
nand U19970 (N_19970,N_19273,N_19230);
or U19971 (N_19971,N_19441,N_19251);
nor U19972 (N_19972,N_19420,N_19337);
nand U19973 (N_19973,N_19453,N_19068);
and U19974 (N_19974,N_19473,N_19339);
nand U19975 (N_19975,N_19345,N_19046);
or U19976 (N_19976,N_19150,N_19341);
nor U19977 (N_19977,N_19236,N_19057);
and U19978 (N_19978,N_19043,N_19034);
or U19979 (N_19979,N_19014,N_19011);
and U19980 (N_19980,N_19473,N_19043);
nor U19981 (N_19981,N_19335,N_19468);
and U19982 (N_19982,N_19395,N_19343);
or U19983 (N_19983,N_19175,N_19130);
nand U19984 (N_19984,N_19036,N_19338);
nand U19985 (N_19985,N_19186,N_19309);
or U19986 (N_19986,N_19499,N_19228);
nand U19987 (N_19987,N_19080,N_19206);
nand U19988 (N_19988,N_19071,N_19008);
nor U19989 (N_19989,N_19083,N_19216);
and U19990 (N_19990,N_19186,N_19429);
and U19991 (N_19991,N_19110,N_19134);
and U19992 (N_19992,N_19255,N_19193);
nor U19993 (N_19993,N_19005,N_19408);
or U19994 (N_19994,N_19152,N_19493);
and U19995 (N_19995,N_19270,N_19245);
nor U19996 (N_19996,N_19087,N_19471);
nor U19997 (N_19997,N_19323,N_19206);
nand U19998 (N_19998,N_19076,N_19409);
nand U19999 (N_19999,N_19104,N_19059);
nor UO_0 (O_0,N_19984,N_19973);
or UO_1 (O_1,N_19866,N_19502);
nor UO_2 (O_2,N_19954,N_19903);
and UO_3 (O_3,N_19615,N_19743);
nand UO_4 (O_4,N_19588,N_19914);
nor UO_5 (O_5,N_19891,N_19970);
nand UO_6 (O_6,N_19799,N_19688);
or UO_7 (O_7,N_19907,N_19992);
nor UO_8 (O_8,N_19553,N_19854);
nor UO_9 (O_9,N_19978,N_19771);
xnor UO_10 (O_10,N_19845,N_19796);
and UO_11 (O_11,N_19751,N_19892);
or UO_12 (O_12,N_19780,N_19597);
or UO_13 (O_13,N_19718,N_19506);
xnor UO_14 (O_14,N_19749,N_19721);
and UO_15 (O_15,N_19827,N_19856);
or UO_16 (O_16,N_19852,N_19693);
nand UO_17 (O_17,N_19662,N_19871);
or UO_18 (O_18,N_19608,N_19574);
nand UO_19 (O_19,N_19637,N_19929);
or UO_20 (O_20,N_19791,N_19740);
nor UO_21 (O_21,N_19863,N_19556);
nand UO_22 (O_22,N_19772,N_19858);
nor UO_23 (O_23,N_19724,N_19834);
or UO_24 (O_24,N_19777,N_19619);
or UO_25 (O_25,N_19513,N_19938);
or UO_26 (O_26,N_19756,N_19861);
or UO_27 (O_27,N_19561,N_19514);
or UO_28 (O_28,N_19562,N_19638);
and UO_29 (O_29,N_19889,N_19609);
or UO_30 (O_30,N_19813,N_19784);
nand UO_31 (O_31,N_19642,N_19682);
nand UO_32 (O_32,N_19744,N_19872);
nor UO_33 (O_33,N_19501,N_19713);
nand UO_34 (O_34,N_19580,N_19916);
nand UO_35 (O_35,N_19648,N_19905);
nand UO_36 (O_36,N_19729,N_19764);
or UO_37 (O_37,N_19692,N_19899);
nor UO_38 (O_38,N_19516,N_19686);
or UO_39 (O_39,N_19994,N_19860);
nor UO_40 (O_40,N_19599,N_19538);
xnor UO_41 (O_41,N_19699,N_19928);
nor UO_42 (O_42,N_19723,N_19785);
nand UO_43 (O_43,N_19865,N_19656);
and UO_44 (O_44,N_19618,N_19974);
nand UO_45 (O_45,N_19894,N_19714);
and UO_46 (O_46,N_19816,N_19635);
and UO_47 (O_47,N_19893,N_19874);
and UO_48 (O_48,N_19951,N_19802);
xnor UO_49 (O_49,N_19722,N_19590);
nor UO_50 (O_50,N_19977,N_19946);
or UO_51 (O_51,N_19783,N_19947);
or UO_52 (O_52,N_19843,N_19508);
nand UO_53 (O_53,N_19825,N_19917);
nor UO_54 (O_54,N_19848,N_19939);
nand UO_55 (O_55,N_19518,N_19776);
nor UO_56 (O_56,N_19684,N_19525);
nand UO_57 (O_57,N_19696,N_19617);
and UO_58 (O_58,N_19822,N_19655);
or UO_59 (O_59,N_19697,N_19775);
and UO_60 (O_60,N_19896,N_19633);
nor UO_61 (O_61,N_19587,N_19622);
or UO_62 (O_62,N_19812,N_19541);
nand UO_63 (O_63,N_19959,N_19924);
nor UO_64 (O_64,N_19968,N_19997);
xor UO_65 (O_65,N_19647,N_19624);
nand UO_66 (O_66,N_19906,N_19673);
nor UO_67 (O_67,N_19550,N_19880);
and UO_68 (O_68,N_19826,N_19859);
or UO_69 (O_69,N_19850,N_19639);
nor UO_70 (O_70,N_19991,N_19895);
and UO_71 (O_71,N_19794,N_19763);
nor UO_72 (O_72,N_19629,N_19886);
or UO_73 (O_73,N_19593,N_19643);
or UO_74 (O_74,N_19930,N_19942);
nor UO_75 (O_75,N_19671,N_19793);
or UO_76 (O_76,N_19566,N_19922);
and UO_77 (O_77,N_19702,N_19589);
nand UO_78 (O_78,N_19950,N_19870);
nand UO_79 (O_79,N_19909,N_19654);
xnor UO_80 (O_80,N_19512,N_19757);
nand UO_81 (O_81,N_19890,N_19980);
nand UO_82 (O_82,N_19539,N_19831);
nor UO_83 (O_83,N_19604,N_19517);
nand UO_84 (O_84,N_19705,N_19641);
and UO_85 (O_85,N_19613,N_19944);
nand UO_86 (O_86,N_19616,N_19990);
or UO_87 (O_87,N_19754,N_19681);
nor UO_88 (O_88,N_19547,N_19811);
and UO_89 (O_89,N_19703,N_19867);
nor UO_90 (O_90,N_19943,N_19901);
nor UO_91 (O_91,N_19979,N_19701);
nor UO_92 (O_92,N_19555,N_19717);
nand UO_93 (O_93,N_19611,N_19962);
and UO_94 (O_94,N_19601,N_19592);
or UO_95 (O_95,N_19832,N_19864);
or UO_96 (O_96,N_19948,N_19623);
and UO_97 (O_97,N_19996,N_19716);
nand UO_98 (O_98,N_19570,N_19885);
nor UO_99 (O_99,N_19698,N_19529);
or UO_100 (O_100,N_19934,N_19963);
nor UO_101 (O_101,N_19847,N_19900);
nor UO_102 (O_102,N_19505,N_19614);
or UO_103 (O_103,N_19746,N_19607);
xor UO_104 (O_104,N_19621,N_19840);
nand UO_105 (O_105,N_19603,N_19790);
nor UO_106 (O_106,N_19683,N_19748);
and UO_107 (O_107,N_19511,N_19519);
or UO_108 (O_108,N_19690,N_19732);
and UO_109 (O_109,N_19591,N_19659);
or UO_110 (O_110,N_19988,N_19846);
nor UO_111 (O_111,N_19773,N_19857);
or UO_112 (O_112,N_19704,N_19798);
and UO_113 (O_113,N_19500,N_19810);
nand UO_114 (O_114,N_19760,N_19600);
and UO_115 (O_115,N_19595,N_19919);
and UO_116 (O_116,N_19975,N_19883);
nand UO_117 (O_117,N_19564,N_19868);
and UO_118 (O_118,N_19920,N_19602);
and UO_119 (O_119,N_19554,N_19809);
nor UO_120 (O_120,N_19630,N_19685);
nor UO_121 (O_121,N_19726,N_19657);
nand UO_122 (O_122,N_19528,N_19869);
nor UO_123 (O_123,N_19884,N_19540);
nand UO_124 (O_124,N_19817,N_19913);
and UO_125 (O_125,N_19879,N_19645);
nand UO_126 (O_126,N_19762,N_19830);
nor UO_127 (O_127,N_19819,N_19522);
nor UO_128 (O_128,N_19842,N_19709);
nor UO_129 (O_129,N_19730,N_19935);
nand UO_130 (O_130,N_19694,N_19806);
and UO_131 (O_131,N_19753,N_19755);
nor UO_132 (O_132,N_19814,N_19627);
nand UO_133 (O_133,N_19952,N_19520);
or UO_134 (O_134,N_19958,N_19768);
xor UO_135 (O_135,N_19808,N_19918);
nand UO_136 (O_136,N_19571,N_19807);
or UO_137 (O_137,N_19912,N_19969);
and UO_138 (O_138,N_19558,N_19949);
nand UO_139 (O_139,N_19653,N_19537);
or UO_140 (O_140,N_19815,N_19745);
or UO_141 (O_141,N_19583,N_19961);
and UO_142 (O_142,N_19829,N_19527);
or UO_143 (O_143,N_19982,N_19679);
or UO_144 (O_144,N_19569,N_19544);
or UO_145 (O_145,N_19786,N_19770);
nand UO_146 (O_146,N_19711,N_19898);
and UO_147 (O_147,N_19851,N_19560);
nand UO_148 (O_148,N_19995,N_19972);
xor UO_149 (O_149,N_19534,N_19572);
or UO_150 (O_150,N_19695,N_19908);
nor UO_151 (O_151,N_19670,N_19971);
or UO_152 (O_152,N_19981,N_19833);
or UO_153 (O_153,N_19792,N_19649);
nand UO_154 (O_154,N_19707,N_19650);
nor UO_155 (O_155,N_19720,N_19549);
or UO_156 (O_156,N_19708,N_19628);
and UO_157 (O_157,N_19552,N_19535);
or UO_158 (O_158,N_19546,N_19680);
and UO_159 (O_159,N_19620,N_19503);
nor UO_160 (O_160,N_19734,N_19735);
nand UO_161 (O_161,N_19582,N_19521);
xnor UO_162 (O_162,N_19965,N_19769);
nor UO_163 (O_163,N_19677,N_19844);
xor UO_164 (O_164,N_19634,N_19551);
and UO_165 (O_165,N_19956,N_19937);
and UO_166 (O_166,N_19636,N_19594);
nand UO_167 (O_167,N_19651,N_19823);
nand UO_168 (O_168,N_19876,N_19646);
nand UO_169 (O_169,N_19976,N_19902);
or UO_170 (O_170,N_19678,N_19668);
or UO_171 (O_171,N_19765,N_19849);
nand UO_172 (O_172,N_19835,N_19644);
and UO_173 (O_173,N_19736,N_19774);
and UO_174 (O_174,N_19836,N_19706);
xor UO_175 (O_175,N_19855,N_19828);
or UO_176 (O_176,N_19789,N_19605);
or UO_177 (O_177,N_19691,N_19563);
nand UO_178 (O_178,N_19779,N_19761);
xnor UO_179 (O_179,N_19676,N_19742);
and UO_180 (O_180,N_19803,N_19873);
and UO_181 (O_181,N_19663,N_19526);
and UO_182 (O_182,N_19941,N_19925);
and UO_183 (O_183,N_19966,N_19999);
nor UO_184 (O_184,N_19586,N_19741);
or UO_185 (O_185,N_19581,N_19933);
nand UO_186 (O_186,N_19759,N_19565);
nand UO_187 (O_187,N_19824,N_19675);
nor UO_188 (O_188,N_19945,N_19640);
nand UO_189 (O_189,N_19993,N_19667);
nand UO_190 (O_190,N_19985,N_19737);
or UO_191 (O_191,N_19986,N_19664);
xor UO_192 (O_192,N_19838,N_19987);
and UO_193 (O_193,N_19758,N_19610);
or UO_194 (O_194,N_19778,N_19559);
nand UO_195 (O_195,N_19936,N_19548);
nor UO_196 (O_196,N_19665,N_19953);
and UO_197 (O_197,N_19575,N_19533);
or UO_198 (O_198,N_19875,N_19577);
nor UO_199 (O_199,N_19881,N_19719);
and UO_200 (O_200,N_19509,N_19804);
and UO_201 (O_201,N_19658,N_19523);
and UO_202 (O_202,N_19878,N_19725);
and UO_203 (O_203,N_19989,N_19877);
nand UO_204 (O_204,N_19964,N_19576);
nand UO_205 (O_205,N_19882,N_19652);
or UO_206 (O_206,N_19957,N_19960);
or UO_207 (O_207,N_19578,N_19738);
xor UO_208 (O_208,N_19931,N_19897);
nor UO_209 (O_209,N_19801,N_19747);
or UO_210 (O_210,N_19787,N_19557);
nand UO_211 (O_211,N_19666,N_19632);
nand UO_212 (O_212,N_19669,N_19568);
and UO_213 (O_213,N_19584,N_19612);
nor UO_214 (O_214,N_19926,N_19606);
and UO_215 (O_215,N_19573,N_19750);
and UO_216 (O_216,N_19940,N_19631);
or UO_217 (O_217,N_19781,N_19674);
or UO_218 (O_218,N_19579,N_19766);
nand UO_219 (O_219,N_19862,N_19921);
nor UO_220 (O_220,N_19661,N_19689);
nor UO_221 (O_221,N_19504,N_19927);
and UO_222 (O_222,N_19510,N_19596);
xnor UO_223 (O_223,N_19805,N_19687);
nor UO_224 (O_224,N_19731,N_19545);
or UO_225 (O_225,N_19797,N_19887);
nor UO_226 (O_226,N_19853,N_19531);
nand UO_227 (O_227,N_19585,N_19727);
nor UO_228 (O_228,N_19660,N_19626);
nor UO_229 (O_229,N_19818,N_19752);
and UO_230 (O_230,N_19567,N_19767);
or UO_231 (O_231,N_19712,N_19532);
or UO_232 (O_232,N_19788,N_19543);
nor UO_233 (O_233,N_19800,N_19923);
and UO_234 (O_234,N_19728,N_19672);
or UO_235 (O_235,N_19524,N_19598);
nor UO_236 (O_236,N_19967,N_19710);
and UO_237 (O_237,N_19536,N_19983);
xnor UO_238 (O_238,N_19888,N_19915);
xnor UO_239 (O_239,N_19932,N_19821);
nor UO_240 (O_240,N_19530,N_19715);
or UO_241 (O_241,N_19625,N_19542);
nor UO_242 (O_242,N_19782,N_19839);
nand UO_243 (O_243,N_19507,N_19841);
or UO_244 (O_244,N_19910,N_19998);
and UO_245 (O_245,N_19820,N_19904);
nor UO_246 (O_246,N_19515,N_19955);
nand UO_247 (O_247,N_19700,N_19911);
or UO_248 (O_248,N_19739,N_19837);
or UO_249 (O_249,N_19733,N_19795);
nor UO_250 (O_250,N_19772,N_19564);
or UO_251 (O_251,N_19602,N_19512);
nand UO_252 (O_252,N_19522,N_19942);
or UO_253 (O_253,N_19626,N_19957);
nand UO_254 (O_254,N_19638,N_19510);
or UO_255 (O_255,N_19926,N_19793);
nand UO_256 (O_256,N_19666,N_19979);
or UO_257 (O_257,N_19824,N_19680);
nor UO_258 (O_258,N_19536,N_19728);
nand UO_259 (O_259,N_19967,N_19623);
xor UO_260 (O_260,N_19848,N_19666);
and UO_261 (O_261,N_19766,N_19677);
or UO_262 (O_262,N_19935,N_19714);
and UO_263 (O_263,N_19902,N_19825);
nand UO_264 (O_264,N_19668,N_19584);
nor UO_265 (O_265,N_19917,N_19863);
nand UO_266 (O_266,N_19879,N_19666);
and UO_267 (O_267,N_19684,N_19611);
nand UO_268 (O_268,N_19911,N_19692);
nor UO_269 (O_269,N_19836,N_19885);
nand UO_270 (O_270,N_19947,N_19723);
and UO_271 (O_271,N_19933,N_19741);
or UO_272 (O_272,N_19824,N_19903);
nand UO_273 (O_273,N_19868,N_19996);
and UO_274 (O_274,N_19503,N_19802);
or UO_275 (O_275,N_19679,N_19685);
nand UO_276 (O_276,N_19921,N_19541);
and UO_277 (O_277,N_19953,N_19525);
nand UO_278 (O_278,N_19932,N_19601);
and UO_279 (O_279,N_19715,N_19841);
or UO_280 (O_280,N_19696,N_19836);
nor UO_281 (O_281,N_19661,N_19928);
nand UO_282 (O_282,N_19998,N_19630);
and UO_283 (O_283,N_19826,N_19623);
nor UO_284 (O_284,N_19684,N_19806);
and UO_285 (O_285,N_19972,N_19542);
or UO_286 (O_286,N_19554,N_19962);
and UO_287 (O_287,N_19935,N_19509);
and UO_288 (O_288,N_19932,N_19565);
and UO_289 (O_289,N_19610,N_19547);
and UO_290 (O_290,N_19899,N_19893);
nand UO_291 (O_291,N_19689,N_19586);
and UO_292 (O_292,N_19981,N_19873);
and UO_293 (O_293,N_19954,N_19728);
nand UO_294 (O_294,N_19622,N_19506);
nor UO_295 (O_295,N_19598,N_19753);
nand UO_296 (O_296,N_19876,N_19778);
nor UO_297 (O_297,N_19912,N_19956);
or UO_298 (O_298,N_19584,N_19749);
nand UO_299 (O_299,N_19675,N_19740);
nor UO_300 (O_300,N_19800,N_19687);
nand UO_301 (O_301,N_19758,N_19680);
xnor UO_302 (O_302,N_19938,N_19738);
nor UO_303 (O_303,N_19552,N_19958);
nor UO_304 (O_304,N_19637,N_19922);
or UO_305 (O_305,N_19683,N_19751);
nor UO_306 (O_306,N_19580,N_19687);
nand UO_307 (O_307,N_19791,N_19952);
nor UO_308 (O_308,N_19530,N_19545);
nand UO_309 (O_309,N_19764,N_19527);
nor UO_310 (O_310,N_19533,N_19790);
or UO_311 (O_311,N_19777,N_19602);
nand UO_312 (O_312,N_19526,N_19606);
nor UO_313 (O_313,N_19805,N_19552);
xor UO_314 (O_314,N_19928,N_19604);
nand UO_315 (O_315,N_19568,N_19883);
and UO_316 (O_316,N_19830,N_19533);
or UO_317 (O_317,N_19953,N_19708);
and UO_318 (O_318,N_19923,N_19939);
nor UO_319 (O_319,N_19854,N_19569);
xor UO_320 (O_320,N_19576,N_19567);
or UO_321 (O_321,N_19592,N_19559);
and UO_322 (O_322,N_19942,N_19525);
xor UO_323 (O_323,N_19903,N_19533);
and UO_324 (O_324,N_19951,N_19873);
or UO_325 (O_325,N_19717,N_19597);
and UO_326 (O_326,N_19962,N_19898);
or UO_327 (O_327,N_19947,N_19852);
and UO_328 (O_328,N_19715,N_19979);
nand UO_329 (O_329,N_19907,N_19751);
or UO_330 (O_330,N_19569,N_19923);
nand UO_331 (O_331,N_19512,N_19869);
nor UO_332 (O_332,N_19897,N_19887);
and UO_333 (O_333,N_19706,N_19632);
nand UO_334 (O_334,N_19507,N_19540);
nand UO_335 (O_335,N_19819,N_19623);
nor UO_336 (O_336,N_19796,N_19620);
nor UO_337 (O_337,N_19698,N_19830);
nand UO_338 (O_338,N_19801,N_19933);
nor UO_339 (O_339,N_19726,N_19963);
nand UO_340 (O_340,N_19590,N_19745);
and UO_341 (O_341,N_19604,N_19806);
xnor UO_342 (O_342,N_19934,N_19834);
nor UO_343 (O_343,N_19987,N_19649);
nand UO_344 (O_344,N_19645,N_19630);
nand UO_345 (O_345,N_19778,N_19561);
and UO_346 (O_346,N_19859,N_19992);
nand UO_347 (O_347,N_19504,N_19713);
nor UO_348 (O_348,N_19951,N_19650);
and UO_349 (O_349,N_19705,N_19952);
and UO_350 (O_350,N_19563,N_19693);
nor UO_351 (O_351,N_19964,N_19737);
nor UO_352 (O_352,N_19751,N_19825);
and UO_353 (O_353,N_19821,N_19938);
nor UO_354 (O_354,N_19863,N_19662);
and UO_355 (O_355,N_19834,N_19741);
nor UO_356 (O_356,N_19755,N_19684);
nor UO_357 (O_357,N_19639,N_19991);
and UO_358 (O_358,N_19799,N_19678);
or UO_359 (O_359,N_19750,N_19570);
and UO_360 (O_360,N_19908,N_19939);
xnor UO_361 (O_361,N_19952,N_19649);
nand UO_362 (O_362,N_19844,N_19949);
nand UO_363 (O_363,N_19852,N_19820);
and UO_364 (O_364,N_19570,N_19566);
or UO_365 (O_365,N_19874,N_19907);
nor UO_366 (O_366,N_19900,N_19979);
or UO_367 (O_367,N_19549,N_19979);
or UO_368 (O_368,N_19947,N_19579);
nor UO_369 (O_369,N_19738,N_19544);
nand UO_370 (O_370,N_19812,N_19898);
and UO_371 (O_371,N_19559,N_19606);
nor UO_372 (O_372,N_19954,N_19637);
nor UO_373 (O_373,N_19529,N_19646);
nor UO_374 (O_374,N_19847,N_19755);
nor UO_375 (O_375,N_19980,N_19539);
or UO_376 (O_376,N_19853,N_19867);
nand UO_377 (O_377,N_19540,N_19542);
or UO_378 (O_378,N_19894,N_19529);
and UO_379 (O_379,N_19708,N_19933);
nand UO_380 (O_380,N_19960,N_19667);
nor UO_381 (O_381,N_19606,N_19647);
nand UO_382 (O_382,N_19544,N_19906);
or UO_383 (O_383,N_19830,N_19525);
and UO_384 (O_384,N_19530,N_19597);
or UO_385 (O_385,N_19548,N_19634);
nor UO_386 (O_386,N_19531,N_19638);
or UO_387 (O_387,N_19906,N_19619);
and UO_388 (O_388,N_19695,N_19919);
nor UO_389 (O_389,N_19571,N_19921);
nor UO_390 (O_390,N_19971,N_19826);
nand UO_391 (O_391,N_19550,N_19940);
or UO_392 (O_392,N_19975,N_19520);
and UO_393 (O_393,N_19710,N_19608);
nand UO_394 (O_394,N_19536,N_19542);
and UO_395 (O_395,N_19614,N_19850);
nor UO_396 (O_396,N_19755,N_19903);
nor UO_397 (O_397,N_19633,N_19968);
nor UO_398 (O_398,N_19575,N_19694);
nand UO_399 (O_399,N_19526,N_19514);
nand UO_400 (O_400,N_19833,N_19915);
or UO_401 (O_401,N_19935,N_19995);
and UO_402 (O_402,N_19764,N_19726);
and UO_403 (O_403,N_19812,N_19729);
nand UO_404 (O_404,N_19623,N_19524);
xnor UO_405 (O_405,N_19753,N_19765);
or UO_406 (O_406,N_19924,N_19868);
nand UO_407 (O_407,N_19827,N_19701);
and UO_408 (O_408,N_19874,N_19839);
and UO_409 (O_409,N_19824,N_19548);
nor UO_410 (O_410,N_19886,N_19576);
nor UO_411 (O_411,N_19596,N_19659);
or UO_412 (O_412,N_19653,N_19610);
or UO_413 (O_413,N_19989,N_19632);
nor UO_414 (O_414,N_19581,N_19674);
nand UO_415 (O_415,N_19805,N_19683);
or UO_416 (O_416,N_19550,N_19872);
and UO_417 (O_417,N_19971,N_19891);
and UO_418 (O_418,N_19983,N_19947);
nor UO_419 (O_419,N_19627,N_19976);
and UO_420 (O_420,N_19911,N_19961);
nor UO_421 (O_421,N_19741,N_19663);
nand UO_422 (O_422,N_19990,N_19745);
or UO_423 (O_423,N_19645,N_19853);
or UO_424 (O_424,N_19933,N_19823);
and UO_425 (O_425,N_19725,N_19612);
or UO_426 (O_426,N_19707,N_19649);
or UO_427 (O_427,N_19952,N_19931);
nor UO_428 (O_428,N_19577,N_19979);
nand UO_429 (O_429,N_19753,N_19796);
nand UO_430 (O_430,N_19512,N_19803);
nand UO_431 (O_431,N_19635,N_19846);
and UO_432 (O_432,N_19665,N_19656);
or UO_433 (O_433,N_19704,N_19510);
nor UO_434 (O_434,N_19884,N_19814);
and UO_435 (O_435,N_19945,N_19526);
nor UO_436 (O_436,N_19542,N_19940);
and UO_437 (O_437,N_19875,N_19989);
nor UO_438 (O_438,N_19796,N_19595);
nand UO_439 (O_439,N_19876,N_19589);
and UO_440 (O_440,N_19774,N_19630);
nor UO_441 (O_441,N_19850,N_19519);
or UO_442 (O_442,N_19922,N_19862);
or UO_443 (O_443,N_19945,N_19714);
and UO_444 (O_444,N_19718,N_19705);
or UO_445 (O_445,N_19682,N_19546);
nand UO_446 (O_446,N_19673,N_19869);
and UO_447 (O_447,N_19719,N_19841);
or UO_448 (O_448,N_19744,N_19870);
nor UO_449 (O_449,N_19602,N_19547);
and UO_450 (O_450,N_19984,N_19710);
nor UO_451 (O_451,N_19655,N_19938);
or UO_452 (O_452,N_19562,N_19632);
nand UO_453 (O_453,N_19814,N_19975);
nand UO_454 (O_454,N_19966,N_19845);
xnor UO_455 (O_455,N_19639,N_19546);
nand UO_456 (O_456,N_19969,N_19718);
nand UO_457 (O_457,N_19822,N_19665);
or UO_458 (O_458,N_19777,N_19799);
xnor UO_459 (O_459,N_19899,N_19985);
nor UO_460 (O_460,N_19585,N_19575);
and UO_461 (O_461,N_19917,N_19968);
nand UO_462 (O_462,N_19511,N_19828);
and UO_463 (O_463,N_19680,N_19671);
and UO_464 (O_464,N_19973,N_19700);
or UO_465 (O_465,N_19897,N_19556);
nand UO_466 (O_466,N_19784,N_19761);
and UO_467 (O_467,N_19638,N_19771);
and UO_468 (O_468,N_19508,N_19919);
nand UO_469 (O_469,N_19837,N_19596);
or UO_470 (O_470,N_19637,N_19844);
nand UO_471 (O_471,N_19860,N_19660);
nand UO_472 (O_472,N_19660,N_19901);
nand UO_473 (O_473,N_19891,N_19788);
nor UO_474 (O_474,N_19669,N_19691);
nor UO_475 (O_475,N_19823,N_19799);
nand UO_476 (O_476,N_19750,N_19822);
or UO_477 (O_477,N_19625,N_19786);
and UO_478 (O_478,N_19680,N_19898);
xor UO_479 (O_479,N_19680,N_19779);
or UO_480 (O_480,N_19913,N_19828);
and UO_481 (O_481,N_19780,N_19649);
or UO_482 (O_482,N_19531,N_19741);
nor UO_483 (O_483,N_19707,N_19762);
and UO_484 (O_484,N_19687,N_19873);
nor UO_485 (O_485,N_19977,N_19816);
and UO_486 (O_486,N_19818,N_19521);
nand UO_487 (O_487,N_19731,N_19766);
nor UO_488 (O_488,N_19731,N_19774);
and UO_489 (O_489,N_19501,N_19666);
nand UO_490 (O_490,N_19831,N_19756);
or UO_491 (O_491,N_19939,N_19773);
nor UO_492 (O_492,N_19879,N_19596);
nor UO_493 (O_493,N_19809,N_19517);
nor UO_494 (O_494,N_19504,N_19847);
or UO_495 (O_495,N_19565,N_19968);
and UO_496 (O_496,N_19882,N_19892);
or UO_497 (O_497,N_19560,N_19631);
nand UO_498 (O_498,N_19852,N_19945);
and UO_499 (O_499,N_19922,N_19825);
and UO_500 (O_500,N_19842,N_19658);
nand UO_501 (O_501,N_19997,N_19746);
nor UO_502 (O_502,N_19567,N_19520);
or UO_503 (O_503,N_19860,N_19562);
nand UO_504 (O_504,N_19681,N_19565);
and UO_505 (O_505,N_19755,N_19506);
and UO_506 (O_506,N_19787,N_19912);
and UO_507 (O_507,N_19710,N_19515);
nor UO_508 (O_508,N_19686,N_19757);
nand UO_509 (O_509,N_19572,N_19900);
nand UO_510 (O_510,N_19981,N_19982);
nand UO_511 (O_511,N_19747,N_19768);
and UO_512 (O_512,N_19859,N_19596);
nor UO_513 (O_513,N_19957,N_19783);
and UO_514 (O_514,N_19915,N_19823);
or UO_515 (O_515,N_19912,N_19928);
or UO_516 (O_516,N_19659,N_19655);
nand UO_517 (O_517,N_19659,N_19559);
nor UO_518 (O_518,N_19792,N_19548);
and UO_519 (O_519,N_19588,N_19540);
nor UO_520 (O_520,N_19852,N_19563);
nor UO_521 (O_521,N_19548,N_19810);
or UO_522 (O_522,N_19961,N_19546);
nand UO_523 (O_523,N_19729,N_19761);
nor UO_524 (O_524,N_19597,N_19751);
and UO_525 (O_525,N_19597,N_19653);
nor UO_526 (O_526,N_19741,N_19822);
or UO_527 (O_527,N_19628,N_19959);
and UO_528 (O_528,N_19836,N_19703);
and UO_529 (O_529,N_19916,N_19711);
or UO_530 (O_530,N_19603,N_19914);
and UO_531 (O_531,N_19912,N_19861);
or UO_532 (O_532,N_19929,N_19653);
nand UO_533 (O_533,N_19606,N_19886);
or UO_534 (O_534,N_19789,N_19863);
nand UO_535 (O_535,N_19909,N_19967);
nor UO_536 (O_536,N_19823,N_19789);
or UO_537 (O_537,N_19674,N_19765);
and UO_538 (O_538,N_19536,N_19758);
or UO_539 (O_539,N_19714,N_19810);
and UO_540 (O_540,N_19740,N_19748);
nor UO_541 (O_541,N_19640,N_19775);
nand UO_542 (O_542,N_19825,N_19940);
or UO_543 (O_543,N_19503,N_19968);
xnor UO_544 (O_544,N_19657,N_19975);
or UO_545 (O_545,N_19743,N_19552);
xor UO_546 (O_546,N_19522,N_19516);
and UO_547 (O_547,N_19815,N_19570);
nor UO_548 (O_548,N_19566,N_19627);
or UO_549 (O_549,N_19725,N_19846);
and UO_550 (O_550,N_19756,N_19915);
nand UO_551 (O_551,N_19516,N_19823);
or UO_552 (O_552,N_19879,N_19554);
or UO_553 (O_553,N_19789,N_19709);
or UO_554 (O_554,N_19517,N_19500);
and UO_555 (O_555,N_19566,N_19608);
and UO_556 (O_556,N_19981,N_19928);
and UO_557 (O_557,N_19800,N_19982);
and UO_558 (O_558,N_19787,N_19788);
or UO_559 (O_559,N_19568,N_19512);
and UO_560 (O_560,N_19957,N_19580);
and UO_561 (O_561,N_19514,N_19933);
and UO_562 (O_562,N_19579,N_19719);
nor UO_563 (O_563,N_19863,N_19938);
nand UO_564 (O_564,N_19942,N_19873);
or UO_565 (O_565,N_19519,N_19564);
nand UO_566 (O_566,N_19757,N_19989);
nand UO_567 (O_567,N_19728,N_19840);
nor UO_568 (O_568,N_19895,N_19512);
and UO_569 (O_569,N_19990,N_19536);
nand UO_570 (O_570,N_19981,N_19501);
or UO_571 (O_571,N_19557,N_19976);
and UO_572 (O_572,N_19674,N_19734);
nor UO_573 (O_573,N_19567,N_19952);
xor UO_574 (O_574,N_19541,N_19548);
nand UO_575 (O_575,N_19946,N_19904);
nor UO_576 (O_576,N_19762,N_19938);
nor UO_577 (O_577,N_19892,N_19995);
or UO_578 (O_578,N_19554,N_19595);
and UO_579 (O_579,N_19725,N_19890);
nand UO_580 (O_580,N_19915,N_19879);
nor UO_581 (O_581,N_19696,N_19782);
nand UO_582 (O_582,N_19577,N_19786);
nand UO_583 (O_583,N_19787,N_19774);
or UO_584 (O_584,N_19524,N_19796);
and UO_585 (O_585,N_19506,N_19503);
nor UO_586 (O_586,N_19757,N_19600);
or UO_587 (O_587,N_19988,N_19811);
nand UO_588 (O_588,N_19824,N_19816);
or UO_589 (O_589,N_19847,N_19731);
nor UO_590 (O_590,N_19617,N_19926);
or UO_591 (O_591,N_19746,N_19778);
and UO_592 (O_592,N_19926,N_19801);
nand UO_593 (O_593,N_19908,N_19768);
nor UO_594 (O_594,N_19689,N_19935);
or UO_595 (O_595,N_19633,N_19945);
or UO_596 (O_596,N_19802,N_19979);
or UO_597 (O_597,N_19832,N_19504);
nand UO_598 (O_598,N_19706,N_19788);
and UO_599 (O_599,N_19805,N_19958);
and UO_600 (O_600,N_19501,N_19772);
nor UO_601 (O_601,N_19683,N_19564);
nor UO_602 (O_602,N_19713,N_19540);
nor UO_603 (O_603,N_19796,N_19818);
or UO_604 (O_604,N_19580,N_19572);
nand UO_605 (O_605,N_19726,N_19584);
and UO_606 (O_606,N_19826,N_19957);
nand UO_607 (O_607,N_19828,N_19518);
and UO_608 (O_608,N_19829,N_19656);
nand UO_609 (O_609,N_19964,N_19717);
or UO_610 (O_610,N_19652,N_19862);
nor UO_611 (O_611,N_19558,N_19856);
or UO_612 (O_612,N_19746,N_19675);
or UO_613 (O_613,N_19794,N_19762);
or UO_614 (O_614,N_19526,N_19641);
nor UO_615 (O_615,N_19766,N_19581);
nor UO_616 (O_616,N_19585,N_19704);
nor UO_617 (O_617,N_19861,N_19820);
nor UO_618 (O_618,N_19893,N_19933);
nand UO_619 (O_619,N_19781,N_19714);
and UO_620 (O_620,N_19715,N_19591);
or UO_621 (O_621,N_19603,N_19986);
nor UO_622 (O_622,N_19919,N_19523);
and UO_623 (O_623,N_19695,N_19859);
nand UO_624 (O_624,N_19829,N_19726);
nor UO_625 (O_625,N_19649,N_19943);
and UO_626 (O_626,N_19524,N_19894);
and UO_627 (O_627,N_19848,N_19834);
and UO_628 (O_628,N_19808,N_19527);
and UO_629 (O_629,N_19599,N_19686);
or UO_630 (O_630,N_19804,N_19610);
nor UO_631 (O_631,N_19832,N_19903);
and UO_632 (O_632,N_19982,N_19925);
nor UO_633 (O_633,N_19638,N_19950);
nand UO_634 (O_634,N_19764,N_19746);
nand UO_635 (O_635,N_19763,N_19890);
nand UO_636 (O_636,N_19799,N_19934);
nor UO_637 (O_637,N_19519,N_19640);
nor UO_638 (O_638,N_19545,N_19529);
nand UO_639 (O_639,N_19555,N_19681);
or UO_640 (O_640,N_19776,N_19886);
and UO_641 (O_641,N_19656,N_19977);
or UO_642 (O_642,N_19521,N_19762);
xor UO_643 (O_643,N_19596,N_19720);
nand UO_644 (O_644,N_19898,N_19629);
and UO_645 (O_645,N_19831,N_19513);
nor UO_646 (O_646,N_19587,N_19591);
nand UO_647 (O_647,N_19789,N_19775);
or UO_648 (O_648,N_19663,N_19714);
and UO_649 (O_649,N_19938,N_19884);
nor UO_650 (O_650,N_19607,N_19626);
nand UO_651 (O_651,N_19679,N_19594);
or UO_652 (O_652,N_19701,N_19587);
or UO_653 (O_653,N_19978,N_19820);
nor UO_654 (O_654,N_19965,N_19960);
and UO_655 (O_655,N_19636,N_19938);
or UO_656 (O_656,N_19626,N_19721);
nor UO_657 (O_657,N_19916,N_19700);
or UO_658 (O_658,N_19761,N_19792);
nor UO_659 (O_659,N_19568,N_19640);
nand UO_660 (O_660,N_19559,N_19527);
and UO_661 (O_661,N_19612,N_19916);
nor UO_662 (O_662,N_19595,N_19680);
nand UO_663 (O_663,N_19839,N_19877);
nor UO_664 (O_664,N_19940,N_19570);
nor UO_665 (O_665,N_19979,N_19967);
or UO_666 (O_666,N_19851,N_19695);
and UO_667 (O_667,N_19688,N_19657);
or UO_668 (O_668,N_19574,N_19985);
and UO_669 (O_669,N_19996,N_19912);
nor UO_670 (O_670,N_19617,N_19821);
and UO_671 (O_671,N_19983,N_19750);
and UO_672 (O_672,N_19820,N_19897);
nor UO_673 (O_673,N_19777,N_19547);
and UO_674 (O_674,N_19602,N_19557);
and UO_675 (O_675,N_19995,N_19628);
and UO_676 (O_676,N_19710,N_19712);
nand UO_677 (O_677,N_19954,N_19981);
and UO_678 (O_678,N_19999,N_19594);
and UO_679 (O_679,N_19658,N_19818);
nor UO_680 (O_680,N_19561,N_19570);
or UO_681 (O_681,N_19788,N_19911);
nor UO_682 (O_682,N_19941,N_19691);
or UO_683 (O_683,N_19527,N_19637);
xor UO_684 (O_684,N_19847,N_19958);
and UO_685 (O_685,N_19681,N_19582);
or UO_686 (O_686,N_19632,N_19766);
nor UO_687 (O_687,N_19940,N_19607);
and UO_688 (O_688,N_19551,N_19754);
nand UO_689 (O_689,N_19616,N_19729);
or UO_690 (O_690,N_19617,N_19827);
and UO_691 (O_691,N_19891,N_19929);
nor UO_692 (O_692,N_19630,N_19657);
xor UO_693 (O_693,N_19526,N_19965);
or UO_694 (O_694,N_19769,N_19704);
nor UO_695 (O_695,N_19807,N_19912);
nor UO_696 (O_696,N_19632,N_19759);
xor UO_697 (O_697,N_19765,N_19549);
nor UO_698 (O_698,N_19505,N_19678);
or UO_699 (O_699,N_19552,N_19636);
nor UO_700 (O_700,N_19790,N_19853);
and UO_701 (O_701,N_19558,N_19672);
nor UO_702 (O_702,N_19613,N_19527);
or UO_703 (O_703,N_19552,N_19952);
and UO_704 (O_704,N_19953,N_19673);
xor UO_705 (O_705,N_19917,N_19537);
and UO_706 (O_706,N_19871,N_19544);
nand UO_707 (O_707,N_19977,N_19883);
and UO_708 (O_708,N_19860,N_19930);
nor UO_709 (O_709,N_19531,N_19547);
nor UO_710 (O_710,N_19948,N_19754);
nor UO_711 (O_711,N_19775,N_19559);
or UO_712 (O_712,N_19769,N_19602);
nand UO_713 (O_713,N_19605,N_19816);
nor UO_714 (O_714,N_19949,N_19976);
and UO_715 (O_715,N_19559,N_19647);
nor UO_716 (O_716,N_19696,N_19881);
and UO_717 (O_717,N_19822,N_19748);
nand UO_718 (O_718,N_19824,N_19562);
or UO_719 (O_719,N_19585,N_19741);
nor UO_720 (O_720,N_19697,N_19954);
or UO_721 (O_721,N_19717,N_19543);
and UO_722 (O_722,N_19828,N_19836);
or UO_723 (O_723,N_19773,N_19836);
and UO_724 (O_724,N_19741,N_19562);
nor UO_725 (O_725,N_19998,N_19604);
nand UO_726 (O_726,N_19802,N_19985);
nor UO_727 (O_727,N_19541,N_19502);
or UO_728 (O_728,N_19769,N_19584);
xnor UO_729 (O_729,N_19681,N_19830);
xor UO_730 (O_730,N_19924,N_19947);
nand UO_731 (O_731,N_19586,N_19884);
and UO_732 (O_732,N_19607,N_19790);
and UO_733 (O_733,N_19605,N_19841);
nand UO_734 (O_734,N_19770,N_19613);
and UO_735 (O_735,N_19789,N_19803);
nor UO_736 (O_736,N_19841,N_19877);
or UO_737 (O_737,N_19976,N_19789);
and UO_738 (O_738,N_19863,N_19808);
nand UO_739 (O_739,N_19825,N_19719);
nand UO_740 (O_740,N_19656,N_19585);
and UO_741 (O_741,N_19612,N_19852);
nor UO_742 (O_742,N_19654,N_19898);
nor UO_743 (O_743,N_19628,N_19666);
nor UO_744 (O_744,N_19583,N_19824);
nor UO_745 (O_745,N_19797,N_19697);
and UO_746 (O_746,N_19588,N_19520);
or UO_747 (O_747,N_19690,N_19586);
and UO_748 (O_748,N_19766,N_19712);
or UO_749 (O_749,N_19964,N_19726);
nor UO_750 (O_750,N_19829,N_19588);
and UO_751 (O_751,N_19801,N_19699);
and UO_752 (O_752,N_19920,N_19716);
or UO_753 (O_753,N_19665,N_19940);
nor UO_754 (O_754,N_19987,N_19643);
and UO_755 (O_755,N_19884,N_19598);
or UO_756 (O_756,N_19767,N_19912);
and UO_757 (O_757,N_19747,N_19787);
or UO_758 (O_758,N_19843,N_19979);
nor UO_759 (O_759,N_19538,N_19742);
and UO_760 (O_760,N_19530,N_19510);
nand UO_761 (O_761,N_19542,N_19617);
nor UO_762 (O_762,N_19997,N_19844);
nand UO_763 (O_763,N_19687,N_19725);
or UO_764 (O_764,N_19736,N_19808);
or UO_765 (O_765,N_19899,N_19644);
or UO_766 (O_766,N_19556,N_19680);
and UO_767 (O_767,N_19796,N_19660);
and UO_768 (O_768,N_19903,N_19914);
and UO_769 (O_769,N_19675,N_19932);
nor UO_770 (O_770,N_19906,N_19798);
nand UO_771 (O_771,N_19942,N_19841);
nor UO_772 (O_772,N_19679,N_19859);
nor UO_773 (O_773,N_19776,N_19562);
or UO_774 (O_774,N_19807,N_19515);
nor UO_775 (O_775,N_19901,N_19504);
and UO_776 (O_776,N_19706,N_19738);
or UO_777 (O_777,N_19962,N_19968);
nor UO_778 (O_778,N_19886,N_19814);
nand UO_779 (O_779,N_19912,N_19575);
and UO_780 (O_780,N_19515,N_19759);
nor UO_781 (O_781,N_19804,N_19563);
and UO_782 (O_782,N_19528,N_19755);
or UO_783 (O_783,N_19859,N_19670);
or UO_784 (O_784,N_19955,N_19690);
and UO_785 (O_785,N_19725,N_19801);
or UO_786 (O_786,N_19978,N_19935);
and UO_787 (O_787,N_19683,N_19980);
and UO_788 (O_788,N_19775,N_19694);
nor UO_789 (O_789,N_19545,N_19926);
or UO_790 (O_790,N_19551,N_19772);
or UO_791 (O_791,N_19744,N_19660);
and UO_792 (O_792,N_19889,N_19723);
nand UO_793 (O_793,N_19611,N_19931);
or UO_794 (O_794,N_19689,N_19745);
and UO_795 (O_795,N_19983,N_19538);
nor UO_796 (O_796,N_19774,N_19530);
nand UO_797 (O_797,N_19521,N_19831);
nand UO_798 (O_798,N_19503,N_19500);
nand UO_799 (O_799,N_19742,N_19985);
or UO_800 (O_800,N_19701,N_19765);
or UO_801 (O_801,N_19996,N_19674);
and UO_802 (O_802,N_19579,N_19715);
nand UO_803 (O_803,N_19536,N_19809);
and UO_804 (O_804,N_19640,N_19621);
and UO_805 (O_805,N_19659,N_19755);
nor UO_806 (O_806,N_19551,N_19796);
nor UO_807 (O_807,N_19747,N_19837);
nor UO_808 (O_808,N_19842,N_19666);
nor UO_809 (O_809,N_19821,N_19520);
or UO_810 (O_810,N_19846,N_19995);
nand UO_811 (O_811,N_19962,N_19974);
and UO_812 (O_812,N_19614,N_19567);
nand UO_813 (O_813,N_19899,N_19733);
or UO_814 (O_814,N_19656,N_19948);
nand UO_815 (O_815,N_19789,N_19752);
nor UO_816 (O_816,N_19502,N_19832);
or UO_817 (O_817,N_19917,N_19628);
or UO_818 (O_818,N_19581,N_19709);
and UO_819 (O_819,N_19919,N_19806);
nor UO_820 (O_820,N_19717,N_19524);
and UO_821 (O_821,N_19656,N_19854);
nor UO_822 (O_822,N_19646,N_19739);
and UO_823 (O_823,N_19889,N_19942);
or UO_824 (O_824,N_19692,N_19981);
nand UO_825 (O_825,N_19919,N_19933);
nor UO_826 (O_826,N_19536,N_19997);
or UO_827 (O_827,N_19968,N_19545);
xnor UO_828 (O_828,N_19579,N_19904);
and UO_829 (O_829,N_19965,N_19843);
xor UO_830 (O_830,N_19552,N_19629);
nor UO_831 (O_831,N_19808,N_19575);
and UO_832 (O_832,N_19652,N_19784);
nand UO_833 (O_833,N_19735,N_19966);
nor UO_834 (O_834,N_19799,N_19776);
nand UO_835 (O_835,N_19984,N_19759);
or UO_836 (O_836,N_19574,N_19821);
nand UO_837 (O_837,N_19594,N_19670);
and UO_838 (O_838,N_19594,N_19567);
or UO_839 (O_839,N_19936,N_19772);
nand UO_840 (O_840,N_19895,N_19760);
nor UO_841 (O_841,N_19966,N_19791);
or UO_842 (O_842,N_19851,N_19691);
nand UO_843 (O_843,N_19591,N_19530);
and UO_844 (O_844,N_19615,N_19573);
or UO_845 (O_845,N_19775,N_19704);
nor UO_846 (O_846,N_19976,N_19568);
or UO_847 (O_847,N_19973,N_19753);
or UO_848 (O_848,N_19930,N_19609);
nand UO_849 (O_849,N_19874,N_19984);
nand UO_850 (O_850,N_19739,N_19604);
nand UO_851 (O_851,N_19779,N_19772);
nor UO_852 (O_852,N_19774,N_19975);
nand UO_853 (O_853,N_19810,N_19583);
nor UO_854 (O_854,N_19824,N_19651);
nand UO_855 (O_855,N_19997,N_19709);
nand UO_856 (O_856,N_19650,N_19968);
and UO_857 (O_857,N_19599,N_19921);
and UO_858 (O_858,N_19922,N_19872);
nor UO_859 (O_859,N_19956,N_19644);
and UO_860 (O_860,N_19734,N_19740);
nor UO_861 (O_861,N_19851,N_19936);
and UO_862 (O_862,N_19896,N_19637);
and UO_863 (O_863,N_19779,N_19809);
and UO_864 (O_864,N_19508,N_19720);
or UO_865 (O_865,N_19729,N_19588);
and UO_866 (O_866,N_19891,N_19855);
nand UO_867 (O_867,N_19881,N_19792);
and UO_868 (O_868,N_19597,N_19845);
nor UO_869 (O_869,N_19760,N_19823);
and UO_870 (O_870,N_19513,N_19508);
nor UO_871 (O_871,N_19712,N_19861);
and UO_872 (O_872,N_19856,N_19738);
nor UO_873 (O_873,N_19598,N_19967);
and UO_874 (O_874,N_19660,N_19580);
and UO_875 (O_875,N_19578,N_19789);
nand UO_876 (O_876,N_19941,N_19743);
nor UO_877 (O_877,N_19563,N_19529);
nand UO_878 (O_878,N_19971,N_19866);
xnor UO_879 (O_879,N_19927,N_19881);
and UO_880 (O_880,N_19561,N_19584);
nor UO_881 (O_881,N_19777,N_19529);
and UO_882 (O_882,N_19791,N_19638);
or UO_883 (O_883,N_19560,N_19546);
xnor UO_884 (O_884,N_19585,N_19696);
nor UO_885 (O_885,N_19538,N_19680);
nor UO_886 (O_886,N_19850,N_19597);
or UO_887 (O_887,N_19924,N_19563);
or UO_888 (O_888,N_19957,N_19675);
nand UO_889 (O_889,N_19989,N_19839);
nor UO_890 (O_890,N_19870,N_19547);
or UO_891 (O_891,N_19738,N_19838);
nor UO_892 (O_892,N_19544,N_19941);
nor UO_893 (O_893,N_19772,N_19828);
or UO_894 (O_894,N_19573,N_19842);
or UO_895 (O_895,N_19885,N_19893);
nor UO_896 (O_896,N_19882,N_19733);
and UO_897 (O_897,N_19651,N_19842);
nor UO_898 (O_898,N_19934,N_19782);
nand UO_899 (O_899,N_19848,N_19656);
or UO_900 (O_900,N_19964,N_19612);
and UO_901 (O_901,N_19986,N_19793);
and UO_902 (O_902,N_19901,N_19973);
and UO_903 (O_903,N_19676,N_19723);
nor UO_904 (O_904,N_19876,N_19889);
or UO_905 (O_905,N_19679,N_19769);
and UO_906 (O_906,N_19506,N_19961);
or UO_907 (O_907,N_19864,N_19714);
and UO_908 (O_908,N_19800,N_19673);
nor UO_909 (O_909,N_19954,N_19861);
or UO_910 (O_910,N_19788,N_19728);
or UO_911 (O_911,N_19574,N_19911);
nor UO_912 (O_912,N_19869,N_19833);
nor UO_913 (O_913,N_19506,N_19627);
and UO_914 (O_914,N_19846,N_19897);
and UO_915 (O_915,N_19769,N_19609);
nand UO_916 (O_916,N_19905,N_19748);
and UO_917 (O_917,N_19823,N_19582);
nand UO_918 (O_918,N_19601,N_19962);
or UO_919 (O_919,N_19638,N_19590);
or UO_920 (O_920,N_19827,N_19680);
nor UO_921 (O_921,N_19710,N_19973);
and UO_922 (O_922,N_19900,N_19739);
and UO_923 (O_923,N_19757,N_19715);
or UO_924 (O_924,N_19999,N_19770);
and UO_925 (O_925,N_19554,N_19642);
nand UO_926 (O_926,N_19812,N_19928);
nor UO_927 (O_927,N_19823,N_19695);
and UO_928 (O_928,N_19833,N_19762);
or UO_929 (O_929,N_19894,N_19719);
nor UO_930 (O_930,N_19912,N_19825);
and UO_931 (O_931,N_19922,N_19881);
and UO_932 (O_932,N_19999,N_19983);
and UO_933 (O_933,N_19533,N_19922);
nor UO_934 (O_934,N_19565,N_19807);
nand UO_935 (O_935,N_19724,N_19929);
nand UO_936 (O_936,N_19719,N_19563);
or UO_937 (O_937,N_19870,N_19703);
nand UO_938 (O_938,N_19695,N_19868);
nand UO_939 (O_939,N_19540,N_19876);
nand UO_940 (O_940,N_19580,N_19822);
and UO_941 (O_941,N_19920,N_19916);
and UO_942 (O_942,N_19887,N_19821);
or UO_943 (O_943,N_19995,N_19852);
nand UO_944 (O_944,N_19808,N_19699);
nand UO_945 (O_945,N_19789,N_19822);
nand UO_946 (O_946,N_19674,N_19846);
and UO_947 (O_947,N_19883,N_19705);
or UO_948 (O_948,N_19771,N_19968);
nand UO_949 (O_949,N_19828,N_19834);
nor UO_950 (O_950,N_19770,N_19926);
nand UO_951 (O_951,N_19830,N_19678);
nor UO_952 (O_952,N_19795,N_19975);
nand UO_953 (O_953,N_19777,N_19790);
and UO_954 (O_954,N_19577,N_19522);
nor UO_955 (O_955,N_19506,N_19948);
or UO_956 (O_956,N_19955,N_19708);
nor UO_957 (O_957,N_19893,N_19628);
nand UO_958 (O_958,N_19659,N_19704);
nand UO_959 (O_959,N_19898,N_19892);
or UO_960 (O_960,N_19677,N_19957);
nor UO_961 (O_961,N_19825,N_19859);
nand UO_962 (O_962,N_19512,N_19916);
and UO_963 (O_963,N_19547,N_19657);
nor UO_964 (O_964,N_19895,N_19972);
nor UO_965 (O_965,N_19856,N_19596);
or UO_966 (O_966,N_19854,N_19761);
and UO_967 (O_967,N_19946,N_19659);
nor UO_968 (O_968,N_19939,N_19643);
or UO_969 (O_969,N_19688,N_19993);
nor UO_970 (O_970,N_19803,N_19882);
nand UO_971 (O_971,N_19884,N_19898);
and UO_972 (O_972,N_19841,N_19943);
nor UO_973 (O_973,N_19854,N_19927);
and UO_974 (O_974,N_19884,N_19575);
xor UO_975 (O_975,N_19637,N_19721);
or UO_976 (O_976,N_19597,N_19747);
nor UO_977 (O_977,N_19824,N_19764);
and UO_978 (O_978,N_19916,N_19701);
nor UO_979 (O_979,N_19733,N_19574);
nor UO_980 (O_980,N_19819,N_19593);
nor UO_981 (O_981,N_19993,N_19672);
nand UO_982 (O_982,N_19775,N_19837);
and UO_983 (O_983,N_19833,N_19755);
nor UO_984 (O_984,N_19510,N_19968);
and UO_985 (O_985,N_19982,N_19683);
or UO_986 (O_986,N_19669,N_19500);
nor UO_987 (O_987,N_19683,N_19566);
nand UO_988 (O_988,N_19965,N_19785);
or UO_989 (O_989,N_19816,N_19802);
and UO_990 (O_990,N_19902,N_19621);
and UO_991 (O_991,N_19646,N_19981);
nand UO_992 (O_992,N_19873,N_19565);
and UO_993 (O_993,N_19801,N_19715);
or UO_994 (O_994,N_19777,N_19862);
or UO_995 (O_995,N_19662,N_19697);
and UO_996 (O_996,N_19639,N_19597);
nand UO_997 (O_997,N_19544,N_19534);
nor UO_998 (O_998,N_19931,N_19898);
nor UO_999 (O_999,N_19975,N_19876);
nor UO_1000 (O_1000,N_19831,N_19520);
nor UO_1001 (O_1001,N_19591,N_19674);
nor UO_1002 (O_1002,N_19517,N_19685);
or UO_1003 (O_1003,N_19967,N_19841);
and UO_1004 (O_1004,N_19754,N_19621);
nor UO_1005 (O_1005,N_19866,N_19753);
or UO_1006 (O_1006,N_19555,N_19724);
or UO_1007 (O_1007,N_19988,N_19771);
or UO_1008 (O_1008,N_19968,N_19774);
nand UO_1009 (O_1009,N_19752,N_19902);
or UO_1010 (O_1010,N_19991,N_19690);
nor UO_1011 (O_1011,N_19640,N_19869);
nor UO_1012 (O_1012,N_19857,N_19658);
and UO_1013 (O_1013,N_19724,N_19813);
or UO_1014 (O_1014,N_19581,N_19819);
and UO_1015 (O_1015,N_19997,N_19503);
and UO_1016 (O_1016,N_19569,N_19582);
nor UO_1017 (O_1017,N_19692,N_19536);
nor UO_1018 (O_1018,N_19529,N_19531);
and UO_1019 (O_1019,N_19883,N_19687);
and UO_1020 (O_1020,N_19884,N_19700);
or UO_1021 (O_1021,N_19735,N_19881);
nor UO_1022 (O_1022,N_19574,N_19503);
or UO_1023 (O_1023,N_19851,N_19584);
nor UO_1024 (O_1024,N_19805,N_19888);
and UO_1025 (O_1025,N_19754,N_19763);
nand UO_1026 (O_1026,N_19518,N_19824);
and UO_1027 (O_1027,N_19829,N_19585);
nand UO_1028 (O_1028,N_19956,N_19833);
and UO_1029 (O_1029,N_19951,N_19607);
nor UO_1030 (O_1030,N_19952,N_19773);
nand UO_1031 (O_1031,N_19518,N_19601);
or UO_1032 (O_1032,N_19979,N_19957);
or UO_1033 (O_1033,N_19976,N_19706);
or UO_1034 (O_1034,N_19964,N_19972);
nand UO_1035 (O_1035,N_19508,N_19806);
and UO_1036 (O_1036,N_19876,N_19515);
nand UO_1037 (O_1037,N_19907,N_19880);
nand UO_1038 (O_1038,N_19926,N_19737);
and UO_1039 (O_1039,N_19883,N_19727);
nand UO_1040 (O_1040,N_19660,N_19715);
nor UO_1041 (O_1041,N_19515,N_19869);
or UO_1042 (O_1042,N_19826,N_19653);
and UO_1043 (O_1043,N_19801,N_19681);
nor UO_1044 (O_1044,N_19973,N_19906);
nor UO_1045 (O_1045,N_19940,N_19686);
nand UO_1046 (O_1046,N_19743,N_19964);
nor UO_1047 (O_1047,N_19876,N_19967);
nor UO_1048 (O_1048,N_19589,N_19705);
nand UO_1049 (O_1049,N_19935,N_19613);
or UO_1050 (O_1050,N_19618,N_19837);
nor UO_1051 (O_1051,N_19779,N_19667);
nor UO_1052 (O_1052,N_19791,N_19698);
and UO_1053 (O_1053,N_19865,N_19711);
nand UO_1054 (O_1054,N_19619,N_19564);
nand UO_1055 (O_1055,N_19523,N_19604);
nor UO_1056 (O_1056,N_19727,N_19862);
nand UO_1057 (O_1057,N_19732,N_19500);
or UO_1058 (O_1058,N_19912,N_19508);
or UO_1059 (O_1059,N_19556,N_19699);
nor UO_1060 (O_1060,N_19709,N_19795);
nor UO_1061 (O_1061,N_19740,N_19602);
nand UO_1062 (O_1062,N_19577,N_19782);
or UO_1063 (O_1063,N_19858,N_19797);
nand UO_1064 (O_1064,N_19805,N_19657);
or UO_1065 (O_1065,N_19562,N_19680);
nor UO_1066 (O_1066,N_19857,N_19516);
or UO_1067 (O_1067,N_19684,N_19717);
nor UO_1068 (O_1068,N_19799,N_19752);
or UO_1069 (O_1069,N_19503,N_19704);
nor UO_1070 (O_1070,N_19567,N_19812);
or UO_1071 (O_1071,N_19899,N_19826);
and UO_1072 (O_1072,N_19662,N_19559);
nor UO_1073 (O_1073,N_19747,N_19765);
nand UO_1074 (O_1074,N_19503,N_19544);
and UO_1075 (O_1075,N_19712,N_19827);
and UO_1076 (O_1076,N_19530,N_19979);
or UO_1077 (O_1077,N_19886,N_19678);
and UO_1078 (O_1078,N_19688,N_19682);
nand UO_1079 (O_1079,N_19959,N_19629);
or UO_1080 (O_1080,N_19504,N_19700);
nor UO_1081 (O_1081,N_19764,N_19725);
and UO_1082 (O_1082,N_19913,N_19689);
or UO_1083 (O_1083,N_19884,N_19773);
xnor UO_1084 (O_1084,N_19844,N_19720);
nor UO_1085 (O_1085,N_19707,N_19798);
nand UO_1086 (O_1086,N_19501,N_19558);
xnor UO_1087 (O_1087,N_19575,N_19609);
nand UO_1088 (O_1088,N_19535,N_19728);
nor UO_1089 (O_1089,N_19921,N_19735);
nand UO_1090 (O_1090,N_19879,N_19836);
nor UO_1091 (O_1091,N_19932,N_19580);
or UO_1092 (O_1092,N_19647,N_19683);
nor UO_1093 (O_1093,N_19893,N_19956);
and UO_1094 (O_1094,N_19875,N_19817);
or UO_1095 (O_1095,N_19907,N_19730);
nand UO_1096 (O_1096,N_19872,N_19501);
or UO_1097 (O_1097,N_19973,N_19957);
or UO_1098 (O_1098,N_19688,N_19897);
nand UO_1099 (O_1099,N_19557,N_19705);
nor UO_1100 (O_1100,N_19502,N_19814);
nor UO_1101 (O_1101,N_19815,N_19883);
nand UO_1102 (O_1102,N_19880,N_19651);
nand UO_1103 (O_1103,N_19744,N_19673);
and UO_1104 (O_1104,N_19891,N_19529);
or UO_1105 (O_1105,N_19847,N_19951);
and UO_1106 (O_1106,N_19834,N_19761);
nand UO_1107 (O_1107,N_19745,N_19750);
and UO_1108 (O_1108,N_19683,N_19550);
or UO_1109 (O_1109,N_19810,N_19599);
and UO_1110 (O_1110,N_19732,N_19982);
nor UO_1111 (O_1111,N_19702,N_19632);
nand UO_1112 (O_1112,N_19968,N_19880);
nand UO_1113 (O_1113,N_19918,N_19805);
nand UO_1114 (O_1114,N_19915,N_19789);
nand UO_1115 (O_1115,N_19646,N_19806);
nand UO_1116 (O_1116,N_19842,N_19670);
nand UO_1117 (O_1117,N_19743,N_19982);
nor UO_1118 (O_1118,N_19819,N_19747);
and UO_1119 (O_1119,N_19933,N_19529);
nor UO_1120 (O_1120,N_19562,N_19629);
and UO_1121 (O_1121,N_19830,N_19548);
nor UO_1122 (O_1122,N_19618,N_19883);
nand UO_1123 (O_1123,N_19931,N_19536);
or UO_1124 (O_1124,N_19984,N_19689);
nor UO_1125 (O_1125,N_19723,N_19561);
or UO_1126 (O_1126,N_19560,N_19777);
nand UO_1127 (O_1127,N_19978,N_19642);
and UO_1128 (O_1128,N_19972,N_19851);
nand UO_1129 (O_1129,N_19636,N_19695);
or UO_1130 (O_1130,N_19779,N_19688);
or UO_1131 (O_1131,N_19753,N_19891);
or UO_1132 (O_1132,N_19899,N_19825);
nand UO_1133 (O_1133,N_19995,N_19933);
nand UO_1134 (O_1134,N_19939,N_19835);
nand UO_1135 (O_1135,N_19673,N_19735);
or UO_1136 (O_1136,N_19842,N_19777);
and UO_1137 (O_1137,N_19939,N_19678);
nor UO_1138 (O_1138,N_19614,N_19631);
or UO_1139 (O_1139,N_19816,N_19587);
and UO_1140 (O_1140,N_19973,N_19920);
or UO_1141 (O_1141,N_19881,N_19716);
or UO_1142 (O_1142,N_19818,N_19975);
or UO_1143 (O_1143,N_19558,N_19981);
or UO_1144 (O_1144,N_19519,N_19744);
nand UO_1145 (O_1145,N_19970,N_19819);
or UO_1146 (O_1146,N_19991,N_19751);
nand UO_1147 (O_1147,N_19827,N_19509);
or UO_1148 (O_1148,N_19859,N_19671);
nand UO_1149 (O_1149,N_19767,N_19710);
and UO_1150 (O_1150,N_19559,N_19740);
nand UO_1151 (O_1151,N_19619,N_19929);
or UO_1152 (O_1152,N_19989,N_19893);
or UO_1153 (O_1153,N_19671,N_19635);
or UO_1154 (O_1154,N_19901,N_19802);
or UO_1155 (O_1155,N_19979,N_19554);
nand UO_1156 (O_1156,N_19979,N_19573);
or UO_1157 (O_1157,N_19962,N_19578);
and UO_1158 (O_1158,N_19614,N_19714);
nand UO_1159 (O_1159,N_19781,N_19872);
or UO_1160 (O_1160,N_19891,N_19942);
nand UO_1161 (O_1161,N_19877,N_19649);
xor UO_1162 (O_1162,N_19705,N_19620);
nor UO_1163 (O_1163,N_19737,N_19873);
nand UO_1164 (O_1164,N_19565,N_19732);
nand UO_1165 (O_1165,N_19547,N_19609);
nor UO_1166 (O_1166,N_19882,N_19678);
xor UO_1167 (O_1167,N_19889,N_19531);
nand UO_1168 (O_1168,N_19994,N_19930);
or UO_1169 (O_1169,N_19619,N_19624);
or UO_1170 (O_1170,N_19626,N_19511);
nor UO_1171 (O_1171,N_19548,N_19646);
nor UO_1172 (O_1172,N_19859,N_19974);
and UO_1173 (O_1173,N_19916,N_19934);
xnor UO_1174 (O_1174,N_19645,N_19519);
nand UO_1175 (O_1175,N_19990,N_19981);
nand UO_1176 (O_1176,N_19788,N_19954);
or UO_1177 (O_1177,N_19618,N_19535);
nand UO_1178 (O_1178,N_19736,N_19922);
and UO_1179 (O_1179,N_19886,N_19515);
nor UO_1180 (O_1180,N_19979,N_19570);
nand UO_1181 (O_1181,N_19882,N_19671);
nand UO_1182 (O_1182,N_19551,N_19871);
and UO_1183 (O_1183,N_19539,N_19706);
or UO_1184 (O_1184,N_19753,N_19636);
nor UO_1185 (O_1185,N_19707,N_19621);
nand UO_1186 (O_1186,N_19673,N_19698);
and UO_1187 (O_1187,N_19823,N_19810);
and UO_1188 (O_1188,N_19941,N_19662);
and UO_1189 (O_1189,N_19933,N_19588);
or UO_1190 (O_1190,N_19926,N_19815);
nor UO_1191 (O_1191,N_19655,N_19981);
nand UO_1192 (O_1192,N_19714,N_19822);
nand UO_1193 (O_1193,N_19914,N_19977);
nor UO_1194 (O_1194,N_19639,N_19728);
nand UO_1195 (O_1195,N_19560,N_19604);
or UO_1196 (O_1196,N_19736,N_19951);
and UO_1197 (O_1197,N_19508,N_19692);
and UO_1198 (O_1198,N_19846,N_19780);
and UO_1199 (O_1199,N_19500,N_19882);
nand UO_1200 (O_1200,N_19510,N_19691);
or UO_1201 (O_1201,N_19619,N_19743);
or UO_1202 (O_1202,N_19752,N_19530);
and UO_1203 (O_1203,N_19631,N_19622);
or UO_1204 (O_1204,N_19545,N_19549);
nand UO_1205 (O_1205,N_19513,N_19614);
nor UO_1206 (O_1206,N_19513,N_19742);
xnor UO_1207 (O_1207,N_19607,N_19514);
nor UO_1208 (O_1208,N_19502,N_19600);
nand UO_1209 (O_1209,N_19533,N_19968);
nand UO_1210 (O_1210,N_19981,N_19539);
nand UO_1211 (O_1211,N_19823,N_19867);
or UO_1212 (O_1212,N_19555,N_19668);
nand UO_1213 (O_1213,N_19920,N_19748);
nor UO_1214 (O_1214,N_19745,N_19693);
nand UO_1215 (O_1215,N_19921,N_19509);
nor UO_1216 (O_1216,N_19662,N_19676);
or UO_1217 (O_1217,N_19676,N_19593);
and UO_1218 (O_1218,N_19783,N_19633);
xor UO_1219 (O_1219,N_19763,N_19616);
nand UO_1220 (O_1220,N_19844,N_19928);
and UO_1221 (O_1221,N_19727,N_19852);
nor UO_1222 (O_1222,N_19856,N_19536);
or UO_1223 (O_1223,N_19624,N_19938);
and UO_1224 (O_1224,N_19985,N_19604);
or UO_1225 (O_1225,N_19920,N_19838);
or UO_1226 (O_1226,N_19935,N_19820);
or UO_1227 (O_1227,N_19870,N_19588);
and UO_1228 (O_1228,N_19810,N_19693);
nand UO_1229 (O_1229,N_19583,N_19596);
nand UO_1230 (O_1230,N_19671,N_19823);
and UO_1231 (O_1231,N_19817,N_19638);
nor UO_1232 (O_1232,N_19882,N_19689);
or UO_1233 (O_1233,N_19901,N_19615);
or UO_1234 (O_1234,N_19905,N_19847);
and UO_1235 (O_1235,N_19565,N_19886);
or UO_1236 (O_1236,N_19563,N_19612);
nor UO_1237 (O_1237,N_19549,N_19855);
or UO_1238 (O_1238,N_19643,N_19557);
nand UO_1239 (O_1239,N_19837,N_19996);
or UO_1240 (O_1240,N_19754,N_19617);
and UO_1241 (O_1241,N_19909,N_19938);
and UO_1242 (O_1242,N_19967,N_19521);
nor UO_1243 (O_1243,N_19870,N_19520);
nor UO_1244 (O_1244,N_19795,N_19826);
or UO_1245 (O_1245,N_19756,N_19887);
or UO_1246 (O_1246,N_19728,N_19501);
nand UO_1247 (O_1247,N_19725,N_19902);
nor UO_1248 (O_1248,N_19584,N_19671);
xnor UO_1249 (O_1249,N_19711,N_19639);
nand UO_1250 (O_1250,N_19846,N_19770);
or UO_1251 (O_1251,N_19549,N_19970);
or UO_1252 (O_1252,N_19801,N_19979);
nor UO_1253 (O_1253,N_19984,N_19546);
and UO_1254 (O_1254,N_19790,N_19739);
nor UO_1255 (O_1255,N_19783,N_19942);
nand UO_1256 (O_1256,N_19815,N_19504);
nor UO_1257 (O_1257,N_19598,N_19977);
and UO_1258 (O_1258,N_19761,N_19981);
nand UO_1259 (O_1259,N_19866,N_19975);
and UO_1260 (O_1260,N_19689,N_19714);
or UO_1261 (O_1261,N_19668,N_19616);
and UO_1262 (O_1262,N_19853,N_19515);
and UO_1263 (O_1263,N_19529,N_19802);
nor UO_1264 (O_1264,N_19990,N_19805);
nand UO_1265 (O_1265,N_19734,N_19849);
nor UO_1266 (O_1266,N_19525,N_19775);
nor UO_1267 (O_1267,N_19860,N_19798);
and UO_1268 (O_1268,N_19893,N_19753);
nand UO_1269 (O_1269,N_19938,N_19879);
and UO_1270 (O_1270,N_19773,N_19599);
and UO_1271 (O_1271,N_19787,N_19932);
nor UO_1272 (O_1272,N_19787,N_19952);
and UO_1273 (O_1273,N_19928,N_19535);
nand UO_1274 (O_1274,N_19513,N_19955);
or UO_1275 (O_1275,N_19741,N_19595);
nor UO_1276 (O_1276,N_19886,N_19920);
nor UO_1277 (O_1277,N_19789,N_19828);
nor UO_1278 (O_1278,N_19756,N_19713);
nand UO_1279 (O_1279,N_19534,N_19786);
nand UO_1280 (O_1280,N_19736,N_19757);
and UO_1281 (O_1281,N_19608,N_19706);
nor UO_1282 (O_1282,N_19971,N_19596);
nand UO_1283 (O_1283,N_19760,N_19880);
xnor UO_1284 (O_1284,N_19699,N_19749);
and UO_1285 (O_1285,N_19673,N_19506);
and UO_1286 (O_1286,N_19736,N_19655);
or UO_1287 (O_1287,N_19710,N_19547);
and UO_1288 (O_1288,N_19662,N_19982);
or UO_1289 (O_1289,N_19502,N_19568);
or UO_1290 (O_1290,N_19772,N_19769);
and UO_1291 (O_1291,N_19988,N_19637);
and UO_1292 (O_1292,N_19813,N_19578);
nor UO_1293 (O_1293,N_19534,N_19614);
nor UO_1294 (O_1294,N_19793,N_19615);
and UO_1295 (O_1295,N_19760,N_19691);
nor UO_1296 (O_1296,N_19892,N_19753);
nor UO_1297 (O_1297,N_19682,N_19990);
nor UO_1298 (O_1298,N_19644,N_19834);
or UO_1299 (O_1299,N_19977,N_19746);
nor UO_1300 (O_1300,N_19737,N_19884);
or UO_1301 (O_1301,N_19785,N_19701);
or UO_1302 (O_1302,N_19517,N_19611);
nand UO_1303 (O_1303,N_19970,N_19928);
and UO_1304 (O_1304,N_19702,N_19623);
nor UO_1305 (O_1305,N_19580,N_19898);
nand UO_1306 (O_1306,N_19618,N_19797);
or UO_1307 (O_1307,N_19750,N_19550);
or UO_1308 (O_1308,N_19886,N_19642);
nor UO_1309 (O_1309,N_19944,N_19602);
nand UO_1310 (O_1310,N_19866,N_19884);
and UO_1311 (O_1311,N_19896,N_19929);
or UO_1312 (O_1312,N_19787,N_19706);
and UO_1313 (O_1313,N_19810,N_19880);
nor UO_1314 (O_1314,N_19906,N_19557);
and UO_1315 (O_1315,N_19602,N_19679);
or UO_1316 (O_1316,N_19543,N_19762);
and UO_1317 (O_1317,N_19516,N_19948);
nor UO_1318 (O_1318,N_19946,N_19662);
or UO_1319 (O_1319,N_19920,N_19552);
nor UO_1320 (O_1320,N_19854,N_19758);
and UO_1321 (O_1321,N_19810,N_19889);
nor UO_1322 (O_1322,N_19618,N_19589);
and UO_1323 (O_1323,N_19513,N_19561);
or UO_1324 (O_1324,N_19870,N_19702);
and UO_1325 (O_1325,N_19666,N_19901);
nand UO_1326 (O_1326,N_19957,N_19770);
nor UO_1327 (O_1327,N_19696,N_19811);
nor UO_1328 (O_1328,N_19972,N_19569);
and UO_1329 (O_1329,N_19718,N_19866);
nor UO_1330 (O_1330,N_19575,N_19563);
or UO_1331 (O_1331,N_19727,N_19782);
and UO_1332 (O_1332,N_19714,N_19635);
nor UO_1333 (O_1333,N_19692,N_19926);
or UO_1334 (O_1334,N_19736,N_19931);
nor UO_1335 (O_1335,N_19709,N_19684);
or UO_1336 (O_1336,N_19569,N_19776);
and UO_1337 (O_1337,N_19515,N_19762);
nand UO_1338 (O_1338,N_19725,N_19737);
or UO_1339 (O_1339,N_19866,N_19655);
nand UO_1340 (O_1340,N_19694,N_19739);
and UO_1341 (O_1341,N_19974,N_19588);
nand UO_1342 (O_1342,N_19877,N_19827);
nand UO_1343 (O_1343,N_19624,N_19880);
nor UO_1344 (O_1344,N_19664,N_19585);
and UO_1345 (O_1345,N_19698,N_19910);
and UO_1346 (O_1346,N_19972,N_19815);
and UO_1347 (O_1347,N_19886,N_19955);
or UO_1348 (O_1348,N_19725,N_19893);
or UO_1349 (O_1349,N_19569,N_19942);
nor UO_1350 (O_1350,N_19500,N_19968);
and UO_1351 (O_1351,N_19868,N_19750);
and UO_1352 (O_1352,N_19999,N_19600);
nand UO_1353 (O_1353,N_19990,N_19907);
nor UO_1354 (O_1354,N_19529,N_19795);
and UO_1355 (O_1355,N_19937,N_19814);
nand UO_1356 (O_1356,N_19979,N_19658);
or UO_1357 (O_1357,N_19938,N_19828);
nor UO_1358 (O_1358,N_19966,N_19955);
nand UO_1359 (O_1359,N_19744,N_19566);
or UO_1360 (O_1360,N_19762,N_19694);
nand UO_1361 (O_1361,N_19698,N_19605);
and UO_1362 (O_1362,N_19552,N_19611);
nor UO_1363 (O_1363,N_19892,N_19796);
and UO_1364 (O_1364,N_19614,N_19503);
and UO_1365 (O_1365,N_19774,N_19839);
or UO_1366 (O_1366,N_19903,N_19567);
nor UO_1367 (O_1367,N_19612,N_19665);
nor UO_1368 (O_1368,N_19737,N_19870);
and UO_1369 (O_1369,N_19671,N_19551);
or UO_1370 (O_1370,N_19615,N_19989);
and UO_1371 (O_1371,N_19637,N_19918);
nor UO_1372 (O_1372,N_19740,N_19623);
and UO_1373 (O_1373,N_19891,N_19743);
nand UO_1374 (O_1374,N_19757,N_19891);
and UO_1375 (O_1375,N_19816,N_19961);
nand UO_1376 (O_1376,N_19731,N_19720);
and UO_1377 (O_1377,N_19873,N_19580);
nor UO_1378 (O_1378,N_19913,N_19537);
nand UO_1379 (O_1379,N_19881,N_19912);
or UO_1380 (O_1380,N_19730,N_19531);
nand UO_1381 (O_1381,N_19552,N_19964);
or UO_1382 (O_1382,N_19982,N_19680);
nand UO_1383 (O_1383,N_19611,N_19935);
and UO_1384 (O_1384,N_19642,N_19710);
or UO_1385 (O_1385,N_19850,N_19845);
nand UO_1386 (O_1386,N_19551,N_19523);
nand UO_1387 (O_1387,N_19732,N_19979);
and UO_1388 (O_1388,N_19896,N_19652);
xor UO_1389 (O_1389,N_19509,N_19860);
and UO_1390 (O_1390,N_19788,N_19811);
nand UO_1391 (O_1391,N_19764,N_19710);
nand UO_1392 (O_1392,N_19830,N_19952);
nor UO_1393 (O_1393,N_19967,N_19566);
nor UO_1394 (O_1394,N_19602,N_19693);
nand UO_1395 (O_1395,N_19913,N_19746);
nor UO_1396 (O_1396,N_19725,N_19584);
or UO_1397 (O_1397,N_19543,N_19800);
nor UO_1398 (O_1398,N_19873,N_19548);
xor UO_1399 (O_1399,N_19537,N_19982);
or UO_1400 (O_1400,N_19864,N_19516);
nand UO_1401 (O_1401,N_19831,N_19584);
or UO_1402 (O_1402,N_19944,N_19994);
and UO_1403 (O_1403,N_19950,N_19991);
and UO_1404 (O_1404,N_19943,N_19894);
nor UO_1405 (O_1405,N_19569,N_19568);
and UO_1406 (O_1406,N_19650,N_19884);
and UO_1407 (O_1407,N_19837,N_19825);
nor UO_1408 (O_1408,N_19646,N_19736);
nand UO_1409 (O_1409,N_19977,N_19667);
and UO_1410 (O_1410,N_19909,N_19554);
nand UO_1411 (O_1411,N_19711,N_19745);
nand UO_1412 (O_1412,N_19925,N_19924);
and UO_1413 (O_1413,N_19989,N_19712);
and UO_1414 (O_1414,N_19697,N_19766);
nand UO_1415 (O_1415,N_19782,N_19974);
or UO_1416 (O_1416,N_19687,N_19868);
nor UO_1417 (O_1417,N_19544,N_19894);
nand UO_1418 (O_1418,N_19971,N_19510);
or UO_1419 (O_1419,N_19793,N_19580);
nand UO_1420 (O_1420,N_19667,N_19671);
nor UO_1421 (O_1421,N_19651,N_19991);
and UO_1422 (O_1422,N_19710,N_19993);
nand UO_1423 (O_1423,N_19839,N_19546);
nor UO_1424 (O_1424,N_19752,N_19826);
and UO_1425 (O_1425,N_19676,N_19814);
and UO_1426 (O_1426,N_19782,N_19527);
nand UO_1427 (O_1427,N_19555,N_19698);
nor UO_1428 (O_1428,N_19724,N_19814);
nand UO_1429 (O_1429,N_19608,N_19659);
or UO_1430 (O_1430,N_19571,N_19630);
nand UO_1431 (O_1431,N_19624,N_19565);
xor UO_1432 (O_1432,N_19820,N_19765);
nand UO_1433 (O_1433,N_19976,N_19845);
nand UO_1434 (O_1434,N_19976,N_19602);
or UO_1435 (O_1435,N_19696,N_19590);
or UO_1436 (O_1436,N_19995,N_19905);
and UO_1437 (O_1437,N_19633,N_19795);
and UO_1438 (O_1438,N_19771,N_19925);
and UO_1439 (O_1439,N_19617,N_19998);
nand UO_1440 (O_1440,N_19857,N_19744);
nor UO_1441 (O_1441,N_19619,N_19851);
and UO_1442 (O_1442,N_19812,N_19673);
and UO_1443 (O_1443,N_19655,N_19801);
or UO_1444 (O_1444,N_19935,N_19984);
or UO_1445 (O_1445,N_19728,N_19830);
nand UO_1446 (O_1446,N_19641,N_19842);
nand UO_1447 (O_1447,N_19540,N_19503);
xnor UO_1448 (O_1448,N_19713,N_19768);
nand UO_1449 (O_1449,N_19845,N_19533);
xor UO_1450 (O_1450,N_19696,N_19766);
nand UO_1451 (O_1451,N_19709,N_19882);
and UO_1452 (O_1452,N_19701,N_19537);
and UO_1453 (O_1453,N_19607,N_19969);
nor UO_1454 (O_1454,N_19837,N_19766);
nand UO_1455 (O_1455,N_19986,N_19692);
and UO_1456 (O_1456,N_19853,N_19615);
nand UO_1457 (O_1457,N_19996,N_19643);
nand UO_1458 (O_1458,N_19668,N_19928);
nor UO_1459 (O_1459,N_19925,N_19717);
and UO_1460 (O_1460,N_19917,N_19524);
nor UO_1461 (O_1461,N_19625,N_19771);
and UO_1462 (O_1462,N_19703,N_19517);
and UO_1463 (O_1463,N_19709,N_19504);
or UO_1464 (O_1464,N_19567,N_19507);
nor UO_1465 (O_1465,N_19795,N_19678);
nand UO_1466 (O_1466,N_19662,N_19720);
nand UO_1467 (O_1467,N_19853,N_19802);
nor UO_1468 (O_1468,N_19796,N_19793);
nand UO_1469 (O_1469,N_19952,N_19690);
and UO_1470 (O_1470,N_19611,N_19869);
nand UO_1471 (O_1471,N_19602,N_19895);
nor UO_1472 (O_1472,N_19611,N_19785);
nor UO_1473 (O_1473,N_19555,N_19640);
nand UO_1474 (O_1474,N_19811,N_19753);
or UO_1475 (O_1475,N_19671,N_19701);
nor UO_1476 (O_1476,N_19566,N_19628);
or UO_1477 (O_1477,N_19543,N_19513);
nand UO_1478 (O_1478,N_19664,N_19576);
nor UO_1479 (O_1479,N_19846,N_19981);
nor UO_1480 (O_1480,N_19631,N_19987);
nand UO_1481 (O_1481,N_19891,N_19996);
or UO_1482 (O_1482,N_19787,N_19649);
and UO_1483 (O_1483,N_19590,N_19915);
nand UO_1484 (O_1484,N_19661,N_19871);
or UO_1485 (O_1485,N_19509,N_19570);
and UO_1486 (O_1486,N_19832,N_19973);
or UO_1487 (O_1487,N_19664,N_19949);
nor UO_1488 (O_1488,N_19693,N_19995);
nor UO_1489 (O_1489,N_19529,N_19953);
nand UO_1490 (O_1490,N_19981,N_19991);
and UO_1491 (O_1491,N_19805,N_19551);
xor UO_1492 (O_1492,N_19971,N_19566);
nand UO_1493 (O_1493,N_19988,N_19964);
nor UO_1494 (O_1494,N_19962,N_19736);
nor UO_1495 (O_1495,N_19630,N_19593);
nor UO_1496 (O_1496,N_19773,N_19946);
nand UO_1497 (O_1497,N_19709,N_19804);
or UO_1498 (O_1498,N_19838,N_19591);
nand UO_1499 (O_1499,N_19624,N_19719);
and UO_1500 (O_1500,N_19738,N_19958);
nor UO_1501 (O_1501,N_19803,N_19685);
and UO_1502 (O_1502,N_19880,N_19521);
and UO_1503 (O_1503,N_19772,N_19898);
nor UO_1504 (O_1504,N_19673,N_19779);
nand UO_1505 (O_1505,N_19875,N_19586);
nor UO_1506 (O_1506,N_19665,N_19522);
nor UO_1507 (O_1507,N_19911,N_19519);
nand UO_1508 (O_1508,N_19758,N_19992);
and UO_1509 (O_1509,N_19666,N_19927);
and UO_1510 (O_1510,N_19752,N_19622);
nor UO_1511 (O_1511,N_19768,N_19786);
nor UO_1512 (O_1512,N_19943,N_19710);
or UO_1513 (O_1513,N_19783,N_19851);
and UO_1514 (O_1514,N_19801,N_19726);
nor UO_1515 (O_1515,N_19819,N_19714);
nor UO_1516 (O_1516,N_19659,N_19985);
nand UO_1517 (O_1517,N_19819,N_19685);
and UO_1518 (O_1518,N_19523,N_19712);
nand UO_1519 (O_1519,N_19705,N_19624);
or UO_1520 (O_1520,N_19708,N_19928);
and UO_1521 (O_1521,N_19885,N_19544);
and UO_1522 (O_1522,N_19811,N_19962);
nand UO_1523 (O_1523,N_19603,N_19558);
nor UO_1524 (O_1524,N_19609,N_19659);
nand UO_1525 (O_1525,N_19936,N_19519);
nand UO_1526 (O_1526,N_19696,N_19987);
or UO_1527 (O_1527,N_19679,N_19697);
and UO_1528 (O_1528,N_19590,N_19791);
nand UO_1529 (O_1529,N_19952,N_19838);
nor UO_1530 (O_1530,N_19862,N_19507);
or UO_1531 (O_1531,N_19724,N_19803);
nor UO_1532 (O_1532,N_19996,N_19794);
nor UO_1533 (O_1533,N_19982,N_19841);
nand UO_1534 (O_1534,N_19654,N_19893);
and UO_1535 (O_1535,N_19680,N_19515);
or UO_1536 (O_1536,N_19604,N_19506);
or UO_1537 (O_1537,N_19687,N_19936);
or UO_1538 (O_1538,N_19761,N_19862);
or UO_1539 (O_1539,N_19548,N_19898);
nor UO_1540 (O_1540,N_19789,N_19762);
or UO_1541 (O_1541,N_19686,N_19589);
or UO_1542 (O_1542,N_19953,N_19913);
xnor UO_1543 (O_1543,N_19968,N_19675);
or UO_1544 (O_1544,N_19835,N_19542);
nand UO_1545 (O_1545,N_19891,N_19618);
and UO_1546 (O_1546,N_19989,N_19742);
nand UO_1547 (O_1547,N_19771,N_19819);
nand UO_1548 (O_1548,N_19757,N_19596);
nand UO_1549 (O_1549,N_19935,N_19629);
or UO_1550 (O_1550,N_19839,N_19583);
and UO_1551 (O_1551,N_19556,N_19687);
nand UO_1552 (O_1552,N_19703,N_19616);
and UO_1553 (O_1553,N_19998,N_19628);
or UO_1554 (O_1554,N_19664,N_19853);
nor UO_1555 (O_1555,N_19633,N_19727);
or UO_1556 (O_1556,N_19593,N_19737);
nor UO_1557 (O_1557,N_19524,N_19563);
and UO_1558 (O_1558,N_19797,N_19757);
nand UO_1559 (O_1559,N_19985,N_19831);
nor UO_1560 (O_1560,N_19663,N_19702);
nor UO_1561 (O_1561,N_19603,N_19664);
or UO_1562 (O_1562,N_19560,N_19892);
nand UO_1563 (O_1563,N_19816,N_19748);
nor UO_1564 (O_1564,N_19696,N_19856);
or UO_1565 (O_1565,N_19879,N_19658);
or UO_1566 (O_1566,N_19957,N_19551);
nor UO_1567 (O_1567,N_19700,N_19888);
and UO_1568 (O_1568,N_19579,N_19803);
nor UO_1569 (O_1569,N_19966,N_19901);
nand UO_1570 (O_1570,N_19912,N_19907);
or UO_1571 (O_1571,N_19939,N_19637);
and UO_1572 (O_1572,N_19575,N_19861);
nand UO_1573 (O_1573,N_19938,N_19865);
and UO_1574 (O_1574,N_19829,N_19761);
xnor UO_1575 (O_1575,N_19854,N_19908);
and UO_1576 (O_1576,N_19822,N_19641);
or UO_1577 (O_1577,N_19832,N_19853);
nor UO_1578 (O_1578,N_19806,N_19564);
and UO_1579 (O_1579,N_19710,N_19918);
and UO_1580 (O_1580,N_19958,N_19767);
and UO_1581 (O_1581,N_19536,N_19729);
nand UO_1582 (O_1582,N_19663,N_19817);
and UO_1583 (O_1583,N_19792,N_19720);
or UO_1584 (O_1584,N_19771,N_19504);
and UO_1585 (O_1585,N_19854,N_19863);
nand UO_1586 (O_1586,N_19563,N_19553);
and UO_1587 (O_1587,N_19955,N_19981);
or UO_1588 (O_1588,N_19808,N_19999);
and UO_1589 (O_1589,N_19889,N_19962);
and UO_1590 (O_1590,N_19552,N_19846);
or UO_1591 (O_1591,N_19768,N_19781);
and UO_1592 (O_1592,N_19823,N_19857);
nand UO_1593 (O_1593,N_19583,N_19741);
and UO_1594 (O_1594,N_19956,N_19646);
or UO_1595 (O_1595,N_19955,N_19882);
and UO_1596 (O_1596,N_19582,N_19664);
xor UO_1597 (O_1597,N_19516,N_19560);
nand UO_1598 (O_1598,N_19899,N_19925);
and UO_1599 (O_1599,N_19678,N_19974);
and UO_1600 (O_1600,N_19943,N_19834);
or UO_1601 (O_1601,N_19740,N_19763);
and UO_1602 (O_1602,N_19814,N_19958);
nand UO_1603 (O_1603,N_19689,N_19717);
nor UO_1604 (O_1604,N_19681,N_19857);
and UO_1605 (O_1605,N_19979,N_19542);
nor UO_1606 (O_1606,N_19720,N_19937);
and UO_1607 (O_1607,N_19527,N_19804);
nor UO_1608 (O_1608,N_19948,N_19688);
xnor UO_1609 (O_1609,N_19642,N_19584);
and UO_1610 (O_1610,N_19961,N_19809);
nand UO_1611 (O_1611,N_19560,N_19811);
nand UO_1612 (O_1612,N_19924,N_19773);
or UO_1613 (O_1613,N_19782,N_19508);
nand UO_1614 (O_1614,N_19611,N_19822);
nor UO_1615 (O_1615,N_19561,N_19781);
or UO_1616 (O_1616,N_19877,N_19699);
or UO_1617 (O_1617,N_19580,N_19573);
and UO_1618 (O_1618,N_19649,N_19757);
nor UO_1619 (O_1619,N_19509,N_19604);
nor UO_1620 (O_1620,N_19721,N_19820);
and UO_1621 (O_1621,N_19728,N_19865);
or UO_1622 (O_1622,N_19917,N_19541);
or UO_1623 (O_1623,N_19987,N_19580);
nor UO_1624 (O_1624,N_19606,N_19963);
or UO_1625 (O_1625,N_19791,N_19871);
or UO_1626 (O_1626,N_19757,N_19611);
or UO_1627 (O_1627,N_19764,N_19680);
nor UO_1628 (O_1628,N_19861,N_19904);
or UO_1629 (O_1629,N_19559,N_19572);
or UO_1630 (O_1630,N_19707,N_19595);
nor UO_1631 (O_1631,N_19744,N_19938);
nor UO_1632 (O_1632,N_19926,N_19688);
and UO_1633 (O_1633,N_19534,N_19801);
nor UO_1634 (O_1634,N_19910,N_19989);
or UO_1635 (O_1635,N_19581,N_19632);
and UO_1636 (O_1636,N_19815,N_19531);
and UO_1637 (O_1637,N_19602,N_19790);
or UO_1638 (O_1638,N_19536,N_19986);
or UO_1639 (O_1639,N_19825,N_19900);
nor UO_1640 (O_1640,N_19735,N_19793);
or UO_1641 (O_1641,N_19595,N_19815);
or UO_1642 (O_1642,N_19673,N_19554);
nand UO_1643 (O_1643,N_19712,N_19740);
nor UO_1644 (O_1644,N_19788,N_19764);
nor UO_1645 (O_1645,N_19586,N_19788);
or UO_1646 (O_1646,N_19720,N_19577);
and UO_1647 (O_1647,N_19960,N_19735);
and UO_1648 (O_1648,N_19613,N_19761);
nor UO_1649 (O_1649,N_19652,N_19565);
and UO_1650 (O_1650,N_19601,N_19564);
nor UO_1651 (O_1651,N_19874,N_19941);
nand UO_1652 (O_1652,N_19550,N_19597);
nor UO_1653 (O_1653,N_19603,N_19948);
or UO_1654 (O_1654,N_19809,N_19986);
nor UO_1655 (O_1655,N_19763,N_19879);
nand UO_1656 (O_1656,N_19815,N_19763);
and UO_1657 (O_1657,N_19813,N_19506);
nand UO_1658 (O_1658,N_19649,N_19524);
nand UO_1659 (O_1659,N_19658,N_19569);
and UO_1660 (O_1660,N_19942,N_19632);
nor UO_1661 (O_1661,N_19765,N_19916);
nor UO_1662 (O_1662,N_19553,N_19605);
nand UO_1663 (O_1663,N_19841,N_19968);
nand UO_1664 (O_1664,N_19539,N_19860);
and UO_1665 (O_1665,N_19859,N_19605);
nand UO_1666 (O_1666,N_19714,N_19657);
or UO_1667 (O_1667,N_19683,N_19848);
nand UO_1668 (O_1668,N_19894,N_19557);
nor UO_1669 (O_1669,N_19686,N_19658);
and UO_1670 (O_1670,N_19570,N_19913);
nor UO_1671 (O_1671,N_19571,N_19782);
nor UO_1672 (O_1672,N_19818,N_19535);
nand UO_1673 (O_1673,N_19514,N_19678);
nor UO_1674 (O_1674,N_19511,N_19973);
nand UO_1675 (O_1675,N_19832,N_19979);
or UO_1676 (O_1676,N_19671,N_19593);
nor UO_1677 (O_1677,N_19995,N_19676);
and UO_1678 (O_1678,N_19849,N_19974);
or UO_1679 (O_1679,N_19925,N_19867);
and UO_1680 (O_1680,N_19843,N_19725);
nand UO_1681 (O_1681,N_19706,N_19545);
and UO_1682 (O_1682,N_19749,N_19632);
nor UO_1683 (O_1683,N_19730,N_19772);
and UO_1684 (O_1684,N_19785,N_19771);
nor UO_1685 (O_1685,N_19965,N_19658);
and UO_1686 (O_1686,N_19585,N_19967);
nor UO_1687 (O_1687,N_19747,N_19547);
nand UO_1688 (O_1688,N_19808,N_19552);
and UO_1689 (O_1689,N_19695,N_19516);
and UO_1690 (O_1690,N_19986,N_19796);
or UO_1691 (O_1691,N_19833,N_19676);
nor UO_1692 (O_1692,N_19841,N_19510);
nor UO_1693 (O_1693,N_19787,N_19551);
or UO_1694 (O_1694,N_19944,N_19625);
or UO_1695 (O_1695,N_19903,N_19882);
nand UO_1696 (O_1696,N_19887,N_19743);
nand UO_1697 (O_1697,N_19544,N_19671);
and UO_1698 (O_1698,N_19887,N_19826);
nor UO_1699 (O_1699,N_19963,N_19883);
or UO_1700 (O_1700,N_19612,N_19784);
and UO_1701 (O_1701,N_19671,N_19715);
nor UO_1702 (O_1702,N_19990,N_19795);
or UO_1703 (O_1703,N_19800,N_19928);
nor UO_1704 (O_1704,N_19575,N_19738);
nor UO_1705 (O_1705,N_19988,N_19809);
and UO_1706 (O_1706,N_19552,N_19896);
or UO_1707 (O_1707,N_19611,N_19929);
or UO_1708 (O_1708,N_19883,N_19867);
xor UO_1709 (O_1709,N_19801,N_19735);
nor UO_1710 (O_1710,N_19529,N_19723);
and UO_1711 (O_1711,N_19876,N_19746);
or UO_1712 (O_1712,N_19685,N_19668);
nand UO_1713 (O_1713,N_19648,N_19919);
or UO_1714 (O_1714,N_19586,N_19946);
and UO_1715 (O_1715,N_19637,N_19963);
nand UO_1716 (O_1716,N_19533,N_19667);
or UO_1717 (O_1717,N_19928,N_19728);
and UO_1718 (O_1718,N_19791,N_19759);
and UO_1719 (O_1719,N_19836,N_19997);
nor UO_1720 (O_1720,N_19565,N_19766);
and UO_1721 (O_1721,N_19946,N_19573);
and UO_1722 (O_1722,N_19510,N_19675);
nor UO_1723 (O_1723,N_19815,N_19770);
and UO_1724 (O_1724,N_19574,N_19955);
xor UO_1725 (O_1725,N_19764,N_19594);
or UO_1726 (O_1726,N_19948,N_19899);
or UO_1727 (O_1727,N_19530,N_19985);
nor UO_1728 (O_1728,N_19567,N_19777);
nor UO_1729 (O_1729,N_19525,N_19569);
and UO_1730 (O_1730,N_19959,N_19746);
nor UO_1731 (O_1731,N_19909,N_19865);
nand UO_1732 (O_1732,N_19876,N_19755);
nor UO_1733 (O_1733,N_19541,N_19988);
and UO_1734 (O_1734,N_19598,N_19711);
or UO_1735 (O_1735,N_19899,N_19850);
or UO_1736 (O_1736,N_19612,N_19684);
and UO_1737 (O_1737,N_19749,N_19509);
or UO_1738 (O_1738,N_19653,N_19909);
and UO_1739 (O_1739,N_19790,N_19553);
xor UO_1740 (O_1740,N_19950,N_19879);
nand UO_1741 (O_1741,N_19715,N_19951);
and UO_1742 (O_1742,N_19766,N_19681);
nor UO_1743 (O_1743,N_19554,N_19670);
or UO_1744 (O_1744,N_19951,N_19545);
or UO_1745 (O_1745,N_19674,N_19891);
nand UO_1746 (O_1746,N_19629,N_19754);
or UO_1747 (O_1747,N_19673,N_19802);
nand UO_1748 (O_1748,N_19511,N_19567);
nand UO_1749 (O_1749,N_19891,N_19568);
nor UO_1750 (O_1750,N_19768,N_19901);
nand UO_1751 (O_1751,N_19902,N_19762);
and UO_1752 (O_1752,N_19742,N_19674);
and UO_1753 (O_1753,N_19717,N_19983);
nor UO_1754 (O_1754,N_19529,N_19756);
or UO_1755 (O_1755,N_19509,N_19659);
nor UO_1756 (O_1756,N_19572,N_19575);
nand UO_1757 (O_1757,N_19963,N_19572);
nor UO_1758 (O_1758,N_19613,N_19656);
nand UO_1759 (O_1759,N_19562,N_19635);
or UO_1760 (O_1760,N_19857,N_19758);
and UO_1761 (O_1761,N_19520,N_19556);
and UO_1762 (O_1762,N_19619,N_19716);
and UO_1763 (O_1763,N_19810,N_19814);
or UO_1764 (O_1764,N_19571,N_19751);
or UO_1765 (O_1765,N_19909,N_19843);
nand UO_1766 (O_1766,N_19606,N_19842);
nand UO_1767 (O_1767,N_19920,N_19948);
or UO_1768 (O_1768,N_19643,N_19539);
and UO_1769 (O_1769,N_19632,N_19566);
or UO_1770 (O_1770,N_19783,N_19600);
nor UO_1771 (O_1771,N_19895,N_19697);
nor UO_1772 (O_1772,N_19842,N_19857);
or UO_1773 (O_1773,N_19625,N_19961);
nor UO_1774 (O_1774,N_19697,N_19863);
nor UO_1775 (O_1775,N_19654,N_19978);
nor UO_1776 (O_1776,N_19648,N_19594);
or UO_1777 (O_1777,N_19928,N_19849);
nor UO_1778 (O_1778,N_19610,N_19741);
or UO_1779 (O_1779,N_19742,N_19559);
nand UO_1780 (O_1780,N_19633,N_19616);
xor UO_1781 (O_1781,N_19854,N_19963);
or UO_1782 (O_1782,N_19989,N_19873);
and UO_1783 (O_1783,N_19941,N_19538);
or UO_1784 (O_1784,N_19686,N_19784);
and UO_1785 (O_1785,N_19832,N_19653);
nor UO_1786 (O_1786,N_19759,N_19944);
nor UO_1787 (O_1787,N_19578,N_19865);
nor UO_1788 (O_1788,N_19624,N_19903);
xnor UO_1789 (O_1789,N_19755,N_19814);
and UO_1790 (O_1790,N_19956,N_19939);
and UO_1791 (O_1791,N_19632,N_19832);
nand UO_1792 (O_1792,N_19597,N_19796);
nand UO_1793 (O_1793,N_19629,N_19547);
or UO_1794 (O_1794,N_19703,N_19654);
nand UO_1795 (O_1795,N_19888,N_19631);
nor UO_1796 (O_1796,N_19577,N_19518);
and UO_1797 (O_1797,N_19771,N_19911);
and UO_1798 (O_1798,N_19685,N_19593);
and UO_1799 (O_1799,N_19730,N_19872);
nand UO_1800 (O_1800,N_19531,N_19979);
and UO_1801 (O_1801,N_19901,N_19670);
or UO_1802 (O_1802,N_19510,N_19608);
and UO_1803 (O_1803,N_19688,N_19693);
nand UO_1804 (O_1804,N_19551,N_19777);
nand UO_1805 (O_1805,N_19771,N_19513);
nor UO_1806 (O_1806,N_19846,N_19602);
nand UO_1807 (O_1807,N_19502,N_19856);
and UO_1808 (O_1808,N_19647,N_19799);
and UO_1809 (O_1809,N_19552,N_19596);
and UO_1810 (O_1810,N_19528,N_19887);
and UO_1811 (O_1811,N_19714,N_19632);
and UO_1812 (O_1812,N_19711,N_19543);
nor UO_1813 (O_1813,N_19781,N_19816);
and UO_1814 (O_1814,N_19604,N_19563);
nand UO_1815 (O_1815,N_19805,N_19531);
or UO_1816 (O_1816,N_19832,N_19974);
nand UO_1817 (O_1817,N_19860,N_19556);
nand UO_1818 (O_1818,N_19524,N_19659);
nor UO_1819 (O_1819,N_19801,N_19528);
or UO_1820 (O_1820,N_19888,N_19926);
xnor UO_1821 (O_1821,N_19527,N_19531);
nand UO_1822 (O_1822,N_19539,N_19904);
nand UO_1823 (O_1823,N_19922,N_19654);
or UO_1824 (O_1824,N_19723,N_19603);
nand UO_1825 (O_1825,N_19918,N_19739);
nor UO_1826 (O_1826,N_19953,N_19830);
nand UO_1827 (O_1827,N_19659,N_19724);
nand UO_1828 (O_1828,N_19950,N_19590);
and UO_1829 (O_1829,N_19955,N_19506);
nand UO_1830 (O_1830,N_19635,N_19601);
or UO_1831 (O_1831,N_19762,N_19783);
nand UO_1832 (O_1832,N_19797,N_19648);
or UO_1833 (O_1833,N_19596,N_19723);
or UO_1834 (O_1834,N_19891,N_19663);
and UO_1835 (O_1835,N_19578,N_19591);
nor UO_1836 (O_1836,N_19836,N_19765);
and UO_1837 (O_1837,N_19763,N_19687);
nand UO_1838 (O_1838,N_19682,N_19805);
nor UO_1839 (O_1839,N_19567,N_19765);
nor UO_1840 (O_1840,N_19654,N_19529);
nand UO_1841 (O_1841,N_19520,N_19930);
nand UO_1842 (O_1842,N_19650,N_19930);
or UO_1843 (O_1843,N_19814,N_19686);
and UO_1844 (O_1844,N_19776,N_19657);
or UO_1845 (O_1845,N_19736,N_19540);
and UO_1846 (O_1846,N_19695,N_19941);
and UO_1847 (O_1847,N_19542,N_19697);
nor UO_1848 (O_1848,N_19754,N_19799);
or UO_1849 (O_1849,N_19709,N_19537);
nand UO_1850 (O_1850,N_19575,N_19751);
nor UO_1851 (O_1851,N_19851,N_19764);
nand UO_1852 (O_1852,N_19635,N_19662);
nor UO_1853 (O_1853,N_19786,N_19927);
nand UO_1854 (O_1854,N_19886,N_19852);
or UO_1855 (O_1855,N_19569,N_19883);
nand UO_1856 (O_1856,N_19959,N_19634);
or UO_1857 (O_1857,N_19645,N_19875);
nand UO_1858 (O_1858,N_19633,N_19661);
and UO_1859 (O_1859,N_19764,N_19645);
nor UO_1860 (O_1860,N_19724,N_19575);
or UO_1861 (O_1861,N_19636,N_19568);
nand UO_1862 (O_1862,N_19905,N_19593);
and UO_1863 (O_1863,N_19708,N_19923);
or UO_1864 (O_1864,N_19927,N_19532);
and UO_1865 (O_1865,N_19791,N_19549);
nand UO_1866 (O_1866,N_19525,N_19804);
nor UO_1867 (O_1867,N_19973,N_19848);
nor UO_1868 (O_1868,N_19523,N_19952);
and UO_1869 (O_1869,N_19983,N_19605);
nand UO_1870 (O_1870,N_19514,N_19853);
nor UO_1871 (O_1871,N_19731,N_19578);
nor UO_1872 (O_1872,N_19829,N_19860);
nor UO_1873 (O_1873,N_19588,N_19922);
or UO_1874 (O_1874,N_19818,N_19809);
nor UO_1875 (O_1875,N_19564,N_19522);
nand UO_1876 (O_1876,N_19674,N_19834);
nor UO_1877 (O_1877,N_19526,N_19686);
or UO_1878 (O_1878,N_19627,N_19841);
or UO_1879 (O_1879,N_19884,N_19891);
nand UO_1880 (O_1880,N_19843,N_19556);
and UO_1881 (O_1881,N_19606,N_19875);
nor UO_1882 (O_1882,N_19749,N_19814);
nor UO_1883 (O_1883,N_19899,N_19770);
and UO_1884 (O_1884,N_19840,N_19847);
nor UO_1885 (O_1885,N_19907,N_19816);
nand UO_1886 (O_1886,N_19758,N_19795);
and UO_1887 (O_1887,N_19670,N_19797);
nand UO_1888 (O_1888,N_19929,N_19853);
or UO_1889 (O_1889,N_19545,N_19633);
or UO_1890 (O_1890,N_19636,N_19787);
or UO_1891 (O_1891,N_19651,N_19734);
nor UO_1892 (O_1892,N_19713,N_19535);
nand UO_1893 (O_1893,N_19837,N_19712);
nand UO_1894 (O_1894,N_19761,N_19530);
and UO_1895 (O_1895,N_19986,N_19833);
or UO_1896 (O_1896,N_19869,N_19860);
nand UO_1897 (O_1897,N_19645,N_19883);
and UO_1898 (O_1898,N_19714,N_19963);
nand UO_1899 (O_1899,N_19623,N_19795);
and UO_1900 (O_1900,N_19542,N_19715);
or UO_1901 (O_1901,N_19539,N_19711);
nand UO_1902 (O_1902,N_19649,N_19752);
xor UO_1903 (O_1903,N_19815,N_19796);
and UO_1904 (O_1904,N_19644,N_19692);
and UO_1905 (O_1905,N_19579,N_19536);
and UO_1906 (O_1906,N_19914,N_19540);
or UO_1907 (O_1907,N_19852,N_19749);
and UO_1908 (O_1908,N_19928,N_19967);
and UO_1909 (O_1909,N_19689,N_19782);
nor UO_1910 (O_1910,N_19571,N_19757);
or UO_1911 (O_1911,N_19680,N_19807);
nand UO_1912 (O_1912,N_19701,N_19534);
and UO_1913 (O_1913,N_19771,N_19755);
and UO_1914 (O_1914,N_19576,N_19833);
and UO_1915 (O_1915,N_19881,N_19673);
xnor UO_1916 (O_1916,N_19506,N_19919);
nor UO_1917 (O_1917,N_19665,N_19830);
or UO_1918 (O_1918,N_19687,N_19637);
and UO_1919 (O_1919,N_19671,N_19601);
nand UO_1920 (O_1920,N_19970,N_19663);
nand UO_1921 (O_1921,N_19979,N_19521);
nor UO_1922 (O_1922,N_19794,N_19926);
and UO_1923 (O_1923,N_19579,N_19964);
nand UO_1924 (O_1924,N_19615,N_19508);
nor UO_1925 (O_1925,N_19880,N_19569);
nor UO_1926 (O_1926,N_19782,N_19952);
and UO_1927 (O_1927,N_19869,N_19835);
or UO_1928 (O_1928,N_19928,N_19665);
nor UO_1929 (O_1929,N_19729,N_19683);
or UO_1930 (O_1930,N_19719,N_19969);
or UO_1931 (O_1931,N_19535,N_19897);
and UO_1932 (O_1932,N_19897,N_19909);
nor UO_1933 (O_1933,N_19728,N_19739);
and UO_1934 (O_1934,N_19901,N_19993);
or UO_1935 (O_1935,N_19540,N_19684);
nor UO_1936 (O_1936,N_19811,N_19834);
or UO_1937 (O_1937,N_19892,N_19731);
and UO_1938 (O_1938,N_19500,N_19507);
nand UO_1939 (O_1939,N_19666,N_19583);
nor UO_1940 (O_1940,N_19758,N_19905);
or UO_1941 (O_1941,N_19831,N_19824);
nand UO_1942 (O_1942,N_19751,N_19568);
and UO_1943 (O_1943,N_19901,N_19593);
or UO_1944 (O_1944,N_19627,N_19834);
nand UO_1945 (O_1945,N_19727,N_19868);
and UO_1946 (O_1946,N_19847,N_19561);
or UO_1947 (O_1947,N_19529,N_19927);
nand UO_1948 (O_1948,N_19759,N_19952);
nand UO_1949 (O_1949,N_19801,N_19927);
or UO_1950 (O_1950,N_19707,N_19851);
nor UO_1951 (O_1951,N_19642,N_19560);
and UO_1952 (O_1952,N_19808,N_19939);
nor UO_1953 (O_1953,N_19530,N_19941);
or UO_1954 (O_1954,N_19858,N_19997);
or UO_1955 (O_1955,N_19678,N_19878);
or UO_1956 (O_1956,N_19554,N_19729);
or UO_1957 (O_1957,N_19957,N_19710);
or UO_1958 (O_1958,N_19903,N_19571);
and UO_1959 (O_1959,N_19991,N_19862);
nand UO_1960 (O_1960,N_19884,N_19816);
nor UO_1961 (O_1961,N_19741,N_19921);
xor UO_1962 (O_1962,N_19507,N_19624);
or UO_1963 (O_1963,N_19844,N_19944);
nor UO_1964 (O_1964,N_19800,N_19841);
nand UO_1965 (O_1965,N_19836,N_19654);
nand UO_1966 (O_1966,N_19556,N_19858);
nor UO_1967 (O_1967,N_19687,N_19768);
nor UO_1968 (O_1968,N_19524,N_19960);
nor UO_1969 (O_1969,N_19862,N_19547);
or UO_1970 (O_1970,N_19808,N_19888);
or UO_1971 (O_1971,N_19654,N_19903);
nand UO_1972 (O_1972,N_19838,N_19771);
nand UO_1973 (O_1973,N_19616,N_19972);
and UO_1974 (O_1974,N_19932,N_19828);
nand UO_1975 (O_1975,N_19625,N_19984);
nand UO_1976 (O_1976,N_19521,N_19800);
or UO_1977 (O_1977,N_19704,N_19940);
or UO_1978 (O_1978,N_19840,N_19554);
or UO_1979 (O_1979,N_19531,N_19769);
nor UO_1980 (O_1980,N_19582,N_19660);
nand UO_1981 (O_1981,N_19670,N_19512);
or UO_1982 (O_1982,N_19953,N_19768);
and UO_1983 (O_1983,N_19708,N_19515);
nand UO_1984 (O_1984,N_19660,N_19982);
and UO_1985 (O_1985,N_19542,N_19790);
or UO_1986 (O_1986,N_19735,N_19578);
nand UO_1987 (O_1987,N_19885,N_19759);
or UO_1988 (O_1988,N_19525,N_19970);
nor UO_1989 (O_1989,N_19724,N_19567);
nand UO_1990 (O_1990,N_19798,N_19742);
nand UO_1991 (O_1991,N_19836,N_19659);
nor UO_1992 (O_1992,N_19804,N_19835);
and UO_1993 (O_1993,N_19684,N_19628);
and UO_1994 (O_1994,N_19738,N_19646);
or UO_1995 (O_1995,N_19938,N_19633);
nand UO_1996 (O_1996,N_19904,N_19649);
nor UO_1997 (O_1997,N_19681,N_19627);
or UO_1998 (O_1998,N_19889,N_19885);
nor UO_1999 (O_1999,N_19514,N_19918);
nor UO_2000 (O_2000,N_19958,N_19659);
nor UO_2001 (O_2001,N_19718,N_19684);
nand UO_2002 (O_2002,N_19602,N_19630);
nor UO_2003 (O_2003,N_19730,N_19615);
and UO_2004 (O_2004,N_19657,N_19519);
or UO_2005 (O_2005,N_19837,N_19957);
nor UO_2006 (O_2006,N_19938,N_19998);
nor UO_2007 (O_2007,N_19731,N_19724);
xnor UO_2008 (O_2008,N_19964,N_19754);
and UO_2009 (O_2009,N_19840,N_19646);
nand UO_2010 (O_2010,N_19697,N_19666);
nand UO_2011 (O_2011,N_19743,N_19835);
or UO_2012 (O_2012,N_19791,N_19907);
or UO_2013 (O_2013,N_19958,N_19623);
nor UO_2014 (O_2014,N_19983,N_19502);
or UO_2015 (O_2015,N_19705,N_19635);
nor UO_2016 (O_2016,N_19706,N_19526);
and UO_2017 (O_2017,N_19812,N_19939);
xor UO_2018 (O_2018,N_19781,N_19847);
and UO_2019 (O_2019,N_19972,N_19954);
nand UO_2020 (O_2020,N_19858,N_19931);
or UO_2021 (O_2021,N_19986,N_19722);
nand UO_2022 (O_2022,N_19759,N_19692);
nand UO_2023 (O_2023,N_19652,N_19877);
or UO_2024 (O_2024,N_19541,N_19529);
nand UO_2025 (O_2025,N_19913,N_19528);
nand UO_2026 (O_2026,N_19883,N_19519);
nand UO_2027 (O_2027,N_19619,N_19635);
nand UO_2028 (O_2028,N_19677,N_19551);
nand UO_2029 (O_2029,N_19988,N_19702);
or UO_2030 (O_2030,N_19660,N_19636);
and UO_2031 (O_2031,N_19520,N_19680);
nand UO_2032 (O_2032,N_19980,N_19949);
or UO_2033 (O_2033,N_19767,N_19518);
and UO_2034 (O_2034,N_19803,N_19693);
or UO_2035 (O_2035,N_19998,N_19511);
nor UO_2036 (O_2036,N_19696,N_19840);
nor UO_2037 (O_2037,N_19805,N_19529);
nor UO_2038 (O_2038,N_19605,N_19800);
and UO_2039 (O_2039,N_19696,N_19958);
nor UO_2040 (O_2040,N_19714,N_19763);
or UO_2041 (O_2041,N_19581,N_19700);
nand UO_2042 (O_2042,N_19837,N_19976);
nand UO_2043 (O_2043,N_19582,N_19987);
or UO_2044 (O_2044,N_19733,N_19541);
or UO_2045 (O_2045,N_19679,N_19524);
nand UO_2046 (O_2046,N_19960,N_19936);
and UO_2047 (O_2047,N_19984,N_19712);
or UO_2048 (O_2048,N_19606,N_19693);
and UO_2049 (O_2049,N_19757,N_19822);
nand UO_2050 (O_2050,N_19723,N_19530);
nor UO_2051 (O_2051,N_19768,N_19732);
or UO_2052 (O_2052,N_19670,N_19528);
or UO_2053 (O_2053,N_19897,N_19517);
and UO_2054 (O_2054,N_19647,N_19578);
and UO_2055 (O_2055,N_19921,N_19764);
nor UO_2056 (O_2056,N_19931,N_19716);
and UO_2057 (O_2057,N_19629,N_19663);
nor UO_2058 (O_2058,N_19989,N_19848);
nor UO_2059 (O_2059,N_19749,N_19599);
nor UO_2060 (O_2060,N_19837,N_19953);
or UO_2061 (O_2061,N_19656,N_19817);
or UO_2062 (O_2062,N_19670,N_19574);
nand UO_2063 (O_2063,N_19791,N_19942);
and UO_2064 (O_2064,N_19574,N_19775);
and UO_2065 (O_2065,N_19720,N_19700);
and UO_2066 (O_2066,N_19856,N_19563);
nand UO_2067 (O_2067,N_19845,N_19502);
and UO_2068 (O_2068,N_19604,N_19938);
nor UO_2069 (O_2069,N_19995,N_19925);
or UO_2070 (O_2070,N_19943,N_19838);
nand UO_2071 (O_2071,N_19714,N_19608);
nor UO_2072 (O_2072,N_19532,N_19801);
nor UO_2073 (O_2073,N_19915,N_19534);
and UO_2074 (O_2074,N_19601,N_19981);
or UO_2075 (O_2075,N_19511,N_19698);
nand UO_2076 (O_2076,N_19898,N_19648);
and UO_2077 (O_2077,N_19772,N_19853);
and UO_2078 (O_2078,N_19573,N_19944);
nor UO_2079 (O_2079,N_19759,N_19802);
nor UO_2080 (O_2080,N_19905,N_19778);
and UO_2081 (O_2081,N_19595,N_19600);
or UO_2082 (O_2082,N_19727,N_19683);
nor UO_2083 (O_2083,N_19869,N_19954);
and UO_2084 (O_2084,N_19925,N_19605);
or UO_2085 (O_2085,N_19659,N_19556);
and UO_2086 (O_2086,N_19765,N_19903);
and UO_2087 (O_2087,N_19744,N_19831);
nand UO_2088 (O_2088,N_19955,N_19530);
and UO_2089 (O_2089,N_19716,N_19970);
nand UO_2090 (O_2090,N_19706,N_19502);
or UO_2091 (O_2091,N_19968,N_19587);
xnor UO_2092 (O_2092,N_19903,N_19831);
nor UO_2093 (O_2093,N_19517,N_19929);
xnor UO_2094 (O_2094,N_19899,N_19895);
nor UO_2095 (O_2095,N_19887,N_19736);
or UO_2096 (O_2096,N_19578,N_19911);
nand UO_2097 (O_2097,N_19640,N_19638);
and UO_2098 (O_2098,N_19703,N_19879);
or UO_2099 (O_2099,N_19765,N_19776);
and UO_2100 (O_2100,N_19651,N_19591);
nand UO_2101 (O_2101,N_19979,N_19997);
xor UO_2102 (O_2102,N_19737,N_19763);
and UO_2103 (O_2103,N_19976,N_19911);
nor UO_2104 (O_2104,N_19997,N_19714);
xnor UO_2105 (O_2105,N_19723,N_19897);
or UO_2106 (O_2106,N_19542,N_19583);
or UO_2107 (O_2107,N_19907,N_19643);
xor UO_2108 (O_2108,N_19720,N_19732);
nand UO_2109 (O_2109,N_19508,N_19886);
nor UO_2110 (O_2110,N_19882,N_19828);
xnor UO_2111 (O_2111,N_19556,N_19622);
nor UO_2112 (O_2112,N_19659,N_19888);
nand UO_2113 (O_2113,N_19807,N_19805);
nor UO_2114 (O_2114,N_19879,N_19830);
or UO_2115 (O_2115,N_19709,N_19750);
and UO_2116 (O_2116,N_19932,N_19904);
nor UO_2117 (O_2117,N_19820,N_19998);
nand UO_2118 (O_2118,N_19524,N_19680);
nand UO_2119 (O_2119,N_19644,N_19772);
nand UO_2120 (O_2120,N_19796,N_19969);
nor UO_2121 (O_2121,N_19587,N_19809);
nand UO_2122 (O_2122,N_19525,N_19905);
nor UO_2123 (O_2123,N_19815,N_19556);
and UO_2124 (O_2124,N_19574,N_19944);
nor UO_2125 (O_2125,N_19883,N_19685);
and UO_2126 (O_2126,N_19704,N_19988);
or UO_2127 (O_2127,N_19870,N_19644);
or UO_2128 (O_2128,N_19870,N_19620);
or UO_2129 (O_2129,N_19867,N_19551);
xnor UO_2130 (O_2130,N_19947,N_19523);
xor UO_2131 (O_2131,N_19957,N_19558);
nor UO_2132 (O_2132,N_19998,N_19749);
nand UO_2133 (O_2133,N_19627,N_19832);
or UO_2134 (O_2134,N_19694,N_19971);
or UO_2135 (O_2135,N_19545,N_19700);
or UO_2136 (O_2136,N_19566,N_19698);
nand UO_2137 (O_2137,N_19646,N_19607);
nand UO_2138 (O_2138,N_19900,N_19704);
nor UO_2139 (O_2139,N_19698,N_19921);
and UO_2140 (O_2140,N_19974,N_19890);
nand UO_2141 (O_2141,N_19779,N_19695);
nand UO_2142 (O_2142,N_19796,N_19555);
nand UO_2143 (O_2143,N_19653,N_19941);
nor UO_2144 (O_2144,N_19826,N_19586);
or UO_2145 (O_2145,N_19928,N_19821);
or UO_2146 (O_2146,N_19854,N_19720);
and UO_2147 (O_2147,N_19856,N_19623);
xnor UO_2148 (O_2148,N_19558,N_19733);
nand UO_2149 (O_2149,N_19537,N_19905);
nand UO_2150 (O_2150,N_19891,N_19932);
or UO_2151 (O_2151,N_19713,N_19677);
or UO_2152 (O_2152,N_19756,N_19704);
or UO_2153 (O_2153,N_19667,N_19749);
and UO_2154 (O_2154,N_19677,N_19837);
or UO_2155 (O_2155,N_19569,N_19797);
nor UO_2156 (O_2156,N_19935,N_19603);
and UO_2157 (O_2157,N_19879,N_19563);
nand UO_2158 (O_2158,N_19859,N_19869);
nor UO_2159 (O_2159,N_19553,N_19689);
nor UO_2160 (O_2160,N_19721,N_19954);
and UO_2161 (O_2161,N_19826,N_19548);
and UO_2162 (O_2162,N_19506,N_19749);
or UO_2163 (O_2163,N_19693,N_19808);
nand UO_2164 (O_2164,N_19987,N_19645);
nand UO_2165 (O_2165,N_19586,N_19815);
and UO_2166 (O_2166,N_19800,N_19602);
or UO_2167 (O_2167,N_19659,N_19530);
nand UO_2168 (O_2168,N_19699,N_19959);
and UO_2169 (O_2169,N_19663,N_19694);
or UO_2170 (O_2170,N_19519,N_19758);
nor UO_2171 (O_2171,N_19663,N_19542);
nand UO_2172 (O_2172,N_19991,N_19577);
xnor UO_2173 (O_2173,N_19538,N_19662);
or UO_2174 (O_2174,N_19848,N_19564);
and UO_2175 (O_2175,N_19919,N_19794);
and UO_2176 (O_2176,N_19738,N_19630);
nand UO_2177 (O_2177,N_19549,N_19980);
nor UO_2178 (O_2178,N_19905,N_19661);
nor UO_2179 (O_2179,N_19596,N_19722);
or UO_2180 (O_2180,N_19865,N_19502);
nand UO_2181 (O_2181,N_19574,N_19990);
xor UO_2182 (O_2182,N_19638,N_19973);
nand UO_2183 (O_2183,N_19677,N_19514);
or UO_2184 (O_2184,N_19745,N_19942);
and UO_2185 (O_2185,N_19935,N_19584);
or UO_2186 (O_2186,N_19724,N_19611);
nor UO_2187 (O_2187,N_19928,N_19582);
nand UO_2188 (O_2188,N_19830,N_19755);
or UO_2189 (O_2189,N_19886,N_19588);
or UO_2190 (O_2190,N_19648,N_19770);
or UO_2191 (O_2191,N_19528,N_19724);
nor UO_2192 (O_2192,N_19768,N_19507);
nand UO_2193 (O_2193,N_19991,N_19770);
nand UO_2194 (O_2194,N_19636,N_19991);
nand UO_2195 (O_2195,N_19524,N_19898);
or UO_2196 (O_2196,N_19684,N_19674);
nor UO_2197 (O_2197,N_19616,N_19872);
or UO_2198 (O_2198,N_19786,N_19523);
nand UO_2199 (O_2199,N_19679,N_19981);
and UO_2200 (O_2200,N_19730,N_19933);
or UO_2201 (O_2201,N_19939,N_19519);
nor UO_2202 (O_2202,N_19507,N_19573);
nor UO_2203 (O_2203,N_19760,N_19617);
nand UO_2204 (O_2204,N_19749,N_19888);
nand UO_2205 (O_2205,N_19610,N_19821);
nand UO_2206 (O_2206,N_19539,N_19650);
nand UO_2207 (O_2207,N_19942,N_19955);
and UO_2208 (O_2208,N_19841,N_19821);
nor UO_2209 (O_2209,N_19876,N_19620);
and UO_2210 (O_2210,N_19556,N_19848);
nand UO_2211 (O_2211,N_19823,N_19548);
and UO_2212 (O_2212,N_19792,N_19805);
nand UO_2213 (O_2213,N_19841,N_19584);
and UO_2214 (O_2214,N_19529,N_19750);
nand UO_2215 (O_2215,N_19868,N_19975);
and UO_2216 (O_2216,N_19517,N_19840);
or UO_2217 (O_2217,N_19707,N_19776);
and UO_2218 (O_2218,N_19526,N_19679);
and UO_2219 (O_2219,N_19673,N_19771);
nor UO_2220 (O_2220,N_19810,N_19738);
nor UO_2221 (O_2221,N_19965,N_19529);
xor UO_2222 (O_2222,N_19810,N_19989);
or UO_2223 (O_2223,N_19737,N_19553);
nor UO_2224 (O_2224,N_19713,N_19667);
and UO_2225 (O_2225,N_19841,N_19917);
nor UO_2226 (O_2226,N_19934,N_19737);
nand UO_2227 (O_2227,N_19559,N_19774);
and UO_2228 (O_2228,N_19786,N_19947);
or UO_2229 (O_2229,N_19948,N_19968);
nand UO_2230 (O_2230,N_19758,N_19986);
nor UO_2231 (O_2231,N_19794,N_19765);
nor UO_2232 (O_2232,N_19693,N_19914);
nand UO_2233 (O_2233,N_19579,N_19830);
and UO_2234 (O_2234,N_19603,N_19657);
and UO_2235 (O_2235,N_19559,N_19895);
and UO_2236 (O_2236,N_19506,N_19990);
nand UO_2237 (O_2237,N_19724,N_19714);
and UO_2238 (O_2238,N_19955,N_19825);
nor UO_2239 (O_2239,N_19738,N_19807);
or UO_2240 (O_2240,N_19503,N_19560);
or UO_2241 (O_2241,N_19667,N_19726);
and UO_2242 (O_2242,N_19772,N_19745);
or UO_2243 (O_2243,N_19530,N_19771);
or UO_2244 (O_2244,N_19897,N_19702);
nand UO_2245 (O_2245,N_19890,N_19975);
or UO_2246 (O_2246,N_19792,N_19594);
nand UO_2247 (O_2247,N_19880,N_19806);
nor UO_2248 (O_2248,N_19522,N_19614);
nor UO_2249 (O_2249,N_19621,N_19855);
or UO_2250 (O_2250,N_19960,N_19949);
nor UO_2251 (O_2251,N_19709,N_19623);
nand UO_2252 (O_2252,N_19595,N_19649);
nand UO_2253 (O_2253,N_19712,N_19550);
nand UO_2254 (O_2254,N_19538,N_19965);
nor UO_2255 (O_2255,N_19703,N_19714);
nand UO_2256 (O_2256,N_19578,N_19568);
nor UO_2257 (O_2257,N_19792,N_19895);
or UO_2258 (O_2258,N_19598,N_19973);
or UO_2259 (O_2259,N_19817,N_19595);
nand UO_2260 (O_2260,N_19808,N_19525);
and UO_2261 (O_2261,N_19723,N_19559);
or UO_2262 (O_2262,N_19950,N_19937);
and UO_2263 (O_2263,N_19854,N_19609);
nand UO_2264 (O_2264,N_19819,N_19680);
or UO_2265 (O_2265,N_19931,N_19937);
and UO_2266 (O_2266,N_19644,N_19580);
nand UO_2267 (O_2267,N_19927,N_19549);
nor UO_2268 (O_2268,N_19778,N_19523);
nand UO_2269 (O_2269,N_19736,N_19696);
or UO_2270 (O_2270,N_19827,N_19926);
or UO_2271 (O_2271,N_19560,N_19878);
and UO_2272 (O_2272,N_19625,N_19995);
or UO_2273 (O_2273,N_19575,N_19816);
nor UO_2274 (O_2274,N_19891,N_19590);
nand UO_2275 (O_2275,N_19549,N_19701);
or UO_2276 (O_2276,N_19694,N_19692);
and UO_2277 (O_2277,N_19809,N_19702);
nor UO_2278 (O_2278,N_19928,N_19647);
and UO_2279 (O_2279,N_19995,N_19746);
nand UO_2280 (O_2280,N_19951,N_19825);
or UO_2281 (O_2281,N_19620,N_19874);
or UO_2282 (O_2282,N_19640,N_19564);
or UO_2283 (O_2283,N_19736,N_19502);
nand UO_2284 (O_2284,N_19971,N_19640);
nand UO_2285 (O_2285,N_19987,N_19673);
and UO_2286 (O_2286,N_19876,N_19841);
and UO_2287 (O_2287,N_19575,N_19657);
or UO_2288 (O_2288,N_19806,N_19814);
nor UO_2289 (O_2289,N_19936,N_19715);
nor UO_2290 (O_2290,N_19674,N_19644);
or UO_2291 (O_2291,N_19729,N_19837);
nand UO_2292 (O_2292,N_19879,N_19877);
and UO_2293 (O_2293,N_19779,N_19560);
and UO_2294 (O_2294,N_19541,N_19669);
or UO_2295 (O_2295,N_19515,N_19642);
nand UO_2296 (O_2296,N_19748,N_19598);
and UO_2297 (O_2297,N_19889,N_19870);
and UO_2298 (O_2298,N_19853,N_19745);
nand UO_2299 (O_2299,N_19805,N_19824);
nor UO_2300 (O_2300,N_19852,N_19532);
or UO_2301 (O_2301,N_19751,N_19697);
and UO_2302 (O_2302,N_19583,N_19916);
or UO_2303 (O_2303,N_19733,N_19906);
and UO_2304 (O_2304,N_19760,N_19595);
or UO_2305 (O_2305,N_19590,N_19989);
nand UO_2306 (O_2306,N_19956,N_19930);
nor UO_2307 (O_2307,N_19528,N_19862);
or UO_2308 (O_2308,N_19578,N_19844);
or UO_2309 (O_2309,N_19992,N_19819);
and UO_2310 (O_2310,N_19748,N_19578);
or UO_2311 (O_2311,N_19550,N_19996);
or UO_2312 (O_2312,N_19616,N_19855);
and UO_2313 (O_2313,N_19591,N_19616);
and UO_2314 (O_2314,N_19501,N_19622);
nand UO_2315 (O_2315,N_19874,N_19603);
nand UO_2316 (O_2316,N_19560,N_19633);
nand UO_2317 (O_2317,N_19705,N_19507);
and UO_2318 (O_2318,N_19942,N_19779);
and UO_2319 (O_2319,N_19959,N_19969);
nor UO_2320 (O_2320,N_19817,N_19558);
or UO_2321 (O_2321,N_19789,N_19594);
or UO_2322 (O_2322,N_19652,N_19772);
nand UO_2323 (O_2323,N_19629,N_19749);
xor UO_2324 (O_2324,N_19685,N_19652);
nor UO_2325 (O_2325,N_19652,N_19898);
xor UO_2326 (O_2326,N_19782,N_19677);
or UO_2327 (O_2327,N_19668,N_19897);
nand UO_2328 (O_2328,N_19959,N_19788);
nand UO_2329 (O_2329,N_19713,N_19716);
nor UO_2330 (O_2330,N_19647,N_19512);
and UO_2331 (O_2331,N_19852,N_19927);
and UO_2332 (O_2332,N_19570,N_19837);
and UO_2333 (O_2333,N_19931,N_19687);
nor UO_2334 (O_2334,N_19526,N_19542);
nor UO_2335 (O_2335,N_19908,N_19784);
and UO_2336 (O_2336,N_19928,N_19528);
or UO_2337 (O_2337,N_19644,N_19948);
and UO_2338 (O_2338,N_19520,N_19560);
nor UO_2339 (O_2339,N_19585,N_19549);
and UO_2340 (O_2340,N_19573,N_19995);
and UO_2341 (O_2341,N_19583,N_19915);
nor UO_2342 (O_2342,N_19673,N_19791);
or UO_2343 (O_2343,N_19924,N_19987);
and UO_2344 (O_2344,N_19809,N_19579);
and UO_2345 (O_2345,N_19595,N_19745);
nor UO_2346 (O_2346,N_19645,N_19802);
and UO_2347 (O_2347,N_19516,N_19881);
and UO_2348 (O_2348,N_19724,N_19616);
and UO_2349 (O_2349,N_19714,N_19555);
or UO_2350 (O_2350,N_19725,N_19776);
nor UO_2351 (O_2351,N_19861,N_19988);
xnor UO_2352 (O_2352,N_19540,N_19544);
or UO_2353 (O_2353,N_19767,N_19729);
nor UO_2354 (O_2354,N_19908,N_19567);
or UO_2355 (O_2355,N_19897,N_19674);
nor UO_2356 (O_2356,N_19858,N_19876);
or UO_2357 (O_2357,N_19787,N_19898);
or UO_2358 (O_2358,N_19528,N_19674);
nand UO_2359 (O_2359,N_19668,N_19816);
or UO_2360 (O_2360,N_19585,N_19636);
or UO_2361 (O_2361,N_19833,N_19770);
and UO_2362 (O_2362,N_19731,N_19564);
and UO_2363 (O_2363,N_19642,N_19885);
nor UO_2364 (O_2364,N_19816,N_19716);
xor UO_2365 (O_2365,N_19976,N_19690);
nand UO_2366 (O_2366,N_19575,N_19562);
or UO_2367 (O_2367,N_19601,N_19684);
or UO_2368 (O_2368,N_19942,N_19971);
or UO_2369 (O_2369,N_19762,N_19984);
nor UO_2370 (O_2370,N_19931,N_19623);
nand UO_2371 (O_2371,N_19665,N_19814);
or UO_2372 (O_2372,N_19919,N_19832);
nand UO_2373 (O_2373,N_19612,N_19582);
nand UO_2374 (O_2374,N_19502,N_19563);
nand UO_2375 (O_2375,N_19685,N_19925);
nand UO_2376 (O_2376,N_19509,N_19625);
nand UO_2377 (O_2377,N_19899,N_19989);
and UO_2378 (O_2378,N_19853,N_19942);
and UO_2379 (O_2379,N_19815,N_19740);
nand UO_2380 (O_2380,N_19837,N_19853);
nor UO_2381 (O_2381,N_19591,N_19936);
nand UO_2382 (O_2382,N_19679,N_19582);
and UO_2383 (O_2383,N_19768,N_19739);
nor UO_2384 (O_2384,N_19830,N_19529);
nor UO_2385 (O_2385,N_19713,N_19891);
or UO_2386 (O_2386,N_19744,N_19593);
nand UO_2387 (O_2387,N_19911,N_19802);
nand UO_2388 (O_2388,N_19761,N_19966);
nor UO_2389 (O_2389,N_19536,N_19970);
nand UO_2390 (O_2390,N_19661,N_19687);
and UO_2391 (O_2391,N_19722,N_19918);
nand UO_2392 (O_2392,N_19869,N_19573);
nor UO_2393 (O_2393,N_19696,N_19959);
nand UO_2394 (O_2394,N_19686,N_19709);
nor UO_2395 (O_2395,N_19953,N_19897);
or UO_2396 (O_2396,N_19535,N_19553);
and UO_2397 (O_2397,N_19858,N_19581);
or UO_2398 (O_2398,N_19505,N_19644);
nand UO_2399 (O_2399,N_19705,N_19616);
nand UO_2400 (O_2400,N_19695,N_19761);
or UO_2401 (O_2401,N_19774,N_19593);
nand UO_2402 (O_2402,N_19746,N_19960);
nand UO_2403 (O_2403,N_19848,N_19776);
nor UO_2404 (O_2404,N_19925,N_19680);
and UO_2405 (O_2405,N_19917,N_19732);
nor UO_2406 (O_2406,N_19964,N_19713);
nor UO_2407 (O_2407,N_19562,N_19627);
nand UO_2408 (O_2408,N_19535,N_19869);
and UO_2409 (O_2409,N_19616,N_19868);
or UO_2410 (O_2410,N_19542,N_19666);
nand UO_2411 (O_2411,N_19667,N_19906);
and UO_2412 (O_2412,N_19760,N_19580);
nand UO_2413 (O_2413,N_19649,N_19613);
or UO_2414 (O_2414,N_19624,N_19904);
and UO_2415 (O_2415,N_19556,N_19889);
and UO_2416 (O_2416,N_19684,N_19591);
and UO_2417 (O_2417,N_19564,N_19752);
nand UO_2418 (O_2418,N_19987,N_19680);
and UO_2419 (O_2419,N_19818,N_19936);
nor UO_2420 (O_2420,N_19696,N_19893);
nor UO_2421 (O_2421,N_19781,N_19766);
and UO_2422 (O_2422,N_19515,N_19730);
nand UO_2423 (O_2423,N_19515,N_19908);
nor UO_2424 (O_2424,N_19857,N_19818);
nand UO_2425 (O_2425,N_19511,N_19561);
and UO_2426 (O_2426,N_19915,N_19818);
nand UO_2427 (O_2427,N_19752,N_19816);
nor UO_2428 (O_2428,N_19668,N_19527);
xnor UO_2429 (O_2429,N_19504,N_19998);
and UO_2430 (O_2430,N_19847,N_19734);
or UO_2431 (O_2431,N_19870,N_19561);
or UO_2432 (O_2432,N_19565,N_19950);
nand UO_2433 (O_2433,N_19877,N_19669);
nand UO_2434 (O_2434,N_19810,N_19538);
or UO_2435 (O_2435,N_19770,N_19964);
nor UO_2436 (O_2436,N_19654,N_19586);
and UO_2437 (O_2437,N_19572,N_19938);
nand UO_2438 (O_2438,N_19960,N_19836);
nand UO_2439 (O_2439,N_19765,N_19691);
nor UO_2440 (O_2440,N_19655,N_19603);
or UO_2441 (O_2441,N_19571,N_19504);
and UO_2442 (O_2442,N_19518,N_19610);
or UO_2443 (O_2443,N_19826,N_19904);
or UO_2444 (O_2444,N_19522,N_19510);
and UO_2445 (O_2445,N_19617,N_19627);
nor UO_2446 (O_2446,N_19967,N_19797);
and UO_2447 (O_2447,N_19644,N_19751);
nor UO_2448 (O_2448,N_19644,N_19957);
nand UO_2449 (O_2449,N_19521,N_19690);
nor UO_2450 (O_2450,N_19947,N_19658);
nand UO_2451 (O_2451,N_19873,N_19513);
nor UO_2452 (O_2452,N_19860,N_19895);
and UO_2453 (O_2453,N_19516,N_19812);
or UO_2454 (O_2454,N_19944,N_19673);
nor UO_2455 (O_2455,N_19587,N_19858);
or UO_2456 (O_2456,N_19738,N_19869);
nand UO_2457 (O_2457,N_19892,N_19725);
nand UO_2458 (O_2458,N_19613,N_19740);
or UO_2459 (O_2459,N_19792,N_19755);
nor UO_2460 (O_2460,N_19689,N_19802);
and UO_2461 (O_2461,N_19578,N_19622);
nor UO_2462 (O_2462,N_19533,N_19552);
nor UO_2463 (O_2463,N_19559,N_19824);
or UO_2464 (O_2464,N_19930,N_19826);
and UO_2465 (O_2465,N_19834,N_19611);
nor UO_2466 (O_2466,N_19755,N_19601);
nand UO_2467 (O_2467,N_19518,N_19719);
nand UO_2468 (O_2468,N_19720,N_19754);
nor UO_2469 (O_2469,N_19508,N_19939);
nand UO_2470 (O_2470,N_19530,N_19525);
nand UO_2471 (O_2471,N_19742,N_19528);
and UO_2472 (O_2472,N_19581,N_19950);
and UO_2473 (O_2473,N_19849,N_19599);
and UO_2474 (O_2474,N_19652,N_19669);
or UO_2475 (O_2475,N_19519,N_19700);
nand UO_2476 (O_2476,N_19539,N_19948);
and UO_2477 (O_2477,N_19880,N_19906);
or UO_2478 (O_2478,N_19795,N_19585);
nand UO_2479 (O_2479,N_19902,N_19599);
nand UO_2480 (O_2480,N_19624,N_19539);
nand UO_2481 (O_2481,N_19656,N_19882);
nand UO_2482 (O_2482,N_19552,N_19575);
nor UO_2483 (O_2483,N_19572,N_19594);
and UO_2484 (O_2484,N_19805,N_19797);
or UO_2485 (O_2485,N_19823,N_19595);
or UO_2486 (O_2486,N_19800,N_19644);
and UO_2487 (O_2487,N_19880,N_19927);
nand UO_2488 (O_2488,N_19645,N_19847);
and UO_2489 (O_2489,N_19937,N_19996);
nor UO_2490 (O_2490,N_19854,N_19709);
and UO_2491 (O_2491,N_19522,N_19600);
nor UO_2492 (O_2492,N_19710,N_19972);
or UO_2493 (O_2493,N_19645,N_19679);
or UO_2494 (O_2494,N_19827,N_19951);
xor UO_2495 (O_2495,N_19706,N_19695);
nor UO_2496 (O_2496,N_19541,N_19935);
nand UO_2497 (O_2497,N_19753,N_19764);
nor UO_2498 (O_2498,N_19924,N_19869);
or UO_2499 (O_2499,N_19894,N_19665);
endmodule