module basic_3000_30000_3500_100_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_1875,In_860);
and U1 (N_1,In_2258,In_1371);
nor U2 (N_2,In_2370,In_1242);
nor U3 (N_3,In_64,In_577);
nand U4 (N_4,In_1800,In_2894);
nor U5 (N_5,In_1446,In_2244);
or U6 (N_6,In_1085,In_2467);
or U7 (N_7,In_2914,In_2193);
nor U8 (N_8,In_1305,In_316);
and U9 (N_9,In_2725,In_230);
xnor U10 (N_10,In_2334,In_932);
or U11 (N_11,In_826,In_720);
or U12 (N_12,In_2132,In_1577);
nand U13 (N_13,In_1665,In_540);
nand U14 (N_14,In_1496,In_806);
or U15 (N_15,In_2508,In_2947);
or U16 (N_16,In_2367,In_2336);
nand U17 (N_17,In_2602,In_466);
or U18 (N_18,In_2918,In_1428);
nand U19 (N_19,In_2450,In_1781);
and U20 (N_20,In_382,In_2466);
xor U21 (N_21,In_1862,In_2391);
and U22 (N_22,In_1080,In_752);
nand U23 (N_23,In_239,In_2523);
or U24 (N_24,In_134,In_521);
nand U25 (N_25,In_2591,In_642);
nor U26 (N_26,In_2317,In_2231);
or U27 (N_27,In_1547,In_1576);
and U28 (N_28,In_2384,In_449);
nand U29 (N_29,In_2506,In_1290);
xor U30 (N_30,In_2026,In_1895);
xnor U31 (N_31,In_2489,In_2011);
or U32 (N_32,In_2456,In_200);
or U33 (N_33,In_1565,In_1769);
or U34 (N_34,In_266,In_1350);
nor U35 (N_35,In_1937,In_2048);
and U36 (N_36,In_131,In_2409);
nor U37 (N_37,In_2668,In_46);
and U38 (N_38,In_690,In_640);
xnor U39 (N_39,In_2779,In_572);
and U40 (N_40,In_498,In_499);
xnor U41 (N_41,In_324,In_1135);
nand U42 (N_42,In_997,In_581);
xor U43 (N_43,In_2598,In_805);
or U44 (N_44,In_2388,In_2975);
nor U45 (N_45,In_280,In_42);
nand U46 (N_46,In_579,In_2039);
or U47 (N_47,In_1345,In_2123);
xnor U48 (N_48,In_2962,In_950);
xor U49 (N_49,In_2061,In_1266);
xor U50 (N_50,In_842,In_320);
nand U51 (N_51,In_2178,In_592);
nor U52 (N_52,In_1819,In_1293);
nand U53 (N_53,In_2457,In_2646);
and U54 (N_54,In_1891,In_162);
nand U55 (N_55,In_881,In_2511);
nor U56 (N_56,In_969,In_991);
nor U57 (N_57,In_1997,In_768);
and U58 (N_58,In_686,In_2066);
or U59 (N_59,In_666,In_451);
and U60 (N_60,In_1578,In_1921);
or U61 (N_61,In_2690,In_1210);
nand U62 (N_62,In_1200,In_2618);
nand U63 (N_63,In_2912,In_1562);
or U64 (N_64,In_1698,In_861);
nor U65 (N_65,In_1880,In_1344);
and U66 (N_66,In_2593,In_2895);
xor U67 (N_67,In_1431,In_1391);
and U68 (N_68,In_2143,In_2605);
nand U69 (N_69,In_2509,In_2294);
xnor U70 (N_70,In_1035,In_1464);
nor U71 (N_71,In_786,In_2485);
nor U72 (N_72,In_1491,In_2741);
xor U73 (N_73,In_1814,In_2966);
xor U74 (N_74,In_458,In_776);
or U75 (N_75,In_2746,In_623);
or U76 (N_76,In_2371,In_2562);
xnor U77 (N_77,In_1870,In_485);
nor U78 (N_78,In_1911,In_393);
nand U79 (N_79,In_664,In_2539);
and U80 (N_80,In_2328,In_2880);
xor U81 (N_81,In_1883,In_2907);
or U82 (N_82,In_2337,In_1955);
and U83 (N_83,In_2643,In_2145);
nor U84 (N_84,In_440,In_441);
and U85 (N_85,In_680,In_377);
or U86 (N_86,In_1585,In_2869);
and U87 (N_87,In_2327,In_246);
and U88 (N_88,In_1207,In_1936);
xnor U89 (N_89,In_1269,In_2475);
xnor U90 (N_90,In_2465,In_1501);
or U91 (N_91,In_2196,In_259);
nor U92 (N_92,In_1668,In_1091);
nor U93 (N_93,In_346,In_1700);
nand U94 (N_94,In_2846,In_2096);
nand U95 (N_95,In_2799,In_2205);
and U96 (N_96,In_1587,In_1477);
or U97 (N_97,In_1904,In_1012);
xor U98 (N_98,In_1555,In_1570);
or U99 (N_99,In_2028,In_272);
nand U100 (N_100,In_1897,In_1497);
or U101 (N_101,In_240,In_2341);
and U102 (N_102,In_2872,In_130);
nor U103 (N_103,In_1796,In_439);
or U104 (N_104,In_819,In_107);
and U105 (N_105,In_282,In_670);
nand U106 (N_106,In_1368,In_2683);
and U107 (N_107,In_1826,In_29);
or U108 (N_108,In_2012,In_2524);
and U109 (N_109,In_65,In_502);
nor U110 (N_110,In_658,In_1910);
nor U111 (N_111,In_1486,In_764);
nand U112 (N_112,In_934,In_2261);
nor U113 (N_113,In_2599,In_2108);
xnor U114 (N_114,In_1600,In_1941);
or U115 (N_115,In_1945,In_2971);
nand U116 (N_116,In_467,In_1327);
or U117 (N_117,In_305,In_2778);
or U118 (N_118,In_948,In_2463);
nand U119 (N_119,In_2688,In_1334);
or U120 (N_120,In_311,In_2249);
xnor U121 (N_121,In_2442,In_1201);
or U122 (N_122,In_68,In_2674);
or U123 (N_123,In_2394,In_613);
nor U124 (N_124,In_2978,In_1525);
nor U125 (N_125,In_2216,In_1098);
or U126 (N_126,In_2252,In_344);
nor U127 (N_127,In_1901,In_2941);
nand U128 (N_128,In_545,In_1443);
nand U129 (N_129,In_2322,In_2641);
nor U130 (N_130,In_1573,In_2232);
and U131 (N_131,In_2279,In_494);
nand U132 (N_132,In_49,In_977);
xnor U133 (N_133,In_2512,In_1773);
or U134 (N_134,In_2520,In_2136);
and U135 (N_135,In_2316,In_1251);
nand U136 (N_136,In_337,In_2927);
xor U137 (N_137,In_1337,In_937);
nand U138 (N_138,In_303,In_2424);
nand U139 (N_139,In_1332,In_1149);
nor U140 (N_140,In_2002,In_2118);
and U141 (N_141,In_2365,In_1124);
nor U142 (N_142,In_2762,In_892);
and U143 (N_143,In_733,In_2528);
nand U144 (N_144,In_392,In_1173);
or U145 (N_145,In_2493,In_527);
nand U146 (N_146,In_957,In_2732);
nor U147 (N_147,In_2204,In_2537);
xor U148 (N_148,In_812,In_1718);
and U149 (N_149,In_2560,In_2590);
or U150 (N_150,In_22,In_2967);
and U151 (N_151,In_1393,In_1390);
nor U152 (N_152,In_2949,In_2468);
or U153 (N_153,In_1185,In_2472);
or U154 (N_154,In_517,In_886);
nor U155 (N_155,In_1719,In_2168);
nand U156 (N_156,In_799,In_2154);
nand U157 (N_157,In_1946,In_2780);
xnor U158 (N_158,In_359,In_2400);
xor U159 (N_159,In_1320,In_1836);
or U160 (N_160,In_358,In_2961);
nand U161 (N_161,In_1925,In_1864);
nand U162 (N_162,In_1268,In_253);
nor U163 (N_163,In_227,In_1508);
or U164 (N_164,In_194,In_2661);
xnor U165 (N_165,In_857,In_372);
nand U166 (N_166,In_852,In_1657);
and U167 (N_167,In_1061,In_2733);
nor U168 (N_168,In_557,In_2504);
and U169 (N_169,In_427,In_2818);
nor U170 (N_170,In_2936,In_1247);
and U171 (N_171,In_2901,In_2785);
nand U172 (N_172,In_772,In_2478);
xor U173 (N_173,In_1140,In_2530);
nor U174 (N_174,In_2151,In_1510);
nor U175 (N_175,In_556,In_612);
nor U176 (N_176,In_1026,In_181);
nand U177 (N_177,In_2025,In_855);
xor U178 (N_178,In_1952,In_168);
nor U179 (N_179,In_1615,In_2019);
or U180 (N_180,In_1662,In_1152);
or U181 (N_181,In_941,In_1704);
nor U182 (N_182,In_1723,In_1004);
nor U183 (N_183,In_769,In_638);
nor U184 (N_184,In_1916,In_1358);
nand U185 (N_185,In_2979,In_1063);
or U186 (N_186,In_483,In_1228);
and U187 (N_187,In_2623,In_357);
or U188 (N_188,In_2666,In_900);
and U189 (N_189,In_851,In_205);
and U190 (N_190,In_126,In_2042);
nand U191 (N_191,In_2223,In_402);
nor U192 (N_192,In_2859,In_2285);
nor U193 (N_193,In_2345,In_2831);
nor U194 (N_194,In_120,In_1130);
and U195 (N_195,In_2808,In_1889);
xnor U196 (N_196,In_1859,In_1301);
and U197 (N_197,In_164,In_224);
nor U198 (N_198,In_428,In_476);
or U199 (N_199,In_574,In_1123);
and U200 (N_200,In_1892,In_1328);
and U201 (N_201,In_870,In_2325);
xor U202 (N_202,In_637,In_1583);
nand U203 (N_203,In_2611,In_1404);
nand U204 (N_204,In_8,In_229);
xnor U205 (N_205,In_2813,In_1774);
nor U206 (N_206,In_1351,In_1436);
nor U207 (N_207,In_2738,In_2995);
xor U208 (N_208,In_73,In_871);
nand U209 (N_209,In_814,In_982);
or U210 (N_210,In_1473,In_460);
nor U211 (N_211,In_1867,In_1265);
or U212 (N_212,In_2302,In_1482);
nor U213 (N_213,In_2844,In_1956);
and U214 (N_214,In_910,In_1579);
nand U215 (N_215,In_509,In_55);
and U216 (N_216,In_180,In_2101);
and U217 (N_217,In_2046,In_185);
and U218 (N_218,In_949,In_1561);
or U219 (N_219,In_1273,In_2597);
nor U220 (N_220,In_2853,In_1281);
and U221 (N_221,In_511,In_1352);
and U222 (N_222,In_2210,In_946);
and U223 (N_223,In_1229,In_1416);
xnor U224 (N_224,In_1392,In_1693);
nor U225 (N_225,In_1324,In_2516);
nand U226 (N_226,In_1394,In_2787);
and U227 (N_227,In_1630,In_2273);
nand U228 (N_228,In_2527,In_844);
or U229 (N_229,In_2405,In_1089);
nand U230 (N_230,In_2320,In_154);
and U231 (N_231,In_782,In_2037);
xor U232 (N_232,In_1746,In_371);
nand U233 (N_233,In_504,In_464);
and U234 (N_234,In_966,In_2270);
nand U235 (N_235,In_1049,In_2968);
nand U236 (N_236,In_986,In_115);
or U237 (N_237,In_1567,In_2129);
nor U238 (N_238,In_905,In_939);
nand U239 (N_239,In_1346,In_2801);
and U240 (N_240,In_1364,In_2536);
and U241 (N_241,In_1882,In_2404);
nand U242 (N_242,In_1742,In_2563);
nor U243 (N_243,In_813,In_487);
xnor U244 (N_244,In_2669,In_47);
nor U245 (N_245,In_2705,In_1975);
xnor U246 (N_246,In_1258,In_268);
nor U247 (N_247,In_1223,In_285);
or U248 (N_248,In_790,In_146);
or U249 (N_249,In_437,In_13);
and U250 (N_250,In_1823,In_1526);
nor U251 (N_251,In_1214,In_1276);
and U252 (N_252,In_1489,In_193);
nand U253 (N_253,In_2575,In_2679);
or U254 (N_254,In_705,In_532);
and U255 (N_255,In_1254,In_473);
and U256 (N_256,In_2559,In_2542);
or U257 (N_257,In_2960,In_2934);
or U258 (N_258,In_1740,In_1453);
nand U259 (N_259,In_2974,In_406);
nand U260 (N_260,In_762,In_1658);
xnor U261 (N_261,In_2849,In_698);
xor U262 (N_262,In_656,In_2021);
xor U263 (N_263,In_2697,In_2374);
or U264 (N_264,In_1913,In_215);
or U265 (N_265,In_2079,In_2877);
and U266 (N_266,In_2418,In_1602);
nor U267 (N_267,In_1167,In_1705);
or U268 (N_268,In_2209,In_2295);
xnor U269 (N_269,In_114,In_2868);
and U270 (N_270,In_1537,In_231);
and U271 (N_271,In_2141,In_644);
nor U272 (N_272,In_2237,In_385);
and U273 (N_273,In_195,In_548);
xnor U274 (N_274,In_70,In_1843);
nand U275 (N_275,In_1783,In_2546);
or U276 (N_276,In_1888,In_763);
and U277 (N_277,In_1960,In_2517);
nand U278 (N_278,In_2604,In_2900);
or U279 (N_279,In_1631,In_2634);
nor U280 (N_280,In_40,In_866);
nand U281 (N_281,In_167,In_2375);
or U282 (N_282,In_1447,In_105);
and U283 (N_283,In_933,In_2488);
and U284 (N_284,In_155,In_2554);
and U285 (N_285,In_56,In_2988);
nand U286 (N_286,In_766,In_235);
xnor U287 (N_287,In_2689,In_1241);
xor U288 (N_288,In_1260,In_961);
nand U289 (N_289,In_2099,In_2724);
nor U290 (N_290,In_2981,In_1974);
xor U291 (N_291,In_2191,In_2699);
or U292 (N_292,In_331,In_1772);
xnor U293 (N_293,In_1756,In_2293);
nor U294 (N_294,In_955,In_2749);
nor U295 (N_295,In_2329,In_2942);
nand U296 (N_296,In_523,In_1995);
xor U297 (N_297,In_1831,In_2126);
nand U298 (N_298,In_1230,In_480);
nor U299 (N_299,In_1126,In_2581);
nand U300 (N_300,In_2878,In_1192);
and U301 (N_301,In_2612,In_108);
nand U302 (N_302,N_109,In_928);
xor U303 (N_303,In_1060,In_2825);
xnor U304 (N_304,In_2832,In_1655);
xnor U305 (N_305,In_2086,In_1499);
nor U306 (N_306,N_259,In_308);
nor U307 (N_307,In_1425,In_1855);
xnor U308 (N_308,In_1161,In_2432);
or U309 (N_309,In_2522,In_1440);
nand U310 (N_310,In_10,In_823);
or U311 (N_311,In_1986,In_1580);
and U312 (N_312,In_26,In_1847);
nand U313 (N_313,In_536,In_784);
nor U314 (N_314,In_1808,In_2201);
or U315 (N_315,In_1953,In_32);
and U316 (N_316,In_1,In_226);
xnor U317 (N_317,In_864,In_2502);
or U318 (N_318,In_1038,In_1967);
and U319 (N_319,In_2430,In_2969);
nand U320 (N_320,In_2071,In_2410);
nand U321 (N_321,In_2954,In_1374);
or U322 (N_322,In_2284,In_1732);
nor U323 (N_323,In_919,In_2972);
nand U324 (N_324,In_952,In_2567);
xnor U325 (N_325,In_1617,In_1353);
xnor U326 (N_326,In_828,In_514);
or U327 (N_327,In_152,In_1551);
and U328 (N_328,In_2529,In_1777);
or U329 (N_329,In_1158,In_2212);
nor U330 (N_330,In_833,N_224);
nor U331 (N_331,In_551,In_2416);
nand U332 (N_332,In_2095,In_2251);
and U333 (N_333,N_245,In_599);
nor U334 (N_334,In_2338,In_2033);
xor U335 (N_335,In_51,In_1779);
nand U336 (N_336,In_1935,In_2695);
or U337 (N_337,In_204,In_921);
or U338 (N_338,In_158,In_2871);
xnor U339 (N_339,In_2739,In_2897);
or U340 (N_340,In_1377,N_59);
nor U341 (N_341,In_2845,In_1382);
and U342 (N_342,In_796,In_113);
xnor U343 (N_343,In_667,In_522);
or U344 (N_344,In_1183,In_2617);
and U345 (N_345,In_50,In_2481);
nand U346 (N_346,N_61,N_103);
and U347 (N_347,In_893,In_2881);
nand U348 (N_348,N_12,N_4);
nand U349 (N_349,In_1156,In_1412);
and U350 (N_350,In_212,In_2800);
nor U351 (N_351,In_2189,N_145);
and U352 (N_352,In_1817,In_877);
or U353 (N_353,In_503,In_1025);
xnor U354 (N_354,In_1461,In_1488);
nand U355 (N_355,In_1726,In_156);
or U356 (N_356,In_742,N_64);
or U357 (N_357,In_386,In_1994);
nand U358 (N_358,In_317,In_2497);
or U359 (N_359,In_199,In_1076);
and U360 (N_360,In_2991,In_2133);
xnor U361 (N_361,In_2862,In_1144);
and U362 (N_362,In_211,In_2519);
or U363 (N_363,N_231,In_53);
nor U364 (N_364,In_707,In_2161);
xnor U365 (N_365,In_1262,In_2913);
and U366 (N_366,In_795,In_1900);
xnor U367 (N_367,In_179,In_1786);
nand U368 (N_368,In_261,In_1968);
xor U369 (N_369,In_1236,In_2176);
nor U370 (N_370,In_1839,In_1816);
xnor U371 (N_371,In_767,N_65);
xor U372 (N_372,In_618,In_54);
and U373 (N_373,In_2063,In_2218);
xor U374 (N_374,In_315,In_2097);
and U375 (N_375,In_2834,In_571);
and U376 (N_376,In_515,In_2272);
and U377 (N_377,In_434,In_963);
or U378 (N_378,In_1078,In_2483);
or U379 (N_379,In_2946,In_868);
and U380 (N_380,In_301,In_622);
nand U381 (N_381,In_2436,In_1159);
nor U382 (N_382,In_1217,In_1625);
xnor U383 (N_383,In_2181,In_2993);
and U384 (N_384,In_2268,In_2074);
and U385 (N_385,In_2632,N_97);
or U386 (N_386,In_479,In_628);
xor U387 (N_387,In_1679,In_2750);
and U388 (N_388,In_1102,In_147);
nor U389 (N_389,In_2510,N_123);
nor U390 (N_390,N_113,In_2073);
or U391 (N_391,In_1743,In_2970);
nand U392 (N_392,In_455,In_474);
xor U393 (N_393,In_926,In_174);
and U394 (N_394,N_13,In_2501);
nor U395 (N_395,In_2582,In_183);
xnor U396 (N_396,In_1639,In_968);
nor U397 (N_397,In_94,In_1589);
nor U398 (N_398,In_1445,In_1065);
and U399 (N_399,In_1611,In_1557);
and U400 (N_400,N_199,In_2356);
or U401 (N_401,In_1829,In_1691);
and U402 (N_402,In_2239,In_602);
xor U403 (N_403,In_1692,In_1370);
xnor U404 (N_404,In_1950,In_2162);
or U405 (N_405,In_2751,In_1275);
nand U406 (N_406,In_1502,In_150);
xnor U407 (N_407,N_56,In_388);
nor U408 (N_408,In_2435,In_366);
xnor U409 (N_409,In_2446,N_229);
or U410 (N_410,In_188,In_1329);
nor U411 (N_411,In_1225,N_20);
and U412 (N_412,In_1789,In_1457);
or U413 (N_413,N_158,N_216);
nand U414 (N_414,In_739,In_500);
or U415 (N_415,In_535,In_74);
xor U416 (N_416,In_850,In_141);
xnor U417 (N_417,In_334,N_112);
xor U418 (N_418,In_1634,In_2735);
or U419 (N_419,In_2874,In_1234);
nand U420 (N_420,In_289,In_1448);
xnor U421 (N_421,In_1681,In_1079);
nor U422 (N_422,In_379,In_2297);
or U423 (N_423,In_560,In_1044);
xor U424 (N_424,In_1381,In_1113);
or U425 (N_425,In_2809,In_2112);
and U426 (N_426,In_2875,In_2155);
nand U427 (N_427,In_1768,In_2087);
nand U428 (N_428,In_1930,In_1070);
nand U429 (N_429,In_1531,In_1702);
nor U430 (N_430,N_240,In_484);
nand U431 (N_431,In_2438,In_23);
or U432 (N_432,In_575,In_875);
nor U433 (N_433,In_1965,In_723);
nor U434 (N_434,In_216,In_726);
nand U435 (N_435,In_2761,In_2928);
or U436 (N_436,In_1683,In_2023);
and U437 (N_437,In_2248,In_2072);
nor U438 (N_438,N_186,In_187);
and U439 (N_439,In_1552,In_2429);
nor U440 (N_440,In_890,In_1354);
nand U441 (N_441,In_273,In_652);
or U442 (N_442,In_1176,In_2022);
or U443 (N_443,In_1199,N_57);
and U444 (N_444,In_990,In_853);
nor U445 (N_445,In_271,N_225);
nor U446 (N_446,N_134,N_191);
nor U447 (N_447,In_489,In_537);
nor U448 (N_448,In_2908,In_2412);
nand U449 (N_449,In_1543,In_1030);
nor U450 (N_450,In_2004,In_591);
and U451 (N_451,In_2083,In_1310);
xnor U452 (N_452,In_944,In_1541);
xor U453 (N_453,N_91,In_620);
and U454 (N_454,In_376,In_2125);
xnor U455 (N_455,In_2107,In_2029);
and U456 (N_456,In_2199,In_2100);
or U457 (N_457,In_2377,In_2982);
nor U458 (N_458,In_725,In_433);
nand U459 (N_459,In_2745,In_914);
nand U460 (N_460,In_1338,In_953);
or U461 (N_461,In_1856,In_1666);
nor U462 (N_462,In_576,In_1643);
and U463 (N_463,In_192,In_2243);
or U464 (N_464,N_133,In_197);
nor U465 (N_465,N_162,In_1278);
or U466 (N_466,In_2333,In_267);
and U467 (N_467,In_2228,In_2943);
xnor U468 (N_468,In_1898,In_2860);
or U469 (N_469,In_482,In_0);
nor U470 (N_470,In_2380,N_181);
nor U471 (N_471,In_911,In_1471);
or U472 (N_472,In_1421,In_2775);
nor U473 (N_473,In_879,In_1942);
nor U474 (N_474,In_1021,In_2389);
and U475 (N_475,In_347,N_275);
nand U476 (N_476,N_246,In_876);
xor U477 (N_477,In_1010,In_958);
nor U478 (N_478,In_874,In_631);
nand U479 (N_479,In_2676,In_738);
xnor U480 (N_480,In_2130,In_2451);
nand U481 (N_481,In_2959,In_843);
xor U482 (N_482,N_135,In_2001);
and U483 (N_483,In_327,In_309);
nor U484 (N_484,In_728,In_2142);
nand U485 (N_485,In_438,In_711);
nor U486 (N_486,In_1333,In_2588);
nand U487 (N_487,In_75,In_2889);
nand U488 (N_488,N_171,In_552);
nand U489 (N_489,In_1710,In_2360);
or U490 (N_490,In_1735,In_1006);
and U491 (N_491,In_2180,In_1194);
or U492 (N_492,In_2464,In_3);
xnor U493 (N_493,In_1738,In_880);
nand U494 (N_494,In_1188,In_2771);
nand U495 (N_495,In_816,In_2188);
nand U496 (N_496,In_1476,In_4);
nor U497 (N_497,In_959,In_1429);
nand U498 (N_498,In_291,In_744);
xor U499 (N_499,In_1616,N_60);
nor U500 (N_500,In_2712,In_2372);
nand U501 (N_501,In_634,In_2213);
and U502 (N_502,In_821,In_1401);
nor U503 (N_503,In_646,In_2447);
nor U504 (N_504,In_998,In_153);
and U505 (N_505,In_2525,In_854);
and U506 (N_506,In_516,In_299);
or U507 (N_507,In_2565,In_409);
nand U508 (N_508,In_2923,N_284);
nor U509 (N_509,In_1684,In_368);
xnor U510 (N_510,In_1951,In_1253);
nor U511 (N_511,In_1564,In_2702);
xor U512 (N_512,N_152,N_42);
xnor U513 (N_513,In_2549,N_77);
nor U514 (N_514,In_1650,In_2376);
xnor U515 (N_515,In_1599,In_935);
and U516 (N_516,In_668,In_1127);
and U517 (N_517,In_1081,In_2027);
and U518 (N_518,In_462,In_2230);
nand U519 (N_519,In_595,In_1717);
nand U520 (N_520,In_1107,In_989);
xnor U521 (N_521,In_2090,In_2802);
nor U522 (N_522,In_381,In_1481);
and U523 (N_523,In_2177,In_729);
nor U524 (N_524,In_354,In_1043);
xnor U525 (N_525,In_2064,In_43);
nand U526 (N_526,In_247,In_415);
and U527 (N_527,N_126,In_1964);
nand U528 (N_528,In_2402,In_306);
nor U529 (N_529,In_1538,In_887);
nand U530 (N_530,In_1733,In_793);
or U531 (N_531,In_2113,In_2558);
nand U532 (N_532,In_475,N_172);
or U533 (N_533,In_2514,In_558);
nand U534 (N_534,In_1097,N_148);
nand U535 (N_535,In_411,In_374);
or U536 (N_536,In_39,N_235);
or U537 (N_537,In_297,N_67);
and U538 (N_538,In_1820,N_89);
nor U539 (N_539,In_1170,In_1944);
nor U540 (N_540,In_2227,In_994);
nor U541 (N_541,In_1046,In_9);
and U542 (N_542,In_28,In_2765);
nor U543 (N_543,In_2434,In_132);
nor U544 (N_544,In_2773,In_1857);
or U545 (N_545,In_1271,In_2584);
xor U546 (N_546,In_836,In_2851);
nand U547 (N_547,In_2837,In_730);
and U548 (N_548,In_2036,In_1782);
and U549 (N_549,In_1558,In_1584);
or U550 (N_550,N_280,In_2873);
xnor U551 (N_551,In_2202,In_2940);
and U552 (N_552,In_2964,In_2983);
nand U553 (N_553,In_1179,In_2401);
and U554 (N_554,In_121,In_2693);
or U555 (N_555,N_46,In_1315);
xor U556 (N_556,N_272,In_1760);
and U557 (N_557,In_1569,In_2764);
or U558 (N_558,In_1292,In_846);
xnor U559 (N_559,In_2006,In_2459);
and U560 (N_560,In_390,In_48);
nor U561 (N_561,In_2980,In_1145);
nor U562 (N_562,In_2552,In_1540);
nor U563 (N_563,In_1629,In_672);
xor U564 (N_564,In_746,In_1850);
or U565 (N_565,In_222,In_116);
and U566 (N_566,In_217,In_993);
nor U567 (N_567,N_267,N_63);
nand U568 (N_568,In_1095,In_2956);
nor U569 (N_569,In_984,In_1514);
nor U570 (N_570,In_678,In_1915);
or U571 (N_571,In_2276,In_2636);
or U572 (N_572,In_747,In_2572);
and U573 (N_573,In_2743,In_1770);
and U574 (N_574,In_648,In_1178);
nand U575 (N_575,In_243,In_2156);
and U576 (N_576,In_2052,In_2867);
and U577 (N_577,In_1110,In_779);
nand U578 (N_578,In_559,In_1545);
and U579 (N_579,In_2596,In_248);
xor U580 (N_580,In_1191,In_908);
or U581 (N_581,In_2452,In_260);
xor U582 (N_582,In_2480,In_569);
or U583 (N_583,In_352,In_1678);
or U584 (N_584,In_639,In_103);
or U585 (N_585,In_2321,In_2672);
nand U586 (N_586,In_2009,In_2620);
and U587 (N_587,In_25,N_3);
nor U588 (N_588,In_1610,In_609);
xor U589 (N_589,In_251,In_2044);
nor U590 (N_590,N_220,In_1886);
xor U591 (N_591,In_149,In_2242);
or U592 (N_592,N_175,In_2233);
and U593 (N_593,In_1688,In_967);
xor U594 (N_594,In_643,In_57);
xnor U595 (N_595,N_141,N_294);
nor U596 (N_596,In_2476,In_930);
nand U597 (N_597,In_1748,In_175);
xor U598 (N_598,In_636,In_2453);
and U599 (N_599,In_2076,In_2518);
xor U600 (N_600,In_2262,In_862);
nand U601 (N_601,N_49,In_2902);
nor U602 (N_602,In_1593,In_829);
nand U603 (N_603,In_2111,In_2214);
nor U604 (N_604,In_2287,N_336);
and U605 (N_605,In_1264,N_335);
xor U606 (N_606,In_1142,In_84);
xnor U607 (N_607,In_2305,In_2658);
or U608 (N_608,N_338,In_1517);
nor U609 (N_609,In_491,In_1434);
or U610 (N_610,N_300,In_1852);
or U611 (N_611,In_109,N_316);
or U612 (N_612,N_576,In_1018);
and U613 (N_613,In_2622,In_1905);
xnor U614 (N_614,In_1343,In_811);
xnor U615 (N_615,In_1979,In_923);
nor U616 (N_616,N_522,In_1656);
xor U617 (N_617,In_2840,In_1058);
and U618 (N_618,N_485,In_1674);
or U619 (N_619,N_306,In_832);
and U620 (N_620,In_1902,In_1532);
nand U621 (N_621,In_624,N_398);
or U622 (N_622,In_1086,In_2170);
xor U623 (N_623,N_412,In_1914);
nor U624 (N_624,In_1403,In_2192);
nand U625 (N_625,In_845,In_355);
and U626 (N_626,N_381,In_996);
or U627 (N_627,In_2730,In_760);
nand U628 (N_628,N_174,N_111);
nor U629 (N_629,In_1009,In_2535);
nor U630 (N_630,In_1809,In_751);
or U631 (N_631,In_95,In_2626);
nor U632 (N_632,In_2496,In_2713);
or U633 (N_633,N_467,In_1549);
nor U634 (N_634,In_2606,N_493);
xnor U635 (N_635,In_2944,In_82);
nand U636 (N_636,In_1226,In_2185);
and U637 (N_637,In_709,In_2754);
xor U638 (N_638,N_329,In_1865);
nor U639 (N_639,In_2120,In_2260);
or U640 (N_640,In_665,In_1799);
nand U641 (N_641,In_615,In_1507);
nand U642 (N_642,In_1771,N_169);
nand U643 (N_643,In_1879,N_293);
xor U644 (N_644,In_2734,In_461);
nor U645 (N_645,In_1171,N_36);
and U646 (N_646,In_2533,N_102);
nand U647 (N_647,In_654,In_2673);
and U648 (N_648,In_2989,In_2441);
and U649 (N_649,In_318,In_1727);
or U650 (N_650,In_214,N_472);
or U651 (N_651,In_2049,N_34);
or U652 (N_652,N_263,In_2638);
nor U653 (N_653,In_2015,In_1792);
nor U654 (N_654,In_1074,In_1114);
xor U655 (N_655,In_1302,N_262);
and U656 (N_656,N_170,In_869);
nand U657 (N_657,In_2777,In_1237);
nand U658 (N_658,N_98,In_898);
and U659 (N_659,N_47,In_1190);
and U660 (N_660,In_2557,In_173);
or U661 (N_661,In_321,In_510);
nor U662 (N_662,In_2290,N_84);
nand U663 (N_663,In_1387,In_2433);
nor U664 (N_664,In_980,In_329);
xor U665 (N_665,In_2828,In_1745);
xnor U666 (N_666,In_1155,In_2138);
or U667 (N_667,In_2610,In_2031);
xnor U668 (N_668,In_671,In_119);
nand U669 (N_669,In_478,N_295);
and U670 (N_670,N_205,N_369);
and U671 (N_671,In_2310,In_281);
xnor U672 (N_672,N_178,In_176);
nor U673 (N_673,N_87,N_208);
xor U674 (N_674,In_1833,In_506);
nand U675 (N_675,In_414,N_242);
and U676 (N_676,In_1331,In_2383);
nor U677 (N_677,In_394,In_430);
and U678 (N_678,N_340,In_562);
nand U679 (N_679,In_973,In_448);
nand U680 (N_680,In_203,In_446);
xor U681 (N_681,In_2931,In_2924);
nand U682 (N_682,In_2190,In_2891);
xnor U683 (N_683,In_547,In_2335);
nand U684 (N_684,In_1581,In_2791);
or U685 (N_685,In_794,In_1785);
xnor U686 (N_686,In_2896,In_2399);
nand U687 (N_687,In_1988,In_1677);
nand U688 (N_688,N_587,In_1279);
xor U689 (N_689,In_2500,In_341);
and U690 (N_690,In_163,In_1608);
or U691 (N_691,In_1039,N_238);
xnor U692 (N_692,In_258,In_2406);
xor U693 (N_693,In_1591,In_2919);
nand U694 (N_694,N_62,N_70);
or U695 (N_695,N_516,In_196);
nand U696 (N_696,N_213,In_2105);
and U697 (N_697,In_1177,In_2449);
xnor U698 (N_698,In_2093,In_999);
and U699 (N_699,In_1136,N_210);
xor U700 (N_700,In_2737,In_2576);
nand U701 (N_701,N_598,In_454);
xnor U702 (N_702,In_2339,In_2783);
xor U703 (N_703,In_1776,In_2035);
nor U704 (N_704,N_298,In_734);
nand U705 (N_705,In_1554,In_431);
or U706 (N_706,In_2241,N_498);
nor U707 (N_707,In_2652,In_2444);
or U708 (N_708,In_1291,In_1483);
nor U709 (N_709,In_718,In_1686);
nand U710 (N_710,In_1563,N_211);
xnor U711 (N_711,In_1148,In_2494);
nand U712 (N_712,In_67,In_1664);
and U713 (N_713,In_2601,N_234);
nor U714 (N_714,In_2379,In_71);
or U715 (N_715,In_2926,N_26);
nor U716 (N_716,In_2215,In_1970);
and U717 (N_717,In_2579,N_553);
or U718 (N_718,In_1378,In_1927);
xor U719 (N_719,In_987,In_2945);
nor U720 (N_720,In_1642,In_1014);
or U721 (N_721,In_1062,In_2759);
xnor U722 (N_722,N_182,In_436);
nand U723 (N_723,In_2054,N_289);
nor U724 (N_724,In_2300,In_78);
and U725 (N_725,In_159,In_1969);
nand U726 (N_726,In_1811,In_1840);
and U727 (N_727,In_2811,In_777);
or U728 (N_728,In_2694,In_2700);
nand U729 (N_729,In_1307,N_142);
or U730 (N_730,In_77,In_1294);
xnor U731 (N_731,N_480,In_129);
and U732 (N_732,N_78,In_2657);
nor U733 (N_733,In_1981,In_2930);
nor U734 (N_734,In_2870,In_630);
or U735 (N_735,In_2131,In_883);
nor U736 (N_736,In_649,In_1592);
or U737 (N_737,In_1244,In_2116);
and U738 (N_738,In_669,In_2526);
and U739 (N_739,N_473,N_120);
and U740 (N_740,In_293,In_2578);
or U741 (N_741,In_1550,In_1724);
or U742 (N_742,In_83,In_697);
nor U743 (N_743,In_1092,In_1052);
xnor U744 (N_744,In_1894,N_387);
and U745 (N_745,In_971,In_979);
or U746 (N_746,N_439,N_6);
and U747 (N_747,In_653,In_753);
xnor U748 (N_748,In_112,In_2271);
nor U749 (N_749,In_2817,In_2304);
nor U750 (N_750,In_2318,In_929);
and U751 (N_751,In_2361,N_8);
xor U752 (N_752,In_1973,In_1871);
or U753 (N_753,N_582,In_79);
and U754 (N_754,In_2667,In_2171);
nand U755 (N_755,In_2723,In_755);
and U756 (N_756,N_318,In_1017);
nand U757 (N_757,In_2682,N_226);
or U758 (N_758,In_1985,N_19);
nor U759 (N_759,In_1408,In_2443);
nor U760 (N_760,N_40,In_859);
nand U761 (N_761,In_774,In_807);
nand U762 (N_762,In_978,In_2841);
nor U763 (N_763,In_18,In_2179);
or U764 (N_764,N_198,In_1042);
xor U765 (N_765,In_694,N_419);
nor U766 (N_766,In_2353,In_2309);
nand U767 (N_767,In_2637,N_462);
nor U768 (N_768,In_287,In_1909);
nand U769 (N_769,In_626,In_459);
or U770 (N_770,In_92,In_117);
and U771 (N_771,N_592,In_1184);
or U772 (N_772,In_1628,In_36);
nand U773 (N_773,In_2543,In_1984);
nand U774 (N_774,In_425,In_1484);
xnor U775 (N_775,In_555,In_1487);
and U776 (N_776,In_1881,In_849);
nor U777 (N_777,In_1641,In_2194);
xnor U778 (N_778,In_1860,In_1224);
nor U779 (N_779,In_570,In_1635);
nor U780 (N_780,N_434,In_284);
nor U781 (N_781,N_481,In_645);
or U782 (N_782,In_655,In_86);
nand U783 (N_783,In_629,N_33);
or U784 (N_784,In_481,In_2747);
and U785 (N_785,In_1807,In_2187);
or U786 (N_786,In_896,In_865);
xnor U787 (N_787,In_2714,N_183);
nand U788 (N_788,In_2521,In_1438);
or U789 (N_789,N_580,N_416);
nand U790 (N_790,In_2283,In_1118);
nor U791 (N_791,In_721,N_413);
and U792 (N_792,In_2906,N_461);
and U793 (N_793,In_2104,In_250);
xor U794 (N_794,N_105,In_2760);
nor U795 (N_795,In_2008,In_1186);
xor U796 (N_796,In_210,In_1759);
and U797 (N_797,In_1806,In_2140);
or U798 (N_798,N_144,N_588);
xor U799 (N_799,In_1504,N_489);
or U800 (N_800,N_313,N_433);
and U801 (N_801,In_1966,N_151);
and U802 (N_802,N_303,N_254);
and U803 (N_803,In_423,In_2220);
and U804 (N_804,In_650,In_1521);
nand U805 (N_805,In_1649,N_44);
and U806 (N_806,In_1546,In_2091);
and U807 (N_807,In_1736,N_312);
nand U808 (N_808,In_1494,N_358);
and U809 (N_809,In_2299,N_486);
nor U810 (N_810,In_1876,In_2303);
xnor U811 (N_811,In_2014,In_223);
or U812 (N_812,In_2225,In_1519);
xor U813 (N_813,In_1325,In_1059);
nand U814 (N_814,In_916,In_1365);
xor U815 (N_815,In_1906,In_2586);
xnor U816 (N_816,N_476,In_2957);
nand U817 (N_817,In_1866,In_1139);
or U818 (N_818,In_2266,In_2413);
nand U819 (N_819,In_2013,In_1115);
xor U820 (N_820,N_180,N_227);
and U821 (N_821,N_265,In_1492);
or U822 (N_822,In_1606,In_2753);
or U823 (N_823,In_1000,In_2445);
and U824 (N_824,In_1853,N_518);
nor U825 (N_825,In_765,In_815);
nand U826 (N_826,In_104,N_195);
nand U827 (N_827,In_1202,In_2792);
nor U828 (N_828,In_137,In_909);
and U829 (N_829,In_1841,N_400);
nand U830 (N_830,In_2647,N_310);
nor U831 (N_831,N_521,In_2041);
or U832 (N_832,In_1069,In_1267);
xnor U833 (N_833,In_6,N_375);
and U834 (N_834,N_217,In_1064);
nor U835 (N_835,In_529,In_2440);
or U836 (N_836,In_2137,In_1485);
nand U837 (N_837,In_1087,N_405);
nor U838 (N_838,In_2540,In_1084);
or U839 (N_839,In_302,N_560);
nand U840 (N_840,In_142,In_66);
nor U841 (N_841,In_405,In_1797);
and U842 (N_842,In_2381,In_2382);
nand U843 (N_843,In_2246,In_2807);
nand U844 (N_844,In_596,In_2551);
xnor U845 (N_845,N_373,In_2550);
nand U846 (N_846,N_586,In_563);
and U847 (N_847,In_20,In_1590);
or U848 (N_848,N_269,In_2574);
nand U849 (N_849,In_310,In_1854);
or U850 (N_850,In_218,In_2890);
nand U851 (N_851,N_204,In_237);
and U852 (N_852,In_236,In_800);
xnor U853 (N_853,In_872,In_2280);
nand U854 (N_854,In_1435,In_2686);
or U855 (N_855,In_882,In_122);
nand U856 (N_856,In_647,In_312);
nor U857 (N_857,N_326,In_335);
or U858 (N_858,N_243,In_143);
and U859 (N_859,N_50,In_1755);
xnor U860 (N_860,In_339,In_683);
xnor U861 (N_861,In_2806,In_2255);
nor U862 (N_862,In_1120,In_1940);
nand U863 (N_863,In_2986,N_589);
xor U864 (N_864,N_547,In_1758);
xor U865 (N_865,In_625,In_1215);
xor U866 (N_866,In_918,In_2088);
xnor U867 (N_867,In_463,In_2253);
xnor U868 (N_868,In_891,N_428);
nand U869 (N_869,In_1335,N_458);
xnor U870 (N_870,N_278,In_1366);
nor U871 (N_871,In_1015,In_604);
nor U872 (N_872,In_954,In_1256);
or U873 (N_873,N_282,In_736);
or U874 (N_874,In_1845,In_1765);
xnor U875 (N_875,In_902,In_2803);
xnor U876 (N_876,In_1181,In_663);
nor U877 (N_877,N_96,In_538);
or U878 (N_878,N_590,In_2645);
xnor U879 (N_879,In_912,In_1775);
nand U880 (N_880,N_92,In_2169);
xnor U881 (N_881,N_5,In_202);
nor U882 (N_882,In_1595,In_2793);
nor U883 (N_883,In_408,In_2217);
nand U884 (N_884,N_161,In_895);
nand U885 (N_885,In_1803,In_580);
or U886 (N_886,In_818,In_1121);
xor U887 (N_887,In_1105,In_1023);
or U888 (N_888,In_387,N_429);
nor U889 (N_889,In_1348,N_350);
or U890 (N_890,In_512,In_1313);
nand U891 (N_891,N_555,In_674);
and U892 (N_892,N_363,In_52);
and U893 (N_893,N_530,In_1689);
xor U894 (N_894,In_756,In_2267);
xor U895 (N_895,N_519,In_1959);
xnor U896 (N_896,In_1289,In_2059);
and U897 (N_897,N_212,In_659);
nor U898 (N_898,In_254,In_2256);
and U899 (N_899,In_2997,In_899);
or U900 (N_900,In_2810,In_897);
or U901 (N_901,In_27,In_565);
nor U902 (N_902,N_661,In_2939);
xnor U903 (N_903,In_1614,N_426);
nand U904 (N_904,In_1534,N_797);
and U905 (N_905,N_477,In_1821);
nor U906 (N_906,N_726,N_713);
and U907 (N_907,In_1410,N_675);
and U908 (N_908,In_378,N_688);
nor U909 (N_909,N_256,In_2766);
xor U910 (N_910,In_761,N_130);
nor U911 (N_911,N_526,N_847);
xor U912 (N_912,In_2397,N_370);
nand U913 (N_913,N_711,In_160);
or U914 (N_914,In_2395,In_2043);
nand U915 (N_915,N_332,In_792);
and U916 (N_916,In_706,In_338);
nor U917 (N_917,In_590,N_389);
nor U918 (N_918,N_349,In_2603);
nor U919 (N_919,In_594,N_892);
nor U920 (N_920,N_478,In_1433);
or U921 (N_921,In_1713,N_658);
or U922 (N_922,In_2684,In_1153);
nand U923 (N_923,In_1597,In_2084);
nand U924 (N_924,N_500,In_2633);
xnor U925 (N_925,In_123,In_1013);
xor U926 (N_926,N_497,N_888);
and U927 (N_927,In_1330,In_2263);
xor U928 (N_928,N_642,In_2075);
xnor U929 (N_929,In_2660,In_356);
nor U930 (N_930,N_828,In_1227);
or U931 (N_931,In_1028,In_2352);
nor U932 (N_932,N_292,In_1699);
nor U933 (N_933,N_571,In_835);
or U934 (N_934,N_746,N_418);
nand U935 (N_935,In_1652,N_315);
or U936 (N_936,In_1638,In_1762);
and U937 (N_937,In_520,N_787);
or U938 (N_938,In_1648,In_1961);
nand U939 (N_939,In_361,In_1669);
and U940 (N_940,N_861,In_1356);
nor U941 (N_941,N_837,In_809);
nand U942 (N_942,In_965,In_2503);
and U943 (N_943,N_859,In_1572);
nor U944 (N_944,In_1982,In_2910);
nor U945 (N_945,In_1863,N_346);
nand U946 (N_946,In_1437,In_1716);
and U947 (N_947,N_495,In_1586);
xnor U948 (N_948,In_2386,N_743);
or U949 (N_949,In_773,N_855);
nand U950 (N_950,N_602,N_348);
or U951 (N_951,In_2865,In_724);
nor U952 (N_952,In_942,In_1825);
nand U953 (N_953,In_413,In_2173);
or U954 (N_954,In_1423,In_2829);
nand U955 (N_955,In_2653,In_322);
nand U956 (N_956,N_873,N_817);
nand U957 (N_957,In_364,In_924);
xor U958 (N_958,N_803,In_265);
xnor U959 (N_959,N_705,N_784);
nor U960 (N_960,In_2744,In_2323);
and U961 (N_961,In_14,In_2307);
and U962 (N_962,In_1588,In_1116);
or U963 (N_963,In_2153,In_1037);
nor U964 (N_964,In_848,N_425);
nand U965 (N_965,In_447,In_2756);
and U966 (N_966,N_722,In_539);
nor U967 (N_967,In_2135,In_2426);
and U968 (N_968,N_769,In_2990);
nor U969 (N_969,N_549,N_830);
and U970 (N_970,In_1728,In_2729);
xor U971 (N_971,In_2040,In_2609);
nor U972 (N_972,In_597,In_2755);
and U973 (N_973,N_324,N_512);
and U974 (N_974,In_808,N_376);
and U975 (N_975,In_533,In_827);
and U976 (N_976,N_727,In_2017);
nor U977 (N_977,N_14,N_501);
and U978 (N_978,In_1539,In_2731);
xnor U979 (N_979,N_625,In_1622);
and U980 (N_980,In_2933,In_1463);
and U981 (N_981,In_2007,In_992);
xnor U982 (N_982,In_399,In_616);
and U983 (N_983,In_830,N_643);
xor U984 (N_984,In_1270,In_2062);
or U985 (N_985,In_783,N_684);
and U986 (N_986,In_2034,N_758);
and U987 (N_987,N_634,In_2691);
nor U988 (N_988,In_2876,N_449);
nand U989 (N_989,In_1468,In_727);
nand U990 (N_990,In_2102,N_157);
nor U991 (N_991,In_803,In_2640);
xnor U992 (N_992,N_159,In_1872);
or U993 (N_993,In_2146,N_520);
nand U994 (N_994,In_2359,In_2313);
and U995 (N_995,In_525,N_465);
or U996 (N_996,N_621,N_341);
and U997 (N_997,In_2748,In_587);
or U998 (N_998,N_510,In_2477);
nor U999 (N_999,N_409,N_680);
and U1000 (N_1000,N_708,N_583);
and U1001 (N_1001,In_1609,In_2005);
xnor U1002 (N_1002,In_600,In_1993);
xor U1003 (N_1003,N_557,In_2134);
and U1004 (N_1004,N_552,In_1180);
and U1005 (N_1005,N_786,In_1106);
xnor U1006 (N_1006,In_2592,In_1646);
nand U1007 (N_1007,N_774,In_2577);
xnor U1008 (N_1008,N_424,N_763);
xnor U1009 (N_1009,In_2758,In_201);
nand U1010 (N_1010,N_836,N_41);
or U1011 (N_1011,In_2769,In_2182);
nor U1012 (N_1012,N_606,N_755);
or U1013 (N_1013,In_1788,In_389);
or U1014 (N_1014,In_1150,N_435);
or U1015 (N_1015,In_858,In_758);
nor U1016 (N_1016,In_443,In_264);
nor U1017 (N_1017,In_810,N_484);
and U1018 (N_1018,In_2916,In_704);
or U1019 (N_1019,N_559,In_2768);
or U1020 (N_1020,In_34,In_96);
xor U1021 (N_1021,In_17,N_452);
or U1022 (N_1022,N_514,N_783);
xor U1023 (N_1023,N_647,In_608);
and U1024 (N_1024,In_518,In_1355);
nor U1025 (N_1025,In_1119,N_185);
nor U1026 (N_1026,N_683,In_2915);
nor U1027 (N_1027,In_1341,N_206);
and U1028 (N_1028,In_396,In_1100);
nor U1029 (N_1029,N_445,In_2115);
nor U1030 (N_1030,In_1413,In_970);
or U1031 (N_1031,In_2385,In_332);
or U1032 (N_1032,N_406,In_370);
nand U1033 (N_1033,In_1462,In_584);
nand U1034 (N_1034,N_394,N_532);
nor U1035 (N_1035,N_868,In_2727);
nor U1036 (N_1036,In_1928,In_1885);
nand U1037 (N_1037,In_225,N_357);
nand U1038 (N_1038,In_2863,N_95);
and U1039 (N_1039,In_839,N_155);
and U1040 (N_1040,In_12,In_1721);
nor U1041 (N_1041,In_1601,In_2884);
and U1042 (N_1042,N_648,N_832);
nand U1043 (N_1043,N_678,N_890);
nand U1044 (N_1044,N_566,In_1096);
xnor U1045 (N_1045,N_599,In_2798);
or U1046 (N_1046,In_2183,In_1931);
and U1047 (N_1047,In_2556,In_1671);
nor U1048 (N_1048,N_575,In_2553);
nand U1049 (N_1049,In_2587,In_2369);
or U1050 (N_1050,In_1389,In_1383);
or U1051 (N_1051,In_2663,N_407);
nand U1052 (N_1052,In_85,N_851);
xor U1053 (N_1053,N_591,In_1221);
or U1054 (N_1054,In_1938,N_454);
or U1055 (N_1055,In_2644,In_342);
and U1056 (N_1056,In_1286,In_770);
or U1057 (N_1057,N_444,In_610);
nor U1058 (N_1058,In_732,In_1322);
xnor U1059 (N_1059,N_443,In_1205);
nand U1060 (N_1060,In_1131,N_569);
nor U1061 (N_1061,N_739,In_2236);
and U1062 (N_1062,N_192,In_867);
and U1063 (N_1063,In_1469,In_675);
or U1064 (N_1064,N_456,In_1169);
xor U1065 (N_1065,In_2032,In_319);
nand U1066 (N_1066,In_2486,In_1238);
xnor U1067 (N_1067,N_117,N_10);
or U1068 (N_1068,In_401,In_2240);
or U1069 (N_1069,In_2719,N_704);
and U1070 (N_1070,In_2286,N_618);
nor U1071 (N_1071,In_505,In_2848);
xor U1072 (N_1072,N_184,N_664);
xor U1073 (N_1073,N_649,In_2580);
nand U1074 (N_1074,In_2479,N_490);
or U1075 (N_1075,In_1947,In_1470);
xor U1076 (N_1076,In_2920,N_731);
nand U1077 (N_1077,In_1321,N_160);
xnor U1078 (N_1078,In_157,In_1751);
nand U1079 (N_1079,In_2222,In_951);
nand U1080 (N_1080,N_534,In_2544);
or U1081 (N_1081,In_1466,In_442);
nor U1082 (N_1082,N_574,N_796);
nand U1083 (N_1083,N_115,In_804);
nand U1084 (N_1084,N_251,In_1529);
nor U1085 (N_1085,N_561,In_2883);
xor U1086 (N_1086,In_1603,In_2794);
nor U1087 (N_1087,In_1068,In_566);
nand U1088 (N_1088,In_2571,In_1780);
or U1089 (N_1089,In_1731,In_2615);
nor U1090 (N_1090,N_760,In_2886);
or U1091 (N_1091,In_1409,In_350);
nor U1092 (N_1092,N_753,In_1067);
or U1093 (N_1093,In_2319,In_741);
nor U1094 (N_1094,In_189,In_798);
and U1095 (N_1095,In_1376,In_1432);
nor U1096 (N_1096,N_750,In_1239);
xor U1097 (N_1097,N_43,In_1133);
nand U1098 (N_1098,In_2836,In_917);
nand U1099 (N_1099,In_88,In_2471);
xnor U1100 (N_1100,In_1022,In_2833);
nor U1101 (N_1101,N_149,In_2330);
or U1102 (N_1102,N_18,In_2821);
nand U1103 (N_1103,In_2150,In_685);
nand U1104 (N_1104,N_247,In_528);
xnor U1105 (N_1105,In_2538,N_9);
and U1106 (N_1106,N_321,In_789);
and U1107 (N_1107,N_468,In_1367);
or U1108 (N_1108,In_1088,In_781);
or U1109 (N_1109,N_624,N_228);
nor U1110 (N_1110,N_197,N_127);
nor U1111 (N_1111,In_2685,In_2158);
or U1112 (N_1112,In_1362,In_1243);
or U1113 (N_1113,In_1094,In_2343);
xor U1114 (N_1114,In_878,N_201);
nor U1115 (N_1115,In_2515,N_30);
or U1116 (N_1116,In_2976,In_208);
or U1117 (N_1117,In_1524,In_1108);
xor U1118 (N_1118,N_728,In_422);
xnor U1119 (N_1119,N_464,In_1132);
or U1120 (N_1120,N_322,In_349);
and U1121 (N_1121,N_432,In_632);
nand U1122 (N_1122,N_250,N_535);
xnor U1123 (N_1123,In_1386,N_898);
or U1124 (N_1124,N_23,In_2929);
or U1125 (N_1125,In_296,N_878);
nand U1126 (N_1126,In_2635,N_483);
or U1127 (N_1127,In_395,N_471);
nand U1128 (N_1128,In_2439,N_706);
nand U1129 (N_1129,In_676,N_687);
nand U1130 (N_1130,In_825,N_367);
or U1131 (N_1131,In_1734,N_820);
nand U1132 (N_1132,In_2639,In_98);
xor U1133 (N_1133,In_295,In_1375);
and U1134 (N_1134,In_1535,N_167);
or U1135 (N_1135,In_1388,N_276);
nand U1136 (N_1136,In_2717,In_228);
xnor U1137 (N_1137,In_2357,In_15);
and U1138 (N_1138,In_1877,In_2938);
or U1139 (N_1139,In_2425,In_1849);
or U1140 (N_1140,In_1007,In_1449);
and U1141 (N_1141,In_841,N_114);
nor U1142 (N_1142,In_888,N_273);
nand U1143 (N_1143,In_1066,In_1295);
nor U1144 (N_1144,In_2473,N_66);
or U1145 (N_1145,In_1996,In_2419);
or U1146 (N_1146,In_716,In_1209);
or U1147 (N_1147,N_857,In_2681);
xnor U1148 (N_1148,N_882,In_2080);
or U1149 (N_1149,In_1047,In_1041);
nand U1150 (N_1150,In_2600,In_2206);
and U1151 (N_1151,N_399,In_714);
xor U1152 (N_1152,N_58,N_674);
nor U1153 (N_1153,N_347,In_1903);
or U1154 (N_1154,N_382,In_1878);
and U1155 (N_1155,In_1893,In_2269);
xnor U1156 (N_1156,In_1990,In_1240);
or U1157 (N_1157,In_1757,N_320);
or U1158 (N_1158,In_2312,In_2655);
nand U1159 (N_1159,N_646,In_1125);
or U1160 (N_1160,In_404,N_378);
nor U1161 (N_1161,In_2774,In_2167);
xnor U1162 (N_1162,N_697,In_1766);
nor U1163 (N_1163,In_2614,In_507);
xnor U1164 (N_1164,N_74,N_177);
and U1165 (N_1165,In_2703,In_976);
nand U1166 (N_1166,N_551,N_756);
nor U1167 (N_1167,In_1868,In_279);
nor U1168 (N_1168,In_501,N_437);
nor U1169 (N_1169,In_1533,In_605);
and U1170 (N_1170,In_713,In_383);
or U1171 (N_1171,In_2184,N_345);
nand U1172 (N_1172,N_427,In_410);
xnor U1173 (N_1173,In_44,In_745);
or U1174 (N_1174,N_867,In_1162);
nand U1175 (N_1175,In_641,N_511);
xnor U1176 (N_1176,N_296,N_301);
xnor U1177 (N_1177,N_99,N_11);
nand U1178 (N_1178,In_1695,In_2985);
and U1179 (N_1179,N_362,N_368);
and U1180 (N_1180,In_1943,In_1624);
and U1181 (N_1181,In_1036,In_1613);
nand U1182 (N_1182,N_866,In_1598);
and U1183 (N_1183,In_80,In_1165);
or U1184 (N_1184,In_1051,N_266);
nor U1185 (N_1185,N_359,N_258);
nand U1186 (N_1186,In_695,In_1714);
and U1187 (N_1187,In_526,N_253);
nor U1188 (N_1188,In_824,N_422);
nor U1189 (N_1189,In_611,In_884);
or U1190 (N_1190,In_1164,N_702);
nand U1191 (N_1191,N_872,In_2350);
xnor U1192 (N_1192,N_430,In_2721);
or U1193 (N_1193,N_811,In_913);
xor U1194 (N_1194,In_1932,In_719);
or U1195 (N_1195,N_773,In_2788);
xor U1196 (N_1196,In_2569,In_583);
xor U1197 (N_1197,In_118,In_206);
nand U1198 (N_1198,N_81,In_269);
and U1199 (N_1199,In_403,N_654);
nand U1200 (N_1200,In_2678,In_995);
and U1201 (N_1201,In_19,In_127);
nand U1202 (N_1202,In_1323,In_1455);
nor U1203 (N_1203,In_2415,In_1512);
nor U1204 (N_1204,In_972,N_938);
xor U1205 (N_1205,N_546,N_239);
or U1206 (N_1206,N_805,In_2159);
nand U1207 (N_1207,In_1020,In_1948);
nand U1208 (N_1208,In_519,N_692);
and U1209 (N_1209,In_1907,N_264);
or U1210 (N_1210,N_460,In_601);
or U1211 (N_1211,N_798,In_2470);
or U1212 (N_1212,N_790,In_277);
and U1213 (N_1213,N_309,N_118);
or U1214 (N_1214,N_952,In_1274);
or U1215 (N_1215,N_488,N_83);
or U1216 (N_1216,N_333,N_865);
nand U1217 (N_1217,In_1134,N_441);
xor U1218 (N_1218,In_1427,In_2342);
xnor U1219 (N_1219,In_2119,N_563);
or U1220 (N_1220,N_923,N_655);
and U1221 (N_1221,N_810,N_1054);
and U1222 (N_1222,N_420,In_985);
nor U1223 (N_1223,N_813,N_408);
and U1224 (N_1224,N_390,N_189);
or U1225 (N_1225,In_2186,N_355);
nand U1226 (N_1226,N_730,N_288);
xor U1227 (N_1227,In_288,In_593);
nand U1228 (N_1228,In_1189,In_1627);
nand U1229 (N_1229,In_801,In_1805);
and U1230 (N_1230,In_2257,N_344);
nor U1231 (N_1231,N_1044,In_708);
or U1232 (N_1232,N_327,In_1182);
nand U1233 (N_1233,In_1093,N_106);
and U1234 (N_1234,In_1794,In_2573);
xnor U1235 (N_1235,N_679,N_353);
xnor U1236 (N_1236,In_2958,In_1206);
and U1237 (N_1237,N_966,In_99);
nor U1238 (N_1238,In_1203,In_1031);
and U1239 (N_1239,In_1619,N_1067);
or U1240 (N_1240,In_543,N_261);
xnor U1241 (N_1241,N_165,N_1159);
nand U1242 (N_1242,In_139,In_1971);
xnor U1243 (N_1243,In_2368,In_564);
and U1244 (N_1244,N_794,N_116);
xor U1245 (N_1245,N_523,In_1198);
or U1246 (N_1246,In_1640,N_1079);
xnor U1247 (N_1247,In_1002,In_2911);
nor U1248 (N_1248,N_1055,In_2786);
xnor U1249 (N_1249,In_1103,N_759);
nor U1250 (N_1250,N_936,In_524);
nand U1251 (N_1251,In_2534,In_2235);
nand U1252 (N_1252,N_749,In_1848);
nor U1253 (N_1253,In_452,In_2757);
xnor U1254 (N_1254,N_668,In_1372);
and U1255 (N_1255,In_2000,In_1245);
xor U1256 (N_1256,In_2812,In_220);
xor U1257 (N_1257,In_2629,In_2491);
or U1258 (N_1258,In_1962,N_568);
nand U1259 (N_1259,N_470,N_1008);
nor U1260 (N_1260,N_37,In_2354);
and U1261 (N_1261,In_1999,N_187);
xor U1262 (N_1262,In_1138,In_2057);
or U1263 (N_1263,In_1208,N_685);
or U1264 (N_1264,In_2707,In_2234);
nand U1265 (N_1265,N_383,N_1018);
and U1266 (N_1266,N_856,In_2555);
or U1267 (N_1267,In_1406,In_2200);
nor U1268 (N_1268,In_696,N_970);
or U1269 (N_1269,N_319,N_1);
nand U1270 (N_1270,In_2089,In_1053);
nor U1271 (N_1271,In_1122,N_22);
and U1272 (N_1272,In_2772,In_2770);
nand U1273 (N_1273,In_1620,N_980);
and U1274 (N_1274,In_444,N_1023);
xnor U1275 (N_1275,N_920,In_323);
or U1276 (N_1276,N_1107,In_2999);
nor U1277 (N_1277,N_1006,N_955);
nor U1278 (N_1278,In_1163,In_2835);
xor U1279 (N_1279,In_1442,In_2051);
xor U1280 (N_1280,In_1284,N_987);
or U1281 (N_1281,In_2172,In_136);
xnor U1282 (N_1282,In_2654,In_1632);
nor U1283 (N_1283,In_1308,N_281);
nor U1284 (N_1284,In_2998,In_2431);
and U1285 (N_1285,In_2157,In_2701);
nand U1286 (N_1286,N_1030,In_2796);
nor U1287 (N_1287,N_1191,In_81);
or U1288 (N_1288,N_388,In_2340);
nand U1289 (N_1289,In_31,N_1140);
nor U1290 (N_1290,N_237,N_806);
or U1291 (N_1291,In_1795,In_110);
xor U1292 (N_1292,N_874,In_1071);
or U1293 (N_1293,In_2720,In_190);
xnor U1294 (N_1294,N_799,In_1032);
xnor U1295 (N_1295,In_582,N_173);
xor U1296 (N_1296,N_125,In_426);
xor U1297 (N_1297,N_932,In_1929);
nand U1298 (N_1298,In_2,In_1802);
nand U1299 (N_1299,N_1152,In_1417);
or U1300 (N_1300,In_453,In_1272);
nand U1301 (N_1301,In_1111,In_681);
xor U1302 (N_1302,In_2454,In_2585);
nor U1303 (N_1303,N_48,N_883);
nand U1304 (N_1304,N_985,In_2198);
and U1305 (N_1305,N_79,N_1021);
nor U1306 (N_1306,In_182,N_913);
nor U1307 (N_1307,N_463,N_75);
and U1308 (N_1308,N_1164,In_2819);
xnor U1309 (N_1309,N_506,N_1129);
and U1310 (N_1310,In_2805,N_507);
nand U1311 (N_1311,In_1715,In_940);
and U1312 (N_1312,N_248,In_2885);
or U1313 (N_1313,N_1015,In_2047);
and U1314 (N_1314,In_1659,In_1493);
nor U1315 (N_1315,In_2247,N_986);
xnor U1316 (N_1316,In_257,N_491);
xor U1317 (N_1317,N_732,In_1336);
nand U1318 (N_1318,In_90,N_627);
or U1319 (N_1319,N_287,N_7);
and U1320 (N_1320,N_1150,In_2324);
nor U1321 (N_1321,N_639,N_354);
nand U1322 (N_1322,In_151,In_419);
xnor U1323 (N_1323,In_2838,N_785);
nor U1324 (N_1324,In_2776,In_2211);
and U1325 (N_1325,N_834,N_1065);
or U1326 (N_1326,In_1219,In_1834);
or U1327 (N_1327,N_781,N_651);
nor U1328 (N_1328,In_493,In_1858);
or U1329 (N_1329,In_775,N_1011);
and U1330 (N_1330,In_1073,N_1082);
or U1331 (N_1331,In_1441,In_58);
nand U1332 (N_1332,In_1231,N_525);
nor U1333 (N_1333,In_1316,In_1694);
nand U1334 (N_1334,In_184,N_122);
or U1335 (N_1335,In_1983,N_0);
or U1336 (N_1336,N_976,In_1846);
nor U1337 (N_1337,N_707,In_492);
nor U1338 (N_1338,N_630,N_714);
or U1339 (N_1339,N_25,N_734);
xnor U1340 (N_1340,In_1478,N_603);
and U1341 (N_1341,In_1218,In_2106);
nor U1342 (N_1342,In_2018,In_1787);
nand U1343 (N_1343,In_797,In_1739);
xnor U1344 (N_1344,N_585,N_995);
nor U1345 (N_1345,N_1132,N_457);
nor U1346 (N_1346,N_1185,In_567);
nand U1347 (N_1347,In_351,In_1460);
and U1348 (N_1348,N_906,N_824);
nor U1349 (N_1349,In_2344,N_2);
nand U1350 (N_1350,In_1972,In_2082);
nor U1351 (N_1351,In_170,In_2278);
nor U1352 (N_1352,In_2165,In_33);
or U1353 (N_1353,N_1042,N_143);
nor U1354 (N_1354,In_407,N_567);
nand U1355 (N_1355,N_804,N_870);
nor U1356 (N_1356,N_842,N_818);
and U1357 (N_1357,N_918,In_938);
and U1358 (N_1358,N_885,In_1607);
xor U1359 (N_1359,In_1887,In_983);
xnor U1360 (N_1360,In_468,In_1920);
xnor U1361 (N_1361,N_751,In_2854);
nand U1362 (N_1362,N_748,N_1092);
nor U1363 (N_1363,In_2373,In_471);
and U1364 (N_1364,N_945,In_2704);
nand U1365 (N_1365,In_2532,In_603);
nor U1366 (N_1366,In_209,N_570);
nand U1367 (N_1367,In_2055,N_601);
or U1368 (N_1368,In_398,In_1277);
xor U1369 (N_1369,In_1384,In_1764);
or U1370 (N_1370,N_789,In_2827);
and U1371 (N_1371,In_2417,N_931);
and U1372 (N_1372,In_1357,In_1306);
nand U1373 (N_1373,N_843,N_741);
or U1374 (N_1374,N_221,In_550);
xnor U1375 (N_1375,N_949,N_297);
xnor U1376 (N_1376,In_2950,In_2662);
nand U1377 (N_1377,N_343,N_1102);
nand U1378 (N_1378,In_495,N_1167);
nand U1379 (N_1379,N_733,N_641);
nor U1380 (N_1380,In_2020,N_137);
nand U1381 (N_1381,N_39,In_2203);
nand U1382 (N_1382,In_102,In_549);
and U1383 (N_1383,N_482,N_241);
xnor U1384 (N_1384,In_962,N_1005);
nand U1385 (N_1385,In_1099,In_2857);
or U1386 (N_1386,N_610,In_542);
or U1387 (N_1387,N_629,N_608);
nor U1388 (N_1388,N_17,N_1004);
and U1389 (N_1389,In_1340,N_645);
xor U1390 (N_1390,N_821,In_1197);
and U1391 (N_1391,In_1687,In_2387);
or U1392 (N_1392,N_128,In_1987);
and U1393 (N_1393,In_1195,In_2282);
nand U1394 (N_1394,In_262,In_945);
xor U1395 (N_1395,N_1075,In_2887);
or U1396 (N_1396,N_176,In_76);
xor U1397 (N_1397,In_456,N_101);
nor U1398 (N_1398,In_353,N_822);
xnor U1399 (N_1399,N_930,N_776);
and U1400 (N_1400,N_1038,In_1706);
nor U1401 (N_1401,In_1318,N_397);
nor U1402 (N_1402,In_2056,In_534);
xor U1403 (N_1403,In_2784,N_812);
nand U1404 (N_1404,In_133,N_988);
or U1405 (N_1405,N_1144,In_2164);
nand U1406 (N_1406,N_1177,In_2010);
and U1407 (N_1407,N_660,N_916);
or U1408 (N_1408,In_1998,In_166);
or U1409 (N_1409,In_1604,In_960);
xnor U1410 (N_1410,N_941,In_2147);
or U1411 (N_1411,In_1527,N_778);
nor U1412 (N_1412,N_360,In_424);
xnor U1413 (N_1413,In_544,N_479);
nand U1414 (N_1414,In_1654,N_1016);
or U1415 (N_1415,N_1033,N_665);
and U1416 (N_1416,In_1418,N_508);
nor U1417 (N_1417,In_2631,In_1804);
xor U1418 (N_1418,In_633,N_1062);
or U1419 (N_1419,N_948,N_997);
nand U1420 (N_1420,In_2081,In_1618);
nand U1421 (N_1421,N_31,In_2098);
nand U1422 (N_1422,In_244,In_1451);
xnor U1423 (N_1423,N_912,N_415);
and U1424 (N_1424,In_328,N_352);
nor U1425 (N_1425,In_2583,N_527);
and U1426 (N_1426,N_717,In_2038);
or U1427 (N_1427,In_1958,In_2548);
nand U1428 (N_1428,N_992,In_822);
xor U1429 (N_1429,In_69,In_787);
nor U1430 (N_1430,N_110,N_640);
nand U1431 (N_1431,In_2856,N_891);
nand U1432 (N_1432,In_2163,N_100);
and U1433 (N_1433,In_1922,N_894);
nand U1434 (N_1434,In_1685,In_1083);
xnor U1435 (N_1435,In_2670,N_154);
xnor U1436 (N_1436,In_2789,In_242);
xnor U1437 (N_1437,N_517,In_1568);
xor U1438 (N_1438,N_971,In_2362);
nand U1439 (N_1439,N_1048,In_2197);
or U1440 (N_1440,N_1149,In_135);
nand U1441 (N_1441,N_1074,In_1419);
and U1442 (N_1442,N_255,In_400);
and U1443 (N_1443,In_2495,N_351);
nor U1444 (N_1444,In_2696,In_2363);
xnor U1445 (N_1445,N_1151,In_627);
and U1446 (N_1446,N_1088,In_238);
or U1447 (N_1447,In_1730,In_1707);
xor U1448 (N_1448,N_807,In_1426);
nand U1449 (N_1449,N_163,N_232);
nor U1450 (N_1450,In_2782,In_684);
and U1451 (N_1451,In_1992,N_862);
xnor U1452 (N_1452,N_1130,In_35);
and U1453 (N_1453,In_700,In_2951);
xor U1454 (N_1454,In_1663,N_1168);
or U1455 (N_1455,In_1414,N_1162);
nand U1456 (N_1456,N_1073,N_544);
and U1457 (N_1457,N_1039,N_15);
nand U1458 (N_1458,N_541,N_1097);
and U1459 (N_1459,N_131,In_1405);
nand U1460 (N_1460,In_2103,In_1711);
or U1461 (N_1461,N_401,N_27);
or U1462 (N_1462,In_1542,In_343);
or U1463 (N_1463,In_1749,N_835);
nand U1464 (N_1464,In_2298,In_1257);
and U1465 (N_1465,In_207,N_849);
or U1466 (N_1466,In_677,N_356);
nand U1467 (N_1467,In_1396,N_32);
and U1468 (N_1468,N_223,N_942);
or U1469 (N_1469,N_1158,N_21);
and U1470 (N_1470,In_2094,In_496);
nor U1471 (N_1471,In_2045,N_440);
nor U1472 (N_1472,N_777,In_1977);
xnor U1473 (N_1473,In_975,In_802);
nor U1474 (N_1474,N_1064,In_831);
or U1475 (N_1475,In_1869,In_1444);
nand U1476 (N_1476,In_2332,N_676);
nand U1477 (N_1477,N_994,In_1838);
or U1478 (N_1478,In_2492,In_2715);
nor U1479 (N_1479,In_1299,In_2804);
or U1480 (N_1480,N_919,N_45);
and U1481 (N_1481,In_2937,In_232);
or U1482 (N_1482,N_937,N_1115);
xnor U1483 (N_1483,N_1083,N_615);
nor U1484 (N_1484,In_191,In_2814);
xnor U1485 (N_1485,In_276,N_1133);
xnor U1486 (N_1486,In_2752,In_2109);
or U1487 (N_1487,In_2740,In_699);
xor U1488 (N_1488,N_209,In_2274);
or U1489 (N_1489,In_553,In_1003);
nor U1490 (N_1490,N_219,In_367);
xnor U1491 (N_1491,N_747,In_1560);
and U1492 (N_1492,In_936,N_203);
xnor U1493 (N_1493,N_436,In_435);
nor U1494 (N_1494,N_474,N_164);
or U1495 (N_1495,In_2642,In_1174);
nor U1496 (N_1496,In_2349,N_168);
nor U1497 (N_1497,In_717,In_1842);
xor U1498 (N_1498,N_914,N_1003);
or U1499 (N_1499,N_698,N_1032);
xor U1500 (N_1500,N_1146,N_1181);
nand U1501 (N_1501,In_1034,N_983);
or U1502 (N_1502,N_1324,N_927);
xor U1503 (N_1503,In_722,N_723);
or U1504 (N_1504,N_626,In_21);
xnor U1505 (N_1505,N_494,In_313);
nand U1506 (N_1506,In_2531,N_720);
nand U1507 (N_1507,N_1499,In_1605);
and U1508 (N_1508,N_76,N_939);
nand U1509 (N_1509,N_1411,N_917);
nor U1510 (N_1510,In_450,N_1301);
nor U1511 (N_1511,N_533,N_984);
xnor U1512 (N_1512,In_1763,In_546);
or U1513 (N_1513,N_1470,N_1256);
or U1514 (N_1514,In_470,In_682);
xnor U1515 (N_1515,N_782,In_1518);
xor U1516 (N_1516,N_1287,N_121);
or U1517 (N_1517,In_336,N_1255);
xnor U1518 (N_1518,N_1077,In_2624);
and U1519 (N_1519,In_144,N_450);
nor U1520 (N_1520,N_600,In_1703);
and U1521 (N_1521,N_1496,N_1456);
nand U1522 (N_1522,In_5,In_2393);
nor U1523 (N_1523,N_1135,N_1172);
nor U1524 (N_1524,In_1213,N_1087);
nor U1525 (N_1525,In_2498,In_256);
xor U1526 (N_1526,N_1022,N_1441);
xnor U1527 (N_1527,In_2166,In_2378);
nor U1528 (N_1528,N_384,In_1490);
nor U1529 (N_1529,N_1113,N_826);
or U1530 (N_1530,In_1933,In_2953);
nand U1531 (N_1531,In_660,In_1259);
nor U1532 (N_1532,N_691,N_1174);
xor U1533 (N_1533,N_1413,In_1456);
xor U1534 (N_1534,N_1436,In_1157);
nand U1535 (N_1535,N_1027,In_2224);
xor U1536 (N_1536,N_93,N_1235);
nor U1537 (N_1537,N_1222,N_693);
or U1538 (N_1538,N_1455,N_207);
nand U1539 (N_1539,In_111,In_63);
nor U1540 (N_1540,In_1235,N_222);
or U1541 (N_1541,N_1045,N_1229);
xnor U1542 (N_1542,N_1420,N_1217);
nor U1543 (N_1543,In_2820,N_673);
or U1544 (N_1544,N_879,N_597);
nor U1545 (N_1545,N_1468,N_513);
nor U1546 (N_1546,In_2077,In_138);
and U1547 (N_1547,N_1344,In_2541);
xor U1548 (N_1548,N_1213,N_1376);
xor U1549 (N_1549,N_1463,N_1365);
or U1550 (N_1550,In_1193,N_218);
xor U1551 (N_1551,N_1120,N_780);
nand U1552 (N_1552,In_1029,In_2823);
nand U1553 (N_1553,N_1053,N_689);
or U1554 (N_1554,In_2265,In_2888);
and U1555 (N_1555,N_663,In_904);
and U1556 (N_1556,In_2708,In_1813);
nand U1557 (N_1557,In_314,In_1653);
or U1558 (N_1558,N_1368,N_537);
and U1559 (N_1559,N_1050,In_2058);
nor U1560 (N_1560,N_1184,In_418);
xor U1561 (N_1561,N_703,N_1173);
and U1562 (N_1562,N_1443,N_314);
and U1563 (N_1563,In_1815,N_963);
nor U1564 (N_1564,N_841,N_1002);
xor U1565 (N_1565,N_696,N_1085);
nand U1566 (N_1566,In_2955,In_1075);
nor U1567 (N_1567,N_72,In_2882);
nor U1568 (N_1568,N_1300,N_853);
nor U1569 (N_1569,N_1116,In_585);
and U1570 (N_1570,In_1248,N_631);
or U1571 (N_1571,N_762,In_1548);
nand U1572 (N_1572,N_1442,In_2680);
xor U1573 (N_1573,In_2070,N_1498);
xnor U1574 (N_1574,N_957,N_233);
and U1575 (N_1575,N_1347,In_1280);
and U1576 (N_1576,N_1469,N_90);
nand U1577 (N_1577,N_1291,In_2437);
or U1578 (N_1578,In_1798,N_492);
or U1579 (N_1579,In_274,N_850);
nand U1580 (N_1580,N_978,N_1335);
and U1581 (N_1581,In_2564,In_712);
and U1582 (N_1582,N_1364,In_2977);
xor U1583 (N_1583,N_908,N_24);
nor U1584 (N_1584,In_330,N_1247);
and U1585 (N_1585,In_1752,In_1623);
and U1586 (N_1586,In_1288,In_2996);
nand U1587 (N_1587,In_701,N_140);
xor U1588 (N_1588,N_1169,In_2219);
xor U1589 (N_1589,N_119,In_1861);
nand U1590 (N_1590,In_59,In_508);
nor U1591 (N_1591,N_1138,N_1266);
or U1592 (N_1592,N_1351,In_1830);
nand U1593 (N_1593,N_718,In_693);
xnor U1594 (N_1594,N_1313,N_1471);
or U1595 (N_1595,N_1190,N_1063);
nand U1596 (N_1596,In_2948,N_1261);
xnor U1597 (N_1597,In_161,N_1282);
xnor U1598 (N_1598,In_1559,N_1398);
xor U1599 (N_1599,In_2016,N_323);
and U1600 (N_1600,In_1249,N_1497);
nand U1601 (N_1601,N_1267,In_2364);
or U1602 (N_1602,In_2921,N_453);
nor U1603 (N_1603,N_1476,In_348);
and U1604 (N_1604,N_1086,N_1195);
nor U1605 (N_1605,N_1387,In_1767);
and U1606 (N_1606,N_1165,N_431);
and U1607 (N_1607,N_304,In_1027);
or U1608 (N_1608,N_757,N_921);
and U1609 (N_1609,In_2067,N_35);
nand U1610 (N_1610,In_1874,In_2030);
or U1611 (N_1611,N_1484,N_1345);
xnor U1612 (N_1612,In_1896,In_661);
nand U1613 (N_1613,N_844,N_814);
or U1614 (N_1614,In_578,In_743);
xor U1615 (N_1615,In_2824,N_1350);
xor U1616 (N_1616,N_257,N_1249);
nor U1617 (N_1617,N_1487,In_1339);
xnor U1618 (N_1618,N_442,N_136);
or U1619 (N_1619,In_169,In_2608);
or U1620 (N_1620,In_1750,In_2763);
and U1621 (N_1621,In_87,In_2861);
and U1622 (N_1622,N_1105,In_1523);
or U1623 (N_1623,N_951,In_2864);
or U1624 (N_1624,N_524,N_1379);
xnor U1625 (N_1625,In_2952,N_1052);
nor U1626 (N_1626,N_372,N_947);
xor U1627 (N_1627,In_1309,N_1098);
xor U1628 (N_1628,N_1481,N_1417);
nor U1629 (N_1629,In_2053,In_1312);
nand U1630 (N_1630,N_1205,N_1349);
xor U1631 (N_1631,N_1435,In_771);
xor U1632 (N_1632,N_1357,N_1355);
or U1633 (N_1633,N_1041,N_469);
xnor U1634 (N_1634,In_1422,In_1644);
nor U1635 (N_1635,In_513,In_1204);
and U1636 (N_1636,N_1253,N_1360);
xnor U1637 (N_1637,In_2893,N_1094);
or U1638 (N_1638,N_138,N_1114);
or U1639 (N_1639,N_1112,N_564);
nand U1640 (N_1640,In_1645,In_1917);
and U1641 (N_1641,N_392,In_1832);
nand U1642 (N_1642,N_735,N_633);
xnor U1643 (N_1643,N_1219,N_290);
or U1644 (N_1644,In_1690,N_1307);
xor U1645 (N_1645,In_60,In_1495);
xor U1646 (N_1646,N_943,In_2347);
xor U1647 (N_1647,N_380,In_1574);
and U1648 (N_1648,In_1285,In_1151);
nor U1649 (N_1649,N_1446,N_1012);
nor U1650 (N_1650,N_531,In_1458);
xor U1651 (N_1651,In_2892,In_1480);
and U1652 (N_1652,In_1296,N_578);
nor U1653 (N_1653,N_975,N_1148);
and U1654 (N_1654,In_2277,N_1367);
nand U1655 (N_1655,In_1024,N_573);
nor U1656 (N_1656,N_579,In_61);
nand U1657 (N_1657,N_1143,In_178);
nand U1658 (N_1658,N_965,In_2117);
nand U1659 (N_1659,In_541,In_2698);
nor U1660 (N_1660,N_1483,N_636);
or U1661 (N_1661,In_1314,In_1976);
xor U1662 (N_1662,In_307,N_925);
or U1663 (N_1663,N_1464,In_2487);
and U1664 (N_1664,In_657,N_833);
nor U1665 (N_1665,N_740,In_286);
nand U1666 (N_1666,N_1251,N_459);
nand U1667 (N_1667,In_925,In_1220);
nor U1668 (N_1668,N_1128,In_2716);
nor U1669 (N_1669,In_885,In_1553);
and U1670 (N_1670,N_1421,In_2650);
xor U1671 (N_1671,N_391,N_1068);
nand U1672 (N_1672,In_89,N_637);
nand U1673 (N_1673,N_1166,N_672);
nor U1674 (N_1674,In_2709,In_2403);
nor U1675 (N_1675,In_292,N_1200);
and U1676 (N_1676,In_1232,In_1520);
and U1677 (N_1677,In_906,N_249);
nor U1678 (N_1678,In_477,In_2490);
nand U1679 (N_1679,In_947,In_1509);
or U1680 (N_1680,N_765,In_172);
xnor U1681 (N_1681,N_1258,In_2973);
nor U1682 (N_1682,In_673,N_1170);
nor U1683 (N_1683,N_1099,In_1141);
nor U1684 (N_1684,N_1466,N_51);
and U1685 (N_1685,N_1163,N_1273);
or U1686 (N_1686,N_1202,N_451);
or U1687 (N_1687,In_757,In_1319);
or U1688 (N_1688,In_901,N_396);
and U1689 (N_1689,N_1059,In_2898);
and U1690 (N_1690,In_2710,In_2965);
nand U1691 (N_1691,In_2651,In_1626);
xor U1692 (N_1692,In_1778,N_802);
and U1693 (N_1693,In_1452,N_1378);
nand U1694 (N_1694,N_28,In_2221);
and U1695 (N_1695,In_691,N_1119);
or U1696 (N_1696,N_1269,In_2830);
nand U1697 (N_1697,N_1288,N_969);
nand U1698 (N_1698,In_1761,N_893);
xor U1699 (N_1699,N_529,In_2460);
xnor U1700 (N_1700,N_1066,In_1369);
nor U1701 (N_1701,N_1211,N_1397);
nor U1702 (N_1702,N_1333,N_1391);
or U1703 (N_1703,In_2458,In_1147);
and U1704 (N_1704,N_1248,In_1154);
and U1705 (N_1705,In_1287,N_1458);
nand U1706 (N_1706,In_1980,N_1321);
or U1707 (N_1707,N_1416,In_469);
nand U1708 (N_1708,N_1141,In_2616);
nor U1709 (N_1709,N_339,In_1566);
nand U1710 (N_1710,N_1450,N_230);
and U1711 (N_1711,In_2314,In_1923);
xor U1712 (N_1712,N_1192,N_845);
nor U1713 (N_1713,In_1741,N_504);
nor U1714 (N_1714,N_699,N_1366);
xnor U1715 (N_1715,N_1069,N_364);
or U1716 (N_1716,N_710,N_1106);
or U1717 (N_1717,N_1126,N_179);
nand U1718 (N_1718,N_1438,N_1204);
nor U1719 (N_1719,N_1459,In_2852);
nand U1720 (N_1720,N_1154,In_1536);
and U1721 (N_1721,N_1406,N_1244);
nor U1722 (N_1722,In_2326,In_363);
or U1723 (N_1723,N_619,In_1175);
xor U1724 (N_1724,In_1282,N_1024);
nor U1725 (N_1725,N_308,In_662);
or U1726 (N_1726,In_530,In_2427);
and U1727 (N_1727,N_1100,N_1134);
xnor U1728 (N_1728,N_1036,N_869);
xor U1729 (N_1729,N_1276,In_2607);
xnor U1730 (N_1730,In_735,In_1439);
nand U1731 (N_1731,In_1395,In_1246);
or U1732 (N_1732,N_1315,In_2065);
and U1733 (N_1733,In_2905,N_880);
nor U1734 (N_1734,In_1361,In_2545);
and U1735 (N_1735,In_2866,N_1326);
nor U1736 (N_1736,In_834,N_1254);
and U1737 (N_1737,N_496,N_277);
or U1738 (N_1738,N_215,N_554);
or U1739 (N_1739,N_829,In_1008);
nand U1740 (N_1740,N_1312,N_448);
nand U1741 (N_1741,N_1109,N_1359);
or U1742 (N_1742,N_1203,N_1156);
or U1743 (N_1743,N_669,N_1445);
nor U1744 (N_1744,In_1474,In_221);
nand U1745 (N_1745,N_1225,In_2411);
or U1746 (N_1746,In_1670,In_1575);
and U1747 (N_1747,In_791,In_1844);
nor U1748 (N_1748,In_1304,N_55);
xnor U1749 (N_1749,N_671,N_1241);
xor U1750 (N_1750,In_373,N_1189);
or U1751 (N_1751,N_124,N_611);
or U1752 (N_1752,In_943,N_614);
and U1753 (N_1753,N_628,In_325);
nand U1754 (N_1754,N_1084,N_1305);
nand U1755 (N_1755,In_2414,In_635);
nand U1756 (N_1756,In_2507,In_1912);
or U1757 (N_1757,N_1444,In_333);
nand U1758 (N_1758,In_2665,In_1918);
and U1759 (N_1759,In_2621,In_2229);
and U1760 (N_1760,In_2469,N_1475);
xor U1761 (N_1761,N_1304,N_904);
and U1762 (N_1762,In_2692,N_1299);
nor U1763 (N_1763,N_876,N_766);
nand U1764 (N_1764,N_1216,N_944);
nor U1765 (N_1765,N_1081,N_132);
xnor U1766 (N_1766,N_1310,N_1331);
or U1767 (N_1767,In_245,In_1919);
or U1768 (N_1768,N_752,In_2308);
and U1769 (N_1769,In_1963,In_2296);
nand U1770 (N_1770,In_2570,N_1412);
and U1771 (N_1771,In_1498,N_1199);
or U1772 (N_1772,N_838,N_317);
and U1773 (N_1773,In_412,In_1363);
and U1774 (N_1774,In_1515,N_475);
or U1775 (N_1775,In_2687,N_808);
and U1776 (N_1776,N_71,In_2144);
and U1777 (N_1777,N_371,N_361);
xnor U1778 (N_1778,In_1311,N_395);
nand U1779 (N_1779,N_1293,In_1187);
or U1780 (N_1780,N_889,In_1424);
and U1781 (N_1781,N_846,In_1989);
nor U1782 (N_1782,N_403,N_1329);
and U1783 (N_1783,N_1123,In_1812);
or U1784 (N_1784,N_190,In_2850);
and U1785 (N_1785,N_1494,N_1488);
nor U1786 (N_1786,In_702,N_286);
nand U1787 (N_1787,N_1096,In_2291);
nand U1788 (N_1788,In_1530,In_1211);
nor U1789 (N_1789,N_147,N_366);
and U1790 (N_1790,In_1380,N_202);
or U1791 (N_1791,N_1139,In_2050);
or U1792 (N_1792,In_2121,In_981);
nor U1793 (N_1793,N_1390,In_263);
nand U1794 (N_1794,N_1415,N_279);
and U1795 (N_1795,N_881,N_1402);
or U1796 (N_1796,In_785,N_771);
or U1797 (N_1797,In_1708,N_594);
and U1798 (N_1798,N_622,N_1262);
xnor U1799 (N_1799,N_1194,In_1045);
nand U1800 (N_1800,In_1137,N_1792);
xor U1801 (N_1801,In_1415,In_369);
xor U1802 (N_1802,N_404,N_1233);
or U1803 (N_1803,In_1398,N_1779);
nand U1804 (N_1804,N_1049,N_1673);
nor U1805 (N_1805,N_1284,In_2847);
or U1806 (N_1806,In_1791,N_1095);
and U1807 (N_1807,N_271,In_554);
xor U1808 (N_1808,In_2462,N_1252);
or U1809 (N_1809,In_2245,N_1452);
nor U1810 (N_1810,N_1396,N_260);
xor U1811 (N_1811,N_1394,N_1728);
and U1812 (N_1812,N_1669,N_858);
xnor U1813 (N_1813,In_2152,N_1401);
or U1814 (N_1814,N_1479,In_1660);
xnor U1815 (N_1815,N_1731,N_1573);
and U1816 (N_1816,N_1523,In_2925);
and U1817 (N_1817,In_171,N_438);
nor U1818 (N_1818,In_420,N_107);
nand U1819 (N_1819,N_884,N_1206);
or U1820 (N_1820,N_1389,In_1300);
xnor U1821 (N_1821,N_1670,In_340);
or U1822 (N_1822,N_1755,In_759);
xnor U1823 (N_1823,N_1652,N_650);
and U1824 (N_1824,In_561,In_589);
nand U1825 (N_1825,N_1533,In_740);
and U1826 (N_1826,In_1400,N_1374);
nand U1827 (N_1827,N_809,In_817);
nor U1828 (N_1828,N_1210,N_736);
nor U1829 (N_1829,In_2656,In_2355);
nor U1830 (N_1830,In_1057,N_1734);
and U1831 (N_1831,N_1514,N_1770);
or U1832 (N_1832,N_848,In_754);
xnor U1833 (N_1833,N_1188,In_2160);
nand U1834 (N_1834,N_1791,N_1794);
and U1835 (N_1835,In_1828,N_1302);
nand U1836 (N_1836,In_2315,In_490);
and U1837 (N_1837,In_1633,N_1597);
xor U1838 (N_1838,N_1090,N_1457);
nand U1839 (N_1839,N_1624,N_1623);
nor U1840 (N_1840,N_831,In_1596);
or U1841 (N_1841,In_1954,N_1362);
nand U1842 (N_1842,N_1622,In_1822);
or U1843 (N_1843,N_1716,N_1545);
or U1844 (N_1844,In_1001,In_124);
nor U1845 (N_1845,In_1801,In_927);
xnor U1846 (N_1846,N_328,N_411);
nor U1847 (N_1847,N_410,N_772);
nand U1848 (N_1848,In_1522,N_1593);
nor U1849 (N_1849,N_1619,In_2195);
nor U1850 (N_1850,N_1528,N_1711);
or U1851 (N_1851,N_1550,N_1182);
xor U1852 (N_1852,In_894,N_973);
or U1853 (N_1853,In_2630,N_1474);
nor U1854 (N_1854,N_1117,N_1263);
xnor U1855 (N_1855,In_365,In_1503);
xnor U1856 (N_1856,N_1574,N_1317);
xnor U1857 (N_1857,N_1684,N_194);
nor U1858 (N_1858,In_1430,In_2903);
nand U1859 (N_1859,N_1308,N_934);
nor U1860 (N_1860,In_651,N_1043);
xor U1861 (N_1861,In_1851,In_1873);
or U1862 (N_1862,In_2664,N_1664);
nor U1863 (N_1863,N_1715,In_2858);
and U1864 (N_1864,In_145,In_1033);
nor U1865 (N_1865,N_414,N_1603);
nand U1866 (N_1866,In_345,In_2122);
xnor U1867 (N_1867,N_1736,In_1233);
nand U1868 (N_1868,N_1517,N_742);
nor U1869 (N_1869,N_1020,N_815);
nor U1870 (N_1870,N_1554,N_1316);
xnor U1871 (N_1871,In_1697,N_1680);
and U1872 (N_1872,N_1692,N_1482);
and U1873 (N_1873,N_1384,N_509);
or U1874 (N_1874,In_93,N_1453);
nor U1875 (N_1875,N_311,N_1493);
and U1876 (N_1876,N_1581,In_2677);
nor U1877 (N_1877,In_2264,In_1077);
xnor U1878 (N_1878,N_1538,In_2259);
nor U1879 (N_1879,N_1592,N_365);
xnor U1880 (N_1880,N_1589,N_446);
nand U1881 (N_1881,In_889,In_1250);
or U1882 (N_1882,N_1682,In_1255);
nand U1883 (N_1883,In_219,N_1607);
xor U1884 (N_1884,In_2238,In_1737);
or U1885 (N_1885,In_255,N_1314);
nand U1886 (N_1886,N_455,N_1558);
and U1887 (N_1887,N_1672,N_1334);
or U1888 (N_1888,N_150,N_1646);
xnor U1889 (N_1889,In_2408,N_1275);
or U1890 (N_1890,N_721,N_1051);
and U1891 (N_1891,N_1201,N_982);
or U1892 (N_1892,N_1512,N_1260);
and U1893 (N_1893,N_1578,N_795);
xor U1894 (N_1894,N_325,N_1289);
xnor U1895 (N_1895,N_1358,N_1691);
and U1896 (N_1896,N_792,N_1245);
or U1897 (N_1897,In_2932,N_1555);
or U1898 (N_1898,In_1556,N_1242);
and U1899 (N_1899,In_1128,N_972);
nor U1900 (N_1900,N_1566,N_1013);
nand U1901 (N_1901,In_1379,N_1093);
xor U1902 (N_1902,In_2781,In_1747);
nor U1903 (N_1903,N_1230,N_1510);
or U1904 (N_1904,N_1626,N_68);
and U1905 (N_1905,N_1294,In_2826);
xnor U1906 (N_1906,N_1681,N_556);
nor U1907 (N_1907,N_69,N_1576);
nand U1908 (N_1908,N_447,N_1658);
or U1909 (N_1909,In_2594,In_1454);
and U1910 (N_1910,N_1695,In_748);
nand U1911 (N_1911,N_1577,N_1186);
and U1912 (N_1912,N_270,N_816);
nand U1913 (N_1913,In_1373,N_1409);
nand U1914 (N_1914,N_1635,N_989);
and U1915 (N_1915,In_1342,N_1764);
or U1916 (N_1916,N_1552,In_1949);
nand U1917 (N_1917,In_213,N_1381);
and U1918 (N_1918,N_1103,In_2722);
nor U1919 (N_1919,In_2627,In_445);
nor U1920 (N_1920,N_1704,N_1636);
or U1921 (N_1921,N_716,In_1399);
xor U1922 (N_1922,In_2613,N_909);
xnor U1923 (N_1923,N_1585,N_166);
nor U1924 (N_1924,N_1587,N_1477);
nand U1925 (N_1925,N_1580,In_300);
xor U1926 (N_1926,N_1214,N_196);
nand U1927 (N_1927,N_1506,N_1354);
xnor U1928 (N_1928,In_731,N_1608);
xnor U1929 (N_1929,N_1383,In_62);
and U1930 (N_1930,N_1648,N_1789);
xnor U1931 (N_1931,N_1525,N_1583);
and U1932 (N_1932,In_2499,N_791);
and U1933 (N_1933,N_1687,N_1318);
or U1934 (N_1934,In_1055,N_1407);
nor U1935 (N_1935,In_1837,N_1616);
nand U1936 (N_1936,N_1429,N_1797);
nand U1937 (N_1937,N_1600,In_2092);
nor U1938 (N_1938,N_1215,In_2816);
nor U1939 (N_1939,N_1604,N_1238);
nor U1940 (N_1940,N_104,In_2292);
and U1941 (N_1941,N_1787,N_193);
or U1942 (N_1942,N_1752,N_605);
nor U1943 (N_1943,In_1050,In_1621);
xnor U1944 (N_1944,N_662,N_1257);
or U1945 (N_1945,In_2994,N_1678);
nand U1946 (N_1946,N_1208,In_749);
nand U1947 (N_1947,N_505,In_1168);
nor U1948 (N_1948,N_1642,N_1428);
xor U1949 (N_1949,In_294,N_1564);
or U1950 (N_1950,N_1788,N_1741);
xnor U1951 (N_1951,In_1528,N_1671);
or U1952 (N_1952,In_30,N_933);
xor U1953 (N_1953,N_1072,N_1584);
xnor U1954 (N_1954,In_2625,In_198);
nand U1955 (N_1955,N_1614,In_573);
nand U1956 (N_1956,N_73,N_1693);
nor U1957 (N_1957,In_2899,N_1615);
xor U1958 (N_1958,N_545,In_2474);
and U1959 (N_1959,In_621,N_1071);
nor U1960 (N_1960,In_241,N_823);
or U1961 (N_1961,N_1056,N_1515);
or U1962 (N_1962,N_825,N_1183);
and U1963 (N_1963,In_1252,N_1675);
nand U1964 (N_1964,N_1239,N_502);
and U1965 (N_1965,In_2619,In_2728);
xor U1966 (N_1966,In_1784,In_2568);
and U1967 (N_1967,N_558,In_1924);
xnor U1968 (N_1968,In_2566,N_686);
or U1969 (N_1969,N_1423,N_377);
or U1970 (N_1970,In_614,In_2726);
nand U1971 (N_1971,N_1618,N_1611);
nor U1972 (N_1972,N_1388,In_283);
xnor U1973 (N_1973,N_946,In_1908);
nor U1974 (N_1974,N_188,N_1509);
and U1975 (N_1975,In_2843,N_1155);
xnor U1976 (N_1976,In_2649,In_391);
or U1977 (N_1977,N_1586,In_1676);
nor U1978 (N_1978,N_682,N_1026);
nor U1979 (N_1979,N_1270,N_385);
xor U1980 (N_1980,In_1991,N_1460);
nand U1981 (N_1981,N_738,N_991);
xnor U1982 (N_1982,N_1410,N_1320);
nor U1983 (N_1983,N_1724,N_274);
nand U1984 (N_1984,In_679,N_745);
nand U1985 (N_1985,In_1673,In_715);
or U1986 (N_1986,N_775,N_1370);
or U1987 (N_1987,N_1224,N_1040);
nand U1988 (N_1988,N_577,N_1432);
and U1989 (N_1989,N_935,N_1111);
xor U1990 (N_1990,N_1057,N_595);
or U1991 (N_1991,N_536,N_681);
nor U1992 (N_1992,N_1562,N_1649);
and U1993 (N_1993,In_100,N_1490);
nand U1994 (N_1994,In_2114,N_1010);
and U1995 (N_1995,N_1110,In_2148);
and U1996 (N_1996,In_2396,In_1016);
nor U1997 (N_1997,In_956,N_1274);
nor U1998 (N_1998,N_911,N_1557);
or U1999 (N_1999,In_1810,N_981);
or U2000 (N_2000,N_1757,In_2301);
xnor U2001 (N_2001,N_1547,N_1746);
nor U2002 (N_2002,N_1793,N_305);
xnor U2003 (N_2003,In_1544,N_1480);
or U2004 (N_2004,N_1234,N_1240);
and U2005 (N_2005,N_1372,In_2706);
nor U2006 (N_2006,In_1720,In_1298);
nand U2007 (N_2007,N_1567,In_128);
or U2008 (N_2008,In_1222,In_1744);
nor U2009 (N_2009,In_380,In_1040);
or U2010 (N_2010,N_285,N_1283);
or U2011 (N_2011,N_1754,N_1651);
nor U2012 (N_2012,In_1005,N_1532);
and U2013 (N_2013,N_1582,In_1160);
nand U2014 (N_2014,N_899,N_1061);
and U2015 (N_2015,N_1575,N_1414);
nand U2016 (N_2016,In_2675,N_996);
and U2017 (N_2017,N_612,In_1884);
nand U2018 (N_2018,In_1957,N_1590);
or U2019 (N_2019,N_1014,N_770);
or U2020 (N_2020,N_1633,N_1323);
nor U2021 (N_2021,N_1766,N_337);
nor U2022 (N_2022,N_593,N_1029);
nand U2023 (N_2023,N_1246,N_800);
nand U2024 (N_2024,N_1076,N_895);
nor U2025 (N_2025,In_1082,In_1506);
nand U2026 (N_2026,In_488,N_1403);
nor U2027 (N_2027,N_236,In_1048);
nor U2028 (N_2028,In_1143,N_1655);
or U2029 (N_2029,In_2790,N_1382);
xor U2030 (N_2030,In_2358,N_1422);
or U2031 (N_2031,N_1303,N_670);
nand U2032 (N_2032,N_1679,N_768);
nand U2033 (N_2033,In_619,In_568);
and U2034 (N_2034,N_1454,N_725);
nand U2035 (N_2035,N_1579,N_1196);
or U2036 (N_2036,N_528,N_1009);
and U2037 (N_2037,N_1676,In_1360);
xor U2038 (N_2038,N_1781,In_778);
xor U2039 (N_2039,N_1718,In_974);
nand U2040 (N_2040,N_1361,N_538);
and U2041 (N_2041,N_793,N_950);
nand U2042 (N_2042,N_1773,N_617);
nand U2043 (N_2043,In_72,N_694);
nand U2044 (N_2044,N_1426,N_1209);
nor U2045 (N_2045,N_700,N_487);
and U2046 (N_2046,N_1227,N_1259);
xnor U2047 (N_2047,In_2175,In_1582);
or U2048 (N_2048,N_53,N_1124);
xor U2049 (N_2049,N_1404,N_1501);
or U2050 (N_2050,N_1690,N_1104);
and U2051 (N_2051,N_827,In_2671);
xor U2052 (N_2052,In_1661,In_486);
nor U2053 (N_2053,N_1527,In_2306);
nand U2054 (N_2054,In_2124,N_656);
or U2055 (N_2055,N_607,N_1758);
nor U2056 (N_2056,N_1047,N_690);
xor U2057 (N_2057,N_1434,In_2068);
and U2058 (N_2058,N_1601,In_840);
nor U2059 (N_2059,N_596,N_1627);
and U2060 (N_2060,N_1546,N_1572);
nor U2061 (N_2061,N_423,N_1540);
xnor U2062 (N_2062,N_1491,N_1145);
or U2063 (N_2063,N_1427,N_1521);
nand U2064 (N_2064,N_1786,In_2139);
or U2065 (N_2065,In_298,N_1720);
nor U2066 (N_2066,N_1553,In_2311);
and U2067 (N_2067,N_268,N_1748);
or U2068 (N_2068,N_581,N_709);
nor U2069 (N_2069,N_1265,In_148);
and U2070 (N_2070,N_864,In_1701);
xor U2071 (N_2071,N_1000,In_1680);
nand U2072 (N_2072,N_1236,N_1701);
and U2073 (N_2073,N_1700,N_1131);
xor U2074 (N_2074,In_988,N_1534);
nor U2075 (N_2075,In_2281,In_465);
nand U2076 (N_2076,In_1516,N_954);
or U2077 (N_2077,N_1689,In_2024);
and U2078 (N_2078,N_724,N_1462);
xor U2079 (N_2079,In_7,N_897);
or U2080 (N_2080,N_1727,N_1686);
xnor U2081 (N_2081,N_1461,In_2348);
or U2082 (N_2082,N_1631,In_598);
xor U2083 (N_2083,N_1001,N_616);
or U2084 (N_2084,N_999,N_754);
nand U2085 (N_2085,In_687,N_1017);
nor U2086 (N_2086,In_2984,N_1272);
and U2087 (N_2087,N_1765,In_2174);
nor U2088 (N_2088,N_1243,N_1264);
and U2089 (N_2089,N_1588,In_1212);
or U2090 (N_2090,In_1818,N_1723);
xnor U2091 (N_2091,In_2904,N_1743);
and U2092 (N_2092,N_839,N_1025);
nand U2093 (N_2093,In_2628,In_2922);
or U2094 (N_2094,N_1035,N_572);
nor U2095 (N_2095,N_1760,N_503);
nor U2096 (N_2096,In_1696,N_638);
nand U2097 (N_2097,N_604,In_2595);
xor U2098 (N_2098,In_1475,N_1430);
xor U2099 (N_2099,In_2839,N_613);
nor U2100 (N_2100,N_1825,In_375);
or U2101 (N_2101,In_1729,N_1037);
and U2102 (N_2102,N_1279,N_1726);
xnor U2103 (N_2103,In_2455,In_2659);
nor U2104 (N_2104,N_2025,N_1898);
nor U2105 (N_2105,N_1800,N_1160);
or U2106 (N_2106,N_1978,N_1767);
xor U2107 (N_2107,N_1660,N_342);
xnor U2108 (N_2108,N_1939,In_1672);
and U2109 (N_2109,N_1778,N_2077);
xnor U2110 (N_2110,N_1993,N_2095);
nand U2111 (N_2111,N_1994,N_1725);
or U2112 (N_2112,N_1883,N_1911);
nand U2113 (N_2113,N_283,N_2054);
and U2114 (N_2114,N_1817,In_964);
nand U2115 (N_2115,N_875,N_1844);
nand U2116 (N_2116,N_1336,N_1865);
and U2117 (N_2117,In_1072,N_1495);
nand U2118 (N_2118,In_421,N_2099);
nand U2119 (N_2119,N_887,N_959);
and U2120 (N_2120,N_1296,N_1418);
and U2121 (N_2121,N_1280,N_1796);
or U2122 (N_2122,N_905,N_38);
xnor U2123 (N_2123,In_2742,N_1903);
nor U2124 (N_2124,N_2030,In_847);
and U2125 (N_2125,N_1891,In_2648);
or U2126 (N_2126,N_2069,N_2086);
nand U2127 (N_2127,N_2027,In_1636);
xor U2128 (N_2128,N_1985,N_1940);
or U2129 (N_2129,In_1513,N_2084);
nor U2130 (N_2130,In_2423,N_1226);
or U2131 (N_2131,N_1568,N_1371);
nor U2132 (N_2132,In_1500,N_2022);
nor U2133 (N_2133,N_1870,In_915);
xnor U2134 (N_2134,N_2067,N_667);
and U2135 (N_2135,N_1972,N_998);
and U2136 (N_2136,N_1395,N_967);
or U2137 (N_2137,In_2822,N_1879);
or U2138 (N_2138,In_1594,N_139);
nand U2139 (N_2139,In_106,In_2078);
and U2140 (N_2140,N_1089,In_2547);
nor U2141 (N_2141,N_1161,In_1835);
xor U2142 (N_2142,N_924,N_1625);
or U2143 (N_2143,N_2014,N_1620);
xor U2144 (N_2144,N_2065,N_1888);
and U2145 (N_2145,In_1402,N_1070);
nor U2146 (N_2146,N_1889,N_1685);
nand U2147 (N_2147,N_1892,N_1657);
and U2148 (N_2148,N_1425,N_1223);
nor U2149 (N_2149,N_1846,N_896);
nand U2150 (N_2150,N_1768,N_1730);
and U2151 (N_2151,N_331,N_1212);
or U2152 (N_2152,N_1630,N_1740);
or U2153 (N_2153,N_540,N_871);
and U2154 (N_2154,N_1941,N_863);
nand U2155 (N_2155,N_1271,N_1543);
or U2156 (N_2156,N_2003,In_1407);
nor U2157 (N_2157,N_1197,N_1176);
xnor U2158 (N_2158,N_334,N_962);
or U2159 (N_2159,In_1411,N_1489);
or U2160 (N_2160,In_750,In_1326);
nand U2161 (N_2161,N_1924,N_1617);
nand U2162 (N_2162,N_958,In_863);
and U2163 (N_2163,N_1448,In_2909);
and U2164 (N_2164,In_2505,N_1744);
nor U2165 (N_2165,N_2032,N_1309);
nand U2166 (N_2166,In_233,In_1117);
nor U2167 (N_2167,N_1500,N_1824);
and U2168 (N_2168,In_856,N_1845);
xnor U2169 (N_2169,In_2407,N_2066);
nand U2170 (N_2170,In_2069,In_41);
nor U2171 (N_2171,N_1850,In_45);
or U2172 (N_2172,N_922,N_1228);
nor U2173 (N_2173,N_1842,N_1136);
nor U2174 (N_2174,N_1854,N_1717);
and U2175 (N_2175,N_1877,N_2010);
and U2176 (N_2176,N_1918,N_1707);
or U2177 (N_2177,N_788,N_1551);
nor U2178 (N_2178,N_1602,In_1420);
and U2179 (N_2179,In_1651,In_417);
and U2180 (N_2180,In_1297,N_1544);
xor U2181 (N_2181,N_1714,N_2000);
nor U2182 (N_2182,N_584,N_2090);
or U2183 (N_2183,N_974,In_2561);
xnor U2184 (N_2184,N_779,In_607);
nand U2185 (N_2185,N_977,N_852);
nor U2186 (N_2186,N_1956,In_2461);
or U2187 (N_2187,N_417,In_1511);
xnor U2188 (N_2188,In_1637,N_94);
and U2189 (N_2189,N_1769,N_1946);
or U2190 (N_2190,N_1465,N_900);
or U2191 (N_2191,N_1542,N_1995);
nor U2192 (N_2192,In_177,N_2001);
nor U2193 (N_2193,N_1772,N_1999);
or U2194 (N_2194,N_1876,In_2879);
or U2195 (N_2195,In_2346,N_1832);
xnor U2196 (N_2196,N_1836,N_1812);
or U2197 (N_2197,N_1221,N_1080);
nor U2198 (N_2198,N_1881,N_1899);
nor U2199 (N_2199,N_1900,N_915);
or U2200 (N_2200,N_1840,N_1118);
xnor U2201 (N_2201,N_1902,N_1996);
nor U2202 (N_2202,N_968,N_1713);
xor U2203 (N_2203,N_1277,N_302);
nand U2204 (N_2204,N_1613,N_2041);
and U2205 (N_2205,In_1827,N_2059);
and U2206 (N_2206,N_2033,N_1609);
nand U2207 (N_2207,In_1753,N_1815);
nor U2208 (N_2208,N_666,In_1459);
or U2209 (N_2209,N_1231,N_1751);
or U2210 (N_2210,N_1847,N_1386);
nor U2211 (N_2211,N_1439,N_1920);
nand U2212 (N_2212,N_1019,N_1322);
xnor U2213 (N_2213,N_1864,N_1187);
xnor U2214 (N_2214,N_108,In_278);
or U2215 (N_2215,N_1831,N_644);
nor U2216 (N_2216,N_819,N_953);
xor U2217 (N_2217,N_2058,N_1638);
nand U2218 (N_2218,N_2028,N_1522);
xnor U2219 (N_2219,N_1935,N_1640);
nor U2220 (N_2220,N_2006,N_1505);
xnor U2221 (N_2221,N_1091,N_2018);
and U2222 (N_2222,N_1571,N_1774);
xnor U2223 (N_2223,N_1703,N_1708);
or U2224 (N_2224,N_1833,N_1803);
and U2225 (N_2225,N_146,N_2064);
nor U2226 (N_2226,N_200,N_1340);
nand U2227 (N_2227,In_2484,N_1777);
and U2228 (N_2228,N_1656,N_926);
or U2229 (N_2229,N_1369,N_1157);
nor U2230 (N_2230,In_703,In_2085);
and U2231 (N_2231,N_1997,In_920);
and U2232 (N_2232,In_922,N_1869);
and U2233 (N_2233,N_2085,N_1915);
nor U2234 (N_2234,N_1775,N_761);
nand U2235 (N_2235,In_290,N_2051);
xor U2236 (N_2236,In_1754,N_1712);
nand U2237 (N_2237,N_1218,N_1424);
nand U2238 (N_2238,N_2087,N_2092);
nor U2239 (N_2239,N_1702,N_928);
xnor U2240 (N_2240,N_1268,N_1560);
or U2241 (N_2241,N_2053,N_1868);
nor U2242 (N_2242,N_1771,N_1810);
or U2243 (N_2243,N_1882,N_2088);
nand U2244 (N_2244,N_907,N_1776);
or U2245 (N_2245,N_1922,N_1809);
or U2246 (N_2246,In_360,N_956);
nor U2247 (N_2247,N_1629,N_1983);
and U2248 (N_2248,N_1598,N_1802);
nor U2249 (N_2249,In_2797,In_2992);
or U2250 (N_2250,N_1122,N_1986);
xnor U2251 (N_2251,N_1659,N_2073);
xor U2252 (N_2252,N_1950,N_1818);
nand U2253 (N_2253,N_1433,N_860);
nor U2254 (N_2254,N_1286,N_1440);
and U2255 (N_2255,In_1647,N_1549);
nand U2256 (N_2256,N_1873,N_1859);
nor U2257 (N_2257,N_1508,N_1867);
xor U2258 (N_2258,N_1694,N_386);
nand U2259 (N_2259,N_2016,N_2011);
and U2260 (N_2260,N_374,N_715);
xor U2261 (N_2261,N_1292,N_1529);
and U2262 (N_2262,In_416,In_2421);
nor U2263 (N_2263,N_252,N_1356);
or U2264 (N_2264,N_1662,N_1934);
nand U2265 (N_2265,N_1807,N_1851);
nor U2266 (N_2266,N_960,N_1153);
xor U2267 (N_2267,N_1565,N_1298);
nor U2268 (N_2268,In_1978,N_1060);
or U2269 (N_2269,N_635,N_2043);
and U2270 (N_2270,N_1628,In_1725);
and U2271 (N_2271,In_907,N_1874);
nor U2272 (N_2272,In_1939,N_940);
or U2273 (N_2273,N_1949,N_1431);
or U2274 (N_2274,N_1951,N_307);
or U2275 (N_2275,N_1937,In_2935);
or U2276 (N_2276,In_1722,N_1722);
nand U2277 (N_2277,N_1909,N_1805);
and U2278 (N_2278,In_788,N_744);
xnor U2279 (N_2279,N_2049,In_497);
or U2280 (N_2280,N_1175,In_2226);
nand U2281 (N_2281,N_1699,N_2050);
xor U2282 (N_2282,N_1830,In_2736);
nand U2283 (N_2283,N_2072,In_2351);
nand U2284 (N_2284,N_1897,N_1856);
nor U2285 (N_2285,N_2004,N_86);
and U2286 (N_2286,N_2002,N_1826);
xor U2287 (N_2287,N_1127,In_1571);
nor U2288 (N_2288,N_1346,N_2097);
nor U2289 (N_2289,N_877,N_1929);
xnor U2290 (N_2290,N_2015,N_1666);
or U2291 (N_2291,In_2855,N_1977);
nand U2292 (N_2292,N_1894,In_2149);
and U2293 (N_2293,N_1606,N_1790);
nand U2294 (N_2294,In_24,N_1732);
and U2295 (N_2295,N_1804,In_710);
xnor U2296 (N_2296,N_1377,N_2045);
nand U2297 (N_2297,In_2127,N_2047);
xnor U2298 (N_2298,N_1955,N_1973);
and U2299 (N_2299,N_1981,N_2031);
and U2300 (N_2300,N_1393,N_2019);
or U2301 (N_2301,N_1337,N_1643);
or U2302 (N_2302,N_1871,N_1814);
or U2303 (N_2303,N_2012,N_1875);
and U2304 (N_2304,In_384,N_402);
or U2305 (N_2305,N_1976,In_2060);
nor U2306 (N_2306,N_1896,N_1989);
xnor U2307 (N_2307,N_1599,N_1785);
nor U2308 (N_2308,N_1964,N_2096);
nand U2309 (N_2309,N_1518,In_2275);
and U2310 (N_2310,In_838,N_1795);
or U2311 (N_2311,N_1539,In_2390);
xor U2312 (N_2312,N_1605,N_393);
and U2313 (N_2313,N_1967,N_1531);
and U2314 (N_2314,N_1537,N_1841);
nand U2315 (N_2315,In_1899,N_2074);
and U2316 (N_2316,N_1668,In_1054);
nor U2317 (N_2317,N_82,N_2056);
or U2318 (N_2318,N_1594,N_1966);
xnor U2319 (N_2319,N_1987,N_1385);
and U2320 (N_2320,N_2055,N_2021);
and U2321 (N_2321,In_2398,N_1862);
or U2322 (N_2322,N_1848,N_677);
and U2323 (N_2323,N_2026,N_562);
and U2324 (N_2324,N_801,N_1419);
nand U2325 (N_2325,N_1405,N_1998);
nor U2326 (N_2326,N_1968,In_1347);
nand U2327 (N_2327,N_652,N_1895);
nand U2328 (N_2328,N_515,N_1342);
or U2329 (N_2329,N_1974,N_88);
and U2330 (N_2330,N_1843,N_1932);
nor U2331 (N_2331,In_1682,N_1207);
and U2332 (N_2332,N_979,In_1261);
and U2333 (N_2333,N_1893,In_1397);
or U2334 (N_2334,In_429,In_2711);
or U2335 (N_2335,N_1634,N_1697);
or U2336 (N_2336,In_2254,N_291);
or U2337 (N_2337,N_1147,N_2040);
nor U2338 (N_2338,N_767,N_1739);
nor U2339 (N_2339,N_1853,N_1838);
xor U2340 (N_2340,N_2082,N_2038);
xnor U2341 (N_2341,N_1721,N_1948);
and U2342 (N_2342,N_1819,N_1928);
xor U2343 (N_2343,N_29,N_1278);
nor U2344 (N_2344,In_1790,N_1753);
or U2345 (N_2345,N_1696,In_140);
nor U2346 (N_2346,N_1121,N_1559);
and U2347 (N_2347,N_1325,N_2008);
nor U2348 (N_2348,N_620,N_657);
nor U2349 (N_2349,N_542,In_1129);
nor U2350 (N_2350,N_1958,N_1828);
and U2351 (N_2351,N_2034,N_1811);
nor U2352 (N_2352,In_1166,In_586);
xor U2353 (N_2353,N_1485,N_609);
xor U2354 (N_2354,In_249,N_2063);
nand U2355 (N_2355,N_1905,In_1317);
nor U2356 (N_2356,N_964,N_1904);
or U2357 (N_2357,N_1467,N_2061);
xnor U2358 (N_2358,N_1511,N_1306);
xnor U2359 (N_2359,N_153,N_1408);
or U2360 (N_2360,N_1193,In_326);
nor U2361 (N_2361,In_2392,In_780);
or U2362 (N_2362,N_1991,N_1281);
and U2363 (N_2363,N_1988,N_1343);
or U2364 (N_2364,N_214,N_2044);
xor U2365 (N_2365,N_1644,N_1813);
nor U2366 (N_2366,N_1962,N_539);
or U2367 (N_2367,In_11,N_1400);
nand U2368 (N_2368,N_1965,N_1971);
nand U2369 (N_2369,N_737,In_1101);
xor U2370 (N_2370,N_1908,In_737);
and U2371 (N_2371,In_1385,N_1563);
and U2372 (N_2372,In_2331,In_1146);
xnor U2373 (N_2373,N_1232,N_1610);
xnor U2374 (N_2374,N_1311,N_1885);
nand U2375 (N_2375,N_1947,In_275);
or U2376 (N_2376,In_903,N_1179);
or U2377 (N_2377,N_1352,N_1399);
xnor U2378 (N_2378,In_165,N_903);
or U2379 (N_2379,N_1990,N_2060);
nor U2380 (N_2380,In_1934,N_1749);
nor U2381 (N_2381,N_701,N_1926);
xnor U2382 (N_2382,N_1919,N_1953);
xor U2383 (N_2383,In_1926,N_886);
and U2384 (N_2384,N_1220,In_2128);
nor U2385 (N_2385,N_1548,N_1887);
nor U2386 (N_2386,N_2098,N_1290);
nor U2387 (N_2387,N_1938,N_1852);
or U2388 (N_2388,In_97,N_1667);
xor U2389 (N_2389,In_432,In_1505);
nor U2390 (N_2390,In_1667,N_1858);
nor U2391 (N_2391,In_101,N_2071);
nor U2392 (N_2392,N_499,In_688);
nor U2393 (N_2393,N_1783,N_543);
or U2394 (N_2394,N_1519,N_1507);
and U2395 (N_2395,N_1837,N_1654);
or U2396 (N_2396,N_2068,N_1437);
and U2397 (N_2397,In_1112,In_531);
xnor U2398 (N_2398,N_1719,N_2078);
or U2399 (N_2399,In_1216,N_1763);
or U2400 (N_2400,N_1927,N_2233);
and U2401 (N_2401,In_1675,N_2035);
nor U2402 (N_2402,N_1954,N_2288);
or U2403 (N_2403,N_1945,N_2354);
xor U2404 (N_2404,N_2114,N_2136);
nor U2405 (N_2405,N_2239,In_931);
and U2406 (N_2406,N_129,N_1237);
nand U2407 (N_2407,In_2366,N_1561);
nand U2408 (N_2408,In_1283,N_632);
nand U2409 (N_2409,N_156,N_2176);
and U2410 (N_2410,N_2188,N_2365);
nor U2411 (N_2411,N_1353,N_1806);
nand U2412 (N_2412,N_2310,N_2332);
or U2413 (N_2413,In_820,N_2159);
nor U2414 (N_2414,N_2240,N_2146);
nor U2415 (N_2415,N_1756,N_854);
xor U2416 (N_2416,N_1472,N_2161);
nand U2417 (N_2417,N_2165,N_2057);
nand U2418 (N_2418,In_1467,N_2234);
and U2419 (N_2419,N_1952,N_1982);
xnor U2420 (N_2420,N_2091,N_1750);
and U2421 (N_2421,N_2276,N_2163);
or U2422 (N_2422,In_2250,N_2383);
nand U2423 (N_2423,N_2363,In_1359);
xnor U2424 (N_2424,N_1822,N_1665);
and U2425 (N_2425,N_2388,N_2156);
nand U2426 (N_2426,N_1647,N_1034);
and U2427 (N_2427,N_2384,N_2315);
nand U2428 (N_2428,N_2218,N_1980);
xor U2429 (N_2429,N_2141,N_1984);
nor U2430 (N_2430,N_2201,In_606);
nand U2431 (N_2431,N_2120,N_1661);
nand U2432 (N_2432,N_2186,N_2135);
or U2433 (N_2433,N_1198,In_2003);
nand U2434 (N_2434,N_1478,In_37);
and U2435 (N_2435,N_2075,N_2164);
xor U2436 (N_2436,In_16,N_2337);
nand U2437 (N_2437,N_2269,N_2263);
xnor U2438 (N_2438,In_1196,N_2245);
and U2439 (N_2439,N_2265,N_2268);
nor U2440 (N_2440,N_1556,N_1663);
xnor U2441 (N_2441,N_1880,N_2349);
and U2442 (N_2442,N_2373,N_2364);
nand U2443 (N_2443,N_2301,N_1526);
or U2444 (N_2444,N_2181,In_1465);
or U2445 (N_2445,N_2118,In_2767);
xnor U2446 (N_2446,N_929,N_1520);
nor U2447 (N_2447,N_1503,N_2214);
xor U2448 (N_2448,N_1348,N_2376);
nor U2449 (N_2449,N_2148,N_2316);
and U2450 (N_2450,N_2295,In_1479);
or U2451 (N_2451,N_2361,N_2255);
and U2452 (N_2452,N_2359,N_1878);
or U2453 (N_2453,N_2122,N_2121);
or U2454 (N_2454,N_2370,N_2261);
and U2455 (N_2455,N_299,N_2331);
xnor U2456 (N_2456,N_1782,N_2282);
and U2457 (N_2457,N_2293,N_2138);
and U2458 (N_2458,N_1979,N_2129);
xnor U2459 (N_2459,N_2323,N_2119);
or U2460 (N_2460,N_2385,N_1944);
xor U2461 (N_2461,N_2113,N_2220);
xnor U2462 (N_2462,N_2101,N_1963);
nand U2463 (N_2463,In_2428,N_2329);
xor U2464 (N_2464,N_1936,N_2346);
nor U2465 (N_2465,In_2842,N_2298);
nand U2466 (N_2466,N_1570,N_2251);
nand U2467 (N_2467,N_2105,N_2274);
xnor U2468 (N_2468,In_2420,N_1046);
nand U2469 (N_2469,N_1808,N_1747);
xor U2470 (N_2470,N_2109,In_1263);
or U2471 (N_2471,N_1849,N_2250);
nand U2472 (N_2472,N_2302,N_52);
or U2473 (N_2473,N_1780,N_2149);
or U2474 (N_2474,N_1784,In_2917);
or U2475 (N_2475,N_1473,N_840);
or U2476 (N_2476,N_1839,In_1104);
or U2477 (N_2477,N_2017,N_2290);
xor U2478 (N_2478,In_2422,N_1688);
and U2479 (N_2479,N_2048,N_2184);
xnor U2480 (N_2480,N_1729,N_1486);
nand U2481 (N_2481,N_2052,N_1860);
nor U2482 (N_2482,N_1295,N_2154);
and U2483 (N_2483,N_2333,N_2371);
and U2484 (N_2484,N_54,In_1019);
nor U2485 (N_2485,N_1142,In_2815);
nand U2486 (N_2486,N_659,N_2352);
nand U2487 (N_2487,N_2398,N_2173);
and U2488 (N_2488,In_1712,N_2213);
nor U2489 (N_2489,N_1492,N_1961);
xor U2490 (N_2490,N_2039,N_2024);
and U2491 (N_2491,N_2142,N_1341);
nand U2492 (N_2492,N_2020,In_1109);
nor U2493 (N_2493,N_1330,N_2286);
or U2494 (N_2494,N_2351,N_2238);
and U2495 (N_2495,N_1524,N_1942);
xnor U2496 (N_2496,N_2179,In_2110);
nor U2497 (N_2497,N_2046,N_2382);
or U2498 (N_2498,N_1742,N_2387);
nand U2499 (N_2499,N_1970,N_2336);
or U2500 (N_2500,N_1957,N_729);
nand U2501 (N_2501,N_2104,N_1513);
xnor U2502 (N_2502,N_1674,N_695);
and U2503 (N_2503,N_910,N_2093);
or U2504 (N_2504,N_902,N_2131);
nand U2505 (N_2505,N_2247,N_1890);
nor U2506 (N_2506,N_2172,N_2244);
nand U2507 (N_2507,N_2262,N_2128);
nor U2508 (N_2508,N_2228,N_2076);
xnor U2509 (N_2509,In_1612,N_2378);
or U2510 (N_2510,N_2079,N_2236);
nor U2511 (N_2511,N_2253,N_1710);
or U2512 (N_2512,N_2264,N_2356);
nor U2513 (N_2513,N_2227,N_2219);
or U2514 (N_2514,N_2080,N_2116);
nor U2515 (N_2515,N_2209,N_2100);
nor U2516 (N_2516,N_2372,N_1137);
and U2517 (N_2517,N_2241,N_2198);
nor U2518 (N_2518,N_2144,N_1931);
or U2519 (N_2519,N_2283,N_2249);
and U2520 (N_2520,N_2182,N_1698);
nor U2521 (N_2521,N_2350,N_2399);
xnor U2522 (N_2522,N_2013,N_2360);
xor U2523 (N_2523,N_244,N_2111);
xor U2524 (N_2524,N_2243,N_2127);
and U2525 (N_2525,N_2192,N_2103);
nand U2526 (N_2526,N_2152,N_1798);
nor U2527 (N_2527,N_2225,N_1866);
or U2528 (N_2528,N_2235,N_1992);
and U2529 (N_2529,N_2217,N_1451);
and U2530 (N_2530,N_2190,N_1380);
xor U2531 (N_2531,N_2258,N_2393);
nand U2532 (N_2532,N_2277,N_1705);
or U2533 (N_2533,In_1793,N_2291);
nor U2534 (N_2534,In_2448,N_2089);
nor U2535 (N_2535,N_2299,N_2115);
or U2536 (N_2536,N_548,N_1180);
or U2537 (N_2537,N_2348,N_2366);
nand U2538 (N_2538,N_2205,N_2125);
and U2539 (N_2539,N_1677,N_2311);
nor U2540 (N_2540,N_2260,N_2143);
or U2541 (N_2541,N_1596,N_2394);
or U2542 (N_2542,N_2390,N_2312);
or U2543 (N_2543,N_2195,N_2223);
nor U2544 (N_2544,N_2194,N_1933);
xor U2545 (N_2545,N_1901,N_2343);
xnor U2546 (N_2546,N_2232,N_1595);
and U2547 (N_2547,N_2203,N_2275);
xnor U2548 (N_2548,N_1917,In_270);
xor U2549 (N_2549,N_2177,N_2324);
xnor U2550 (N_2550,In_2963,N_2380);
nand U2551 (N_2551,N_2221,N_1907);
nor U2552 (N_2552,N_1884,N_1285);
or U2553 (N_2553,N_2147,N_1906);
xnor U2554 (N_2554,N_1827,N_1516);
or U2555 (N_2555,N_2229,N_2197);
or U2556 (N_2556,N_1621,N_1058);
or U2557 (N_2557,N_2222,N_2369);
and U2558 (N_2558,In_1890,N_1530);
or U2559 (N_2559,N_2306,N_2254);
nand U2560 (N_2560,In_1172,In_1472);
or U2561 (N_2561,N_2397,N_2355);
and U2562 (N_2562,N_2180,N_1449);
xnor U2563 (N_2563,N_85,N_2117);
and U2564 (N_2564,N_1969,N_565);
nor U2565 (N_2565,N_1943,N_1504);
or U2566 (N_2566,N_1916,N_2327);
nor U2567 (N_2567,N_2377,N_16);
nor U2568 (N_2568,In_1824,N_2320);
or U2569 (N_2569,N_2313,N_2279);
or U2570 (N_2570,N_2110,N_550);
and U2571 (N_2571,N_2167,N_379);
and U2572 (N_2572,N_2292,In_873);
xnor U2573 (N_2573,N_2157,N_2335);
and U2574 (N_2574,In_1090,N_2153);
and U2575 (N_2575,N_1683,N_1332);
nand U2576 (N_2576,N_2208,N_2340);
and U2577 (N_2577,N_2169,N_2183);
or U2578 (N_2578,N_2166,N_2112);
nand U2579 (N_2579,N_1031,In_2482);
and U2580 (N_2580,N_2170,N_993);
xnor U2581 (N_2581,N_2391,N_1641);
nor U2582 (N_2582,In_2513,N_2357);
xor U2583 (N_2583,N_2155,In_91);
nand U2584 (N_2584,N_1250,N_1861);
xor U2585 (N_2585,N_2133,N_2392);
and U2586 (N_2586,N_2191,In_186);
xor U2587 (N_2587,N_1108,N_1737);
nand U2588 (N_2588,N_1738,N_719);
and U2589 (N_2589,N_2326,N_2271);
nor U2590 (N_2590,N_2341,N_2362);
nor U2591 (N_2591,N_2139,N_2273);
or U2592 (N_2592,N_2389,N_2081);
xor U2593 (N_2593,N_2285,N_2102);
nor U2594 (N_2594,N_2037,N_2330);
xnor U2595 (N_2595,N_961,N_1541);
xnor U2596 (N_2596,N_1375,N_1078);
nand U2597 (N_2597,In_472,N_901);
xor U2598 (N_2598,N_2137,N_2266);
or U2599 (N_2599,N_2374,N_1799);
nor U2600 (N_2600,In_2795,In_397);
nor U2601 (N_2601,In_2207,In_2718);
xor U2602 (N_2602,N_2130,N_2325);
and U2603 (N_2603,N_2237,N_1975);
xor U2604 (N_2604,N_2178,In_1303);
nand U2605 (N_2605,N_1569,In_2289);
xor U2606 (N_2606,N_2319,N_2224);
or U2607 (N_2607,N_2029,N_2210);
nand U2608 (N_2608,N_2353,N_2296);
nand U2609 (N_2609,In_1056,N_1821);
xor U2610 (N_2610,In_1349,N_2160);
and U2611 (N_2611,N_2174,N_1706);
and U2612 (N_2612,N_2193,N_2257);
nor U2613 (N_2613,N_2338,N_1373);
xnor U2614 (N_2614,N_2309,N_2070);
and U2615 (N_2615,N_1823,N_2185);
and U2616 (N_2616,N_1536,N_2256);
nand U2617 (N_2617,N_2140,N_2322);
nand U2618 (N_2618,N_1759,N_1910);
nand U2619 (N_2619,N_2145,N_2287);
nand U2620 (N_2620,N_1007,N_2328);
or U2621 (N_2621,N_1921,N_2083);
xnor U2622 (N_2622,N_2036,In_125);
nor U2623 (N_2623,N_764,N_2005);
and U2624 (N_2624,N_1028,N_1327);
or U2625 (N_2625,N_1632,N_1829);
and U2626 (N_2626,N_1653,N_2395);
nand U2627 (N_2627,N_990,N_2207);
xor U2628 (N_2628,N_2007,N_1171);
nand U2629 (N_2629,N_1319,N_2151);
nand U2630 (N_2630,N_1591,N_2300);
nor U2631 (N_2631,N_330,N_2305);
nor U2632 (N_2632,N_1447,N_623);
nand U2633 (N_2633,N_1914,N_653);
xor U2634 (N_2634,N_2307,N_2196);
nor U2635 (N_2635,N_2278,N_2200);
or U2636 (N_2636,N_1886,N_2062);
and U2637 (N_2637,N_2206,N_2199);
xor U2638 (N_2638,N_2248,N_2368);
xor U2639 (N_2639,N_2270,N_2267);
or U2640 (N_2640,N_2342,N_1297);
nor U2641 (N_2641,N_1535,In_1011);
nand U2642 (N_2642,N_2231,N_2280);
nand U2643 (N_2643,N_1959,N_1733);
and U2644 (N_2644,N_1363,N_1645);
and U2645 (N_2645,In_1450,N_2281);
or U2646 (N_2646,N_1338,N_2272);
nor U2647 (N_2647,N_1834,N_2124);
xor U2648 (N_2648,N_2230,N_2168);
nand U2649 (N_2649,N_1855,In_38);
and U2650 (N_2650,N_1125,N_2107);
xor U2651 (N_2651,N_2303,N_2202);
xnor U2652 (N_2652,N_2150,N_2246);
nand U2653 (N_2653,In_252,N_1709);
nand U2654 (N_2654,N_2344,N_1925);
or U2655 (N_2655,N_1745,N_2171);
or U2656 (N_2656,N_1857,N_2162);
nor U2657 (N_2657,N_1930,N_421);
and U2658 (N_2658,N_1835,N_1502);
and U2659 (N_2659,N_466,N_2108);
xor U2660 (N_2660,In_1709,N_1735);
and U2661 (N_2661,N_2381,N_1178);
or U2662 (N_2662,N_1639,N_2321);
nor U2663 (N_2663,N_2347,N_2314);
or U2664 (N_2664,N_1637,N_2187);
or U2665 (N_2665,N_2317,N_2386);
or U2666 (N_2666,N_1912,N_2226);
and U2667 (N_2667,N_1339,In_362);
nand U2668 (N_2668,N_2242,N_2304);
xor U2669 (N_2669,In_234,N_2204);
nor U2670 (N_2670,N_2297,N_2134);
or U2671 (N_2671,N_80,N_2106);
and U2672 (N_2672,N_2158,In_457);
nor U2673 (N_2673,N_1863,N_1328);
or U2674 (N_2674,N_2308,In_2589);
xnor U2675 (N_2675,N_2211,N_1650);
or U2676 (N_2676,In_837,In_689);
xnor U2677 (N_2677,N_2215,N_1101);
nand U2678 (N_2678,N_2175,N_2123);
nand U2679 (N_2679,N_712,N_2289);
xnor U2680 (N_2680,N_1960,N_1761);
and U2681 (N_2681,N_2345,N_2126);
and U2682 (N_2682,N_1392,In_588);
nor U2683 (N_2683,N_2396,N_2216);
or U2684 (N_2684,N_2189,N_2023);
and U2685 (N_2685,N_1816,In_2288);
nand U2686 (N_2686,N_1872,N_2375);
xnor U2687 (N_2687,In_617,In_304);
nor U2688 (N_2688,N_2358,N_1923);
nand U2689 (N_2689,N_1913,N_2318);
or U2690 (N_2690,N_2334,N_2094);
or U2691 (N_2691,N_1801,N_1762);
xor U2692 (N_2692,N_2339,N_2212);
xor U2693 (N_2693,N_2252,N_2379);
or U2694 (N_2694,N_1612,N_2132);
and U2695 (N_2695,N_2042,N_1820);
nor U2696 (N_2696,N_2284,In_2987);
xor U2697 (N_2697,N_2294,N_2367);
xor U2698 (N_2698,N_2009,N_2259);
nand U2699 (N_2699,In_2208,In_692);
nand U2700 (N_2700,N_2402,N_2416);
nor U2701 (N_2701,N_2610,N_2462);
nor U2702 (N_2702,N_2656,N_2546);
nand U2703 (N_2703,N_2404,N_2513);
and U2704 (N_2704,N_2699,N_2526);
and U2705 (N_2705,N_2599,N_2470);
or U2706 (N_2706,N_2529,N_2620);
nor U2707 (N_2707,N_2647,N_2433);
nor U2708 (N_2708,N_2411,N_2458);
nor U2709 (N_2709,N_2447,N_2648);
nor U2710 (N_2710,N_2577,N_2615);
nand U2711 (N_2711,N_2540,N_2500);
nor U2712 (N_2712,N_2669,N_2479);
nor U2713 (N_2713,N_2641,N_2562);
and U2714 (N_2714,N_2486,N_2437);
xnor U2715 (N_2715,N_2473,N_2440);
nor U2716 (N_2716,N_2649,N_2681);
nand U2717 (N_2717,N_2607,N_2482);
or U2718 (N_2718,N_2525,N_2695);
nand U2719 (N_2719,N_2467,N_2468);
nand U2720 (N_2720,N_2679,N_2569);
nor U2721 (N_2721,N_2408,N_2658);
xor U2722 (N_2722,N_2521,N_2603);
nor U2723 (N_2723,N_2630,N_2680);
xor U2724 (N_2724,N_2629,N_2661);
xor U2725 (N_2725,N_2545,N_2466);
nor U2726 (N_2726,N_2444,N_2427);
and U2727 (N_2727,N_2561,N_2475);
nand U2728 (N_2728,N_2530,N_2512);
nand U2729 (N_2729,N_2657,N_2697);
nand U2730 (N_2730,N_2520,N_2481);
and U2731 (N_2731,N_2614,N_2509);
and U2732 (N_2732,N_2622,N_2464);
nand U2733 (N_2733,N_2413,N_2651);
nor U2734 (N_2734,N_2590,N_2635);
nand U2735 (N_2735,N_2452,N_2556);
or U2736 (N_2736,N_2628,N_2508);
or U2737 (N_2737,N_2484,N_2650);
or U2738 (N_2738,N_2598,N_2636);
and U2739 (N_2739,N_2499,N_2535);
and U2740 (N_2740,N_2673,N_2548);
and U2741 (N_2741,N_2469,N_2686);
or U2742 (N_2742,N_2426,N_2496);
nor U2743 (N_2743,N_2584,N_2559);
and U2744 (N_2744,N_2445,N_2631);
or U2745 (N_2745,N_2688,N_2563);
xor U2746 (N_2746,N_2660,N_2595);
nand U2747 (N_2747,N_2684,N_2687);
nand U2748 (N_2748,N_2642,N_2483);
nor U2749 (N_2749,N_2528,N_2517);
nor U2750 (N_2750,N_2410,N_2471);
xor U2751 (N_2751,N_2676,N_2572);
or U2752 (N_2752,N_2461,N_2438);
nor U2753 (N_2753,N_2672,N_2685);
nand U2754 (N_2754,N_2503,N_2538);
xnor U2755 (N_2755,N_2534,N_2533);
nand U2756 (N_2756,N_2576,N_2618);
xnor U2757 (N_2757,N_2409,N_2608);
nor U2758 (N_2758,N_2566,N_2507);
and U2759 (N_2759,N_2459,N_2574);
xor U2760 (N_2760,N_2463,N_2627);
or U2761 (N_2761,N_2449,N_2532);
nor U2762 (N_2762,N_2612,N_2417);
xor U2763 (N_2763,N_2544,N_2518);
nand U2764 (N_2764,N_2698,N_2455);
or U2765 (N_2765,N_2439,N_2543);
nor U2766 (N_2766,N_2653,N_2412);
nand U2767 (N_2767,N_2550,N_2575);
nor U2768 (N_2768,N_2609,N_2665);
and U2769 (N_2769,N_2527,N_2693);
or U2770 (N_2770,N_2583,N_2474);
xor U2771 (N_2771,N_2565,N_2425);
and U2772 (N_2772,N_2604,N_2493);
xor U2773 (N_2773,N_2505,N_2696);
xor U2774 (N_2774,N_2446,N_2616);
nand U2775 (N_2775,N_2586,N_2519);
and U2776 (N_2776,N_2560,N_2515);
xor U2777 (N_2777,N_2654,N_2621);
xnor U2778 (N_2778,N_2625,N_2571);
and U2779 (N_2779,N_2578,N_2597);
nor U2780 (N_2780,N_2516,N_2542);
nand U2781 (N_2781,N_2451,N_2549);
or U2782 (N_2782,N_2663,N_2429);
nor U2783 (N_2783,N_2624,N_2644);
or U2784 (N_2784,N_2420,N_2659);
nor U2785 (N_2785,N_2555,N_2585);
nand U2786 (N_2786,N_2454,N_2547);
nand U2787 (N_2787,N_2558,N_2593);
nor U2788 (N_2788,N_2421,N_2567);
and U2789 (N_2789,N_2424,N_2442);
nand U2790 (N_2790,N_2587,N_2457);
nor U2791 (N_2791,N_2692,N_2683);
nand U2792 (N_2792,N_2623,N_2606);
and U2793 (N_2793,N_2668,N_2406);
and U2794 (N_2794,N_2418,N_2589);
or U2795 (N_2795,N_2490,N_2489);
nand U2796 (N_2796,N_2662,N_2436);
or U2797 (N_2797,N_2579,N_2634);
nor U2798 (N_2798,N_2605,N_2403);
xnor U2799 (N_2799,N_2419,N_2594);
nand U2800 (N_2800,N_2472,N_2645);
nand U2801 (N_2801,N_2637,N_2480);
xnor U2802 (N_2802,N_2638,N_2477);
xor U2803 (N_2803,N_2422,N_2655);
nand U2804 (N_2804,N_2643,N_2450);
nand U2805 (N_2805,N_2488,N_2691);
or U2806 (N_2806,N_2553,N_2510);
xnor U2807 (N_2807,N_2431,N_2689);
or U2808 (N_2808,N_2580,N_2570);
and U2809 (N_2809,N_2582,N_2539);
or U2810 (N_2810,N_2491,N_2476);
or U2811 (N_2811,N_2423,N_2494);
nand U2812 (N_2812,N_2667,N_2541);
nand U2813 (N_2813,N_2531,N_2448);
xnor U2814 (N_2814,N_2405,N_2573);
or U2815 (N_2815,N_2497,N_2675);
xnor U2816 (N_2816,N_2504,N_2485);
or U2817 (N_2817,N_2511,N_2495);
nor U2818 (N_2818,N_2600,N_2588);
nand U2819 (N_2819,N_2492,N_2407);
or U2820 (N_2820,N_2524,N_2602);
nand U2821 (N_2821,N_2460,N_2428);
nand U2822 (N_2822,N_2677,N_2487);
and U2823 (N_2823,N_2498,N_2694);
nand U2824 (N_2824,N_2537,N_2557);
or U2825 (N_2825,N_2523,N_2554);
nor U2826 (N_2826,N_2581,N_2453);
nor U2827 (N_2827,N_2666,N_2400);
and U2828 (N_2828,N_2502,N_2639);
nand U2829 (N_2829,N_2674,N_2592);
nand U2830 (N_2830,N_2617,N_2611);
and U2831 (N_2831,N_2670,N_2664);
xnor U2832 (N_2832,N_2551,N_2646);
xor U2833 (N_2833,N_2632,N_2441);
xor U2834 (N_2834,N_2678,N_2430);
nor U2835 (N_2835,N_2613,N_2478);
and U2836 (N_2836,N_2601,N_2568);
or U2837 (N_2837,N_2506,N_2522);
or U2838 (N_2838,N_2652,N_2640);
nand U2839 (N_2839,N_2414,N_2633);
or U2840 (N_2840,N_2514,N_2619);
nand U2841 (N_2841,N_2465,N_2536);
nor U2842 (N_2842,N_2552,N_2456);
or U2843 (N_2843,N_2415,N_2671);
nand U2844 (N_2844,N_2682,N_2434);
or U2845 (N_2845,N_2596,N_2432);
xor U2846 (N_2846,N_2591,N_2501);
nor U2847 (N_2847,N_2443,N_2626);
nand U2848 (N_2848,N_2564,N_2690);
nand U2849 (N_2849,N_2435,N_2401);
or U2850 (N_2850,N_2565,N_2505);
nor U2851 (N_2851,N_2405,N_2559);
nor U2852 (N_2852,N_2552,N_2448);
and U2853 (N_2853,N_2500,N_2632);
and U2854 (N_2854,N_2626,N_2552);
xnor U2855 (N_2855,N_2643,N_2675);
nand U2856 (N_2856,N_2544,N_2548);
nor U2857 (N_2857,N_2695,N_2424);
or U2858 (N_2858,N_2664,N_2409);
nor U2859 (N_2859,N_2461,N_2626);
xnor U2860 (N_2860,N_2592,N_2465);
or U2861 (N_2861,N_2535,N_2599);
xnor U2862 (N_2862,N_2575,N_2437);
or U2863 (N_2863,N_2566,N_2683);
and U2864 (N_2864,N_2401,N_2476);
nand U2865 (N_2865,N_2666,N_2459);
xnor U2866 (N_2866,N_2634,N_2420);
nor U2867 (N_2867,N_2406,N_2631);
xor U2868 (N_2868,N_2458,N_2416);
or U2869 (N_2869,N_2615,N_2423);
nor U2870 (N_2870,N_2524,N_2650);
or U2871 (N_2871,N_2607,N_2630);
and U2872 (N_2872,N_2494,N_2536);
and U2873 (N_2873,N_2516,N_2683);
nand U2874 (N_2874,N_2527,N_2628);
and U2875 (N_2875,N_2415,N_2610);
nor U2876 (N_2876,N_2451,N_2479);
and U2877 (N_2877,N_2521,N_2674);
xnor U2878 (N_2878,N_2651,N_2650);
or U2879 (N_2879,N_2614,N_2667);
xor U2880 (N_2880,N_2541,N_2699);
nor U2881 (N_2881,N_2593,N_2420);
nor U2882 (N_2882,N_2648,N_2468);
xnor U2883 (N_2883,N_2541,N_2542);
xor U2884 (N_2884,N_2592,N_2478);
xnor U2885 (N_2885,N_2483,N_2631);
nor U2886 (N_2886,N_2402,N_2548);
nand U2887 (N_2887,N_2566,N_2620);
xnor U2888 (N_2888,N_2540,N_2453);
nor U2889 (N_2889,N_2481,N_2460);
and U2890 (N_2890,N_2429,N_2445);
or U2891 (N_2891,N_2489,N_2625);
xnor U2892 (N_2892,N_2617,N_2484);
nand U2893 (N_2893,N_2590,N_2425);
and U2894 (N_2894,N_2607,N_2605);
nand U2895 (N_2895,N_2534,N_2498);
and U2896 (N_2896,N_2429,N_2624);
or U2897 (N_2897,N_2635,N_2489);
xor U2898 (N_2898,N_2413,N_2541);
nor U2899 (N_2899,N_2540,N_2609);
nand U2900 (N_2900,N_2498,N_2616);
nor U2901 (N_2901,N_2582,N_2619);
nor U2902 (N_2902,N_2689,N_2684);
and U2903 (N_2903,N_2424,N_2562);
nor U2904 (N_2904,N_2615,N_2470);
nor U2905 (N_2905,N_2618,N_2449);
xor U2906 (N_2906,N_2555,N_2531);
nand U2907 (N_2907,N_2483,N_2461);
nor U2908 (N_2908,N_2692,N_2558);
or U2909 (N_2909,N_2404,N_2549);
xor U2910 (N_2910,N_2563,N_2419);
xor U2911 (N_2911,N_2643,N_2455);
and U2912 (N_2912,N_2508,N_2632);
xnor U2913 (N_2913,N_2470,N_2488);
nor U2914 (N_2914,N_2532,N_2621);
nor U2915 (N_2915,N_2419,N_2647);
nand U2916 (N_2916,N_2568,N_2624);
nor U2917 (N_2917,N_2600,N_2580);
or U2918 (N_2918,N_2407,N_2538);
and U2919 (N_2919,N_2546,N_2445);
and U2920 (N_2920,N_2519,N_2649);
nand U2921 (N_2921,N_2588,N_2581);
and U2922 (N_2922,N_2512,N_2422);
or U2923 (N_2923,N_2530,N_2532);
xor U2924 (N_2924,N_2532,N_2614);
nor U2925 (N_2925,N_2419,N_2645);
nor U2926 (N_2926,N_2510,N_2551);
nor U2927 (N_2927,N_2594,N_2549);
nand U2928 (N_2928,N_2516,N_2531);
or U2929 (N_2929,N_2560,N_2493);
or U2930 (N_2930,N_2642,N_2502);
nand U2931 (N_2931,N_2579,N_2556);
xor U2932 (N_2932,N_2434,N_2618);
xor U2933 (N_2933,N_2615,N_2655);
and U2934 (N_2934,N_2451,N_2561);
nand U2935 (N_2935,N_2476,N_2568);
and U2936 (N_2936,N_2503,N_2604);
nor U2937 (N_2937,N_2422,N_2522);
xor U2938 (N_2938,N_2603,N_2450);
xor U2939 (N_2939,N_2500,N_2669);
nand U2940 (N_2940,N_2464,N_2646);
nor U2941 (N_2941,N_2607,N_2489);
or U2942 (N_2942,N_2452,N_2431);
nand U2943 (N_2943,N_2664,N_2579);
xnor U2944 (N_2944,N_2661,N_2653);
nor U2945 (N_2945,N_2530,N_2680);
and U2946 (N_2946,N_2650,N_2515);
nand U2947 (N_2947,N_2655,N_2577);
nor U2948 (N_2948,N_2409,N_2651);
and U2949 (N_2949,N_2472,N_2427);
xor U2950 (N_2950,N_2442,N_2560);
xnor U2951 (N_2951,N_2691,N_2652);
and U2952 (N_2952,N_2412,N_2662);
and U2953 (N_2953,N_2515,N_2574);
xor U2954 (N_2954,N_2585,N_2611);
xnor U2955 (N_2955,N_2548,N_2497);
nand U2956 (N_2956,N_2535,N_2451);
and U2957 (N_2957,N_2427,N_2699);
and U2958 (N_2958,N_2428,N_2513);
nand U2959 (N_2959,N_2643,N_2565);
nor U2960 (N_2960,N_2585,N_2580);
nand U2961 (N_2961,N_2410,N_2652);
or U2962 (N_2962,N_2600,N_2613);
nor U2963 (N_2963,N_2588,N_2455);
xor U2964 (N_2964,N_2582,N_2418);
nor U2965 (N_2965,N_2501,N_2695);
nor U2966 (N_2966,N_2574,N_2640);
and U2967 (N_2967,N_2456,N_2545);
xor U2968 (N_2968,N_2578,N_2689);
nand U2969 (N_2969,N_2677,N_2475);
or U2970 (N_2970,N_2502,N_2521);
xor U2971 (N_2971,N_2595,N_2470);
nor U2972 (N_2972,N_2438,N_2531);
nand U2973 (N_2973,N_2508,N_2676);
xnor U2974 (N_2974,N_2631,N_2646);
or U2975 (N_2975,N_2642,N_2449);
xor U2976 (N_2976,N_2524,N_2578);
nand U2977 (N_2977,N_2448,N_2618);
xnor U2978 (N_2978,N_2427,N_2428);
or U2979 (N_2979,N_2507,N_2668);
and U2980 (N_2980,N_2624,N_2527);
xor U2981 (N_2981,N_2471,N_2554);
xnor U2982 (N_2982,N_2407,N_2576);
nand U2983 (N_2983,N_2400,N_2527);
and U2984 (N_2984,N_2555,N_2642);
or U2985 (N_2985,N_2504,N_2558);
or U2986 (N_2986,N_2479,N_2617);
nor U2987 (N_2987,N_2620,N_2674);
and U2988 (N_2988,N_2464,N_2641);
and U2989 (N_2989,N_2675,N_2582);
nor U2990 (N_2990,N_2624,N_2581);
nor U2991 (N_2991,N_2594,N_2555);
xnor U2992 (N_2992,N_2530,N_2667);
and U2993 (N_2993,N_2528,N_2651);
nand U2994 (N_2994,N_2445,N_2515);
nand U2995 (N_2995,N_2696,N_2467);
xor U2996 (N_2996,N_2524,N_2451);
nor U2997 (N_2997,N_2567,N_2653);
or U2998 (N_2998,N_2656,N_2557);
nor U2999 (N_2999,N_2444,N_2682);
nand U3000 (N_3000,N_2986,N_2997);
xnor U3001 (N_3001,N_2809,N_2745);
nand U3002 (N_3002,N_2941,N_2749);
nor U3003 (N_3003,N_2895,N_2803);
xor U3004 (N_3004,N_2978,N_2816);
and U3005 (N_3005,N_2922,N_2714);
xor U3006 (N_3006,N_2929,N_2826);
nor U3007 (N_3007,N_2884,N_2717);
xnor U3008 (N_3008,N_2709,N_2973);
xor U3009 (N_3009,N_2873,N_2733);
nor U3010 (N_3010,N_2737,N_2950);
nor U3011 (N_3011,N_2930,N_2847);
nor U3012 (N_3012,N_2976,N_2833);
nand U3013 (N_3013,N_2940,N_2876);
nor U3014 (N_3014,N_2837,N_2964);
and U3015 (N_3015,N_2993,N_2947);
and U3016 (N_3016,N_2741,N_2901);
and U3017 (N_3017,N_2788,N_2701);
nor U3018 (N_3018,N_2914,N_2946);
nand U3019 (N_3019,N_2753,N_2731);
or U3020 (N_3020,N_2888,N_2920);
and U3021 (N_3021,N_2766,N_2834);
and U3022 (N_3022,N_2751,N_2711);
and U3023 (N_3023,N_2878,N_2892);
xnor U3024 (N_3024,N_2750,N_2921);
and U3025 (N_3025,N_2814,N_2805);
or U3026 (N_3026,N_2704,N_2974);
nand U3027 (N_3027,N_2867,N_2724);
xor U3028 (N_3028,N_2813,N_2938);
nand U3029 (N_3029,N_2860,N_2885);
xor U3030 (N_3030,N_2861,N_2829);
nor U3031 (N_3031,N_2739,N_2736);
xor U3032 (N_3032,N_2807,N_2850);
nor U3033 (N_3033,N_2913,N_2996);
nor U3034 (N_3034,N_2721,N_2952);
and U3035 (N_3035,N_2783,N_2735);
nand U3036 (N_3036,N_2887,N_2911);
nand U3037 (N_3037,N_2866,N_2747);
or U3038 (N_3038,N_2726,N_2728);
and U3039 (N_3039,N_2894,N_2916);
nor U3040 (N_3040,N_2848,N_2907);
nand U3041 (N_3041,N_2754,N_2810);
xnor U3042 (N_3042,N_2982,N_2835);
nand U3043 (N_3043,N_2919,N_2971);
nor U3044 (N_3044,N_2994,N_2980);
nor U3045 (N_3045,N_2933,N_2825);
xnor U3046 (N_3046,N_2725,N_2801);
and U3047 (N_3047,N_2937,N_2862);
and U3048 (N_3048,N_2778,N_2927);
xor U3049 (N_3049,N_2798,N_2926);
nand U3050 (N_3050,N_2961,N_2792);
nor U3051 (N_3051,N_2968,N_2932);
or U3052 (N_3052,N_2991,N_2757);
nand U3053 (N_3053,N_2943,N_2705);
and U3054 (N_3054,N_2794,N_2820);
and U3055 (N_3055,N_2975,N_2761);
or U3056 (N_3056,N_2874,N_2967);
and U3057 (N_3057,N_2984,N_2910);
or U3058 (N_3058,N_2791,N_2954);
nor U3059 (N_3059,N_2990,N_2746);
and U3060 (N_3060,N_2918,N_2828);
nor U3061 (N_3061,N_2729,N_2905);
and U3062 (N_3062,N_2955,N_2844);
nand U3063 (N_3063,N_2995,N_2708);
or U3064 (N_3064,N_2858,N_2845);
nor U3065 (N_3065,N_2893,N_2908);
or U3066 (N_3066,N_2896,N_2945);
and U3067 (N_3067,N_2942,N_2793);
nand U3068 (N_3068,N_2832,N_2843);
xor U3069 (N_3069,N_2883,N_2764);
nand U3070 (N_3070,N_2868,N_2912);
xor U3071 (N_3071,N_2979,N_2966);
xnor U3072 (N_3072,N_2956,N_2902);
or U3073 (N_3073,N_2931,N_2999);
or U3074 (N_3074,N_2738,N_2727);
nand U3075 (N_3075,N_2981,N_2762);
xor U3076 (N_3076,N_2758,N_2957);
nand U3077 (N_3077,N_2806,N_2787);
and U3078 (N_3078,N_2872,N_2768);
nand U3079 (N_3079,N_2742,N_2821);
nor U3080 (N_3080,N_2871,N_2998);
nor U3081 (N_3081,N_2811,N_2881);
nor U3082 (N_3082,N_2812,N_2859);
nor U3083 (N_3083,N_2772,N_2935);
xnor U3084 (N_3084,N_2877,N_2953);
or U3085 (N_3085,N_2818,N_2795);
and U3086 (N_3086,N_2780,N_2886);
xor U3087 (N_3087,N_2936,N_2989);
or U3088 (N_3088,N_2863,N_2889);
xnor U3089 (N_3089,N_2836,N_2944);
and U3090 (N_3090,N_2804,N_2734);
or U3091 (N_3091,N_2934,N_2775);
nor U3092 (N_3092,N_2962,N_2924);
xnor U3093 (N_3093,N_2959,N_2915);
or U3094 (N_3094,N_2857,N_2760);
or U3095 (N_3095,N_2906,N_2700);
nor U3096 (N_3096,N_2853,N_2917);
or U3097 (N_3097,N_2819,N_2838);
nand U3098 (N_3098,N_2909,N_2713);
or U3099 (N_3099,N_2904,N_2782);
or U3100 (N_3100,N_2827,N_2707);
or U3101 (N_3101,N_2800,N_2903);
nor U3102 (N_3102,N_2824,N_2846);
or U3103 (N_3103,N_2732,N_2744);
nor U3104 (N_3104,N_2965,N_2719);
nor U3105 (N_3105,N_2992,N_2756);
or U3106 (N_3106,N_2988,N_2797);
and U3107 (N_3107,N_2770,N_2856);
and U3108 (N_3108,N_2808,N_2755);
nor U3109 (N_3109,N_2928,N_2703);
nor U3110 (N_3110,N_2712,N_2958);
or U3111 (N_3111,N_2785,N_2784);
xor U3112 (N_3112,N_2900,N_2830);
nor U3113 (N_3113,N_2875,N_2702);
nand U3114 (N_3114,N_2977,N_2939);
and U3115 (N_3115,N_2983,N_2779);
or U3116 (N_3116,N_2822,N_2969);
and U3117 (N_3117,N_2882,N_2718);
or U3118 (N_3118,N_2752,N_2865);
or U3119 (N_3119,N_2972,N_2716);
and U3120 (N_3120,N_2951,N_2852);
nor U3121 (N_3121,N_2715,N_2786);
nor U3122 (N_3122,N_2817,N_2765);
and U3123 (N_3123,N_2773,N_2781);
nand U3124 (N_3124,N_2767,N_2851);
nand U3125 (N_3125,N_2854,N_2710);
nand U3126 (N_3126,N_2855,N_2763);
and U3127 (N_3127,N_2899,N_2796);
and U3128 (N_3128,N_2880,N_2777);
or U3129 (N_3129,N_2864,N_2831);
and U3130 (N_3130,N_2730,N_2963);
nand U3131 (N_3131,N_2740,N_2890);
nand U3132 (N_3132,N_2960,N_2970);
xor U3133 (N_3133,N_2769,N_2841);
xor U3134 (N_3134,N_2985,N_2925);
nor U3135 (N_3135,N_2923,N_2840);
nand U3136 (N_3136,N_2723,N_2774);
and U3137 (N_3137,N_2789,N_2790);
and U3138 (N_3138,N_2799,N_2815);
and U3139 (N_3139,N_2948,N_2879);
nand U3140 (N_3140,N_2748,N_2759);
or U3141 (N_3141,N_2849,N_2823);
or U3142 (N_3142,N_2870,N_2720);
nand U3143 (N_3143,N_2743,N_2897);
xnor U3144 (N_3144,N_2949,N_2771);
xnor U3145 (N_3145,N_2869,N_2842);
nor U3146 (N_3146,N_2898,N_2891);
or U3147 (N_3147,N_2722,N_2987);
and U3148 (N_3148,N_2839,N_2706);
or U3149 (N_3149,N_2776,N_2802);
nor U3150 (N_3150,N_2874,N_2896);
nor U3151 (N_3151,N_2989,N_2789);
or U3152 (N_3152,N_2833,N_2766);
nand U3153 (N_3153,N_2735,N_2766);
nor U3154 (N_3154,N_2862,N_2748);
or U3155 (N_3155,N_2916,N_2783);
or U3156 (N_3156,N_2903,N_2746);
and U3157 (N_3157,N_2998,N_2939);
xnor U3158 (N_3158,N_2820,N_2972);
nand U3159 (N_3159,N_2855,N_2912);
nor U3160 (N_3160,N_2932,N_2739);
nor U3161 (N_3161,N_2766,N_2975);
nand U3162 (N_3162,N_2937,N_2796);
nor U3163 (N_3163,N_2706,N_2937);
nand U3164 (N_3164,N_2985,N_2710);
nor U3165 (N_3165,N_2724,N_2896);
and U3166 (N_3166,N_2899,N_2731);
nand U3167 (N_3167,N_2853,N_2739);
nor U3168 (N_3168,N_2878,N_2893);
and U3169 (N_3169,N_2836,N_2805);
nor U3170 (N_3170,N_2949,N_2883);
and U3171 (N_3171,N_2974,N_2789);
or U3172 (N_3172,N_2723,N_2769);
and U3173 (N_3173,N_2905,N_2828);
xnor U3174 (N_3174,N_2767,N_2849);
nor U3175 (N_3175,N_2730,N_2907);
and U3176 (N_3176,N_2770,N_2837);
or U3177 (N_3177,N_2925,N_2926);
xor U3178 (N_3178,N_2900,N_2793);
xnor U3179 (N_3179,N_2724,N_2768);
nand U3180 (N_3180,N_2973,N_2896);
nor U3181 (N_3181,N_2867,N_2953);
nand U3182 (N_3182,N_2845,N_2976);
and U3183 (N_3183,N_2850,N_2761);
nand U3184 (N_3184,N_2863,N_2898);
nand U3185 (N_3185,N_2899,N_2950);
nand U3186 (N_3186,N_2807,N_2952);
nand U3187 (N_3187,N_2882,N_2856);
or U3188 (N_3188,N_2766,N_2888);
xnor U3189 (N_3189,N_2905,N_2983);
and U3190 (N_3190,N_2990,N_2887);
nor U3191 (N_3191,N_2770,N_2815);
xor U3192 (N_3192,N_2707,N_2746);
nor U3193 (N_3193,N_2746,N_2957);
or U3194 (N_3194,N_2986,N_2896);
nor U3195 (N_3195,N_2813,N_2994);
xor U3196 (N_3196,N_2834,N_2748);
or U3197 (N_3197,N_2959,N_2969);
or U3198 (N_3198,N_2928,N_2895);
nor U3199 (N_3199,N_2730,N_2742);
xnor U3200 (N_3200,N_2980,N_2768);
and U3201 (N_3201,N_2792,N_2763);
xor U3202 (N_3202,N_2788,N_2923);
nand U3203 (N_3203,N_2735,N_2846);
or U3204 (N_3204,N_2813,N_2708);
nor U3205 (N_3205,N_2752,N_2819);
and U3206 (N_3206,N_2775,N_2982);
nand U3207 (N_3207,N_2885,N_2927);
or U3208 (N_3208,N_2877,N_2755);
nand U3209 (N_3209,N_2719,N_2912);
xor U3210 (N_3210,N_2846,N_2832);
or U3211 (N_3211,N_2985,N_2984);
or U3212 (N_3212,N_2718,N_2901);
and U3213 (N_3213,N_2711,N_2748);
nor U3214 (N_3214,N_2706,N_2741);
xor U3215 (N_3215,N_2788,N_2723);
nand U3216 (N_3216,N_2765,N_2814);
xnor U3217 (N_3217,N_2785,N_2888);
nor U3218 (N_3218,N_2908,N_2729);
xnor U3219 (N_3219,N_2972,N_2885);
nor U3220 (N_3220,N_2914,N_2981);
and U3221 (N_3221,N_2838,N_2902);
and U3222 (N_3222,N_2817,N_2755);
and U3223 (N_3223,N_2818,N_2733);
and U3224 (N_3224,N_2956,N_2986);
and U3225 (N_3225,N_2895,N_2850);
or U3226 (N_3226,N_2818,N_2808);
nand U3227 (N_3227,N_2725,N_2719);
xnor U3228 (N_3228,N_2934,N_2935);
nor U3229 (N_3229,N_2945,N_2844);
nand U3230 (N_3230,N_2838,N_2709);
nand U3231 (N_3231,N_2745,N_2724);
nor U3232 (N_3232,N_2853,N_2795);
nand U3233 (N_3233,N_2967,N_2737);
or U3234 (N_3234,N_2720,N_2996);
nor U3235 (N_3235,N_2944,N_2733);
nand U3236 (N_3236,N_2820,N_2808);
or U3237 (N_3237,N_2818,N_2888);
or U3238 (N_3238,N_2999,N_2799);
or U3239 (N_3239,N_2979,N_2793);
and U3240 (N_3240,N_2976,N_2703);
or U3241 (N_3241,N_2884,N_2804);
nor U3242 (N_3242,N_2722,N_2768);
nand U3243 (N_3243,N_2765,N_2977);
and U3244 (N_3244,N_2836,N_2708);
nand U3245 (N_3245,N_2884,N_2993);
and U3246 (N_3246,N_2811,N_2720);
and U3247 (N_3247,N_2909,N_2750);
nor U3248 (N_3248,N_2731,N_2901);
and U3249 (N_3249,N_2982,N_2985);
nor U3250 (N_3250,N_2907,N_2773);
and U3251 (N_3251,N_2709,N_2948);
xor U3252 (N_3252,N_2750,N_2726);
xnor U3253 (N_3253,N_2731,N_2963);
nand U3254 (N_3254,N_2768,N_2932);
xor U3255 (N_3255,N_2704,N_2894);
or U3256 (N_3256,N_2802,N_2865);
nand U3257 (N_3257,N_2716,N_2747);
xor U3258 (N_3258,N_2874,N_2773);
nor U3259 (N_3259,N_2768,N_2785);
and U3260 (N_3260,N_2765,N_2797);
nand U3261 (N_3261,N_2715,N_2858);
and U3262 (N_3262,N_2954,N_2914);
or U3263 (N_3263,N_2971,N_2710);
or U3264 (N_3264,N_2808,N_2863);
nand U3265 (N_3265,N_2846,N_2742);
and U3266 (N_3266,N_2805,N_2968);
or U3267 (N_3267,N_2834,N_2746);
nor U3268 (N_3268,N_2984,N_2874);
xor U3269 (N_3269,N_2939,N_2875);
nor U3270 (N_3270,N_2861,N_2745);
nor U3271 (N_3271,N_2844,N_2757);
xor U3272 (N_3272,N_2970,N_2832);
nand U3273 (N_3273,N_2789,N_2959);
or U3274 (N_3274,N_2925,N_2817);
xor U3275 (N_3275,N_2937,N_2991);
and U3276 (N_3276,N_2869,N_2935);
or U3277 (N_3277,N_2813,N_2982);
or U3278 (N_3278,N_2949,N_2956);
xor U3279 (N_3279,N_2846,N_2758);
nand U3280 (N_3280,N_2785,N_2710);
and U3281 (N_3281,N_2808,N_2790);
and U3282 (N_3282,N_2876,N_2916);
nor U3283 (N_3283,N_2796,N_2983);
nor U3284 (N_3284,N_2857,N_2873);
or U3285 (N_3285,N_2883,N_2973);
nor U3286 (N_3286,N_2741,N_2784);
and U3287 (N_3287,N_2786,N_2992);
nand U3288 (N_3288,N_2709,N_2837);
or U3289 (N_3289,N_2877,N_2775);
or U3290 (N_3290,N_2747,N_2711);
nand U3291 (N_3291,N_2753,N_2996);
nor U3292 (N_3292,N_2835,N_2705);
and U3293 (N_3293,N_2889,N_2834);
xor U3294 (N_3294,N_2849,N_2740);
and U3295 (N_3295,N_2874,N_2720);
and U3296 (N_3296,N_2904,N_2743);
nand U3297 (N_3297,N_2824,N_2819);
nor U3298 (N_3298,N_2780,N_2904);
nor U3299 (N_3299,N_2879,N_2838);
nand U3300 (N_3300,N_3263,N_3206);
xor U3301 (N_3301,N_3167,N_3141);
and U3302 (N_3302,N_3181,N_3293);
nor U3303 (N_3303,N_3104,N_3267);
nand U3304 (N_3304,N_3113,N_3053);
or U3305 (N_3305,N_3004,N_3028);
or U3306 (N_3306,N_3086,N_3117);
and U3307 (N_3307,N_3207,N_3173);
or U3308 (N_3308,N_3059,N_3144);
nand U3309 (N_3309,N_3220,N_3123);
xnor U3310 (N_3310,N_3175,N_3080);
nand U3311 (N_3311,N_3229,N_3067);
nand U3312 (N_3312,N_3023,N_3275);
or U3313 (N_3313,N_3024,N_3231);
nand U3314 (N_3314,N_3218,N_3076);
nor U3315 (N_3315,N_3255,N_3165);
xor U3316 (N_3316,N_3073,N_3202);
nor U3317 (N_3317,N_3066,N_3283);
nor U3318 (N_3318,N_3217,N_3014);
nor U3319 (N_3319,N_3243,N_3057);
nand U3320 (N_3320,N_3156,N_3044);
and U3321 (N_3321,N_3169,N_3171);
or U3322 (N_3322,N_3237,N_3034);
nand U3323 (N_3323,N_3108,N_3159);
nand U3324 (N_3324,N_3046,N_3025);
and U3325 (N_3325,N_3155,N_3258);
nor U3326 (N_3326,N_3128,N_3008);
nor U3327 (N_3327,N_3278,N_3092);
xor U3328 (N_3328,N_3042,N_3016);
nand U3329 (N_3329,N_3257,N_3051);
or U3330 (N_3330,N_3048,N_3249);
and U3331 (N_3331,N_3285,N_3027);
nand U3332 (N_3332,N_3158,N_3195);
or U3333 (N_3333,N_3287,N_3070);
nor U3334 (N_3334,N_3199,N_3238);
and U3335 (N_3335,N_3244,N_3031);
or U3336 (N_3336,N_3127,N_3193);
nor U3337 (N_3337,N_3242,N_3094);
and U3338 (N_3338,N_3083,N_3132);
xor U3339 (N_3339,N_3182,N_3029);
nor U3340 (N_3340,N_3254,N_3111);
nand U3341 (N_3341,N_3105,N_3277);
and U3342 (N_3342,N_3147,N_3078);
or U3343 (N_3343,N_3134,N_3178);
and U3344 (N_3344,N_3118,N_3272);
nor U3345 (N_3345,N_3280,N_3087);
xnor U3346 (N_3346,N_3019,N_3266);
xnor U3347 (N_3347,N_3114,N_3268);
xnor U3348 (N_3348,N_3174,N_3055);
or U3349 (N_3349,N_3216,N_3071);
xor U3350 (N_3350,N_3191,N_3219);
and U3351 (N_3351,N_3299,N_3115);
nand U3352 (N_3352,N_3192,N_3126);
nand U3353 (N_3353,N_3274,N_3183);
and U3354 (N_3354,N_3098,N_3050);
xor U3355 (N_3355,N_3200,N_3194);
and U3356 (N_3356,N_3101,N_3236);
nand U3357 (N_3357,N_3136,N_3125);
and U3358 (N_3358,N_3010,N_3106);
nand U3359 (N_3359,N_3011,N_3168);
or U3360 (N_3360,N_3210,N_3061);
nor U3361 (N_3361,N_3189,N_3045);
nor U3362 (N_3362,N_3110,N_3228);
nor U3363 (N_3363,N_3058,N_3079);
and U3364 (N_3364,N_3140,N_3063);
nand U3365 (N_3365,N_3120,N_3259);
nand U3366 (N_3366,N_3157,N_3065);
nor U3367 (N_3367,N_3163,N_3099);
and U3368 (N_3368,N_3121,N_3291);
or U3369 (N_3369,N_3021,N_3253);
or U3370 (N_3370,N_3064,N_3166);
and U3371 (N_3371,N_3172,N_3222);
nand U3372 (N_3372,N_3088,N_3139);
and U3373 (N_3373,N_3015,N_3124);
and U3374 (N_3374,N_3143,N_3007);
nor U3375 (N_3375,N_3142,N_3116);
and U3376 (N_3376,N_3233,N_3035);
xnor U3377 (N_3377,N_3271,N_3074);
and U3378 (N_3378,N_3187,N_3091);
and U3379 (N_3379,N_3264,N_3054);
xor U3380 (N_3380,N_3049,N_3234);
nor U3381 (N_3381,N_3138,N_3164);
nand U3382 (N_3382,N_3020,N_3224);
or U3383 (N_3383,N_3297,N_3112);
xnor U3384 (N_3384,N_3043,N_3246);
nor U3385 (N_3385,N_3282,N_3060);
nor U3386 (N_3386,N_3241,N_3056);
or U3387 (N_3387,N_3081,N_3265);
nand U3388 (N_3388,N_3018,N_3072);
or U3389 (N_3389,N_3270,N_3288);
nand U3390 (N_3390,N_3284,N_3204);
or U3391 (N_3391,N_3279,N_3290);
xor U3392 (N_3392,N_3030,N_3221);
xor U3393 (N_3393,N_3149,N_3240);
xnor U3394 (N_3394,N_3036,N_3069);
or U3395 (N_3395,N_3040,N_3000);
nand U3396 (N_3396,N_3033,N_3214);
nor U3397 (N_3397,N_3145,N_3198);
or U3398 (N_3398,N_3184,N_3269);
nor U3399 (N_3399,N_3102,N_3235);
or U3400 (N_3400,N_3245,N_3292);
nor U3401 (N_3401,N_3012,N_3131);
nor U3402 (N_3402,N_3013,N_3135);
xor U3403 (N_3403,N_3185,N_3090);
nand U3404 (N_3404,N_3032,N_3026);
nand U3405 (N_3405,N_3154,N_3006);
or U3406 (N_3406,N_3262,N_3153);
xnor U3407 (N_3407,N_3068,N_3089);
or U3408 (N_3408,N_3225,N_3203);
nand U3409 (N_3409,N_3186,N_3211);
or U3410 (N_3410,N_3295,N_3205);
nor U3411 (N_3411,N_3130,N_3075);
xor U3412 (N_3412,N_3129,N_3232);
and U3413 (N_3413,N_3190,N_3085);
nor U3414 (N_3414,N_3002,N_3215);
and U3415 (N_3415,N_3096,N_3146);
nand U3416 (N_3416,N_3151,N_3084);
xor U3417 (N_3417,N_3095,N_3247);
nor U3418 (N_3418,N_3180,N_3097);
nor U3419 (N_3419,N_3152,N_3005);
nor U3420 (N_3420,N_3041,N_3286);
xnor U3421 (N_3421,N_3093,N_3294);
and U3422 (N_3422,N_3230,N_3226);
nand U3423 (N_3423,N_3122,N_3197);
xnor U3424 (N_3424,N_3261,N_3188);
nand U3425 (N_3425,N_3296,N_3298);
nand U3426 (N_3426,N_3150,N_3227);
nand U3427 (N_3427,N_3201,N_3209);
nand U3428 (N_3428,N_3208,N_3022);
or U3429 (N_3429,N_3289,N_3223);
or U3430 (N_3430,N_3179,N_3119);
xnor U3431 (N_3431,N_3103,N_3037);
or U3432 (N_3432,N_3212,N_3177);
nand U3433 (N_3433,N_3047,N_3148);
nor U3434 (N_3434,N_3137,N_3170);
nor U3435 (N_3435,N_3009,N_3251);
nand U3436 (N_3436,N_3213,N_3038);
nand U3437 (N_3437,N_3176,N_3107);
or U3438 (N_3438,N_3276,N_3109);
or U3439 (N_3439,N_3052,N_3281);
xor U3440 (N_3440,N_3133,N_3250);
or U3441 (N_3441,N_3248,N_3273);
nand U3442 (N_3442,N_3003,N_3260);
and U3443 (N_3443,N_3162,N_3001);
nand U3444 (N_3444,N_3252,N_3256);
and U3445 (N_3445,N_3196,N_3161);
nand U3446 (N_3446,N_3039,N_3062);
or U3447 (N_3447,N_3100,N_3017);
and U3448 (N_3448,N_3077,N_3239);
or U3449 (N_3449,N_3082,N_3160);
nor U3450 (N_3450,N_3134,N_3299);
nor U3451 (N_3451,N_3255,N_3091);
and U3452 (N_3452,N_3069,N_3284);
or U3453 (N_3453,N_3066,N_3209);
and U3454 (N_3454,N_3258,N_3049);
or U3455 (N_3455,N_3007,N_3049);
xor U3456 (N_3456,N_3042,N_3052);
and U3457 (N_3457,N_3024,N_3067);
nand U3458 (N_3458,N_3103,N_3226);
xor U3459 (N_3459,N_3033,N_3161);
xor U3460 (N_3460,N_3274,N_3122);
and U3461 (N_3461,N_3036,N_3285);
xor U3462 (N_3462,N_3014,N_3072);
xnor U3463 (N_3463,N_3169,N_3184);
or U3464 (N_3464,N_3039,N_3033);
or U3465 (N_3465,N_3102,N_3247);
and U3466 (N_3466,N_3068,N_3036);
and U3467 (N_3467,N_3099,N_3279);
xor U3468 (N_3468,N_3289,N_3158);
or U3469 (N_3469,N_3099,N_3206);
and U3470 (N_3470,N_3042,N_3144);
nor U3471 (N_3471,N_3201,N_3258);
nor U3472 (N_3472,N_3095,N_3293);
and U3473 (N_3473,N_3049,N_3179);
or U3474 (N_3474,N_3153,N_3022);
xnor U3475 (N_3475,N_3044,N_3130);
nor U3476 (N_3476,N_3175,N_3114);
and U3477 (N_3477,N_3267,N_3011);
or U3478 (N_3478,N_3267,N_3182);
nand U3479 (N_3479,N_3197,N_3258);
xor U3480 (N_3480,N_3197,N_3027);
xnor U3481 (N_3481,N_3174,N_3204);
xnor U3482 (N_3482,N_3261,N_3277);
nor U3483 (N_3483,N_3157,N_3012);
xor U3484 (N_3484,N_3271,N_3050);
nor U3485 (N_3485,N_3165,N_3278);
nand U3486 (N_3486,N_3108,N_3144);
nand U3487 (N_3487,N_3138,N_3141);
nor U3488 (N_3488,N_3003,N_3169);
and U3489 (N_3489,N_3205,N_3266);
xnor U3490 (N_3490,N_3126,N_3045);
or U3491 (N_3491,N_3193,N_3137);
nor U3492 (N_3492,N_3272,N_3140);
xor U3493 (N_3493,N_3203,N_3227);
or U3494 (N_3494,N_3283,N_3208);
nand U3495 (N_3495,N_3131,N_3093);
xnor U3496 (N_3496,N_3127,N_3185);
xnor U3497 (N_3497,N_3050,N_3026);
nor U3498 (N_3498,N_3013,N_3109);
nand U3499 (N_3499,N_3098,N_3099);
or U3500 (N_3500,N_3243,N_3123);
nand U3501 (N_3501,N_3052,N_3070);
and U3502 (N_3502,N_3141,N_3214);
xor U3503 (N_3503,N_3141,N_3225);
and U3504 (N_3504,N_3187,N_3060);
nand U3505 (N_3505,N_3022,N_3027);
and U3506 (N_3506,N_3261,N_3152);
or U3507 (N_3507,N_3057,N_3028);
nor U3508 (N_3508,N_3205,N_3007);
or U3509 (N_3509,N_3153,N_3264);
nor U3510 (N_3510,N_3249,N_3065);
and U3511 (N_3511,N_3007,N_3233);
or U3512 (N_3512,N_3118,N_3038);
xor U3513 (N_3513,N_3059,N_3015);
nor U3514 (N_3514,N_3280,N_3278);
or U3515 (N_3515,N_3177,N_3129);
nand U3516 (N_3516,N_3187,N_3228);
or U3517 (N_3517,N_3249,N_3204);
nand U3518 (N_3518,N_3270,N_3063);
and U3519 (N_3519,N_3134,N_3042);
or U3520 (N_3520,N_3259,N_3072);
and U3521 (N_3521,N_3165,N_3169);
xor U3522 (N_3522,N_3123,N_3151);
nor U3523 (N_3523,N_3105,N_3057);
nand U3524 (N_3524,N_3200,N_3088);
or U3525 (N_3525,N_3058,N_3060);
or U3526 (N_3526,N_3284,N_3299);
nor U3527 (N_3527,N_3149,N_3262);
nor U3528 (N_3528,N_3266,N_3136);
nand U3529 (N_3529,N_3077,N_3126);
nand U3530 (N_3530,N_3298,N_3051);
xnor U3531 (N_3531,N_3083,N_3124);
xnor U3532 (N_3532,N_3234,N_3035);
and U3533 (N_3533,N_3121,N_3032);
and U3534 (N_3534,N_3290,N_3153);
nor U3535 (N_3535,N_3287,N_3158);
xnor U3536 (N_3536,N_3104,N_3226);
nand U3537 (N_3537,N_3054,N_3107);
or U3538 (N_3538,N_3251,N_3255);
nor U3539 (N_3539,N_3091,N_3188);
and U3540 (N_3540,N_3082,N_3011);
xnor U3541 (N_3541,N_3256,N_3090);
or U3542 (N_3542,N_3006,N_3232);
or U3543 (N_3543,N_3174,N_3201);
and U3544 (N_3544,N_3000,N_3138);
nand U3545 (N_3545,N_3287,N_3131);
or U3546 (N_3546,N_3117,N_3280);
nand U3547 (N_3547,N_3103,N_3101);
and U3548 (N_3548,N_3203,N_3165);
xnor U3549 (N_3549,N_3056,N_3201);
nand U3550 (N_3550,N_3081,N_3023);
and U3551 (N_3551,N_3146,N_3082);
nand U3552 (N_3552,N_3071,N_3048);
and U3553 (N_3553,N_3136,N_3261);
or U3554 (N_3554,N_3055,N_3284);
nand U3555 (N_3555,N_3142,N_3164);
xnor U3556 (N_3556,N_3102,N_3025);
nor U3557 (N_3557,N_3223,N_3192);
and U3558 (N_3558,N_3107,N_3018);
nor U3559 (N_3559,N_3117,N_3243);
and U3560 (N_3560,N_3161,N_3107);
nand U3561 (N_3561,N_3042,N_3164);
xnor U3562 (N_3562,N_3054,N_3267);
or U3563 (N_3563,N_3257,N_3086);
nand U3564 (N_3564,N_3039,N_3294);
or U3565 (N_3565,N_3067,N_3079);
or U3566 (N_3566,N_3071,N_3106);
nor U3567 (N_3567,N_3195,N_3230);
nor U3568 (N_3568,N_3067,N_3225);
nor U3569 (N_3569,N_3100,N_3153);
xnor U3570 (N_3570,N_3128,N_3087);
nor U3571 (N_3571,N_3180,N_3212);
or U3572 (N_3572,N_3185,N_3188);
or U3573 (N_3573,N_3052,N_3116);
nand U3574 (N_3574,N_3038,N_3260);
nand U3575 (N_3575,N_3264,N_3272);
nor U3576 (N_3576,N_3056,N_3293);
xnor U3577 (N_3577,N_3107,N_3285);
xor U3578 (N_3578,N_3108,N_3210);
and U3579 (N_3579,N_3198,N_3107);
nand U3580 (N_3580,N_3080,N_3166);
nand U3581 (N_3581,N_3112,N_3064);
or U3582 (N_3582,N_3078,N_3246);
nor U3583 (N_3583,N_3135,N_3180);
or U3584 (N_3584,N_3111,N_3019);
and U3585 (N_3585,N_3164,N_3178);
or U3586 (N_3586,N_3095,N_3164);
nor U3587 (N_3587,N_3154,N_3265);
xor U3588 (N_3588,N_3243,N_3197);
xnor U3589 (N_3589,N_3225,N_3267);
or U3590 (N_3590,N_3074,N_3257);
or U3591 (N_3591,N_3159,N_3229);
nor U3592 (N_3592,N_3239,N_3044);
and U3593 (N_3593,N_3175,N_3211);
nand U3594 (N_3594,N_3181,N_3254);
xnor U3595 (N_3595,N_3288,N_3141);
nand U3596 (N_3596,N_3170,N_3254);
nor U3597 (N_3597,N_3031,N_3233);
and U3598 (N_3598,N_3158,N_3070);
xor U3599 (N_3599,N_3190,N_3001);
and U3600 (N_3600,N_3446,N_3457);
or U3601 (N_3601,N_3364,N_3490);
nand U3602 (N_3602,N_3318,N_3383);
nand U3603 (N_3603,N_3437,N_3333);
and U3604 (N_3604,N_3576,N_3548);
nor U3605 (N_3605,N_3420,N_3435);
xor U3606 (N_3606,N_3581,N_3355);
nand U3607 (N_3607,N_3413,N_3365);
nand U3608 (N_3608,N_3380,N_3505);
or U3609 (N_3609,N_3352,N_3343);
nand U3610 (N_3610,N_3478,N_3554);
or U3611 (N_3611,N_3479,N_3449);
nand U3612 (N_3612,N_3533,N_3538);
and U3613 (N_3613,N_3304,N_3350);
and U3614 (N_3614,N_3378,N_3376);
nand U3615 (N_3615,N_3509,N_3463);
nor U3616 (N_3616,N_3426,N_3442);
xnor U3617 (N_3617,N_3403,N_3521);
or U3618 (N_3618,N_3444,N_3360);
nand U3619 (N_3619,N_3312,N_3382);
or U3620 (N_3620,N_3408,N_3445);
nand U3621 (N_3621,N_3441,N_3329);
nor U3622 (N_3622,N_3520,N_3472);
nor U3623 (N_3623,N_3432,N_3402);
nand U3624 (N_3624,N_3356,N_3386);
nor U3625 (N_3625,N_3592,N_3323);
and U3626 (N_3626,N_3575,N_3315);
nand U3627 (N_3627,N_3436,N_3465);
nor U3628 (N_3628,N_3572,N_3341);
xor U3629 (N_3629,N_3532,N_3433);
or U3630 (N_3630,N_3443,N_3428);
and U3631 (N_3631,N_3307,N_3518);
and U3632 (N_3632,N_3534,N_3596);
nor U3633 (N_3633,N_3526,N_3547);
nor U3634 (N_3634,N_3543,N_3502);
xor U3635 (N_3635,N_3303,N_3394);
nand U3636 (N_3636,N_3368,N_3396);
or U3637 (N_3637,N_3302,N_3540);
xor U3638 (N_3638,N_3586,N_3527);
and U3639 (N_3639,N_3384,N_3359);
and U3640 (N_3640,N_3568,N_3473);
nor U3641 (N_3641,N_3489,N_3559);
nor U3642 (N_3642,N_3468,N_3392);
nand U3643 (N_3643,N_3582,N_3555);
and U3644 (N_3644,N_3460,N_3519);
nand U3645 (N_3645,N_3462,N_3504);
and U3646 (N_3646,N_3510,N_3499);
nand U3647 (N_3647,N_3388,N_3379);
nor U3648 (N_3648,N_3590,N_3390);
and U3649 (N_3649,N_3539,N_3372);
or U3650 (N_3650,N_3565,N_3567);
or U3651 (N_3651,N_3481,N_3599);
nor U3652 (N_3652,N_3589,N_3373);
or U3653 (N_3653,N_3497,N_3566);
nor U3654 (N_3654,N_3399,N_3531);
nor U3655 (N_3655,N_3588,N_3541);
nand U3656 (N_3656,N_3458,N_3546);
nand U3657 (N_3657,N_3471,N_3345);
and U3658 (N_3658,N_3553,N_3451);
or U3659 (N_3659,N_3366,N_3371);
and U3660 (N_3660,N_3524,N_3571);
xnor U3661 (N_3661,N_3484,N_3535);
nand U3662 (N_3662,N_3562,N_3339);
nor U3663 (N_3663,N_3337,N_3330);
nor U3664 (N_3664,N_3338,N_3585);
xnor U3665 (N_3665,N_3577,N_3529);
or U3666 (N_3666,N_3561,N_3331);
xnor U3667 (N_3667,N_3401,N_3453);
nand U3668 (N_3668,N_3447,N_3528);
nand U3669 (N_3669,N_3448,N_3503);
nand U3670 (N_3670,N_3459,N_3300);
or U3671 (N_3671,N_3517,N_3580);
xor U3672 (N_3672,N_3357,N_3421);
xor U3673 (N_3673,N_3557,N_3344);
xnor U3674 (N_3674,N_3369,N_3393);
or U3675 (N_3675,N_3439,N_3347);
and U3676 (N_3676,N_3487,N_3466);
nor U3677 (N_3677,N_3346,N_3310);
nor U3678 (N_3678,N_3370,N_3410);
xor U3679 (N_3679,N_3595,N_3507);
nand U3680 (N_3680,N_3587,N_3349);
and U3681 (N_3681,N_3563,N_3556);
nand U3682 (N_3682,N_3430,N_3573);
or U3683 (N_3683,N_3511,N_3427);
and U3684 (N_3684,N_3516,N_3361);
nor U3685 (N_3685,N_3407,N_3363);
nand U3686 (N_3686,N_3314,N_3486);
or U3687 (N_3687,N_3464,N_3354);
nand U3688 (N_3688,N_3501,N_3334);
nor U3689 (N_3689,N_3362,N_3377);
nand U3690 (N_3690,N_3498,N_3381);
and U3691 (N_3691,N_3415,N_3579);
nor U3692 (N_3692,N_3597,N_3305);
xor U3693 (N_3693,N_3313,N_3574);
xnor U3694 (N_3694,N_3508,N_3454);
nand U3695 (N_3695,N_3494,N_3391);
and U3696 (N_3696,N_3523,N_3308);
xor U3697 (N_3697,N_3423,N_3536);
nor U3698 (N_3698,N_3405,N_3429);
or U3699 (N_3699,N_3434,N_3340);
and U3700 (N_3700,N_3594,N_3422);
xor U3701 (N_3701,N_3450,N_3500);
or U3702 (N_3702,N_3467,N_3414);
nand U3703 (N_3703,N_3475,N_3438);
nand U3704 (N_3704,N_3584,N_3409);
or U3705 (N_3705,N_3456,N_3469);
or U3706 (N_3706,N_3316,N_3387);
xnor U3707 (N_3707,N_3431,N_3474);
xnor U3708 (N_3708,N_3375,N_3406);
or U3709 (N_3709,N_3425,N_3542);
xnor U3710 (N_3710,N_3358,N_3417);
or U3711 (N_3711,N_3322,N_3496);
xnor U3712 (N_3712,N_3424,N_3537);
xor U3713 (N_3713,N_3558,N_3353);
xnor U3714 (N_3714,N_3560,N_3514);
nor U3715 (N_3715,N_3583,N_3351);
xor U3716 (N_3716,N_3327,N_3335);
xor U3717 (N_3717,N_3564,N_3591);
nand U3718 (N_3718,N_3321,N_3477);
xor U3719 (N_3719,N_3480,N_3492);
nand U3720 (N_3720,N_3326,N_3495);
nor U3721 (N_3721,N_3404,N_3512);
nor U3722 (N_3722,N_3549,N_3325);
xnor U3723 (N_3723,N_3385,N_3530);
or U3724 (N_3724,N_3395,N_3348);
or U3725 (N_3725,N_3455,N_3522);
xnor U3726 (N_3726,N_3398,N_3389);
nor U3727 (N_3727,N_3342,N_3470);
or U3728 (N_3728,N_3461,N_3570);
nor U3729 (N_3729,N_3476,N_3452);
xnor U3730 (N_3730,N_3598,N_3515);
nor U3731 (N_3731,N_3552,N_3306);
and U3732 (N_3732,N_3400,N_3419);
nand U3733 (N_3733,N_3488,N_3317);
and U3734 (N_3734,N_3411,N_3491);
or U3735 (N_3735,N_3506,N_3569);
or U3736 (N_3736,N_3544,N_3550);
or U3737 (N_3737,N_3324,N_3336);
nor U3738 (N_3738,N_3309,N_3513);
xnor U3739 (N_3739,N_3367,N_3551);
or U3740 (N_3740,N_3482,N_3483);
nand U3741 (N_3741,N_3412,N_3525);
xnor U3742 (N_3742,N_3320,N_3332);
nor U3743 (N_3743,N_3397,N_3418);
xnor U3744 (N_3744,N_3416,N_3493);
and U3745 (N_3745,N_3485,N_3319);
or U3746 (N_3746,N_3440,N_3328);
or U3747 (N_3747,N_3578,N_3301);
and U3748 (N_3748,N_3545,N_3374);
and U3749 (N_3749,N_3593,N_3311);
and U3750 (N_3750,N_3507,N_3445);
and U3751 (N_3751,N_3480,N_3376);
nor U3752 (N_3752,N_3574,N_3358);
or U3753 (N_3753,N_3492,N_3439);
xnor U3754 (N_3754,N_3565,N_3410);
or U3755 (N_3755,N_3455,N_3490);
xor U3756 (N_3756,N_3320,N_3457);
xor U3757 (N_3757,N_3326,N_3456);
or U3758 (N_3758,N_3482,N_3540);
nor U3759 (N_3759,N_3492,N_3420);
and U3760 (N_3760,N_3536,N_3508);
and U3761 (N_3761,N_3530,N_3401);
xor U3762 (N_3762,N_3560,N_3583);
nor U3763 (N_3763,N_3425,N_3308);
nor U3764 (N_3764,N_3478,N_3580);
nand U3765 (N_3765,N_3570,N_3474);
nand U3766 (N_3766,N_3433,N_3472);
and U3767 (N_3767,N_3571,N_3331);
xor U3768 (N_3768,N_3301,N_3415);
xnor U3769 (N_3769,N_3553,N_3324);
and U3770 (N_3770,N_3488,N_3593);
xor U3771 (N_3771,N_3454,N_3450);
xnor U3772 (N_3772,N_3469,N_3569);
and U3773 (N_3773,N_3523,N_3427);
xnor U3774 (N_3774,N_3537,N_3577);
nor U3775 (N_3775,N_3368,N_3385);
xor U3776 (N_3776,N_3544,N_3362);
or U3777 (N_3777,N_3476,N_3418);
nand U3778 (N_3778,N_3408,N_3337);
xor U3779 (N_3779,N_3572,N_3411);
xor U3780 (N_3780,N_3553,N_3466);
nor U3781 (N_3781,N_3326,N_3413);
or U3782 (N_3782,N_3382,N_3483);
xnor U3783 (N_3783,N_3506,N_3459);
nor U3784 (N_3784,N_3504,N_3527);
nor U3785 (N_3785,N_3338,N_3535);
and U3786 (N_3786,N_3486,N_3302);
nand U3787 (N_3787,N_3386,N_3588);
or U3788 (N_3788,N_3529,N_3512);
nand U3789 (N_3789,N_3472,N_3490);
or U3790 (N_3790,N_3596,N_3360);
xnor U3791 (N_3791,N_3344,N_3551);
or U3792 (N_3792,N_3478,N_3352);
nor U3793 (N_3793,N_3563,N_3536);
nand U3794 (N_3794,N_3499,N_3408);
nor U3795 (N_3795,N_3514,N_3326);
and U3796 (N_3796,N_3452,N_3482);
nor U3797 (N_3797,N_3320,N_3474);
or U3798 (N_3798,N_3406,N_3337);
nor U3799 (N_3799,N_3578,N_3472);
nand U3800 (N_3800,N_3313,N_3514);
nor U3801 (N_3801,N_3362,N_3457);
nor U3802 (N_3802,N_3552,N_3323);
xor U3803 (N_3803,N_3317,N_3309);
nand U3804 (N_3804,N_3410,N_3481);
nor U3805 (N_3805,N_3494,N_3434);
and U3806 (N_3806,N_3391,N_3589);
or U3807 (N_3807,N_3578,N_3548);
or U3808 (N_3808,N_3450,N_3425);
and U3809 (N_3809,N_3498,N_3517);
or U3810 (N_3810,N_3567,N_3458);
and U3811 (N_3811,N_3401,N_3576);
and U3812 (N_3812,N_3329,N_3497);
and U3813 (N_3813,N_3421,N_3380);
xnor U3814 (N_3814,N_3349,N_3483);
nor U3815 (N_3815,N_3517,N_3578);
nor U3816 (N_3816,N_3327,N_3546);
xnor U3817 (N_3817,N_3368,N_3540);
or U3818 (N_3818,N_3429,N_3430);
xor U3819 (N_3819,N_3441,N_3492);
or U3820 (N_3820,N_3302,N_3307);
xor U3821 (N_3821,N_3313,N_3441);
nand U3822 (N_3822,N_3337,N_3516);
nor U3823 (N_3823,N_3596,N_3586);
xor U3824 (N_3824,N_3486,N_3329);
and U3825 (N_3825,N_3453,N_3593);
xnor U3826 (N_3826,N_3317,N_3346);
and U3827 (N_3827,N_3442,N_3369);
nand U3828 (N_3828,N_3567,N_3405);
nor U3829 (N_3829,N_3318,N_3561);
nor U3830 (N_3830,N_3465,N_3406);
xor U3831 (N_3831,N_3539,N_3475);
xnor U3832 (N_3832,N_3507,N_3348);
and U3833 (N_3833,N_3378,N_3362);
xnor U3834 (N_3834,N_3433,N_3465);
nand U3835 (N_3835,N_3486,N_3434);
or U3836 (N_3836,N_3405,N_3562);
or U3837 (N_3837,N_3352,N_3494);
or U3838 (N_3838,N_3520,N_3459);
or U3839 (N_3839,N_3571,N_3552);
nand U3840 (N_3840,N_3530,N_3333);
nand U3841 (N_3841,N_3301,N_3549);
xnor U3842 (N_3842,N_3564,N_3460);
xor U3843 (N_3843,N_3535,N_3417);
nand U3844 (N_3844,N_3379,N_3361);
nor U3845 (N_3845,N_3303,N_3467);
nand U3846 (N_3846,N_3533,N_3458);
xor U3847 (N_3847,N_3325,N_3302);
xor U3848 (N_3848,N_3393,N_3555);
nand U3849 (N_3849,N_3495,N_3450);
xnor U3850 (N_3850,N_3488,N_3520);
nand U3851 (N_3851,N_3419,N_3350);
xnor U3852 (N_3852,N_3521,N_3390);
and U3853 (N_3853,N_3508,N_3426);
or U3854 (N_3854,N_3513,N_3486);
xor U3855 (N_3855,N_3306,N_3533);
nor U3856 (N_3856,N_3365,N_3524);
nor U3857 (N_3857,N_3393,N_3423);
nor U3858 (N_3858,N_3404,N_3380);
nor U3859 (N_3859,N_3515,N_3358);
xnor U3860 (N_3860,N_3371,N_3421);
nor U3861 (N_3861,N_3569,N_3594);
or U3862 (N_3862,N_3393,N_3501);
xnor U3863 (N_3863,N_3438,N_3391);
nor U3864 (N_3864,N_3527,N_3339);
xor U3865 (N_3865,N_3312,N_3585);
or U3866 (N_3866,N_3375,N_3508);
nand U3867 (N_3867,N_3470,N_3567);
nand U3868 (N_3868,N_3452,N_3395);
and U3869 (N_3869,N_3391,N_3428);
or U3870 (N_3870,N_3409,N_3427);
or U3871 (N_3871,N_3546,N_3308);
nand U3872 (N_3872,N_3313,N_3579);
or U3873 (N_3873,N_3525,N_3508);
nand U3874 (N_3874,N_3533,N_3570);
or U3875 (N_3875,N_3309,N_3349);
and U3876 (N_3876,N_3350,N_3556);
xor U3877 (N_3877,N_3565,N_3341);
and U3878 (N_3878,N_3599,N_3431);
xor U3879 (N_3879,N_3445,N_3406);
or U3880 (N_3880,N_3417,N_3368);
or U3881 (N_3881,N_3568,N_3575);
xnor U3882 (N_3882,N_3506,N_3524);
or U3883 (N_3883,N_3426,N_3399);
nand U3884 (N_3884,N_3477,N_3560);
nor U3885 (N_3885,N_3590,N_3395);
or U3886 (N_3886,N_3349,N_3550);
nor U3887 (N_3887,N_3354,N_3381);
and U3888 (N_3888,N_3388,N_3501);
or U3889 (N_3889,N_3459,N_3492);
and U3890 (N_3890,N_3456,N_3510);
nor U3891 (N_3891,N_3476,N_3539);
nor U3892 (N_3892,N_3391,N_3317);
xnor U3893 (N_3893,N_3399,N_3582);
xnor U3894 (N_3894,N_3407,N_3316);
and U3895 (N_3895,N_3370,N_3408);
xnor U3896 (N_3896,N_3457,N_3385);
xor U3897 (N_3897,N_3425,N_3443);
nor U3898 (N_3898,N_3412,N_3476);
xnor U3899 (N_3899,N_3515,N_3487);
and U3900 (N_3900,N_3661,N_3683);
and U3901 (N_3901,N_3721,N_3863);
xor U3902 (N_3902,N_3899,N_3797);
nor U3903 (N_3903,N_3849,N_3764);
or U3904 (N_3904,N_3763,N_3774);
xnor U3905 (N_3905,N_3719,N_3673);
nand U3906 (N_3906,N_3823,N_3881);
and U3907 (N_3907,N_3613,N_3716);
nand U3908 (N_3908,N_3704,N_3884);
and U3909 (N_3909,N_3694,N_3648);
nand U3910 (N_3910,N_3846,N_3800);
xnor U3911 (N_3911,N_3713,N_3795);
or U3912 (N_3912,N_3816,N_3814);
or U3913 (N_3913,N_3640,N_3853);
and U3914 (N_3914,N_3778,N_3844);
nor U3915 (N_3915,N_3717,N_3618);
nor U3916 (N_3916,N_3788,N_3867);
and U3917 (N_3917,N_3865,N_3631);
nand U3918 (N_3918,N_3862,N_3799);
or U3919 (N_3919,N_3645,N_3748);
or U3920 (N_3920,N_3866,N_3610);
nor U3921 (N_3921,N_3670,N_3776);
nor U3922 (N_3922,N_3824,N_3883);
xor U3923 (N_3923,N_3811,N_3808);
nand U3924 (N_3924,N_3680,N_3761);
nand U3925 (N_3925,N_3890,N_3607);
nor U3926 (N_3926,N_3871,N_3681);
nor U3927 (N_3927,N_3757,N_3747);
or U3928 (N_3928,N_3741,N_3665);
nand U3929 (N_3929,N_3635,N_3619);
or U3930 (N_3930,N_3633,N_3718);
nor U3931 (N_3931,N_3767,N_3662);
or U3932 (N_3932,N_3813,N_3664);
xor U3933 (N_3933,N_3628,N_3622);
or U3934 (N_3934,N_3655,N_3775);
nor U3935 (N_3935,N_3707,N_3609);
xor U3936 (N_3936,N_3892,N_3700);
or U3937 (N_3937,N_3732,N_3627);
or U3938 (N_3938,N_3658,N_3620);
or U3939 (N_3939,N_3724,N_3705);
nor U3940 (N_3940,N_3897,N_3818);
or U3941 (N_3941,N_3854,N_3752);
or U3942 (N_3942,N_3848,N_3789);
or U3943 (N_3943,N_3603,N_3843);
nand U3944 (N_3944,N_3829,N_3838);
and U3945 (N_3945,N_3787,N_3750);
nor U3946 (N_3946,N_3731,N_3698);
or U3947 (N_3947,N_3817,N_3842);
nand U3948 (N_3948,N_3668,N_3671);
nand U3949 (N_3949,N_3855,N_3651);
xor U3950 (N_3950,N_3638,N_3803);
and U3951 (N_3951,N_3807,N_3879);
or U3952 (N_3952,N_3793,N_3687);
or U3953 (N_3953,N_3647,N_3674);
nand U3954 (N_3954,N_3754,N_3758);
or U3955 (N_3955,N_3784,N_3737);
xor U3956 (N_3956,N_3768,N_3790);
or U3957 (N_3957,N_3804,N_3659);
nand U3958 (N_3958,N_3637,N_3765);
nand U3959 (N_3959,N_3669,N_3735);
and U3960 (N_3960,N_3749,N_3895);
nand U3961 (N_3961,N_3810,N_3812);
nor U3962 (N_3962,N_3692,N_3682);
and U3963 (N_3963,N_3623,N_3828);
xnor U3964 (N_3964,N_3699,N_3860);
xnor U3965 (N_3965,N_3835,N_3714);
nand U3966 (N_3966,N_3891,N_3760);
and U3967 (N_3967,N_3792,N_3858);
or U3968 (N_3968,N_3887,N_3825);
nand U3969 (N_3969,N_3771,N_3832);
and U3970 (N_3970,N_3857,N_3781);
nor U3971 (N_3971,N_3802,N_3880);
nand U3972 (N_3972,N_3872,N_3801);
or U3973 (N_3973,N_3606,N_3734);
nor U3974 (N_3974,N_3755,N_3690);
or U3975 (N_3975,N_3696,N_3739);
and U3976 (N_3976,N_3822,N_3675);
nand U3977 (N_3977,N_3644,N_3605);
or U3978 (N_3978,N_3614,N_3753);
nor U3979 (N_3979,N_3723,N_3710);
nand U3980 (N_3980,N_3695,N_3602);
and U3981 (N_3981,N_3646,N_3746);
nand U3982 (N_3982,N_3634,N_3851);
and U3983 (N_3983,N_3679,N_3780);
nand U3984 (N_3984,N_3888,N_3654);
and U3985 (N_3985,N_3821,N_3621);
or U3986 (N_3986,N_3666,N_3685);
and U3987 (N_3987,N_3702,N_3672);
and U3988 (N_3988,N_3629,N_3711);
or U3989 (N_3989,N_3736,N_3726);
and U3990 (N_3990,N_3762,N_3641);
xor U3991 (N_3991,N_3684,N_3738);
and U3992 (N_3992,N_3625,N_3652);
and U3993 (N_3993,N_3712,N_3770);
nand U3994 (N_3994,N_3691,N_3756);
nand U3995 (N_3995,N_3663,N_3894);
nand U3996 (N_3996,N_3727,N_3820);
xnor U3997 (N_3997,N_3831,N_3836);
nor U3998 (N_3998,N_3861,N_3678);
nor U3999 (N_3999,N_3882,N_3885);
nor U4000 (N_4000,N_3677,N_3856);
and U4001 (N_4001,N_3751,N_3656);
and U4002 (N_4002,N_3773,N_3786);
nand U4003 (N_4003,N_3772,N_3600);
and U4004 (N_4004,N_3850,N_3722);
nand U4005 (N_4005,N_3688,N_3777);
nor U4006 (N_4006,N_3632,N_3604);
nor U4007 (N_4007,N_3834,N_3859);
and U4008 (N_4008,N_3745,N_3806);
or U4009 (N_4009,N_3870,N_3794);
or U4010 (N_4010,N_3759,N_3798);
xnor U4011 (N_4011,N_3611,N_3877);
nor U4012 (N_4012,N_3733,N_3676);
nor U4013 (N_4013,N_3827,N_3782);
xor U4014 (N_4014,N_3624,N_3839);
xnor U4015 (N_4015,N_3686,N_3689);
nand U4016 (N_4016,N_3706,N_3819);
or U4017 (N_4017,N_3608,N_3601);
or U4018 (N_4018,N_3805,N_3630);
nand U4019 (N_4019,N_3626,N_3657);
nand U4020 (N_4020,N_3660,N_3703);
nor U4021 (N_4021,N_3869,N_3649);
xor U4022 (N_4022,N_3639,N_3725);
or U4023 (N_4023,N_3876,N_3616);
xor U4024 (N_4024,N_3868,N_3847);
xnor U4025 (N_4025,N_3667,N_3833);
nand U4026 (N_4026,N_3837,N_3715);
and U4027 (N_4027,N_3809,N_3896);
nand U4028 (N_4028,N_3728,N_3643);
and U4029 (N_4029,N_3785,N_3766);
xnor U4030 (N_4030,N_3612,N_3815);
or U4031 (N_4031,N_3653,N_3796);
and U4032 (N_4032,N_3791,N_3893);
or U4033 (N_4033,N_3873,N_3840);
nand U4034 (N_4034,N_3886,N_3742);
xnor U4035 (N_4035,N_3701,N_3898);
nor U4036 (N_4036,N_3642,N_3779);
nor U4037 (N_4037,N_3830,N_3720);
or U4038 (N_4038,N_3709,N_3878);
nor U4039 (N_4039,N_3617,N_3615);
nor U4040 (N_4040,N_3852,N_3783);
or U4041 (N_4041,N_3743,N_3889);
nand U4042 (N_4042,N_3826,N_3845);
or U4043 (N_4043,N_3730,N_3693);
and U4044 (N_4044,N_3864,N_3650);
or U4045 (N_4045,N_3708,N_3636);
and U4046 (N_4046,N_3769,N_3740);
xnor U4047 (N_4047,N_3875,N_3874);
nor U4048 (N_4048,N_3744,N_3729);
nor U4049 (N_4049,N_3697,N_3841);
or U4050 (N_4050,N_3698,N_3773);
nand U4051 (N_4051,N_3821,N_3798);
nor U4052 (N_4052,N_3862,N_3711);
xnor U4053 (N_4053,N_3850,N_3710);
and U4054 (N_4054,N_3792,N_3896);
or U4055 (N_4055,N_3677,N_3704);
nand U4056 (N_4056,N_3855,N_3742);
nand U4057 (N_4057,N_3611,N_3710);
or U4058 (N_4058,N_3864,N_3758);
and U4059 (N_4059,N_3899,N_3729);
nor U4060 (N_4060,N_3645,N_3847);
and U4061 (N_4061,N_3832,N_3702);
and U4062 (N_4062,N_3846,N_3657);
nand U4063 (N_4063,N_3825,N_3765);
and U4064 (N_4064,N_3601,N_3665);
or U4065 (N_4065,N_3676,N_3768);
xor U4066 (N_4066,N_3691,N_3840);
or U4067 (N_4067,N_3892,N_3720);
and U4068 (N_4068,N_3888,N_3866);
nand U4069 (N_4069,N_3713,N_3658);
or U4070 (N_4070,N_3607,N_3809);
and U4071 (N_4071,N_3803,N_3766);
or U4072 (N_4072,N_3861,N_3892);
xnor U4073 (N_4073,N_3750,N_3756);
and U4074 (N_4074,N_3650,N_3860);
nand U4075 (N_4075,N_3621,N_3778);
nand U4076 (N_4076,N_3851,N_3659);
nor U4077 (N_4077,N_3734,N_3615);
nand U4078 (N_4078,N_3621,N_3653);
nand U4079 (N_4079,N_3802,N_3734);
and U4080 (N_4080,N_3714,N_3754);
or U4081 (N_4081,N_3706,N_3767);
xor U4082 (N_4082,N_3830,N_3600);
and U4083 (N_4083,N_3658,N_3663);
and U4084 (N_4084,N_3730,N_3867);
and U4085 (N_4085,N_3899,N_3845);
xnor U4086 (N_4086,N_3840,N_3693);
nand U4087 (N_4087,N_3880,N_3623);
and U4088 (N_4088,N_3883,N_3859);
nor U4089 (N_4089,N_3844,N_3638);
or U4090 (N_4090,N_3717,N_3870);
nor U4091 (N_4091,N_3700,N_3756);
nor U4092 (N_4092,N_3806,N_3835);
xor U4093 (N_4093,N_3628,N_3738);
nor U4094 (N_4094,N_3773,N_3751);
or U4095 (N_4095,N_3831,N_3601);
nand U4096 (N_4096,N_3867,N_3702);
and U4097 (N_4097,N_3785,N_3869);
xor U4098 (N_4098,N_3749,N_3636);
nand U4099 (N_4099,N_3680,N_3853);
xnor U4100 (N_4100,N_3658,N_3714);
nor U4101 (N_4101,N_3789,N_3697);
and U4102 (N_4102,N_3883,N_3664);
xor U4103 (N_4103,N_3819,N_3862);
and U4104 (N_4104,N_3822,N_3793);
or U4105 (N_4105,N_3691,N_3634);
nand U4106 (N_4106,N_3887,N_3737);
and U4107 (N_4107,N_3748,N_3740);
and U4108 (N_4108,N_3604,N_3667);
nand U4109 (N_4109,N_3760,N_3658);
and U4110 (N_4110,N_3773,N_3772);
nor U4111 (N_4111,N_3651,N_3657);
nand U4112 (N_4112,N_3821,N_3667);
or U4113 (N_4113,N_3788,N_3896);
nand U4114 (N_4114,N_3740,N_3760);
xnor U4115 (N_4115,N_3886,N_3633);
nand U4116 (N_4116,N_3848,N_3752);
xor U4117 (N_4117,N_3804,N_3747);
xor U4118 (N_4118,N_3813,N_3889);
xor U4119 (N_4119,N_3788,N_3636);
or U4120 (N_4120,N_3867,N_3843);
xnor U4121 (N_4121,N_3770,N_3703);
nor U4122 (N_4122,N_3736,N_3660);
and U4123 (N_4123,N_3779,N_3657);
and U4124 (N_4124,N_3764,N_3795);
and U4125 (N_4125,N_3835,N_3821);
or U4126 (N_4126,N_3777,N_3840);
nor U4127 (N_4127,N_3867,N_3736);
nand U4128 (N_4128,N_3685,N_3778);
or U4129 (N_4129,N_3648,N_3722);
xor U4130 (N_4130,N_3747,N_3845);
or U4131 (N_4131,N_3635,N_3627);
nand U4132 (N_4132,N_3899,N_3791);
xor U4133 (N_4133,N_3844,N_3741);
nor U4134 (N_4134,N_3683,N_3868);
or U4135 (N_4135,N_3877,N_3886);
nand U4136 (N_4136,N_3801,N_3847);
or U4137 (N_4137,N_3798,N_3823);
and U4138 (N_4138,N_3791,N_3753);
or U4139 (N_4139,N_3778,N_3704);
and U4140 (N_4140,N_3663,N_3784);
nor U4141 (N_4141,N_3735,N_3653);
nor U4142 (N_4142,N_3710,N_3738);
nor U4143 (N_4143,N_3723,N_3747);
xnor U4144 (N_4144,N_3602,N_3786);
and U4145 (N_4145,N_3611,N_3640);
xnor U4146 (N_4146,N_3692,N_3697);
or U4147 (N_4147,N_3637,N_3790);
nor U4148 (N_4148,N_3848,N_3763);
and U4149 (N_4149,N_3636,N_3772);
and U4150 (N_4150,N_3653,N_3650);
nand U4151 (N_4151,N_3679,N_3880);
nand U4152 (N_4152,N_3866,N_3648);
and U4153 (N_4153,N_3670,N_3881);
or U4154 (N_4154,N_3674,N_3778);
and U4155 (N_4155,N_3796,N_3728);
nor U4156 (N_4156,N_3632,N_3819);
xor U4157 (N_4157,N_3634,N_3619);
nor U4158 (N_4158,N_3755,N_3833);
xnor U4159 (N_4159,N_3689,N_3632);
nor U4160 (N_4160,N_3812,N_3642);
and U4161 (N_4161,N_3610,N_3879);
and U4162 (N_4162,N_3808,N_3616);
nor U4163 (N_4163,N_3721,N_3643);
and U4164 (N_4164,N_3739,N_3769);
and U4165 (N_4165,N_3772,N_3778);
or U4166 (N_4166,N_3801,N_3677);
or U4167 (N_4167,N_3750,N_3614);
and U4168 (N_4168,N_3852,N_3881);
and U4169 (N_4169,N_3876,N_3728);
xnor U4170 (N_4170,N_3706,N_3638);
and U4171 (N_4171,N_3702,N_3857);
xor U4172 (N_4172,N_3827,N_3847);
or U4173 (N_4173,N_3682,N_3777);
and U4174 (N_4174,N_3782,N_3751);
and U4175 (N_4175,N_3605,N_3870);
nand U4176 (N_4176,N_3633,N_3637);
or U4177 (N_4177,N_3808,N_3845);
nor U4178 (N_4178,N_3844,N_3801);
or U4179 (N_4179,N_3633,N_3846);
and U4180 (N_4180,N_3704,N_3782);
nand U4181 (N_4181,N_3897,N_3867);
nand U4182 (N_4182,N_3656,N_3607);
nor U4183 (N_4183,N_3871,N_3683);
or U4184 (N_4184,N_3839,N_3674);
or U4185 (N_4185,N_3894,N_3849);
and U4186 (N_4186,N_3620,N_3731);
xnor U4187 (N_4187,N_3752,N_3755);
xor U4188 (N_4188,N_3810,N_3641);
and U4189 (N_4189,N_3705,N_3804);
nor U4190 (N_4190,N_3810,N_3808);
xnor U4191 (N_4191,N_3744,N_3609);
and U4192 (N_4192,N_3655,N_3761);
xnor U4193 (N_4193,N_3723,N_3813);
xnor U4194 (N_4194,N_3692,N_3647);
nor U4195 (N_4195,N_3669,N_3706);
nand U4196 (N_4196,N_3786,N_3802);
nand U4197 (N_4197,N_3748,N_3791);
and U4198 (N_4198,N_3635,N_3755);
or U4199 (N_4199,N_3827,N_3710);
and U4200 (N_4200,N_4194,N_4034);
and U4201 (N_4201,N_4106,N_4042);
nand U4202 (N_4202,N_3977,N_4171);
nor U4203 (N_4203,N_3922,N_3991);
nor U4204 (N_4204,N_4158,N_4015);
nand U4205 (N_4205,N_4109,N_3947);
nand U4206 (N_4206,N_4146,N_3913);
or U4207 (N_4207,N_4011,N_4001);
nand U4208 (N_4208,N_4067,N_4073);
nand U4209 (N_4209,N_3924,N_3934);
xnor U4210 (N_4210,N_3933,N_3952);
nor U4211 (N_4211,N_4174,N_3910);
and U4212 (N_4212,N_4163,N_3902);
nor U4213 (N_4213,N_4177,N_4003);
nor U4214 (N_4214,N_3918,N_3937);
nand U4215 (N_4215,N_4130,N_4120);
xnor U4216 (N_4216,N_3945,N_4085);
xnor U4217 (N_4217,N_4184,N_3905);
and U4218 (N_4218,N_4033,N_4024);
nand U4219 (N_4219,N_4028,N_3917);
nor U4220 (N_4220,N_4164,N_3983);
xor U4221 (N_4221,N_4172,N_4114);
nand U4222 (N_4222,N_3981,N_3916);
and U4223 (N_4223,N_3963,N_3968);
nand U4224 (N_4224,N_4117,N_4064);
xnor U4225 (N_4225,N_3969,N_4013);
and U4226 (N_4226,N_4105,N_4099);
and U4227 (N_4227,N_3962,N_4111);
nand U4228 (N_4228,N_4090,N_3985);
nor U4229 (N_4229,N_4144,N_4168);
nand U4230 (N_4230,N_4170,N_4197);
nor U4231 (N_4231,N_4190,N_4176);
or U4232 (N_4232,N_4062,N_4089);
nand U4233 (N_4233,N_3966,N_3976);
or U4234 (N_4234,N_4094,N_4103);
xnor U4235 (N_4235,N_3992,N_3927);
nor U4236 (N_4236,N_3928,N_4093);
or U4237 (N_4237,N_4151,N_4128);
and U4238 (N_4238,N_3919,N_4022);
nand U4239 (N_4239,N_4101,N_3939);
and U4240 (N_4240,N_4083,N_3958);
and U4241 (N_4241,N_4155,N_3929);
nor U4242 (N_4242,N_3989,N_4115);
nor U4243 (N_4243,N_4084,N_3950);
and U4244 (N_4244,N_3948,N_4110);
xnor U4245 (N_4245,N_3974,N_4178);
or U4246 (N_4246,N_3996,N_4020);
xnor U4247 (N_4247,N_3954,N_4188);
nand U4248 (N_4248,N_4167,N_3912);
nand U4249 (N_4249,N_3904,N_3941);
and U4250 (N_4250,N_4199,N_4198);
nor U4251 (N_4251,N_3970,N_4021);
nand U4252 (N_4252,N_3923,N_4100);
and U4253 (N_4253,N_4157,N_4133);
xor U4254 (N_4254,N_4112,N_4162);
nor U4255 (N_4255,N_4192,N_4107);
and U4256 (N_4256,N_3907,N_4012);
nor U4257 (N_4257,N_4060,N_4049);
nor U4258 (N_4258,N_4180,N_4179);
or U4259 (N_4259,N_4145,N_3959);
or U4260 (N_4260,N_4082,N_4059);
nand U4261 (N_4261,N_4023,N_4029);
xnor U4262 (N_4262,N_4113,N_4087);
nand U4263 (N_4263,N_4069,N_4074);
and U4264 (N_4264,N_3926,N_3901);
or U4265 (N_4265,N_3932,N_4196);
nand U4266 (N_4266,N_4104,N_4159);
nand U4267 (N_4267,N_4027,N_4143);
xor U4268 (N_4268,N_4142,N_3957);
or U4269 (N_4269,N_4102,N_3915);
nand U4270 (N_4270,N_4149,N_4131);
nor U4271 (N_4271,N_4035,N_4005);
nand U4272 (N_4272,N_4169,N_4116);
and U4273 (N_4273,N_4135,N_4006);
xor U4274 (N_4274,N_4019,N_3984);
and U4275 (N_4275,N_4055,N_4056);
and U4276 (N_4276,N_3925,N_3909);
nor U4277 (N_4277,N_3956,N_4129);
nor U4278 (N_4278,N_3990,N_4095);
or U4279 (N_4279,N_4193,N_4044);
xor U4280 (N_4280,N_4008,N_4123);
xnor U4281 (N_4281,N_3982,N_4191);
or U4282 (N_4282,N_3936,N_3942);
and U4283 (N_4283,N_3906,N_4124);
nor U4284 (N_4284,N_3972,N_3949);
and U4285 (N_4285,N_4000,N_3980);
and U4286 (N_4286,N_4092,N_3999);
xnor U4287 (N_4287,N_4004,N_4166);
or U4288 (N_4288,N_4052,N_3943);
nand U4289 (N_4289,N_4010,N_4043);
nand U4290 (N_4290,N_4121,N_3979);
nor U4291 (N_4291,N_3995,N_4160);
or U4292 (N_4292,N_4076,N_4061);
nor U4293 (N_4293,N_3944,N_3965);
nor U4294 (N_4294,N_4071,N_3993);
and U4295 (N_4295,N_4014,N_4185);
xor U4296 (N_4296,N_3997,N_4016);
xnor U4297 (N_4297,N_4119,N_4081);
and U4298 (N_4298,N_4031,N_3971);
nand U4299 (N_4299,N_4118,N_4195);
nor U4300 (N_4300,N_3908,N_4141);
and U4301 (N_4301,N_3987,N_4053);
nand U4302 (N_4302,N_4097,N_4039);
nand U4303 (N_4303,N_4054,N_4173);
nand U4304 (N_4304,N_3994,N_4091);
and U4305 (N_4305,N_4108,N_4136);
nor U4306 (N_4306,N_3903,N_3955);
nor U4307 (N_4307,N_3986,N_3938);
xor U4308 (N_4308,N_4078,N_4080);
and U4309 (N_4309,N_4048,N_4046);
nand U4310 (N_4310,N_4051,N_4018);
nand U4311 (N_4311,N_4009,N_4150);
nand U4312 (N_4312,N_3960,N_4189);
nand U4313 (N_4313,N_3911,N_4047);
xor U4314 (N_4314,N_4086,N_3940);
nor U4315 (N_4315,N_3935,N_4139);
nor U4316 (N_4316,N_4077,N_4138);
nand U4317 (N_4317,N_3998,N_3921);
and U4318 (N_4318,N_4068,N_4122);
nor U4319 (N_4319,N_3914,N_4137);
xnor U4320 (N_4320,N_4079,N_4058);
xnor U4321 (N_4321,N_4187,N_4057);
or U4322 (N_4322,N_4147,N_4183);
nor U4323 (N_4323,N_3953,N_4007);
nand U4324 (N_4324,N_4026,N_4030);
and U4325 (N_4325,N_4127,N_4156);
nor U4326 (N_4326,N_4072,N_3978);
nor U4327 (N_4327,N_3900,N_3973);
or U4328 (N_4328,N_3946,N_4140);
nand U4329 (N_4329,N_4037,N_4025);
and U4330 (N_4330,N_4125,N_4041);
xnor U4331 (N_4331,N_4066,N_4161);
or U4332 (N_4332,N_4098,N_4132);
nor U4333 (N_4333,N_3967,N_4070);
and U4334 (N_4334,N_4134,N_4050);
and U4335 (N_4335,N_4126,N_4154);
xnor U4336 (N_4336,N_4065,N_4088);
and U4337 (N_4337,N_4038,N_4148);
or U4338 (N_4338,N_4096,N_3961);
nor U4339 (N_4339,N_4040,N_3975);
and U4340 (N_4340,N_4165,N_3951);
and U4341 (N_4341,N_4186,N_4153);
nand U4342 (N_4342,N_4182,N_4002);
xor U4343 (N_4343,N_4036,N_3988);
nor U4344 (N_4344,N_4175,N_4017);
nor U4345 (N_4345,N_3920,N_3930);
nand U4346 (N_4346,N_4045,N_4152);
xnor U4347 (N_4347,N_4075,N_4063);
xor U4348 (N_4348,N_4032,N_3964);
or U4349 (N_4349,N_3931,N_4181);
and U4350 (N_4350,N_4045,N_4005);
or U4351 (N_4351,N_3943,N_4194);
nand U4352 (N_4352,N_3982,N_3938);
xor U4353 (N_4353,N_4170,N_4116);
xor U4354 (N_4354,N_4048,N_4042);
xor U4355 (N_4355,N_4000,N_4083);
and U4356 (N_4356,N_4062,N_3942);
or U4357 (N_4357,N_3961,N_3995);
or U4358 (N_4358,N_4141,N_4105);
nand U4359 (N_4359,N_4111,N_3993);
or U4360 (N_4360,N_4032,N_4195);
or U4361 (N_4361,N_4091,N_4182);
and U4362 (N_4362,N_3900,N_4153);
nor U4363 (N_4363,N_3915,N_4008);
or U4364 (N_4364,N_3927,N_4136);
and U4365 (N_4365,N_4060,N_3910);
nand U4366 (N_4366,N_3975,N_4094);
nor U4367 (N_4367,N_4056,N_3978);
or U4368 (N_4368,N_4045,N_4017);
and U4369 (N_4369,N_3972,N_4129);
nor U4370 (N_4370,N_4011,N_3986);
or U4371 (N_4371,N_4049,N_4145);
nand U4372 (N_4372,N_4167,N_4154);
and U4373 (N_4373,N_4042,N_4139);
xnor U4374 (N_4374,N_4096,N_4163);
nor U4375 (N_4375,N_4055,N_4142);
or U4376 (N_4376,N_4125,N_4127);
nand U4377 (N_4377,N_3917,N_4157);
nand U4378 (N_4378,N_4032,N_3956);
nand U4379 (N_4379,N_4093,N_4120);
and U4380 (N_4380,N_4092,N_4193);
or U4381 (N_4381,N_4091,N_3995);
or U4382 (N_4382,N_4166,N_3918);
xor U4383 (N_4383,N_3902,N_4026);
nor U4384 (N_4384,N_4037,N_3903);
and U4385 (N_4385,N_3905,N_4039);
nor U4386 (N_4386,N_4055,N_4166);
and U4387 (N_4387,N_4135,N_4169);
and U4388 (N_4388,N_4170,N_3930);
nand U4389 (N_4389,N_3971,N_3966);
nor U4390 (N_4390,N_4113,N_4121);
nor U4391 (N_4391,N_4158,N_3996);
or U4392 (N_4392,N_4131,N_3919);
and U4393 (N_4393,N_3992,N_4053);
xnor U4394 (N_4394,N_4132,N_4161);
nor U4395 (N_4395,N_4057,N_4190);
and U4396 (N_4396,N_4146,N_4095);
nor U4397 (N_4397,N_4014,N_4028);
nand U4398 (N_4398,N_3986,N_4114);
and U4399 (N_4399,N_3908,N_4195);
nand U4400 (N_4400,N_4072,N_3986);
and U4401 (N_4401,N_4198,N_4190);
or U4402 (N_4402,N_4128,N_3918);
and U4403 (N_4403,N_4068,N_4069);
nor U4404 (N_4404,N_4068,N_4046);
and U4405 (N_4405,N_4083,N_4163);
nor U4406 (N_4406,N_3926,N_4149);
or U4407 (N_4407,N_4050,N_3947);
xnor U4408 (N_4408,N_4100,N_3994);
nor U4409 (N_4409,N_4028,N_3911);
nand U4410 (N_4410,N_4187,N_4145);
nand U4411 (N_4411,N_4084,N_4053);
and U4412 (N_4412,N_4192,N_3905);
nor U4413 (N_4413,N_4155,N_4055);
nand U4414 (N_4414,N_4188,N_4037);
and U4415 (N_4415,N_4192,N_4026);
nor U4416 (N_4416,N_3984,N_3952);
xnor U4417 (N_4417,N_4036,N_3900);
nand U4418 (N_4418,N_3983,N_4045);
nor U4419 (N_4419,N_3992,N_4159);
nor U4420 (N_4420,N_4140,N_4002);
nand U4421 (N_4421,N_4085,N_3944);
nor U4422 (N_4422,N_4076,N_4006);
or U4423 (N_4423,N_4160,N_3917);
and U4424 (N_4424,N_4123,N_4109);
nand U4425 (N_4425,N_4193,N_4174);
or U4426 (N_4426,N_4158,N_4140);
nor U4427 (N_4427,N_4047,N_4064);
nor U4428 (N_4428,N_4162,N_4100);
nand U4429 (N_4429,N_3948,N_4059);
xnor U4430 (N_4430,N_3983,N_3994);
xor U4431 (N_4431,N_4111,N_4070);
nand U4432 (N_4432,N_3994,N_4157);
nand U4433 (N_4433,N_4024,N_4111);
xnor U4434 (N_4434,N_3988,N_3902);
or U4435 (N_4435,N_4061,N_4040);
xor U4436 (N_4436,N_3991,N_4158);
xor U4437 (N_4437,N_4011,N_4049);
nor U4438 (N_4438,N_4086,N_4176);
xnor U4439 (N_4439,N_4117,N_4055);
and U4440 (N_4440,N_4189,N_3955);
and U4441 (N_4441,N_3948,N_3925);
or U4442 (N_4442,N_4046,N_4051);
or U4443 (N_4443,N_4028,N_3932);
xnor U4444 (N_4444,N_3941,N_3988);
nand U4445 (N_4445,N_4087,N_4190);
or U4446 (N_4446,N_4028,N_4136);
xnor U4447 (N_4447,N_4010,N_4167);
nand U4448 (N_4448,N_4048,N_4041);
and U4449 (N_4449,N_3980,N_4190);
or U4450 (N_4450,N_4113,N_4079);
and U4451 (N_4451,N_3982,N_3901);
nand U4452 (N_4452,N_4112,N_3929);
xnor U4453 (N_4453,N_3995,N_3945);
and U4454 (N_4454,N_4171,N_3989);
or U4455 (N_4455,N_4053,N_4139);
and U4456 (N_4456,N_3971,N_4138);
or U4457 (N_4457,N_4130,N_3930);
nand U4458 (N_4458,N_3908,N_4183);
nor U4459 (N_4459,N_4137,N_4075);
and U4460 (N_4460,N_4158,N_4020);
or U4461 (N_4461,N_4026,N_3915);
nor U4462 (N_4462,N_4138,N_4072);
and U4463 (N_4463,N_4176,N_4130);
or U4464 (N_4464,N_4101,N_4026);
nand U4465 (N_4465,N_4178,N_3927);
nor U4466 (N_4466,N_4056,N_3945);
nor U4467 (N_4467,N_3994,N_4168);
or U4468 (N_4468,N_3981,N_3917);
and U4469 (N_4469,N_4076,N_4002);
or U4470 (N_4470,N_4149,N_3986);
or U4471 (N_4471,N_4104,N_4122);
nor U4472 (N_4472,N_3990,N_4190);
nor U4473 (N_4473,N_4056,N_4107);
or U4474 (N_4474,N_3951,N_4008);
and U4475 (N_4475,N_4041,N_4167);
nand U4476 (N_4476,N_4117,N_4077);
xor U4477 (N_4477,N_4047,N_4049);
or U4478 (N_4478,N_4049,N_4101);
xor U4479 (N_4479,N_4140,N_3961);
xnor U4480 (N_4480,N_4092,N_3958);
nand U4481 (N_4481,N_4021,N_4030);
or U4482 (N_4482,N_3975,N_3900);
or U4483 (N_4483,N_4192,N_3975);
and U4484 (N_4484,N_3933,N_4077);
nor U4485 (N_4485,N_3939,N_3922);
nor U4486 (N_4486,N_4143,N_3972);
nor U4487 (N_4487,N_4097,N_4138);
or U4488 (N_4488,N_4070,N_4179);
or U4489 (N_4489,N_4058,N_4097);
xor U4490 (N_4490,N_4151,N_4084);
nor U4491 (N_4491,N_3916,N_4147);
nor U4492 (N_4492,N_4071,N_4120);
nor U4493 (N_4493,N_4042,N_4075);
or U4494 (N_4494,N_4190,N_4149);
xnor U4495 (N_4495,N_4188,N_4030);
nor U4496 (N_4496,N_4198,N_4116);
or U4497 (N_4497,N_4135,N_3949);
nor U4498 (N_4498,N_3990,N_3988);
xnor U4499 (N_4499,N_4007,N_3970);
or U4500 (N_4500,N_4370,N_4478);
nor U4501 (N_4501,N_4279,N_4423);
and U4502 (N_4502,N_4448,N_4496);
or U4503 (N_4503,N_4300,N_4245);
nand U4504 (N_4504,N_4379,N_4359);
nand U4505 (N_4505,N_4497,N_4434);
and U4506 (N_4506,N_4320,N_4425);
nand U4507 (N_4507,N_4254,N_4253);
nand U4508 (N_4508,N_4429,N_4399);
or U4509 (N_4509,N_4480,N_4221);
nor U4510 (N_4510,N_4476,N_4266);
or U4511 (N_4511,N_4283,N_4489);
or U4512 (N_4512,N_4347,N_4224);
or U4513 (N_4513,N_4335,N_4269);
or U4514 (N_4514,N_4459,N_4303);
nor U4515 (N_4515,N_4299,N_4210);
or U4516 (N_4516,N_4212,N_4403);
or U4517 (N_4517,N_4220,N_4402);
xnor U4518 (N_4518,N_4318,N_4435);
nor U4519 (N_4519,N_4329,N_4331);
and U4520 (N_4520,N_4377,N_4244);
xnor U4521 (N_4521,N_4345,N_4207);
or U4522 (N_4522,N_4404,N_4414);
nor U4523 (N_4523,N_4427,N_4219);
xnor U4524 (N_4524,N_4289,N_4317);
and U4525 (N_4525,N_4374,N_4201);
nor U4526 (N_4526,N_4360,N_4225);
nor U4527 (N_4527,N_4366,N_4341);
xor U4528 (N_4528,N_4275,N_4388);
xnor U4529 (N_4529,N_4230,N_4250);
and U4530 (N_4530,N_4463,N_4492);
or U4531 (N_4531,N_4306,N_4452);
and U4532 (N_4532,N_4421,N_4413);
xnor U4533 (N_4533,N_4213,N_4292);
or U4534 (N_4534,N_4256,N_4324);
nor U4535 (N_4535,N_4323,N_4419);
xnor U4536 (N_4536,N_4396,N_4348);
nor U4537 (N_4537,N_4386,N_4484);
nor U4538 (N_4538,N_4385,N_4475);
xor U4539 (N_4539,N_4354,N_4298);
nand U4540 (N_4540,N_4200,N_4491);
nand U4541 (N_4541,N_4450,N_4276);
and U4542 (N_4542,N_4390,N_4357);
or U4543 (N_4543,N_4321,N_4342);
nor U4544 (N_4544,N_4235,N_4268);
and U4545 (N_4545,N_4297,N_4285);
xnor U4546 (N_4546,N_4286,N_4454);
nor U4547 (N_4547,N_4352,N_4499);
xor U4548 (N_4548,N_4490,N_4365);
and U4549 (N_4549,N_4486,N_4251);
and U4550 (N_4550,N_4319,N_4401);
or U4551 (N_4551,N_4238,N_4305);
nand U4552 (N_4552,N_4485,N_4458);
or U4553 (N_4553,N_4392,N_4308);
and U4554 (N_4554,N_4255,N_4314);
xor U4555 (N_4555,N_4264,N_4466);
and U4556 (N_4556,N_4481,N_4280);
nand U4557 (N_4557,N_4330,N_4234);
and U4558 (N_4558,N_4407,N_4364);
or U4559 (N_4559,N_4265,N_4227);
and U4560 (N_4560,N_4239,N_4311);
xnor U4561 (N_4561,N_4397,N_4443);
or U4562 (N_4562,N_4209,N_4483);
or U4563 (N_4563,N_4494,N_4441);
and U4564 (N_4564,N_4247,N_4334);
xnor U4565 (N_4565,N_4204,N_4217);
and U4566 (N_4566,N_4249,N_4442);
and U4567 (N_4567,N_4270,N_4465);
nor U4568 (N_4568,N_4322,N_4284);
nand U4569 (N_4569,N_4432,N_4336);
and U4570 (N_4570,N_4428,N_4228);
and U4571 (N_4571,N_4358,N_4461);
xnor U4572 (N_4572,N_4216,N_4240);
xnor U4573 (N_4573,N_4363,N_4468);
or U4574 (N_4574,N_4472,N_4437);
and U4575 (N_4575,N_4393,N_4451);
or U4576 (N_4576,N_4355,N_4222);
and U4577 (N_4577,N_4383,N_4426);
or U4578 (N_4578,N_4373,N_4202);
and U4579 (N_4579,N_4444,N_4367);
nor U4580 (N_4580,N_4293,N_4315);
xor U4581 (N_4581,N_4462,N_4333);
or U4582 (N_4582,N_4498,N_4471);
nor U4583 (N_4583,N_4327,N_4262);
and U4584 (N_4584,N_4416,N_4350);
nand U4585 (N_4585,N_4464,N_4361);
or U4586 (N_4586,N_4487,N_4260);
xnor U4587 (N_4587,N_4446,N_4460);
and U4588 (N_4588,N_4467,N_4353);
nand U4589 (N_4589,N_4325,N_4274);
or U4590 (N_4590,N_4391,N_4438);
nor U4591 (N_4591,N_4436,N_4326);
nand U4592 (N_4592,N_4271,N_4312);
nor U4593 (N_4593,N_4422,N_4440);
nand U4594 (N_4594,N_4316,N_4338);
xnor U4595 (N_4595,N_4420,N_4307);
and U4596 (N_4596,N_4282,N_4433);
xor U4597 (N_4597,N_4208,N_4394);
or U4598 (N_4598,N_4493,N_4304);
nor U4599 (N_4599,N_4295,N_4371);
and U4600 (N_4600,N_4457,N_4237);
nand U4601 (N_4601,N_4231,N_4445);
or U4602 (N_4602,N_4206,N_4349);
xnor U4603 (N_4603,N_4372,N_4455);
and U4604 (N_4604,N_4406,N_4453);
nor U4605 (N_4605,N_4380,N_4281);
and U4606 (N_4606,N_4368,N_4477);
and U4607 (N_4607,N_4469,N_4405);
nor U4608 (N_4608,N_4415,N_4203);
and U4609 (N_4609,N_4339,N_4313);
or U4610 (N_4610,N_4449,N_4278);
nor U4611 (N_4611,N_4439,N_4229);
or U4612 (N_4612,N_4309,N_4273);
nor U4613 (N_4613,N_4205,N_4257);
or U4614 (N_4614,N_4369,N_4447);
nor U4615 (N_4615,N_4470,N_4412);
and U4616 (N_4616,N_4236,N_4259);
nor U4617 (N_4617,N_4346,N_4302);
xnor U4618 (N_4618,N_4288,N_4218);
nand U4619 (N_4619,N_4291,N_4243);
nor U4620 (N_4620,N_4344,N_4242);
xnor U4621 (N_4621,N_4246,N_4328);
nand U4622 (N_4622,N_4351,N_4395);
and U4623 (N_4623,N_4263,N_4332);
or U4624 (N_4624,N_4389,N_4410);
xor U4625 (N_4625,N_4362,N_4474);
or U4626 (N_4626,N_4290,N_4409);
or U4627 (N_4627,N_4248,N_4310);
or U4628 (N_4628,N_4398,N_4378);
and U4629 (N_4629,N_4261,N_4340);
nor U4630 (N_4630,N_4252,N_4267);
and U4631 (N_4631,N_4430,N_4408);
xor U4632 (N_4632,N_4431,N_4223);
nor U4633 (N_4633,N_4232,N_4418);
xor U4634 (N_4634,N_4356,N_4387);
nor U4635 (N_4635,N_4296,N_4473);
nand U4636 (N_4636,N_4214,N_4211);
and U4637 (N_4637,N_4294,N_4233);
nor U4638 (N_4638,N_4375,N_4241);
nor U4639 (N_4639,N_4343,N_4384);
xor U4640 (N_4640,N_4417,N_4226);
nor U4641 (N_4641,N_4479,N_4482);
xor U4642 (N_4642,N_4215,N_4258);
and U4643 (N_4643,N_4277,N_4272);
nor U4644 (N_4644,N_4376,N_4400);
xor U4645 (N_4645,N_4337,N_4287);
xor U4646 (N_4646,N_4456,N_4488);
nor U4647 (N_4647,N_4495,N_4301);
xor U4648 (N_4648,N_4382,N_4411);
nor U4649 (N_4649,N_4381,N_4424);
or U4650 (N_4650,N_4423,N_4257);
or U4651 (N_4651,N_4308,N_4263);
nand U4652 (N_4652,N_4296,N_4334);
xor U4653 (N_4653,N_4307,N_4321);
xnor U4654 (N_4654,N_4236,N_4254);
xor U4655 (N_4655,N_4244,N_4478);
or U4656 (N_4656,N_4328,N_4217);
and U4657 (N_4657,N_4309,N_4418);
nand U4658 (N_4658,N_4477,N_4210);
nor U4659 (N_4659,N_4270,N_4281);
nor U4660 (N_4660,N_4232,N_4213);
and U4661 (N_4661,N_4408,N_4427);
nand U4662 (N_4662,N_4360,N_4208);
nor U4663 (N_4663,N_4376,N_4282);
and U4664 (N_4664,N_4460,N_4350);
and U4665 (N_4665,N_4495,N_4317);
nor U4666 (N_4666,N_4204,N_4395);
or U4667 (N_4667,N_4481,N_4380);
nand U4668 (N_4668,N_4467,N_4492);
nor U4669 (N_4669,N_4383,N_4412);
and U4670 (N_4670,N_4205,N_4297);
and U4671 (N_4671,N_4335,N_4434);
and U4672 (N_4672,N_4243,N_4469);
or U4673 (N_4673,N_4278,N_4203);
nor U4674 (N_4674,N_4424,N_4316);
or U4675 (N_4675,N_4282,N_4273);
nor U4676 (N_4676,N_4382,N_4293);
and U4677 (N_4677,N_4272,N_4450);
xnor U4678 (N_4678,N_4498,N_4408);
xnor U4679 (N_4679,N_4455,N_4284);
xor U4680 (N_4680,N_4388,N_4270);
nand U4681 (N_4681,N_4206,N_4468);
nand U4682 (N_4682,N_4224,N_4226);
or U4683 (N_4683,N_4212,N_4340);
and U4684 (N_4684,N_4301,N_4478);
nand U4685 (N_4685,N_4253,N_4289);
or U4686 (N_4686,N_4218,N_4209);
and U4687 (N_4687,N_4257,N_4463);
or U4688 (N_4688,N_4234,N_4313);
or U4689 (N_4689,N_4334,N_4405);
and U4690 (N_4690,N_4227,N_4406);
or U4691 (N_4691,N_4268,N_4417);
xor U4692 (N_4692,N_4242,N_4443);
and U4693 (N_4693,N_4427,N_4248);
or U4694 (N_4694,N_4476,N_4369);
nand U4695 (N_4695,N_4240,N_4205);
or U4696 (N_4696,N_4353,N_4307);
nand U4697 (N_4697,N_4216,N_4413);
or U4698 (N_4698,N_4395,N_4274);
xnor U4699 (N_4699,N_4355,N_4477);
or U4700 (N_4700,N_4247,N_4440);
or U4701 (N_4701,N_4380,N_4420);
and U4702 (N_4702,N_4203,N_4214);
and U4703 (N_4703,N_4259,N_4495);
or U4704 (N_4704,N_4364,N_4479);
and U4705 (N_4705,N_4472,N_4444);
nor U4706 (N_4706,N_4351,N_4447);
and U4707 (N_4707,N_4297,N_4273);
nor U4708 (N_4708,N_4416,N_4389);
nand U4709 (N_4709,N_4208,N_4439);
or U4710 (N_4710,N_4247,N_4475);
nor U4711 (N_4711,N_4416,N_4281);
nand U4712 (N_4712,N_4364,N_4454);
nand U4713 (N_4713,N_4228,N_4322);
and U4714 (N_4714,N_4421,N_4311);
and U4715 (N_4715,N_4202,N_4334);
nand U4716 (N_4716,N_4331,N_4262);
nor U4717 (N_4717,N_4348,N_4251);
nor U4718 (N_4718,N_4347,N_4489);
and U4719 (N_4719,N_4269,N_4394);
or U4720 (N_4720,N_4275,N_4276);
nor U4721 (N_4721,N_4201,N_4381);
nand U4722 (N_4722,N_4359,N_4202);
or U4723 (N_4723,N_4328,N_4348);
nor U4724 (N_4724,N_4239,N_4476);
nor U4725 (N_4725,N_4225,N_4423);
and U4726 (N_4726,N_4203,N_4460);
nor U4727 (N_4727,N_4294,N_4408);
and U4728 (N_4728,N_4417,N_4412);
xor U4729 (N_4729,N_4325,N_4393);
and U4730 (N_4730,N_4430,N_4457);
and U4731 (N_4731,N_4277,N_4360);
nand U4732 (N_4732,N_4204,N_4259);
nand U4733 (N_4733,N_4463,N_4296);
nand U4734 (N_4734,N_4393,N_4302);
xnor U4735 (N_4735,N_4337,N_4341);
nor U4736 (N_4736,N_4309,N_4490);
xor U4737 (N_4737,N_4208,N_4330);
and U4738 (N_4738,N_4242,N_4239);
xor U4739 (N_4739,N_4389,N_4434);
and U4740 (N_4740,N_4408,N_4366);
nor U4741 (N_4741,N_4389,N_4298);
nand U4742 (N_4742,N_4491,N_4306);
nand U4743 (N_4743,N_4383,N_4333);
nor U4744 (N_4744,N_4433,N_4322);
and U4745 (N_4745,N_4450,N_4264);
nor U4746 (N_4746,N_4480,N_4205);
nand U4747 (N_4747,N_4430,N_4217);
or U4748 (N_4748,N_4255,N_4394);
and U4749 (N_4749,N_4488,N_4219);
nand U4750 (N_4750,N_4419,N_4328);
nor U4751 (N_4751,N_4434,N_4202);
xor U4752 (N_4752,N_4492,N_4477);
nand U4753 (N_4753,N_4408,N_4326);
nand U4754 (N_4754,N_4417,N_4339);
xor U4755 (N_4755,N_4457,N_4462);
and U4756 (N_4756,N_4294,N_4466);
nand U4757 (N_4757,N_4304,N_4470);
and U4758 (N_4758,N_4494,N_4484);
and U4759 (N_4759,N_4396,N_4274);
nand U4760 (N_4760,N_4345,N_4338);
xor U4761 (N_4761,N_4274,N_4403);
xor U4762 (N_4762,N_4320,N_4340);
nor U4763 (N_4763,N_4314,N_4381);
xnor U4764 (N_4764,N_4227,N_4317);
or U4765 (N_4765,N_4347,N_4286);
nor U4766 (N_4766,N_4380,N_4214);
xor U4767 (N_4767,N_4473,N_4294);
nand U4768 (N_4768,N_4217,N_4389);
nor U4769 (N_4769,N_4270,N_4437);
nor U4770 (N_4770,N_4309,N_4414);
nor U4771 (N_4771,N_4375,N_4283);
or U4772 (N_4772,N_4477,N_4321);
xnor U4773 (N_4773,N_4283,N_4210);
and U4774 (N_4774,N_4451,N_4360);
nand U4775 (N_4775,N_4207,N_4386);
or U4776 (N_4776,N_4321,N_4454);
and U4777 (N_4777,N_4244,N_4371);
nand U4778 (N_4778,N_4373,N_4313);
xnor U4779 (N_4779,N_4300,N_4394);
nand U4780 (N_4780,N_4486,N_4488);
xor U4781 (N_4781,N_4214,N_4431);
nor U4782 (N_4782,N_4454,N_4317);
nand U4783 (N_4783,N_4437,N_4330);
or U4784 (N_4784,N_4327,N_4440);
nand U4785 (N_4785,N_4336,N_4280);
and U4786 (N_4786,N_4334,N_4383);
or U4787 (N_4787,N_4313,N_4334);
nor U4788 (N_4788,N_4210,N_4201);
nand U4789 (N_4789,N_4310,N_4422);
xnor U4790 (N_4790,N_4421,N_4450);
xor U4791 (N_4791,N_4209,N_4212);
or U4792 (N_4792,N_4272,N_4211);
nand U4793 (N_4793,N_4359,N_4276);
nand U4794 (N_4794,N_4311,N_4372);
nor U4795 (N_4795,N_4411,N_4392);
xor U4796 (N_4796,N_4267,N_4295);
xnor U4797 (N_4797,N_4404,N_4264);
and U4798 (N_4798,N_4297,N_4339);
or U4799 (N_4799,N_4416,N_4431);
and U4800 (N_4800,N_4711,N_4636);
nand U4801 (N_4801,N_4786,N_4662);
xor U4802 (N_4802,N_4560,N_4655);
nand U4803 (N_4803,N_4550,N_4607);
or U4804 (N_4804,N_4631,N_4597);
nand U4805 (N_4805,N_4630,N_4531);
and U4806 (N_4806,N_4663,N_4744);
or U4807 (N_4807,N_4731,N_4618);
and U4808 (N_4808,N_4626,N_4559);
and U4809 (N_4809,N_4545,N_4608);
nor U4810 (N_4810,N_4503,N_4682);
xor U4811 (N_4811,N_4654,N_4622);
nor U4812 (N_4812,N_4722,N_4688);
and U4813 (N_4813,N_4639,N_4793);
and U4814 (N_4814,N_4653,N_4527);
nand U4815 (N_4815,N_4652,N_4641);
or U4816 (N_4816,N_4667,N_4792);
nor U4817 (N_4817,N_4536,N_4727);
nand U4818 (N_4818,N_4543,N_4554);
xnor U4819 (N_4819,N_4742,N_4574);
and U4820 (N_4820,N_4704,N_4657);
nand U4821 (N_4821,N_4528,N_4557);
nand U4822 (N_4822,N_4569,N_4646);
or U4823 (N_4823,N_4635,N_4587);
nor U4824 (N_4824,N_4678,N_4782);
xnor U4825 (N_4825,N_4714,N_4519);
nand U4826 (N_4826,N_4596,N_4796);
nand U4827 (N_4827,N_4666,N_4748);
or U4828 (N_4828,N_4552,N_4583);
or U4829 (N_4829,N_4617,N_4585);
nor U4830 (N_4830,N_4791,N_4717);
and U4831 (N_4831,N_4763,N_4577);
nor U4832 (N_4832,N_4650,N_4575);
nor U4833 (N_4833,N_4625,N_4677);
and U4834 (N_4834,N_4563,N_4774);
xor U4835 (N_4835,N_4707,N_4627);
and U4836 (N_4836,N_4721,N_4609);
nor U4837 (N_4837,N_4773,N_4522);
xor U4838 (N_4838,N_4532,N_4725);
nand U4839 (N_4839,N_4765,N_4787);
or U4840 (N_4840,N_4570,N_4584);
or U4841 (N_4841,N_4517,N_4753);
and U4842 (N_4842,N_4743,N_4592);
or U4843 (N_4843,N_4740,N_4789);
nor U4844 (N_4844,N_4526,N_4561);
nand U4845 (N_4845,N_4565,N_4612);
nand U4846 (N_4846,N_4757,N_4647);
nor U4847 (N_4847,N_4708,N_4593);
nor U4848 (N_4848,N_4735,N_4761);
xnor U4849 (N_4849,N_4610,N_4656);
xnor U4850 (N_4850,N_4555,N_4785);
or U4851 (N_4851,N_4643,N_4611);
nor U4852 (N_4852,N_4673,N_4568);
nor U4853 (N_4853,N_4718,N_4694);
nand U4854 (N_4854,N_4524,N_4598);
nor U4855 (N_4855,N_4799,N_4695);
or U4856 (N_4856,N_4573,N_4516);
nand U4857 (N_4857,N_4776,N_4648);
or U4858 (N_4858,N_4542,N_4778);
nor U4859 (N_4859,N_4693,N_4540);
nor U4860 (N_4860,N_4798,N_4750);
and U4861 (N_4861,N_4586,N_4779);
and U4862 (N_4862,N_4615,N_4692);
or U4863 (N_4863,N_4589,N_4502);
and U4864 (N_4864,N_4566,N_4614);
nor U4865 (N_4865,N_4747,N_4600);
nor U4866 (N_4866,N_4723,N_4613);
or U4867 (N_4867,N_4665,N_4534);
nor U4868 (N_4868,N_4661,N_4705);
nor U4869 (N_4869,N_4701,N_4697);
and U4870 (N_4870,N_4762,N_4752);
xor U4871 (N_4871,N_4637,N_4576);
nand U4872 (N_4872,N_4685,N_4706);
or U4873 (N_4873,N_4755,N_4681);
nor U4874 (N_4874,N_4518,N_4741);
nand U4875 (N_4875,N_4670,N_4700);
nor U4876 (N_4876,N_4501,N_4766);
and U4877 (N_4877,N_4749,N_4726);
nor U4878 (N_4878,N_4515,N_4724);
xor U4879 (N_4879,N_4764,N_4633);
nor U4880 (N_4880,N_4572,N_4732);
nand U4881 (N_4881,N_4745,N_4671);
nor U4882 (N_4882,N_4702,N_4571);
nor U4883 (N_4883,N_4538,N_4523);
xnor U4884 (N_4884,N_4760,N_4664);
xnor U4885 (N_4885,N_4530,N_4709);
nand U4886 (N_4886,N_4780,N_4621);
nand U4887 (N_4887,N_4508,N_4590);
nor U4888 (N_4888,N_4553,N_4734);
nand U4889 (N_4889,N_4513,N_4698);
nand U4890 (N_4890,N_4603,N_4767);
xnor U4891 (N_4891,N_4544,N_4602);
nand U4892 (N_4892,N_4730,N_4795);
and U4893 (N_4893,N_4712,N_4736);
or U4894 (N_4894,N_4507,N_4537);
nor U4895 (N_4895,N_4772,N_4506);
or U4896 (N_4896,N_4746,N_4649);
nor U4897 (N_4897,N_4771,N_4505);
or U4898 (N_4898,N_4719,N_4684);
nand U4899 (N_4899,N_4541,N_4710);
or U4900 (N_4900,N_4616,N_4728);
nor U4901 (N_4901,N_4558,N_4642);
and U4902 (N_4902,N_4713,N_4686);
xor U4903 (N_4903,N_4674,N_4659);
nor U4904 (N_4904,N_4556,N_4605);
or U4905 (N_4905,N_4514,N_4788);
nand U4906 (N_4906,N_4546,N_4567);
and U4907 (N_4907,N_4521,N_4783);
nand U4908 (N_4908,N_4738,N_4510);
nand U4909 (N_4909,N_4683,N_4720);
nand U4910 (N_4910,N_4638,N_4751);
and U4911 (N_4911,N_4511,N_4781);
or U4912 (N_4912,N_4651,N_4672);
xor U4913 (N_4913,N_4580,N_4624);
xnor U4914 (N_4914,N_4769,N_4595);
and U4915 (N_4915,N_4690,N_4581);
nand U4916 (N_4916,N_4628,N_4620);
nand U4917 (N_4917,N_4759,N_4691);
xor U4918 (N_4918,N_4591,N_4588);
nand U4919 (N_4919,N_4629,N_4551);
nor U4920 (N_4920,N_4645,N_4582);
nor U4921 (N_4921,N_4784,N_4512);
xnor U4922 (N_4922,N_4562,N_4634);
nand U4923 (N_4923,N_4716,N_4794);
and U4924 (N_4924,N_4715,N_4500);
nor U4925 (N_4925,N_4601,N_4777);
nand U4926 (N_4926,N_4739,N_4564);
nand U4927 (N_4927,N_4604,N_4790);
and U4928 (N_4928,N_4775,N_4549);
nand U4929 (N_4929,N_4539,N_4623);
or U4930 (N_4930,N_4504,N_4689);
nand U4931 (N_4931,N_4533,N_4525);
nor U4932 (N_4932,N_4680,N_4548);
nand U4933 (N_4933,N_4547,N_4644);
or U4934 (N_4934,N_4768,N_4579);
and U4935 (N_4935,N_4640,N_4754);
and U4936 (N_4936,N_4599,N_4797);
nand U4937 (N_4937,N_4668,N_4660);
or U4938 (N_4938,N_4529,N_4679);
and U4939 (N_4939,N_4737,N_4770);
nor U4940 (N_4940,N_4675,N_4729);
xnor U4941 (N_4941,N_4687,N_4520);
nand U4942 (N_4942,N_4756,N_4606);
nand U4943 (N_4943,N_4699,N_4733);
nand U4944 (N_4944,N_4703,N_4696);
nor U4945 (N_4945,N_4578,N_4658);
nor U4946 (N_4946,N_4619,N_4669);
or U4947 (N_4947,N_4535,N_4676);
xnor U4948 (N_4948,N_4594,N_4509);
nand U4949 (N_4949,N_4632,N_4758);
and U4950 (N_4950,N_4517,N_4598);
nor U4951 (N_4951,N_4657,N_4503);
nor U4952 (N_4952,N_4585,N_4798);
or U4953 (N_4953,N_4765,N_4577);
and U4954 (N_4954,N_4706,N_4750);
xor U4955 (N_4955,N_4683,N_4714);
xnor U4956 (N_4956,N_4689,N_4714);
xnor U4957 (N_4957,N_4793,N_4561);
or U4958 (N_4958,N_4683,N_4577);
or U4959 (N_4959,N_4611,N_4539);
or U4960 (N_4960,N_4783,N_4519);
xor U4961 (N_4961,N_4647,N_4790);
nor U4962 (N_4962,N_4500,N_4716);
nand U4963 (N_4963,N_4653,N_4543);
nor U4964 (N_4964,N_4718,N_4623);
nor U4965 (N_4965,N_4735,N_4683);
nand U4966 (N_4966,N_4630,N_4725);
or U4967 (N_4967,N_4640,N_4791);
and U4968 (N_4968,N_4530,N_4591);
or U4969 (N_4969,N_4601,N_4774);
nand U4970 (N_4970,N_4553,N_4670);
xor U4971 (N_4971,N_4505,N_4656);
nand U4972 (N_4972,N_4774,N_4678);
xnor U4973 (N_4973,N_4668,N_4571);
nand U4974 (N_4974,N_4556,N_4693);
nand U4975 (N_4975,N_4652,N_4670);
or U4976 (N_4976,N_4549,N_4757);
xor U4977 (N_4977,N_4751,N_4781);
nand U4978 (N_4978,N_4632,N_4607);
nor U4979 (N_4979,N_4779,N_4581);
nor U4980 (N_4980,N_4595,N_4642);
nand U4981 (N_4981,N_4790,N_4613);
nand U4982 (N_4982,N_4753,N_4633);
nor U4983 (N_4983,N_4508,N_4519);
and U4984 (N_4984,N_4641,N_4619);
and U4985 (N_4985,N_4578,N_4600);
nor U4986 (N_4986,N_4658,N_4612);
nand U4987 (N_4987,N_4679,N_4686);
xnor U4988 (N_4988,N_4541,N_4622);
or U4989 (N_4989,N_4539,N_4557);
xor U4990 (N_4990,N_4597,N_4608);
nand U4991 (N_4991,N_4784,N_4518);
nor U4992 (N_4992,N_4567,N_4591);
nand U4993 (N_4993,N_4534,N_4619);
or U4994 (N_4994,N_4753,N_4528);
nand U4995 (N_4995,N_4703,N_4727);
and U4996 (N_4996,N_4631,N_4642);
nand U4997 (N_4997,N_4735,N_4540);
nand U4998 (N_4998,N_4760,N_4570);
or U4999 (N_4999,N_4731,N_4747);
nand U5000 (N_5000,N_4651,N_4677);
nand U5001 (N_5001,N_4541,N_4752);
nor U5002 (N_5002,N_4600,N_4530);
nand U5003 (N_5003,N_4680,N_4638);
nand U5004 (N_5004,N_4545,N_4750);
and U5005 (N_5005,N_4567,N_4790);
nor U5006 (N_5006,N_4761,N_4698);
nand U5007 (N_5007,N_4607,N_4662);
and U5008 (N_5008,N_4790,N_4562);
and U5009 (N_5009,N_4533,N_4666);
or U5010 (N_5010,N_4646,N_4653);
and U5011 (N_5011,N_4665,N_4755);
or U5012 (N_5012,N_4670,N_4671);
or U5013 (N_5013,N_4531,N_4598);
xor U5014 (N_5014,N_4523,N_4792);
nand U5015 (N_5015,N_4517,N_4626);
nor U5016 (N_5016,N_4710,N_4577);
nand U5017 (N_5017,N_4723,N_4587);
nor U5018 (N_5018,N_4752,N_4512);
nand U5019 (N_5019,N_4529,N_4671);
xor U5020 (N_5020,N_4577,N_4725);
nand U5021 (N_5021,N_4697,N_4773);
and U5022 (N_5022,N_4559,N_4545);
xor U5023 (N_5023,N_4768,N_4646);
or U5024 (N_5024,N_4570,N_4550);
xnor U5025 (N_5025,N_4644,N_4554);
and U5026 (N_5026,N_4567,N_4778);
xor U5027 (N_5027,N_4606,N_4724);
and U5028 (N_5028,N_4690,N_4582);
nor U5029 (N_5029,N_4584,N_4666);
or U5030 (N_5030,N_4767,N_4634);
nor U5031 (N_5031,N_4538,N_4577);
and U5032 (N_5032,N_4762,N_4707);
nand U5033 (N_5033,N_4713,N_4797);
xor U5034 (N_5034,N_4630,N_4720);
nor U5035 (N_5035,N_4541,N_4774);
or U5036 (N_5036,N_4525,N_4734);
nand U5037 (N_5037,N_4770,N_4634);
and U5038 (N_5038,N_4644,N_4608);
and U5039 (N_5039,N_4585,N_4580);
nand U5040 (N_5040,N_4690,N_4547);
and U5041 (N_5041,N_4676,N_4622);
nand U5042 (N_5042,N_4654,N_4787);
nand U5043 (N_5043,N_4760,N_4517);
nor U5044 (N_5044,N_4545,N_4760);
and U5045 (N_5045,N_4784,N_4545);
and U5046 (N_5046,N_4630,N_4609);
nand U5047 (N_5047,N_4510,N_4785);
xor U5048 (N_5048,N_4643,N_4631);
and U5049 (N_5049,N_4548,N_4513);
and U5050 (N_5050,N_4730,N_4653);
nand U5051 (N_5051,N_4785,N_4558);
nor U5052 (N_5052,N_4542,N_4652);
nand U5053 (N_5053,N_4704,N_4769);
and U5054 (N_5054,N_4581,N_4589);
and U5055 (N_5055,N_4721,N_4507);
xor U5056 (N_5056,N_4711,N_4716);
or U5057 (N_5057,N_4655,N_4645);
nor U5058 (N_5058,N_4755,N_4692);
or U5059 (N_5059,N_4565,N_4658);
xor U5060 (N_5060,N_4681,N_4536);
nand U5061 (N_5061,N_4788,N_4606);
or U5062 (N_5062,N_4742,N_4630);
nor U5063 (N_5063,N_4641,N_4500);
and U5064 (N_5064,N_4755,N_4683);
nand U5065 (N_5065,N_4760,N_4709);
nand U5066 (N_5066,N_4603,N_4571);
nand U5067 (N_5067,N_4598,N_4652);
or U5068 (N_5068,N_4676,N_4708);
nand U5069 (N_5069,N_4642,N_4609);
xor U5070 (N_5070,N_4749,N_4676);
nand U5071 (N_5071,N_4676,N_4743);
or U5072 (N_5072,N_4728,N_4617);
nand U5073 (N_5073,N_4593,N_4552);
nor U5074 (N_5074,N_4741,N_4566);
or U5075 (N_5075,N_4619,N_4584);
and U5076 (N_5076,N_4765,N_4629);
nand U5077 (N_5077,N_4574,N_4528);
and U5078 (N_5078,N_4723,N_4583);
and U5079 (N_5079,N_4590,N_4505);
xor U5080 (N_5080,N_4612,N_4525);
or U5081 (N_5081,N_4626,N_4551);
nor U5082 (N_5082,N_4561,N_4773);
and U5083 (N_5083,N_4706,N_4770);
nand U5084 (N_5084,N_4592,N_4656);
or U5085 (N_5085,N_4687,N_4654);
and U5086 (N_5086,N_4635,N_4515);
nand U5087 (N_5087,N_4552,N_4647);
nor U5088 (N_5088,N_4710,N_4513);
nor U5089 (N_5089,N_4766,N_4790);
or U5090 (N_5090,N_4681,N_4606);
and U5091 (N_5091,N_4675,N_4771);
and U5092 (N_5092,N_4592,N_4757);
nor U5093 (N_5093,N_4554,N_4506);
or U5094 (N_5094,N_4554,N_4660);
and U5095 (N_5095,N_4629,N_4613);
nand U5096 (N_5096,N_4733,N_4618);
nor U5097 (N_5097,N_4657,N_4646);
nor U5098 (N_5098,N_4712,N_4658);
nand U5099 (N_5099,N_4717,N_4605);
nand U5100 (N_5100,N_4816,N_5074);
nor U5101 (N_5101,N_5015,N_5070);
xor U5102 (N_5102,N_4944,N_4863);
xor U5103 (N_5103,N_5029,N_4838);
and U5104 (N_5104,N_4836,N_4986);
nand U5105 (N_5105,N_4834,N_4820);
or U5106 (N_5106,N_4806,N_4801);
and U5107 (N_5107,N_5087,N_4891);
nand U5108 (N_5108,N_4884,N_4919);
and U5109 (N_5109,N_4954,N_5068);
xor U5110 (N_5110,N_4952,N_4930);
xnor U5111 (N_5111,N_4821,N_4865);
nand U5112 (N_5112,N_4953,N_5004);
nand U5113 (N_5113,N_4909,N_5088);
xnor U5114 (N_5114,N_5064,N_5007);
or U5115 (N_5115,N_5017,N_4847);
nand U5116 (N_5116,N_4921,N_4845);
or U5117 (N_5117,N_4914,N_5002);
or U5118 (N_5118,N_4990,N_5075);
xnor U5119 (N_5119,N_4984,N_5080);
and U5120 (N_5120,N_4974,N_4866);
and U5121 (N_5121,N_4880,N_5052);
and U5122 (N_5122,N_4886,N_5025);
or U5123 (N_5123,N_4889,N_5092);
and U5124 (N_5124,N_4902,N_4818);
or U5125 (N_5125,N_4811,N_4911);
nand U5126 (N_5126,N_4965,N_4927);
or U5127 (N_5127,N_4808,N_4802);
nand U5128 (N_5128,N_4904,N_4991);
or U5129 (N_5129,N_4841,N_5035);
or U5130 (N_5130,N_5060,N_5038);
nor U5131 (N_5131,N_4971,N_5079);
nand U5132 (N_5132,N_4924,N_4829);
or U5133 (N_5133,N_4917,N_4885);
nand U5134 (N_5134,N_4853,N_4882);
xor U5135 (N_5135,N_5051,N_5076);
nor U5136 (N_5136,N_4926,N_4903);
or U5137 (N_5137,N_4852,N_5026);
nor U5138 (N_5138,N_5021,N_5050);
xnor U5139 (N_5139,N_4942,N_4810);
nor U5140 (N_5140,N_4878,N_4812);
xnor U5141 (N_5141,N_4955,N_4868);
or U5142 (N_5142,N_5043,N_4985);
nor U5143 (N_5143,N_4839,N_4981);
nor U5144 (N_5144,N_4950,N_4840);
nand U5145 (N_5145,N_4996,N_4947);
or U5146 (N_5146,N_5063,N_5001);
or U5147 (N_5147,N_5047,N_4893);
xnor U5148 (N_5148,N_4905,N_4867);
and U5149 (N_5149,N_4949,N_4823);
and U5150 (N_5150,N_5083,N_4896);
nor U5151 (N_5151,N_4993,N_4923);
or U5152 (N_5152,N_4945,N_5023);
xnor U5153 (N_5153,N_4895,N_4931);
xnor U5154 (N_5154,N_4804,N_5081);
xnor U5155 (N_5155,N_4872,N_4928);
and U5156 (N_5156,N_4883,N_4830);
xor U5157 (N_5157,N_4910,N_4846);
or U5158 (N_5158,N_5031,N_4957);
or U5159 (N_5159,N_4828,N_4961);
xnor U5160 (N_5160,N_5020,N_5024);
and U5161 (N_5161,N_5089,N_4862);
nor U5162 (N_5162,N_4900,N_4912);
or U5163 (N_5163,N_5053,N_4887);
or U5164 (N_5164,N_4915,N_4843);
nand U5165 (N_5165,N_4807,N_4875);
and U5166 (N_5166,N_4835,N_4998);
xnor U5167 (N_5167,N_5078,N_5040);
or U5168 (N_5168,N_4892,N_5030);
and U5169 (N_5169,N_4994,N_4855);
nand U5170 (N_5170,N_5032,N_5094);
or U5171 (N_5171,N_4825,N_4813);
and U5172 (N_5172,N_4881,N_4934);
and U5173 (N_5173,N_4857,N_4951);
or U5174 (N_5174,N_5012,N_4879);
nand U5175 (N_5175,N_5058,N_4869);
or U5176 (N_5176,N_5013,N_4890);
xor U5177 (N_5177,N_4918,N_5018);
xnor U5178 (N_5178,N_5085,N_5049);
nand U5179 (N_5179,N_5069,N_4908);
and U5180 (N_5180,N_4817,N_4939);
or U5181 (N_5181,N_4963,N_4913);
nand U5182 (N_5182,N_4854,N_4929);
nor U5183 (N_5183,N_4848,N_4975);
nand U5184 (N_5184,N_4859,N_4803);
nand U5185 (N_5185,N_4874,N_5041);
nand U5186 (N_5186,N_5044,N_4831);
nand U5187 (N_5187,N_5071,N_5000);
xnor U5188 (N_5188,N_4966,N_4959);
nand U5189 (N_5189,N_4860,N_4956);
nand U5190 (N_5190,N_4844,N_4907);
xnor U5191 (N_5191,N_5096,N_4962);
or U5192 (N_5192,N_4983,N_4943);
and U5193 (N_5193,N_4969,N_4851);
nand U5194 (N_5194,N_4978,N_5036);
and U5195 (N_5195,N_5066,N_4960);
and U5196 (N_5196,N_4970,N_5093);
xor U5197 (N_5197,N_5065,N_4877);
nor U5198 (N_5198,N_5034,N_4809);
nand U5199 (N_5199,N_4894,N_4898);
or U5200 (N_5200,N_4979,N_5045);
nor U5201 (N_5201,N_4973,N_5082);
xnor U5202 (N_5202,N_5062,N_4856);
nand U5203 (N_5203,N_5097,N_5055);
nor U5204 (N_5204,N_4873,N_4870);
xnor U5205 (N_5205,N_4925,N_4995);
xor U5206 (N_5206,N_4864,N_4964);
xnor U5207 (N_5207,N_4826,N_4837);
or U5208 (N_5208,N_5090,N_5054);
or U5209 (N_5209,N_4832,N_4968);
or U5210 (N_5210,N_4850,N_5056);
xor U5211 (N_5211,N_4937,N_4819);
and U5212 (N_5212,N_4920,N_4980);
nor U5213 (N_5213,N_5067,N_4815);
and U5214 (N_5214,N_5016,N_5091);
xor U5215 (N_5215,N_5014,N_4824);
nor U5216 (N_5216,N_5022,N_4982);
nor U5217 (N_5217,N_5061,N_5077);
xnor U5218 (N_5218,N_4992,N_4805);
nand U5219 (N_5219,N_4946,N_5008);
nand U5220 (N_5220,N_4999,N_4997);
or U5221 (N_5221,N_4987,N_5027);
and U5222 (N_5222,N_4871,N_4842);
nand U5223 (N_5223,N_4833,N_4899);
nand U5224 (N_5224,N_5005,N_4876);
nand U5225 (N_5225,N_5042,N_5072);
xor U5226 (N_5226,N_4897,N_4861);
nor U5227 (N_5227,N_4932,N_5048);
nor U5228 (N_5228,N_5086,N_5099);
xor U5229 (N_5229,N_4958,N_4938);
and U5230 (N_5230,N_5003,N_4977);
nand U5231 (N_5231,N_5073,N_5039);
and U5232 (N_5232,N_4933,N_4972);
or U5233 (N_5233,N_5059,N_4822);
and U5234 (N_5234,N_4935,N_4906);
and U5235 (N_5235,N_4941,N_5037);
nand U5236 (N_5236,N_5019,N_4976);
xnor U5237 (N_5237,N_5046,N_5057);
nor U5238 (N_5238,N_5095,N_5084);
and U5239 (N_5239,N_4948,N_4988);
or U5240 (N_5240,N_5006,N_5011);
nor U5241 (N_5241,N_4967,N_5098);
nor U5242 (N_5242,N_4901,N_4849);
or U5243 (N_5243,N_5028,N_4922);
nor U5244 (N_5244,N_4800,N_4989);
and U5245 (N_5245,N_4814,N_5010);
or U5246 (N_5246,N_4827,N_4936);
and U5247 (N_5247,N_4888,N_5009);
xnor U5248 (N_5248,N_4916,N_5033);
and U5249 (N_5249,N_4858,N_4940);
xor U5250 (N_5250,N_4806,N_4963);
and U5251 (N_5251,N_4951,N_4928);
nor U5252 (N_5252,N_5056,N_5006);
xor U5253 (N_5253,N_4847,N_5059);
nor U5254 (N_5254,N_4839,N_5009);
xor U5255 (N_5255,N_4956,N_5005);
nor U5256 (N_5256,N_5075,N_4984);
and U5257 (N_5257,N_5039,N_4917);
and U5258 (N_5258,N_4871,N_5087);
or U5259 (N_5259,N_4836,N_5025);
and U5260 (N_5260,N_4973,N_5063);
xor U5261 (N_5261,N_5071,N_4845);
nor U5262 (N_5262,N_4827,N_4913);
and U5263 (N_5263,N_5098,N_4932);
and U5264 (N_5264,N_5061,N_4992);
xor U5265 (N_5265,N_4803,N_5031);
nand U5266 (N_5266,N_5005,N_5075);
xnor U5267 (N_5267,N_4970,N_4808);
xor U5268 (N_5268,N_4973,N_5017);
xnor U5269 (N_5269,N_4950,N_5000);
and U5270 (N_5270,N_5044,N_4824);
nand U5271 (N_5271,N_4805,N_4936);
nor U5272 (N_5272,N_4881,N_4906);
nor U5273 (N_5273,N_4873,N_4898);
or U5274 (N_5274,N_4879,N_4912);
and U5275 (N_5275,N_5024,N_4974);
nand U5276 (N_5276,N_4887,N_4954);
nor U5277 (N_5277,N_4940,N_5025);
nor U5278 (N_5278,N_4837,N_5042);
nor U5279 (N_5279,N_4938,N_4808);
nor U5280 (N_5280,N_5062,N_5020);
xnor U5281 (N_5281,N_4916,N_4969);
nor U5282 (N_5282,N_4910,N_5097);
xnor U5283 (N_5283,N_4854,N_4924);
xor U5284 (N_5284,N_4992,N_5085);
nand U5285 (N_5285,N_4868,N_5093);
and U5286 (N_5286,N_4980,N_4963);
nand U5287 (N_5287,N_5091,N_5045);
and U5288 (N_5288,N_5040,N_5071);
and U5289 (N_5289,N_4983,N_4954);
nor U5290 (N_5290,N_4929,N_4920);
nor U5291 (N_5291,N_4990,N_4800);
xor U5292 (N_5292,N_5009,N_4987);
nor U5293 (N_5293,N_5019,N_5008);
xnor U5294 (N_5294,N_5077,N_4978);
nor U5295 (N_5295,N_4960,N_5094);
xnor U5296 (N_5296,N_4842,N_4881);
xnor U5297 (N_5297,N_4958,N_4867);
nand U5298 (N_5298,N_4883,N_4995);
or U5299 (N_5299,N_4993,N_4922);
nand U5300 (N_5300,N_4826,N_4875);
xnor U5301 (N_5301,N_5002,N_4827);
or U5302 (N_5302,N_4897,N_4913);
or U5303 (N_5303,N_4886,N_5090);
or U5304 (N_5304,N_4867,N_4896);
and U5305 (N_5305,N_4857,N_5019);
nor U5306 (N_5306,N_5001,N_4813);
xnor U5307 (N_5307,N_4832,N_4838);
or U5308 (N_5308,N_4973,N_5075);
nand U5309 (N_5309,N_5042,N_5064);
nand U5310 (N_5310,N_4884,N_4853);
nor U5311 (N_5311,N_4927,N_4892);
nand U5312 (N_5312,N_5077,N_5076);
or U5313 (N_5313,N_4993,N_4943);
or U5314 (N_5314,N_4890,N_5042);
nor U5315 (N_5315,N_4907,N_5031);
nand U5316 (N_5316,N_4937,N_4996);
or U5317 (N_5317,N_5023,N_4886);
nand U5318 (N_5318,N_4914,N_5024);
nor U5319 (N_5319,N_4969,N_4879);
and U5320 (N_5320,N_4807,N_4942);
nand U5321 (N_5321,N_4905,N_4872);
or U5322 (N_5322,N_5029,N_4829);
nor U5323 (N_5323,N_4853,N_4891);
nand U5324 (N_5324,N_4964,N_4832);
nor U5325 (N_5325,N_4907,N_5052);
xor U5326 (N_5326,N_4882,N_4822);
xor U5327 (N_5327,N_5009,N_4805);
nor U5328 (N_5328,N_5018,N_4815);
nand U5329 (N_5329,N_4982,N_5039);
nand U5330 (N_5330,N_4935,N_4897);
nand U5331 (N_5331,N_5052,N_5084);
or U5332 (N_5332,N_4903,N_5059);
nor U5333 (N_5333,N_5082,N_4856);
and U5334 (N_5334,N_4839,N_4848);
nor U5335 (N_5335,N_5045,N_5011);
and U5336 (N_5336,N_4924,N_5043);
or U5337 (N_5337,N_4940,N_4816);
nor U5338 (N_5338,N_5058,N_5090);
and U5339 (N_5339,N_5099,N_4843);
nor U5340 (N_5340,N_4889,N_4913);
xor U5341 (N_5341,N_4888,N_4818);
xnor U5342 (N_5342,N_4906,N_5004);
xor U5343 (N_5343,N_4944,N_5058);
and U5344 (N_5344,N_4972,N_4913);
or U5345 (N_5345,N_4886,N_4809);
or U5346 (N_5346,N_4820,N_5067);
nor U5347 (N_5347,N_5071,N_4855);
and U5348 (N_5348,N_4820,N_5023);
xor U5349 (N_5349,N_4891,N_4821);
and U5350 (N_5350,N_4877,N_4859);
or U5351 (N_5351,N_4892,N_4822);
and U5352 (N_5352,N_4943,N_4801);
or U5353 (N_5353,N_4882,N_4987);
nand U5354 (N_5354,N_5000,N_4938);
and U5355 (N_5355,N_5076,N_4983);
xnor U5356 (N_5356,N_4886,N_5095);
xor U5357 (N_5357,N_4889,N_4860);
and U5358 (N_5358,N_4845,N_5088);
or U5359 (N_5359,N_5085,N_4933);
nor U5360 (N_5360,N_4905,N_4961);
and U5361 (N_5361,N_4985,N_5033);
nor U5362 (N_5362,N_4837,N_4975);
or U5363 (N_5363,N_5093,N_4888);
nor U5364 (N_5364,N_4932,N_4872);
nor U5365 (N_5365,N_5049,N_5020);
xor U5366 (N_5366,N_5013,N_4945);
nor U5367 (N_5367,N_4974,N_4868);
nor U5368 (N_5368,N_4947,N_5041);
nor U5369 (N_5369,N_5053,N_5082);
and U5370 (N_5370,N_5099,N_4897);
and U5371 (N_5371,N_5021,N_4941);
nand U5372 (N_5372,N_4815,N_4812);
nand U5373 (N_5373,N_4832,N_4860);
nor U5374 (N_5374,N_5005,N_4858);
xnor U5375 (N_5375,N_4990,N_4874);
nor U5376 (N_5376,N_4971,N_5091);
and U5377 (N_5377,N_5097,N_4988);
xor U5378 (N_5378,N_4965,N_5048);
nor U5379 (N_5379,N_4964,N_4908);
and U5380 (N_5380,N_4940,N_5033);
and U5381 (N_5381,N_4811,N_5061);
and U5382 (N_5382,N_5041,N_4851);
and U5383 (N_5383,N_4805,N_4850);
xor U5384 (N_5384,N_4853,N_5097);
nor U5385 (N_5385,N_4879,N_4818);
nor U5386 (N_5386,N_5053,N_5005);
nand U5387 (N_5387,N_5028,N_4824);
xnor U5388 (N_5388,N_4862,N_4913);
nor U5389 (N_5389,N_4878,N_4936);
or U5390 (N_5390,N_5042,N_5023);
nand U5391 (N_5391,N_4862,N_4966);
and U5392 (N_5392,N_4840,N_4866);
xnor U5393 (N_5393,N_4838,N_5065);
xnor U5394 (N_5394,N_5095,N_4854);
xor U5395 (N_5395,N_5060,N_4997);
and U5396 (N_5396,N_4837,N_5061);
nand U5397 (N_5397,N_5040,N_5083);
and U5398 (N_5398,N_5041,N_4808);
xnor U5399 (N_5399,N_4985,N_4901);
xor U5400 (N_5400,N_5312,N_5129);
or U5401 (N_5401,N_5158,N_5236);
and U5402 (N_5402,N_5109,N_5152);
xor U5403 (N_5403,N_5208,N_5139);
nand U5404 (N_5404,N_5348,N_5136);
or U5405 (N_5405,N_5321,N_5227);
nor U5406 (N_5406,N_5183,N_5249);
and U5407 (N_5407,N_5345,N_5188);
nand U5408 (N_5408,N_5194,N_5241);
nor U5409 (N_5409,N_5195,N_5127);
nand U5410 (N_5410,N_5354,N_5113);
or U5411 (N_5411,N_5147,N_5137);
nor U5412 (N_5412,N_5198,N_5215);
and U5413 (N_5413,N_5211,N_5336);
and U5414 (N_5414,N_5165,N_5294);
nor U5415 (N_5415,N_5234,N_5190);
nand U5416 (N_5416,N_5269,N_5161);
xnor U5417 (N_5417,N_5355,N_5128);
xnor U5418 (N_5418,N_5191,N_5143);
nand U5419 (N_5419,N_5180,N_5101);
nor U5420 (N_5420,N_5105,N_5142);
and U5421 (N_5421,N_5289,N_5248);
nor U5422 (N_5422,N_5299,N_5373);
nand U5423 (N_5423,N_5134,N_5357);
xnor U5424 (N_5424,N_5376,N_5398);
xor U5425 (N_5425,N_5393,N_5245);
or U5426 (N_5426,N_5392,N_5209);
and U5427 (N_5427,N_5155,N_5196);
nor U5428 (N_5428,N_5146,N_5169);
nand U5429 (N_5429,N_5253,N_5154);
nor U5430 (N_5430,N_5316,N_5347);
nor U5431 (N_5431,N_5233,N_5261);
nor U5432 (N_5432,N_5157,N_5112);
and U5433 (N_5433,N_5213,N_5349);
nand U5434 (N_5434,N_5259,N_5362);
xor U5435 (N_5435,N_5186,N_5121);
nor U5436 (N_5436,N_5118,N_5371);
and U5437 (N_5437,N_5212,N_5315);
or U5438 (N_5438,N_5330,N_5167);
nand U5439 (N_5439,N_5162,N_5337);
nand U5440 (N_5440,N_5384,N_5228);
or U5441 (N_5441,N_5344,N_5148);
xnor U5442 (N_5442,N_5232,N_5184);
or U5443 (N_5443,N_5331,N_5322);
xor U5444 (N_5444,N_5358,N_5138);
xor U5445 (N_5445,N_5107,N_5181);
xor U5446 (N_5446,N_5296,N_5395);
or U5447 (N_5447,N_5356,N_5334);
xor U5448 (N_5448,N_5319,N_5173);
and U5449 (N_5449,N_5262,N_5230);
nand U5450 (N_5450,N_5237,N_5323);
and U5451 (N_5451,N_5303,N_5126);
nand U5452 (N_5452,N_5368,N_5290);
or U5453 (N_5453,N_5279,N_5166);
and U5454 (N_5454,N_5175,N_5171);
nand U5455 (N_5455,N_5199,N_5329);
nand U5456 (N_5456,N_5313,N_5268);
nor U5457 (N_5457,N_5131,N_5282);
nand U5458 (N_5458,N_5178,N_5133);
nor U5459 (N_5459,N_5267,N_5244);
xnor U5460 (N_5460,N_5201,N_5111);
xor U5461 (N_5461,N_5350,N_5122);
nand U5462 (N_5462,N_5177,N_5285);
nand U5463 (N_5463,N_5260,N_5189);
or U5464 (N_5464,N_5272,N_5295);
nand U5465 (N_5465,N_5204,N_5256);
and U5466 (N_5466,N_5264,N_5219);
nor U5467 (N_5467,N_5207,N_5339);
xor U5468 (N_5468,N_5104,N_5359);
nor U5469 (N_5469,N_5399,N_5251);
nand U5470 (N_5470,N_5242,N_5153);
and U5471 (N_5471,N_5305,N_5385);
xor U5472 (N_5472,N_5317,N_5270);
or U5473 (N_5473,N_5388,N_5389);
nand U5474 (N_5474,N_5281,N_5324);
nand U5475 (N_5475,N_5218,N_5221);
or U5476 (N_5476,N_5130,N_5116);
nand U5477 (N_5477,N_5397,N_5110);
or U5478 (N_5478,N_5366,N_5263);
nor U5479 (N_5479,N_5308,N_5123);
nor U5480 (N_5480,N_5182,N_5370);
xnor U5481 (N_5481,N_5170,N_5226);
nand U5482 (N_5482,N_5159,N_5205);
xnor U5483 (N_5483,N_5246,N_5378);
nand U5484 (N_5484,N_5302,N_5274);
nor U5485 (N_5485,N_5247,N_5287);
xnor U5486 (N_5486,N_5108,N_5225);
nor U5487 (N_5487,N_5379,N_5117);
nor U5488 (N_5488,N_5377,N_5163);
and U5489 (N_5489,N_5187,N_5149);
or U5490 (N_5490,N_5333,N_5367);
nand U5491 (N_5491,N_5318,N_5346);
xnor U5492 (N_5492,N_5174,N_5306);
and U5493 (N_5493,N_5200,N_5325);
nor U5494 (N_5494,N_5192,N_5327);
and U5495 (N_5495,N_5100,N_5206);
xor U5496 (N_5496,N_5220,N_5203);
nand U5497 (N_5497,N_5120,N_5286);
nand U5498 (N_5498,N_5114,N_5375);
or U5499 (N_5499,N_5254,N_5164);
nand U5500 (N_5500,N_5224,N_5374);
xor U5501 (N_5501,N_5342,N_5360);
nand U5502 (N_5502,N_5222,N_5176);
or U5503 (N_5503,N_5301,N_5396);
nand U5504 (N_5504,N_5298,N_5103);
nand U5505 (N_5505,N_5140,N_5202);
xnor U5506 (N_5506,N_5390,N_5156);
nand U5507 (N_5507,N_5193,N_5258);
xnor U5508 (N_5508,N_5106,N_5292);
and U5509 (N_5509,N_5277,N_5210);
nand U5510 (N_5510,N_5266,N_5102);
nor U5511 (N_5511,N_5273,N_5320);
or U5512 (N_5512,N_5235,N_5255);
and U5513 (N_5513,N_5328,N_5293);
nor U5514 (N_5514,N_5151,N_5223);
xor U5515 (N_5515,N_5144,N_5297);
and U5516 (N_5516,N_5280,N_5283);
nand U5517 (N_5517,N_5145,N_5278);
nor U5518 (N_5518,N_5326,N_5338);
or U5519 (N_5519,N_5351,N_5300);
xnor U5520 (N_5520,N_5243,N_5150);
and U5521 (N_5521,N_5386,N_5387);
nor U5522 (N_5522,N_5288,N_5343);
xor U5523 (N_5523,N_5394,N_5363);
nor U5524 (N_5524,N_5304,N_5275);
nand U5525 (N_5525,N_5252,N_5309);
or U5526 (N_5526,N_5135,N_5341);
nor U5527 (N_5527,N_5172,N_5276);
xnor U5528 (N_5528,N_5291,N_5168);
and U5529 (N_5529,N_5365,N_5311);
nor U5530 (N_5530,N_5185,N_5214);
nand U5531 (N_5531,N_5217,N_5238);
nor U5532 (N_5532,N_5361,N_5335);
xor U5533 (N_5533,N_5271,N_5179);
xor U5534 (N_5534,N_5380,N_5332);
nor U5535 (N_5535,N_5381,N_5250);
nor U5536 (N_5536,N_5124,N_5372);
xnor U5537 (N_5537,N_5125,N_5132);
or U5538 (N_5538,N_5352,N_5231);
or U5539 (N_5539,N_5257,N_5369);
xor U5540 (N_5540,N_5240,N_5141);
and U5541 (N_5541,N_5391,N_5115);
nor U5542 (N_5542,N_5383,N_5382);
xor U5543 (N_5543,N_5229,N_5307);
nor U5544 (N_5544,N_5353,N_5265);
xnor U5545 (N_5545,N_5239,N_5197);
and U5546 (N_5546,N_5364,N_5284);
xor U5547 (N_5547,N_5314,N_5216);
and U5548 (N_5548,N_5119,N_5340);
nand U5549 (N_5549,N_5160,N_5310);
and U5550 (N_5550,N_5102,N_5353);
or U5551 (N_5551,N_5198,N_5373);
nor U5552 (N_5552,N_5399,N_5281);
and U5553 (N_5553,N_5277,N_5264);
nand U5554 (N_5554,N_5169,N_5247);
nor U5555 (N_5555,N_5300,N_5332);
nand U5556 (N_5556,N_5294,N_5110);
nor U5557 (N_5557,N_5154,N_5182);
and U5558 (N_5558,N_5167,N_5325);
nor U5559 (N_5559,N_5134,N_5331);
and U5560 (N_5560,N_5225,N_5262);
or U5561 (N_5561,N_5311,N_5383);
or U5562 (N_5562,N_5319,N_5391);
nor U5563 (N_5563,N_5377,N_5231);
nand U5564 (N_5564,N_5150,N_5335);
and U5565 (N_5565,N_5380,N_5182);
xnor U5566 (N_5566,N_5326,N_5342);
or U5567 (N_5567,N_5212,N_5205);
xor U5568 (N_5568,N_5159,N_5160);
nor U5569 (N_5569,N_5395,N_5336);
nand U5570 (N_5570,N_5352,N_5131);
xnor U5571 (N_5571,N_5387,N_5319);
nor U5572 (N_5572,N_5174,N_5142);
nand U5573 (N_5573,N_5344,N_5240);
xor U5574 (N_5574,N_5120,N_5242);
nand U5575 (N_5575,N_5227,N_5324);
nand U5576 (N_5576,N_5129,N_5127);
and U5577 (N_5577,N_5295,N_5350);
or U5578 (N_5578,N_5299,N_5276);
or U5579 (N_5579,N_5220,N_5267);
or U5580 (N_5580,N_5132,N_5127);
or U5581 (N_5581,N_5244,N_5329);
nand U5582 (N_5582,N_5105,N_5115);
nand U5583 (N_5583,N_5191,N_5360);
nand U5584 (N_5584,N_5386,N_5375);
nand U5585 (N_5585,N_5230,N_5148);
nand U5586 (N_5586,N_5149,N_5238);
nor U5587 (N_5587,N_5166,N_5208);
xnor U5588 (N_5588,N_5148,N_5308);
and U5589 (N_5589,N_5397,N_5232);
xor U5590 (N_5590,N_5246,N_5279);
and U5591 (N_5591,N_5215,N_5153);
nand U5592 (N_5592,N_5376,N_5319);
xor U5593 (N_5593,N_5367,N_5142);
or U5594 (N_5594,N_5217,N_5276);
and U5595 (N_5595,N_5159,N_5183);
xor U5596 (N_5596,N_5131,N_5285);
and U5597 (N_5597,N_5196,N_5154);
or U5598 (N_5598,N_5249,N_5198);
and U5599 (N_5599,N_5117,N_5331);
and U5600 (N_5600,N_5235,N_5202);
nor U5601 (N_5601,N_5312,N_5232);
and U5602 (N_5602,N_5378,N_5159);
or U5603 (N_5603,N_5216,N_5372);
nor U5604 (N_5604,N_5181,N_5288);
and U5605 (N_5605,N_5115,N_5314);
xnor U5606 (N_5606,N_5252,N_5375);
nand U5607 (N_5607,N_5328,N_5308);
xnor U5608 (N_5608,N_5110,N_5295);
nor U5609 (N_5609,N_5141,N_5198);
xor U5610 (N_5610,N_5194,N_5324);
nand U5611 (N_5611,N_5363,N_5327);
xnor U5612 (N_5612,N_5172,N_5367);
or U5613 (N_5613,N_5373,N_5351);
xnor U5614 (N_5614,N_5237,N_5316);
xor U5615 (N_5615,N_5207,N_5136);
xnor U5616 (N_5616,N_5290,N_5250);
nand U5617 (N_5617,N_5186,N_5323);
and U5618 (N_5618,N_5125,N_5345);
xor U5619 (N_5619,N_5236,N_5153);
nand U5620 (N_5620,N_5322,N_5187);
or U5621 (N_5621,N_5247,N_5378);
nor U5622 (N_5622,N_5254,N_5259);
xor U5623 (N_5623,N_5140,N_5350);
nor U5624 (N_5624,N_5158,N_5196);
nand U5625 (N_5625,N_5150,N_5285);
and U5626 (N_5626,N_5179,N_5366);
xor U5627 (N_5627,N_5174,N_5237);
nor U5628 (N_5628,N_5289,N_5399);
xnor U5629 (N_5629,N_5325,N_5146);
or U5630 (N_5630,N_5106,N_5351);
nand U5631 (N_5631,N_5364,N_5237);
nor U5632 (N_5632,N_5103,N_5332);
nor U5633 (N_5633,N_5285,N_5237);
nand U5634 (N_5634,N_5187,N_5347);
nand U5635 (N_5635,N_5231,N_5149);
nand U5636 (N_5636,N_5234,N_5142);
nand U5637 (N_5637,N_5210,N_5147);
or U5638 (N_5638,N_5111,N_5186);
and U5639 (N_5639,N_5349,N_5210);
or U5640 (N_5640,N_5371,N_5144);
or U5641 (N_5641,N_5335,N_5302);
and U5642 (N_5642,N_5174,N_5252);
nor U5643 (N_5643,N_5292,N_5325);
and U5644 (N_5644,N_5181,N_5195);
and U5645 (N_5645,N_5285,N_5116);
and U5646 (N_5646,N_5321,N_5247);
or U5647 (N_5647,N_5140,N_5242);
and U5648 (N_5648,N_5248,N_5245);
nor U5649 (N_5649,N_5145,N_5300);
and U5650 (N_5650,N_5331,N_5136);
or U5651 (N_5651,N_5224,N_5167);
nor U5652 (N_5652,N_5395,N_5283);
or U5653 (N_5653,N_5246,N_5292);
and U5654 (N_5654,N_5119,N_5189);
nand U5655 (N_5655,N_5342,N_5348);
nor U5656 (N_5656,N_5249,N_5110);
or U5657 (N_5657,N_5126,N_5392);
or U5658 (N_5658,N_5367,N_5177);
or U5659 (N_5659,N_5313,N_5358);
nand U5660 (N_5660,N_5333,N_5159);
xnor U5661 (N_5661,N_5297,N_5199);
nor U5662 (N_5662,N_5262,N_5376);
nand U5663 (N_5663,N_5332,N_5273);
xnor U5664 (N_5664,N_5216,N_5388);
nand U5665 (N_5665,N_5137,N_5211);
xnor U5666 (N_5666,N_5318,N_5128);
nand U5667 (N_5667,N_5277,N_5253);
xor U5668 (N_5668,N_5326,N_5345);
xnor U5669 (N_5669,N_5167,N_5301);
and U5670 (N_5670,N_5125,N_5154);
and U5671 (N_5671,N_5237,N_5391);
and U5672 (N_5672,N_5279,N_5127);
and U5673 (N_5673,N_5362,N_5338);
xor U5674 (N_5674,N_5255,N_5214);
xor U5675 (N_5675,N_5196,N_5352);
nand U5676 (N_5676,N_5233,N_5124);
xor U5677 (N_5677,N_5340,N_5375);
nand U5678 (N_5678,N_5199,N_5393);
nor U5679 (N_5679,N_5113,N_5159);
or U5680 (N_5680,N_5353,N_5338);
or U5681 (N_5681,N_5354,N_5399);
and U5682 (N_5682,N_5247,N_5382);
xnor U5683 (N_5683,N_5226,N_5116);
and U5684 (N_5684,N_5332,N_5105);
nand U5685 (N_5685,N_5119,N_5293);
and U5686 (N_5686,N_5309,N_5105);
or U5687 (N_5687,N_5298,N_5349);
xor U5688 (N_5688,N_5177,N_5266);
nand U5689 (N_5689,N_5146,N_5151);
nand U5690 (N_5690,N_5152,N_5399);
xnor U5691 (N_5691,N_5268,N_5284);
xnor U5692 (N_5692,N_5167,N_5221);
xnor U5693 (N_5693,N_5178,N_5249);
xor U5694 (N_5694,N_5144,N_5190);
xnor U5695 (N_5695,N_5262,N_5131);
or U5696 (N_5696,N_5300,N_5344);
nand U5697 (N_5697,N_5311,N_5267);
xnor U5698 (N_5698,N_5326,N_5132);
nor U5699 (N_5699,N_5173,N_5265);
or U5700 (N_5700,N_5573,N_5482);
nand U5701 (N_5701,N_5524,N_5404);
xnor U5702 (N_5702,N_5557,N_5452);
and U5703 (N_5703,N_5442,N_5505);
xnor U5704 (N_5704,N_5409,N_5607);
and U5705 (N_5705,N_5475,N_5476);
nor U5706 (N_5706,N_5533,N_5610);
xor U5707 (N_5707,N_5497,N_5599);
and U5708 (N_5708,N_5558,N_5665);
nor U5709 (N_5709,N_5537,N_5652);
and U5710 (N_5710,N_5683,N_5563);
xnor U5711 (N_5711,N_5477,N_5565);
or U5712 (N_5712,N_5642,N_5414);
nand U5713 (N_5713,N_5663,N_5602);
nand U5714 (N_5714,N_5536,N_5673);
xnor U5715 (N_5715,N_5680,N_5647);
and U5716 (N_5716,N_5454,N_5681);
or U5717 (N_5717,N_5521,N_5440);
nor U5718 (N_5718,N_5567,N_5639);
and U5719 (N_5719,N_5522,N_5624);
or U5720 (N_5720,N_5616,N_5636);
and U5721 (N_5721,N_5572,N_5595);
nor U5722 (N_5722,N_5553,N_5604);
xnor U5723 (N_5723,N_5523,N_5662);
nor U5724 (N_5724,N_5597,N_5643);
or U5725 (N_5725,N_5661,N_5532);
nor U5726 (N_5726,N_5658,N_5619);
nor U5727 (N_5727,N_5552,N_5686);
or U5728 (N_5728,N_5418,N_5594);
and U5729 (N_5729,N_5578,N_5691);
nor U5730 (N_5730,N_5517,N_5588);
nor U5731 (N_5731,N_5651,N_5659);
xor U5732 (N_5732,N_5500,N_5462);
or U5733 (N_5733,N_5492,N_5504);
nand U5734 (N_5734,N_5582,N_5484);
and U5735 (N_5735,N_5612,N_5628);
xnor U5736 (N_5736,N_5623,N_5592);
xnor U5737 (N_5737,N_5650,N_5530);
or U5738 (N_5738,N_5626,N_5422);
xor U5739 (N_5739,N_5687,N_5561);
nor U5740 (N_5740,N_5640,N_5645);
or U5741 (N_5741,N_5449,N_5549);
nor U5742 (N_5742,N_5515,N_5471);
nor U5743 (N_5743,N_5554,N_5406);
nand U5744 (N_5744,N_5556,N_5506);
xor U5745 (N_5745,N_5575,N_5603);
nand U5746 (N_5746,N_5605,N_5544);
nor U5747 (N_5747,N_5466,N_5633);
nor U5748 (N_5748,N_5480,N_5421);
nor U5749 (N_5749,N_5630,N_5596);
nor U5750 (N_5750,N_5581,N_5423);
nor U5751 (N_5751,N_5496,N_5420);
nor U5752 (N_5752,N_5463,N_5412);
or U5753 (N_5753,N_5668,N_5540);
nor U5754 (N_5754,N_5618,N_5631);
xnor U5755 (N_5755,N_5456,N_5459);
xnor U5756 (N_5756,N_5694,N_5473);
nor U5757 (N_5757,N_5656,N_5550);
nand U5758 (N_5758,N_5629,N_5699);
and U5759 (N_5759,N_5614,N_5591);
nor U5760 (N_5760,N_5675,N_5613);
or U5761 (N_5761,N_5520,N_5510);
nor U5762 (N_5762,N_5405,N_5568);
nor U5763 (N_5763,N_5525,N_5627);
and U5764 (N_5764,N_5489,N_5464);
xor U5765 (N_5765,N_5589,N_5541);
nor U5766 (N_5766,N_5432,N_5411);
xnor U5767 (N_5767,N_5419,N_5601);
nor U5768 (N_5768,N_5664,N_5534);
nor U5769 (N_5769,N_5527,N_5427);
and U5770 (N_5770,N_5685,N_5543);
or U5771 (N_5771,N_5483,N_5696);
and U5772 (N_5772,N_5660,N_5415);
nand U5773 (N_5773,N_5470,N_5564);
nand U5774 (N_5774,N_5569,N_5439);
or U5775 (N_5775,N_5511,N_5438);
nor U5776 (N_5776,N_5674,N_5402);
and U5777 (N_5777,N_5450,N_5695);
and U5778 (N_5778,N_5469,N_5431);
xnor U5779 (N_5779,N_5494,N_5407);
nor U5780 (N_5780,N_5467,N_5598);
xor U5781 (N_5781,N_5649,N_5493);
and U5782 (N_5782,N_5555,N_5474);
nand U5783 (N_5783,N_5417,N_5670);
or U5784 (N_5784,N_5667,N_5637);
nor U5785 (N_5785,N_5646,N_5655);
nand U5786 (N_5786,N_5583,N_5512);
nand U5787 (N_5787,N_5451,N_5539);
nor U5788 (N_5788,N_5508,N_5571);
and U5789 (N_5789,N_5617,N_5485);
and U5790 (N_5790,N_5429,N_5408);
or U5791 (N_5791,N_5657,N_5446);
and U5792 (N_5792,N_5545,N_5546);
or U5793 (N_5793,N_5410,N_5559);
and U5794 (N_5794,N_5580,N_5608);
xor U5795 (N_5795,N_5453,N_5455);
xnor U5796 (N_5796,N_5577,N_5579);
nor U5797 (N_5797,N_5513,N_5606);
xor U5798 (N_5798,N_5562,N_5503);
nor U5799 (N_5799,N_5416,N_5570);
nor U5800 (N_5800,N_5516,N_5501);
and U5801 (N_5801,N_5547,N_5635);
nand U5802 (N_5802,N_5698,N_5400);
nor U5803 (N_5803,N_5528,N_5433);
and U5804 (N_5804,N_5499,N_5625);
nand U5805 (N_5805,N_5697,N_5666);
xnor U5806 (N_5806,N_5441,N_5507);
nor U5807 (N_5807,N_5529,N_5478);
nor U5808 (N_5808,N_5531,N_5479);
and U5809 (N_5809,N_5632,N_5654);
nor U5810 (N_5810,N_5689,N_5586);
or U5811 (N_5811,N_5434,N_5413);
nor U5812 (N_5812,N_5444,N_5472);
and U5813 (N_5813,N_5679,N_5600);
xnor U5814 (N_5814,N_5574,N_5488);
nor U5815 (N_5815,N_5671,N_5502);
and U5816 (N_5816,N_5535,N_5443);
nand U5817 (N_5817,N_5435,N_5678);
nand U5818 (N_5818,N_5437,N_5693);
or U5819 (N_5819,N_5430,N_5622);
xor U5820 (N_5820,N_5447,N_5584);
or U5821 (N_5821,N_5609,N_5428);
or U5822 (N_5822,N_5425,N_5620);
or U5823 (N_5823,N_5682,N_5458);
xor U5824 (N_5824,N_5486,N_5514);
nor U5825 (N_5825,N_5638,N_5587);
and U5826 (N_5826,N_5611,N_5548);
and U5827 (N_5827,N_5615,N_5672);
nor U5828 (N_5828,N_5576,N_5641);
or U5829 (N_5829,N_5490,N_5538);
or U5830 (N_5830,N_5457,N_5644);
xnor U5831 (N_5831,N_5436,N_5690);
or U5832 (N_5832,N_5426,N_5560);
or U5833 (N_5833,N_5634,N_5518);
xnor U5834 (N_5834,N_5487,N_5648);
or U5835 (N_5835,N_5465,N_5566);
or U5836 (N_5836,N_5519,N_5669);
or U5837 (N_5837,N_5653,N_5677);
xor U5838 (N_5838,N_5401,N_5509);
nand U5839 (N_5839,N_5688,N_5684);
xnor U5840 (N_5840,N_5491,N_5495);
nand U5841 (N_5841,N_5692,N_5621);
xnor U5842 (N_5842,N_5448,N_5542);
nand U5843 (N_5843,N_5460,N_5526);
xnor U5844 (N_5844,N_5551,N_5403);
and U5845 (N_5845,N_5593,N_5676);
or U5846 (N_5846,N_5461,N_5481);
and U5847 (N_5847,N_5468,N_5585);
nand U5848 (N_5848,N_5445,N_5424);
and U5849 (N_5849,N_5498,N_5590);
nor U5850 (N_5850,N_5696,N_5450);
or U5851 (N_5851,N_5500,N_5474);
or U5852 (N_5852,N_5643,N_5585);
nand U5853 (N_5853,N_5547,N_5562);
xnor U5854 (N_5854,N_5578,N_5686);
and U5855 (N_5855,N_5560,N_5580);
xnor U5856 (N_5856,N_5597,N_5606);
nand U5857 (N_5857,N_5668,N_5693);
xnor U5858 (N_5858,N_5450,N_5518);
and U5859 (N_5859,N_5430,N_5685);
nand U5860 (N_5860,N_5636,N_5604);
nand U5861 (N_5861,N_5656,N_5484);
or U5862 (N_5862,N_5480,N_5442);
xnor U5863 (N_5863,N_5459,N_5440);
and U5864 (N_5864,N_5686,N_5667);
and U5865 (N_5865,N_5653,N_5662);
xnor U5866 (N_5866,N_5402,N_5625);
and U5867 (N_5867,N_5573,N_5511);
nand U5868 (N_5868,N_5545,N_5553);
xor U5869 (N_5869,N_5628,N_5655);
or U5870 (N_5870,N_5466,N_5467);
or U5871 (N_5871,N_5575,N_5664);
or U5872 (N_5872,N_5611,N_5574);
nor U5873 (N_5873,N_5448,N_5420);
and U5874 (N_5874,N_5599,N_5494);
xor U5875 (N_5875,N_5610,N_5509);
nor U5876 (N_5876,N_5503,N_5576);
xor U5877 (N_5877,N_5577,N_5434);
or U5878 (N_5878,N_5449,N_5518);
nand U5879 (N_5879,N_5619,N_5600);
xnor U5880 (N_5880,N_5577,N_5422);
nor U5881 (N_5881,N_5446,N_5479);
nand U5882 (N_5882,N_5405,N_5461);
xor U5883 (N_5883,N_5665,N_5435);
and U5884 (N_5884,N_5408,N_5636);
nand U5885 (N_5885,N_5661,N_5494);
xnor U5886 (N_5886,N_5400,N_5568);
nand U5887 (N_5887,N_5525,N_5431);
nand U5888 (N_5888,N_5641,N_5684);
or U5889 (N_5889,N_5533,N_5553);
or U5890 (N_5890,N_5504,N_5582);
nand U5891 (N_5891,N_5574,N_5595);
nor U5892 (N_5892,N_5558,N_5529);
nor U5893 (N_5893,N_5548,N_5527);
xnor U5894 (N_5894,N_5489,N_5499);
nor U5895 (N_5895,N_5443,N_5623);
nor U5896 (N_5896,N_5664,N_5544);
nand U5897 (N_5897,N_5540,N_5697);
and U5898 (N_5898,N_5604,N_5404);
or U5899 (N_5899,N_5469,N_5602);
or U5900 (N_5900,N_5466,N_5411);
or U5901 (N_5901,N_5694,N_5638);
nor U5902 (N_5902,N_5409,N_5641);
nor U5903 (N_5903,N_5576,N_5630);
nor U5904 (N_5904,N_5438,N_5583);
and U5905 (N_5905,N_5658,N_5450);
or U5906 (N_5906,N_5566,N_5659);
or U5907 (N_5907,N_5622,N_5541);
or U5908 (N_5908,N_5527,N_5580);
or U5909 (N_5909,N_5463,N_5565);
nand U5910 (N_5910,N_5422,N_5592);
nand U5911 (N_5911,N_5462,N_5533);
or U5912 (N_5912,N_5692,N_5468);
xor U5913 (N_5913,N_5441,N_5446);
nand U5914 (N_5914,N_5578,N_5547);
and U5915 (N_5915,N_5612,N_5501);
nand U5916 (N_5916,N_5631,N_5601);
or U5917 (N_5917,N_5668,N_5503);
nand U5918 (N_5918,N_5496,N_5578);
nand U5919 (N_5919,N_5490,N_5504);
and U5920 (N_5920,N_5652,N_5603);
and U5921 (N_5921,N_5439,N_5551);
xor U5922 (N_5922,N_5439,N_5601);
xnor U5923 (N_5923,N_5598,N_5613);
nand U5924 (N_5924,N_5691,N_5470);
or U5925 (N_5925,N_5611,N_5530);
xor U5926 (N_5926,N_5562,N_5410);
or U5927 (N_5927,N_5645,N_5550);
nor U5928 (N_5928,N_5504,N_5643);
xnor U5929 (N_5929,N_5688,N_5485);
and U5930 (N_5930,N_5554,N_5479);
and U5931 (N_5931,N_5677,N_5643);
nor U5932 (N_5932,N_5489,N_5423);
and U5933 (N_5933,N_5473,N_5470);
or U5934 (N_5934,N_5596,N_5478);
xor U5935 (N_5935,N_5638,N_5407);
and U5936 (N_5936,N_5509,N_5697);
nand U5937 (N_5937,N_5660,N_5464);
and U5938 (N_5938,N_5527,N_5600);
xnor U5939 (N_5939,N_5455,N_5437);
or U5940 (N_5940,N_5636,N_5575);
or U5941 (N_5941,N_5576,N_5541);
or U5942 (N_5942,N_5613,N_5491);
or U5943 (N_5943,N_5493,N_5618);
xor U5944 (N_5944,N_5418,N_5443);
nand U5945 (N_5945,N_5419,N_5545);
nand U5946 (N_5946,N_5517,N_5434);
xnor U5947 (N_5947,N_5579,N_5597);
nor U5948 (N_5948,N_5511,N_5653);
and U5949 (N_5949,N_5641,N_5575);
nand U5950 (N_5950,N_5579,N_5529);
xnor U5951 (N_5951,N_5451,N_5643);
nand U5952 (N_5952,N_5600,N_5698);
nand U5953 (N_5953,N_5519,N_5620);
and U5954 (N_5954,N_5560,N_5438);
or U5955 (N_5955,N_5514,N_5455);
nand U5956 (N_5956,N_5536,N_5460);
nand U5957 (N_5957,N_5627,N_5662);
and U5958 (N_5958,N_5471,N_5609);
nand U5959 (N_5959,N_5497,N_5675);
nor U5960 (N_5960,N_5461,N_5451);
nor U5961 (N_5961,N_5431,N_5669);
nor U5962 (N_5962,N_5656,N_5591);
nor U5963 (N_5963,N_5584,N_5508);
and U5964 (N_5964,N_5520,N_5630);
or U5965 (N_5965,N_5548,N_5539);
or U5966 (N_5966,N_5425,N_5468);
and U5967 (N_5967,N_5493,N_5686);
or U5968 (N_5968,N_5664,N_5675);
or U5969 (N_5969,N_5633,N_5593);
and U5970 (N_5970,N_5636,N_5436);
xnor U5971 (N_5971,N_5524,N_5528);
xor U5972 (N_5972,N_5619,N_5693);
or U5973 (N_5973,N_5526,N_5531);
xor U5974 (N_5974,N_5625,N_5483);
or U5975 (N_5975,N_5505,N_5413);
nor U5976 (N_5976,N_5589,N_5512);
nor U5977 (N_5977,N_5677,N_5648);
and U5978 (N_5978,N_5471,N_5590);
or U5979 (N_5979,N_5616,N_5499);
xnor U5980 (N_5980,N_5458,N_5509);
and U5981 (N_5981,N_5452,N_5544);
or U5982 (N_5982,N_5529,N_5580);
and U5983 (N_5983,N_5569,N_5662);
or U5984 (N_5984,N_5675,N_5472);
nor U5985 (N_5985,N_5442,N_5479);
xor U5986 (N_5986,N_5601,N_5422);
and U5987 (N_5987,N_5459,N_5563);
nand U5988 (N_5988,N_5555,N_5621);
nor U5989 (N_5989,N_5653,N_5638);
nand U5990 (N_5990,N_5531,N_5683);
nor U5991 (N_5991,N_5631,N_5585);
or U5992 (N_5992,N_5699,N_5462);
nor U5993 (N_5993,N_5603,N_5596);
nor U5994 (N_5994,N_5630,N_5664);
or U5995 (N_5995,N_5564,N_5589);
xor U5996 (N_5996,N_5415,N_5646);
xnor U5997 (N_5997,N_5679,N_5560);
xor U5998 (N_5998,N_5607,N_5500);
nand U5999 (N_5999,N_5504,N_5557);
nor U6000 (N_6000,N_5798,N_5966);
or U6001 (N_6001,N_5864,N_5813);
xnor U6002 (N_6002,N_5987,N_5846);
nor U6003 (N_6003,N_5869,N_5965);
xor U6004 (N_6004,N_5716,N_5859);
or U6005 (N_6005,N_5794,N_5911);
nor U6006 (N_6006,N_5816,N_5978);
nor U6007 (N_6007,N_5962,N_5909);
xor U6008 (N_6008,N_5845,N_5931);
or U6009 (N_6009,N_5944,N_5988);
nand U6010 (N_6010,N_5884,N_5760);
xnor U6011 (N_6011,N_5995,N_5939);
nor U6012 (N_6012,N_5810,N_5873);
and U6013 (N_6013,N_5901,N_5967);
or U6014 (N_6014,N_5743,N_5889);
xor U6015 (N_6015,N_5914,N_5976);
or U6016 (N_6016,N_5842,N_5768);
or U6017 (N_6017,N_5817,N_5999);
or U6018 (N_6018,N_5941,N_5996);
and U6019 (N_6019,N_5828,N_5740);
and U6020 (N_6020,N_5912,N_5910);
or U6021 (N_6021,N_5879,N_5839);
or U6022 (N_6022,N_5757,N_5748);
or U6023 (N_6023,N_5886,N_5756);
nor U6024 (N_6024,N_5936,N_5770);
nand U6025 (N_6025,N_5858,N_5727);
xor U6026 (N_6026,N_5706,N_5904);
xor U6027 (N_6027,N_5883,N_5733);
nand U6028 (N_6028,N_5862,N_5834);
and U6029 (N_6029,N_5829,N_5715);
and U6030 (N_6030,N_5782,N_5949);
or U6031 (N_6031,N_5826,N_5942);
and U6032 (N_6032,N_5735,N_5890);
nor U6033 (N_6033,N_5950,N_5796);
nand U6034 (N_6034,N_5855,N_5710);
xor U6035 (N_6035,N_5778,N_5811);
nor U6036 (N_6036,N_5970,N_5874);
or U6037 (N_6037,N_5744,N_5801);
nor U6038 (N_6038,N_5948,N_5878);
nand U6039 (N_6039,N_5924,N_5713);
nor U6040 (N_6040,N_5865,N_5892);
or U6041 (N_6041,N_5926,N_5933);
xnor U6042 (N_6042,N_5762,N_5902);
and U6043 (N_6043,N_5785,N_5986);
and U6044 (N_6044,N_5788,N_5885);
nor U6045 (N_6045,N_5871,N_5791);
or U6046 (N_6046,N_5860,N_5827);
nor U6047 (N_6047,N_5964,N_5849);
nor U6048 (N_6048,N_5711,N_5701);
and U6049 (N_6049,N_5998,N_5705);
or U6050 (N_6050,N_5857,N_5917);
or U6051 (N_6051,N_5887,N_5900);
and U6052 (N_6052,N_5784,N_5968);
nor U6053 (N_6053,N_5803,N_5937);
and U6054 (N_6054,N_5983,N_5877);
nand U6055 (N_6055,N_5905,N_5702);
nand U6056 (N_6056,N_5763,N_5789);
and U6057 (N_6057,N_5835,N_5891);
nor U6058 (N_6058,N_5809,N_5847);
or U6059 (N_6059,N_5730,N_5831);
nor U6060 (N_6060,N_5940,N_5844);
and U6061 (N_6061,N_5703,N_5752);
nor U6062 (N_6062,N_5928,N_5707);
xor U6063 (N_6063,N_5738,N_5975);
xor U6064 (N_6064,N_5749,N_5758);
nor U6065 (N_6065,N_5704,N_5938);
and U6066 (N_6066,N_5822,N_5898);
and U6067 (N_6067,N_5896,N_5807);
or U6068 (N_6068,N_5766,N_5908);
nand U6069 (N_6069,N_5947,N_5952);
xor U6070 (N_6070,N_5830,N_5991);
and U6071 (N_6071,N_5953,N_5870);
nor U6072 (N_6072,N_5951,N_5843);
nand U6073 (N_6073,N_5802,N_5765);
and U6074 (N_6074,N_5754,N_5872);
and U6075 (N_6075,N_5934,N_5919);
and U6076 (N_6076,N_5994,N_5806);
and U6077 (N_6077,N_5804,N_5927);
or U6078 (N_6078,N_5774,N_5984);
or U6079 (N_6079,N_5741,N_5981);
or U6080 (N_6080,N_5915,N_5814);
nor U6081 (N_6081,N_5923,N_5974);
nand U6082 (N_6082,N_5786,N_5720);
nand U6083 (N_6083,N_5742,N_5734);
and U6084 (N_6084,N_5880,N_5840);
nor U6085 (N_6085,N_5795,N_5866);
or U6086 (N_6086,N_5867,N_5719);
nand U6087 (N_6087,N_5850,N_5812);
and U6088 (N_6088,N_5722,N_5751);
nand U6089 (N_6089,N_5989,N_5985);
nand U6090 (N_6090,N_5956,N_5815);
and U6091 (N_6091,N_5781,N_5990);
xor U6092 (N_6092,N_5980,N_5709);
and U6093 (N_6093,N_5777,N_5712);
and U6094 (N_6094,N_5750,N_5838);
nand U6095 (N_6095,N_5739,N_5856);
nor U6096 (N_6096,N_5775,N_5823);
nor U6097 (N_6097,N_5893,N_5776);
or U6098 (N_6098,N_5800,N_5783);
nor U6099 (N_6099,N_5961,N_5745);
or U6100 (N_6100,N_5755,N_5818);
nor U6101 (N_6101,N_5841,N_5759);
or U6102 (N_6102,N_5913,N_5851);
nand U6103 (N_6103,N_5888,N_5824);
nor U6104 (N_6104,N_5725,N_5767);
and U6105 (N_6105,N_5921,N_5732);
and U6106 (N_6106,N_5746,N_5821);
or U6107 (N_6107,N_5916,N_5932);
and U6108 (N_6108,N_5979,N_5906);
or U6109 (N_6109,N_5882,N_5971);
and U6110 (N_6110,N_5929,N_5922);
nor U6111 (N_6111,N_5875,N_5997);
xnor U6112 (N_6112,N_5772,N_5714);
and U6113 (N_6113,N_5779,N_5832);
xor U6114 (N_6114,N_5700,N_5769);
nor U6115 (N_6115,N_5761,N_5868);
nand U6116 (N_6116,N_5805,N_5993);
or U6117 (N_6117,N_5957,N_5881);
and U6118 (N_6118,N_5854,N_5895);
nor U6119 (N_6119,N_5771,N_5920);
or U6120 (N_6120,N_5819,N_5946);
xor U6121 (N_6121,N_5973,N_5897);
xnor U6122 (N_6122,N_5736,N_5969);
and U6123 (N_6123,N_5861,N_5797);
and U6124 (N_6124,N_5992,N_5925);
xnor U6125 (N_6125,N_5787,N_5836);
and U6126 (N_6126,N_5708,N_5825);
nor U6127 (N_6127,N_5930,N_5721);
xor U6128 (N_6128,N_5780,N_5753);
nand U6129 (N_6129,N_5955,N_5833);
and U6130 (N_6130,N_5729,N_5863);
xnor U6131 (N_6131,N_5737,N_5899);
or U6132 (N_6132,N_5731,N_5977);
nand U6133 (N_6133,N_5960,N_5958);
nand U6134 (N_6134,N_5790,N_5907);
and U6135 (N_6135,N_5728,N_5853);
nand U6136 (N_6136,N_5718,N_5852);
and U6137 (N_6137,N_5723,N_5959);
nor U6138 (N_6138,N_5945,N_5972);
xnor U6139 (N_6139,N_5837,N_5726);
xor U6140 (N_6140,N_5792,N_5935);
nor U6141 (N_6141,N_5876,N_5982);
and U6142 (N_6142,N_5820,N_5773);
and U6143 (N_6143,N_5918,N_5894);
nor U6144 (N_6144,N_5808,N_5764);
xor U6145 (N_6145,N_5963,N_5799);
or U6146 (N_6146,N_5717,N_5724);
xor U6147 (N_6147,N_5943,N_5848);
xnor U6148 (N_6148,N_5793,N_5903);
or U6149 (N_6149,N_5954,N_5747);
nor U6150 (N_6150,N_5981,N_5797);
nand U6151 (N_6151,N_5975,N_5954);
nor U6152 (N_6152,N_5731,N_5914);
xnor U6153 (N_6153,N_5857,N_5950);
nor U6154 (N_6154,N_5974,N_5903);
or U6155 (N_6155,N_5925,N_5759);
nand U6156 (N_6156,N_5928,N_5730);
nand U6157 (N_6157,N_5741,N_5885);
xor U6158 (N_6158,N_5818,N_5840);
nand U6159 (N_6159,N_5906,N_5970);
and U6160 (N_6160,N_5857,N_5821);
and U6161 (N_6161,N_5875,N_5756);
nand U6162 (N_6162,N_5895,N_5887);
or U6163 (N_6163,N_5891,N_5904);
nor U6164 (N_6164,N_5996,N_5851);
xor U6165 (N_6165,N_5862,N_5926);
nand U6166 (N_6166,N_5815,N_5979);
and U6167 (N_6167,N_5769,N_5992);
and U6168 (N_6168,N_5993,N_5938);
or U6169 (N_6169,N_5905,N_5874);
and U6170 (N_6170,N_5843,N_5960);
xnor U6171 (N_6171,N_5969,N_5959);
nand U6172 (N_6172,N_5823,N_5751);
nor U6173 (N_6173,N_5966,N_5726);
or U6174 (N_6174,N_5717,N_5854);
nor U6175 (N_6175,N_5893,N_5768);
xor U6176 (N_6176,N_5973,N_5910);
or U6177 (N_6177,N_5799,N_5826);
or U6178 (N_6178,N_5911,N_5820);
xor U6179 (N_6179,N_5966,N_5789);
nand U6180 (N_6180,N_5733,N_5752);
xor U6181 (N_6181,N_5779,N_5796);
and U6182 (N_6182,N_5833,N_5952);
nor U6183 (N_6183,N_5773,N_5899);
nand U6184 (N_6184,N_5934,N_5766);
xnor U6185 (N_6185,N_5971,N_5972);
nand U6186 (N_6186,N_5789,N_5856);
nor U6187 (N_6187,N_5998,N_5997);
or U6188 (N_6188,N_5900,N_5782);
or U6189 (N_6189,N_5921,N_5816);
nor U6190 (N_6190,N_5756,N_5732);
or U6191 (N_6191,N_5960,N_5982);
nor U6192 (N_6192,N_5846,N_5713);
nand U6193 (N_6193,N_5860,N_5858);
xnor U6194 (N_6194,N_5984,N_5828);
nor U6195 (N_6195,N_5878,N_5763);
xnor U6196 (N_6196,N_5776,N_5996);
xnor U6197 (N_6197,N_5708,N_5796);
xnor U6198 (N_6198,N_5846,N_5764);
nand U6199 (N_6199,N_5717,N_5888);
nor U6200 (N_6200,N_5807,N_5799);
nand U6201 (N_6201,N_5844,N_5809);
or U6202 (N_6202,N_5915,N_5864);
nor U6203 (N_6203,N_5987,N_5978);
nand U6204 (N_6204,N_5845,N_5727);
and U6205 (N_6205,N_5736,N_5741);
xnor U6206 (N_6206,N_5940,N_5814);
and U6207 (N_6207,N_5824,N_5959);
and U6208 (N_6208,N_5927,N_5875);
and U6209 (N_6209,N_5929,N_5703);
nor U6210 (N_6210,N_5730,N_5742);
nor U6211 (N_6211,N_5820,N_5883);
or U6212 (N_6212,N_5960,N_5767);
nor U6213 (N_6213,N_5977,N_5849);
and U6214 (N_6214,N_5718,N_5784);
nor U6215 (N_6215,N_5901,N_5960);
nand U6216 (N_6216,N_5942,N_5748);
nor U6217 (N_6217,N_5755,N_5854);
and U6218 (N_6218,N_5813,N_5769);
or U6219 (N_6219,N_5922,N_5830);
nand U6220 (N_6220,N_5846,N_5916);
nand U6221 (N_6221,N_5789,N_5880);
and U6222 (N_6222,N_5787,N_5811);
or U6223 (N_6223,N_5785,N_5788);
nor U6224 (N_6224,N_5843,N_5954);
nor U6225 (N_6225,N_5969,N_5719);
nand U6226 (N_6226,N_5803,N_5879);
xnor U6227 (N_6227,N_5749,N_5844);
nand U6228 (N_6228,N_5899,N_5722);
xnor U6229 (N_6229,N_5780,N_5978);
nor U6230 (N_6230,N_5919,N_5861);
nor U6231 (N_6231,N_5771,N_5923);
nand U6232 (N_6232,N_5977,N_5752);
nor U6233 (N_6233,N_5829,N_5951);
or U6234 (N_6234,N_5761,N_5839);
and U6235 (N_6235,N_5844,N_5801);
xnor U6236 (N_6236,N_5955,N_5904);
nor U6237 (N_6237,N_5823,N_5707);
and U6238 (N_6238,N_5945,N_5941);
nor U6239 (N_6239,N_5801,N_5991);
xor U6240 (N_6240,N_5747,N_5851);
nor U6241 (N_6241,N_5763,N_5952);
nand U6242 (N_6242,N_5930,N_5966);
or U6243 (N_6243,N_5744,N_5931);
and U6244 (N_6244,N_5986,N_5963);
xor U6245 (N_6245,N_5913,N_5827);
nor U6246 (N_6246,N_5716,N_5732);
nand U6247 (N_6247,N_5932,N_5994);
or U6248 (N_6248,N_5844,N_5776);
xor U6249 (N_6249,N_5790,N_5903);
nand U6250 (N_6250,N_5859,N_5976);
xnor U6251 (N_6251,N_5959,N_5924);
and U6252 (N_6252,N_5890,N_5745);
xnor U6253 (N_6253,N_5774,N_5803);
nor U6254 (N_6254,N_5808,N_5757);
xnor U6255 (N_6255,N_5863,N_5908);
nor U6256 (N_6256,N_5712,N_5799);
xnor U6257 (N_6257,N_5961,N_5920);
xor U6258 (N_6258,N_5995,N_5857);
and U6259 (N_6259,N_5965,N_5807);
nor U6260 (N_6260,N_5917,N_5833);
or U6261 (N_6261,N_5884,N_5942);
nor U6262 (N_6262,N_5958,N_5795);
or U6263 (N_6263,N_5921,N_5712);
and U6264 (N_6264,N_5962,N_5925);
xor U6265 (N_6265,N_5888,N_5848);
and U6266 (N_6266,N_5942,N_5789);
or U6267 (N_6267,N_5859,N_5840);
nor U6268 (N_6268,N_5772,N_5747);
and U6269 (N_6269,N_5756,N_5791);
xnor U6270 (N_6270,N_5932,N_5998);
xor U6271 (N_6271,N_5852,N_5767);
nand U6272 (N_6272,N_5898,N_5792);
xnor U6273 (N_6273,N_5884,N_5951);
and U6274 (N_6274,N_5983,N_5882);
nand U6275 (N_6275,N_5745,N_5928);
xnor U6276 (N_6276,N_5886,N_5718);
nand U6277 (N_6277,N_5992,N_5777);
and U6278 (N_6278,N_5969,N_5979);
or U6279 (N_6279,N_5814,N_5762);
xnor U6280 (N_6280,N_5707,N_5869);
nand U6281 (N_6281,N_5909,N_5812);
and U6282 (N_6282,N_5864,N_5887);
nand U6283 (N_6283,N_5792,N_5745);
xnor U6284 (N_6284,N_5791,N_5984);
nand U6285 (N_6285,N_5912,N_5972);
and U6286 (N_6286,N_5862,N_5785);
xnor U6287 (N_6287,N_5914,N_5902);
and U6288 (N_6288,N_5708,N_5788);
nand U6289 (N_6289,N_5795,N_5995);
xnor U6290 (N_6290,N_5705,N_5720);
nor U6291 (N_6291,N_5923,N_5755);
or U6292 (N_6292,N_5742,N_5861);
nor U6293 (N_6293,N_5901,N_5702);
nand U6294 (N_6294,N_5825,N_5743);
nand U6295 (N_6295,N_5888,N_5940);
or U6296 (N_6296,N_5807,N_5732);
xor U6297 (N_6297,N_5772,N_5818);
nand U6298 (N_6298,N_5862,N_5767);
xnor U6299 (N_6299,N_5873,N_5869);
nor U6300 (N_6300,N_6122,N_6108);
nand U6301 (N_6301,N_6261,N_6061);
nor U6302 (N_6302,N_6299,N_6185);
nor U6303 (N_6303,N_6014,N_6000);
or U6304 (N_6304,N_6234,N_6175);
or U6305 (N_6305,N_6111,N_6093);
nor U6306 (N_6306,N_6121,N_6103);
xor U6307 (N_6307,N_6079,N_6206);
nor U6308 (N_6308,N_6073,N_6054);
nor U6309 (N_6309,N_6156,N_6126);
or U6310 (N_6310,N_6099,N_6065);
or U6311 (N_6311,N_6159,N_6056);
xnor U6312 (N_6312,N_6050,N_6043);
or U6313 (N_6313,N_6124,N_6030);
nand U6314 (N_6314,N_6135,N_6214);
or U6315 (N_6315,N_6213,N_6114);
or U6316 (N_6316,N_6259,N_6171);
and U6317 (N_6317,N_6033,N_6205);
or U6318 (N_6318,N_6026,N_6128);
and U6319 (N_6319,N_6029,N_6215);
and U6320 (N_6320,N_6230,N_6285);
or U6321 (N_6321,N_6109,N_6177);
nand U6322 (N_6322,N_6264,N_6241);
xor U6323 (N_6323,N_6148,N_6019);
nand U6324 (N_6324,N_6203,N_6252);
xnor U6325 (N_6325,N_6157,N_6196);
nor U6326 (N_6326,N_6219,N_6134);
or U6327 (N_6327,N_6199,N_6220);
xor U6328 (N_6328,N_6039,N_6211);
nand U6329 (N_6329,N_6223,N_6036);
nand U6330 (N_6330,N_6074,N_6001);
xnor U6331 (N_6331,N_6145,N_6044);
xor U6332 (N_6332,N_6201,N_6105);
xor U6333 (N_6333,N_6077,N_6191);
and U6334 (N_6334,N_6198,N_6067);
nand U6335 (N_6335,N_6084,N_6282);
nor U6336 (N_6336,N_6080,N_6060);
and U6337 (N_6337,N_6130,N_6286);
nor U6338 (N_6338,N_6270,N_6104);
xnor U6339 (N_6339,N_6020,N_6255);
or U6340 (N_6340,N_6218,N_6209);
xor U6341 (N_6341,N_6257,N_6140);
nand U6342 (N_6342,N_6064,N_6151);
or U6343 (N_6343,N_6256,N_6042);
and U6344 (N_6344,N_6136,N_6069);
or U6345 (N_6345,N_6047,N_6132);
nand U6346 (N_6346,N_6266,N_6248);
or U6347 (N_6347,N_6155,N_6166);
nand U6348 (N_6348,N_6150,N_6037);
and U6349 (N_6349,N_6202,N_6267);
nor U6350 (N_6350,N_6070,N_6072);
and U6351 (N_6351,N_6032,N_6193);
and U6352 (N_6352,N_6028,N_6189);
or U6353 (N_6353,N_6051,N_6129);
or U6354 (N_6354,N_6204,N_6007);
xor U6355 (N_6355,N_6058,N_6127);
nor U6356 (N_6356,N_6002,N_6228);
xnor U6357 (N_6357,N_6290,N_6237);
xor U6358 (N_6358,N_6287,N_6115);
or U6359 (N_6359,N_6279,N_6097);
nor U6360 (N_6360,N_6227,N_6200);
xor U6361 (N_6361,N_6053,N_6249);
or U6362 (N_6362,N_6003,N_6005);
nand U6363 (N_6363,N_6146,N_6075);
and U6364 (N_6364,N_6041,N_6260);
nand U6365 (N_6365,N_6207,N_6018);
or U6366 (N_6366,N_6046,N_6123);
and U6367 (N_6367,N_6274,N_6263);
or U6368 (N_6368,N_6294,N_6055);
and U6369 (N_6369,N_6226,N_6297);
and U6370 (N_6370,N_6068,N_6147);
and U6371 (N_6371,N_6245,N_6008);
nand U6372 (N_6372,N_6078,N_6288);
or U6373 (N_6373,N_6062,N_6182);
xnor U6374 (N_6374,N_6141,N_6293);
or U6375 (N_6375,N_6277,N_6106);
and U6376 (N_6376,N_6035,N_6283);
nor U6377 (N_6377,N_6059,N_6027);
nor U6378 (N_6378,N_6164,N_6197);
nor U6379 (N_6379,N_6083,N_6246);
and U6380 (N_6380,N_6170,N_6125);
nor U6381 (N_6381,N_6190,N_6243);
nor U6382 (N_6382,N_6173,N_6268);
and U6383 (N_6383,N_6149,N_6269);
or U6384 (N_6384,N_6284,N_6253);
xor U6385 (N_6385,N_6210,N_6165);
or U6386 (N_6386,N_6112,N_6242);
xnor U6387 (N_6387,N_6162,N_6212);
and U6388 (N_6388,N_6086,N_6233);
and U6389 (N_6389,N_6089,N_6231);
nor U6390 (N_6390,N_6119,N_6280);
or U6391 (N_6391,N_6222,N_6172);
xnor U6392 (N_6392,N_6240,N_6163);
and U6393 (N_6393,N_6031,N_6258);
and U6394 (N_6394,N_6076,N_6013);
nor U6395 (N_6395,N_6009,N_6022);
nand U6396 (N_6396,N_6038,N_6120);
nor U6397 (N_6397,N_6102,N_6006);
or U6398 (N_6398,N_6158,N_6271);
or U6399 (N_6399,N_6168,N_6094);
nor U6400 (N_6400,N_6152,N_6217);
nand U6401 (N_6401,N_6278,N_6281);
nor U6402 (N_6402,N_6088,N_6116);
nand U6403 (N_6403,N_6138,N_6174);
and U6404 (N_6404,N_6092,N_6024);
or U6405 (N_6405,N_6265,N_6110);
xor U6406 (N_6406,N_6133,N_6034);
and U6407 (N_6407,N_6161,N_6023);
or U6408 (N_6408,N_6186,N_6160);
or U6409 (N_6409,N_6082,N_6250);
and U6410 (N_6410,N_6276,N_6113);
xor U6411 (N_6411,N_6180,N_6183);
xnor U6412 (N_6412,N_6131,N_6272);
nand U6413 (N_6413,N_6224,N_6187);
and U6414 (N_6414,N_6154,N_6045);
nand U6415 (N_6415,N_6235,N_6063);
nor U6416 (N_6416,N_6225,N_6275);
or U6417 (N_6417,N_6291,N_6208);
nor U6418 (N_6418,N_6236,N_6244);
and U6419 (N_6419,N_6012,N_6017);
and U6420 (N_6420,N_6100,N_6107);
or U6421 (N_6421,N_6081,N_6021);
or U6422 (N_6422,N_6239,N_6167);
xnor U6423 (N_6423,N_6296,N_6048);
nor U6424 (N_6424,N_6262,N_6101);
or U6425 (N_6425,N_6025,N_6091);
and U6426 (N_6426,N_6142,N_6085);
and U6427 (N_6427,N_6137,N_6143);
xor U6428 (N_6428,N_6216,N_6251);
nand U6429 (N_6429,N_6153,N_6016);
nor U6430 (N_6430,N_6178,N_6071);
and U6431 (N_6431,N_6188,N_6169);
and U6432 (N_6432,N_6117,N_6176);
and U6433 (N_6433,N_6295,N_6004);
nand U6434 (N_6434,N_6049,N_6232);
nor U6435 (N_6435,N_6221,N_6098);
and U6436 (N_6436,N_6040,N_6192);
nand U6437 (N_6437,N_6057,N_6010);
or U6438 (N_6438,N_6179,N_6144);
xnor U6439 (N_6439,N_6087,N_6118);
nand U6440 (N_6440,N_6254,N_6052);
nor U6441 (N_6441,N_6011,N_6298);
xnor U6442 (N_6442,N_6139,N_6238);
or U6443 (N_6443,N_6090,N_6181);
and U6444 (N_6444,N_6292,N_6247);
and U6445 (N_6445,N_6015,N_6195);
or U6446 (N_6446,N_6096,N_6194);
nand U6447 (N_6447,N_6184,N_6095);
and U6448 (N_6448,N_6289,N_6229);
or U6449 (N_6449,N_6273,N_6066);
xnor U6450 (N_6450,N_6027,N_6186);
and U6451 (N_6451,N_6098,N_6274);
nand U6452 (N_6452,N_6104,N_6250);
xnor U6453 (N_6453,N_6234,N_6118);
nand U6454 (N_6454,N_6188,N_6281);
and U6455 (N_6455,N_6059,N_6055);
nor U6456 (N_6456,N_6171,N_6057);
xnor U6457 (N_6457,N_6135,N_6050);
and U6458 (N_6458,N_6023,N_6053);
nand U6459 (N_6459,N_6289,N_6104);
or U6460 (N_6460,N_6008,N_6274);
xnor U6461 (N_6461,N_6056,N_6198);
and U6462 (N_6462,N_6166,N_6022);
or U6463 (N_6463,N_6163,N_6281);
nor U6464 (N_6464,N_6010,N_6211);
xnor U6465 (N_6465,N_6121,N_6021);
or U6466 (N_6466,N_6057,N_6262);
xnor U6467 (N_6467,N_6212,N_6236);
xnor U6468 (N_6468,N_6007,N_6225);
and U6469 (N_6469,N_6215,N_6025);
nor U6470 (N_6470,N_6298,N_6201);
nor U6471 (N_6471,N_6098,N_6242);
xnor U6472 (N_6472,N_6186,N_6019);
or U6473 (N_6473,N_6173,N_6262);
xor U6474 (N_6474,N_6161,N_6147);
and U6475 (N_6475,N_6247,N_6171);
nand U6476 (N_6476,N_6248,N_6141);
xnor U6477 (N_6477,N_6111,N_6187);
nor U6478 (N_6478,N_6180,N_6193);
xnor U6479 (N_6479,N_6119,N_6203);
nor U6480 (N_6480,N_6184,N_6024);
nor U6481 (N_6481,N_6172,N_6272);
or U6482 (N_6482,N_6089,N_6060);
nand U6483 (N_6483,N_6131,N_6012);
xor U6484 (N_6484,N_6174,N_6226);
nor U6485 (N_6485,N_6114,N_6277);
nand U6486 (N_6486,N_6105,N_6196);
or U6487 (N_6487,N_6282,N_6115);
nand U6488 (N_6488,N_6290,N_6182);
nor U6489 (N_6489,N_6251,N_6069);
nand U6490 (N_6490,N_6001,N_6283);
and U6491 (N_6491,N_6237,N_6226);
nand U6492 (N_6492,N_6251,N_6126);
xor U6493 (N_6493,N_6242,N_6106);
nor U6494 (N_6494,N_6144,N_6160);
nand U6495 (N_6495,N_6142,N_6101);
nand U6496 (N_6496,N_6116,N_6006);
xor U6497 (N_6497,N_6262,N_6066);
and U6498 (N_6498,N_6055,N_6147);
nand U6499 (N_6499,N_6083,N_6182);
xnor U6500 (N_6500,N_6067,N_6294);
nand U6501 (N_6501,N_6215,N_6287);
or U6502 (N_6502,N_6104,N_6111);
nor U6503 (N_6503,N_6236,N_6050);
and U6504 (N_6504,N_6022,N_6014);
or U6505 (N_6505,N_6069,N_6111);
or U6506 (N_6506,N_6189,N_6008);
or U6507 (N_6507,N_6189,N_6123);
or U6508 (N_6508,N_6192,N_6234);
nor U6509 (N_6509,N_6048,N_6119);
xnor U6510 (N_6510,N_6129,N_6265);
nand U6511 (N_6511,N_6214,N_6208);
or U6512 (N_6512,N_6254,N_6128);
and U6513 (N_6513,N_6154,N_6293);
or U6514 (N_6514,N_6151,N_6234);
and U6515 (N_6515,N_6132,N_6095);
or U6516 (N_6516,N_6152,N_6006);
nand U6517 (N_6517,N_6205,N_6079);
xor U6518 (N_6518,N_6118,N_6031);
and U6519 (N_6519,N_6096,N_6279);
or U6520 (N_6520,N_6146,N_6053);
and U6521 (N_6521,N_6193,N_6249);
nor U6522 (N_6522,N_6007,N_6065);
nor U6523 (N_6523,N_6106,N_6132);
or U6524 (N_6524,N_6024,N_6025);
or U6525 (N_6525,N_6123,N_6108);
nor U6526 (N_6526,N_6255,N_6191);
or U6527 (N_6527,N_6018,N_6210);
nor U6528 (N_6528,N_6259,N_6060);
nor U6529 (N_6529,N_6229,N_6017);
nand U6530 (N_6530,N_6186,N_6116);
nand U6531 (N_6531,N_6053,N_6126);
nand U6532 (N_6532,N_6167,N_6016);
nand U6533 (N_6533,N_6064,N_6037);
xor U6534 (N_6534,N_6049,N_6203);
and U6535 (N_6535,N_6019,N_6164);
and U6536 (N_6536,N_6138,N_6103);
or U6537 (N_6537,N_6164,N_6045);
nor U6538 (N_6538,N_6143,N_6130);
or U6539 (N_6539,N_6072,N_6098);
nor U6540 (N_6540,N_6007,N_6032);
xnor U6541 (N_6541,N_6205,N_6255);
and U6542 (N_6542,N_6257,N_6214);
nand U6543 (N_6543,N_6033,N_6042);
and U6544 (N_6544,N_6183,N_6250);
xor U6545 (N_6545,N_6252,N_6022);
or U6546 (N_6546,N_6231,N_6026);
xor U6547 (N_6547,N_6179,N_6184);
and U6548 (N_6548,N_6136,N_6235);
xor U6549 (N_6549,N_6206,N_6184);
nor U6550 (N_6550,N_6037,N_6090);
xnor U6551 (N_6551,N_6065,N_6059);
and U6552 (N_6552,N_6049,N_6075);
xor U6553 (N_6553,N_6000,N_6242);
or U6554 (N_6554,N_6272,N_6151);
xor U6555 (N_6555,N_6132,N_6068);
or U6556 (N_6556,N_6225,N_6260);
xor U6557 (N_6557,N_6098,N_6150);
and U6558 (N_6558,N_6066,N_6246);
nor U6559 (N_6559,N_6180,N_6151);
or U6560 (N_6560,N_6081,N_6214);
nor U6561 (N_6561,N_6066,N_6239);
xor U6562 (N_6562,N_6132,N_6185);
nand U6563 (N_6563,N_6140,N_6077);
or U6564 (N_6564,N_6094,N_6073);
or U6565 (N_6565,N_6111,N_6058);
and U6566 (N_6566,N_6294,N_6206);
nand U6567 (N_6567,N_6289,N_6262);
nor U6568 (N_6568,N_6235,N_6203);
or U6569 (N_6569,N_6270,N_6224);
or U6570 (N_6570,N_6192,N_6103);
nand U6571 (N_6571,N_6140,N_6149);
xor U6572 (N_6572,N_6284,N_6266);
and U6573 (N_6573,N_6175,N_6040);
nor U6574 (N_6574,N_6098,N_6086);
nor U6575 (N_6575,N_6178,N_6112);
nor U6576 (N_6576,N_6109,N_6265);
or U6577 (N_6577,N_6169,N_6099);
and U6578 (N_6578,N_6291,N_6072);
nand U6579 (N_6579,N_6164,N_6013);
and U6580 (N_6580,N_6279,N_6024);
nor U6581 (N_6581,N_6241,N_6080);
nand U6582 (N_6582,N_6241,N_6061);
nand U6583 (N_6583,N_6237,N_6299);
or U6584 (N_6584,N_6172,N_6028);
xnor U6585 (N_6585,N_6116,N_6264);
or U6586 (N_6586,N_6086,N_6204);
xor U6587 (N_6587,N_6044,N_6027);
or U6588 (N_6588,N_6133,N_6115);
or U6589 (N_6589,N_6046,N_6184);
and U6590 (N_6590,N_6107,N_6244);
xnor U6591 (N_6591,N_6297,N_6064);
nor U6592 (N_6592,N_6053,N_6228);
nor U6593 (N_6593,N_6290,N_6055);
or U6594 (N_6594,N_6206,N_6203);
nor U6595 (N_6595,N_6191,N_6270);
nand U6596 (N_6596,N_6025,N_6262);
nand U6597 (N_6597,N_6022,N_6111);
xnor U6598 (N_6598,N_6120,N_6272);
or U6599 (N_6599,N_6299,N_6071);
and U6600 (N_6600,N_6372,N_6353);
nor U6601 (N_6601,N_6468,N_6497);
xor U6602 (N_6602,N_6474,N_6364);
nand U6603 (N_6603,N_6525,N_6338);
nand U6604 (N_6604,N_6379,N_6383);
and U6605 (N_6605,N_6333,N_6324);
and U6606 (N_6606,N_6439,N_6515);
xnor U6607 (N_6607,N_6530,N_6445);
xor U6608 (N_6608,N_6553,N_6577);
nand U6609 (N_6609,N_6581,N_6342);
xor U6610 (N_6610,N_6412,N_6352);
and U6611 (N_6611,N_6355,N_6340);
nor U6612 (N_6612,N_6398,N_6453);
and U6613 (N_6613,N_6387,N_6572);
or U6614 (N_6614,N_6366,N_6421);
or U6615 (N_6615,N_6509,N_6307);
xor U6616 (N_6616,N_6409,N_6531);
or U6617 (N_6617,N_6332,N_6496);
or U6618 (N_6618,N_6423,N_6305);
and U6619 (N_6619,N_6586,N_6442);
nor U6620 (N_6620,N_6403,N_6417);
or U6621 (N_6621,N_6546,N_6476);
nand U6622 (N_6622,N_6330,N_6571);
or U6623 (N_6623,N_6527,N_6351);
nor U6624 (N_6624,N_6431,N_6323);
nand U6625 (N_6625,N_6511,N_6341);
and U6626 (N_6626,N_6493,N_6494);
or U6627 (N_6627,N_6460,N_6549);
xnor U6628 (N_6628,N_6433,N_6504);
or U6629 (N_6629,N_6430,N_6432);
nor U6630 (N_6630,N_6405,N_6545);
and U6631 (N_6631,N_6344,N_6518);
and U6632 (N_6632,N_6516,N_6590);
xnor U6633 (N_6633,N_6579,N_6346);
xnor U6634 (N_6634,N_6477,N_6552);
nor U6635 (N_6635,N_6569,N_6374);
or U6636 (N_6636,N_6303,N_6555);
or U6637 (N_6637,N_6304,N_6537);
xor U6638 (N_6638,N_6534,N_6401);
xnor U6639 (N_6639,N_6416,N_6559);
and U6640 (N_6640,N_6470,N_6473);
nor U6641 (N_6641,N_6574,N_6359);
nor U6642 (N_6642,N_6487,N_6436);
nor U6643 (N_6643,N_6566,N_6311);
nor U6644 (N_6644,N_6337,N_6319);
nand U6645 (N_6645,N_6402,N_6539);
xor U6646 (N_6646,N_6459,N_6587);
xnor U6647 (N_6647,N_6514,N_6373);
xor U6648 (N_6648,N_6541,N_6316);
nor U6649 (N_6649,N_6513,N_6594);
or U6650 (N_6650,N_6375,N_6321);
nand U6651 (N_6651,N_6326,N_6413);
and U6652 (N_6652,N_6310,N_6302);
nor U6653 (N_6653,N_6596,N_6486);
and U6654 (N_6654,N_6396,N_6523);
nor U6655 (N_6655,N_6595,N_6576);
xnor U6656 (N_6656,N_6535,N_6526);
xor U6657 (N_6657,N_6394,N_6507);
xor U6658 (N_6658,N_6503,N_6519);
nand U6659 (N_6659,N_6455,N_6484);
nand U6660 (N_6660,N_6454,N_6588);
or U6661 (N_6661,N_6415,N_6481);
nand U6662 (N_6662,N_6567,N_6389);
xor U6663 (N_6663,N_6457,N_6306);
nand U6664 (N_6664,N_6528,N_6358);
or U6665 (N_6665,N_6369,N_6472);
nor U6666 (N_6666,N_6501,N_6591);
or U6667 (N_6667,N_6483,N_6585);
or U6668 (N_6668,N_6367,N_6466);
nor U6669 (N_6669,N_6573,N_6510);
and U6670 (N_6670,N_6300,N_6322);
xnor U6671 (N_6671,N_6438,N_6557);
xnor U6672 (N_6672,N_6381,N_6584);
or U6673 (N_6673,N_6400,N_6388);
xor U6674 (N_6674,N_6498,N_6397);
nand U6675 (N_6675,N_6318,N_6325);
and U6676 (N_6676,N_6551,N_6540);
and U6677 (N_6677,N_6478,N_6522);
and U6678 (N_6678,N_6425,N_6391);
and U6679 (N_6679,N_6465,N_6544);
xnor U6680 (N_6680,N_6538,N_6532);
xor U6681 (N_6681,N_6392,N_6570);
or U6682 (N_6682,N_6349,N_6368);
or U6683 (N_6683,N_6565,N_6406);
or U6684 (N_6684,N_6376,N_6314);
nand U6685 (N_6685,N_6428,N_6598);
or U6686 (N_6686,N_6562,N_6464);
and U6687 (N_6687,N_6427,N_6301);
nand U6688 (N_6688,N_6365,N_6410);
nor U6689 (N_6689,N_6578,N_6554);
xor U6690 (N_6690,N_6429,N_6434);
xor U6691 (N_6691,N_6482,N_6480);
or U6692 (N_6692,N_6395,N_6435);
or U6693 (N_6693,N_6593,N_6560);
xnor U6694 (N_6694,N_6450,N_6357);
nor U6695 (N_6695,N_6350,N_6354);
or U6696 (N_6696,N_6536,N_6463);
or U6697 (N_6697,N_6456,N_6471);
xnor U6698 (N_6698,N_6488,N_6317);
nor U6699 (N_6699,N_6561,N_6583);
nor U6700 (N_6700,N_6345,N_6408);
nand U6701 (N_6701,N_6437,N_6424);
nor U6702 (N_6702,N_6356,N_6491);
nand U6703 (N_6703,N_6461,N_6362);
nand U6704 (N_6704,N_6599,N_6575);
or U6705 (N_6705,N_6378,N_6390);
nor U6706 (N_6706,N_6512,N_6309);
and U6707 (N_6707,N_6441,N_6377);
nand U6708 (N_6708,N_6343,N_6458);
or U6709 (N_6709,N_6517,N_6580);
xor U6710 (N_6710,N_6380,N_6521);
nand U6711 (N_6711,N_6543,N_6399);
nor U6712 (N_6712,N_6542,N_6446);
nand U6713 (N_6713,N_6347,N_6370);
xor U6714 (N_6714,N_6589,N_6469);
nor U6715 (N_6715,N_6582,N_6550);
and U6716 (N_6716,N_6462,N_6414);
and U6717 (N_6717,N_6407,N_6385);
and U6718 (N_6718,N_6485,N_6500);
xor U6719 (N_6719,N_6331,N_6564);
xor U6720 (N_6720,N_6426,N_6520);
nor U6721 (N_6721,N_6479,N_6492);
and U6722 (N_6722,N_6419,N_6449);
nand U6723 (N_6723,N_6506,N_6505);
or U6724 (N_6724,N_6336,N_6490);
or U6725 (N_6725,N_6361,N_6444);
nand U6726 (N_6726,N_6334,N_6393);
or U6727 (N_6727,N_6597,N_6440);
or U6728 (N_6728,N_6547,N_6329);
nand U6729 (N_6729,N_6335,N_6327);
or U6730 (N_6730,N_6467,N_6568);
or U6731 (N_6731,N_6495,N_6411);
nor U6732 (N_6732,N_6420,N_6320);
nor U6733 (N_6733,N_6548,N_6524);
xnor U6734 (N_6734,N_6475,N_6348);
xnor U6735 (N_6735,N_6404,N_6360);
or U6736 (N_6736,N_6489,N_6447);
or U6737 (N_6737,N_6384,N_6452);
xnor U6738 (N_6738,N_6382,N_6363);
nand U6739 (N_6739,N_6313,N_6448);
xnor U6740 (N_6740,N_6451,N_6592);
xnor U6741 (N_6741,N_6499,N_6502);
or U6742 (N_6742,N_6508,N_6386);
xor U6743 (N_6743,N_6328,N_6339);
or U6744 (N_6744,N_6418,N_6422);
nand U6745 (N_6745,N_6312,N_6315);
nor U6746 (N_6746,N_6529,N_6533);
or U6747 (N_6747,N_6443,N_6371);
nand U6748 (N_6748,N_6556,N_6563);
and U6749 (N_6749,N_6558,N_6308);
or U6750 (N_6750,N_6439,N_6379);
xnor U6751 (N_6751,N_6320,N_6362);
xor U6752 (N_6752,N_6548,N_6390);
or U6753 (N_6753,N_6340,N_6481);
and U6754 (N_6754,N_6301,N_6506);
xnor U6755 (N_6755,N_6323,N_6527);
nor U6756 (N_6756,N_6486,N_6353);
and U6757 (N_6757,N_6571,N_6471);
nand U6758 (N_6758,N_6539,N_6314);
xor U6759 (N_6759,N_6486,N_6573);
and U6760 (N_6760,N_6503,N_6471);
or U6761 (N_6761,N_6368,N_6559);
or U6762 (N_6762,N_6585,N_6514);
and U6763 (N_6763,N_6549,N_6563);
nor U6764 (N_6764,N_6528,N_6565);
and U6765 (N_6765,N_6489,N_6510);
and U6766 (N_6766,N_6439,N_6581);
nor U6767 (N_6767,N_6412,N_6415);
nor U6768 (N_6768,N_6349,N_6478);
and U6769 (N_6769,N_6319,N_6417);
nand U6770 (N_6770,N_6511,N_6443);
or U6771 (N_6771,N_6424,N_6318);
nand U6772 (N_6772,N_6347,N_6328);
and U6773 (N_6773,N_6415,N_6363);
nand U6774 (N_6774,N_6537,N_6340);
nor U6775 (N_6775,N_6435,N_6397);
or U6776 (N_6776,N_6309,N_6516);
xor U6777 (N_6777,N_6367,N_6573);
xnor U6778 (N_6778,N_6322,N_6566);
nand U6779 (N_6779,N_6511,N_6422);
nor U6780 (N_6780,N_6431,N_6519);
and U6781 (N_6781,N_6583,N_6399);
xor U6782 (N_6782,N_6532,N_6549);
or U6783 (N_6783,N_6488,N_6329);
nor U6784 (N_6784,N_6492,N_6424);
nor U6785 (N_6785,N_6304,N_6350);
or U6786 (N_6786,N_6478,N_6491);
and U6787 (N_6787,N_6448,N_6583);
nand U6788 (N_6788,N_6490,N_6550);
nor U6789 (N_6789,N_6349,N_6400);
or U6790 (N_6790,N_6331,N_6409);
or U6791 (N_6791,N_6400,N_6493);
nor U6792 (N_6792,N_6475,N_6438);
or U6793 (N_6793,N_6480,N_6475);
nor U6794 (N_6794,N_6414,N_6322);
nor U6795 (N_6795,N_6329,N_6307);
and U6796 (N_6796,N_6567,N_6416);
or U6797 (N_6797,N_6452,N_6378);
or U6798 (N_6798,N_6330,N_6543);
nor U6799 (N_6799,N_6511,N_6523);
nand U6800 (N_6800,N_6488,N_6353);
and U6801 (N_6801,N_6515,N_6584);
xnor U6802 (N_6802,N_6317,N_6561);
xnor U6803 (N_6803,N_6510,N_6380);
nand U6804 (N_6804,N_6350,N_6538);
nand U6805 (N_6805,N_6318,N_6544);
xor U6806 (N_6806,N_6357,N_6400);
nand U6807 (N_6807,N_6383,N_6512);
and U6808 (N_6808,N_6486,N_6390);
or U6809 (N_6809,N_6491,N_6535);
or U6810 (N_6810,N_6420,N_6449);
nand U6811 (N_6811,N_6424,N_6407);
and U6812 (N_6812,N_6552,N_6445);
nor U6813 (N_6813,N_6345,N_6570);
xnor U6814 (N_6814,N_6529,N_6406);
nand U6815 (N_6815,N_6569,N_6571);
nand U6816 (N_6816,N_6373,N_6374);
and U6817 (N_6817,N_6498,N_6324);
nor U6818 (N_6818,N_6492,N_6485);
and U6819 (N_6819,N_6550,N_6430);
nand U6820 (N_6820,N_6561,N_6429);
or U6821 (N_6821,N_6540,N_6331);
xnor U6822 (N_6822,N_6301,N_6315);
nand U6823 (N_6823,N_6366,N_6568);
and U6824 (N_6824,N_6396,N_6351);
xor U6825 (N_6825,N_6591,N_6416);
or U6826 (N_6826,N_6553,N_6567);
xnor U6827 (N_6827,N_6552,N_6460);
nand U6828 (N_6828,N_6394,N_6367);
or U6829 (N_6829,N_6527,N_6584);
xnor U6830 (N_6830,N_6517,N_6523);
or U6831 (N_6831,N_6474,N_6314);
and U6832 (N_6832,N_6386,N_6402);
xor U6833 (N_6833,N_6311,N_6357);
nand U6834 (N_6834,N_6578,N_6401);
nor U6835 (N_6835,N_6568,N_6307);
or U6836 (N_6836,N_6420,N_6514);
xnor U6837 (N_6837,N_6555,N_6395);
and U6838 (N_6838,N_6324,N_6365);
nor U6839 (N_6839,N_6451,N_6515);
and U6840 (N_6840,N_6438,N_6446);
or U6841 (N_6841,N_6537,N_6528);
xnor U6842 (N_6842,N_6395,N_6389);
nand U6843 (N_6843,N_6318,N_6435);
or U6844 (N_6844,N_6587,N_6421);
xnor U6845 (N_6845,N_6539,N_6546);
and U6846 (N_6846,N_6546,N_6580);
xor U6847 (N_6847,N_6414,N_6439);
nand U6848 (N_6848,N_6484,N_6594);
xnor U6849 (N_6849,N_6565,N_6442);
nand U6850 (N_6850,N_6514,N_6562);
or U6851 (N_6851,N_6323,N_6579);
and U6852 (N_6852,N_6479,N_6469);
xor U6853 (N_6853,N_6419,N_6496);
and U6854 (N_6854,N_6572,N_6369);
nor U6855 (N_6855,N_6569,N_6398);
nor U6856 (N_6856,N_6410,N_6548);
xnor U6857 (N_6857,N_6317,N_6430);
xnor U6858 (N_6858,N_6311,N_6483);
or U6859 (N_6859,N_6377,N_6447);
nor U6860 (N_6860,N_6509,N_6360);
xor U6861 (N_6861,N_6338,N_6585);
or U6862 (N_6862,N_6348,N_6588);
xnor U6863 (N_6863,N_6517,N_6539);
xnor U6864 (N_6864,N_6505,N_6571);
xnor U6865 (N_6865,N_6587,N_6402);
nor U6866 (N_6866,N_6529,N_6388);
nand U6867 (N_6867,N_6452,N_6401);
nand U6868 (N_6868,N_6464,N_6576);
nand U6869 (N_6869,N_6576,N_6448);
nand U6870 (N_6870,N_6355,N_6302);
nand U6871 (N_6871,N_6575,N_6325);
and U6872 (N_6872,N_6483,N_6595);
xnor U6873 (N_6873,N_6437,N_6588);
xor U6874 (N_6874,N_6580,N_6445);
nand U6875 (N_6875,N_6446,N_6457);
xnor U6876 (N_6876,N_6398,N_6509);
and U6877 (N_6877,N_6394,N_6504);
and U6878 (N_6878,N_6404,N_6429);
xnor U6879 (N_6879,N_6346,N_6382);
or U6880 (N_6880,N_6362,N_6556);
or U6881 (N_6881,N_6571,N_6591);
or U6882 (N_6882,N_6560,N_6548);
nor U6883 (N_6883,N_6573,N_6428);
xor U6884 (N_6884,N_6571,N_6312);
xnor U6885 (N_6885,N_6384,N_6369);
and U6886 (N_6886,N_6431,N_6367);
nand U6887 (N_6887,N_6390,N_6558);
nand U6888 (N_6888,N_6345,N_6491);
nor U6889 (N_6889,N_6463,N_6419);
or U6890 (N_6890,N_6392,N_6443);
nor U6891 (N_6891,N_6301,N_6351);
and U6892 (N_6892,N_6306,N_6564);
xnor U6893 (N_6893,N_6530,N_6443);
xnor U6894 (N_6894,N_6507,N_6516);
or U6895 (N_6895,N_6501,N_6573);
nand U6896 (N_6896,N_6381,N_6406);
xnor U6897 (N_6897,N_6580,N_6586);
nor U6898 (N_6898,N_6350,N_6486);
nor U6899 (N_6899,N_6389,N_6364);
or U6900 (N_6900,N_6746,N_6744);
xnor U6901 (N_6901,N_6876,N_6621);
nand U6902 (N_6902,N_6884,N_6847);
nand U6903 (N_6903,N_6871,N_6687);
or U6904 (N_6904,N_6637,N_6769);
nor U6905 (N_6905,N_6670,N_6872);
nand U6906 (N_6906,N_6700,N_6776);
and U6907 (N_6907,N_6681,N_6679);
nor U6908 (N_6908,N_6719,N_6866);
and U6909 (N_6909,N_6780,N_6655);
xor U6910 (N_6910,N_6628,N_6813);
xor U6911 (N_6911,N_6882,N_6678);
and U6912 (N_6912,N_6873,N_6717);
or U6913 (N_6913,N_6755,N_6714);
or U6914 (N_6914,N_6781,N_6630);
nor U6915 (N_6915,N_6836,N_6777);
or U6916 (N_6916,N_6839,N_6688);
xnor U6917 (N_6917,N_6863,N_6737);
or U6918 (N_6918,N_6821,N_6827);
or U6919 (N_6919,N_6853,N_6680);
nand U6920 (N_6920,N_6823,N_6773);
and U6921 (N_6921,N_6765,N_6715);
nand U6922 (N_6922,N_6728,N_6788);
xor U6923 (N_6923,N_6733,N_6812);
and U6924 (N_6924,N_6638,N_6881);
nor U6925 (N_6925,N_6686,N_6610);
and U6926 (N_6926,N_6811,N_6726);
nand U6927 (N_6927,N_6732,N_6694);
xnor U6928 (N_6928,N_6880,N_6609);
and U6929 (N_6929,N_6622,N_6674);
nand U6930 (N_6930,N_6656,N_6711);
xnor U6931 (N_6931,N_6826,N_6707);
or U6932 (N_6932,N_6627,N_6838);
nand U6933 (N_6933,N_6867,N_6830);
nand U6934 (N_6934,N_6607,N_6846);
or U6935 (N_6935,N_6774,N_6874);
xnor U6936 (N_6936,N_6664,N_6742);
xnor U6937 (N_6937,N_6759,N_6785);
or U6938 (N_6938,N_6615,N_6659);
and U6939 (N_6939,N_6756,N_6752);
xnor U6940 (N_6940,N_6894,N_6779);
xnor U6941 (N_6941,N_6851,N_6825);
xor U6942 (N_6942,N_6635,N_6648);
or U6943 (N_6943,N_6891,N_6834);
and U6944 (N_6944,N_6745,N_6602);
nor U6945 (N_6945,N_6848,N_6682);
xnor U6946 (N_6946,N_6632,N_6662);
nand U6947 (N_6947,N_6721,N_6605);
xor U6948 (N_6948,N_6870,N_6684);
nor U6949 (N_6949,N_6604,N_6722);
nand U6950 (N_6950,N_6748,N_6818);
and U6951 (N_6951,N_6723,N_6819);
nor U6952 (N_6952,N_6676,N_6783);
and U6953 (N_6953,N_6766,N_6690);
nand U6954 (N_6954,N_6730,N_6668);
nand U6955 (N_6955,N_6801,N_6683);
or U6956 (N_6956,N_6640,N_6718);
and U6957 (N_6957,N_6789,N_6887);
or U6958 (N_6958,N_6835,N_6852);
nor U6959 (N_6959,N_6810,N_6753);
and U6960 (N_6960,N_6631,N_6747);
nor U6961 (N_6961,N_6868,N_6832);
nand U6962 (N_6962,N_6724,N_6639);
xnor U6963 (N_6963,N_6691,N_6771);
nor U6964 (N_6964,N_6654,N_6661);
and U6965 (N_6965,N_6800,N_6650);
nor U6966 (N_6966,N_6896,N_6701);
or U6967 (N_6967,N_6697,N_6725);
or U6968 (N_6968,N_6603,N_6828);
and U6969 (N_6969,N_6854,N_6849);
nor U6970 (N_6970,N_6862,N_6763);
or U6971 (N_6971,N_6820,N_6841);
xor U6972 (N_6972,N_6762,N_6815);
nor U6973 (N_6973,N_6734,N_6888);
nor U6974 (N_6974,N_6877,N_6875);
and U6975 (N_6975,N_6806,N_6642);
and U6976 (N_6976,N_6646,N_6614);
nand U6977 (N_6977,N_6667,N_6750);
or U6978 (N_6978,N_6705,N_6751);
xor U6979 (N_6979,N_6669,N_6816);
and U6980 (N_6980,N_6833,N_6651);
nand U6981 (N_6981,N_6786,N_6802);
and U6982 (N_6982,N_6652,N_6814);
and U6983 (N_6983,N_6695,N_6768);
and U6984 (N_6984,N_6807,N_6885);
and U6985 (N_6985,N_6658,N_6624);
nor U6986 (N_6986,N_6796,N_6649);
xor U6987 (N_6987,N_6665,N_6611);
xor U6988 (N_6988,N_6808,N_6601);
and U6989 (N_6989,N_6675,N_6699);
xor U6990 (N_6990,N_6754,N_6720);
nor U6991 (N_6991,N_6764,N_6660);
nand U6992 (N_6992,N_6770,N_6727);
or U6993 (N_6993,N_6729,N_6898);
nand U6994 (N_6994,N_6893,N_6619);
nand U6995 (N_6995,N_6889,N_6616);
nor U6996 (N_6996,N_6878,N_6817);
or U6997 (N_6997,N_6620,N_6842);
or U6998 (N_6998,N_6738,N_6865);
and U6999 (N_6999,N_6740,N_6743);
or U7000 (N_7000,N_6799,N_6673);
nand U7001 (N_7001,N_6600,N_6677);
or U7002 (N_7002,N_6689,N_6634);
nand U7003 (N_7003,N_6804,N_6775);
xnor U7004 (N_7004,N_6837,N_6692);
xor U7005 (N_7005,N_6716,N_6757);
or U7006 (N_7006,N_6794,N_6787);
nor U7007 (N_7007,N_6805,N_6663);
and U7008 (N_7008,N_6767,N_6824);
nand U7009 (N_7009,N_6861,N_6672);
or U7010 (N_7010,N_6803,N_6749);
and U7011 (N_7011,N_6731,N_6844);
nor U7012 (N_7012,N_6895,N_6736);
and U7013 (N_7013,N_6644,N_6706);
and U7014 (N_7014,N_6708,N_6758);
and U7015 (N_7015,N_6840,N_6657);
or U7016 (N_7016,N_6857,N_6831);
xor U7017 (N_7017,N_6625,N_6886);
xor U7018 (N_7018,N_6859,N_6892);
xor U7019 (N_7019,N_6829,N_6879);
or U7020 (N_7020,N_6704,N_6698);
nor U7021 (N_7021,N_6890,N_6685);
or U7022 (N_7022,N_6822,N_6629);
nor U7023 (N_7023,N_6739,N_6703);
nand U7024 (N_7024,N_6897,N_6845);
and U7025 (N_7025,N_6606,N_6671);
or U7026 (N_7026,N_6693,N_6856);
or U7027 (N_7027,N_6696,N_6850);
xnor U7028 (N_7028,N_6641,N_6843);
or U7029 (N_7029,N_6784,N_6761);
nand U7030 (N_7030,N_6864,N_6791);
and U7031 (N_7031,N_6643,N_6778);
and U7032 (N_7032,N_6809,N_6798);
nor U7033 (N_7033,N_6860,N_6617);
nor U7034 (N_7034,N_6772,N_6782);
nor U7035 (N_7035,N_6712,N_6702);
xor U7036 (N_7036,N_6735,N_6612);
xnor U7037 (N_7037,N_6636,N_6709);
nand U7038 (N_7038,N_6760,N_6710);
xnor U7039 (N_7039,N_6858,N_6899);
or U7040 (N_7040,N_6713,N_6633);
or U7041 (N_7041,N_6608,N_6645);
nor U7042 (N_7042,N_6790,N_6613);
nand U7043 (N_7043,N_6855,N_6792);
or U7044 (N_7044,N_6793,N_6741);
nand U7045 (N_7045,N_6647,N_6618);
nand U7046 (N_7046,N_6869,N_6666);
nand U7047 (N_7047,N_6623,N_6797);
nand U7048 (N_7048,N_6626,N_6653);
nand U7049 (N_7049,N_6883,N_6795);
nand U7050 (N_7050,N_6820,N_6884);
or U7051 (N_7051,N_6829,N_6763);
nor U7052 (N_7052,N_6845,N_6662);
nand U7053 (N_7053,N_6807,N_6802);
xnor U7054 (N_7054,N_6628,N_6705);
and U7055 (N_7055,N_6671,N_6736);
nor U7056 (N_7056,N_6701,N_6729);
xnor U7057 (N_7057,N_6781,N_6612);
or U7058 (N_7058,N_6623,N_6672);
nor U7059 (N_7059,N_6660,N_6678);
nand U7060 (N_7060,N_6850,N_6706);
nand U7061 (N_7061,N_6711,N_6765);
or U7062 (N_7062,N_6600,N_6657);
and U7063 (N_7063,N_6741,N_6872);
xor U7064 (N_7064,N_6793,N_6731);
nand U7065 (N_7065,N_6801,N_6718);
xor U7066 (N_7066,N_6671,N_6788);
and U7067 (N_7067,N_6650,N_6710);
nor U7068 (N_7068,N_6732,N_6781);
and U7069 (N_7069,N_6662,N_6655);
nand U7070 (N_7070,N_6861,N_6647);
nand U7071 (N_7071,N_6838,N_6625);
xor U7072 (N_7072,N_6895,N_6614);
or U7073 (N_7073,N_6689,N_6721);
nor U7074 (N_7074,N_6736,N_6720);
and U7075 (N_7075,N_6895,N_6742);
nand U7076 (N_7076,N_6812,N_6625);
and U7077 (N_7077,N_6605,N_6686);
xor U7078 (N_7078,N_6605,N_6746);
nand U7079 (N_7079,N_6857,N_6671);
or U7080 (N_7080,N_6627,N_6741);
xnor U7081 (N_7081,N_6815,N_6744);
xor U7082 (N_7082,N_6809,N_6896);
or U7083 (N_7083,N_6714,N_6625);
nor U7084 (N_7084,N_6602,N_6795);
nand U7085 (N_7085,N_6737,N_6639);
or U7086 (N_7086,N_6602,N_6619);
and U7087 (N_7087,N_6702,N_6728);
or U7088 (N_7088,N_6704,N_6846);
and U7089 (N_7089,N_6866,N_6892);
or U7090 (N_7090,N_6883,N_6611);
or U7091 (N_7091,N_6647,N_6609);
xnor U7092 (N_7092,N_6672,N_6847);
or U7093 (N_7093,N_6796,N_6627);
and U7094 (N_7094,N_6645,N_6808);
nor U7095 (N_7095,N_6863,N_6615);
xor U7096 (N_7096,N_6854,N_6893);
nand U7097 (N_7097,N_6697,N_6862);
and U7098 (N_7098,N_6728,N_6818);
nand U7099 (N_7099,N_6898,N_6814);
nand U7100 (N_7100,N_6754,N_6895);
or U7101 (N_7101,N_6671,N_6732);
xor U7102 (N_7102,N_6854,N_6773);
xnor U7103 (N_7103,N_6884,N_6896);
nor U7104 (N_7104,N_6887,N_6671);
nand U7105 (N_7105,N_6789,N_6707);
xor U7106 (N_7106,N_6697,N_6836);
and U7107 (N_7107,N_6604,N_6757);
and U7108 (N_7108,N_6712,N_6682);
nand U7109 (N_7109,N_6633,N_6842);
and U7110 (N_7110,N_6647,N_6889);
nor U7111 (N_7111,N_6760,N_6719);
nand U7112 (N_7112,N_6687,N_6787);
or U7113 (N_7113,N_6737,N_6717);
or U7114 (N_7114,N_6859,N_6871);
or U7115 (N_7115,N_6669,N_6744);
nor U7116 (N_7116,N_6696,N_6843);
and U7117 (N_7117,N_6669,N_6827);
or U7118 (N_7118,N_6665,N_6754);
nor U7119 (N_7119,N_6863,N_6857);
xnor U7120 (N_7120,N_6772,N_6617);
or U7121 (N_7121,N_6632,N_6608);
xor U7122 (N_7122,N_6833,N_6650);
nand U7123 (N_7123,N_6802,N_6608);
xnor U7124 (N_7124,N_6646,N_6752);
xnor U7125 (N_7125,N_6720,N_6833);
or U7126 (N_7126,N_6866,N_6647);
nor U7127 (N_7127,N_6600,N_6750);
nand U7128 (N_7128,N_6646,N_6790);
nand U7129 (N_7129,N_6662,N_6653);
xnor U7130 (N_7130,N_6633,N_6698);
nand U7131 (N_7131,N_6749,N_6673);
xnor U7132 (N_7132,N_6720,N_6876);
xor U7133 (N_7133,N_6721,N_6820);
nand U7134 (N_7134,N_6892,N_6781);
nor U7135 (N_7135,N_6616,N_6649);
xnor U7136 (N_7136,N_6678,N_6879);
nor U7137 (N_7137,N_6745,N_6616);
xor U7138 (N_7138,N_6618,N_6753);
and U7139 (N_7139,N_6883,N_6658);
nand U7140 (N_7140,N_6784,N_6719);
xor U7141 (N_7141,N_6846,N_6683);
nor U7142 (N_7142,N_6678,N_6711);
xnor U7143 (N_7143,N_6789,N_6600);
xnor U7144 (N_7144,N_6617,N_6653);
and U7145 (N_7145,N_6756,N_6866);
nor U7146 (N_7146,N_6700,N_6647);
or U7147 (N_7147,N_6606,N_6659);
xor U7148 (N_7148,N_6892,N_6852);
nand U7149 (N_7149,N_6891,N_6853);
xnor U7150 (N_7150,N_6899,N_6845);
xnor U7151 (N_7151,N_6691,N_6628);
nor U7152 (N_7152,N_6607,N_6824);
nor U7153 (N_7153,N_6699,N_6804);
nor U7154 (N_7154,N_6787,N_6619);
xnor U7155 (N_7155,N_6720,N_6889);
xnor U7156 (N_7156,N_6712,N_6798);
nor U7157 (N_7157,N_6770,N_6838);
xnor U7158 (N_7158,N_6623,N_6723);
nand U7159 (N_7159,N_6779,N_6728);
or U7160 (N_7160,N_6885,N_6646);
nand U7161 (N_7161,N_6886,N_6770);
and U7162 (N_7162,N_6787,N_6749);
nand U7163 (N_7163,N_6850,N_6851);
and U7164 (N_7164,N_6780,N_6751);
nand U7165 (N_7165,N_6646,N_6797);
xor U7166 (N_7166,N_6609,N_6886);
nand U7167 (N_7167,N_6723,N_6651);
nand U7168 (N_7168,N_6849,N_6653);
or U7169 (N_7169,N_6707,N_6604);
or U7170 (N_7170,N_6815,N_6839);
and U7171 (N_7171,N_6695,N_6711);
and U7172 (N_7172,N_6613,N_6616);
and U7173 (N_7173,N_6823,N_6755);
xor U7174 (N_7174,N_6880,N_6769);
nand U7175 (N_7175,N_6840,N_6889);
nand U7176 (N_7176,N_6615,N_6848);
nand U7177 (N_7177,N_6816,N_6679);
nand U7178 (N_7178,N_6818,N_6601);
and U7179 (N_7179,N_6688,N_6796);
nand U7180 (N_7180,N_6603,N_6635);
nand U7181 (N_7181,N_6687,N_6796);
and U7182 (N_7182,N_6688,N_6739);
nand U7183 (N_7183,N_6832,N_6822);
and U7184 (N_7184,N_6637,N_6877);
xor U7185 (N_7185,N_6644,N_6673);
and U7186 (N_7186,N_6644,N_6696);
nand U7187 (N_7187,N_6834,N_6610);
and U7188 (N_7188,N_6861,N_6873);
nor U7189 (N_7189,N_6629,N_6772);
nand U7190 (N_7190,N_6829,N_6693);
or U7191 (N_7191,N_6646,N_6607);
and U7192 (N_7192,N_6816,N_6706);
nand U7193 (N_7193,N_6677,N_6762);
nand U7194 (N_7194,N_6619,N_6865);
and U7195 (N_7195,N_6814,N_6692);
and U7196 (N_7196,N_6600,N_6697);
or U7197 (N_7197,N_6687,N_6669);
nor U7198 (N_7198,N_6751,N_6708);
xnor U7199 (N_7199,N_6886,N_6663);
or U7200 (N_7200,N_7147,N_7101);
and U7201 (N_7201,N_7060,N_7148);
nor U7202 (N_7202,N_7196,N_7019);
nand U7203 (N_7203,N_6970,N_7023);
and U7204 (N_7204,N_7142,N_7004);
nand U7205 (N_7205,N_7176,N_7159);
nand U7206 (N_7206,N_7099,N_6940);
xor U7207 (N_7207,N_7040,N_7098);
xnor U7208 (N_7208,N_7097,N_7030);
nand U7209 (N_7209,N_7191,N_7050);
nor U7210 (N_7210,N_7143,N_7003);
or U7211 (N_7211,N_7039,N_6994);
nand U7212 (N_7212,N_6978,N_7192);
or U7213 (N_7213,N_7083,N_6922);
and U7214 (N_7214,N_6923,N_7120);
xnor U7215 (N_7215,N_7032,N_7199);
nand U7216 (N_7216,N_7072,N_6915);
and U7217 (N_7217,N_7088,N_7153);
and U7218 (N_7218,N_7074,N_7036);
and U7219 (N_7219,N_7131,N_7041);
or U7220 (N_7220,N_6980,N_7085);
nor U7221 (N_7221,N_7010,N_6981);
and U7222 (N_7222,N_7089,N_6901);
nand U7223 (N_7223,N_7095,N_7157);
and U7224 (N_7224,N_7110,N_7035);
nor U7225 (N_7225,N_7045,N_6920);
nand U7226 (N_7226,N_6931,N_7141);
nand U7227 (N_7227,N_7184,N_7130);
nor U7228 (N_7228,N_7049,N_7092);
or U7229 (N_7229,N_6930,N_7014);
nor U7230 (N_7230,N_7154,N_7042);
or U7231 (N_7231,N_6987,N_7077);
and U7232 (N_7232,N_7044,N_7053);
nand U7233 (N_7233,N_6917,N_7047);
xnor U7234 (N_7234,N_7028,N_7122);
nand U7235 (N_7235,N_7128,N_6996);
nand U7236 (N_7236,N_6948,N_7001);
nand U7237 (N_7237,N_6965,N_7057);
xnor U7238 (N_7238,N_7055,N_6961);
nor U7239 (N_7239,N_7013,N_7084);
or U7240 (N_7240,N_7174,N_6986);
nand U7241 (N_7241,N_7158,N_6903);
nor U7242 (N_7242,N_7114,N_7104);
and U7243 (N_7243,N_7046,N_6997);
nor U7244 (N_7244,N_7108,N_6902);
nand U7245 (N_7245,N_6914,N_6910);
nor U7246 (N_7246,N_7024,N_7166);
and U7247 (N_7247,N_7165,N_6949);
nand U7248 (N_7248,N_7155,N_7070);
nand U7249 (N_7249,N_6945,N_7094);
or U7250 (N_7250,N_7167,N_7116);
or U7251 (N_7251,N_7109,N_7056);
or U7252 (N_7252,N_6905,N_7115);
nor U7253 (N_7253,N_6943,N_7194);
and U7254 (N_7254,N_7171,N_6936);
nand U7255 (N_7255,N_6968,N_6937);
nand U7256 (N_7256,N_6959,N_7016);
nor U7257 (N_7257,N_7179,N_7182);
nor U7258 (N_7258,N_6951,N_6927);
and U7259 (N_7259,N_7076,N_7107);
xor U7260 (N_7260,N_7058,N_7091);
nor U7261 (N_7261,N_7172,N_7123);
xor U7262 (N_7262,N_7081,N_6999);
and U7263 (N_7263,N_7135,N_6918);
xor U7264 (N_7264,N_7008,N_6946);
nand U7265 (N_7265,N_7164,N_7082);
or U7266 (N_7266,N_7038,N_6900);
nand U7267 (N_7267,N_6958,N_7073);
xor U7268 (N_7268,N_7161,N_7173);
xnor U7269 (N_7269,N_7133,N_7065);
xnor U7270 (N_7270,N_7071,N_7087);
and U7271 (N_7271,N_6964,N_6908);
nand U7272 (N_7272,N_7005,N_7193);
or U7273 (N_7273,N_6911,N_7129);
nand U7274 (N_7274,N_6977,N_7051);
and U7275 (N_7275,N_7197,N_6957);
and U7276 (N_7276,N_6982,N_6983);
or U7277 (N_7277,N_6990,N_7183);
nand U7278 (N_7278,N_7127,N_6942);
nor U7279 (N_7279,N_6976,N_7150);
nand U7280 (N_7280,N_7029,N_7170);
and U7281 (N_7281,N_7119,N_6933);
nand U7282 (N_7282,N_6919,N_7124);
xnor U7283 (N_7283,N_6984,N_7079);
nor U7284 (N_7284,N_7054,N_6925);
xor U7285 (N_7285,N_7009,N_7113);
and U7286 (N_7286,N_7111,N_6993);
nand U7287 (N_7287,N_7187,N_7006);
xnor U7288 (N_7288,N_6909,N_7067);
nor U7289 (N_7289,N_7156,N_7132);
nand U7290 (N_7290,N_7169,N_6995);
nand U7291 (N_7291,N_6912,N_7002);
nand U7292 (N_7292,N_7027,N_6952);
xor U7293 (N_7293,N_7017,N_7080);
or U7294 (N_7294,N_6974,N_7175);
and U7295 (N_7295,N_6991,N_7061);
nand U7296 (N_7296,N_7064,N_6992);
and U7297 (N_7297,N_7007,N_7100);
and U7298 (N_7298,N_6955,N_7198);
nor U7299 (N_7299,N_7031,N_7140);
xor U7300 (N_7300,N_7086,N_6926);
nor U7301 (N_7301,N_6929,N_7068);
xnor U7302 (N_7302,N_7152,N_7063);
nor U7303 (N_7303,N_6921,N_7103);
nand U7304 (N_7304,N_7093,N_6998);
nand U7305 (N_7305,N_7048,N_7102);
xor U7306 (N_7306,N_6939,N_7181);
nand U7307 (N_7307,N_6966,N_6934);
xor U7308 (N_7308,N_6985,N_7022);
and U7309 (N_7309,N_7020,N_6944);
and U7310 (N_7310,N_6950,N_6907);
nor U7311 (N_7311,N_6932,N_6972);
nor U7312 (N_7312,N_7000,N_6938);
and U7313 (N_7313,N_7190,N_7075);
nand U7314 (N_7314,N_6904,N_7138);
xor U7315 (N_7315,N_7011,N_7043);
and U7316 (N_7316,N_6954,N_7034);
and U7317 (N_7317,N_6962,N_7118);
nand U7318 (N_7318,N_7021,N_7018);
or U7319 (N_7319,N_7144,N_6971);
nand U7320 (N_7320,N_7117,N_6973);
xnor U7321 (N_7321,N_7139,N_7025);
xor U7322 (N_7322,N_7136,N_7069);
nor U7323 (N_7323,N_7059,N_6969);
nor U7324 (N_7324,N_7186,N_7121);
or U7325 (N_7325,N_7078,N_7146);
or U7326 (N_7326,N_7015,N_7106);
nor U7327 (N_7327,N_7096,N_7178);
nor U7328 (N_7328,N_6975,N_7149);
or U7329 (N_7329,N_7195,N_7177);
or U7330 (N_7330,N_6953,N_6913);
and U7331 (N_7331,N_7090,N_7137);
nand U7332 (N_7332,N_6906,N_6935);
nor U7333 (N_7333,N_7033,N_7160);
and U7334 (N_7334,N_6916,N_6979);
and U7335 (N_7335,N_7189,N_7105);
or U7336 (N_7336,N_7188,N_6956);
xnor U7337 (N_7337,N_6967,N_7180);
xor U7338 (N_7338,N_6928,N_7037);
nand U7339 (N_7339,N_7168,N_7185);
or U7340 (N_7340,N_7112,N_7066);
and U7341 (N_7341,N_6988,N_6947);
or U7342 (N_7342,N_6989,N_7126);
and U7343 (N_7343,N_7062,N_7052);
or U7344 (N_7344,N_7134,N_7125);
and U7345 (N_7345,N_7145,N_6941);
or U7346 (N_7346,N_6963,N_7163);
nand U7347 (N_7347,N_7162,N_7151);
xor U7348 (N_7348,N_7026,N_6960);
or U7349 (N_7349,N_6924,N_7012);
nor U7350 (N_7350,N_6940,N_6936);
or U7351 (N_7351,N_6990,N_7069);
and U7352 (N_7352,N_7010,N_7194);
and U7353 (N_7353,N_6945,N_6901);
or U7354 (N_7354,N_7154,N_7160);
and U7355 (N_7355,N_7114,N_7019);
nand U7356 (N_7356,N_7152,N_7059);
or U7357 (N_7357,N_7117,N_7128);
and U7358 (N_7358,N_7146,N_6936);
and U7359 (N_7359,N_7160,N_6941);
xnor U7360 (N_7360,N_6926,N_7116);
and U7361 (N_7361,N_7031,N_7088);
and U7362 (N_7362,N_6989,N_7036);
nand U7363 (N_7363,N_7139,N_6986);
xor U7364 (N_7364,N_7064,N_7054);
nor U7365 (N_7365,N_7142,N_6933);
and U7366 (N_7366,N_6982,N_7183);
nand U7367 (N_7367,N_7061,N_7062);
or U7368 (N_7368,N_7141,N_7166);
nand U7369 (N_7369,N_7100,N_6966);
xor U7370 (N_7370,N_6919,N_7006);
and U7371 (N_7371,N_7010,N_7164);
and U7372 (N_7372,N_7081,N_7059);
or U7373 (N_7373,N_6997,N_6932);
nand U7374 (N_7374,N_6956,N_7191);
nand U7375 (N_7375,N_7024,N_7058);
or U7376 (N_7376,N_7129,N_7082);
and U7377 (N_7377,N_6995,N_7126);
nor U7378 (N_7378,N_7002,N_7036);
xor U7379 (N_7379,N_6999,N_7103);
nor U7380 (N_7380,N_6966,N_7135);
nand U7381 (N_7381,N_7007,N_6948);
nor U7382 (N_7382,N_6999,N_6917);
and U7383 (N_7383,N_6974,N_6986);
and U7384 (N_7384,N_6927,N_7106);
nor U7385 (N_7385,N_7144,N_6935);
and U7386 (N_7386,N_7095,N_7098);
and U7387 (N_7387,N_6960,N_7048);
and U7388 (N_7388,N_7161,N_6959);
or U7389 (N_7389,N_7092,N_7094);
or U7390 (N_7390,N_7080,N_7028);
and U7391 (N_7391,N_7108,N_7154);
nand U7392 (N_7392,N_7100,N_7152);
xor U7393 (N_7393,N_6926,N_7173);
or U7394 (N_7394,N_6966,N_7116);
xor U7395 (N_7395,N_7066,N_7170);
and U7396 (N_7396,N_6949,N_6900);
nand U7397 (N_7397,N_7175,N_7016);
and U7398 (N_7398,N_7016,N_7012);
nor U7399 (N_7399,N_6980,N_7063);
nand U7400 (N_7400,N_7089,N_7176);
nor U7401 (N_7401,N_7126,N_7100);
nor U7402 (N_7402,N_7157,N_7119);
xor U7403 (N_7403,N_7149,N_6995);
nor U7404 (N_7404,N_6958,N_7121);
nor U7405 (N_7405,N_7118,N_7105);
xor U7406 (N_7406,N_7053,N_7045);
xor U7407 (N_7407,N_6903,N_7172);
or U7408 (N_7408,N_6979,N_7079);
xnor U7409 (N_7409,N_6904,N_6977);
or U7410 (N_7410,N_7014,N_6917);
or U7411 (N_7411,N_7198,N_7123);
nor U7412 (N_7412,N_7198,N_6972);
or U7413 (N_7413,N_7115,N_7103);
nand U7414 (N_7414,N_7101,N_7082);
nand U7415 (N_7415,N_6964,N_6963);
nor U7416 (N_7416,N_7104,N_7161);
nand U7417 (N_7417,N_6903,N_7104);
nor U7418 (N_7418,N_6966,N_6908);
xnor U7419 (N_7419,N_7173,N_7053);
nor U7420 (N_7420,N_6909,N_6927);
xnor U7421 (N_7421,N_6919,N_7148);
nand U7422 (N_7422,N_7134,N_7017);
xnor U7423 (N_7423,N_7179,N_7009);
xor U7424 (N_7424,N_7036,N_6931);
or U7425 (N_7425,N_7018,N_6920);
nand U7426 (N_7426,N_7076,N_7046);
and U7427 (N_7427,N_7121,N_7176);
nor U7428 (N_7428,N_6918,N_7066);
and U7429 (N_7429,N_7013,N_7137);
nor U7430 (N_7430,N_7063,N_7160);
nand U7431 (N_7431,N_6914,N_6956);
nand U7432 (N_7432,N_7128,N_7013);
or U7433 (N_7433,N_7190,N_7029);
or U7434 (N_7434,N_7072,N_7071);
nand U7435 (N_7435,N_7081,N_7002);
nand U7436 (N_7436,N_6953,N_7055);
nor U7437 (N_7437,N_7154,N_6974);
nor U7438 (N_7438,N_6972,N_7183);
nor U7439 (N_7439,N_7125,N_7170);
or U7440 (N_7440,N_7059,N_6992);
xor U7441 (N_7441,N_7062,N_6918);
nor U7442 (N_7442,N_6985,N_6911);
xnor U7443 (N_7443,N_7060,N_6997);
and U7444 (N_7444,N_6912,N_6983);
nand U7445 (N_7445,N_6924,N_7091);
nor U7446 (N_7446,N_6987,N_7051);
nand U7447 (N_7447,N_7191,N_7098);
and U7448 (N_7448,N_7148,N_7109);
and U7449 (N_7449,N_7057,N_6953);
xor U7450 (N_7450,N_7174,N_7021);
nor U7451 (N_7451,N_7067,N_7170);
nand U7452 (N_7452,N_7073,N_6942);
nand U7453 (N_7453,N_7129,N_7001);
xor U7454 (N_7454,N_7186,N_6990);
or U7455 (N_7455,N_7188,N_6986);
xor U7456 (N_7456,N_7098,N_7084);
nor U7457 (N_7457,N_7003,N_6963);
or U7458 (N_7458,N_7155,N_6902);
xnor U7459 (N_7459,N_6983,N_7135);
and U7460 (N_7460,N_6975,N_7191);
xor U7461 (N_7461,N_7020,N_7118);
nor U7462 (N_7462,N_7085,N_7010);
xor U7463 (N_7463,N_7148,N_7184);
xor U7464 (N_7464,N_6926,N_6983);
xnor U7465 (N_7465,N_7111,N_7153);
nor U7466 (N_7466,N_7158,N_7077);
nand U7467 (N_7467,N_7116,N_7168);
or U7468 (N_7468,N_6955,N_6945);
nand U7469 (N_7469,N_7008,N_6912);
xor U7470 (N_7470,N_7060,N_7113);
xor U7471 (N_7471,N_7127,N_7020);
and U7472 (N_7472,N_7043,N_7189);
xnor U7473 (N_7473,N_7053,N_6908);
and U7474 (N_7474,N_7131,N_7090);
nor U7475 (N_7475,N_7148,N_7138);
xnor U7476 (N_7476,N_7133,N_6901);
xnor U7477 (N_7477,N_7183,N_7062);
xnor U7478 (N_7478,N_6945,N_7060);
nor U7479 (N_7479,N_6946,N_7129);
xnor U7480 (N_7480,N_6902,N_7006);
and U7481 (N_7481,N_6991,N_7093);
and U7482 (N_7482,N_7023,N_6907);
or U7483 (N_7483,N_7143,N_6996);
or U7484 (N_7484,N_7047,N_6956);
or U7485 (N_7485,N_7190,N_7194);
xnor U7486 (N_7486,N_6962,N_7026);
and U7487 (N_7487,N_7180,N_7044);
or U7488 (N_7488,N_6965,N_6921);
nor U7489 (N_7489,N_6982,N_6989);
nor U7490 (N_7490,N_6999,N_6978);
nor U7491 (N_7491,N_7120,N_7105);
and U7492 (N_7492,N_6993,N_7165);
or U7493 (N_7493,N_6948,N_6921);
nor U7494 (N_7494,N_6906,N_7167);
nand U7495 (N_7495,N_7009,N_6996);
or U7496 (N_7496,N_7092,N_7015);
and U7497 (N_7497,N_7082,N_6918);
nor U7498 (N_7498,N_7074,N_7111);
and U7499 (N_7499,N_7131,N_6929);
and U7500 (N_7500,N_7401,N_7455);
xor U7501 (N_7501,N_7289,N_7319);
or U7502 (N_7502,N_7322,N_7353);
nand U7503 (N_7503,N_7463,N_7207);
nand U7504 (N_7504,N_7261,N_7243);
or U7505 (N_7505,N_7350,N_7275);
or U7506 (N_7506,N_7221,N_7390);
nor U7507 (N_7507,N_7254,N_7230);
xnor U7508 (N_7508,N_7364,N_7277);
or U7509 (N_7509,N_7205,N_7303);
xor U7510 (N_7510,N_7325,N_7305);
nor U7511 (N_7511,N_7320,N_7270);
xnor U7512 (N_7512,N_7458,N_7279);
or U7513 (N_7513,N_7404,N_7471);
xnor U7514 (N_7514,N_7371,N_7382);
nor U7515 (N_7515,N_7402,N_7342);
nand U7516 (N_7516,N_7466,N_7233);
nor U7517 (N_7517,N_7328,N_7377);
or U7518 (N_7518,N_7449,N_7400);
xor U7519 (N_7519,N_7271,N_7429);
xor U7520 (N_7520,N_7412,N_7419);
and U7521 (N_7521,N_7389,N_7344);
and U7522 (N_7522,N_7239,N_7286);
nor U7523 (N_7523,N_7487,N_7381);
or U7524 (N_7524,N_7268,N_7385);
or U7525 (N_7525,N_7324,N_7369);
nand U7526 (N_7526,N_7444,N_7365);
xor U7527 (N_7527,N_7311,N_7313);
and U7528 (N_7528,N_7283,N_7329);
and U7529 (N_7529,N_7459,N_7308);
nor U7530 (N_7530,N_7394,N_7301);
nor U7531 (N_7531,N_7264,N_7461);
and U7532 (N_7532,N_7479,N_7440);
xnor U7533 (N_7533,N_7290,N_7464);
and U7534 (N_7534,N_7361,N_7306);
and U7535 (N_7535,N_7240,N_7446);
nand U7536 (N_7536,N_7407,N_7477);
or U7537 (N_7537,N_7293,N_7362);
nor U7538 (N_7538,N_7281,N_7201);
nand U7539 (N_7539,N_7378,N_7409);
or U7540 (N_7540,N_7334,N_7203);
nand U7541 (N_7541,N_7386,N_7476);
nor U7542 (N_7542,N_7478,N_7425);
and U7543 (N_7543,N_7357,N_7310);
and U7544 (N_7544,N_7332,N_7222);
or U7545 (N_7545,N_7421,N_7263);
and U7546 (N_7546,N_7231,N_7383);
xnor U7547 (N_7547,N_7356,N_7349);
nand U7548 (N_7548,N_7360,N_7309);
nand U7549 (N_7549,N_7418,N_7226);
and U7550 (N_7550,N_7292,N_7491);
nor U7551 (N_7551,N_7278,N_7420);
xnor U7552 (N_7552,N_7339,N_7299);
nor U7553 (N_7553,N_7482,N_7341);
or U7554 (N_7554,N_7273,N_7436);
or U7555 (N_7555,N_7314,N_7238);
nor U7556 (N_7556,N_7288,N_7212);
nand U7557 (N_7557,N_7272,N_7416);
and U7558 (N_7558,N_7448,N_7452);
nand U7559 (N_7559,N_7399,N_7225);
xnor U7560 (N_7560,N_7291,N_7468);
and U7561 (N_7561,N_7280,N_7327);
nand U7562 (N_7562,N_7204,N_7200);
xnor U7563 (N_7563,N_7312,N_7375);
and U7564 (N_7564,N_7241,N_7426);
and U7565 (N_7565,N_7331,N_7297);
and U7566 (N_7566,N_7372,N_7494);
xnor U7567 (N_7567,N_7210,N_7257);
nand U7568 (N_7568,N_7262,N_7223);
nand U7569 (N_7569,N_7335,N_7284);
nand U7570 (N_7570,N_7435,N_7247);
and U7571 (N_7571,N_7493,N_7330);
or U7572 (N_7572,N_7411,N_7232);
nand U7573 (N_7573,N_7417,N_7398);
or U7574 (N_7574,N_7220,N_7379);
or U7575 (N_7575,N_7470,N_7216);
xor U7576 (N_7576,N_7498,N_7206);
nand U7577 (N_7577,N_7427,N_7316);
nand U7578 (N_7578,N_7395,N_7246);
nand U7579 (N_7579,N_7408,N_7460);
nand U7580 (N_7580,N_7256,N_7492);
nand U7581 (N_7581,N_7250,N_7454);
nor U7582 (N_7582,N_7323,N_7295);
and U7583 (N_7583,N_7430,N_7218);
and U7584 (N_7584,N_7403,N_7414);
xor U7585 (N_7585,N_7302,N_7442);
and U7586 (N_7586,N_7266,N_7345);
or U7587 (N_7587,N_7433,N_7213);
nor U7588 (N_7588,N_7358,N_7481);
or U7589 (N_7589,N_7431,N_7462);
and U7590 (N_7590,N_7294,N_7483);
nor U7591 (N_7591,N_7488,N_7208);
xor U7592 (N_7592,N_7318,N_7296);
and U7593 (N_7593,N_7443,N_7456);
or U7594 (N_7594,N_7496,N_7287);
xnor U7595 (N_7595,N_7307,N_7260);
and U7596 (N_7596,N_7202,N_7423);
nor U7597 (N_7597,N_7485,N_7392);
or U7598 (N_7598,N_7368,N_7469);
xnor U7599 (N_7599,N_7282,N_7252);
and U7600 (N_7600,N_7234,N_7352);
nor U7601 (N_7601,N_7276,N_7388);
xor U7602 (N_7602,N_7224,N_7317);
or U7603 (N_7603,N_7237,N_7384);
nor U7604 (N_7604,N_7219,N_7450);
or U7605 (N_7605,N_7351,N_7333);
nor U7606 (N_7606,N_7438,N_7336);
nor U7607 (N_7607,N_7391,N_7337);
or U7608 (N_7608,N_7441,N_7214);
nor U7609 (N_7609,N_7253,N_7298);
xor U7610 (N_7610,N_7370,N_7366);
nand U7611 (N_7611,N_7285,N_7367);
xor U7612 (N_7612,N_7248,N_7354);
nor U7613 (N_7613,N_7235,N_7457);
and U7614 (N_7614,N_7413,N_7265);
and U7615 (N_7615,N_7258,N_7359);
or U7616 (N_7616,N_7499,N_7422);
nand U7617 (N_7617,N_7465,N_7405);
or U7618 (N_7618,N_7363,N_7348);
nor U7619 (N_7619,N_7437,N_7236);
nor U7620 (N_7620,N_7259,N_7380);
nor U7621 (N_7621,N_7326,N_7269);
xor U7622 (N_7622,N_7497,N_7484);
xnor U7623 (N_7623,N_7209,N_7267);
or U7624 (N_7624,N_7439,N_7451);
and U7625 (N_7625,N_7393,N_7376);
xor U7626 (N_7626,N_7215,N_7338);
or U7627 (N_7627,N_7227,N_7340);
nand U7628 (N_7628,N_7249,N_7300);
nor U7629 (N_7629,N_7387,N_7467);
nor U7630 (N_7630,N_7406,N_7453);
or U7631 (N_7631,N_7229,N_7490);
nand U7632 (N_7632,N_7374,N_7474);
and U7633 (N_7633,N_7245,N_7415);
or U7634 (N_7634,N_7489,N_7211);
nor U7635 (N_7635,N_7321,N_7217);
nand U7636 (N_7636,N_7473,N_7410);
nor U7637 (N_7637,N_7255,N_7432);
or U7638 (N_7638,N_7396,N_7251);
nor U7639 (N_7639,N_7228,N_7486);
and U7640 (N_7640,N_7424,N_7447);
or U7641 (N_7641,N_7495,N_7315);
nor U7642 (N_7642,N_7355,N_7244);
nand U7643 (N_7643,N_7480,N_7428);
nor U7644 (N_7644,N_7274,N_7346);
and U7645 (N_7645,N_7472,N_7445);
or U7646 (N_7646,N_7373,N_7304);
and U7647 (N_7647,N_7343,N_7434);
nor U7648 (N_7648,N_7347,N_7397);
and U7649 (N_7649,N_7242,N_7475);
or U7650 (N_7650,N_7346,N_7336);
or U7651 (N_7651,N_7288,N_7429);
and U7652 (N_7652,N_7331,N_7308);
nand U7653 (N_7653,N_7259,N_7345);
and U7654 (N_7654,N_7474,N_7436);
or U7655 (N_7655,N_7381,N_7450);
or U7656 (N_7656,N_7413,N_7446);
nand U7657 (N_7657,N_7316,N_7335);
and U7658 (N_7658,N_7240,N_7248);
and U7659 (N_7659,N_7440,N_7225);
nor U7660 (N_7660,N_7484,N_7253);
and U7661 (N_7661,N_7331,N_7479);
or U7662 (N_7662,N_7493,N_7324);
nor U7663 (N_7663,N_7299,N_7234);
nor U7664 (N_7664,N_7463,N_7360);
and U7665 (N_7665,N_7460,N_7272);
nand U7666 (N_7666,N_7463,N_7218);
nand U7667 (N_7667,N_7381,N_7357);
and U7668 (N_7668,N_7338,N_7447);
and U7669 (N_7669,N_7352,N_7423);
xor U7670 (N_7670,N_7324,N_7431);
or U7671 (N_7671,N_7233,N_7369);
and U7672 (N_7672,N_7437,N_7386);
nand U7673 (N_7673,N_7353,N_7355);
and U7674 (N_7674,N_7296,N_7432);
nor U7675 (N_7675,N_7467,N_7232);
xnor U7676 (N_7676,N_7362,N_7220);
nand U7677 (N_7677,N_7266,N_7287);
or U7678 (N_7678,N_7265,N_7280);
and U7679 (N_7679,N_7397,N_7229);
nor U7680 (N_7680,N_7428,N_7403);
or U7681 (N_7681,N_7289,N_7496);
and U7682 (N_7682,N_7274,N_7364);
and U7683 (N_7683,N_7350,N_7408);
nand U7684 (N_7684,N_7426,N_7259);
nor U7685 (N_7685,N_7342,N_7471);
or U7686 (N_7686,N_7280,N_7424);
nor U7687 (N_7687,N_7310,N_7393);
nand U7688 (N_7688,N_7424,N_7217);
or U7689 (N_7689,N_7349,N_7456);
or U7690 (N_7690,N_7360,N_7451);
xnor U7691 (N_7691,N_7467,N_7309);
nor U7692 (N_7692,N_7377,N_7430);
and U7693 (N_7693,N_7218,N_7364);
nand U7694 (N_7694,N_7232,N_7378);
nand U7695 (N_7695,N_7268,N_7371);
and U7696 (N_7696,N_7447,N_7397);
and U7697 (N_7697,N_7424,N_7310);
nand U7698 (N_7698,N_7325,N_7265);
or U7699 (N_7699,N_7327,N_7325);
and U7700 (N_7700,N_7372,N_7269);
nor U7701 (N_7701,N_7487,N_7339);
and U7702 (N_7702,N_7340,N_7463);
nand U7703 (N_7703,N_7359,N_7265);
or U7704 (N_7704,N_7455,N_7233);
or U7705 (N_7705,N_7456,N_7346);
and U7706 (N_7706,N_7413,N_7389);
and U7707 (N_7707,N_7285,N_7303);
nor U7708 (N_7708,N_7475,N_7480);
nor U7709 (N_7709,N_7319,N_7409);
nor U7710 (N_7710,N_7444,N_7368);
xor U7711 (N_7711,N_7434,N_7266);
xnor U7712 (N_7712,N_7292,N_7306);
xnor U7713 (N_7713,N_7404,N_7308);
and U7714 (N_7714,N_7341,N_7246);
and U7715 (N_7715,N_7331,N_7359);
nand U7716 (N_7716,N_7367,N_7427);
nand U7717 (N_7717,N_7467,N_7405);
and U7718 (N_7718,N_7300,N_7460);
nand U7719 (N_7719,N_7294,N_7361);
nand U7720 (N_7720,N_7372,N_7233);
xnor U7721 (N_7721,N_7352,N_7220);
nand U7722 (N_7722,N_7437,N_7384);
nand U7723 (N_7723,N_7267,N_7298);
nand U7724 (N_7724,N_7349,N_7274);
nor U7725 (N_7725,N_7235,N_7450);
xnor U7726 (N_7726,N_7261,N_7331);
nor U7727 (N_7727,N_7389,N_7422);
nand U7728 (N_7728,N_7219,N_7202);
nor U7729 (N_7729,N_7407,N_7301);
nor U7730 (N_7730,N_7348,N_7435);
or U7731 (N_7731,N_7242,N_7443);
or U7732 (N_7732,N_7375,N_7467);
or U7733 (N_7733,N_7246,N_7306);
xnor U7734 (N_7734,N_7291,N_7381);
or U7735 (N_7735,N_7395,N_7350);
xor U7736 (N_7736,N_7469,N_7464);
xor U7737 (N_7737,N_7261,N_7472);
nor U7738 (N_7738,N_7498,N_7304);
or U7739 (N_7739,N_7448,N_7289);
nor U7740 (N_7740,N_7428,N_7408);
and U7741 (N_7741,N_7406,N_7440);
xnor U7742 (N_7742,N_7358,N_7465);
and U7743 (N_7743,N_7233,N_7296);
nand U7744 (N_7744,N_7401,N_7302);
nor U7745 (N_7745,N_7481,N_7280);
and U7746 (N_7746,N_7375,N_7276);
or U7747 (N_7747,N_7408,N_7260);
nor U7748 (N_7748,N_7384,N_7416);
nand U7749 (N_7749,N_7236,N_7249);
xor U7750 (N_7750,N_7491,N_7259);
or U7751 (N_7751,N_7345,N_7249);
xnor U7752 (N_7752,N_7411,N_7287);
nand U7753 (N_7753,N_7373,N_7489);
and U7754 (N_7754,N_7367,N_7310);
nor U7755 (N_7755,N_7251,N_7475);
nor U7756 (N_7756,N_7288,N_7223);
nor U7757 (N_7757,N_7499,N_7232);
nand U7758 (N_7758,N_7322,N_7457);
and U7759 (N_7759,N_7419,N_7443);
nand U7760 (N_7760,N_7430,N_7353);
xor U7761 (N_7761,N_7368,N_7256);
nor U7762 (N_7762,N_7339,N_7375);
nor U7763 (N_7763,N_7349,N_7445);
and U7764 (N_7764,N_7446,N_7350);
xor U7765 (N_7765,N_7302,N_7323);
and U7766 (N_7766,N_7263,N_7468);
nor U7767 (N_7767,N_7347,N_7225);
or U7768 (N_7768,N_7460,N_7223);
or U7769 (N_7769,N_7325,N_7226);
nor U7770 (N_7770,N_7413,N_7436);
nor U7771 (N_7771,N_7302,N_7363);
nor U7772 (N_7772,N_7207,N_7384);
or U7773 (N_7773,N_7465,N_7216);
xor U7774 (N_7774,N_7393,N_7382);
xnor U7775 (N_7775,N_7406,N_7482);
and U7776 (N_7776,N_7387,N_7278);
nor U7777 (N_7777,N_7369,N_7424);
nand U7778 (N_7778,N_7455,N_7319);
and U7779 (N_7779,N_7352,N_7258);
nand U7780 (N_7780,N_7450,N_7392);
and U7781 (N_7781,N_7206,N_7286);
or U7782 (N_7782,N_7218,N_7279);
nand U7783 (N_7783,N_7428,N_7499);
nor U7784 (N_7784,N_7237,N_7278);
nand U7785 (N_7785,N_7476,N_7248);
nor U7786 (N_7786,N_7221,N_7402);
nor U7787 (N_7787,N_7279,N_7399);
nand U7788 (N_7788,N_7363,N_7282);
nand U7789 (N_7789,N_7323,N_7312);
xnor U7790 (N_7790,N_7318,N_7217);
or U7791 (N_7791,N_7291,N_7488);
nor U7792 (N_7792,N_7479,N_7365);
and U7793 (N_7793,N_7348,N_7309);
nor U7794 (N_7794,N_7451,N_7447);
nor U7795 (N_7795,N_7331,N_7419);
and U7796 (N_7796,N_7471,N_7324);
nor U7797 (N_7797,N_7370,N_7453);
or U7798 (N_7798,N_7450,N_7470);
and U7799 (N_7799,N_7264,N_7227);
xor U7800 (N_7800,N_7600,N_7750);
and U7801 (N_7801,N_7714,N_7774);
nor U7802 (N_7802,N_7677,N_7516);
and U7803 (N_7803,N_7503,N_7674);
nor U7804 (N_7804,N_7711,N_7696);
nand U7805 (N_7805,N_7684,N_7785);
nor U7806 (N_7806,N_7584,N_7766);
and U7807 (N_7807,N_7760,N_7756);
xnor U7808 (N_7808,N_7723,N_7567);
and U7809 (N_7809,N_7786,N_7621);
nand U7810 (N_7810,N_7559,N_7616);
and U7811 (N_7811,N_7560,N_7707);
and U7812 (N_7812,N_7724,N_7635);
or U7813 (N_7813,N_7761,N_7783);
nor U7814 (N_7814,N_7590,N_7614);
xnor U7815 (N_7815,N_7619,N_7625);
or U7816 (N_7816,N_7612,N_7541);
or U7817 (N_7817,N_7652,N_7742);
and U7818 (N_7818,N_7535,N_7575);
nand U7819 (N_7819,N_7501,N_7752);
xnor U7820 (N_7820,N_7670,N_7659);
xor U7821 (N_7821,N_7637,N_7609);
xnor U7822 (N_7822,N_7664,N_7610);
xnor U7823 (N_7823,N_7574,N_7645);
or U7824 (N_7824,N_7528,N_7680);
nor U7825 (N_7825,N_7524,N_7613);
nand U7826 (N_7826,N_7718,N_7527);
nand U7827 (N_7827,N_7772,N_7726);
xnor U7828 (N_7828,N_7540,N_7534);
xor U7829 (N_7829,N_7504,N_7639);
nand U7830 (N_7830,N_7626,N_7578);
nor U7831 (N_7831,N_7716,N_7604);
xnor U7832 (N_7832,N_7758,N_7552);
and U7833 (N_7833,N_7517,N_7751);
xnor U7834 (N_7834,N_7562,N_7539);
nor U7835 (N_7835,N_7599,N_7563);
nand U7836 (N_7836,N_7765,N_7569);
nand U7837 (N_7837,N_7520,N_7555);
and U7838 (N_7838,N_7725,N_7721);
nor U7839 (N_7839,N_7530,N_7663);
and U7840 (N_7840,N_7586,N_7737);
nor U7841 (N_7841,N_7757,N_7617);
or U7842 (N_7842,N_7705,N_7576);
and U7843 (N_7843,N_7788,N_7589);
nand U7844 (N_7844,N_7546,N_7717);
nand U7845 (N_7845,N_7722,N_7611);
nand U7846 (N_7846,N_7660,N_7790);
or U7847 (N_7847,N_7633,N_7505);
or U7848 (N_7848,N_7577,N_7720);
nand U7849 (N_7849,N_7697,N_7548);
and U7850 (N_7850,N_7689,N_7566);
or U7851 (N_7851,N_7508,N_7500);
nand U7852 (N_7852,N_7585,N_7688);
nor U7853 (N_7853,N_7671,N_7507);
nor U7854 (N_7854,N_7564,N_7579);
and U7855 (N_7855,N_7768,N_7743);
or U7856 (N_7856,N_7668,N_7654);
xor U7857 (N_7857,N_7525,N_7704);
nand U7858 (N_7858,N_7526,N_7515);
xor U7859 (N_7859,N_7618,N_7657);
nor U7860 (N_7860,N_7538,N_7632);
and U7861 (N_7861,N_7702,N_7665);
and U7862 (N_7862,N_7615,N_7736);
nor U7863 (N_7863,N_7789,N_7588);
nor U7864 (N_7864,N_7506,N_7732);
and U7865 (N_7865,N_7762,N_7798);
or U7866 (N_7866,N_7606,N_7655);
xnor U7867 (N_7867,N_7744,N_7542);
nor U7868 (N_7868,N_7532,N_7636);
or U7869 (N_7869,N_7687,N_7630);
and U7870 (N_7870,N_7767,N_7640);
xor U7871 (N_7871,N_7627,N_7658);
and U7872 (N_7872,N_7690,N_7512);
xor U7873 (N_7873,N_7776,N_7780);
nor U7874 (N_7874,N_7593,N_7691);
nand U7875 (N_7875,N_7649,N_7692);
xor U7876 (N_7876,N_7719,N_7745);
or U7877 (N_7877,N_7667,N_7683);
or U7878 (N_7878,N_7710,N_7675);
and U7879 (N_7879,N_7779,N_7682);
xor U7880 (N_7880,N_7676,N_7746);
and U7881 (N_7881,N_7713,N_7543);
nand U7882 (N_7882,N_7597,N_7522);
and U7883 (N_7883,N_7650,N_7557);
nor U7884 (N_7884,N_7666,N_7729);
and U7885 (N_7885,N_7797,N_7793);
or U7886 (N_7886,N_7608,N_7519);
and U7887 (N_7887,N_7537,N_7603);
or U7888 (N_7888,N_7770,N_7735);
xnor U7889 (N_7889,N_7643,N_7605);
nand U7890 (N_7890,N_7669,N_7741);
xnor U7891 (N_7891,N_7544,N_7749);
xnor U7892 (N_7892,N_7523,N_7738);
or U7893 (N_7893,N_7511,N_7572);
xnor U7894 (N_7894,N_7781,N_7799);
xnor U7895 (N_7895,N_7708,N_7596);
nor U7896 (N_7896,N_7583,N_7554);
or U7897 (N_7897,N_7672,N_7734);
and U7898 (N_7898,N_7698,N_7634);
nor U7899 (N_7899,N_7648,N_7573);
nand U7900 (N_7900,N_7771,N_7775);
or U7901 (N_7901,N_7536,N_7556);
xnor U7902 (N_7902,N_7733,N_7791);
nand U7903 (N_7903,N_7529,N_7518);
nand U7904 (N_7904,N_7551,N_7531);
and U7905 (N_7905,N_7769,N_7792);
and U7906 (N_7906,N_7502,N_7782);
nor U7907 (N_7907,N_7594,N_7715);
nand U7908 (N_7908,N_7582,N_7700);
nand U7909 (N_7909,N_7695,N_7601);
nand U7910 (N_7910,N_7694,N_7784);
nor U7911 (N_7911,N_7623,N_7796);
xor U7912 (N_7912,N_7703,N_7513);
nand U7913 (N_7913,N_7638,N_7685);
and U7914 (N_7914,N_7550,N_7754);
nor U7915 (N_7915,N_7673,N_7509);
or U7916 (N_7916,N_7679,N_7602);
or U7917 (N_7917,N_7701,N_7641);
or U7918 (N_7918,N_7662,N_7607);
nor U7919 (N_7919,N_7709,N_7549);
and U7920 (N_7920,N_7570,N_7624);
nand U7921 (N_7921,N_7739,N_7533);
and U7922 (N_7922,N_7521,N_7706);
or U7923 (N_7923,N_7580,N_7644);
or U7924 (N_7924,N_7545,N_7592);
xor U7925 (N_7925,N_7510,N_7763);
xnor U7926 (N_7926,N_7777,N_7595);
nor U7927 (N_7927,N_7581,N_7755);
and U7928 (N_7928,N_7642,N_7598);
xnor U7929 (N_7929,N_7565,N_7661);
xnor U7930 (N_7930,N_7656,N_7678);
xor U7931 (N_7931,N_7568,N_7686);
or U7932 (N_7932,N_7558,N_7571);
and U7933 (N_7933,N_7727,N_7764);
xor U7934 (N_7934,N_7778,N_7651);
nor U7935 (N_7935,N_7795,N_7728);
or U7936 (N_7936,N_7628,N_7794);
nand U7937 (N_7937,N_7622,N_7553);
or U7938 (N_7938,N_7759,N_7591);
nor U7939 (N_7939,N_7653,N_7631);
nand U7940 (N_7940,N_7629,N_7699);
nand U7941 (N_7941,N_7748,N_7514);
and U7942 (N_7942,N_7773,N_7561);
or U7943 (N_7943,N_7731,N_7712);
nor U7944 (N_7944,N_7681,N_7547);
xnor U7945 (N_7945,N_7753,N_7730);
and U7946 (N_7946,N_7647,N_7646);
and U7947 (N_7947,N_7693,N_7620);
nor U7948 (N_7948,N_7747,N_7787);
nor U7949 (N_7949,N_7587,N_7740);
xnor U7950 (N_7950,N_7543,N_7720);
and U7951 (N_7951,N_7685,N_7599);
nand U7952 (N_7952,N_7524,N_7538);
and U7953 (N_7953,N_7534,N_7787);
xor U7954 (N_7954,N_7788,N_7793);
nand U7955 (N_7955,N_7538,N_7737);
nor U7956 (N_7956,N_7745,N_7715);
and U7957 (N_7957,N_7569,N_7777);
or U7958 (N_7958,N_7538,N_7577);
xnor U7959 (N_7959,N_7537,N_7694);
and U7960 (N_7960,N_7781,N_7694);
and U7961 (N_7961,N_7574,N_7674);
nand U7962 (N_7962,N_7505,N_7683);
nand U7963 (N_7963,N_7793,N_7737);
or U7964 (N_7964,N_7753,N_7740);
nor U7965 (N_7965,N_7772,N_7743);
xnor U7966 (N_7966,N_7556,N_7779);
and U7967 (N_7967,N_7666,N_7694);
nor U7968 (N_7968,N_7596,N_7739);
xnor U7969 (N_7969,N_7537,N_7621);
and U7970 (N_7970,N_7510,N_7757);
nand U7971 (N_7971,N_7640,N_7699);
nor U7972 (N_7972,N_7584,N_7721);
nor U7973 (N_7973,N_7589,N_7687);
or U7974 (N_7974,N_7566,N_7757);
xor U7975 (N_7975,N_7526,N_7662);
nor U7976 (N_7976,N_7640,N_7710);
xor U7977 (N_7977,N_7539,N_7607);
or U7978 (N_7978,N_7752,N_7640);
nand U7979 (N_7979,N_7505,N_7554);
or U7980 (N_7980,N_7658,N_7540);
xnor U7981 (N_7981,N_7691,N_7790);
nor U7982 (N_7982,N_7676,N_7644);
and U7983 (N_7983,N_7693,N_7762);
nand U7984 (N_7984,N_7721,N_7663);
nor U7985 (N_7985,N_7667,N_7678);
and U7986 (N_7986,N_7615,N_7566);
nand U7987 (N_7987,N_7516,N_7573);
xnor U7988 (N_7988,N_7557,N_7786);
nand U7989 (N_7989,N_7502,N_7591);
nor U7990 (N_7990,N_7736,N_7676);
and U7991 (N_7991,N_7509,N_7587);
and U7992 (N_7992,N_7742,N_7703);
nor U7993 (N_7993,N_7570,N_7534);
nor U7994 (N_7994,N_7711,N_7783);
and U7995 (N_7995,N_7687,N_7625);
and U7996 (N_7996,N_7645,N_7650);
and U7997 (N_7997,N_7718,N_7792);
and U7998 (N_7998,N_7643,N_7653);
or U7999 (N_7999,N_7675,N_7683);
and U8000 (N_8000,N_7630,N_7608);
nand U8001 (N_8001,N_7752,N_7581);
xnor U8002 (N_8002,N_7528,N_7621);
nand U8003 (N_8003,N_7735,N_7618);
nand U8004 (N_8004,N_7565,N_7660);
or U8005 (N_8005,N_7591,N_7631);
or U8006 (N_8006,N_7557,N_7552);
nand U8007 (N_8007,N_7738,N_7703);
nand U8008 (N_8008,N_7764,N_7766);
or U8009 (N_8009,N_7515,N_7503);
or U8010 (N_8010,N_7628,N_7780);
nor U8011 (N_8011,N_7726,N_7699);
or U8012 (N_8012,N_7703,N_7629);
or U8013 (N_8013,N_7738,N_7579);
and U8014 (N_8014,N_7529,N_7757);
nand U8015 (N_8015,N_7641,N_7727);
nand U8016 (N_8016,N_7560,N_7712);
xnor U8017 (N_8017,N_7557,N_7762);
or U8018 (N_8018,N_7592,N_7757);
nor U8019 (N_8019,N_7529,N_7750);
nand U8020 (N_8020,N_7589,N_7605);
xor U8021 (N_8021,N_7517,N_7513);
or U8022 (N_8022,N_7606,N_7694);
nand U8023 (N_8023,N_7537,N_7738);
nand U8024 (N_8024,N_7504,N_7720);
and U8025 (N_8025,N_7502,N_7622);
and U8026 (N_8026,N_7521,N_7620);
nand U8027 (N_8027,N_7778,N_7625);
nand U8028 (N_8028,N_7791,N_7501);
xor U8029 (N_8029,N_7591,N_7628);
xor U8030 (N_8030,N_7711,N_7787);
xor U8031 (N_8031,N_7762,N_7531);
nand U8032 (N_8032,N_7552,N_7559);
or U8033 (N_8033,N_7738,N_7633);
nand U8034 (N_8034,N_7536,N_7792);
or U8035 (N_8035,N_7604,N_7602);
and U8036 (N_8036,N_7711,N_7729);
nand U8037 (N_8037,N_7516,N_7660);
nor U8038 (N_8038,N_7763,N_7636);
or U8039 (N_8039,N_7537,N_7569);
nor U8040 (N_8040,N_7723,N_7720);
nor U8041 (N_8041,N_7573,N_7668);
or U8042 (N_8042,N_7503,N_7678);
or U8043 (N_8043,N_7665,N_7522);
nand U8044 (N_8044,N_7789,N_7530);
nand U8045 (N_8045,N_7509,N_7707);
nand U8046 (N_8046,N_7674,N_7597);
nand U8047 (N_8047,N_7608,N_7592);
and U8048 (N_8048,N_7626,N_7730);
and U8049 (N_8049,N_7673,N_7717);
or U8050 (N_8050,N_7735,N_7793);
nand U8051 (N_8051,N_7606,N_7515);
nor U8052 (N_8052,N_7500,N_7705);
nor U8053 (N_8053,N_7701,N_7727);
xnor U8054 (N_8054,N_7503,N_7524);
xnor U8055 (N_8055,N_7736,N_7534);
or U8056 (N_8056,N_7720,N_7785);
and U8057 (N_8057,N_7783,N_7587);
and U8058 (N_8058,N_7693,N_7750);
and U8059 (N_8059,N_7721,N_7733);
xor U8060 (N_8060,N_7722,N_7767);
nor U8061 (N_8061,N_7759,N_7735);
and U8062 (N_8062,N_7765,N_7742);
nand U8063 (N_8063,N_7756,N_7626);
or U8064 (N_8064,N_7753,N_7577);
nor U8065 (N_8065,N_7575,N_7512);
xor U8066 (N_8066,N_7669,N_7660);
nand U8067 (N_8067,N_7506,N_7588);
nor U8068 (N_8068,N_7571,N_7505);
nand U8069 (N_8069,N_7764,N_7796);
nand U8070 (N_8070,N_7614,N_7750);
nor U8071 (N_8071,N_7600,N_7500);
xnor U8072 (N_8072,N_7516,N_7688);
or U8073 (N_8073,N_7626,N_7509);
nand U8074 (N_8074,N_7594,N_7656);
xnor U8075 (N_8075,N_7641,N_7577);
xnor U8076 (N_8076,N_7541,N_7711);
or U8077 (N_8077,N_7772,N_7785);
xnor U8078 (N_8078,N_7679,N_7644);
nand U8079 (N_8079,N_7541,N_7762);
xnor U8080 (N_8080,N_7756,N_7563);
and U8081 (N_8081,N_7747,N_7753);
nand U8082 (N_8082,N_7562,N_7611);
and U8083 (N_8083,N_7558,N_7622);
nor U8084 (N_8084,N_7797,N_7556);
nand U8085 (N_8085,N_7506,N_7673);
and U8086 (N_8086,N_7572,N_7772);
and U8087 (N_8087,N_7639,N_7583);
and U8088 (N_8088,N_7783,N_7674);
and U8089 (N_8089,N_7728,N_7759);
or U8090 (N_8090,N_7710,N_7549);
nor U8091 (N_8091,N_7567,N_7575);
and U8092 (N_8092,N_7529,N_7652);
or U8093 (N_8093,N_7519,N_7515);
nand U8094 (N_8094,N_7663,N_7755);
and U8095 (N_8095,N_7570,N_7663);
xor U8096 (N_8096,N_7749,N_7509);
and U8097 (N_8097,N_7525,N_7787);
and U8098 (N_8098,N_7561,N_7793);
and U8099 (N_8099,N_7734,N_7515);
nand U8100 (N_8100,N_8066,N_8061);
nand U8101 (N_8101,N_7864,N_8078);
nand U8102 (N_8102,N_7803,N_8024);
nor U8103 (N_8103,N_7894,N_7959);
xor U8104 (N_8104,N_7980,N_7833);
nor U8105 (N_8105,N_7891,N_8038);
xor U8106 (N_8106,N_8065,N_7809);
or U8107 (N_8107,N_7879,N_8050);
xor U8108 (N_8108,N_7811,N_7929);
or U8109 (N_8109,N_7848,N_7961);
nor U8110 (N_8110,N_8004,N_7912);
or U8111 (N_8111,N_8032,N_8076);
and U8112 (N_8112,N_8006,N_7883);
or U8113 (N_8113,N_7934,N_8027);
nor U8114 (N_8114,N_7839,N_8011);
and U8115 (N_8115,N_7889,N_8088);
xor U8116 (N_8116,N_7815,N_8068);
or U8117 (N_8117,N_7945,N_8080);
or U8118 (N_8118,N_7899,N_7947);
and U8119 (N_8119,N_7876,N_7994);
nor U8120 (N_8120,N_8072,N_7919);
nand U8121 (N_8121,N_7996,N_7874);
xor U8122 (N_8122,N_7862,N_7953);
nor U8123 (N_8123,N_7946,N_8036);
nand U8124 (N_8124,N_7856,N_7829);
nand U8125 (N_8125,N_8033,N_7855);
nand U8126 (N_8126,N_7888,N_8074);
nand U8127 (N_8127,N_7968,N_8012);
nand U8128 (N_8128,N_7970,N_7927);
or U8129 (N_8129,N_7985,N_7963);
nand U8130 (N_8130,N_7886,N_8093);
nor U8131 (N_8131,N_7906,N_7885);
or U8132 (N_8132,N_7917,N_8060);
or U8133 (N_8133,N_7853,N_8086);
or U8134 (N_8134,N_7974,N_8040);
nor U8135 (N_8135,N_7805,N_7926);
and U8136 (N_8136,N_7863,N_8057);
nand U8137 (N_8137,N_7852,N_7893);
or U8138 (N_8138,N_7903,N_7965);
nor U8139 (N_8139,N_7824,N_7860);
nand U8140 (N_8140,N_8037,N_7958);
or U8141 (N_8141,N_8071,N_7867);
nor U8142 (N_8142,N_7928,N_8089);
nor U8143 (N_8143,N_8022,N_7982);
and U8144 (N_8144,N_8092,N_7827);
nand U8145 (N_8145,N_7924,N_7819);
nand U8146 (N_8146,N_8000,N_8042);
xor U8147 (N_8147,N_8067,N_7804);
xnor U8148 (N_8148,N_7972,N_7964);
xnor U8149 (N_8149,N_8010,N_7909);
nor U8150 (N_8150,N_8025,N_7812);
and U8151 (N_8151,N_8028,N_8070);
nand U8152 (N_8152,N_8069,N_7998);
nand U8153 (N_8153,N_7977,N_7878);
or U8154 (N_8154,N_7845,N_8009);
xor U8155 (N_8155,N_8075,N_7895);
xor U8156 (N_8156,N_7918,N_8083);
xnor U8157 (N_8157,N_7957,N_8023);
and U8158 (N_8158,N_7822,N_8013);
and U8159 (N_8159,N_7941,N_7988);
or U8160 (N_8160,N_7814,N_8098);
nand U8161 (N_8161,N_7887,N_8002);
and U8162 (N_8162,N_7971,N_8087);
nor U8163 (N_8163,N_7841,N_8017);
nor U8164 (N_8164,N_7881,N_7826);
and U8165 (N_8165,N_7849,N_7992);
and U8166 (N_8166,N_7933,N_8016);
xnor U8167 (N_8167,N_7817,N_7984);
and U8168 (N_8168,N_8035,N_7902);
or U8169 (N_8169,N_7806,N_7979);
xnor U8170 (N_8170,N_7956,N_7830);
and U8171 (N_8171,N_8056,N_7935);
nor U8172 (N_8172,N_8019,N_8034);
or U8173 (N_8173,N_7834,N_7844);
nor U8174 (N_8174,N_7859,N_7869);
nand U8175 (N_8175,N_7892,N_7868);
xnor U8176 (N_8176,N_8029,N_7955);
nor U8177 (N_8177,N_7975,N_7914);
nor U8178 (N_8178,N_8084,N_7816);
xnor U8179 (N_8179,N_7991,N_7837);
nor U8180 (N_8180,N_7925,N_7931);
and U8181 (N_8181,N_8064,N_7952);
nor U8182 (N_8182,N_8041,N_8051);
or U8183 (N_8183,N_7904,N_7949);
or U8184 (N_8184,N_7872,N_7801);
nand U8185 (N_8185,N_7897,N_7967);
nand U8186 (N_8186,N_7880,N_7911);
xnor U8187 (N_8187,N_8039,N_8055);
and U8188 (N_8188,N_7978,N_7983);
or U8189 (N_8189,N_7847,N_7989);
nor U8190 (N_8190,N_8096,N_7908);
xor U8191 (N_8191,N_8095,N_7832);
nor U8192 (N_8192,N_7866,N_7937);
or U8193 (N_8193,N_7802,N_7820);
or U8194 (N_8194,N_7901,N_7861);
nand U8195 (N_8195,N_7951,N_7865);
nand U8196 (N_8196,N_8079,N_7884);
nand U8197 (N_8197,N_8059,N_8014);
and U8198 (N_8198,N_8030,N_7896);
nor U8199 (N_8199,N_8044,N_7831);
and U8200 (N_8200,N_8099,N_7843);
xor U8201 (N_8201,N_7943,N_8091);
xor U8202 (N_8202,N_7990,N_7987);
or U8203 (N_8203,N_7916,N_8052);
nand U8204 (N_8204,N_7915,N_8073);
or U8205 (N_8205,N_7840,N_8094);
nor U8206 (N_8206,N_7873,N_7950);
nand U8207 (N_8207,N_7932,N_7942);
nand U8208 (N_8208,N_8021,N_8047);
and U8209 (N_8209,N_7858,N_7923);
nand U8210 (N_8210,N_7821,N_7875);
xnor U8211 (N_8211,N_7810,N_7838);
nand U8212 (N_8212,N_8054,N_8003);
nand U8213 (N_8213,N_8015,N_8082);
nor U8214 (N_8214,N_7940,N_8090);
nand U8215 (N_8215,N_7857,N_7999);
and U8216 (N_8216,N_7939,N_7997);
xnor U8217 (N_8217,N_8081,N_7800);
or U8218 (N_8218,N_7920,N_8043);
or U8219 (N_8219,N_7900,N_7981);
or U8220 (N_8220,N_7944,N_7871);
xnor U8221 (N_8221,N_7973,N_7854);
or U8222 (N_8222,N_7995,N_7823);
nand U8223 (N_8223,N_7910,N_8020);
or U8224 (N_8224,N_8046,N_7969);
and U8225 (N_8225,N_8007,N_7938);
nand U8226 (N_8226,N_8063,N_7846);
xnor U8227 (N_8227,N_7825,N_7818);
nor U8228 (N_8228,N_7808,N_7850);
xor U8229 (N_8229,N_7807,N_7842);
or U8230 (N_8230,N_8026,N_8031);
or U8231 (N_8231,N_7813,N_7960);
nor U8232 (N_8232,N_7890,N_8005);
nand U8233 (N_8233,N_7828,N_8085);
nand U8234 (N_8234,N_7948,N_7835);
and U8235 (N_8235,N_8077,N_8048);
nand U8236 (N_8236,N_7966,N_8018);
or U8237 (N_8237,N_7913,N_8062);
xor U8238 (N_8238,N_7898,N_7936);
and U8239 (N_8239,N_8045,N_7907);
xor U8240 (N_8240,N_7962,N_8001);
or U8241 (N_8241,N_7836,N_8049);
nand U8242 (N_8242,N_7870,N_8053);
or U8243 (N_8243,N_8097,N_7851);
nor U8244 (N_8244,N_8008,N_7986);
xnor U8245 (N_8245,N_7922,N_7930);
or U8246 (N_8246,N_7993,N_7882);
xor U8247 (N_8247,N_7954,N_7976);
or U8248 (N_8248,N_7921,N_7905);
and U8249 (N_8249,N_7877,N_8058);
or U8250 (N_8250,N_7921,N_8019);
and U8251 (N_8251,N_8056,N_7876);
and U8252 (N_8252,N_8058,N_7925);
nor U8253 (N_8253,N_7880,N_8093);
nand U8254 (N_8254,N_7919,N_7909);
xor U8255 (N_8255,N_7889,N_7872);
nor U8256 (N_8256,N_7914,N_8063);
nand U8257 (N_8257,N_7894,N_8072);
nand U8258 (N_8258,N_8058,N_7929);
xnor U8259 (N_8259,N_7984,N_7847);
nor U8260 (N_8260,N_7829,N_7943);
nor U8261 (N_8261,N_7900,N_7920);
or U8262 (N_8262,N_7866,N_7836);
xnor U8263 (N_8263,N_8054,N_7904);
or U8264 (N_8264,N_7830,N_7842);
or U8265 (N_8265,N_7830,N_7849);
nand U8266 (N_8266,N_7992,N_8037);
nor U8267 (N_8267,N_7927,N_7883);
nand U8268 (N_8268,N_7828,N_7807);
or U8269 (N_8269,N_7879,N_7887);
or U8270 (N_8270,N_7881,N_8076);
nor U8271 (N_8271,N_7876,N_7986);
nor U8272 (N_8272,N_7904,N_8033);
nor U8273 (N_8273,N_7816,N_8010);
nor U8274 (N_8274,N_7862,N_7835);
nor U8275 (N_8275,N_8097,N_7981);
nor U8276 (N_8276,N_7849,N_8067);
nor U8277 (N_8277,N_7981,N_7834);
nand U8278 (N_8278,N_8048,N_8071);
and U8279 (N_8279,N_7963,N_8038);
nor U8280 (N_8280,N_7900,N_8012);
nand U8281 (N_8281,N_8082,N_7975);
nor U8282 (N_8282,N_7975,N_7929);
or U8283 (N_8283,N_8017,N_7809);
nand U8284 (N_8284,N_7947,N_8027);
nor U8285 (N_8285,N_7974,N_7812);
nand U8286 (N_8286,N_7984,N_8050);
or U8287 (N_8287,N_8053,N_7910);
nand U8288 (N_8288,N_7999,N_7804);
xnor U8289 (N_8289,N_8081,N_8052);
nand U8290 (N_8290,N_7974,N_8042);
or U8291 (N_8291,N_7853,N_7995);
and U8292 (N_8292,N_7922,N_7820);
and U8293 (N_8293,N_7931,N_8060);
nand U8294 (N_8294,N_7959,N_8022);
nand U8295 (N_8295,N_8092,N_7978);
nor U8296 (N_8296,N_7941,N_7860);
and U8297 (N_8297,N_7834,N_8039);
xor U8298 (N_8298,N_7855,N_8047);
or U8299 (N_8299,N_8002,N_7859);
and U8300 (N_8300,N_8085,N_7823);
xnor U8301 (N_8301,N_8059,N_7860);
and U8302 (N_8302,N_7984,N_7851);
xor U8303 (N_8303,N_7875,N_8092);
or U8304 (N_8304,N_8048,N_8068);
xor U8305 (N_8305,N_7979,N_7893);
xor U8306 (N_8306,N_8050,N_7917);
or U8307 (N_8307,N_7976,N_8076);
nand U8308 (N_8308,N_7987,N_7860);
xnor U8309 (N_8309,N_8094,N_7912);
and U8310 (N_8310,N_7951,N_7880);
nand U8311 (N_8311,N_7900,N_7825);
or U8312 (N_8312,N_8084,N_8092);
nand U8313 (N_8313,N_7968,N_8017);
and U8314 (N_8314,N_8094,N_7917);
and U8315 (N_8315,N_7964,N_7827);
nor U8316 (N_8316,N_7931,N_7854);
xor U8317 (N_8317,N_7933,N_8055);
nor U8318 (N_8318,N_8061,N_7910);
and U8319 (N_8319,N_8049,N_7865);
or U8320 (N_8320,N_7983,N_8045);
nand U8321 (N_8321,N_7884,N_7951);
nand U8322 (N_8322,N_7964,N_7887);
nand U8323 (N_8323,N_7992,N_7913);
nor U8324 (N_8324,N_7880,N_8007);
nor U8325 (N_8325,N_8013,N_7931);
xnor U8326 (N_8326,N_8097,N_7948);
xnor U8327 (N_8327,N_7838,N_7894);
and U8328 (N_8328,N_7876,N_7953);
nor U8329 (N_8329,N_8072,N_7869);
or U8330 (N_8330,N_7954,N_7952);
and U8331 (N_8331,N_8062,N_7897);
nor U8332 (N_8332,N_7888,N_7896);
nor U8333 (N_8333,N_7805,N_8004);
nor U8334 (N_8334,N_8071,N_7830);
nand U8335 (N_8335,N_7875,N_7978);
nand U8336 (N_8336,N_7996,N_7907);
nor U8337 (N_8337,N_8079,N_8089);
nand U8338 (N_8338,N_7933,N_7937);
or U8339 (N_8339,N_7947,N_7951);
nand U8340 (N_8340,N_8058,N_7915);
and U8341 (N_8341,N_7999,N_7888);
xnor U8342 (N_8342,N_7926,N_7995);
nor U8343 (N_8343,N_7847,N_8081);
and U8344 (N_8344,N_7821,N_7918);
xnor U8345 (N_8345,N_7863,N_8058);
nand U8346 (N_8346,N_7869,N_7996);
nor U8347 (N_8347,N_7868,N_7952);
nor U8348 (N_8348,N_8019,N_7875);
nand U8349 (N_8349,N_8074,N_7931);
or U8350 (N_8350,N_7932,N_7871);
xnor U8351 (N_8351,N_8085,N_8035);
and U8352 (N_8352,N_8043,N_8069);
nor U8353 (N_8353,N_7939,N_7803);
nor U8354 (N_8354,N_8068,N_7880);
and U8355 (N_8355,N_8075,N_7850);
nand U8356 (N_8356,N_7835,N_7954);
xor U8357 (N_8357,N_8026,N_8046);
nor U8358 (N_8358,N_7823,N_7876);
or U8359 (N_8359,N_7979,N_8020);
xnor U8360 (N_8360,N_8047,N_7810);
and U8361 (N_8361,N_7963,N_8085);
xor U8362 (N_8362,N_8014,N_8083);
or U8363 (N_8363,N_7916,N_7921);
or U8364 (N_8364,N_8013,N_7846);
xor U8365 (N_8365,N_7843,N_8050);
xnor U8366 (N_8366,N_7985,N_7965);
nand U8367 (N_8367,N_7893,N_8066);
or U8368 (N_8368,N_8087,N_7819);
nor U8369 (N_8369,N_7899,N_8037);
nor U8370 (N_8370,N_7997,N_7974);
nor U8371 (N_8371,N_7909,N_7893);
nand U8372 (N_8372,N_8019,N_7899);
or U8373 (N_8373,N_7995,N_7989);
nand U8374 (N_8374,N_7995,N_8031);
or U8375 (N_8375,N_7861,N_7976);
or U8376 (N_8376,N_8098,N_7948);
nand U8377 (N_8377,N_7912,N_7911);
or U8378 (N_8378,N_7832,N_8019);
or U8379 (N_8379,N_8086,N_7966);
nor U8380 (N_8380,N_7858,N_7978);
or U8381 (N_8381,N_7848,N_7933);
and U8382 (N_8382,N_7912,N_8027);
or U8383 (N_8383,N_7953,N_8033);
nand U8384 (N_8384,N_8017,N_8022);
nor U8385 (N_8385,N_7830,N_7934);
and U8386 (N_8386,N_7946,N_8050);
nand U8387 (N_8387,N_7881,N_8088);
or U8388 (N_8388,N_7920,N_7907);
nand U8389 (N_8389,N_8059,N_8096);
xor U8390 (N_8390,N_7972,N_7879);
nor U8391 (N_8391,N_7883,N_7951);
or U8392 (N_8392,N_7839,N_7874);
nand U8393 (N_8393,N_7811,N_7926);
xnor U8394 (N_8394,N_7922,N_8090);
and U8395 (N_8395,N_7887,N_8067);
or U8396 (N_8396,N_7994,N_8070);
xnor U8397 (N_8397,N_7904,N_7948);
or U8398 (N_8398,N_8081,N_8022);
nor U8399 (N_8399,N_7928,N_7821);
nor U8400 (N_8400,N_8174,N_8349);
nor U8401 (N_8401,N_8242,N_8385);
nand U8402 (N_8402,N_8186,N_8295);
xor U8403 (N_8403,N_8221,N_8289);
or U8404 (N_8404,N_8283,N_8201);
nor U8405 (N_8405,N_8358,N_8264);
xnor U8406 (N_8406,N_8372,N_8311);
nand U8407 (N_8407,N_8388,N_8352);
or U8408 (N_8408,N_8200,N_8184);
nand U8409 (N_8409,N_8206,N_8393);
and U8410 (N_8410,N_8226,N_8116);
or U8411 (N_8411,N_8222,N_8287);
or U8412 (N_8412,N_8111,N_8270);
xnor U8413 (N_8413,N_8110,N_8359);
and U8414 (N_8414,N_8119,N_8371);
xnor U8415 (N_8415,N_8387,N_8175);
xor U8416 (N_8416,N_8165,N_8275);
nor U8417 (N_8417,N_8172,N_8310);
and U8418 (N_8418,N_8229,N_8170);
and U8419 (N_8419,N_8203,N_8292);
or U8420 (N_8420,N_8231,N_8139);
and U8421 (N_8421,N_8301,N_8215);
xnor U8422 (N_8422,N_8339,N_8363);
nand U8423 (N_8423,N_8160,N_8266);
and U8424 (N_8424,N_8317,N_8218);
or U8425 (N_8425,N_8233,N_8282);
nand U8426 (N_8426,N_8183,N_8223);
xor U8427 (N_8427,N_8300,N_8374);
nand U8428 (N_8428,N_8255,N_8258);
and U8429 (N_8429,N_8128,N_8336);
and U8430 (N_8430,N_8152,N_8217);
and U8431 (N_8431,N_8386,N_8316);
xnor U8432 (N_8432,N_8271,N_8357);
nor U8433 (N_8433,N_8296,N_8308);
nand U8434 (N_8434,N_8273,N_8360);
nand U8435 (N_8435,N_8396,N_8199);
nand U8436 (N_8436,N_8168,N_8328);
xor U8437 (N_8437,N_8395,N_8265);
nor U8438 (N_8438,N_8305,N_8190);
and U8439 (N_8439,N_8104,N_8167);
and U8440 (N_8440,N_8241,N_8147);
nor U8441 (N_8441,N_8345,N_8375);
xnor U8442 (N_8442,N_8248,N_8120);
xor U8443 (N_8443,N_8333,N_8319);
nor U8444 (N_8444,N_8114,N_8259);
xor U8445 (N_8445,N_8195,N_8362);
and U8446 (N_8446,N_8234,N_8125);
xnor U8447 (N_8447,N_8324,N_8197);
nor U8448 (N_8448,N_8103,N_8252);
xnor U8449 (N_8449,N_8394,N_8361);
xnor U8450 (N_8450,N_8102,N_8127);
and U8451 (N_8451,N_8318,N_8340);
or U8452 (N_8452,N_8214,N_8192);
or U8453 (N_8453,N_8398,N_8124);
xor U8454 (N_8454,N_8173,N_8341);
nor U8455 (N_8455,N_8299,N_8205);
nand U8456 (N_8456,N_8288,N_8213);
or U8457 (N_8457,N_8159,N_8302);
nor U8458 (N_8458,N_8377,N_8212);
and U8459 (N_8459,N_8101,N_8312);
xor U8460 (N_8460,N_8364,N_8356);
nor U8461 (N_8461,N_8331,N_8198);
or U8462 (N_8462,N_8293,N_8137);
nor U8463 (N_8463,N_8368,N_8251);
xor U8464 (N_8464,N_8244,N_8100);
or U8465 (N_8465,N_8188,N_8237);
and U8466 (N_8466,N_8370,N_8391);
nand U8467 (N_8467,N_8323,N_8381);
nand U8468 (N_8468,N_8144,N_8384);
and U8469 (N_8469,N_8254,N_8366);
and U8470 (N_8470,N_8194,N_8397);
nand U8471 (N_8471,N_8109,N_8353);
nor U8472 (N_8472,N_8278,N_8187);
or U8473 (N_8473,N_8193,N_8150);
or U8474 (N_8474,N_8162,N_8281);
or U8475 (N_8475,N_8228,N_8351);
nand U8476 (N_8476,N_8290,N_8247);
or U8477 (N_8477,N_8269,N_8294);
xnor U8478 (N_8478,N_8344,N_8130);
or U8479 (N_8479,N_8123,N_8141);
nand U8480 (N_8480,N_8304,N_8315);
nor U8481 (N_8481,N_8291,N_8298);
or U8482 (N_8482,N_8327,N_8367);
xnor U8483 (N_8483,N_8179,N_8376);
xnor U8484 (N_8484,N_8240,N_8332);
nor U8485 (N_8485,N_8224,N_8106);
and U8486 (N_8486,N_8121,N_8209);
xnor U8487 (N_8487,N_8325,N_8134);
nor U8488 (N_8488,N_8346,N_8202);
xnor U8489 (N_8489,N_8280,N_8232);
xnor U8490 (N_8490,N_8143,N_8149);
and U8491 (N_8491,N_8338,N_8286);
xor U8492 (N_8492,N_8238,N_8140);
nand U8493 (N_8493,N_8135,N_8354);
nor U8494 (N_8494,N_8256,N_8330);
or U8495 (N_8495,N_8313,N_8274);
and U8496 (N_8496,N_8230,N_8245);
nand U8497 (N_8497,N_8243,N_8322);
and U8498 (N_8498,N_8284,N_8306);
xor U8499 (N_8499,N_8285,N_8161);
or U8500 (N_8500,N_8207,N_8138);
nand U8501 (N_8501,N_8343,N_8335);
xor U8502 (N_8502,N_8276,N_8369);
or U8503 (N_8503,N_8392,N_8383);
nor U8504 (N_8504,N_8334,N_8189);
and U8505 (N_8505,N_8157,N_8262);
nand U8506 (N_8506,N_8191,N_8216);
or U8507 (N_8507,N_8151,N_8380);
nor U8508 (N_8508,N_8155,N_8178);
nor U8509 (N_8509,N_8122,N_8181);
nand U8510 (N_8510,N_8129,N_8177);
or U8511 (N_8511,N_8378,N_8272);
or U8512 (N_8512,N_8148,N_8277);
xor U8513 (N_8513,N_8303,N_8118);
xor U8514 (N_8514,N_8166,N_8350);
or U8515 (N_8515,N_8132,N_8268);
and U8516 (N_8516,N_8107,N_8297);
and U8517 (N_8517,N_8133,N_8236);
nor U8518 (N_8518,N_8365,N_8113);
or U8519 (N_8519,N_8250,N_8257);
nand U8520 (N_8520,N_8267,N_8320);
or U8521 (N_8521,N_8220,N_8342);
nor U8522 (N_8522,N_8182,N_8249);
or U8523 (N_8523,N_8145,N_8105);
nor U8524 (N_8524,N_8390,N_8261);
xnor U8525 (N_8525,N_8235,N_8309);
nor U8526 (N_8526,N_8142,N_8314);
xnor U8527 (N_8527,N_8108,N_8211);
and U8528 (N_8528,N_8185,N_8347);
nand U8529 (N_8529,N_8326,N_8329);
xnor U8530 (N_8530,N_8379,N_8136);
nor U8531 (N_8531,N_8337,N_8117);
nor U8532 (N_8532,N_8382,N_8171);
nor U8533 (N_8533,N_8146,N_8263);
and U8534 (N_8534,N_8204,N_8126);
nor U8535 (N_8535,N_8389,N_8115);
xor U8536 (N_8536,N_8156,N_8196);
nand U8537 (N_8537,N_8253,N_8112);
or U8538 (N_8538,N_8169,N_8260);
or U8539 (N_8539,N_8373,N_8154);
or U8540 (N_8540,N_8355,N_8225);
nand U8541 (N_8541,N_8176,N_8246);
xnor U8542 (N_8542,N_8153,N_8307);
nor U8543 (N_8543,N_8164,N_8208);
nand U8544 (N_8544,N_8227,N_8210);
and U8545 (N_8545,N_8321,N_8163);
nand U8546 (N_8546,N_8348,N_8131);
nand U8547 (N_8547,N_8158,N_8279);
nand U8548 (N_8548,N_8399,N_8239);
nand U8549 (N_8549,N_8180,N_8219);
or U8550 (N_8550,N_8173,N_8246);
and U8551 (N_8551,N_8103,N_8323);
and U8552 (N_8552,N_8227,N_8104);
and U8553 (N_8553,N_8232,N_8142);
nand U8554 (N_8554,N_8179,N_8112);
or U8555 (N_8555,N_8128,N_8337);
and U8556 (N_8556,N_8322,N_8175);
or U8557 (N_8557,N_8308,N_8197);
nor U8558 (N_8558,N_8367,N_8305);
xor U8559 (N_8559,N_8278,N_8363);
or U8560 (N_8560,N_8387,N_8327);
xor U8561 (N_8561,N_8183,N_8366);
and U8562 (N_8562,N_8379,N_8106);
nand U8563 (N_8563,N_8143,N_8298);
xor U8564 (N_8564,N_8244,N_8140);
and U8565 (N_8565,N_8185,N_8243);
or U8566 (N_8566,N_8159,N_8111);
or U8567 (N_8567,N_8182,N_8253);
xor U8568 (N_8568,N_8396,N_8149);
nor U8569 (N_8569,N_8214,N_8398);
xor U8570 (N_8570,N_8325,N_8323);
and U8571 (N_8571,N_8300,N_8396);
nand U8572 (N_8572,N_8239,N_8177);
and U8573 (N_8573,N_8220,N_8119);
nand U8574 (N_8574,N_8172,N_8168);
xor U8575 (N_8575,N_8204,N_8293);
nand U8576 (N_8576,N_8360,N_8397);
nor U8577 (N_8577,N_8294,N_8282);
xor U8578 (N_8578,N_8341,N_8247);
and U8579 (N_8579,N_8190,N_8250);
nand U8580 (N_8580,N_8101,N_8266);
xnor U8581 (N_8581,N_8257,N_8291);
xnor U8582 (N_8582,N_8396,N_8380);
nor U8583 (N_8583,N_8138,N_8224);
or U8584 (N_8584,N_8158,N_8202);
and U8585 (N_8585,N_8101,N_8364);
or U8586 (N_8586,N_8163,N_8146);
nand U8587 (N_8587,N_8270,N_8256);
xor U8588 (N_8588,N_8163,N_8154);
xor U8589 (N_8589,N_8368,N_8136);
nand U8590 (N_8590,N_8342,N_8321);
and U8591 (N_8591,N_8289,N_8262);
and U8592 (N_8592,N_8193,N_8294);
nand U8593 (N_8593,N_8117,N_8125);
xnor U8594 (N_8594,N_8108,N_8371);
xor U8595 (N_8595,N_8114,N_8280);
nand U8596 (N_8596,N_8337,N_8381);
or U8597 (N_8597,N_8207,N_8283);
xor U8598 (N_8598,N_8238,N_8341);
xnor U8599 (N_8599,N_8280,N_8251);
xnor U8600 (N_8600,N_8296,N_8237);
and U8601 (N_8601,N_8122,N_8270);
and U8602 (N_8602,N_8397,N_8119);
nor U8603 (N_8603,N_8339,N_8234);
and U8604 (N_8604,N_8327,N_8283);
and U8605 (N_8605,N_8243,N_8182);
nand U8606 (N_8606,N_8140,N_8258);
nor U8607 (N_8607,N_8116,N_8381);
or U8608 (N_8608,N_8157,N_8379);
xor U8609 (N_8609,N_8317,N_8209);
xor U8610 (N_8610,N_8110,N_8356);
nand U8611 (N_8611,N_8132,N_8133);
or U8612 (N_8612,N_8360,N_8285);
nand U8613 (N_8613,N_8207,N_8308);
xor U8614 (N_8614,N_8280,N_8255);
and U8615 (N_8615,N_8111,N_8175);
xor U8616 (N_8616,N_8261,N_8333);
or U8617 (N_8617,N_8299,N_8103);
or U8618 (N_8618,N_8356,N_8147);
nand U8619 (N_8619,N_8178,N_8118);
nor U8620 (N_8620,N_8167,N_8290);
and U8621 (N_8621,N_8297,N_8203);
and U8622 (N_8622,N_8380,N_8291);
xor U8623 (N_8623,N_8209,N_8352);
nand U8624 (N_8624,N_8209,N_8253);
or U8625 (N_8625,N_8388,N_8196);
nor U8626 (N_8626,N_8354,N_8244);
and U8627 (N_8627,N_8109,N_8326);
xor U8628 (N_8628,N_8368,N_8375);
xor U8629 (N_8629,N_8111,N_8202);
or U8630 (N_8630,N_8175,N_8346);
nor U8631 (N_8631,N_8243,N_8111);
nand U8632 (N_8632,N_8343,N_8225);
nand U8633 (N_8633,N_8169,N_8251);
and U8634 (N_8634,N_8136,N_8372);
nand U8635 (N_8635,N_8181,N_8306);
nand U8636 (N_8636,N_8284,N_8175);
and U8637 (N_8637,N_8166,N_8188);
nor U8638 (N_8638,N_8235,N_8129);
nand U8639 (N_8639,N_8184,N_8130);
and U8640 (N_8640,N_8142,N_8259);
and U8641 (N_8641,N_8215,N_8268);
or U8642 (N_8642,N_8272,N_8231);
nor U8643 (N_8643,N_8270,N_8370);
nor U8644 (N_8644,N_8195,N_8296);
and U8645 (N_8645,N_8215,N_8227);
nor U8646 (N_8646,N_8178,N_8197);
nor U8647 (N_8647,N_8181,N_8141);
nand U8648 (N_8648,N_8322,N_8195);
nand U8649 (N_8649,N_8190,N_8134);
and U8650 (N_8650,N_8384,N_8122);
nor U8651 (N_8651,N_8180,N_8216);
or U8652 (N_8652,N_8360,N_8315);
and U8653 (N_8653,N_8226,N_8107);
xor U8654 (N_8654,N_8148,N_8109);
nand U8655 (N_8655,N_8229,N_8231);
nor U8656 (N_8656,N_8220,N_8223);
nand U8657 (N_8657,N_8394,N_8356);
or U8658 (N_8658,N_8291,N_8253);
nor U8659 (N_8659,N_8346,N_8234);
nand U8660 (N_8660,N_8163,N_8176);
xor U8661 (N_8661,N_8360,N_8251);
nor U8662 (N_8662,N_8104,N_8373);
xor U8663 (N_8663,N_8331,N_8181);
nor U8664 (N_8664,N_8178,N_8233);
and U8665 (N_8665,N_8301,N_8246);
and U8666 (N_8666,N_8392,N_8195);
nor U8667 (N_8667,N_8235,N_8170);
nand U8668 (N_8668,N_8351,N_8125);
nand U8669 (N_8669,N_8194,N_8330);
nor U8670 (N_8670,N_8333,N_8141);
nand U8671 (N_8671,N_8109,N_8272);
nor U8672 (N_8672,N_8107,N_8255);
xnor U8673 (N_8673,N_8232,N_8136);
or U8674 (N_8674,N_8276,N_8244);
nand U8675 (N_8675,N_8379,N_8329);
nor U8676 (N_8676,N_8211,N_8218);
and U8677 (N_8677,N_8249,N_8369);
nor U8678 (N_8678,N_8239,N_8124);
or U8679 (N_8679,N_8199,N_8388);
nor U8680 (N_8680,N_8228,N_8223);
and U8681 (N_8681,N_8134,N_8398);
or U8682 (N_8682,N_8362,N_8342);
nand U8683 (N_8683,N_8367,N_8166);
nor U8684 (N_8684,N_8211,N_8302);
or U8685 (N_8685,N_8309,N_8150);
or U8686 (N_8686,N_8356,N_8163);
nand U8687 (N_8687,N_8285,N_8112);
xor U8688 (N_8688,N_8191,N_8358);
and U8689 (N_8689,N_8278,N_8357);
nand U8690 (N_8690,N_8318,N_8304);
xor U8691 (N_8691,N_8362,N_8117);
nor U8692 (N_8692,N_8203,N_8138);
nand U8693 (N_8693,N_8153,N_8382);
and U8694 (N_8694,N_8154,N_8274);
or U8695 (N_8695,N_8305,N_8360);
nand U8696 (N_8696,N_8122,N_8365);
xor U8697 (N_8697,N_8369,N_8338);
or U8698 (N_8698,N_8197,N_8200);
or U8699 (N_8699,N_8372,N_8289);
or U8700 (N_8700,N_8680,N_8558);
nor U8701 (N_8701,N_8634,N_8505);
nor U8702 (N_8702,N_8688,N_8522);
nor U8703 (N_8703,N_8670,N_8439);
nor U8704 (N_8704,N_8521,N_8659);
xor U8705 (N_8705,N_8466,N_8420);
xor U8706 (N_8706,N_8646,N_8638);
and U8707 (N_8707,N_8470,N_8464);
and U8708 (N_8708,N_8413,N_8624);
nor U8709 (N_8709,N_8673,N_8555);
nand U8710 (N_8710,N_8510,N_8430);
nand U8711 (N_8711,N_8529,N_8553);
nand U8712 (N_8712,N_8465,N_8407);
and U8713 (N_8713,N_8656,N_8660);
nand U8714 (N_8714,N_8604,N_8691);
nor U8715 (N_8715,N_8674,N_8663);
xor U8716 (N_8716,N_8435,N_8473);
or U8717 (N_8717,N_8643,N_8491);
nor U8718 (N_8718,N_8667,N_8446);
xor U8719 (N_8719,N_8409,N_8530);
nor U8720 (N_8720,N_8497,N_8597);
nand U8721 (N_8721,N_8488,N_8619);
or U8722 (N_8722,N_8697,N_8645);
nor U8723 (N_8723,N_8426,N_8432);
xor U8724 (N_8724,N_8441,N_8600);
nand U8725 (N_8725,N_8566,N_8574);
and U8726 (N_8726,N_8481,N_8467);
xnor U8727 (N_8727,N_8605,N_8507);
nand U8728 (N_8728,N_8572,N_8516);
and U8729 (N_8729,N_8696,N_8588);
and U8730 (N_8730,N_8622,N_8463);
xor U8731 (N_8731,N_8649,N_8581);
xnor U8732 (N_8732,N_8436,N_8445);
xnor U8733 (N_8733,N_8517,N_8564);
and U8734 (N_8734,N_8559,N_8595);
nand U8735 (N_8735,N_8582,N_8616);
nor U8736 (N_8736,N_8698,N_8583);
or U8737 (N_8737,N_8661,N_8414);
nand U8738 (N_8738,N_8613,N_8552);
xor U8739 (N_8739,N_8550,N_8669);
and U8740 (N_8740,N_8603,N_8568);
nand U8741 (N_8741,N_8617,N_8417);
and U8742 (N_8742,N_8535,N_8614);
and U8743 (N_8743,N_8524,N_8422);
or U8744 (N_8744,N_8694,N_8699);
xor U8745 (N_8745,N_8685,N_8458);
nor U8746 (N_8746,N_8450,N_8533);
nor U8747 (N_8747,N_8448,N_8684);
and U8748 (N_8748,N_8665,N_8653);
and U8749 (N_8749,N_8615,N_8443);
xor U8750 (N_8750,N_8562,N_8455);
nand U8751 (N_8751,N_8472,N_8598);
xnor U8752 (N_8752,N_8630,N_8502);
nor U8753 (N_8753,N_8462,N_8585);
nand U8754 (N_8754,N_8531,N_8456);
or U8755 (N_8755,N_8644,N_8449);
or U8756 (N_8756,N_8547,N_8418);
and U8757 (N_8757,N_8654,N_8518);
xor U8758 (N_8758,N_8639,N_8536);
nor U8759 (N_8759,N_8628,N_8438);
and U8760 (N_8760,N_8612,N_8411);
nor U8761 (N_8761,N_8623,N_8658);
nor U8762 (N_8762,N_8403,N_8423);
nor U8763 (N_8763,N_8678,N_8651);
and U8764 (N_8764,N_8546,N_8541);
xnor U8765 (N_8765,N_8608,N_8592);
or U8766 (N_8766,N_8416,N_8548);
and U8767 (N_8767,N_8693,N_8631);
nor U8768 (N_8768,N_8509,N_8542);
and U8769 (N_8769,N_8484,N_8650);
or U8770 (N_8770,N_8537,N_8493);
and U8771 (N_8771,N_8561,N_8679);
nand U8772 (N_8772,N_8668,N_8591);
nor U8773 (N_8773,N_8457,N_8690);
nand U8774 (N_8774,N_8499,N_8508);
or U8775 (N_8775,N_8586,N_8440);
xnor U8776 (N_8776,N_8557,N_8618);
xnor U8777 (N_8777,N_8611,N_8675);
and U8778 (N_8778,N_8621,N_8512);
and U8779 (N_8779,N_8648,N_8433);
nand U8780 (N_8780,N_8666,N_8607);
nor U8781 (N_8781,N_8496,N_8682);
or U8782 (N_8782,N_8402,N_8534);
and U8783 (N_8783,N_8429,N_8543);
and U8784 (N_8784,N_8601,N_8434);
and U8785 (N_8785,N_8408,N_8571);
xnor U8786 (N_8786,N_8442,N_8410);
nor U8787 (N_8787,N_8695,N_8655);
and U8788 (N_8788,N_8672,N_8652);
nand U8789 (N_8789,N_8683,N_8635);
nor U8790 (N_8790,N_8437,N_8689);
nor U8791 (N_8791,N_8578,N_8627);
xor U8792 (N_8792,N_8515,N_8573);
and U8793 (N_8793,N_8589,N_8584);
xor U8794 (N_8794,N_8478,N_8474);
nand U8795 (N_8795,N_8647,N_8560);
or U8796 (N_8796,N_8480,N_8453);
xnor U8797 (N_8797,N_8587,N_8594);
and U8798 (N_8798,N_8477,N_8479);
xnor U8799 (N_8799,N_8640,N_8610);
and U8800 (N_8800,N_8527,N_8528);
nand U8801 (N_8801,N_8451,N_8482);
nand U8802 (N_8802,N_8545,N_8520);
or U8803 (N_8803,N_8539,N_8540);
and U8804 (N_8804,N_8506,N_8662);
xnor U8805 (N_8805,N_8580,N_8428);
nor U8806 (N_8806,N_8483,N_8492);
nor U8807 (N_8807,N_8569,N_8565);
nand U8808 (N_8808,N_8625,N_8406);
xnor U8809 (N_8809,N_8503,N_8425);
or U8810 (N_8810,N_8419,N_8526);
nor U8811 (N_8811,N_8489,N_8620);
nand U8812 (N_8812,N_8447,N_8570);
nor U8813 (N_8813,N_8551,N_8421);
nand U8814 (N_8814,N_8664,N_8461);
xor U8815 (N_8815,N_8641,N_8642);
nand U8816 (N_8816,N_8415,N_8401);
or U8817 (N_8817,N_8487,N_8544);
or U8818 (N_8818,N_8538,N_8476);
nand U8819 (N_8819,N_8686,N_8692);
nand U8820 (N_8820,N_8459,N_8677);
nand U8821 (N_8821,N_8475,N_8579);
and U8822 (N_8822,N_8405,N_8556);
nand U8823 (N_8823,N_8498,N_8412);
or U8824 (N_8824,N_8687,N_8404);
or U8825 (N_8825,N_8444,N_8532);
and U8826 (N_8826,N_8632,N_8563);
and U8827 (N_8827,N_8486,N_8454);
and U8828 (N_8828,N_8554,N_8523);
xor U8829 (N_8829,N_8513,N_8494);
nor U8830 (N_8830,N_8460,N_8427);
xnor U8831 (N_8831,N_8495,N_8525);
nand U8832 (N_8832,N_8471,N_8590);
xor U8833 (N_8833,N_8511,N_8504);
xnor U8834 (N_8834,N_8577,N_8567);
and U8835 (N_8835,N_8633,N_8671);
or U8836 (N_8836,N_8424,N_8637);
nor U8837 (N_8837,N_8490,N_8609);
nor U8838 (N_8838,N_8602,N_8593);
or U8839 (N_8839,N_8596,N_8469);
nand U8840 (N_8840,N_8519,N_8599);
xor U8841 (N_8841,N_8452,N_8636);
and U8842 (N_8842,N_8676,N_8606);
and U8843 (N_8843,N_8431,N_8468);
xnor U8844 (N_8844,N_8549,N_8485);
or U8845 (N_8845,N_8575,N_8514);
and U8846 (N_8846,N_8657,N_8576);
or U8847 (N_8847,N_8400,N_8500);
nand U8848 (N_8848,N_8626,N_8501);
nor U8849 (N_8849,N_8629,N_8681);
and U8850 (N_8850,N_8403,N_8638);
xor U8851 (N_8851,N_8635,N_8569);
xnor U8852 (N_8852,N_8683,N_8506);
or U8853 (N_8853,N_8543,N_8546);
and U8854 (N_8854,N_8507,N_8430);
or U8855 (N_8855,N_8559,N_8488);
and U8856 (N_8856,N_8556,N_8458);
nor U8857 (N_8857,N_8586,N_8646);
or U8858 (N_8858,N_8577,N_8672);
xor U8859 (N_8859,N_8549,N_8550);
nor U8860 (N_8860,N_8585,N_8483);
and U8861 (N_8861,N_8646,N_8653);
xnor U8862 (N_8862,N_8515,N_8448);
or U8863 (N_8863,N_8546,N_8419);
and U8864 (N_8864,N_8407,N_8644);
nor U8865 (N_8865,N_8585,N_8480);
nor U8866 (N_8866,N_8607,N_8463);
or U8867 (N_8867,N_8541,N_8650);
nand U8868 (N_8868,N_8433,N_8621);
or U8869 (N_8869,N_8550,N_8463);
and U8870 (N_8870,N_8422,N_8690);
and U8871 (N_8871,N_8649,N_8463);
and U8872 (N_8872,N_8570,N_8622);
and U8873 (N_8873,N_8422,N_8510);
nand U8874 (N_8874,N_8579,N_8531);
xnor U8875 (N_8875,N_8595,N_8495);
nand U8876 (N_8876,N_8458,N_8652);
nor U8877 (N_8877,N_8405,N_8534);
nor U8878 (N_8878,N_8448,N_8508);
and U8879 (N_8879,N_8457,N_8618);
nor U8880 (N_8880,N_8664,N_8494);
or U8881 (N_8881,N_8412,N_8441);
or U8882 (N_8882,N_8682,N_8643);
or U8883 (N_8883,N_8571,N_8665);
xor U8884 (N_8884,N_8529,N_8670);
xor U8885 (N_8885,N_8457,N_8567);
and U8886 (N_8886,N_8570,N_8676);
xnor U8887 (N_8887,N_8432,N_8577);
nand U8888 (N_8888,N_8631,N_8492);
xor U8889 (N_8889,N_8649,N_8545);
nand U8890 (N_8890,N_8595,N_8459);
or U8891 (N_8891,N_8624,N_8482);
and U8892 (N_8892,N_8601,N_8495);
nand U8893 (N_8893,N_8467,N_8598);
xor U8894 (N_8894,N_8528,N_8661);
xor U8895 (N_8895,N_8554,N_8638);
or U8896 (N_8896,N_8545,N_8424);
nor U8897 (N_8897,N_8645,N_8666);
nand U8898 (N_8898,N_8486,N_8424);
nor U8899 (N_8899,N_8695,N_8605);
or U8900 (N_8900,N_8642,N_8499);
nor U8901 (N_8901,N_8433,N_8431);
xor U8902 (N_8902,N_8403,N_8450);
and U8903 (N_8903,N_8671,N_8538);
or U8904 (N_8904,N_8625,N_8639);
nor U8905 (N_8905,N_8432,N_8584);
xor U8906 (N_8906,N_8564,N_8654);
or U8907 (N_8907,N_8447,N_8561);
nor U8908 (N_8908,N_8525,N_8685);
or U8909 (N_8909,N_8437,N_8588);
or U8910 (N_8910,N_8652,N_8497);
nor U8911 (N_8911,N_8406,N_8695);
and U8912 (N_8912,N_8503,N_8477);
nand U8913 (N_8913,N_8411,N_8685);
and U8914 (N_8914,N_8424,N_8613);
xnor U8915 (N_8915,N_8602,N_8662);
nor U8916 (N_8916,N_8540,N_8589);
or U8917 (N_8917,N_8605,N_8454);
and U8918 (N_8918,N_8597,N_8668);
or U8919 (N_8919,N_8496,N_8469);
or U8920 (N_8920,N_8680,N_8661);
and U8921 (N_8921,N_8571,N_8622);
xnor U8922 (N_8922,N_8674,N_8540);
nand U8923 (N_8923,N_8411,N_8686);
nor U8924 (N_8924,N_8404,N_8486);
nor U8925 (N_8925,N_8684,N_8537);
and U8926 (N_8926,N_8538,N_8576);
and U8927 (N_8927,N_8631,N_8412);
or U8928 (N_8928,N_8691,N_8567);
nand U8929 (N_8929,N_8436,N_8692);
nor U8930 (N_8930,N_8587,N_8592);
xor U8931 (N_8931,N_8662,N_8465);
nand U8932 (N_8932,N_8401,N_8649);
xnor U8933 (N_8933,N_8579,N_8580);
nand U8934 (N_8934,N_8428,N_8485);
nor U8935 (N_8935,N_8465,N_8535);
nor U8936 (N_8936,N_8683,N_8520);
or U8937 (N_8937,N_8484,N_8666);
nand U8938 (N_8938,N_8665,N_8560);
or U8939 (N_8939,N_8678,N_8625);
and U8940 (N_8940,N_8492,N_8695);
and U8941 (N_8941,N_8485,N_8661);
or U8942 (N_8942,N_8421,N_8538);
nand U8943 (N_8943,N_8577,N_8548);
or U8944 (N_8944,N_8619,N_8676);
and U8945 (N_8945,N_8624,N_8429);
nand U8946 (N_8946,N_8606,N_8462);
and U8947 (N_8947,N_8492,N_8607);
nor U8948 (N_8948,N_8579,N_8487);
nand U8949 (N_8949,N_8460,N_8504);
and U8950 (N_8950,N_8621,N_8615);
xnor U8951 (N_8951,N_8581,N_8588);
nor U8952 (N_8952,N_8423,N_8515);
nand U8953 (N_8953,N_8576,N_8601);
xnor U8954 (N_8954,N_8525,N_8578);
or U8955 (N_8955,N_8441,N_8456);
nor U8956 (N_8956,N_8614,N_8580);
nor U8957 (N_8957,N_8492,N_8449);
nor U8958 (N_8958,N_8539,N_8480);
and U8959 (N_8959,N_8640,N_8450);
xor U8960 (N_8960,N_8650,N_8596);
nand U8961 (N_8961,N_8435,N_8536);
nand U8962 (N_8962,N_8429,N_8510);
or U8963 (N_8963,N_8612,N_8577);
xnor U8964 (N_8964,N_8599,N_8468);
xnor U8965 (N_8965,N_8517,N_8498);
or U8966 (N_8966,N_8660,N_8511);
and U8967 (N_8967,N_8690,N_8580);
and U8968 (N_8968,N_8680,N_8484);
and U8969 (N_8969,N_8428,N_8607);
nor U8970 (N_8970,N_8461,N_8646);
nand U8971 (N_8971,N_8404,N_8437);
and U8972 (N_8972,N_8427,N_8669);
and U8973 (N_8973,N_8498,N_8521);
or U8974 (N_8974,N_8449,N_8443);
and U8975 (N_8975,N_8528,N_8543);
nor U8976 (N_8976,N_8517,N_8641);
nor U8977 (N_8977,N_8512,N_8525);
or U8978 (N_8978,N_8471,N_8689);
and U8979 (N_8979,N_8577,N_8690);
nor U8980 (N_8980,N_8484,N_8597);
or U8981 (N_8981,N_8660,N_8586);
and U8982 (N_8982,N_8552,N_8640);
xor U8983 (N_8983,N_8445,N_8582);
nor U8984 (N_8984,N_8406,N_8411);
xnor U8985 (N_8985,N_8529,N_8548);
and U8986 (N_8986,N_8685,N_8660);
and U8987 (N_8987,N_8490,N_8697);
or U8988 (N_8988,N_8535,N_8658);
nand U8989 (N_8989,N_8616,N_8656);
or U8990 (N_8990,N_8556,N_8693);
xnor U8991 (N_8991,N_8515,N_8642);
xnor U8992 (N_8992,N_8639,N_8520);
or U8993 (N_8993,N_8505,N_8424);
or U8994 (N_8994,N_8688,N_8444);
nand U8995 (N_8995,N_8444,N_8662);
nand U8996 (N_8996,N_8689,N_8446);
xor U8997 (N_8997,N_8526,N_8662);
nand U8998 (N_8998,N_8624,N_8699);
xor U8999 (N_8999,N_8401,N_8692);
and U9000 (N_9000,N_8988,N_8989);
or U9001 (N_9001,N_8879,N_8833);
xnor U9002 (N_9002,N_8724,N_8710);
nand U9003 (N_9003,N_8828,N_8939);
and U9004 (N_9004,N_8757,N_8764);
and U9005 (N_9005,N_8995,N_8932);
nor U9006 (N_9006,N_8908,N_8812);
nand U9007 (N_9007,N_8743,N_8755);
or U9008 (N_9008,N_8865,N_8918);
nor U9009 (N_9009,N_8930,N_8745);
and U9010 (N_9010,N_8984,N_8844);
or U9011 (N_9011,N_8837,N_8907);
nand U9012 (N_9012,N_8901,N_8974);
and U9013 (N_9013,N_8871,N_8813);
nor U9014 (N_9014,N_8866,N_8840);
xnor U9015 (N_9015,N_8778,N_8889);
nor U9016 (N_9016,N_8963,N_8718);
and U9017 (N_9017,N_8872,N_8969);
or U9018 (N_9018,N_8835,N_8985);
or U9019 (N_9019,N_8714,N_8888);
nor U9020 (N_9020,N_8912,N_8773);
or U9021 (N_9021,N_8829,N_8736);
nand U9022 (N_9022,N_8702,N_8964);
and U9023 (N_9023,N_8793,N_8784);
xor U9024 (N_9024,N_8852,N_8945);
xor U9025 (N_9025,N_8876,N_8786);
nand U9026 (N_9026,N_8892,N_8823);
nand U9027 (N_9027,N_8982,N_8931);
and U9028 (N_9028,N_8814,N_8853);
xnor U9029 (N_9029,N_8781,N_8794);
and U9030 (N_9030,N_8747,N_8834);
and U9031 (N_9031,N_8796,N_8763);
nand U9032 (N_9032,N_8961,N_8787);
or U9033 (N_9033,N_8864,N_8848);
nor U9034 (N_9034,N_8877,N_8999);
or U9035 (N_9035,N_8821,N_8845);
and U9036 (N_9036,N_8830,N_8751);
nor U9037 (N_9037,N_8952,N_8700);
nand U9038 (N_9038,N_8972,N_8949);
xor U9039 (N_9039,N_8849,N_8775);
xor U9040 (N_9040,N_8933,N_8774);
and U9041 (N_9041,N_8827,N_8959);
xnor U9042 (N_9042,N_8976,N_8809);
nor U9043 (N_9043,N_8869,N_8723);
and U9044 (N_9044,N_8944,N_8779);
nor U9045 (N_9045,N_8818,N_8749);
or U9046 (N_9046,N_8756,N_8929);
or U9047 (N_9047,N_8896,N_8922);
nor U9048 (N_9048,N_8968,N_8859);
xnor U9049 (N_9049,N_8948,N_8752);
or U9050 (N_9050,N_8758,N_8903);
nor U9051 (N_9051,N_8916,N_8785);
or U9052 (N_9052,N_8734,N_8898);
nor U9053 (N_9053,N_8966,N_8767);
xnor U9054 (N_9054,N_8762,N_8973);
xnor U9055 (N_9055,N_8719,N_8937);
or U9056 (N_9056,N_8725,N_8788);
and U9057 (N_9057,N_8867,N_8811);
nor U9058 (N_9058,N_8970,N_8727);
nand U9059 (N_9059,N_8816,N_8981);
or U9060 (N_9060,N_8983,N_8957);
and U9061 (N_9061,N_8824,N_8847);
nor U9062 (N_9062,N_8986,N_8706);
xor U9063 (N_9063,N_8910,N_8776);
nor U9064 (N_9064,N_8717,N_8769);
xnor U9065 (N_9065,N_8920,N_8790);
nand U9066 (N_9066,N_8921,N_8800);
and U9067 (N_9067,N_8902,N_8807);
and U9068 (N_9068,N_8713,N_8777);
or U9069 (N_9069,N_8791,N_8941);
and U9070 (N_9070,N_8860,N_8906);
nand U9071 (N_9071,N_8815,N_8801);
or U9072 (N_9072,N_8950,N_8768);
nand U9073 (N_9073,N_8819,N_8861);
nand U9074 (N_9074,N_8942,N_8881);
or U9075 (N_9075,N_8917,N_8980);
nand U9076 (N_9076,N_8956,N_8810);
xnor U9077 (N_9077,N_8730,N_8737);
xor U9078 (N_9078,N_8943,N_8975);
xor U9079 (N_9079,N_8895,N_8946);
xnor U9080 (N_9080,N_8708,N_8978);
nand U9081 (N_9081,N_8760,N_8803);
nand U9082 (N_9082,N_8971,N_8862);
nor U9083 (N_9083,N_8928,N_8831);
nand U9084 (N_9084,N_8897,N_8856);
nand U9085 (N_9085,N_8741,N_8765);
xnor U9086 (N_9086,N_8750,N_8780);
nand U9087 (N_9087,N_8890,N_8887);
or U9088 (N_9088,N_8919,N_8936);
and U9089 (N_9089,N_8893,N_8891);
xor U9090 (N_9090,N_8802,N_8965);
xor U9091 (N_9091,N_8934,N_8817);
xor U9092 (N_9092,N_8716,N_8863);
or U9093 (N_9093,N_8720,N_8924);
or U9094 (N_9094,N_8729,N_8820);
xnor U9095 (N_9095,N_8799,N_8742);
xor U9096 (N_9096,N_8739,N_8977);
xnor U9097 (N_9097,N_8868,N_8954);
nor U9098 (N_9098,N_8870,N_8962);
nand U9099 (N_9099,N_8836,N_8772);
xnor U9100 (N_9100,N_8766,N_8707);
and U9101 (N_9101,N_8992,N_8955);
and U9102 (N_9102,N_8875,N_8997);
xnor U9103 (N_9103,N_8987,N_8940);
or U9104 (N_9104,N_8843,N_8996);
and U9105 (N_9105,N_8880,N_8873);
or U9106 (N_9106,N_8926,N_8740);
nor U9107 (N_9107,N_8909,N_8857);
or U9108 (N_9108,N_8754,N_8792);
nor U9109 (N_9109,N_8771,N_8947);
or U9110 (N_9110,N_8722,N_8967);
nor U9111 (N_9111,N_8846,N_8770);
nor U9112 (N_9112,N_8735,N_8855);
and U9113 (N_9113,N_8782,N_8858);
nor U9114 (N_9114,N_8884,N_8826);
nor U9115 (N_9115,N_8728,N_8991);
and U9116 (N_9116,N_8854,N_8994);
nand U9117 (N_9117,N_8732,N_8753);
or U9118 (N_9118,N_8905,N_8808);
or U9119 (N_9119,N_8904,N_8721);
and U9120 (N_9120,N_8715,N_8915);
xnor U9121 (N_9121,N_8759,N_8705);
nor U9122 (N_9122,N_8838,N_8701);
and U9123 (N_9123,N_8797,N_8703);
nand U9124 (N_9124,N_8738,N_8850);
or U9125 (N_9125,N_8899,N_8806);
or U9126 (N_9126,N_8874,N_8979);
nand U9127 (N_9127,N_8733,N_8958);
nand U9128 (N_9128,N_8804,N_8894);
xnor U9129 (N_9129,N_8711,N_8746);
nand U9130 (N_9130,N_8842,N_8709);
and U9131 (N_9131,N_8748,N_8832);
nor U9132 (N_9132,N_8990,N_8825);
and U9133 (N_9133,N_8878,N_8911);
nand U9134 (N_9134,N_8885,N_8923);
or U9135 (N_9135,N_8914,N_8935);
xnor U9136 (N_9136,N_8886,N_8925);
or U9137 (N_9137,N_8960,N_8726);
xnor U9138 (N_9138,N_8883,N_8798);
and U9139 (N_9139,N_8882,N_8822);
and U9140 (N_9140,N_8953,N_8761);
nand U9141 (N_9141,N_8795,N_8927);
or U9142 (N_9142,N_8731,N_8938);
and U9143 (N_9143,N_8841,N_8900);
nand U9144 (N_9144,N_8789,N_8744);
and U9145 (N_9145,N_8913,N_8712);
xnor U9146 (N_9146,N_8951,N_8851);
nand U9147 (N_9147,N_8993,N_8704);
or U9148 (N_9148,N_8783,N_8998);
xor U9149 (N_9149,N_8839,N_8805);
nor U9150 (N_9150,N_8949,N_8780);
or U9151 (N_9151,N_8762,N_8849);
or U9152 (N_9152,N_8928,N_8838);
nor U9153 (N_9153,N_8774,N_8777);
or U9154 (N_9154,N_8795,N_8964);
or U9155 (N_9155,N_8923,N_8880);
xor U9156 (N_9156,N_8908,N_8801);
xor U9157 (N_9157,N_8821,N_8887);
nand U9158 (N_9158,N_8950,N_8796);
xor U9159 (N_9159,N_8898,N_8855);
or U9160 (N_9160,N_8785,N_8900);
or U9161 (N_9161,N_8842,N_8782);
and U9162 (N_9162,N_8721,N_8801);
xor U9163 (N_9163,N_8878,N_8750);
nor U9164 (N_9164,N_8880,N_8912);
nand U9165 (N_9165,N_8954,N_8816);
or U9166 (N_9166,N_8870,N_8764);
or U9167 (N_9167,N_8877,N_8906);
nor U9168 (N_9168,N_8875,N_8725);
nor U9169 (N_9169,N_8989,N_8818);
nand U9170 (N_9170,N_8863,N_8807);
xnor U9171 (N_9171,N_8951,N_8981);
nand U9172 (N_9172,N_8751,N_8967);
xnor U9173 (N_9173,N_8897,N_8794);
or U9174 (N_9174,N_8718,N_8776);
nand U9175 (N_9175,N_8941,N_8871);
and U9176 (N_9176,N_8743,N_8846);
and U9177 (N_9177,N_8955,N_8786);
xnor U9178 (N_9178,N_8716,N_8925);
and U9179 (N_9179,N_8933,N_8764);
nand U9180 (N_9180,N_8760,N_8922);
nand U9181 (N_9181,N_8909,N_8715);
and U9182 (N_9182,N_8985,N_8950);
nand U9183 (N_9183,N_8978,N_8935);
xor U9184 (N_9184,N_8843,N_8831);
and U9185 (N_9185,N_8828,N_8850);
nor U9186 (N_9186,N_8717,N_8777);
and U9187 (N_9187,N_8923,N_8758);
nor U9188 (N_9188,N_8813,N_8772);
or U9189 (N_9189,N_8831,N_8827);
nand U9190 (N_9190,N_8897,N_8915);
or U9191 (N_9191,N_8736,N_8933);
and U9192 (N_9192,N_8764,N_8910);
nor U9193 (N_9193,N_8799,N_8820);
xor U9194 (N_9194,N_8773,N_8973);
and U9195 (N_9195,N_8705,N_8754);
nor U9196 (N_9196,N_8781,N_8706);
nand U9197 (N_9197,N_8817,N_8987);
nor U9198 (N_9198,N_8937,N_8963);
nand U9199 (N_9199,N_8942,N_8860);
and U9200 (N_9200,N_8961,N_8970);
and U9201 (N_9201,N_8705,N_8981);
or U9202 (N_9202,N_8852,N_8964);
and U9203 (N_9203,N_8725,N_8974);
and U9204 (N_9204,N_8926,N_8746);
nand U9205 (N_9205,N_8788,N_8966);
nor U9206 (N_9206,N_8881,N_8753);
nand U9207 (N_9207,N_8892,N_8810);
or U9208 (N_9208,N_8911,N_8946);
or U9209 (N_9209,N_8823,N_8856);
and U9210 (N_9210,N_8792,N_8853);
or U9211 (N_9211,N_8864,N_8982);
xor U9212 (N_9212,N_8741,N_8858);
nand U9213 (N_9213,N_8704,N_8873);
or U9214 (N_9214,N_8877,N_8998);
and U9215 (N_9215,N_8909,N_8755);
or U9216 (N_9216,N_8772,N_8873);
and U9217 (N_9217,N_8915,N_8979);
and U9218 (N_9218,N_8787,N_8861);
or U9219 (N_9219,N_8981,N_8896);
and U9220 (N_9220,N_8998,N_8981);
nand U9221 (N_9221,N_8908,N_8740);
and U9222 (N_9222,N_8811,N_8776);
nor U9223 (N_9223,N_8946,N_8831);
xor U9224 (N_9224,N_8718,N_8858);
or U9225 (N_9225,N_8802,N_8869);
xnor U9226 (N_9226,N_8780,N_8768);
nor U9227 (N_9227,N_8847,N_8700);
and U9228 (N_9228,N_8765,N_8846);
nor U9229 (N_9229,N_8889,N_8725);
or U9230 (N_9230,N_8975,N_8714);
and U9231 (N_9231,N_8935,N_8843);
xor U9232 (N_9232,N_8736,N_8930);
xor U9233 (N_9233,N_8998,N_8916);
and U9234 (N_9234,N_8786,N_8775);
nand U9235 (N_9235,N_8867,N_8774);
and U9236 (N_9236,N_8877,N_8727);
nor U9237 (N_9237,N_8900,N_8986);
nand U9238 (N_9238,N_8737,N_8998);
nor U9239 (N_9239,N_8974,N_8742);
nand U9240 (N_9240,N_8841,N_8736);
nand U9241 (N_9241,N_8779,N_8967);
xnor U9242 (N_9242,N_8806,N_8991);
or U9243 (N_9243,N_8713,N_8793);
nand U9244 (N_9244,N_8897,N_8896);
or U9245 (N_9245,N_8759,N_8893);
or U9246 (N_9246,N_8856,N_8916);
nor U9247 (N_9247,N_8741,N_8900);
or U9248 (N_9248,N_8951,N_8718);
nor U9249 (N_9249,N_8901,N_8848);
nand U9250 (N_9250,N_8838,N_8780);
xor U9251 (N_9251,N_8959,N_8965);
nor U9252 (N_9252,N_8724,N_8827);
nor U9253 (N_9253,N_8740,N_8911);
nor U9254 (N_9254,N_8784,N_8997);
and U9255 (N_9255,N_8725,N_8736);
and U9256 (N_9256,N_8741,N_8714);
xnor U9257 (N_9257,N_8901,N_8916);
nand U9258 (N_9258,N_8770,N_8898);
xnor U9259 (N_9259,N_8877,N_8863);
or U9260 (N_9260,N_8750,N_8711);
xnor U9261 (N_9261,N_8874,N_8763);
nand U9262 (N_9262,N_8728,N_8810);
or U9263 (N_9263,N_8752,N_8741);
or U9264 (N_9264,N_8901,N_8703);
and U9265 (N_9265,N_8996,N_8985);
and U9266 (N_9266,N_8724,N_8971);
or U9267 (N_9267,N_8921,N_8734);
xor U9268 (N_9268,N_8851,N_8750);
nand U9269 (N_9269,N_8845,N_8853);
and U9270 (N_9270,N_8878,N_8945);
and U9271 (N_9271,N_8954,N_8846);
xnor U9272 (N_9272,N_8850,N_8830);
and U9273 (N_9273,N_8861,N_8829);
xnor U9274 (N_9274,N_8700,N_8736);
nor U9275 (N_9275,N_8717,N_8861);
nand U9276 (N_9276,N_8886,N_8910);
nand U9277 (N_9277,N_8907,N_8720);
or U9278 (N_9278,N_8990,N_8743);
xnor U9279 (N_9279,N_8791,N_8934);
and U9280 (N_9280,N_8878,N_8704);
xor U9281 (N_9281,N_8802,N_8771);
or U9282 (N_9282,N_8766,N_8781);
or U9283 (N_9283,N_8771,N_8893);
and U9284 (N_9284,N_8924,N_8983);
or U9285 (N_9285,N_8786,N_8982);
nor U9286 (N_9286,N_8977,N_8882);
nand U9287 (N_9287,N_8748,N_8758);
nor U9288 (N_9288,N_8709,N_8710);
nand U9289 (N_9289,N_8957,N_8730);
nand U9290 (N_9290,N_8979,N_8787);
nand U9291 (N_9291,N_8912,N_8837);
nand U9292 (N_9292,N_8809,N_8874);
xor U9293 (N_9293,N_8946,N_8881);
nand U9294 (N_9294,N_8858,N_8719);
or U9295 (N_9295,N_8834,N_8823);
and U9296 (N_9296,N_8966,N_8927);
xnor U9297 (N_9297,N_8707,N_8768);
or U9298 (N_9298,N_8980,N_8793);
and U9299 (N_9299,N_8867,N_8767);
nand U9300 (N_9300,N_9124,N_9033);
or U9301 (N_9301,N_9254,N_9178);
nand U9302 (N_9302,N_9245,N_9247);
or U9303 (N_9303,N_9085,N_9070);
nand U9304 (N_9304,N_9134,N_9021);
and U9305 (N_9305,N_9128,N_9189);
and U9306 (N_9306,N_9282,N_9286);
and U9307 (N_9307,N_9080,N_9115);
xnor U9308 (N_9308,N_9154,N_9159);
or U9309 (N_9309,N_9067,N_9288);
or U9310 (N_9310,N_9161,N_9212);
xnor U9311 (N_9311,N_9275,N_9280);
and U9312 (N_9312,N_9294,N_9056);
and U9313 (N_9313,N_9179,N_9263);
or U9314 (N_9314,N_9290,N_9100);
and U9315 (N_9315,N_9277,N_9057);
xnor U9316 (N_9316,N_9034,N_9051);
xnor U9317 (N_9317,N_9127,N_9299);
or U9318 (N_9318,N_9158,N_9096);
nand U9319 (N_9319,N_9196,N_9058);
nand U9320 (N_9320,N_9191,N_9145);
nand U9321 (N_9321,N_9129,N_9244);
and U9322 (N_9322,N_9004,N_9109);
and U9323 (N_9323,N_9024,N_9048);
and U9324 (N_9324,N_9227,N_9181);
xor U9325 (N_9325,N_9125,N_9172);
nor U9326 (N_9326,N_9155,N_9138);
or U9327 (N_9327,N_9182,N_9162);
nor U9328 (N_9328,N_9187,N_9010);
and U9329 (N_9329,N_9193,N_9150);
and U9330 (N_9330,N_9174,N_9169);
xor U9331 (N_9331,N_9269,N_9297);
or U9332 (N_9332,N_9040,N_9092);
and U9333 (N_9333,N_9111,N_9088);
or U9334 (N_9334,N_9079,N_9201);
nand U9335 (N_9335,N_9203,N_9052);
nor U9336 (N_9336,N_9272,N_9170);
xor U9337 (N_9337,N_9011,N_9243);
xnor U9338 (N_9338,N_9218,N_9240);
and U9339 (N_9339,N_9002,N_9241);
and U9340 (N_9340,N_9295,N_9130);
nor U9341 (N_9341,N_9166,N_9121);
nor U9342 (N_9342,N_9110,N_9032);
nand U9343 (N_9343,N_9045,N_9131);
xnor U9344 (N_9344,N_9279,N_9221);
nand U9345 (N_9345,N_9252,N_9224);
nand U9346 (N_9346,N_9207,N_9242);
nand U9347 (N_9347,N_9061,N_9098);
nand U9348 (N_9348,N_9097,N_9060);
or U9349 (N_9349,N_9255,N_9261);
or U9350 (N_9350,N_9152,N_9019);
nor U9351 (N_9351,N_9027,N_9168);
or U9352 (N_9352,N_9046,N_9013);
nor U9353 (N_9353,N_9082,N_9017);
or U9354 (N_9354,N_9005,N_9059);
xnor U9355 (N_9355,N_9190,N_9267);
nor U9356 (N_9356,N_9108,N_9090);
nand U9357 (N_9357,N_9065,N_9132);
and U9358 (N_9358,N_9153,N_9133);
nor U9359 (N_9359,N_9076,N_9236);
and U9360 (N_9360,N_9078,N_9068);
and U9361 (N_9361,N_9265,N_9177);
nand U9362 (N_9362,N_9208,N_9211);
nand U9363 (N_9363,N_9022,N_9194);
xor U9364 (N_9364,N_9106,N_9268);
xor U9365 (N_9365,N_9200,N_9120);
nand U9366 (N_9366,N_9216,N_9163);
or U9367 (N_9367,N_9081,N_9001);
or U9368 (N_9368,N_9015,N_9054);
xor U9369 (N_9369,N_9266,N_9160);
nor U9370 (N_9370,N_9285,N_9102);
or U9371 (N_9371,N_9296,N_9144);
and U9372 (N_9372,N_9149,N_9072);
xor U9373 (N_9373,N_9093,N_9050);
xnor U9374 (N_9374,N_9287,N_9273);
and U9375 (N_9375,N_9270,N_9183);
nand U9376 (N_9376,N_9123,N_9039);
xor U9377 (N_9377,N_9089,N_9043);
xor U9378 (N_9378,N_9003,N_9037);
nand U9379 (N_9379,N_9091,N_9141);
nor U9380 (N_9380,N_9206,N_9256);
and U9381 (N_9381,N_9014,N_9044);
or U9382 (N_9382,N_9104,N_9055);
xor U9383 (N_9383,N_9164,N_9074);
nor U9384 (N_9384,N_9101,N_9049);
or U9385 (N_9385,N_9210,N_9157);
nand U9386 (N_9386,N_9063,N_9007);
nor U9387 (N_9387,N_9250,N_9069);
nor U9388 (N_9388,N_9239,N_9146);
nor U9389 (N_9389,N_9235,N_9292);
nor U9390 (N_9390,N_9156,N_9142);
nor U9391 (N_9391,N_9136,N_9113);
xnor U9392 (N_9392,N_9077,N_9197);
or U9393 (N_9393,N_9249,N_9122);
or U9394 (N_9394,N_9232,N_9148);
nor U9395 (N_9395,N_9213,N_9233);
nand U9396 (N_9396,N_9281,N_9234);
xor U9397 (N_9397,N_9192,N_9000);
or U9398 (N_9398,N_9237,N_9025);
nand U9399 (N_9399,N_9259,N_9204);
nand U9400 (N_9400,N_9231,N_9176);
and U9401 (N_9401,N_9271,N_9031);
xor U9402 (N_9402,N_9165,N_9041);
xor U9403 (N_9403,N_9083,N_9180);
or U9404 (N_9404,N_9035,N_9202);
nand U9405 (N_9405,N_9095,N_9064);
and U9406 (N_9406,N_9217,N_9117);
nor U9407 (N_9407,N_9274,N_9053);
and U9408 (N_9408,N_9167,N_9228);
and U9409 (N_9409,N_9246,N_9225);
xnor U9410 (N_9410,N_9185,N_9188);
nand U9411 (N_9411,N_9278,N_9008);
or U9412 (N_9412,N_9209,N_9114);
nor U9413 (N_9413,N_9291,N_9084);
nor U9414 (N_9414,N_9086,N_9147);
or U9415 (N_9415,N_9103,N_9251);
nor U9416 (N_9416,N_9016,N_9006);
nand U9417 (N_9417,N_9253,N_9038);
xor U9418 (N_9418,N_9284,N_9298);
nor U9419 (N_9419,N_9116,N_9226);
xor U9420 (N_9420,N_9262,N_9248);
nand U9421 (N_9421,N_9293,N_9135);
xor U9422 (N_9422,N_9205,N_9030);
and U9423 (N_9423,N_9137,N_9087);
or U9424 (N_9424,N_9220,N_9173);
and U9425 (N_9425,N_9289,N_9139);
nand U9426 (N_9426,N_9184,N_9257);
nand U9427 (N_9427,N_9229,N_9042);
nor U9428 (N_9428,N_9075,N_9112);
xnor U9429 (N_9429,N_9283,N_9260);
xnor U9430 (N_9430,N_9140,N_9105);
and U9431 (N_9431,N_9028,N_9199);
nand U9432 (N_9432,N_9214,N_9276);
and U9433 (N_9433,N_9071,N_9066);
nor U9434 (N_9434,N_9107,N_9126);
or U9435 (N_9435,N_9198,N_9009);
nor U9436 (N_9436,N_9047,N_9222);
xor U9437 (N_9437,N_9026,N_9023);
and U9438 (N_9438,N_9073,N_9151);
or U9439 (N_9439,N_9119,N_9238);
nor U9440 (N_9440,N_9062,N_9143);
nand U9441 (N_9441,N_9258,N_9171);
xor U9442 (N_9442,N_9223,N_9186);
nor U9443 (N_9443,N_9020,N_9029);
or U9444 (N_9444,N_9118,N_9195);
nand U9445 (N_9445,N_9230,N_9219);
xnor U9446 (N_9446,N_9264,N_9099);
and U9447 (N_9447,N_9018,N_9036);
and U9448 (N_9448,N_9094,N_9175);
and U9449 (N_9449,N_9215,N_9012);
or U9450 (N_9450,N_9270,N_9128);
nor U9451 (N_9451,N_9164,N_9227);
nor U9452 (N_9452,N_9112,N_9183);
nand U9453 (N_9453,N_9105,N_9122);
xnor U9454 (N_9454,N_9172,N_9097);
nand U9455 (N_9455,N_9264,N_9000);
or U9456 (N_9456,N_9257,N_9209);
xnor U9457 (N_9457,N_9187,N_9181);
or U9458 (N_9458,N_9186,N_9072);
nand U9459 (N_9459,N_9179,N_9206);
and U9460 (N_9460,N_9233,N_9231);
xor U9461 (N_9461,N_9053,N_9260);
nand U9462 (N_9462,N_9038,N_9046);
and U9463 (N_9463,N_9004,N_9272);
nand U9464 (N_9464,N_9077,N_9232);
and U9465 (N_9465,N_9121,N_9026);
xnor U9466 (N_9466,N_9250,N_9210);
or U9467 (N_9467,N_9219,N_9161);
nand U9468 (N_9468,N_9059,N_9054);
nand U9469 (N_9469,N_9071,N_9288);
and U9470 (N_9470,N_9009,N_9280);
nor U9471 (N_9471,N_9067,N_9197);
nor U9472 (N_9472,N_9131,N_9256);
xor U9473 (N_9473,N_9274,N_9097);
nand U9474 (N_9474,N_9006,N_9043);
nor U9475 (N_9475,N_9167,N_9089);
and U9476 (N_9476,N_9260,N_9068);
and U9477 (N_9477,N_9174,N_9099);
nor U9478 (N_9478,N_9224,N_9258);
xor U9479 (N_9479,N_9183,N_9178);
and U9480 (N_9480,N_9079,N_9297);
xor U9481 (N_9481,N_9245,N_9125);
nand U9482 (N_9482,N_9196,N_9090);
and U9483 (N_9483,N_9127,N_9189);
and U9484 (N_9484,N_9256,N_9265);
nand U9485 (N_9485,N_9034,N_9173);
nand U9486 (N_9486,N_9013,N_9209);
nand U9487 (N_9487,N_9028,N_9263);
and U9488 (N_9488,N_9149,N_9283);
nor U9489 (N_9489,N_9239,N_9021);
xnor U9490 (N_9490,N_9214,N_9133);
and U9491 (N_9491,N_9196,N_9227);
nor U9492 (N_9492,N_9027,N_9138);
nand U9493 (N_9493,N_9008,N_9057);
nor U9494 (N_9494,N_9057,N_9290);
nand U9495 (N_9495,N_9020,N_9125);
and U9496 (N_9496,N_9188,N_9130);
nand U9497 (N_9497,N_9127,N_9216);
and U9498 (N_9498,N_9270,N_9262);
nand U9499 (N_9499,N_9067,N_9212);
nand U9500 (N_9500,N_9045,N_9203);
nand U9501 (N_9501,N_9074,N_9072);
xor U9502 (N_9502,N_9112,N_9229);
nor U9503 (N_9503,N_9265,N_9130);
xor U9504 (N_9504,N_9108,N_9131);
nor U9505 (N_9505,N_9132,N_9260);
xor U9506 (N_9506,N_9076,N_9222);
nor U9507 (N_9507,N_9154,N_9150);
xor U9508 (N_9508,N_9092,N_9183);
nand U9509 (N_9509,N_9064,N_9077);
xnor U9510 (N_9510,N_9014,N_9291);
xor U9511 (N_9511,N_9111,N_9069);
nand U9512 (N_9512,N_9250,N_9290);
or U9513 (N_9513,N_9289,N_9068);
and U9514 (N_9514,N_9079,N_9214);
xnor U9515 (N_9515,N_9236,N_9106);
and U9516 (N_9516,N_9144,N_9046);
nor U9517 (N_9517,N_9139,N_9256);
or U9518 (N_9518,N_9156,N_9022);
nor U9519 (N_9519,N_9078,N_9071);
and U9520 (N_9520,N_9047,N_9190);
xor U9521 (N_9521,N_9271,N_9101);
xnor U9522 (N_9522,N_9165,N_9288);
nand U9523 (N_9523,N_9200,N_9011);
xnor U9524 (N_9524,N_9127,N_9005);
nand U9525 (N_9525,N_9218,N_9145);
nor U9526 (N_9526,N_9239,N_9177);
nand U9527 (N_9527,N_9283,N_9183);
nand U9528 (N_9528,N_9118,N_9100);
xor U9529 (N_9529,N_9257,N_9142);
nand U9530 (N_9530,N_9000,N_9029);
or U9531 (N_9531,N_9186,N_9084);
or U9532 (N_9532,N_9038,N_9012);
nand U9533 (N_9533,N_9125,N_9116);
nand U9534 (N_9534,N_9292,N_9249);
nand U9535 (N_9535,N_9294,N_9054);
and U9536 (N_9536,N_9181,N_9132);
nand U9537 (N_9537,N_9159,N_9261);
or U9538 (N_9538,N_9066,N_9041);
or U9539 (N_9539,N_9265,N_9006);
or U9540 (N_9540,N_9011,N_9291);
xor U9541 (N_9541,N_9080,N_9089);
nor U9542 (N_9542,N_9100,N_9221);
and U9543 (N_9543,N_9292,N_9273);
nand U9544 (N_9544,N_9240,N_9078);
or U9545 (N_9545,N_9261,N_9207);
nor U9546 (N_9546,N_9026,N_9017);
xnor U9547 (N_9547,N_9134,N_9210);
xnor U9548 (N_9548,N_9277,N_9267);
xnor U9549 (N_9549,N_9001,N_9018);
and U9550 (N_9550,N_9183,N_9021);
nand U9551 (N_9551,N_9253,N_9183);
nor U9552 (N_9552,N_9263,N_9152);
and U9553 (N_9553,N_9128,N_9172);
and U9554 (N_9554,N_9107,N_9192);
or U9555 (N_9555,N_9260,N_9038);
nand U9556 (N_9556,N_9253,N_9100);
nor U9557 (N_9557,N_9293,N_9138);
nor U9558 (N_9558,N_9248,N_9175);
nand U9559 (N_9559,N_9213,N_9296);
and U9560 (N_9560,N_9018,N_9264);
nand U9561 (N_9561,N_9028,N_9230);
xor U9562 (N_9562,N_9232,N_9276);
and U9563 (N_9563,N_9171,N_9087);
nand U9564 (N_9564,N_9207,N_9107);
and U9565 (N_9565,N_9174,N_9228);
nor U9566 (N_9566,N_9276,N_9245);
nand U9567 (N_9567,N_9233,N_9229);
xor U9568 (N_9568,N_9124,N_9025);
or U9569 (N_9569,N_9143,N_9287);
nor U9570 (N_9570,N_9150,N_9026);
or U9571 (N_9571,N_9166,N_9238);
nand U9572 (N_9572,N_9204,N_9218);
xnor U9573 (N_9573,N_9158,N_9014);
nor U9574 (N_9574,N_9262,N_9141);
and U9575 (N_9575,N_9228,N_9291);
nor U9576 (N_9576,N_9206,N_9082);
nor U9577 (N_9577,N_9161,N_9005);
or U9578 (N_9578,N_9158,N_9050);
or U9579 (N_9579,N_9096,N_9105);
xnor U9580 (N_9580,N_9183,N_9055);
or U9581 (N_9581,N_9200,N_9284);
xor U9582 (N_9582,N_9068,N_9111);
or U9583 (N_9583,N_9185,N_9143);
nand U9584 (N_9584,N_9094,N_9023);
nor U9585 (N_9585,N_9080,N_9272);
nor U9586 (N_9586,N_9248,N_9194);
nand U9587 (N_9587,N_9183,N_9109);
and U9588 (N_9588,N_9103,N_9085);
or U9589 (N_9589,N_9208,N_9228);
nor U9590 (N_9590,N_9021,N_9164);
xor U9591 (N_9591,N_9093,N_9108);
nand U9592 (N_9592,N_9051,N_9147);
nor U9593 (N_9593,N_9054,N_9071);
nor U9594 (N_9594,N_9218,N_9260);
and U9595 (N_9595,N_9019,N_9147);
xor U9596 (N_9596,N_9139,N_9236);
nand U9597 (N_9597,N_9208,N_9061);
nor U9598 (N_9598,N_9007,N_9257);
xor U9599 (N_9599,N_9003,N_9162);
xor U9600 (N_9600,N_9355,N_9541);
xor U9601 (N_9601,N_9361,N_9514);
nor U9602 (N_9602,N_9414,N_9515);
nand U9603 (N_9603,N_9468,N_9481);
nor U9604 (N_9604,N_9403,N_9410);
and U9605 (N_9605,N_9376,N_9551);
or U9606 (N_9606,N_9366,N_9463);
nor U9607 (N_9607,N_9378,N_9535);
xor U9608 (N_9608,N_9372,N_9309);
nor U9609 (N_9609,N_9563,N_9335);
or U9610 (N_9610,N_9497,N_9428);
or U9611 (N_9611,N_9461,N_9507);
or U9612 (N_9612,N_9517,N_9446);
or U9613 (N_9613,N_9454,N_9411);
nand U9614 (N_9614,N_9373,N_9333);
xnor U9615 (N_9615,N_9394,N_9437);
xor U9616 (N_9616,N_9576,N_9307);
nor U9617 (N_9617,N_9432,N_9483);
nand U9618 (N_9618,N_9345,N_9529);
or U9619 (N_9619,N_9327,N_9300);
xor U9620 (N_9620,N_9399,N_9451);
and U9621 (N_9621,N_9510,N_9492);
or U9622 (N_9622,N_9533,N_9490);
nor U9623 (N_9623,N_9413,N_9467);
xnor U9624 (N_9624,N_9385,N_9462);
nor U9625 (N_9625,N_9457,N_9342);
nand U9626 (N_9626,N_9475,N_9443);
and U9627 (N_9627,N_9339,N_9306);
or U9628 (N_9628,N_9544,N_9445);
and U9629 (N_9629,N_9397,N_9424);
xor U9630 (N_9630,N_9408,N_9423);
xor U9631 (N_9631,N_9560,N_9386);
or U9632 (N_9632,N_9364,N_9539);
nor U9633 (N_9633,N_9395,N_9485);
and U9634 (N_9634,N_9402,N_9591);
nor U9635 (N_9635,N_9516,N_9405);
xnor U9636 (N_9636,N_9494,N_9564);
nand U9637 (N_9637,N_9469,N_9491);
nor U9638 (N_9638,N_9487,N_9545);
nand U9639 (N_9639,N_9420,N_9547);
nand U9640 (N_9640,N_9417,N_9480);
nand U9641 (N_9641,N_9552,N_9556);
nor U9642 (N_9642,N_9593,N_9512);
and U9643 (N_9643,N_9434,N_9347);
nor U9644 (N_9644,N_9375,N_9573);
or U9645 (N_9645,N_9317,N_9542);
or U9646 (N_9646,N_9572,N_9578);
and U9647 (N_9647,N_9519,N_9441);
nand U9648 (N_9648,N_9599,N_9455);
and U9649 (N_9649,N_9496,N_9555);
xor U9650 (N_9650,N_9370,N_9419);
and U9651 (N_9651,N_9575,N_9574);
xnor U9652 (N_9652,N_9486,N_9587);
or U9653 (N_9653,N_9447,N_9464);
and U9654 (N_9654,N_9525,N_9318);
xnor U9655 (N_9655,N_9416,N_9553);
nor U9656 (N_9656,N_9381,N_9415);
and U9657 (N_9657,N_9508,N_9302);
xor U9658 (N_9658,N_9597,N_9357);
nor U9659 (N_9659,N_9524,N_9334);
and U9660 (N_9660,N_9550,N_9321);
nor U9661 (N_9661,N_9439,N_9543);
or U9662 (N_9662,N_9330,N_9495);
or U9663 (N_9663,N_9577,N_9474);
nor U9664 (N_9664,N_9436,N_9562);
nor U9665 (N_9665,N_9312,N_9374);
xor U9666 (N_9666,N_9350,N_9418);
and U9667 (N_9667,N_9594,N_9592);
nand U9668 (N_9668,N_9584,N_9558);
nand U9669 (N_9669,N_9315,N_9484);
nor U9670 (N_9670,N_9477,N_9581);
nand U9671 (N_9671,N_9588,N_9349);
or U9672 (N_9672,N_9433,N_9459);
xnor U9673 (N_9673,N_9513,N_9323);
xor U9674 (N_9674,N_9389,N_9503);
nor U9675 (N_9675,N_9589,N_9319);
nor U9676 (N_9676,N_9530,N_9353);
xor U9677 (N_9677,N_9412,N_9505);
nand U9678 (N_9678,N_9328,N_9466);
or U9679 (N_9679,N_9470,N_9549);
and U9680 (N_9680,N_9565,N_9362);
nor U9681 (N_9681,N_9383,N_9358);
nor U9682 (N_9682,N_9531,N_9324);
xnor U9683 (N_9683,N_9340,N_9548);
nor U9684 (N_9684,N_9499,N_9569);
nand U9685 (N_9685,N_9393,N_9448);
and U9686 (N_9686,N_9520,N_9528);
or U9687 (N_9687,N_9450,N_9406);
and U9688 (N_9688,N_9427,N_9527);
xor U9689 (N_9689,N_9401,N_9392);
and U9690 (N_9690,N_9396,N_9534);
and U9691 (N_9691,N_9407,N_9346);
and U9692 (N_9692,N_9331,N_9465);
or U9693 (N_9693,N_9438,N_9337);
or U9694 (N_9694,N_9566,N_9532);
xor U9695 (N_9695,N_9301,N_9429);
nor U9696 (N_9696,N_9303,N_9400);
nand U9697 (N_9697,N_9546,N_9580);
nand U9698 (N_9698,N_9479,N_9371);
or U9699 (N_9699,N_9506,N_9311);
or U9700 (N_9700,N_9325,N_9380);
nand U9701 (N_9701,N_9314,N_9360);
nand U9702 (N_9702,N_9310,N_9557);
or U9703 (N_9703,N_9453,N_9568);
nand U9704 (N_9704,N_9368,N_9338);
nor U9705 (N_9705,N_9582,N_9598);
xor U9706 (N_9706,N_9476,N_9567);
xor U9707 (N_9707,N_9460,N_9570);
or U9708 (N_9708,N_9354,N_9518);
xnor U9709 (N_9709,N_9421,N_9536);
or U9710 (N_9710,N_9391,N_9352);
nor U9711 (N_9711,N_9500,N_9387);
nor U9712 (N_9712,N_9472,N_9595);
xnor U9713 (N_9713,N_9489,N_9585);
nand U9714 (N_9714,N_9554,N_9452);
xor U9715 (N_9715,N_9526,N_9379);
or U9716 (N_9716,N_9404,N_9471);
xor U9717 (N_9717,N_9316,N_9422);
xor U9718 (N_9718,N_9341,N_9501);
xor U9719 (N_9719,N_9456,N_9498);
nor U9720 (N_9720,N_9559,N_9351);
nor U9721 (N_9721,N_9377,N_9511);
nor U9722 (N_9722,N_9449,N_9579);
or U9723 (N_9723,N_9442,N_9493);
nand U9724 (N_9724,N_9590,N_9537);
xnor U9725 (N_9725,N_9356,N_9561);
or U9726 (N_9726,N_9329,N_9305);
nand U9727 (N_9727,N_9365,N_9382);
and U9728 (N_9728,N_9430,N_9583);
nand U9729 (N_9729,N_9523,N_9586);
or U9730 (N_9730,N_9478,N_9425);
nand U9731 (N_9731,N_9473,N_9509);
xor U9732 (N_9732,N_9504,N_9409);
nor U9733 (N_9733,N_9435,N_9390);
or U9734 (N_9734,N_9596,N_9482);
nor U9735 (N_9735,N_9348,N_9521);
xor U9736 (N_9736,N_9488,N_9308);
xor U9737 (N_9737,N_9384,N_9343);
or U9738 (N_9738,N_9369,N_9502);
and U9739 (N_9739,N_9344,N_9367);
and U9740 (N_9740,N_9320,N_9440);
xnor U9741 (N_9741,N_9538,N_9336);
or U9742 (N_9742,N_9359,N_9304);
xnor U9743 (N_9743,N_9363,N_9571);
or U9744 (N_9744,N_9322,N_9398);
and U9745 (N_9745,N_9426,N_9431);
or U9746 (N_9746,N_9540,N_9326);
or U9747 (N_9747,N_9313,N_9388);
or U9748 (N_9748,N_9444,N_9332);
and U9749 (N_9749,N_9522,N_9458);
nand U9750 (N_9750,N_9563,N_9584);
nand U9751 (N_9751,N_9548,N_9350);
and U9752 (N_9752,N_9554,N_9539);
and U9753 (N_9753,N_9436,N_9396);
nor U9754 (N_9754,N_9336,N_9480);
nor U9755 (N_9755,N_9517,N_9477);
nor U9756 (N_9756,N_9448,N_9589);
nand U9757 (N_9757,N_9319,N_9577);
xnor U9758 (N_9758,N_9542,N_9561);
and U9759 (N_9759,N_9538,N_9399);
nand U9760 (N_9760,N_9329,N_9493);
nor U9761 (N_9761,N_9514,N_9328);
nand U9762 (N_9762,N_9577,N_9425);
and U9763 (N_9763,N_9549,N_9532);
nand U9764 (N_9764,N_9543,N_9584);
xor U9765 (N_9765,N_9374,N_9542);
and U9766 (N_9766,N_9523,N_9570);
nor U9767 (N_9767,N_9462,N_9322);
nand U9768 (N_9768,N_9529,N_9470);
xnor U9769 (N_9769,N_9340,N_9329);
xor U9770 (N_9770,N_9541,N_9560);
nor U9771 (N_9771,N_9354,N_9511);
xnor U9772 (N_9772,N_9328,N_9425);
and U9773 (N_9773,N_9385,N_9461);
or U9774 (N_9774,N_9503,N_9566);
and U9775 (N_9775,N_9447,N_9549);
xor U9776 (N_9776,N_9380,N_9454);
nand U9777 (N_9777,N_9438,N_9348);
and U9778 (N_9778,N_9315,N_9594);
and U9779 (N_9779,N_9410,N_9319);
xnor U9780 (N_9780,N_9530,N_9387);
and U9781 (N_9781,N_9364,N_9431);
nor U9782 (N_9782,N_9354,N_9410);
or U9783 (N_9783,N_9497,N_9463);
nor U9784 (N_9784,N_9305,N_9514);
nor U9785 (N_9785,N_9397,N_9451);
and U9786 (N_9786,N_9402,N_9572);
and U9787 (N_9787,N_9443,N_9429);
nor U9788 (N_9788,N_9339,N_9327);
and U9789 (N_9789,N_9574,N_9429);
xor U9790 (N_9790,N_9381,N_9521);
or U9791 (N_9791,N_9462,N_9498);
nor U9792 (N_9792,N_9368,N_9552);
and U9793 (N_9793,N_9460,N_9573);
xor U9794 (N_9794,N_9547,N_9333);
nor U9795 (N_9795,N_9539,N_9321);
and U9796 (N_9796,N_9448,N_9545);
xor U9797 (N_9797,N_9556,N_9454);
xor U9798 (N_9798,N_9312,N_9524);
nand U9799 (N_9799,N_9577,N_9558);
or U9800 (N_9800,N_9527,N_9321);
or U9801 (N_9801,N_9502,N_9449);
and U9802 (N_9802,N_9411,N_9503);
nor U9803 (N_9803,N_9552,N_9319);
or U9804 (N_9804,N_9553,N_9361);
and U9805 (N_9805,N_9315,N_9342);
and U9806 (N_9806,N_9508,N_9407);
and U9807 (N_9807,N_9360,N_9522);
nor U9808 (N_9808,N_9436,N_9369);
xor U9809 (N_9809,N_9488,N_9586);
nor U9810 (N_9810,N_9542,N_9496);
nand U9811 (N_9811,N_9469,N_9324);
and U9812 (N_9812,N_9487,N_9594);
xor U9813 (N_9813,N_9438,N_9309);
nor U9814 (N_9814,N_9598,N_9360);
or U9815 (N_9815,N_9311,N_9327);
nor U9816 (N_9816,N_9403,N_9576);
or U9817 (N_9817,N_9480,N_9478);
and U9818 (N_9818,N_9452,N_9403);
or U9819 (N_9819,N_9532,N_9372);
nor U9820 (N_9820,N_9594,N_9528);
or U9821 (N_9821,N_9473,N_9379);
xnor U9822 (N_9822,N_9364,N_9561);
and U9823 (N_9823,N_9471,N_9349);
xnor U9824 (N_9824,N_9423,N_9460);
nand U9825 (N_9825,N_9321,N_9380);
nand U9826 (N_9826,N_9437,N_9490);
nor U9827 (N_9827,N_9344,N_9515);
xor U9828 (N_9828,N_9580,N_9484);
or U9829 (N_9829,N_9370,N_9377);
nor U9830 (N_9830,N_9581,N_9317);
nor U9831 (N_9831,N_9441,N_9384);
and U9832 (N_9832,N_9496,N_9577);
xor U9833 (N_9833,N_9438,N_9378);
and U9834 (N_9834,N_9372,N_9588);
or U9835 (N_9835,N_9596,N_9510);
nand U9836 (N_9836,N_9540,N_9506);
or U9837 (N_9837,N_9533,N_9394);
nand U9838 (N_9838,N_9587,N_9383);
and U9839 (N_9839,N_9381,N_9409);
or U9840 (N_9840,N_9448,N_9597);
xnor U9841 (N_9841,N_9512,N_9474);
or U9842 (N_9842,N_9315,N_9384);
xor U9843 (N_9843,N_9478,N_9374);
and U9844 (N_9844,N_9516,N_9374);
xnor U9845 (N_9845,N_9537,N_9358);
nand U9846 (N_9846,N_9489,N_9513);
and U9847 (N_9847,N_9564,N_9482);
xnor U9848 (N_9848,N_9303,N_9357);
and U9849 (N_9849,N_9514,N_9593);
nor U9850 (N_9850,N_9425,N_9487);
nor U9851 (N_9851,N_9470,N_9322);
nand U9852 (N_9852,N_9425,N_9482);
nor U9853 (N_9853,N_9413,N_9350);
xor U9854 (N_9854,N_9314,N_9495);
nor U9855 (N_9855,N_9405,N_9518);
nand U9856 (N_9856,N_9457,N_9477);
xor U9857 (N_9857,N_9386,N_9471);
and U9858 (N_9858,N_9536,N_9428);
nand U9859 (N_9859,N_9553,N_9467);
nand U9860 (N_9860,N_9402,N_9415);
nand U9861 (N_9861,N_9486,N_9390);
nor U9862 (N_9862,N_9511,N_9462);
and U9863 (N_9863,N_9553,N_9568);
xor U9864 (N_9864,N_9597,N_9349);
and U9865 (N_9865,N_9539,N_9481);
and U9866 (N_9866,N_9325,N_9448);
nor U9867 (N_9867,N_9417,N_9498);
xor U9868 (N_9868,N_9521,N_9520);
nand U9869 (N_9869,N_9364,N_9568);
and U9870 (N_9870,N_9505,N_9536);
nand U9871 (N_9871,N_9414,N_9408);
or U9872 (N_9872,N_9375,N_9526);
nor U9873 (N_9873,N_9485,N_9432);
and U9874 (N_9874,N_9394,N_9368);
and U9875 (N_9875,N_9589,N_9370);
and U9876 (N_9876,N_9390,N_9315);
nand U9877 (N_9877,N_9593,N_9531);
xnor U9878 (N_9878,N_9408,N_9362);
or U9879 (N_9879,N_9532,N_9313);
and U9880 (N_9880,N_9332,N_9578);
nand U9881 (N_9881,N_9459,N_9465);
nor U9882 (N_9882,N_9541,N_9512);
or U9883 (N_9883,N_9531,N_9328);
nand U9884 (N_9884,N_9377,N_9526);
and U9885 (N_9885,N_9345,N_9446);
nand U9886 (N_9886,N_9389,N_9370);
xor U9887 (N_9887,N_9373,N_9357);
nand U9888 (N_9888,N_9446,N_9579);
and U9889 (N_9889,N_9332,N_9448);
nand U9890 (N_9890,N_9430,N_9335);
xnor U9891 (N_9891,N_9426,N_9318);
nor U9892 (N_9892,N_9365,N_9387);
xor U9893 (N_9893,N_9443,N_9352);
nor U9894 (N_9894,N_9437,N_9558);
and U9895 (N_9895,N_9586,N_9344);
xor U9896 (N_9896,N_9455,N_9477);
nor U9897 (N_9897,N_9373,N_9551);
and U9898 (N_9898,N_9338,N_9559);
and U9899 (N_9899,N_9360,N_9409);
nand U9900 (N_9900,N_9663,N_9660);
nand U9901 (N_9901,N_9874,N_9830);
and U9902 (N_9902,N_9645,N_9726);
nor U9903 (N_9903,N_9879,N_9733);
or U9904 (N_9904,N_9678,N_9887);
or U9905 (N_9905,N_9834,N_9842);
nor U9906 (N_9906,N_9739,N_9802);
nor U9907 (N_9907,N_9783,N_9815);
xnor U9908 (N_9908,N_9779,N_9627);
and U9909 (N_9909,N_9870,N_9800);
nor U9910 (N_9910,N_9851,N_9633);
nor U9911 (N_9911,N_9816,N_9799);
or U9912 (N_9912,N_9757,N_9872);
nand U9913 (N_9913,N_9670,N_9692);
nand U9914 (N_9914,N_9616,N_9804);
nor U9915 (N_9915,N_9706,N_9743);
and U9916 (N_9916,N_9658,N_9756);
and U9917 (N_9917,N_9661,N_9632);
or U9918 (N_9918,N_9849,N_9710);
and U9919 (N_9919,N_9676,N_9805);
nor U9920 (N_9920,N_9797,N_9664);
or U9921 (N_9921,N_9636,N_9820);
nand U9922 (N_9922,N_9899,N_9647);
and U9923 (N_9923,N_9693,N_9866);
or U9924 (N_9924,N_9853,N_9701);
nand U9925 (N_9925,N_9723,N_9650);
xor U9926 (N_9926,N_9639,N_9827);
nor U9927 (N_9927,N_9725,N_9886);
and U9928 (N_9928,N_9836,N_9729);
nor U9929 (N_9929,N_9785,N_9705);
or U9930 (N_9930,N_9778,N_9715);
nor U9931 (N_9931,N_9712,N_9727);
and U9932 (N_9932,N_9810,N_9607);
nor U9933 (N_9933,N_9751,N_9737);
nor U9934 (N_9934,N_9606,N_9788);
xnor U9935 (N_9935,N_9792,N_9718);
nor U9936 (N_9936,N_9719,N_9847);
nand U9937 (N_9937,N_9858,N_9690);
nor U9938 (N_9938,N_9686,N_9894);
or U9939 (N_9939,N_9696,N_9646);
xnor U9940 (N_9940,N_9634,N_9776);
or U9941 (N_9941,N_9742,N_9861);
or U9942 (N_9942,N_9709,N_9873);
nor U9943 (N_9943,N_9770,N_9601);
and U9944 (N_9944,N_9652,N_9774);
and U9945 (N_9945,N_9614,N_9669);
nand U9946 (N_9946,N_9608,N_9746);
xnor U9947 (N_9947,N_9612,N_9674);
nor U9948 (N_9948,N_9818,N_9771);
or U9949 (N_9949,N_9855,N_9694);
and U9950 (N_9950,N_9720,N_9624);
xor U9951 (N_9951,N_9837,N_9806);
and U9952 (N_9952,N_9613,N_9611);
nor U9953 (N_9953,N_9898,N_9801);
and U9954 (N_9954,N_9602,N_9666);
nand U9955 (N_9955,N_9654,N_9741);
and U9956 (N_9956,N_9603,N_9825);
or U9957 (N_9957,N_9649,N_9672);
and U9958 (N_9958,N_9782,N_9618);
nand U9959 (N_9959,N_9755,N_9734);
nor U9960 (N_9960,N_9891,N_9713);
or U9961 (N_9961,N_9884,N_9888);
and U9962 (N_9962,N_9772,N_9600);
or U9963 (N_9963,N_9648,N_9609);
and U9964 (N_9964,N_9675,N_9637);
nand U9965 (N_9965,N_9735,N_9644);
nand U9966 (N_9966,N_9716,N_9862);
xor U9967 (N_9967,N_9653,N_9681);
xnor U9968 (N_9968,N_9630,N_9750);
xor U9969 (N_9969,N_9748,N_9688);
nand U9970 (N_9970,N_9813,N_9610);
nor U9971 (N_9971,N_9859,N_9832);
nor U9972 (N_9972,N_9698,N_9795);
and U9973 (N_9973,N_9667,N_9714);
or U9974 (N_9974,N_9895,N_9777);
and U9975 (N_9975,N_9684,N_9761);
or U9976 (N_9976,N_9695,N_9736);
or U9977 (N_9977,N_9848,N_9699);
and U9978 (N_9978,N_9828,N_9821);
or U9979 (N_9979,N_9814,N_9811);
and U9980 (N_9980,N_9864,N_9880);
and U9981 (N_9981,N_9605,N_9626);
and U9982 (N_9982,N_9857,N_9780);
or U9983 (N_9983,N_9683,N_9867);
xnor U9984 (N_9984,N_9728,N_9812);
and U9985 (N_9985,N_9786,N_9789);
nor U9986 (N_9986,N_9856,N_9702);
and U9987 (N_9987,N_9844,N_9680);
nand U9988 (N_9988,N_9892,N_9657);
xnor U9989 (N_9989,N_9707,N_9622);
and U9990 (N_9990,N_9794,N_9835);
nand U9991 (N_9991,N_9691,N_9708);
xnor U9992 (N_9992,N_9869,N_9882);
xnor U9993 (N_9993,N_9717,N_9662);
xor U9994 (N_9994,N_9843,N_9846);
and U9995 (N_9995,N_9865,N_9745);
or U9996 (N_9996,N_9655,N_9787);
xnor U9997 (N_9997,N_9896,N_9885);
nand U9998 (N_9998,N_9700,N_9829);
xnor U9999 (N_9999,N_9833,N_9689);
nor U10000 (N_10000,N_9638,N_9826);
and U10001 (N_10001,N_9781,N_9897);
nor U10002 (N_10002,N_9754,N_9854);
nand U10003 (N_10003,N_9819,N_9831);
or U10004 (N_10004,N_9615,N_9871);
nand U10005 (N_10005,N_9791,N_9752);
or U10006 (N_10006,N_9883,N_9604);
nor U10007 (N_10007,N_9724,N_9641);
xnor U10008 (N_10008,N_9732,N_9822);
or U10009 (N_10009,N_9766,N_9809);
and U10010 (N_10010,N_9763,N_9890);
and U10011 (N_10011,N_9839,N_9807);
xnor U10012 (N_10012,N_9889,N_9640);
xor U10013 (N_10013,N_9659,N_9668);
nor U10014 (N_10014,N_9730,N_9768);
nand U10015 (N_10015,N_9744,N_9628);
or U10016 (N_10016,N_9767,N_9823);
nand U10017 (N_10017,N_9784,N_9685);
and U10018 (N_10018,N_9738,N_9852);
xnor U10019 (N_10019,N_9878,N_9629);
or U10020 (N_10020,N_9620,N_9838);
and U10021 (N_10021,N_9677,N_9642);
nor U10022 (N_10022,N_9711,N_9621);
xnor U10023 (N_10023,N_9840,N_9893);
nor U10024 (N_10024,N_9656,N_9740);
or U10025 (N_10025,N_9773,N_9875);
or U10026 (N_10026,N_9697,N_9673);
or U10027 (N_10027,N_9863,N_9808);
and U10028 (N_10028,N_9703,N_9881);
nand U10029 (N_10029,N_9704,N_9643);
or U10030 (N_10030,N_9860,N_9721);
xnor U10031 (N_10031,N_9671,N_9876);
or U10032 (N_10032,N_9753,N_9764);
or U10033 (N_10033,N_9824,N_9651);
xor U10034 (N_10034,N_9623,N_9762);
xor U10035 (N_10035,N_9760,N_9769);
nor U10036 (N_10036,N_9665,N_9722);
nor U10037 (N_10037,N_9796,N_9631);
or U10038 (N_10038,N_9817,N_9765);
nand U10039 (N_10039,N_9635,N_9759);
nand U10040 (N_10040,N_9850,N_9679);
nand U10041 (N_10041,N_9803,N_9868);
nor U10042 (N_10042,N_9619,N_9775);
nor U10043 (N_10043,N_9877,N_9798);
or U10044 (N_10044,N_9687,N_9793);
nand U10045 (N_10045,N_9790,N_9617);
nor U10046 (N_10046,N_9845,N_9758);
and U10047 (N_10047,N_9682,N_9625);
or U10048 (N_10048,N_9747,N_9749);
xor U10049 (N_10049,N_9841,N_9731);
nand U10050 (N_10050,N_9867,N_9827);
nor U10051 (N_10051,N_9694,N_9693);
or U10052 (N_10052,N_9863,N_9737);
xor U10053 (N_10053,N_9636,N_9734);
nand U10054 (N_10054,N_9880,N_9669);
xnor U10055 (N_10055,N_9656,N_9843);
nand U10056 (N_10056,N_9630,N_9840);
xor U10057 (N_10057,N_9677,N_9638);
nor U10058 (N_10058,N_9749,N_9842);
nand U10059 (N_10059,N_9618,N_9829);
or U10060 (N_10060,N_9852,N_9791);
xor U10061 (N_10061,N_9896,N_9604);
or U10062 (N_10062,N_9727,N_9675);
xor U10063 (N_10063,N_9871,N_9609);
xor U10064 (N_10064,N_9719,N_9834);
xor U10065 (N_10065,N_9828,N_9646);
xor U10066 (N_10066,N_9712,N_9800);
xnor U10067 (N_10067,N_9711,N_9625);
or U10068 (N_10068,N_9770,N_9769);
and U10069 (N_10069,N_9884,N_9645);
or U10070 (N_10070,N_9649,N_9805);
and U10071 (N_10071,N_9818,N_9750);
nor U10072 (N_10072,N_9627,N_9636);
and U10073 (N_10073,N_9605,N_9673);
or U10074 (N_10074,N_9878,N_9742);
or U10075 (N_10075,N_9683,N_9780);
nor U10076 (N_10076,N_9773,N_9627);
and U10077 (N_10077,N_9854,N_9716);
or U10078 (N_10078,N_9797,N_9885);
nor U10079 (N_10079,N_9834,N_9730);
xnor U10080 (N_10080,N_9819,N_9797);
or U10081 (N_10081,N_9797,N_9841);
nor U10082 (N_10082,N_9729,N_9603);
nand U10083 (N_10083,N_9689,N_9662);
nor U10084 (N_10084,N_9796,N_9758);
xnor U10085 (N_10085,N_9763,N_9758);
nor U10086 (N_10086,N_9771,N_9700);
nand U10087 (N_10087,N_9859,N_9714);
xor U10088 (N_10088,N_9616,N_9720);
and U10089 (N_10089,N_9705,N_9653);
nor U10090 (N_10090,N_9838,N_9728);
and U10091 (N_10091,N_9890,N_9847);
or U10092 (N_10092,N_9789,N_9628);
nand U10093 (N_10093,N_9703,N_9673);
nand U10094 (N_10094,N_9741,N_9727);
and U10095 (N_10095,N_9829,N_9729);
nand U10096 (N_10096,N_9629,N_9649);
nand U10097 (N_10097,N_9870,N_9731);
or U10098 (N_10098,N_9879,N_9878);
nand U10099 (N_10099,N_9715,N_9769);
nor U10100 (N_10100,N_9637,N_9756);
xor U10101 (N_10101,N_9665,N_9636);
nand U10102 (N_10102,N_9862,N_9643);
or U10103 (N_10103,N_9612,N_9719);
xnor U10104 (N_10104,N_9737,N_9781);
and U10105 (N_10105,N_9871,N_9755);
nand U10106 (N_10106,N_9678,N_9866);
nand U10107 (N_10107,N_9634,N_9853);
nand U10108 (N_10108,N_9787,N_9890);
nand U10109 (N_10109,N_9758,N_9682);
nor U10110 (N_10110,N_9807,N_9600);
nor U10111 (N_10111,N_9775,N_9891);
xor U10112 (N_10112,N_9713,N_9614);
or U10113 (N_10113,N_9607,N_9637);
or U10114 (N_10114,N_9722,N_9888);
nor U10115 (N_10115,N_9669,N_9760);
or U10116 (N_10116,N_9658,N_9654);
xor U10117 (N_10117,N_9763,N_9785);
nand U10118 (N_10118,N_9641,N_9771);
and U10119 (N_10119,N_9633,N_9876);
xor U10120 (N_10120,N_9666,N_9672);
xor U10121 (N_10121,N_9709,N_9630);
nor U10122 (N_10122,N_9681,N_9890);
xnor U10123 (N_10123,N_9885,N_9637);
or U10124 (N_10124,N_9651,N_9734);
nand U10125 (N_10125,N_9712,N_9757);
xor U10126 (N_10126,N_9753,N_9656);
or U10127 (N_10127,N_9830,N_9689);
and U10128 (N_10128,N_9664,N_9798);
and U10129 (N_10129,N_9767,N_9699);
xnor U10130 (N_10130,N_9661,N_9744);
nand U10131 (N_10131,N_9720,N_9651);
and U10132 (N_10132,N_9778,N_9856);
or U10133 (N_10133,N_9630,N_9605);
nand U10134 (N_10134,N_9634,N_9676);
or U10135 (N_10135,N_9685,N_9763);
xnor U10136 (N_10136,N_9807,N_9730);
xor U10137 (N_10137,N_9875,N_9774);
or U10138 (N_10138,N_9867,N_9618);
xnor U10139 (N_10139,N_9747,N_9683);
or U10140 (N_10140,N_9603,N_9676);
and U10141 (N_10141,N_9877,N_9778);
or U10142 (N_10142,N_9784,N_9655);
and U10143 (N_10143,N_9865,N_9733);
and U10144 (N_10144,N_9763,N_9801);
nor U10145 (N_10145,N_9776,N_9829);
xnor U10146 (N_10146,N_9733,N_9669);
nor U10147 (N_10147,N_9802,N_9749);
nand U10148 (N_10148,N_9849,N_9826);
xnor U10149 (N_10149,N_9757,N_9882);
and U10150 (N_10150,N_9717,N_9893);
nor U10151 (N_10151,N_9888,N_9685);
nand U10152 (N_10152,N_9810,N_9895);
and U10153 (N_10153,N_9840,N_9883);
nand U10154 (N_10154,N_9760,N_9743);
nand U10155 (N_10155,N_9886,N_9728);
and U10156 (N_10156,N_9705,N_9751);
and U10157 (N_10157,N_9715,N_9741);
or U10158 (N_10158,N_9628,N_9687);
nor U10159 (N_10159,N_9705,N_9713);
or U10160 (N_10160,N_9882,N_9791);
xnor U10161 (N_10161,N_9851,N_9655);
nand U10162 (N_10162,N_9600,N_9839);
or U10163 (N_10163,N_9690,N_9715);
nor U10164 (N_10164,N_9646,N_9844);
nor U10165 (N_10165,N_9651,N_9860);
xnor U10166 (N_10166,N_9762,N_9700);
nor U10167 (N_10167,N_9741,N_9810);
nand U10168 (N_10168,N_9853,N_9678);
xor U10169 (N_10169,N_9693,N_9876);
nor U10170 (N_10170,N_9775,N_9641);
xnor U10171 (N_10171,N_9743,N_9625);
and U10172 (N_10172,N_9857,N_9739);
nand U10173 (N_10173,N_9760,N_9697);
xor U10174 (N_10174,N_9659,N_9831);
and U10175 (N_10175,N_9786,N_9625);
or U10176 (N_10176,N_9736,N_9851);
nor U10177 (N_10177,N_9690,N_9779);
xnor U10178 (N_10178,N_9850,N_9788);
xor U10179 (N_10179,N_9805,N_9641);
and U10180 (N_10180,N_9707,N_9667);
nand U10181 (N_10181,N_9656,N_9771);
xnor U10182 (N_10182,N_9673,N_9617);
or U10183 (N_10183,N_9759,N_9838);
nand U10184 (N_10184,N_9827,N_9845);
or U10185 (N_10185,N_9833,N_9655);
xor U10186 (N_10186,N_9714,N_9637);
nand U10187 (N_10187,N_9735,N_9780);
xnor U10188 (N_10188,N_9889,N_9783);
nor U10189 (N_10189,N_9809,N_9820);
nor U10190 (N_10190,N_9667,N_9622);
xnor U10191 (N_10191,N_9667,N_9820);
or U10192 (N_10192,N_9805,N_9798);
nor U10193 (N_10193,N_9622,N_9721);
nor U10194 (N_10194,N_9841,N_9823);
nor U10195 (N_10195,N_9780,N_9662);
nor U10196 (N_10196,N_9714,N_9688);
nor U10197 (N_10197,N_9837,N_9703);
nand U10198 (N_10198,N_9730,N_9689);
and U10199 (N_10199,N_9693,N_9712);
nor U10200 (N_10200,N_10194,N_9909);
and U10201 (N_10201,N_10124,N_10099);
or U10202 (N_10202,N_10106,N_9996);
nor U10203 (N_10203,N_9929,N_10006);
nand U10204 (N_10204,N_9924,N_10191);
nor U10205 (N_10205,N_10011,N_10035);
and U10206 (N_10206,N_10033,N_9920);
nor U10207 (N_10207,N_10160,N_9987);
nand U10208 (N_10208,N_10027,N_10064);
and U10209 (N_10209,N_10116,N_10005);
nand U10210 (N_10210,N_9946,N_10195);
and U10211 (N_10211,N_10135,N_10184);
or U10212 (N_10212,N_10047,N_10082);
nand U10213 (N_10213,N_10058,N_9950);
or U10214 (N_10214,N_10198,N_10010);
nor U10215 (N_10215,N_10022,N_9932);
or U10216 (N_10216,N_9927,N_10147);
xor U10217 (N_10217,N_9925,N_10144);
or U10218 (N_10218,N_10186,N_9978);
nor U10219 (N_10219,N_10055,N_10090);
or U10220 (N_10220,N_9935,N_10165);
or U10221 (N_10221,N_9958,N_10009);
nor U10222 (N_10222,N_9913,N_10016);
nor U10223 (N_10223,N_10134,N_10030);
nand U10224 (N_10224,N_10119,N_9911);
xnor U10225 (N_10225,N_10012,N_10152);
and U10226 (N_10226,N_9965,N_9954);
xor U10227 (N_10227,N_10038,N_10000);
xnor U10228 (N_10228,N_10168,N_9990);
or U10229 (N_10229,N_10042,N_9976);
nor U10230 (N_10230,N_10196,N_10175);
nor U10231 (N_10231,N_9922,N_10133);
nand U10232 (N_10232,N_9986,N_9930);
xnor U10233 (N_10233,N_10032,N_10017);
nand U10234 (N_10234,N_10050,N_9940);
or U10235 (N_10235,N_10182,N_10178);
nor U10236 (N_10236,N_10069,N_10138);
nor U10237 (N_10237,N_9979,N_9989);
nand U10238 (N_10238,N_10077,N_10020);
or U10239 (N_10239,N_9974,N_10072);
or U10240 (N_10240,N_10130,N_10065);
nand U10241 (N_10241,N_10159,N_10048);
or U10242 (N_10242,N_10054,N_10170);
nand U10243 (N_10243,N_10008,N_10105);
or U10244 (N_10244,N_9998,N_10003);
and U10245 (N_10245,N_10150,N_10084);
nor U10246 (N_10246,N_9952,N_10117);
xor U10247 (N_10247,N_9902,N_10101);
nor U10248 (N_10248,N_9942,N_9919);
nand U10249 (N_10249,N_9916,N_10102);
nand U10250 (N_10250,N_10085,N_9988);
and U10251 (N_10251,N_10114,N_10148);
nand U10252 (N_10252,N_9982,N_10031);
nand U10253 (N_10253,N_10163,N_9917);
and U10254 (N_10254,N_10097,N_9951);
nand U10255 (N_10255,N_10068,N_10121);
nor U10256 (N_10256,N_10014,N_10154);
nor U10257 (N_10257,N_10029,N_10060);
or U10258 (N_10258,N_10043,N_9923);
or U10259 (N_10259,N_10081,N_10018);
nand U10260 (N_10260,N_9966,N_10136);
xnor U10261 (N_10261,N_10171,N_10040);
nand U10262 (N_10262,N_10123,N_9901);
nor U10263 (N_10263,N_10128,N_9928);
and U10264 (N_10264,N_10180,N_9997);
nand U10265 (N_10265,N_9949,N_9957);
xnor U10266 (N_10266,N_10070,N_10083);
or U10267 (N_10267,N_9903,N_10164);
nand U10268 (N_10268,N_10001,N_10073);
nor U10269 (N_10269,N_10051,N_9938);
and U10270 (N_10270,N_10122,N_10061);
xor U10271 (N_10271,N_9984,N_10067);
nor U10272 (N_10272,N_10026,N_9918);
xor U10273 (N_10273,N_9972,N_9977);
and U10274 (N_10274,N_10125,N_10110);
nor U10275 (N_10275,N_10062,N_9944);
nand U10276 (N_10276,N_10157,N_10041);
and U10277 (N_10277,N_9926,N_10126);
nand U10278 (N_10278,N_10132,N_10181);
and U10279 (N_10279,N_10078,N_10088);
xnor U10280 (N_10280,N_10100,N_10053);
nor U10281 (N_10281,N_10057,N_10046);
or U10282 (N_10282,N_10197,N_10049);
and U10283 (N_10283,N_10177,N_9955);
or U10284 (N_10284,N_10158,N_10140);
nor U10285 (N_10285,N_10146,N_9995);
nor U10286 (N_10286,N_10019,N_9905);
xnor U10287 (N_10287,N_10066,N_10129);
nor U10288 (N_10288,N_10141,N_9971);
nand U10289 (N_10289,N_10095,N_10059);
or U10290 (N_10290,N_10025,N_10193);
and U10291 (N_10291,N_10076,N_10192);
and U10292 (N_10292,N_9945,N_10172);
and U10293 (N_10293,N_9904,N_10161);
and U10294 (N_10294,N_9985,N_9933);
xnor U10295 (N_10295,N_10063,N_10096);
xor U10296 (N_10296,N_9948,N_9908);
and U10297 (N_10297,N_9943,N_10098);
xor U10298 (N_10298,N_10111,N_10094);
or U10299 (N_10299,N_9969,N_10151);
nand U10300 (N_10300,N_10075,N_10120);
xor U10301 (N_10301,N_9931,N_10023);
and U10302 (N_10302,N_10034,N_10103);
nand U10303 (N_10303,N_9980,N_9999);
or U10304 (N_10304,N_10037,N_10166);
nor U10305 (N_10305,N_9970,N_9921);
nand U10306 (N_10306,N_10039,N_10139);
and U10307 (N_10307,N_10185,N_10007);
nor U10308 (N_10308,N_10115,N_10086);
nand U10309 (N_10309,N_10156,N_10137);
nor U10310 (N_10310,N_10089,N_10169);
xnor U10311 (N_10311,N_10188,N_10021);
nor U10312 (N_10312,N_9936,N_10071);
nor U10313 (N_10313,N_10183,N_10002);
xor U10314 (N_10314,N_10056,N_10199);
xnor U10315 (N_10315,N_10131,N_9910);
nor U10316 (N_10316,N_10104,N_10045);
nor U10317 (N_10317,N_10080,N_10093);
nor U10318 (N_10318,N_9937,N_9953);
nor U10319 (N_10319,N_9934,N_10173);
xnor U10320 (N_10320,N_9956,N_9961);
xnor U10321 (N_10321,N_10176,N_10036);
xnor U10322 (N_10322,N_10079,N_10155);
xnor U10323 (N_10323,N_10087,N_9939);
xnor U10324 (N_10324,N_9914,N_10149);
nand U10325 (N_10325,N_9900,N_10174);
xnor U10326 (N_10326,N_9993,N_10013);
nor U10327 (N_10327,N_9975,N_10113);
or U10328 (N_10328,N_9941,N_9915);
nor U10329 (N_10329,N_9983,N_10109);
or U10330 (N_10330,N_10112,N_9991);
and U10331 (N_10331,N_9963,N_10167);
or U10332 (N_10332,N_10004,N_10153);
nand U10333 (N_10333,N_10143,N_10015);
or U10334 (N_10334,N_10052,N_9973);
or U10335 (N_10335,N_10107,N_9912);
and U10336 (N_10336,N_10190,N_10145);
and U10337 (N_10337,N_9981,N_9907);
xor U10338 (N_10338,N_9962,N_10127);
nand U10339 (N_10339,N_9947,N_10028);
nor U10340 (N_10340,N_9994,N_10189);
nand U10341 (N_10341,N_9960,N_10092);
or U10342 (N_10342,N_10074,N_10024);
xor U10343 (N_10343,N_9964,N_10187);
nor U10344 (N_10344,N_9968,N_10142);
and U10345 (N_10345,N_9967,N_10118);
nor U10346 (N_10346,N_10179,N_9959);
and U10347 (N_10347,N_9906,N_9992);
nand U10348 (N_10348,N_10108,N_10162);
and U10349 (N_10349,N_10044,N_10091);
xor U10350 (N_10350,N_9914,N_10132);
or U10351 (N_10351,N_9927,N_10120);
nand U10352 (N_10352,N_9921,N_10178);
or U10353 (N_10353,N_10131,N_9939);
and U10354 (N_10354,N_9900,N_10097);
or U10355 (N_10355,N_10135,N_10132);
xor U10356 (N_10356,N_10064,N_10118);
xor U10357 (N_10357,N_9950,N_10112);
or U10358 (N_10358,N_9934,N_10190);
and U10359 (N_10359,N_10083,N_10183);
and U10360 (N_10360,N_10029,N_10125);
nand U10361 (N_10361,N_9987,N_10070);
nand U10362 (N_10362,N_9930,N_9976);
nand U10363 (N_10363,N_10197,N_9964);
nand U10364 (N_10364,N_9948,N_9982);
and U10365 (N_10365,N_10162,N_10103);
nor U10366 (N_10366,N_10184,N_9999);
nor U10367 (N_10367,N_10129,N_10117);
nor U10368 (N_10368,N_9921,N_9912);
and U10369 (N_10369,N_9933,N_10051);
and U10370 (N_10370,N_9966,N_10116);
or U10371 (N_10371,N_10026,N_10187);
nand U10372 (N_10372,N_10004,N_10184);
and U10373 (N_10373,N_10092,N_10036);
or U10374 (N_10374,N_10175,N_9969);
nor U10375 (N_10375,N_9981,N_10032);
and U10376 (N_10376,N_10158,N_9963);
nand U10377 (N_10377,N_10024,N_10084);
xnor U10378 (N_10378,N_10048,N_9959);
or U10379 (N_10379,N_9948,N_10014);
nor U10380 (N_10380,N_10096,N_10164);
xnor U10381 (N_10381,N_10086,N_9920);
xnor U10382 (N_10382,N_9933,N_10096);
nor U10383 (N_10383,N_10194,N_10148);
nor U10384 (N_10384,N_9950,N_10068);
xnor U10385 (N_10385,N_10020,N_9956);
xnor U10386 (N_10386,N_10193,N_10143);
xor U10387 (N_10387,N_9913,N_9994);
xnor U10388 (N_10388,N_9986,N_10167);
nor U10389 (N_10389,N_10179,N_10058);
nand U10390 (N_10390,N_10050,N_10163);
xnor U10391 (N_10391,N_9945,N_9947);
nor U10392 (N_10392,N_10006,N_9954);
nand U10393 (N_10393,N_10039,N_9901);
nand U10394 (N_10394,N_9996,N_10089);
or U10395 (N_10395,N_10128,N_9942);
or U10396 (N_10396,N_10187,N_9930);
and U10397 (N_10397,N_9900,N_10165);
and U10398 (N_10398,N_10014,N_9952);
nand U10399 (N_10399,N_9944,N_10089);
nor U10400 (N_10400,N_10117,N_10155);
and U10401 (N_10401,N_10152,N_10149);
nor U10402 (N_10402,N_9922,N_9976);
and U10403 (N_10403,N_10147,N_10055);
and U10404 (N_10404,N_10167,N_10051);
and U10405 (N_10405,N_9967,N_9935);
and U10406 (N_10406,N_9973,N_10056);
nor U10407 (N_10407,N_9993,N_10006);
nor U10408 (N_10408,N_10163,N_10159);
nand U10409 (N_10409,N_9938,N_10072);
and U10410 (N_10410,N_10141,N_10190);
xor U10411 (N_10411,N_10053,N_10144);
nor U10412 (N_10412,N_9914,N_10137);
xor U10413 (N_10413,N_10055,N_10084);
nor U10414 (N_10414,N_9980,N_9916);
or U10415 (N_10415,N_10111,N_9929);
nand U10416 (N_10416,N_10099,N_10193);
or U10417 (N_10417,N_10132,N_10105);
or U10418 (N_10418,N_10047,N_10155);
nand U10419 (N_10419,N_9988,N_10184);
and U10420 (N_10420,N_10045,N_10195);
or U10421 (N_10421,N_9957,N_9915);
nor U10422 (N_10422,N_9986,N_10097);
and U10423 (N_10423,N_9910,N_10045);
or U10424 (N_10424,N_10072,N_10160);
nor U10425 (N_10425,N_9986,N_10115);
xnor U10426 (N_10426,N_10007,N_10086);
nand U10427 (N_10427,N_9998,N_10114);
nor U10428 (N_10428,N_9902,N_10123);
nand U10429 (N_10429,N_9958,N_9914);
and U10430 (N_10430,N_9949,N_10186);
and U10431 (N_10431,N_10084,N_9925);
nand U10432 (N_10432,N_10178,N_9935);
or U10433 (N_10433,N_10122,N_10006);
xnor U10434 (N_10434,N_9927,N_10048);
nand U10435 (N_10435,N_10180,N_10061);
nor U10436 (N_10436,N_9961,N_10031);
xnor U10437 (N_10437,N_9966,N_9961);
nor U10438 (N_10438,N_9926,N_10194);
xnor U10439 (N_10439,N_10069,N_9912);
and U10440 (N_10440,N_9907,N_9952);
nor U10441 (N_10441,N_9953,N_9996);
or U10442 (N_10442,N_10159,N_10108);
or U10443 (N_10443,N_10043,N_10129);
nor U10444 (N_10444,N_9924,N_9925);
nand U10445 (N_10445,N_10173,N_9928);
or U10446 (N_10446,N_10131,N_10137);
and U10447 (N_10447,N_10020,N_10087);
nor U10448 (N_10448,N_10042,N_10032);
and U10449 (N_10449,N_9946,N_9986);
nand U10450 (N_10450,N_10183,N_10119);
nor U10451 (N_10451,N_10032,N_9913);
and U10452 (N_10452,N_10090,N_10109);
nor U10453 (N_10453,N_10061,N_9953);
nand U10454 (N_10454,N_10183,N_9923);
or U10455 (N_10455,N_10098,N_10089);
nor U10456 (N_10456,N_10125,N_10121);
or U10457 (N_10457,N_10130,N_10138);
and U10458 (N_10458,N_9969,N_10147);
or U10459 (N_10459,N_10021,N_10134);
nor U10460 (N_10460,N_10104,N_10135);
nand U10461 (N_10461,N_9939,N_10015);
nor U10462 (N_10462,N_9929,N_10146);
and U10463 (N_10463,N_9900,N_9928);
nand U10464 (N_10464,N_10180,N_9980);
or U10465 (N_10465,N_10124,N_9933);
nor U10466 (N_10466,N_10062,N_10122);
or U10467 (N_10467,N_9940,N_10047);
and U10468 (N_10468,N_10154,N_10167);
and U10469 (N_10469,N_9987,N_10021);
or U10470 (N_10470,N_10007,N_10031);
or U10471 (N_10471,N_10193,N_9971);
or U10472 (N_10472,N_10184,N_10145);
xor U10473 (N_10473,N_10077,N_10074);
or U10474 (N_10474,N_10136,N_9930);
or U10475 (N_10475,N_10138,N_9937);
nor U10476 (N_10476,N_10095,N_10104);
nor U10477 (N_10477,N_9930,N_10163);
xor U10478 (N_10478,N_9904,N_9956);
or U10479 (N_10479,N_10190,N_10131);
or U10480 (N_10480,N_10102,N_10087);
nand U10481 (N_10481,N_9930,N_10074);
nor U10482 (N_10482,N_10179,N_9925);
or U10483 (N_10483,N_10136,N_9991);
or U10484 (N_10484,N_10076,N_10068);
nand U10485 (N_10485,N_10106,N_9981);
or U10486 (N_10486,N_10058,N_10105);
and U10487 (N_10487,N_10196,N_10111);
or U10488 (N_10488,N_9995,N_9933);
and U10489 (N_10489,N_10136,N_9997);
nor U10490 (N_10490,N_9953,N_10034);
xor U10491 (N_10491,N_10064,N_9974);
nor U10492 (N_10492,N_10198,N_10071);
and U10493 (N_10493,N_10108,N_10154);
or U10494 (N_10494,N_10158,N_10054);
xor U10495 (N_10495,N_10095,N_10146);
nand U10496 (N_10496,N_10149,N_10143);
nand U10497 (N_10497,N_10007,N_10152);
or U10498 (N_10498,N_10110,N_10009);
nor U10499 (N_10499,N_9976,N_10155);
xor U10500 (N_10500,N_10292,N_10235);
nand U10501 (N_10501,N_10379,N_10374);
nand U10502 (N_10502,N_10433,N_10453);
xnor U10503 (N_10503,N_10418,N_10388);
or U10504 (N_10504,N_10454,N_10449);
nor U10505 (N_10505,N_10497,N_10356);
xor U10506 (N_10506,N_10441,N_10206);
nand U10507 (N_10507,N_10463,N_10320);
nor U10508 (N_10508,N_10218,N_10373);
xor U10509 (N_10509,N_10483,N_10289);
or U10510 (N_10510,N_10307,N_10305);
nand U10511 (N_10511,N_10347,N_10465);
xnor U10512 (N_10512,N_10428,N_10225);
nor U10513 (N_10513,N_10425,N_10415);
or U10514 (N_10514,N_10499,N_10229);
nand U10515 (N_10515,N_10417,N_10223);
nand U10516 (N_10516,N_10341,N_10215);
or U10517 (N_10517,N_10475,N_10286);
or U10518 (N_10518,N_10321,N_10464);
nor U10519 (N_10519,N_10406,N_10244);
nor U10520 (N_10520,N_10240,N_10348);
xnor U10521 (N_10521,N_10239,N_10477);
xor U10522 (N_10522,N_10359,N_10284);
nand U10523 (N_10523,N_10450,N_10285);
and U10524 (N_10524,N_10455,N_10330);
nand U10525 (N_10525,N_10457,N_10252);
and U10526 (N_10526,N_10443,N_10383);
and U10527 (N_10527,N_10226,N_10291);
or U10528 (N_10528,N_10234,N_10430);
or U10529 (N_10529,N_10259,N_10227);
nor U10530 (N_10530,N_10371,N_10325);
and U10531 (N_10531,N_10385,N_10300);
xor U10532 (N_10532,N_10365,N_10380);
xor U10533 (N_10533,N_10436,N_10427);
or U10534 (N_10534,N_10253,N_10386);
nor U10535 (N_10535,N_10312,N_10261);
nor U10536 (N_10536,N_10423,N_10370);
nor U10537 (N_10537,N_10217,N_10280);
or U10538 (N_10538,N_10279,N_10466);
nand U10539 (N_10539,N_10474,N_10272);
nor U10540 (N_10540,N_10209,N_10316);
or U10541 (N_10541,N_10358,N_10344);
nand U10542 (N_10542,N_10250,N_10322);
xor U10543 (N_10543,N_10339,N_10294);
nor U10544 (N_10544,N_10257,N_10412);
xnor U10545 (N_10545,N_10486,N_10340);
xnor U10546 (N_10546,N_10381,N_10256);
xnor U10547 (N_10547,N_10470,N_10432);
and U10548 (N_10548,N_10458,N_10233);
and U10549 (N_10549,N_10313,N_10243);
or U10550 (N_10550,N_10440,N_10387);
or U10551 (N_10551,N_10476,N_10298);
xor U10552 (N_10552,N_10277,N_10364);
nand U10553 (N_10553,N_10437,N_10489);
nor U10554 (N_10554,N_10404,N_10461);
nand U10555 (N_10555,N_10293,N_10210);
nor U10556 (N_10556,N_10248,N_10480);
and U10557 (N_10557,N_10398,N_10420);
or U10558 (N_10558,N_10262,N_10214);
or U10559 (N_10559,N_10354,N_10408);
nand U10560 (N_10560,N_10376,N_10459);
nor U10561 (N_10561,N_10485,N_10202);
or U10562 (N_10562,N_10336,N_10296);
nor U10563 (N_10563,N_10382,N_10488);
and U10564 (N_10564,N_10472,N_10447);
or U10565 (N_10565,N_10448,N_10343);
and U10566 (N_10566,N_10492,N_10342);
or U10567 (N_10567,N_10274,N_10351);
nor U10568 (N_10568,N_10283,N_10334);
or U10569 (N_10569,N_10290,N_10324);
nor U10570 (N_10570,N_10350,N_10281);
nand U10571 (N_10571,N_10378,N_10241);
and U10572 (N_10572,N_10255,N_10473);
and U10573 (N_10573,N_10328,N_10216);
xnor U10574 (N_10574,N_10419,N_10395);
nand U10575 (N_10575,N_10487,N_10391);
nand U10576 (N_10576,N_10287,N_10212);
nor U10577 (N_10577,N_10399,N_10394);
nand U10578 (N_10578,N_10352,N_10219);
and U10579 (N_10579,N_10236,N_10393);
nand U10580 (N_10580,N_10315,N_10462);
xnor U10581 (N_10581,N_10242,N_10246);
xnor U10582 (N_10582,N_10203,N_10451);
xor U10583 (N_10583,N_10375,N_10349);
xnor U10584 (N_10584,N_10208,N_10366);
nor U10585 (N_10585,N_10377,N_10200);
xor U10586 (N_10586,N_10355,N_10369);
xnor U10587 (N_10587,N_10269,N_10491);
and U10588 (N_10588,N_10360,N_10251);
nand U10589 (N_10589,N_10338,N_10314);
nand U10590 (N_10590,N_10361,N_10362);
or U10591 (N_10591,N_10495,N_10201);
xnor U10592 (N_10592,N_10372,N_10258);
and U10593 (N_10593,N_10438,N_10207);
nand U10594 (N_10594,N_10389,N_10402);
xor U10595 (N_10595,N_10498,N_10230);
nand U10596 (N_10596,N_10442,N_10345);
nand U10597 (N_10597,N_10303,N_10435);
nand U10598 (N_10598,N_10329,N_10392);
nand U10599 (N_10599,N_10318,N_10431);
nand U10600 (N_10600,N_10490,N_10205);
nor U10601 (N_10601,N_10446,N_10301);
nor U10602 (N_10602,N_10434,N_10297);
or U10603 (N_10603,N_10471,N_10396);
and U10604 (N_10604,N_10335,N_10327);
xor U10605 (N_10605,N_10414,N_10228);
and U10606 (N_10606,N_10231,N_10260);
nand U10607 (N_10607,N_10309,N_10468);
xnor U10608 (N_10608,N_10479,N_10278);
nand U10609 (N_10609,N_10310,N_10222);
xnor U10610 (N_10610,N_10238,N_10416);
or U10611 (N_10611,N_10493,N_10496);
xnor U10612 (N_10612,N_10275,N_10400);
or U10613 (N_10613,N_10265,N_10456);
nand U10614 (N_10614,N_10319,N_10221);
nor U10615 (N_10615,N_10333,N_10271);
nor U10616 (N_10616,N_10481,N_10288);
nor U10617 (N_10617,N_10247,N_10295);
nand U10618 (N_10618,N_10452,N_10264);
or U10619 (N_10619,N_10323,N_10422);
or U10620 (N_10620,N_10204,N_10401);
xnor U10621 (N_10621,N_10224,N_10413);
xnor U10622 (N_10622,N_10211,N_10306);
and U10623 (N_10623,N_10424,N_10411);
nand U10624 (N_10624,N_10444,N_10397);
xor U10625 (N_10625,N_10403,N_10213);
nor U10626 (N_10626,N_10429,N_10421);
or U10627 (N_10627,N_10439,N_10282);
xnor U10628 (N_10628,N_10263,N_10407);
or U10629 (N_10629,N_10245,N_10332);
and U10630 (N_10630,N_10494,N_10390);
nor U10631 (N_10631,N_10410,N_10308);
or U10632 (N_10632,N_10326,N_10270);
xor U10633 (N_10633,N_10445,N_10482);
nand U10634 (N_10634,N_10384,N_10237);
nand U10635 (N_10635,N_10311,N_10353);
and U10636 (N_10636,N_10331,N_10405);
and U10637 (N_10637,N_10478,N_10232);
nand U10638 (N_10638,N_10302,N_10460);
and U10639 (N_10639,N_10273,N_10368);
and U10640 (N_10640,N_10299,N_10249);
and U10641 (N_10641,N_10317,N_10469);
nand U10642 (N_10642,N_10363,N_10337);
nor U10643 (N_10643,N_10484,N_10267);
xor U10644 (N_10644,N_10268,N_10254);
or U10645 (N_10645,N_10467,N_10426);
nor U10646 (N_10646,N_10266,N_10357);
and U10647 (N_10647,N_10220,N_10276);
nor U10648 (N_10648,N_10367,N_10304);
or U10649 (N_10649,N_10409,N_10346);
nor U10650 (N_10650,N_10255,N_10457);
and U10651 (N_10651,N_10357,N_10473);
or U10652 (N_10652,N_10489,N_10252);
xor U10653 (N_10653,N_10390,N_10263);
or U10654 (N_10654,N_10357,N_10237);
nand U10655 (N_10655,N_10379,N_10399);
xor U10656 (N_10656,N_10365,N_10350);
nor U10657 (N_10657,N_10225,N_10408);
and U10658 (N_10658,N_10429,N_10402);
xor U10659 (N_10659,N_10429,N_10276);
nor U10660 (N_10660,N_10247,N_10481);
xor U10661 (N_10661,N_10272,N_10395);
and U10662 (N_10662,N_10370,N_10293);
and U10663 (N_10663,N_10274,N_10495);
xnor U10664 (N_10664,N_10317,N_10462);
xor U10665 (N_10665,N_10494,N_10413);
and U10666 (N_10666,N_10326,N_10210);
xor U10667 (N_10667,N_10416,N_10399);
and U10668 (N_10668,N_10269,N_10339);
nor U10669 (N_10669,N_10473,N_10327);
nor U10670 (N_10670,N_10493,N_10453);
and U10671 (N_10671,N_10242,N_10252);
or U10672 (N_10672,N_10473,N_10386);
nor U10673 (N_10673,N_10220,N_10341);
nand U10674 (N_10674,N_10480,N_10445);
nand U10675 (N_10675,N_10391,N_10266);
or U10676 (N_10676,N_10415,N_10384);
nand U10677 (N_10677,N_10361,N_10243);
nand U10678 (N_10678,N_10268,N_10333);
nand U10679 (N_10679,N_10404,N_10250);
nand U10680 (N_10680,N_10324,N_10256);
and U10681 (N_10681,N_10241,N_10212);
and U10682 (N_10682,N_10225,N_10334);
xnor U10683 (N_10683,N_10476,N_10259);
and U10684 (N_10684,N_10398,N_10471);
nor U10685 (N_10685,N_10228,N_10497);
nor U10686 (N_10686,N_10321,N_10409);
nand U10687 (N_10687,N_10222,N_10372);
xor U10688 (N_10688,N_10465,N_10312);
xor U10689 (N_10689,N_10303,N_10265);
xnor U10690 (N_10690,N_10237,N_10404);
or U10691 (N_10691,N_10424,N_10340);
nand U10692 (N_10692,N_10317,N_10446);
and U10693 (N_10693,N_10246,N_10249);
and U10694 (N_10694,N_10292,N_10232);
nor U10695 (N_10695,N_10459,N_10473);
or U10696 (N_10696,N_10299,N_10392);
nor U10697 (N_10697,N_10461,N_10348);
nor U10698 (N_10698,N_10374,N_10340);
nand U10699 (N_10699,N_10352,N_10222);
nand U10700 (N_10700,N_10405,N_10235);
xor U10701 (N_10701,N_10342,N_10319);
and U10702 (N_10702,N_10219,N_10287);
nor U10703 (N_10703,N_10354,N_10444);
xnor U10704 (N_10704,N_10238,N_10441);
and U10705 (N_10705,N_10384,N_10379);
or U10706 (N_10706,N_10443,N_10311);
or U10707 (N_10707,N_10389,N_10456);
xnor U10708 (N_10708,N_10417,N_10291);
and U10709 (N_10709,N_10426,N_10432);
xor U10710 (N_10710,N_10224,N_10367);
xor U10711 (N_10711,N_10342,N_10244);
nor U10712 (N_10712,N_10266,N_10314);
and U10713 (N_10713,N_10421,N_10440);
nor U10714 (N_10714,N_10354,N_10464);
xnor U10715 (N_10715,N_10425,N_10489);
xor U10716 (N_10716,N_10343,N_10408);
xor U10717 (N_10717,N_10262,N_10272);
xor U10718 (N_10718,N_10298,N_10285);
nand U10719 (N_10719,N_10221,N_10226);
and U10720 (N_10720,N_10427,N_10346);
xnor U10721 (N_10721,N_10402,N_10235);
and U10722 (N_10722,N_10338,N_10496);
nand U10723 (N_10723,N_10361,N_10291);
xor U10724 (N_10724,N_10437,N_10331);
and U10725 (N_10725,N_10499,N_10387);
and U10726 (N_10726,N_10415,N_10451);
nor U10727 (N_10727,N_10265,N_10472);
nand U10728 (N_10728,N_10384,N_10324);
nor U10729 (N_10729,N_10486,N_10381);
xnor U10730 (N_10730,N_10447,N_10385);
nor U10731 (N_10731,N_10237,N_10341);
or U10732 (N_10732,N_10426,N_10331);
or U10733 (N_10733,N_10410,N_10242);
nand U10734 (N_10734,N_10219,N_10295);
nand U10735 (N_10735,N_10218,N_10264);
and U10736 (N_10736,N_10453,N_10245);
and U10737 (N_10737,N_10395,N_10262);
nand U10738 (N_10738,N_10377,N_10359);
nand U10739 (N_10739,N_10393,N_10431);
and U10740 (N_10740,N_10375,N_10222);
xnor U10741 (N_10741,N_10370,N_10233);
and U10742 (N_10742,N_10476,N_10438);
nand U10743 (N_10743,N_10483,N_10470);
nand U10744 (N_10744,N_10381,N_10477);
and U10745 (N_10745,N_10366,N_10298);
or U10746 (N_10746,N_10308,N_10497);
or U10747 (N_10747,N_10433,N_10401);
or U10748 (N_10748,N_10460,N_10386);
and U10749 (N_10749,N_10270,N_10271);
and U10750 (N_10750,N_10292,N_10467);
nand U10751 (N_10751,N_10205,N_10300);
nand U10752 (N_10752,N_10380,N_10208);
nor U10753 (N_10753,N_10387,N_10374);
xnor U10754 (N_10754,N_10470,N_10495);
nor U10755 (N_10755,N_10249,N_10281);
xnor U10756 (N_10756,N_10317,N_10213);
nand U10757 (N_10757,N_10204,N_10487);
xnor U10758 (N_10758,N_10298,N_10398);
xor U10759 (N_10759,N_10462,N_10212);
nand U10760 (N_10760,N_10219,N_10393);
nor U10761 (N_10761,N_10284,N_10286);
or U10762 (N_10762,N_10265,N_10427);
nand U10763 (N_10763,N_10265,N_10420);
nor U10764 (N_10764,N_10479,N_10449);
or U10765 (N_10765,N_10251,N_10451);
or U10766 (N_10766,N_10463,N_10221);
nand U10767 (N_10767,N_10436,N_10377);
nand U10768 (N_10768,N_10361,N_10353);
nor U10769 (N_10769,N_10446,N_10257);
or U10770 (N_10770,N_10330,N_10239);
nand U10771 (N_10771,N_10349,N_10334);
xor U10772 (N_10772,N_10248,N_10452);
nor U10773 (N_10773,N_10435,N_10425);
nor U10774 (N_10774,N_10261,N_10469);
xnor U10775 (N_10775,N_10349,N_10396);
nand U10776 (N_10776,N_10232,N_10437);
or U10777 (N_10777,N_10365,N_10267);
or U10778 (N_10778,N_10285,N_10356);
nand U10779 (N_10779,N_10422,N_10408);
and U10780 (N_10780,N_10476,N_10489);
nor U10781 (N_10781,N_10346,N_10312);
or U10782 (N_10782,N_10451,N_10219);
nor U10783 (N_10783,N_10254,N_10211);
xor U10784 (N_10784,N_10258,N_10321);
nand U10785 (N_10785,N_10491,N_10376);
nor U10786 (N_10786,N_10241,N_10490);
xor U10787 (N_10787,N_10292,N_10420);
nor U10788 (N_10788,N_10286,N_10327);
or U10789 (N_10789,N_10333,N_10483);
and U10790 (N_10790,N_10202,N_10371);
and U10791 (N_10791,N_10325,N_10423);
and U10792 (N_10792,N_10350,N_10453);
and U10793 (N_10793,N_10427,N_10352);
nor U10794 (N_10794,N_10398,N_10428);
xor U10795 (N_10795,N_10358,N_10264);
or U10796 (N_10796,N_10261,N_10408);
and U10797 (N_10797,N_10226,N_10425);
nand U10798 (N_10798,N_10469,N_10493);
or U10799 (N_10799,N_10263,N_10373);
xnor U10800 (N_10800,N_10579,N_10774);
or U10801 (N_10801,N_10730,N_10770);
nor U10802 (N_10802,N_10689,N_10562);
nor U10803 (N_10803,N_10655,N_10549);
nor U10804 (N_10804,N_10573,N_10600);
or U10805 (N_10805,N_10508,N_10768);
nor U10806 (N_10806,N_10656,N_10572);
nand U10807 (N_10807,N_10560,N_10668);
xor U10808 (N_10808,N_10649,N_10797);
or U10809 (N_10809,N_10603,N_10758);
nor U10810 (N_10810,N_10721,N_10773);
nand U10811 (N_10811,N_10561,N_10554);
and U10812 (N_10812,N_10651,N_10686);
and U10813 (N_10813,N_10687,N_10597);
and U10814 (N_10814,N_10644,N_10620);
or U10815 (N_10815,N_10747,N_10605);
nor U10816 (N_10816,N_10648,N_10776);
xnor U10817 (N_10817,N_10718,N_10639);
and U10818 (N_10818,N_10506,N_10581);
nand U10819 (N_10819,N_10567,N_10501);
or U10820 (N_10820,N_10624,N_10691);
xor U10821 (N_10821,N_10626,N_10729);
xor U10822 (N_10822,N_10673,N_10681);
nand U10823 (N_10823,N_10745,N_10539);
or U10824 (N_10824,N_10650,N_10688);
xnor U10825 (N_10825,N_10614,N_10515);
and U10826 (N_10826,N_10785,N_10552);
nand U10827 (N_10827,N_10739,N_10502);
xnor U10828 (N_10828,N_10748,N_10666);
xnor U10829 (N_10829,N_10728,N_10734);
and U10830 (N_10830,N_10698,N_10590);
or U10831 (N_10831,N_10667,N_10543);
nor U10832 (N_10832,N_10719,N_10665);
and U10833 (N_10833,N_10535,N_10727);
and U10834 (N_10834,N_10636,N_10680);
nand U10835 (N_10835,N_10537,N_10578);
and U10836 (N_10836,N_10787,N_10577);
or U10837 (N_10837,N_10763,N_10796);
or U10838 (N_10838,N_10596,N_10558);
nor U10839 (N_10839,N_10635,N_10643);
and U10840 (N_10840,N_10653,N_10602);
or U10841 (N_10841,N_10520,N_10557);
or U10842 (N_10842,N_10720,N_10753);
nand U10843 (N_10843,N_10793,N_10713);
nor U10844 (N_10844,N_10752,N_10780);
xor U10845 (N_10845,N_10692,N_10546);
or U10846 (N_10846,N_10791,N_10762);
and U10847 (N_10847,N_10675,N_10771);
nor U10848 (N_10848,N_10764,N_10783);
nor U10849 (N_10849,N_10725,N_10707);
nor U10850 (N_10850,N_10658,N_10664);
xor U10851 (N_10851,N_10786,N_10700);
or U10852 (N_10852,N_10576,N_10555);
nor U10853 (N_10853,N_10723,N_10531);
and U10854 (N_10854,N_10615,N_10732);
xnor U10855 (N_10855,N_10616,N_10663);
xor U10856 (N_10856,N_10659,N_10741);
or U10857 (N_10857,N_10618,N_10674);
or U10858 (N_10858,N_10592,N_10523);
nor U10859 (N_10859,N_10604,N_10799);
nor U10860 (N_10860,N_10740,N_10580);
nor U10861 (N_10861,N_10593,N_10583);
or U10862 (N_10862,N_10599,N_10755);
or U10863 (N_10863,N_10504,N_10622);
or U10864 (N_10864,N_10532,N_10705);
nor U10865 (N_10865,N_10777,N_10756);
nor U10866 (N_10866,N_10529,N_10696);
xnor U10867 (N_10867,N_10559,N_10789);
xor U10868 (N_10868,N_10714,N_10717);
nand U10869 (N_10869,N_10709,N_10566);
nand U10870 (N_10870,N_10556,N_10517);
xor U10871 (N_10871,N_10534,N_10676);
and U10872 (N_10872,N_10790,N_10631);
or U10873 (N_10873,N_10798,N_10574);
xor U10874 (N_10874,N_10536,N_10736);
nor U10875 (N_10875,N_10509,N_10779);
nand U10876 (N_10876,N_10512,N_10695);
or U10877 (N_10877,N_10704,N_10708);
xor U10878 (N_10878,N_10735,N_10570);
nor U10879 (N_10879,N_10661,N_10701);
xnor U10880 (N_10880,N_10652,N_10550);
or U10881 (N_10881,N_10654,N_10722);
nand U10882 (N_10882,N_10607,N_10611);
and U10883 (N_10883,N_10685,N_10519);
nor U10884 (N_10884,N_10571,N_10754);
xnor U10885 (N_10885,N_10724,N_10731);
nand U10886 (N_10886,N_10530,N_10660);
nand U10887 (N_10887,N_10795,N_10759);
and U10888 (N_10888,N_10540,N_10619);
and U10889 (N_10889,N_10778,N_10672);
xor U10890 (N_10890,N_10553,N_10744);
or U10891 (N_10891,N_10679,N_10563);
or U10892 (N_10892,N_10690,N_10684);
or U10893 (N_10893,N_10646,N_10591);
nor U10894 (N_10894,N_10609,N_10505);
nand U10895 (N_10895,N_10629,N_10575);
or U10896 (N_10896,N_10767,N_10595);
or U10897 (N_10897,N_10746,N_10533);
nand U10898 (N_10898,N_10683,N_10769);
xor U10899 (N_10899,N_10757,N_10784);
nand U10900 (N_10900,N_10742,N_10524);
nor U10901 (N_10901,N_10694,N_10706);
or U10902 (N_10902,N_10606,N_10510);
or U10903 (N_10903,N_10584,N_10548);
and U10904 (N_10904,N_10633,N_10640);
xor U10905 (N_10905,N_10612,N_10503);
nor U10906 (N_10906,N_10792,N_10677);
xor U10907 (N_10907,N_10772,N_10647);
nor U10908 (N_10908,N_10726,N_10628);
nand U10909 (N_10909,N_10585,N_10582);
and U10910 (N_10910,N_10551,N_10610);
and U10911 (N_10911,N_10662,N_10669);
or U10912 (N_10912,N_10794,N_10697);
or U10913 (N_10913,N_10547,N_10587);
nor U10914 (N_10914,N_10760,N_10637);
nor U10915 (N_10915,N_10598,N_10500);
nor U10916 (N_10916,N_10516,N_10528);
or U10917 (N_10917,N_10670,N_10613);
nand U10918 (N_10918,N_10711,N_10608);
xnor U10919 (N_10919,N_10627,N_10733);
and U10920 (N_10920,N_10565,N_10589);
nor U10921 (N_10921,N_10568,N_10716);
or U10922 (N_10922,N_10511,N_10541);
nand U10923 (N_10923,N_10586,N_10712);
xnor U10924 (N_10924,N_10751,N_10538);
and U10925 (N_10925,N_10542,N_10738);
nand U10926 (N_10926,N_10527,N_10743);
xor U10927 (N_10927,N_10630,N_10645);
nor U10928 (N_10928,N_10765,N_10678);
or U10929 (N_10929,N_10703,N_10715);
nor U10930 (N_10930,N_10588,N_10632);
nand U10931 (N_10931,N_10518,N_10569);
or U10932 (N_10932,N_10634,N_10710);
nor U10933 (N_10933,N_10625,N_10781);
nor U10934 (N_10934,N_10671,N_10545);
and U10935 (N_10935,N_10641,N_10682);
nor U10936 (N_10936,N_10617,N_10766);
nor U10937 (N_10937,N_10544,N_10514);
and U10938 (N_10938,N_10507,N_10522);
nor U10939 (N_10939,N_10601,N_10564);
nor U10940 (N_10940,N_10526,N_10693);
nand U10941 (N_10941,N_10699,N_10657);
xor U10942 (N_10942,N_10761,N_10750);
or U10943 (N_10943,N_10623,N_10775);
or U10944 (N_10944,N_10788,N_10525);
nor U10945 (N_10945,N_10749,N_10782);
and U10946 (N_10946,N_10702,N_10737);
or U10947 (N_10947,N_10513,N_10521);
and U10948 (N_10948,N_10621,N_10642);
and U10949 (N_10949,N_10638,N_10594);
or U10950 (N_10950,N_10719,N_10555);
and U10951 (N_10951,N_10678,N_10706);
nor U10952 (N_10952,N_10783,N_10665);
and U10953 (N_10953,N_10605,N_10636);
and U10954 (N_10954,N_10530,N_10600);
nor U10955 (N_10955,N_10782,N_10724);
or U10956 (N_10956,N_10525,N_10645);
xor U10957 (N_10957,N_10759,N_10785);
xor U10958 (N_10958,N_10639,N_10679);
nand U10959 (N_10959,N_10785,N_10587);
and U10960 (N_10960,N_10689,N_10592);
and U10961 (N_10961,N_10746,N_10684);
xor U10962 (N_10962,N_10522,N_10599);
or U10963 (N_10963,N_10798,N_10745);
or U10964 (N_10964,N_10758,N_10536);
xor U10965 (N_10965,N_10786,N_10553);
nand U10966 (N_10966,N_10746,N_10719);
nand U10967 (N_10967,N_10799,N_10761);
and U10968 (N_10968,N_10645,N_10585);
nand U10969 (N_10969,N_10591,N_10568);
or U10970 (N_10970,N_10524,N_10792);
and U10971 (N_10971,N_10756,N_10635);
nand U10972 (N_10972,N_10721,N_10650);
and U10973 (N_10973,N_10681,N_10543);
or U10974 (N_10974,N_10680,N_10511);
or U10975 (N_10975,N_10539,N_10709);
xnor U10976 (N_10976,N_10691,N_10611);
or U10977 (N_10977,N_10798,N_10513);
xnor U10978 (N_10978,N_10596,N_10590);
xor U10979 (N_10979,N_10790,N_10578);
xor U10980 (N_10980,N_10688,N_10735);
nor U10981 (N_10981,N_10652,N_10707);
nor U10982 (N_10982,N_10584,N_10596);
and U10983 (N_10983,N_10713,N_10566);
nand U10984 (N_10984,N_10518,N_10655);
nand U10985 (N_10985,N_10519,N_10737);
or U10986 (N_10986,N_10684,N_10572);
nor U10987 (N_10987,N_10685,N_10754);
nor U10988 (N_10988,N_10706,N_10604);
nor U10989 (N_10989,N_10601,N_10786);
nand U10990 (N_10990,N_10536,N_10513);
nand U10991 (N_10991,N_10556,N_10665);
xor U10992 (N_10992,N_10607,N_10676);
or U10993 (N_10993,N_10511,N_10625);
and U10994 (N_10994,N_10639,N_10743);
and U10995 (N_10995,N_10544,N_10538);
nor U10996 (N_10996,N_10581,N_10693);
or U10997 (N_10997,N_10729,N_10617);
nand U10998 (N_10998,N_10652,N_10635);
nand U10999 (N_10999,N_10677,N_10699);
nor U11000 (N_11000,N_10537,N_10583);
nor U11001 (N_11001,N_10729,N_10700);
nor U11002 (N_11002,N_10550,N_10541);
and U11003 (N_11003,N_10771,N_10732);
nor U11004 (N_11004,N_10540,N_10733);
and U11005 (N_11005,N_10660,N_10691);
nor U11006 (N_11006,N_10599,N_10552);
and U11007 (N_11007,N_10695,N_10746);
or U11008 (N_11008,N_10716,N_10629);
and U11009 (N_11009,N_10673,N_10714);
or U11010 (N_11010,N_10706,N_10647);
or U11011 (N_11011,N_10505,N_10522);
and U11012 (N_11012,N_10517,N_10574);
and U11013 (N_11013,N_10684,N_10522);
xnor U11014 (N_11014,N_10702,N_10704);
nor U11015 (N_11015,N_10689,N_10645);
and U11016 (N_11016,N_10553,N_10728);
nor U11017 (N_11017,N_10649,N_10544);
nor U11018 (N_11018,N_10627,N_10796);
nor U11019 (N_11019,N_10537,N_10561);
and U11020 (N_11020,N_10642,N_10682);
xnor U11021 (N_11021,N_10669,N_10722);
or U11022 (N_11022,N_10630,N_10676);
and U11023 (N_11023,N_10681,N_10591);
nor U11024 (N_11024,N_10795,N_10564);
and U11025 (N_11025,N_10738,N_10654);
and U11026 (N_11026,N_10700,N_10792);
nand U11027 (N_11027,N_10501,N_10684);
nor U11028 (N_11028,N_10604,N_10667);
xnor U11029 (N_11029,N_10657,N_10698);
xnor U11030 (N_11030,N_10526,N_10604);
or U11031 (N_11031,N_10608,N_10630);
nor U11032 (N_11032,N_10695,N_10545);
nor U11033 (N_11033,N_10594,N_10781);
nand U11034 (N_11034,N_10777,N_10504);
and U11035 (N_11035,N_10694,N_10521);
or U11036 (N_11036,N_10625,N_10575);
nand U11037 (N_11037,N_10503,N_10798);
nor U11038 (N_11038,N_10785,N_10682);
and U11039 (N_11039,N_10760,N_10575);
or U11040 (N_11040,N_10739,N_10656);
nand U11041 (N_11041,N_10680,N_10790);
xnor U11042 (N_11042,N_10639,N_10750);
and U11043 (N_11043,N_10619,N_10505);
nor U11044 (N_11044,N_10758,N_10557);
nor U11045 (N_11045,N_10758,N_10675);
xor U11046 (N_11046,N_10597,N_10784);
nor U11047 (N_11047,N_10754,N_10769);
and U11048 (N_11048,N_10733,N_10628);
nor U11049 (N_11049,N_10795,N_10619);
nand U11050 (N_11050,N_10587,N_10737);
or U11051 (N_11051,N_10717,N_10536);
xnor U11052 (N_11052,N_10699,N_10547);
nand U11053 (N_11053,N_10528,N_10673);
xor U11054 (N_11054,N_10595,N_10534);
nand U11055 (N_11055,N_10573,N_10700);
nor U11056 (N_11056,N_10510,N_10547);
nor U11057 (N_11057,N_10513,N_10591);
and U11058 (N_11058,N_10542,N_10559);
nor U11059 (N_11059,N_10721,N_10659);
or U11060 (N_11060,N_10604,N_10688);
nand U11061 (N_11061,N_10737,N_10535);
or U11062 (N_11062,N_10518,N_10560);
and U11063 (N_11063,N_10643,N_10589);
nand U11064 (N_11064,N_10586,N_10582);
and U11065 (N_11065,N_10569,N_10661);
xnor U11066 (N_11066,N_10770,N_10502);
nor U11067 (N_11067,N_10573,N_10750);
nor U11068 (N_11068,N_10593,N_10628);
xnor U11069 (N_11069,N_10776,N_10712);
nor U11070 (N_11070,N_10779,N_10656);
or U11071 (N_11071,N_10688,N_10543);
nor U11072 (N_11072,N_10794,N_10656);
nand U11073 (N_11073,N_10662,N_10682);
nand U11074 (N_11074,N_10628,N_10575);
or U11075 (N_11075,N_10699,N_10765);
and U11076 (N_11076,N_10586,N_10754);
or U11077 (N_11077,N_10508,N_10722);
and U11078 (N_11078,N_10563,N_10769);
nand U11079 (N_11079,N_10727,N_10689);
or U11080 (N_11080,N_10615,N_10525);
and U11081 (N_11081,N_10658,N_10524);
and U11082 (N_11082,N_10797,N_10783);
nor U11083 (N_11083,N_10557,N_10787);
xor U11084 (N_11084,N_10760,N_10553);
and U11085 (N_11085,N_10599,N_10505);
xnor U11086 (N_11086,N_10753,N_10700);
nand U11087 (N_11087,N_10771,N_10517);
xnor U11088 (N_11088,N_10676,N_10658);
and U11089 (N_11089,N_10573,N_10641);
nor U11090 (N_11090,N_10781,N_10639);
nor U11091 (N_11091,N_10563,N_10577);
and U11092 (N_11092,N_10539,N_10665);
nor U11093 (N_11093,N_10596,N_10791);
nand U11094 (N_11094,N_10634,N_10760);
and U11095 (N_11095,N_10581,N_10620);
and U11096 (N_11096,N_10765,N_10557);
nor U11097 (N_11097,N_10754,N_10659);
xor U11098 (N_11098,N_10582,N_10652);
nor U11099 (N_11099,N_10516,N_10668);
or U11100 (N_11100,N_10900,N_10952);
xor U11101 (N_11101,N_10846,N_10940);
xnor U11102 (N_11102,N_10841,N_11087);
and U11103 (N_11103,N_10977,N_11042);
xor U11104 (N_11104,N_11099,N_11075);
nor U11105 (N_11105,N_10995,N_11048);
nand U11106 (N_11106,N_11093,N_11058);
nand U11107 (N_11107,N_11022,N_10902);
or U11108 (N_11108,N_10849,N_11019);
xnor U11109 (N_11109,N_10853,N_11068);
nand U11110 (N_11110,N_10811,N_10883);
nor U11111 (N_11111,N_11043,N_11054);
nor U11112 (N_11112,N_10852,N_11066);
xor U11113 (N_11113,N_11079,N_10978);
and U11114 (N_11114,N_11070,N_10869);
or U11115 (N_11115,N_11074,N_11053);
nor U11116 (N_11116,N_10817,N_11050);
or U11117 (N_11117,N_10968,N_10868);
nor U11118 (N_11118,N_11055,N_10971);
nand U11119 (N_11119,N_11085,N_10974);
and U11120 (N_11120,N_10939,N_10864);
or U11121 (N_11121,N_10956,N_11064);
or U11122 (N_11122,N_10930,N_10943);
nand U11123 (N_11123,N_10962,N_10861);
and U11124 (N_11124,N_10865,N_10858);
or U11125 (N_11125,N_10808,N_11098);
nand U11126 (N_11126,N_10907,N_10945);
and U11127 (N_11127,N_10891,N_11045);
and U11128 (N_11128,N_10917,N_11038);
and U11129 (N_11129,N_10910,N_10921);
nor U11130 (N_11130,N_10908,N_11051);
xnor U11131 (N_11131,N_11060,N_11002);
nor U11132 (N_11132,N_11052,N_10965);
nand U11133 (N_11133,N_11044,N_10862);
nand U11134 (N_11134,N_10975,N_10879);
and U11135 (N_11135,N_10827,N_10876);
nor U11136 (N_11136,N_10806,N_10980);
nand U11137 (N_11137,N_10961,N_10816);
xor U11138 (N_11138,N_10922,N_11035);
or U11139 (N_11139,N_11014,N_10923);
nand U11140 (N_11140,N_11011,N_11026);
or U11141 (N_11141,N_10957,N_11057);
and U11142 (N_11142,N_10912,N_11004);
and U11143 (N_11143,N_11006,N_10969);
nand U11144 (N_11144,N_10814,N_11024);
nand U11145 (N_11145,N_10855,N_10958);
and U11146 (N_11146,N_10889,N_11012);
nor U11147 (N_11147,N_11062,N_11061);
and U11148 (N_11148,N_10914,N_11027);
xnor U11149 (N_11149,N_11016,N_10805);
nand U11150 (N_11150,N_10916,N_10938);
or U11151 (N_11151,N_11088,N_10821);
or U11152 (N_11152,N_10898,N_11095);
xor U11153 (N_11153,N_10904,N_10870);
nor U11154 (N_11154,N_10949,N_10990);
xor U11155 (N_11155,N_11056,N_10899);
nand U11156 (N_11156,N_10931,N_10934);
xor U11157 (N_11157,N_11063,N_11037);
and U11158 (N_11158,N_11017,N_10860);
nor U11159 (N_11159,N_10873,N_10982);
xor U11160 (N_11160,N_11008,N_10963);
nand U11161 (N_11161,N_10839,N_10972);
and U11162 (N_11162,N_10925,N_10813);
nand U11163 (N_11163,N_10818,N_11097);
xor U11164 (N_11164,N_10911,N_11072);
xnor U11165 (N_11165,N_10843,N_10913);
and U11166 (N_11166,N_10997,N_10953);
nand U11167 (N_11167,N_11090,N_10906);
nor U11168 (N_11168,N_10820,N_10847);
nor U11169 (N_11169,N_11015,N_10800);
and U11170 (N_11170,N_11029,N_10988);
nand U11171 (N_11171,N_10944,N_11071);
nor U11172 (N_11172,N_10840,N_10823);
xnor U11173 (N_11173,N_10863,N_10915);
nand U11174 (N_11174,N_10802,N_10801);
nor U11175 (N_11175,N_10892,N_11034);
and U11176 (N_11176,N_10881,N_10960);
or U11177 (N_11177,N_10948,N_10896);
nand U11178 (N_11178,N_11080,N_11041);
and U11179 (N_11179,N_11023,N_10893);
xor U11180 (N_11180,N_10959,N_10924);
nand U11181 (N_11181,N_10822,N_10920);
nor U11182 (N_11182,N_10829,N_11078);
nor U11183 (N_11183,N_10973,N_10832);
or U11184 (N_11184,N_10866,N_10828);
nor U11185 (N_11185,N_11081,N_11047);
nand U11186 (N_11186,N_10901,N_10985);
nand U11187 (N_11187,N_10854,N_10897);
nor U11188 (N_11188,N_10935,N_10964);
nand U11189 (N_11189,N_10903,N_10986);
and U11190 (N_11190,N_11036,N_10989);
or U11191 (N_11191,N_10836,N_10880);
and U11192 (N_11192,N_10947,N_10888);
nand U11193 (N_11193,N_10936,N_10951);
and U11194 (N_11194,N_10937,N_10992);
nor U11195 (N_11195,N_10926,N_10838);
or U11196 (N_11196,N_10927,N_11032);
nand U11197 (N_11197,N_11073,N_10842);
or U11198 (N_11198,N_10857,N_10890);
nor U11199 (N_11199,N_10966,N_10812);
nor U11200 (N_11200,N_11028,N_11076);
or U11201 (N_11201,N_11065,N_10918);
or U11202 (N_11202,N_11082,N_11030);
or U11203 (N_11203,N_10983,N_10874);
or U11204 (N_11204,N_10871,N_11086);
and U11205 (N_11205,N_10810,N_11084);
and U11206 (N_11206,N_10875,N_11013);
xor U11207 (N_11207,N_10848,N_10878);
xor U11208 (N_11208,N_10809,N_10844);
nand U11209 (N_11209,N_10885,N_10803);
or U11210 (N_11210,N_10970,N_11067);
nor U11211 (N_11211,N_10877,N_11096);
and U11212 (N_11212,N_10994,N_10967);
xor U11213 (N_11213,N_10942,N_10987);
and U11214 (N_11214,N_11000,N_11005);
and U11215 (N_11215,N_10976,N_10824);
nand U11216 (N_11216,N_11025,N_11094);
and U11217 (N_11217,N_11040,N_10835);
xnor U11218 (N_11218,N_10929,N_10845);
nand U11219 (N_11219,N_10932,N_10950);
or U11220 (N_11220,N_10815,N_10993);
xor U11221 (N_11221,N_11089,N_11033);
or U11222 (N_11222,N_10909,N_11001);
nand U11223 (N_11223,N_11039,N_10946);
nor U11224 (N_11224,N_10928,N_11031);
nand U11225 (N_11225,N_11046,N_10819);
xnor U11226 (N_11226,N_11020,N_10919);
and U11227 (N_11227,N_10984,N_10833);
nor U11228 (N_11228,N_10872,N_10999);
nor U11229 (N_11229,N_10905,N_10882);
xnor U11230 (N_11230,N_10850,N_11059);
or U11231 (N_11231,N_11092,N_11009);
nor U11232 (N_11232,N_11077,N_10834);
xnor U11233 (N_11233,N_11010,N_10886);
nor U11234 (N_11234,N_10837,N_10867);
xor U11235 (N_11235,N_10996,N_10831);
nand U11236 (N_11236,N_10991,N_10933);
nand U11237 (N_11237,N_11007,N_10856);
nor U11238 (N_11238,N_10955,N_10894);
nor U11239 (N_11239,N_10954,N_10830);
nor U11240 (N_11240,N_11049,N_10941);
nor U11241 (N_11241,N_10859,N_10979);
nand U11242 (N_11242,N_11021,N_10851);
nand U11243 (N_11243,N_11069,N_10825);
and U11244 (N_11244,N_10826,N_11091);
and U11245 (N_11245,N_11018,N_11003);
nand U11246 (N_11246,N_10807,N_11083);
xnor U11247 (N_11247,N_10998,N_10887);
xnor U11248 (N_11248,N_10884,N_10804);
nor U11249 (N_11249,N_10981,N_10895);
xor U11250 (N_11250,N_10996,N_10906);
xnor U11251 (N_11251,N_10934,N_10949);
nand U11252 (N_11252,N_10866,N_11043);
xor U11253 (N_11253,N_10933,N_10986);
xnor U11254 (N_11254,N_10891,N_11083);
xnor U11255 (N_11255,N_11010,N_11058);
or U11256 (N_11256,N_10986,N_11022);
nor U11257 (N_11257,N_10931,N_10855);
xor U11258 (N_11258,N_10811,N_11000);
xnor U11259 (N_11259,N_10821,N_10904);
xor U11260 (N_11260,N_11019,N_11010);
xnor U11261 (N_11261,N_11082,N_10807);
and U11262 (N_11262,N_11085,N_10939);
and U11263 (N_11263,N_10873,N_10997);
nand U11264 (N_11264,N_10910,N_10878);
nor U11265 (N_11265,N_10825,N_10952);
xor U11266 (N_11266,N_11034,N_11060);
xnor U11267 (N_11267,N_11033,N_10944);
nand U11268 (N_11268,N_10805,N_10945);
xnor U11269 (N_11269,N_11022,N_10865);
and U11270 (N_11270,N_10983,N_10976);
nand U11271 (N_11271,N_10915,N_10974);
or U11272 (N_11272,N_10934,N_11014);
nand U11273 (N_11273,N_11044,N_10859);
nor U11274 (N_11274,N_10817,N_10937);
xor U11275 (N_11275,N_10812,N_10866);
or U11276 (N_11276,N_10803,N_11068);
or U11277 (N_11277,N_10806,N_10939);
nand U11278 (N_11278,N_10883,N_11023);
nor U11279 (N_11279,N_10811,N_11068);
nor U11280 (N_11280,N_11008,N_10892);
nand U11281 (N_11281,N_11065,N_10870);
and U11282 (N_11282,N_10965,N_11010);
or U11283 (N_11283,N_11057,N_10862);
xnor U11284 (N_11284,N_10990,N_11033);
nand U11285 (N_11285,N_10997,N_10952);
xnor U11286 (N_11286,N_10948,N_10840);
xnor U11287 (N_11287,N_11094,N_11050);
xor U11288 (N_11288,N_10946,N_11090);
or U11289 (N_11289,N_11057,N_10851);
nor U11290 (N_11290,N_10857,N_10930);
nand U11291 (N_11291,N_10828,N_11025);
xnor U11292 (N_11292,N_10943,N_10898);
nor U11293 (N_11293,N_11007,N_11079);
and U11294 (N_11294,N_10910,N_11018);
nor U11295 (N_11295,N_11004,N_11016);
or U11296 (N_11296,N_10999,N_10807);
xnor U11297 (N_11297,N_10843,N_11055);
nand U11298 (N_11298,N_10825,N_10807);
xnor U11299 (N_11299,N_10843,N_11020);
nand U11300 (N_11300,N_10982,N_10999);
xnor U11301 (N_11301,N_10998,N_11002);
xor U11302 (N_11302,N_11061,N_11007);
xnor U11303 (N_11303,N_10820,N_10936);
nor U11304 (N_11304,N_10877,N_10933);
nand U11305 (N_11305,N_10935,N_10841);
nor U11306 (N_11306,N_10966,N_11035);
nor U11307 (N_11307,N_10929,N_10975);
nand U11308 (N_11308,N_10822,N_10917);
or U11309 (N_11309,N_11098,N_10957);
xor U11310 (N_11310,N_10965,N_11065);
and U11311 (N_11311,N_10882,N_10853);
nor U11312 (N_11312,N_10870,N_10960);
and U11313 (N_11313,N_10850,N_10852);
nor U11314 (N_11314,N_10823,N_11004);
nand U11315 (N_11315,N_10958,N_10912);
or U11316 (N_11316,N_10969,N_11067);
nor U11317 (N_11317,N_11024,N_10811);
and U11318 (N_11318,N_11080,N_10958);
and U11319 (N_11319,N_10936,N_10915);
nor U11320 (N_11320,N_10909,N_11044);
nand U11321 (N_11321,N_10866,N_11034);
or U11322 (N_11322,N_10898,N_10855);
or U11323 (N_11323,N_10833,N_11063);
xor U11324 (N_11324,N_11094,N_11083);
nand U11325 (N_11325,N_10852,N_11026);
nor U11326 (N_11326,N_11033,N_10839);
and U11327 (N_11327,N_10823,N_10901);
nor U11328 (N_11328,N_10928,N_10860);
nor U11329 (N_11329,N_11026,N_11028);
and U11330 (N_11330,N_10956,N_10994);
or U11331 (N_11331,N_10843,N_10847);
nand U11332 (N_11332,N_10824,N_11044);
nor U11333 (N_11333,N_10800,N_10950);
and U11334 (N_11334,N_11010,N_11090);
nor U11335 (N_11335,N_10952,N_10884);
nor U11336 (N_11336,N_10806,N_10873);
nor U11337 (N_11337,N_10861,N_10807);
nor U11338 (N_11338,N_11022,N_10834);
or U11339 (N_11339,N_11073,N_10819);
nor U11340 (N_11340,N_10980,N_10894);
xor U11341 (N_11341,N_10945,N_10814);
nor U11342 (N_11342,N_10917,N_10914);
xnor U11343 (N_11343,N_10964,N_11089);
nand U11344 (N_11344,N_11067,N_11018);
nor U11345 (N_11345,N_11034,N_10946);
nand U11346 (N_11346,N_10814,N_11084);
and U11347 (N_11347,N_10851,N_10850);
nor U11348 (N_11348,N_11027,N_10855);
xor U11349 (N_11349,N_10841,N_10902);
nor U11350 (N_11350,N_10922,N_10890);
xor U11351 (N_11351,N_10981,N_10811);
and U11352 (N_11352,N_10867,N_10949);
or U11353 (N_11353,N_11051,N_10869);
nor U11354 (N_11354,N_10832,N_11022);
nor U11355 (N_11355,N_10934,N_11062);
xor U11356 (N_11356,N_10995,N_10868);
or U11357 (N_11357,N_10973,N_10818);
and U11358 (N_11358,N_10902,N_10876);
xnor U11359 (N_11359,N_10850,N_11099);
or U11360 (N_11360,N_11045,N_10874);
or U11361 (N_11361,N_10843,N_11071);
nor U11362 (N_11362,N_10925,N_10820);
nor U11363 (N_11363,N_10969,N_10973);
and U11364 (N_11364,N_10909,N_11024);
xor U11365 (N_11365,N_11098,N_10992);
nor U11366 (N_11366,N_10870,N_10812);
and U11367 (N_11367,N_10981,N_11065);
or U11368 (N_11368,N_10844,N_10945);
nor U11369 (N_11369,N_10932,N_10848);
nand U11370 (N_11370,N_10858,N_11036);
and U11371 (N_11371,N_10857,N_10903);
nor U11372 (N_11372,N_10982,N_10896);
or U11373 (N_11373,N_10833,N_11083);
xor U11374 (N_11374,N_10916,N_10870);
nand U11375 (N_11375,N_11043,N_10964);
nor U11376 (N_11376,N_10995,N_11054);
or U11377 (N_11377,N_10965,N_10852);
nor U11378 (N_11378,N_10822,N_10907);
xnor U11379 (N_11379,N_11092,N_10968);
nand U11380 (N_11380,N_10834,N_10800);
nor U11381 (N_11381,N_10833,N_11068);
nand U11382 (N_11382,N_11051,N_10814);
xnor U11383 (N_11383,N_11011,N_10892);
nor U11384 (N_11384,N_11033,N_10836);
nand U11385 (N_11385,N_11076,N_10931);
nor U11386 (N_11386,N_10951,N_10928);
and U11387 (N_11387,N_10959,N_10929);
xor U11388 (N_11388,N_10892,N_11040);
nor U11389 (N_11389,N_10884,N_10826);
and U11390 (N_11390,N_10850,N_10821);
nor U11391 (N_11391,N_10925,N_10948);
nand U11392 (N_11392,N_11007,N_10939);
nor U11393 (N_11393,N_10942,N_10973);
xnor U11394 (N_11394,N_10871,N_10911);
nand U11395 (N_11395,N_10978,N_10997);
or U11396 (N_11396,N_10927,N_11058);
xor U11397 (N_11397,N_10822,N_10997);
xnor U11398 (N_11398,N_10845,N_10895);
and U11399 (N_11399,N_10990,N_11035);
and U11400 (N_11400,N_11343,N_11393);
xor U11401 (N_11401,N_11316,N_11177);
nand U11402 (N_11402,N_11300,N_11203);
xnor U11403 (N_11403,N_11315,N_11367);
nor U11404 (N_11404,N_11277,N_11171);
nand U11405 (N_11405,N_11180,N_11299);
or U11406 (N_11406,N_11135,N_11115);
nor U11407 (N_11407,N_11149,N_11228);
xor U11408 (N_11408,N_11298,N_11339);
nand U11409 (N_11409,N_11118,N_11244);
nor U11410 (N_11410,N_11133,N_11100);
nand U11411 (N_11411,N_11161,N_11108);
or U11412 (N_11412,N_11188,N_11119);
or U11413 (N_11413,N_11190,N_11282);
nand U11414 (N_11414,N_11385,N_11372);
nand U11415 (N_11415,N_11317,N_11296);
nand U11416 (N_11416,N_11301,N_11327);
nand U11417 (N_11417,N_11205,N_11279);
or U11418 (N_11418,N_11332,N_11304);
nand U11419 (N_11419,N_11318,N_11158);
xnor U11420 (N_11420,N_11348,N_11284);
nor U11421 (N_11421,N_11355,N_11107);
nor U11422 (N_11422,N_11183,N_11346);
nor U11423 (N_11423,N_11261,N_11210);
and U11424 (N_11424,N_11106,N_11379);
nand U11425 (N_11425,N_11237,N_11248);
xnor U11426 (N_11426,N_11249,N_11386);
xor U11427 (N_11427,N_11394,N_11251);
nor U11428 (N_11428,N_11280,N_11159);
and U11429 (N_11429,N_11314,N_11223);
nand U11430 (N_11430,N_11287,N_11169);
nand U11431 (N_11431,N_11303,N_11270);
or U11432 (N_11432,N_11285,N_11233);
and U11433 (N_11433,N_11232,N_11260);
or U11434 (N_11434,N_11306,N_11241);
xor U11435 (N_11435,N_11142,N_11143);
or U11436 (N_11436,N_11396,N_11224);
and U11437 (N_11437,N_11189,N_11139);
and U11438 (N_11438,N_11330,N_11154);
or U11439 (N_11439,N_11112,N_11371);
and U11440 (N_11440,N_11256,N_11365);
or U11441 (N_11441,N_11229,N_11218);
and U11442 (N_11442,N_11352,N_11195);
nor U11443 (N_11443,N_11297,N_11322);
nor U11444 (N_11444,N_11354,N_11212);
and U11445 (N_11445,N_11114,N_11377);
or U11446 (N_11446,N_11311,N_11290);
and U11447 (N_11447,N_11240,N_11364);
and U11448 (N_11448,N_11344,N_11383);
nor U11449 (N_11449,N_11324,N_11321);
nor U11450 (N_11450,N_11333,N_11358);
xnor U11451 (N_11451,N_11312,N_11341);
xnor U11452 (N_11452,N_11391,N_11199);
and U11453 (N_11453,N_11124,N_11225);
and U11454 (N_11454,N_11201,N_11347);
nand U11455 (N_11455,N_11216,N_11234);
nand U11456 (N_11456,N_11144,N_11274);
nand U11457 (N_11457,N_11289,N_11325);
nand U11458 (N_11458,N_11208,N_11313);
xnor U11459 (N_11459,N_11104,N_11271);
nand U11460 (N_11460,N_11126,N_11369);
xor U11461 (N_11461,N_11309,N_11226);
and U11462 (N_11462,N_11121,N_11160);
or U11463 (N_11463,N_11388,N_11227);
or U11464 (N_11464,N_11140,N_11239);
nor U11465 (N_11465,N_11384,N_11141);
xor U11466 (N_11466,N_11340,N_11138);
xor U11467 (N_11467,N_11136,N_11254);
nand U11468 (N_11468,N_11250,N_11310);
xor U11469 (N_11469,N_11191,N_11117);
nor U11470 (N_11470,N_11127,N_11185);
or U11471 (N_11471,N_11276,N_11123);
xnor U11472 (N_11472,N_11157,N_11168);
xnor U11473 (N_11473,N_11389,N_11176);
nand U11474 (N_11474,N_11258,N_11192);
or U11475 (N_11475,N_11302,N_11174);
xnor U11476 (N_11476,N_11231,N_11253);
nand U11477 (N_11477,N_11272,N_11281);
nor U11478 (N_11478,N_11204,N_11334);
and U11479 (N_11479,N_11328,N_11378);
nor U11480 (N_11480,N_11235,N_11266);
nand U11481 (N_11481,N_11246,N_11278);
xor U11482 (N_11482,N_11150,N_11152);
and U11483 (N_11483,N_11375,N_11392);
or U11484 (N_11484,N_11387,N_11214);
or U11485 (N_11485,N_11390,N_11326);
xor U11486 (N_11486,N_11172,N_11398);
xnor U11487 (N_11487,N_11275,N_11202);
or U11488 (N_11488,N_11320,N_11166);
or U11489 (N_11489,N_11292,N_11363);
and U11490 (N_11490,N_11101,N_11353);
nor U11491 (N_11491,N_11103,N_11175);
xnor U11492 (N_11492,N_11257,N_11259);
xnor U11493 (N_11493,N_11220,N_11145);
nand U11494 (N_11494,N_11197,N_11156);
nand U11495 (N_11495,N_11273,N_11360);
and U11496 (N_11496,N_11151,N_11155);
nor U11497 (N_11497,N_11267,N_11213);
xnor U11498 (N_11498,N_11111,N_11336);
xor U11499 (N_11499,N_11230,N_11359);
xnor U11500 (N_11500,N_11295,N_11373);
xnor U11501 (N_11501,N_11262,N_11342);
nand U11502 (N_11502,N_11194,N_11370);
nor U11503 (N_11503,N_11263,N_11397);
xnor U11504 (N_11504,N_11198,N_11288);
and U11505 (N_11505,N_11120,N_11215);
nand U11506 (N_11506,N_11128,N_11366);
or U11507 (N_11507,N_11132,N_11187);
nor U11508 (N_11508,N_11335,N_11293);
xnor U11509 (N_11509,N_11147,N_11247);
nor U11510 (N_11510,N_11178,N_11102);
nand U11511 (N_11511,N_11268,N_11269);
nand U11512 (N_11512,N_11173,N_11125);
nand U11513 (N_11513,N_11146,N_11356);
nand U11514 (N_11514,N_11308,N_11170);
nor U11515 (N_11515,N_11162,N_11362);
nand U11516 (N_11516,N_11376,N_11323);
nand U11517 (N_11517,N_11222,N_11209);
and U11518 (N_11518,N_11129,N_11153);
nor U11519 (N_11519,N_11165,N_11164);
and U11520 (N_11520,N_11167,N_11380);
nor U11521 (N_11521,N_11395,N_11350);
nand U11522 (N_11522,N_11374,N_11345);
nor U11523 (N_11523,N_11184,N_11109);
and U11524 (N_11524,N_11179,N_11105);
xor U11525 (N_11525,N_11148,N_11283);
nor U11526 (N_11526,N_11286,N_11181);
or U11527 (N_11527,N_11245,N_11382);
nand U11528 (N_11528,N_11134,N_11221);
and U11529 (N_11529,N_11338,N_11381);
or U11530 (N_11530,N_11242,N_11329);
nand U11531 (N_11531,N_11130,N_11211);
xnor U11532 (N_11532,N_11264,N_11200);
and U11533 (N_11533,N_11331,N_11243);
nor U11534 (N_11534,N_11294,N_11351);
nor U11535 (N_11535,N_11238,N_11131);
xnor U11536 (N_11536,N_11305,N_11116);
and U11537 (N_11537,N_11113,N_11217);
and U11538 (N_11538,N_11337,N_11207);
nor U11539 (N_11539,N_11255,N_11399);
xnor U11540 (N_11540,N_11110,N_11163);
xnor U11541 (N_11541,N_11252,N_11122);
nand U11542 (N_11542,N_11357,N_11265);
nor U11543 (N_11543,N_11137,N_11186);
xnor U11544 (N_11544,N_11368,N_11307);
nand U11545 (N_11545,N_11193,N_11182);
or U11546 (N_11546,N_11361,N_11206);
and U11547 (N_11547,N_11319,N_11236);
xnor U11548 (N_11548,N_11291,N_11219);
nand U11549 (N_11549,N_11196,N_11349);
xnor U11550 (N_11550,N_11148,N_11274);
or U11551 (N_11551,N_11335,N_11107);
or U11552 (N_11552,N_11305,N_11208);
or U11553 (N_11553,N_11324,N_11137);
or U11554 (N_11554,N_11176,N_11222);
xnor U11555 (N_11555,N_11353,N_11106);
nor U11556 (N_11556,N_11353,N_11189);
nand U11557 (N_11557,N_11203,N_11344);
or U11558 (N_11558,N_11232,N_11175);
xor U11559 (N_11559,N_11174,N_11346);
xor U11560 (N_11560,N_11344,N_11182);
xnor U11561 (N_11561,N_11383,N_11161);
nor U11562 (N_11562,N_11134,N_11114);
nand U11563 (N_11563,N_11382,N_11219);
xnor U11564 (N_11564,N_11256,N_11384);
nor U11565 (N_11565,N_11146,N_11246);
nor U11566 (N_11566,N_11383,N_11146);
and U11567 (N_11567,N_11132,N_11167);
and U11568 (N_11568,N_11333,N_11235);
xor U11569 (N_11569,N_11200,N_11305);
nor U11570 (N_11570,N_11214,N_11393);
and U11571 (N_11571,N_11205,N_11112);
nor U11572 (N_11572,N_11360,N_11315);
xor U11573 (N_11573,N_11334,N_11171);
or U11574 (N_11574,N_11386,N_11217);
xor U11575 (N_11575,N_11272,N_11122);
or U11576 (N_11576,N_11197,N_11200);
or U11577 (N_11577,N_11205,N_11357);
xor U11578 (N_11578,N_11319,N_11198);
and U11579 (N_11579,N_11260,N_11393);
nor U11580 (N_11580,N_11268,N_11368);
and U11581 (N_11581,N_11212,N_11368);
nor U11582 (N_11582,N_11275,N_11390);
nor U11583 (N_11583,N_11357,N_11388);
or U11584 (N_11584,N_11187,N_11314);
and U11585 (N_11585,N_11395,N_11260);
nor U11586 (N_11586,N_11134,N_11212);
xnor U11587 (N_11587,N_11209,N_11298);
nor U11588 (N_11588,N_11323,N_11169);
and U11589 (N_11589,N_11135,N_11298);
xnor U11590 (N_11590,N_11385,N_11388);
xor U11591 (N_11591,N_11174,N_11199);
xnor U11592 (N_11592,N_11302,N_11372);
and U11593 (N_11593,N_11237,N_11311);
nand U11594 (N_11594,N_11275,N_11279);
or U11595 (N_11595,N_11134,N_11346);
xnor U11596 (N_11596,N_11216,N_11248);
and U11597 (N_11597,N_11358,N_11386);
or U11598 (N_11598,N_11167,N_11375);
or U11599 (N_11599,N_11245,N_11160);
xor U11600 (N_11600,N_11178,N_11338);
and U11601 (N_11601,N_11237,N_11280);
xnor U11602 (N_11602,N_11299,N_11268);
and U11603 (N_11603,N_11179,N_11331);
nor U11604 (N_11604,N_11203,N_11272);
xor U11605 (N_11605,N_11362,N_11165);
nand U11606 (N_11606,N_11334,N_11225);
or U11607 (N_11607,N_11143,N_11357);
xor U11608 (N_11608,N_11104,N_11229);
xor U11609 (N_11609,N_11335,N_11238);
nand U11610 (N_11610,N_11202,N_11374);
nand U11611 (N_11611,N_11309,N_11304);
xor U11612 (N_11612,N_11349,N_11383);
and U11613 (N_11613,N_11342,N_11381);
or U11614 (N_11614,N_11240,N_11350);
xor U11615 (N_11615,N_11318,N_11340);
nor U11616 (N_11616,N_11299,N_11110);
and U11617 (N_11617,N_11242,N_11174);
and U11618 (N_11618,N_11148,N_11320);
and U11619 (N_11619,N_11190,N_11208);
nand U11620 (N_11620,N_11270,N_11275);
nor U11621 (N_11621,N_11357,N_11178);
nand U11622 (N_11622,N_11306,N_11138);
xnor U11623 (N_11623,N_11272,N_11278);
and U11624 (N_11624,N_11339,N_11104);
xnor U11625 (N_11625,N_11120,N_11373);
and U11626 (N_11626,N_11130,N_11100);
nor U11627 (N_11627,N_11119,N_11147);
xnor U11628 (N_11628,N_11162,N_11302);
nor U11629 (N_11629,N_11384,N_11207);
and U11630 (N_11630,N_11328,N_11383);
and U11631 (N_11631,N_11342,N_11232);
or U11632 (N_11632,N_11332,N_11242);
or U11633 (N_11633,N_11205,N_11174);
or U11634 (N_11634,N_11274,N_11297);
xor U11635 (N_11635,N_11352,N_11137);
or U11636 (N_11636,N_11354,N_11279);
or U11637 (N_11637,N_11103,N_11257);
nor U11638 (N_11638,N_11345,N_11304);
nor U11639 (N_11639,N_11203,N_11349);
nor U11640 (N_11640,N_11299,N_11363);
nor U11641 (N_11641,N_11354,N_11285);
or U11642 (N_11642,N_11343,N_11134);
nand U11643 (N_11643,N_11237,N_11136);
nor U11644 (N_11644,N_11213,N_11385);
xnor U11645 (N_11645,N_11212,N_11100);
and U11646 (N_11646,N_11137,N_11250);
nor U11647 (N_11647,N_11200,N_11377);
or U11648 (N_11648,N_11322,N_11374);
nand U11649 (N_11649,N_11347,N_11113);
or U11650 (N_11650,N_11134,N_11176);
nand U11651 (N_11651,N_11395,N_11285);
or U11652 (N_11652,N_11364,N_11109);
xnor U11653 (N_11653,N_11327,N_11104);
xor U11654 (N_11654,N_11384,N_11324);
nand U11655 (N_11655,N_11349,N_11174);
nor U11656 (N_11656,N_11103,N_11185);
and U11657 (N_11657,N_11211,N_11143);
and U11658 (N_11658,N_11128,N_11152);
xnor U11659 (N_11659,N_11268,N_11363);
or U11660 (N_11660,N_11145,N_11106);
nand U11661 (N_11661,N_11353,N_11263);
nor U11662 (N_11662,N_11129,N_11319);
nor U11663 (N_11663,N_11214,N_11116);
and U11664 (N_11664,N_11151,N_11222);
or U11665 (N_11665,N_11221,N_11294);
xnor U11666 (N_11666,N_11167,N_11101);
nor U11667 (N_11667,N_11241,N_11356);
or U11668 (N_11668,N_11251,N_11376);
xor U11669 (N_11669,N_11239,N_11376);
or U11670 (N_11670,N_11340,N_11104);
or U11671 (N_11671,N_11129,N_11318);
or U11672 (N_11672,N_11187,N_11159);
or U11673 (N_11673,N_11318,N_11232);
nand U11674 (N_11674,N_11389,N_11390);
xor U11675 (N_11675,N_11187,N_11374);
nor U11676 (N_11676,N_11214,N_11268);
nand U11677 (N_11677,N_11323,N_11191);
xor U11678 (N_11678,N_11322,N_11270);
nor U11679 (N_11679,N_11150,N_11193);
xnor U11680 (N_11680,N_11274,N_11223);
xnor U11681 (N_11681,N_11259,N_11185);
nor U11682 (N_11682,N_11124,N_11303);
and U11683 (N_11683,N_11325,N_11393);
nor U11684 (N_11684,N_11256,N_11101);
or U11685 (N_11685,N_11132,N_11152);
and U11686 (N_11686,N_11295,N_11253);
or U11687 (N_11687,N_11264,N_11361);
nor U11688 (N_11688,N_11348,N_11242);
xnor U11689 (N_11689,N_11252,N_11204);
and U11690 (N_11690,N_11264,N_11151);
nand U11691 (N_11691,N_11333,N_11386);
nand U11692 (N_11692,N_11155,N_11252);
and U11693 (N_11693,N_11377,N_11233);
and U11694 (N_11694,N_11254,N_11288);
or U11695 (N_11695,N_11205,N_11238);
and U11696 (N_11696,N_11293,N_11237);
or U11697 (N_11697,N_11385,N_11145);
and U11698 (N_11698,N_11175,N_11110);
or U11699 (N_11699,N_11238,N_11106);
xnor U11700 (N_11700,N_11631,N_11665);
xor U11701 (N_11701,N_11645,N_11416);
nand U11702 (N_11702,N_11550,N_11411);
and U11703 (N_11703,N_11519,N_11441);
nor U11704 (N_11704,N_11636,N_11696);
nor U11705 (N_11705,N_11470,N_11415);
and U11706 (N_11706,N_11684,N_11567);
nor U11707 (N_11707,N_11449,N_11689);
and U11708 (N_11708,N_11571,N_11431);
and U11709 (N_11709,N_11646,N_11420);
nand U11710 (N_11710,N_11545,N_11452);
nor U11711 (N_11711,N_11474,N_11616);
or U11712 (N_11712,N_11456,N_11419);
nor U11713 (N_11713,N_11609,N_11464);
and U11714 (N_11714,N_11561,N_11598);
and U11715 (N_11715,N_11466,N_11542);
nor U11716 (N_11716,N_11418,N_11403);
nand U11717 (N_11717,N_11534,N_11683);
and U11718 (N_11718,N_11490,N_11435);
nand U11719 (N_11719,N_11507,N_11671);
nand U11720 (N_11720,N_11544,N_11642);
nand U11721 (N_11721,N_11572,N_11543);
and U11722 (N_11722,N_11670,N_11552);
xor U11723 (N_11723,N_11436,N_11607);
or U11724 (N_11724,N_11653,N_11469);
nor U11725 (N_11725,N_11502,N_11667);
and U11726 (N_11726,N_11460,N_11629);
or U11727 (N_11727,N_11639,N_11555);
nor U11728 (N_11728,N_11424,N_11593);
nand U11729 (N_11729,N_11495,N_11663);
or U11730 (N_11730,N_11672,N_11549);
and U11731 (N_11731,N_11638,N_11491);
or U11732 (N_11732,N_11473,N_11658);
or U11733 (N_11733,N_11660,N_11613);
and U11734 (N_11734,N_11486,N_11509);
and U11735 (N_11735,N_11527,N_11581);
nor U11736 (N_11736,N_11566,N_11513);
or U11737 (N_11737,N_11476,N_11569);
xnor U11738 (N_11738,N_11429,N_11493);
and U11739 (N_11739,N_11468,N_11668);
and U11740 (N_11740,N_11654,N_11414);
nand U11741 (N_11741,N_11485,N_11422);
nor U11742 (N_11742,N_11535,N_11676);
and U11743 (N_11743,N_11624,N_11650);
nand U11744 (N_11744,N_11462,N_11536);
nor U11745 (N_11745,N_11632,N_11529);
and U11746 (N_11746,N_11589,N_11582);
nor U11747 (N_11747,N_11587,N_11596);
nor U11748 (N_11748,N_11546,N_11408);
nand U11749 (N_11749,N_11659,N_11517);
nor U11750 (N_11750,N_11506,N_11438);
nand U11751 (N_11751,N_11447,N_11463);
nor U11752 (N_11752,N_11532,N_11677);
nand U11753 (N_11753,N_11565,N_11558);
xnor U11754 (N_11754,N_11608,N_11487);
nand U11755 (N_11755,N_11538,N_11475);
nand U11756 (N_11756,N_11514,N_11649);
or U11757 (N_11757,N_11401,N_11610);
and U11758 (N_11758,N_11526,N_11410);
nand U11759 (N_11759,N_11619,N_11553);
xor U11760 (N_11760,N_11459,N_11691);
xor U11761 (N_11761,N_11568,N_11563);
nand U11762 (N_11762,N_11580,N_11625);
or U11763 (N_11763,N_11597,N_11427);
nand U11764 (N_11764,N_11515,N_11467);
or U11765 (N_11765,N_11407,N_11451);
and U11766 (N_11766,N_11617,N_11477);
nor U11767 (N_11767,N_11655,N_11694);
or U11768 (N_11768,N_11674,N_11405);
nand U11769 (N_11769,N_11461,N_11618);
nand U11770 (N_11770,N_11530,N_11637);
nor U11771 (N_11771,N_11426,N_11522);
nor U11772 (N_11772,N_11564,N_11577);
nand U11773 (N_11773,N_11661,N_11578);
nor U11774 (N_11774,N_11524,N_11400);
xor U11775 (N_11775,N_11453,N_11444);
nor U11776 (N_11776,N_11611,N_11657);
and U11777 (N_11777,N_11479,N_11425);
xor U11778 (N_11778,N_11688,N_11471);
nand U11779 (N_11779,N_11647,N_11521);
nor U11780 (N_11780,N_11409,N_11523);
nor U11781 (N_11781,N_11573,N_11533);
xor U11782 (N_11782,N_11501,N_11525);
and U11783 (N_11783,N_11586,N_11455);
nand U11784 (N_11784,N_11579,N_11628);
nand U11785 (N_11785,N_11559,N_11622);
xnor U11786 (N_11786,N_11627,N_11417);
nand U11787 (N_11787,N_11458,N_11584);
nand U11788 (N_11788,N_11500,N_11504);
xor U11789 (N_11789,N_11432,N_11673);
nand U11790 (N_11790,N_11621,N_11595);
nor U11791 (N_11791,N_11556,N_11472);
or U11792 (N_11792,N_11412,N_11434);
and U11793 (N_11793,N_11592,N_11406);
and U11794 (N_11794,N_11574,N_11454);
xor U11795 (N_11795,N_11531,N_11560);
nand U11796 (N_11796,N_11539,N_11442);
nor U11797 (N_11797,N_11685,N_11600);
and U11798 (N_11798,N_11481,N_11575);
nor U11799 (N_11799,N_11644,N_11602);
nand U11800 (N_11800,N_11433,N_11488);
or U11801 (N_11801,N_11604,N_11465);
nand U11802 (N_11802,N_11623,N_11498);
nand U11803 (N_11803,N_11428,N_11497);
xor U11804 (N_11804,N_11537,N_11499);
or U11805 (N_11805,N_11640,N_11554);
and U11806 (N_11806,N_11496,N_11520);
nor U11807 (N_11807,N_11675,N_11682);
nor U11808 (N_11808,N_11457,N_11570);
or U11809 (N_11809,N_11599,N_11666);
nand U11810 (N_11810,N_11620,N_11615);
nand U11811 (N_11811,N_11430,N_11678);
nand U11812 (N_11812,N_11698,N_11562);
nor U11813 (N_11813,N_11445,N_11695);
or U11814 (N_11814,N_11651,N_11633);
xor U11815 (N_11815,N_11494,N_11512);
xnor U11816 (N_11816,N_11656,N_11478);
nor U11817 (N_11817,N_11503,N_11630);
and U11818 (N_11818,N_11483,N_11489);
xor U11819 (N_11819,N_11635,N_11626);
and U11820 (N_11820,N_11641,N_11583);
nor U11821 (N_11821,N_11541,N_11681);
and U11822 (N_11822,N_11437,N_11585);
nand U11823 (N_11823,N_11505,N_11679);
nand U11824 (N_11824,N_11516,N_11508);
xor U11825 (N_11825,N_11690,N_11606);
nor U11826 (N_11826,N_11557,N_11590);
and U11827 (N_11827,N_11540,N_11551);
and U11828 (N_11828,N_11446,N_11594);
nand U11829 (N_11829,N_11548,N_11612);
and U11830 (N_11830,N_11440,N_11643);
nand U11831 (N_11831,N_11603,N_11680);
or U11832 (N_11832,N_11492,N_11547);
and U11833 (N_11833,N_11413,N_11591);
nor U11834 (N_11834,N_11402,N_11614);
or U11835 (N_11835,N_11511,N_11664);
nor U11836 (N_11836,N_11693,N_11528);
xnor U11837 (N_11837,N_11482,N_11634);
nand U11838 (N_11838,N_11450,N_11648);
xor U11839 (N_11839,N_11448,N_11510);
and U11840 (N_11840,N_11605,N_11443);
and U11841 (N_11841,N_11588,N_11652);
xor U11842 (N_11842,N_11423,N_11480);
or U11843 (N_11843,N_11518,N_11669);
nand U11844 (N_11844,N_11404,N_11697);
nor U11845 (N_11845,N_11662,N_11576);
or U11846 (N_11846,N_11601,N_11687);
xor U11847 (N_11847,N_11421,N_11692);
and U11848 (N_11848,N_11699,N_11439);
nor U11849 (N_11849,N_11484,N_11686);
or U11850 (N_11850,N_11535,N_11599);
nand U11851 (N_11851,N_11573,N_11453);
or U11852 (N_11852,N_11414,N_11466);
nor U11853 (N_11853,N_11475,N_11541);
nor U11854 (N_11854,N_11696,N_11426);
nor U11855 (N_11855,N_11581,N_11562);
or U11856 (N_11856,N_11550,N_11611);
or U11857 (N_11857,N_11570,N_11524);
nor U11858 (N_11858,N_11429,N_11508);
or U11859 (N_11859,N_11445,N_11416);
xnor U11860 (N_11860,N_11506,N_11503);
nor U11861 (N_11861,N_11512,N_11696);
and U11862 (N_11862,N_11552,N_11531);
nand U11863 (N_11863,N_11459,N_11522);
nand U11864 (N_11864,N_11410,N_11532);
or U11865 (N_11865,N_11640,N_11566);
xnor U11866 (N_11866,N_11413,N_11507);
and U11867 (N_11867,N_11530,N_11431);
nand U11868 (N_11868,N_11438,N_11427);
xor U11869 (N_11869,N_11611,N_11671);
nor U11870 (N_11870,N_11580,N_11437);
or U11871 (N_11871,N_11533,N_11652);
nor U11872 (N_11872,N_11522,N_11666);
nand U11873 (N_11873,N_11547,N_11697);
nor U11874 (N_11874,N_11429,N_11635);
xnor U11875 (N_11875,N_11687,N_11491);
nand U11876 (N_11876,N_11582,N_11492);
or U11877 (N_11877,N_11535,N_11409);
and U11878 (N_11878,N_11484,N_11521);
xnor U11879 (N_11879,N_11403,N_11671);
and U11880 (N_11880,N_11405,N_11472);
or U11881 (N_11881,N_11439,N_11592);
or U11882 (N_11882,N_11587,N_11518);
or U11883 (N_11883,N_11601,N_11423);
and U11884 (N_11884,N_11493,N_11578);
or U11885 (N_11885,N_11411,N_11502);
or U11886 (N_11886,N_11486,N_11632);
and U11887 (N_11887,N_11649,N_11486);
and U11888 (N_11888,N_11458,N_11622);
nor U11889 (N_11889,N_11435,N_11508);
and U11890 (N_11890,N_11523,N_11570);
nor U11891 (N_11891,N_11552,N_11527);
nand U11892 (N_11892,N_11687,N_11606);
and U11893 (N_11893,N_11425,N_11609);
or U11894 (N_11894,N_11635,N_11669);
and U11895 (N_11895,N_11688,N_11483);
nor U11896 (N_11896,N_11677,N_11560);
nor U11897 (N_11897,N_11527,N_11490);
xor U11898 (N_11898,N_11604,N_11502);
and U11899 (N_11899,N_11653,N_11486);
or U11900 (N_11900,N_11686,N_11489);
and U11901 (N_11901,N_11597,N_11504);
nand U11902 (N_11902,N_11565,N_11464);
nor U11903 (N_11903,N_11481,N_11441);
xnor U11904 (N_11904,N_11527,N_11548);
and U11905 (N_11905,N_11413,N_11679);
and U11906 (N_11906,N_11517,N_11499);
xor U11907 (N_11907,N_11688,N_11671);
or U11908 (N_11908,N_11680,N_11555);
nand U11909 (N_11909,N_11553,N_11406);
nand U11910 (N_11910,N_11633,N_11496);
and U11911 (N_11911,N_11555,N_11449);
xor U11912 (N_11912,N_11423,N_11422);
or U11913 (N_11913,N_11537,N_11661);
or U11914 (N_11914,N_11640,N_11598);
xor U11915 (N_11915,N_11485,N_11436);
xor U11916 (N_11916,N_11442,N_11555);
nand U11917 (N_11917,N_11513,N_11470);
or U11918 (N_11918,N_11552,N_11623);
and U11919 (N_11919,N_11462,N_11619);
nand U11920 (N_11920,N_11509,N_11687);
nor U11921 (N_11921,N_11418,N_11549);
xnor U11922 (N_11922,N_11583,N_11593);
or U11923 (N_11923,N_11542,N_11515);
nand U11924 (N_11924,N_11410,N_11606);
and U11925 (N_11925,N_11466,N_11640);
nor U11926 (N_11926,N_11453,N_11564);
nand U11927 (N_11927,N_11439,N_11627);
or U11928 (N_11928,N_11552,N_11694);
nand U11929 (N_11929,N_11507,N_11402);
and U11930 (N_11930,N_11412,N_11635);
or U11931 (N_11931,N_11468,N_11436);
nor U11932 (N_11932,N_11643,N_11481);
xnor U11933 (N_11933,N_11517,N_11505);
xnor U11934 (N_11934,N_11579,N_11692);
and U11935 (N_11935,N_11697,N_11458);
nor U11936 (N_11936,N_11443,N_11482);
nand U11937 (N_11937,N_11625,N_11564);
and U11938 (N_11938,N_11412,N_11542);
or U11939 (N_11939,N_11402,N_11669);
xor U11940 (N_11940,N_11629,N_11692);
or U11941 (N_11941,N_11526,N_11541);
nor U11942 (N_11942,N_11473,N_11646);
nor U11943 (N_11943,N_11412,N_11551);
or U11944 (N_11944,N_11688,N_11619);
xor U11945 (N_11945,N_11634,N_11408);
or U11946 (N_11946,N_11468,N_11411);
nor U11947 (N_11947,N_11492,N_11479);
and U11948 (N_11948,N_11639,N_11455);
nor U11949 (N_11949,N_11433,N_11541);
and U11950 (N_11950,N_11602,N_11535);
nand U11951 (N_11951,N_11590,N_11410);
nor U11952 (N_11952,N_11492,N_11659);
nand U11953 (N_11953,N_11562,N_11596);
xor U11954 (N_11954,N_11644,N_11478);
nor U11955 (N_11955,N_11422,N_11547);
xnor U11956 (N_11956,N_11424,N_11451);
and U11957 (N_11957,N_11538,N_11666);
or U11958 (N_11958,N_11416,N_11551);
and U11959 (N_11959,N_11408,N_11667);
xor U11960 (N_11960,N_11526,N_11521);
xnor U11961 (N_11961,N_11521,N_11515);
xor U11962 (N_11962,N_11454,N_11464);
xnor U11963 (N_11963,N_11470,N_11640);
nand U11964 (N_11964,N_11424,N_11646);
or U11965 (N_11965,N_11632,N_11634);
nor U11966 (N_11966,N_11566,N_11647);
xor U11967 (N_11967,N_11643,N_11437);
nand U11968 (N_11968,N_11626,N_11469);
xor U11969 (N_11969,N_11444,N_11508);
nor U11970 (N_11970,N_11419,N_11450);
or U11971 (N_11971,N_11468,N_11646);
or U11972 (N_11972,N_11602,N_11668);
or U11973 (N_11973,N_11650,N_11651);
xnor U11974 (N_11974,N_11546,N_11455);
or U11975 (N_11975,N_11563,N_11670);
nand U11976 (N_11976,N_11467,N_11572);
and U11977 (N_11977,N_11605,N_11634);
nor U11978 (N_11978,N_11473,N_11455);
nor U11979 (N_11979,N_11621,N_11594);
and U11980 (N_11980,N_11427,N_11684);
nor U11981 (N_11981,N_11426,N_11544);
xor U11982 (N_11982,N_11602,N_11481);
or U11983 (N_11983,N_11421,N_11461);
and U11984 (N_11984,N_11649,N_11436);
xor U11985 (N_11985,N_11631,N_11569);
or U11986 (N_11986,N_11675,N_11529);
and U11987 (N_11987,N_11578,N_11481);
nor U11988 (N_11988,N_11495,N_11603);
or U11989 (N_11989,N_11628,N_11402);
and U11990 (N_11990,N_11476,N_11515);
and U11991 (N_11991,N_11551,N_11511);
and U11992 (N_11992,N_11667,N_11498);
nor U11993 (N_11993,N_11575,N_11491);
or U11994 (N_11994,N_11649,N_11414);
or U11995 (N_11995,N_11413,N_11538);
and U11996 (N_11996,N_11524,N_11632);
xor U11997 (N_11997,N_11617,N_11511);
nand U11998 (N_11998,N_11551,N_11554);
xnor U11999 (N_11999,N_11562,N_11552);
xnor U12000 (N_12000,N_11806,N_11874);
xnor U12001 (N_12001,N_11845,N_11733);
nand U12002 (N_12002,N_11794,N_11798);
nor U12003 (N_12003,N_11870,N_11704);
nor U12004 (N_12004,N_11833,N_11951);
nor U12005 (N_12005,N_11722,N_11934);
nand U12006 (N_12006,N_11703,N_11955);
nand U12007 (N_12007,N_11712,N_11884);
nand U12008 (N_12008,N_11911,N_11982);
or U12009 (N_12009,N_11910,N_11867);
and U12010 (N_12010,N_11967,N_11724);
and U12011 (N_12011,N_11888,N_11864);
xor U12012 (N_12012,N_11941,N_11811);
nor U12013 (N_12013,N_11930,N_11745);
and U12014 (N_12014,N_11940,N_11986);
and U12015 (N_12015,N_11840,N_11937);
or U12016 (N_12016,N_11772,N_11970);
nand U12017 (N_12017,N_11735,N_11869);
nand U12018 (N_12018,N_11943,N_11990);
or U12019 (N_12019,N_11879,N_11889);
or U12020 (N_12020,N_11968,N_11732);
xnor U12021 (N_12021,N_11752,N_11979);
and U12022 (N_12022,N_11956,N_11717);
or U12023 (N_12023,N_11853,N_11729);
or U12024 (N_12024,N_11725,N_11927);
nand U12025 (N_12025,N_11932,N_11823);
nand U12026 (N_12026,N_11764,N_11834);
or U12027 (N_12027,N_11714,N_11918);
nor U12028 (N_12028,N_11816,N_11768);
and U12029 (N_12029,N_11915,N_11878);
nand U12030 (N_12030,N_11776,N_11829);
or U12031 (N_12031,N_11756,N_11734);
xor U12032 (N_12032,N_11906,N_11887);
nor U12033 (N_12033,N_11966,N_11877);
nand U12034 (N_12034,N_11942,N_11914);
or U12035 (N_12035,N_11825,N_11813);
and U12036 (N_12036,N_11861,N_11959);
nand U12037 (N_12037,N_11720,N_11983);
nand U12038 (N_12038,N_11849,N_11814);
or U12039 (N_12039,N_11962,N_11999);
nor U12040 (N_12040,N_11846,N_11783);
or U12041 (N_12041,N_11706,N_11753);
nand U12042 (N_12042,N_11715,N_11707);
or U12043 (N_12043,N_11730,N_11796);
nor U12044 (N_12044,N_11969,N_11975);
and U12045 (N_12045,N_11716,N_11862);
nand U12046 (N_12046,N_11963,N_11807);
or U12047 (N_12047,N_11763,N_11789);
or U12048 (N_12048,N_11819,N_11981);
or U12049 (N_12049,N_11863,N_11800);
nor U12050 (N_12050,N_11711,N_11933);
and U12051 (N_12051,N_11821,N_11902);
nand U12052 (N_12052,N_11894,N_11786);
or U12053 (N_12053,N_11944,N_11993);
xor U12054 (N_12054,N_11987,N_11767);
nand U12055 (N_12055,N_11801,N_11890);
nand U12056 (N_12056,N_11857,N_11779);
and U12057 (N_12057,N_11892,N_11936);
xnor U12058 (N_12058,N_11810,N_11770);
xnor U12059 (N_12059,N_11868,N_11923);
nand U12060 (N_12060,N_11971,N_11795);
xor U12061 (N_12061,N_11827,N_11835);
nand U12062 (N_12062,N_11950,N_11782);
nand U12063 (N_12063,N_11713,N_11973);
or U12064 (N_12064,N_11916,N_11850);
xnor U12065 (N_12065,N_11978,N_11952);
nor U12066 (N_12066,N_11908,N_11784);
nand U12067 (N_12067,N_11928,N_11872);
xnor U12068 (N_12068,N_11891,N_11896);
or U12069 (N_12069,N_11964,N_11700);
and U12070 (N_12070,N_11792,N_11995);
nor U12071 (N_12071,N_11728,N_11960);
nor U12072 (N_12072,N_11781,N_11997);
and U12073 (N_12073,N_11804,N_11946);
and U12074 (N_12074,N_11721,N_11965);
and U12075 (N_12075,N_11740,N_11812);
nand U12076 (N_12076,N_11830,N_11949);
nand U12077 (N_12077,N_11921,N_11907);
or U12078 (N_12078,N_11843,N_11788);
and U12079 (N_12079,N_11848,N_11817);
nand U12080 (N_12080,N_11984,N_11954);
nand U12081 (N_12081,N_11885,N_11780);
nand U12082 (N_12082,N_11702,N_11755);
xor U12083 (N_12083,N_11925,N_11769);
or U12084 (N_12084,N_11777,N_11851);
xnor U12085 (N_12085,N_11858,N_11760);
nand U12086 (N_12086,N_11919,N_11790);
xnor U12087 (N_12087,N_11931,N_11882);
or U12088 (N_12088,N_11837,N_11988);
or U12089 (N_12089,N_11876,N_11855);
nor U12090 (N_12090,N_11996,N_11977);
nor U12091 (N_12091,N_11739,N_11909);
or U12092 (N_12092,N_11765,N_11992);
or U12093 (N_12093,N_11748,N_11886);
xnor U12094 (N_12094,N_11945,N_11750);
and U12095 (N_12095,N_11778,N_11935);
and U12096 (N_12096,N_11991,N_11948);
nand U12097 (N_12097,N_11917,N_11880);
and U12098 (N_12098,N_11929,N_11974);
nor U12099 (N_12099,N_11920,N_11976);
and U12100 (N_12100,N_11961,N_11746);
xnor U12101 (N_12101,N_11709,N_11953);
nor U12102 (N_12102,N_11803,N_11898);
nor U12103 (N_12103,N_11985,N_11901);
nand U12104 (N_12104,N_11939,N_11805);
nand U12105 (N_12105,N_11913,N_11736);
or U12106 (N_12106,N_11787,N_11852);
nand U12107 (N_12107,N_11831,N_11771);
nor U12108 (N_12108,N_11836,N_11824);
or U12109 (N_12109,N_11773,N_11873);
nand U12110 (N_12110,N_11922,N_11859);
xnor U12111 (N_12111,N_11912,N_11972);
xor U12112 (N_12112,N_11924,N_11856);
and U12113 (N_12113,N_11998,N_11947);
nand U12114 (N_12114,N_11904,N_11899);
and U12115 (N_12115,N_11926,N_11737);
nor U12116 (N_12116,N_11866,N_11708);
and U12117 (N_12117,N_11815,N_11762);
nor U12118 (N_12118,N_11842,N_11741);
nor U12119 (N_12119,N_11895,N_11797);
nand U12120 (N_12120,N_11980,N_11726);
nor U12121 (N_12121,N_11818,N_11839);
xor U12122 (N_12122,N_11723,N_11994);
or U12123 (N_12123,N_11785,N_11742);
nand U12124 (N_12124,N_11758,N_11838);
and U12125 (N_12125,N_11751,N_11791);
and U12126 (N_12126,N_11841,N_11705);
nor U12127 (N_12127,N_11761,N_11766);
and U12128 (N_12128,N_11719,N_11883);
xnor U12129 (N_12129,N_11820,N_11775);
xnor U12130 (N_12130,N_11793,N_11774);
nor U12131 (N_12131,N_11799,N_11865);
or U12132 (N_12132,N_11828,N_11854);
and U12133 (N_12133,N_11826,N_11731);
or U12134 (N_12134,N_11743,N_11871);
and U12135 (N_12135,N_11893,N_11958);
and U12136 (N_12136,N_11802,N_11701);
and U12137 (N_12137,N_11749,N_11903);
or U12138 (N_12138,N_11809,N_11989);
or U12139 (N_12139,N_11718,N_11759);
and U12140 (N_12140,N_11847,N_11822);
or U12141 (N_12141,N_11754,N_11875);
or U12142 (N_12142,N_11727,N_11744);
xnor U12143 (N_12143,N_11881,N_11738);
and U12144 (N_12144,N_11957,N_11710);
xor U12145 (N_12145,N_11905,N_11844);
nor U12146 (N_12146,N_11757,N_11860);
nand U12147 (N_12147,N_11900,N_11832);
xor U12148 (N_12148,N_11747,N_11897);
nor U12149 (N_12149,N_11808,N_11938);
nand U12150 (N_12150,N_11911,N_11882);
xnor U12151 (N_12151,N_11898,N_11985);
nand U12152 (N_12152,N_11714,N_11855);
or U12153 (N_12153,N_11854,N_11735);
or U12154 (N_12154,N_11948,N_11879);
and U12155 (N_12155,N_11868,N_11846);
or U12156 (N_12156,N_11891,N_11919);
xor U12157 (N_12157,N_11875,N_11983);
or U12158 (N_12158,N_11908,N_11911);
xnor U12159 (N_12159,N_11741,N_11775);
nand U12160 (N_12160,N_11735,N_11902);
nand U12161 (N_12161,N_11930,N_11977);
and U12162 (N_12162,N_11759,N_11741);
or U12163 (N_12163,N_11940,N_11737);
xor U12164 (N_12164,N_11825,N_11739);
nand U12165 (N_12165,N_11993,N_11892);
or U12166 (N_12166,N_11871,N_11721);
nor U12167 (N_12167,N_11707,N_11738);
xnor U12168 (N_12168,N_11800,N_11967);
and U12169 (N_12169,N_11773,N_11769);
nand U12170 (N_12170,N_11892,N_11875);
or U12171 (N_12171,N_11997,N_11769);
or U12172 (N_12172,N_11859,N_11925);
nor U12173 (N_12173,N_11953,N_11966);
or U12174 (N_12174,N_11858,N_11847);
nor U12175 (N_12175,N_11743,N_11711);
nor U12176 (N_12176,N_11814,N_11874);
or U12177 (N_12177,N_11997,N_11991);
and U12178 (N_12178,N_11728,N_11733);
and U12179 (N_12179,N_11952,N_11959);
nor U12180 (N_12180,N_11976,N_11882);
or U12181 (N_12181,N_11955,N_11751);
and U12182 (N_12182,N_11853,N_11957);
nor U12183 (N_12183,N_11984,N_11767);
or U12184 (N_12184,N_11902,N_11707);
xnor U12185 (N_12185,N_11700,N_11856);
xor U12186 (N_12186,N_11980,N_11950);
nor U12187 (N_12187,N_11845,N_11883);
or U12188 (N_12188,N_11881,N_11842);
xnor U12189 (N_12189,N_11954,N_11881);
and U12190 (N_12190,N_11791,N_11834);
or U12191 (N_12191,N_11732,N_11874);
nand U12192 (N_12192,N_11997,N_11883);
nor U12193 (N_12193,N_11701,N_11748);
and U12194 (N_12194,N_11989,N_11755);
or U12195 (N_12195,N_11776,N_11738);
nand U12196 (N_12196,N_11864,N_11815);
nand U12197 (N_12197,N_11940,N_11735);
nor U12198 (N_12198,N_11846,N_11780);
or U12199 (N_12199,N_11813,N_11986);
nand U12200 (N_12200,N_11928,N_11946);
xnor U12201 (N_12201,N_11903,N_11939);
nor U12202 (N_12202,N_11753,N_11866);
and U12203 (N_12203,N_11793,N_11749);
nand U12204 (N_12204,N_11755,N_11830);
nor U12205 (N_12205,N_11998,N_11778);
xor U12206 (N_12206,N_11919,N_11783);
xnor U12207 (N_12207,N_11916,N_11706);
nand U12208 (N_12208,N_11882,N_11722);
nor U12209 (N_12209,N_11959,N_11859);
or U12210 (N_12210,N_11806,N_11976);
xor U12211 (N_12211,N_11951,N_11764);
nand U12212 (N_12212,N_11832,N_11938);
nand U12213 (N_12213,N_11835,N_11702);
or U12214 (N_12214,N_11921,N_11953);
or U12215 (N_12215,N_11755,N_11782);
and U12216 (N_12216,N_11758,N_11822);
nor U12217 (N_12217,N_11939,N_11801);
and U12218 (N_12218,N_11703,N_11847);
nor U12219 (N_12219,N_11716,N_11831);
nor U12220 (N_12220,N_11872,N_11871);
nand U12221 (N_12221,N_11746,N_11747);
xor U12222 (N_12222,N_11809,N_11978);
and U12223 (N_12223,N_11727,N_11990);
and U12224 (N_12224,N_11863,N_11864);
and U12225 (N_12225,N_11974,N_11957);
and U12226 (N_12226,N_11850,N_11941);
nand U12227 (N_12227,N_11753,N_11974);
nor U12228 (N_12228,N_11944,N_11852);
or U12229 (N_12229,N_11918,N_11790);
and U12230 (N_12230,N_11933,N_11790);
xnor U12231 (N_12231,N_11770,N_11827);
or U12232 (N_12232,N_11910,N_11727);
and U12233 (N_12233,N_11730,N_11845);
and U12234 (N_12234,N_11889,N_11952);
or U12235 (N_12235,N_11943,N_11817);
and U12236 (N_12236,N_11860,N_11941);
nor U12237 (N_12237,N_11983,N_11786);
nor U12238 (N_12238,N_11972,N_11729);
xor U12239 (N_12239,N_11954,N_11917);
xor U12240 (N_12240,N_11725,N_11960);
xnor U12241 (N_12241,N_11924,N_11978);
or U12242 (N_12242,N_11906,N_11817);
nand U12243 (N_12243,N_11997,N_11737);
or U12244 (N_12244,N_11926,N_11705);
or U12245 (N_12245,N_11756,N_11926);
nor U12246 (N_12246,N_11766,N_11880);
or U12247 (N_12247,N_11873,N_11784);
xnor U12248 (N_12248,N_11703,N_11851);
nand U12249 (N_12249,N_11874,N_11720);
nor U12250 (N_12250,N_11903,N_11928);
nor U12251 (N_12251,N_11955,N_11804);
or U12252 (N_12252,N_11881,N_11959);
nand U12253 (N_12253,N_11719,N_11993);
or U12254 (N_12254,N_11831,N_11968);
and U12255 (N_12255,N_11778,N_11842);
or U12256 (N_12256,N_11993,N_11703);
nor U12257 (N_12257,N_11705,N_11760);
nand U12258 (N_12258,N_11734,N_11702);
nor U12259 (N_12259,N_11740,N_11970);
and U12260 (N_12260,N_11868,N_11998);
nand U12261 (N_12261,N_11879,N_11917);
and U12262 (N_12262,N_11731,N_11799);
nand U12263 (N_12263,N_11869,N_11936);
xnor U12264 (N_12264,N_11895,N_11801);
or U12265 (N_12265,N_11953,N_11991);
nor U12266 (N_12266,N_11858,N_11922);
xnor U12267 (N_12267,N_11802,N_11790);
xor U12268 (N_12268,N_11908,N_11855);
xnor U12269 (N_12269,N_11873,N_11753);
nand U12270 (N_12270,N_11778,N_11803);
xnor U12271 (N_12271,N_11886,N_11995);
xor U12272 (N_12272,N_11774,N_11998);
and U12273 (N_12273,N_11791,N_11936);
xnor U12274 (N_12274,N_11863,N_11848);
xor U12275 (N_12275,N_11787,N_11781);
or U12276 (N_12276,N_11982,N_11816);
or U12277 (N_12277,N_11766,N_11826);
or U12278 (N_12278,N_11959,N_11895);
xnor U12279 (N_12279,N_11882,N_11981);
xnor U12280 (N_12280,N_11991,N_11732);
nand U12281 (N_12281,N_11847,N_11762);
or U12282 (N_12282,N_11801,N_11824);
nor U12283 (N_12283,N_11770,N_11940);
xnor U12284 (N_12284,N_11834,N_11729);
and U12285 (N_12285,N_11801,N_11874);
nand U12286 (N_12286,N_11989,N_11855);
nand U12287 (N_12287,N_11869,N_11946);
or U12288 (N_12288,N_11803,N_11990);
nor U12289 (N_12289,N_11745,N_11828);
nor U12290 (N_12290,N_11823,N_11722);
nor U12291 (N_12291,N_11955,N_11959);
or U12292 (N_12292,N_11931,N_11992);
or U12293 (N_12293,N_11988,N_11982);
and U12294 (N_12294,N_11707,N_11781);
xor U12295 (N_12295,N_11908,N_11734);
nor U12296 (N_12296,N_11925,N_11883);
or U12297 (N_12297,N_11993,N_11764);
xor U12298 (N_12298,N_11827,N_11787);
or U12299 (N_12299,N_11702,N_11771);
nand U12300 (N_12300,N_12011,N_12203);
nand U12301 (N_12301,N_12259,N_12246);
nand U12302 (N_12302,N_12251,N_12238);
xor U12303 (N_12303,N_12041,N_12146);
xnor U12304 (N_12304,N_12192,N_12147);
nand U12305 (N_12305,N_12233,N_12269);
xnor U12306 (N_12306,N_12110,N_12247);
nand U12307 (N_12307,N_12121,N_12194);
xnor U12308 (N_12308,N_12169,N_12168);
and U12309 (N_12309,N_12025,N_12176);
and U12310 (N_12310,N_12236,N_12007);
and U12311 (N_12311,N_12111,N_12250);
and U12312 (N_12312,N_12114,N_12135);
or U12313 (N_12313,N_12137,N_12024);
nor U12314 (N_12314,N_12214,N_12115);
and U12315 (N_12315,N_12198,N_12086);
nor U12316 (N_12316,N_12260,N_12240);
or U12317 (N_12317,N_12243,N_12093);
or U12318 (N_12318,N_12063,N_12266);
or U12319 (N_12319,N_12188,N_12245);
or U12320 (N_12320,N_12167,N_12087);
and U12321 (N_12321,N_12197,N_12189);
and U12322 (N_12322,N_12280,N_12201);
nor U12323 (N_12323,N_12042,N_12183);
xor U12324 (N_12324,N_12285,N_12090);
xor U12325 (N_12325,N_12255,N_12065);
nand U12326 (N_12326,N_12049,N_12289);
or U12327 (N_12327,N_12180,N_12045);
or U12328 (N_12328,N_12297,N_12278);
nand U12329 (N_12329,N_12195,N_12241);
or U12330 (N_12330,N_12089,N_12116);
nor U12331 (N_12331,N_12258,N_12092);
nand U12332 (N_12332,N_12112,N_12252);
or U12333 (N_12333,N_12181,N_12179);
or U12334 (N_12334,N_12030,N_12070);
and U12335 (N_12335,N_12193,N_12222);
nor U12336 (N_12336,N_12129,N_12082);
nor U12337 (N_12337,N_12215,N_12102);
nand U12338 (N_12338,N_12173,N_12164);
and U12339 (N_12339,N_12154,N_12174);
xnor U12340 (N_12340,N_12133,N_12265);
and U12341 (N_12341,N_12091,N_12066);
xor U12342 (N_12342,N_12064,N_12134);
or U12343 (N_12343,N_12295,N_12299);
or U12344 (N_12344,N_12225,N_12150);
or U12345 (N_12345,N_12142,N_12022);
xor U12346 (N_12346,N_12277,N_12079);
or U12347 (N_12347,N_12058,N_12261);
or U12348 (N_12348,N_12177,N_12230);
nand U12349 (N_12349,N_12264,N_12004);
and U12350 (N_12350,N_12076,N_12032);
xor U12351 (N_12351,N_12149,N_12219);
or U12352 (N_12352,N_12283,N_12253);
and U12353 (N_12353,N_12101,N_12132);
nor U12354 (N_12354,N_12175,N_12153);
and U12355 (N_12355,N_12160,N_12124);
and U12356 (N_12356,N_12248,N_12071);
nor U12357 (N_12357,N_12166,N_12224);
xnor U12358 (N_12358,N_12060,N_12182);
or U12359 (N_12359,N_12163,N_12006);
and U12360 (N_12360,N_12199,N_12159);
nor U12361 (N_12361,N_12069,N_12044);
or U12362 (N_12362,N_12139,N_12262);
and U12363 (N_12363,N_12141,N_12190);
nor U12364 (N_12364,N_12023,N_12205);
and U12365 (N_12365,N_12213,N_12012);
or U12366 (N_12366,N_12254,N_12292);
nor U12367 (N_12367,N_12220,N_12273);
nand U12368 (N_12368,N_12085,N_12062);
and U12369 (N_12369,N_12125,N_12216);
xor U12370 (N_12370,N_12123,N_12016);
xnor U12371 (N_12371,N_12281,N_12155);
nor U12372 (N_12372,N_12196,N_12267);
nand U12373 (N_12373,N_12015,N_12017);
and U12374 (N_12374,N_12104,N_12008);
nor U12375 (N_12375,N_12027,N_12156);
xnor U12376 (N_12376,N_12095,N_12035);
nor U12377 (N_12377,N_12221,N_12239);
and U12378 (N_12378,N_12152,N_12072);
nor U12379 (N_12379,N_12140,N_12067);
or U12380 (N_12380,N_12271,N_12131);
and U12381 (N_12381,N_12158,N_12223);
or U12382 (N_12382,N_12053,N_12191);
and U12383 (N_12383,N_12094,N_12081);
nand U12384 (N_12384,N_12038,N_12013);
or U12385 (N_12385,N_12286,N_12028);
or U12386 (N_12386,N_12206,N_12046);
nor U12387 (N_12387,N_12040,N_12178);
xnor U12388 (N_12388,N_12108,N_12130);
and U12389 (N_12389,N_12296,N_12204);
and U12390 (N_12390,N_12228,N_12096);
or U12391 (N_12391,N_12172,N_12157);
or U12392 (N_12392,N_12298,N_12145);
xnor U12393 (N_12393,N_12294,N_12293);
xor U12394 (N_12394,N_12232,N_12034);
xnor U12395 (N_12395,N_12021,N_12014);
and U12396 (N_12396,N_12217,N_12211);
xor U12397 (N_12397,N_12084,N_12026);
and U12398 (N_12398,N_12287,N_12005);
and U12399 (N_12399,N_12249,N_12276);
nand U12400 (N_12400,N_12052,N_12078);
or U12401 (N_12401,N_12165,N_12151);
nand U12402 (N_12402,N_12161,N_12107);
nor U12403 (N_12403,N_12185,N_12054);
nor U12404 (N_12404,N_12029,N_12018);
xnor U12405 (N_12405,N_12119,N_12227);
and U12406 (N_12406,N_12234,N_12077);
nand U12407 (N_12407,N_12138,N_12083);
and U12408 (N_12408,N_12207,N_12088);
xnor U12409 (N_12409,N_12272,N_12120);
or U12410 (N_12410,N_12170,N_12097);
and U12411 (N_12411,N_12162,N_12109);
nor U12412 (N_12412,N_12268,N_12279);
nor U12413 (N_12413,N_12117,N_12019);
nor U12414 (N_12414,N_12055,N_12020);
nor U12415 (N_12415,N_12113,N_12010);
xor U12416 (N_12416,N_12242,N_12290);
and U12417 (N_12417,N_12231,N_12031);
and U12418 (N_12418,N_12033,N_12002);
and U12419 (N_12419,N_12103,N_12057);
nor U12420 (N_12420,N_12051,N_12200);
nor U12421 (N_12421,N_12226,N_12237);
or U12422 (N_12422,N_12043,N_12074);
xnor U12423 (N_12423,N_12284,N_12073);
xnor U12424 (N_12424,N_12263,N_12039);
or U12425 (N_12425,N_12171,N_12037);
xor U12426 (N_12426,N_12118,N_12036);
nand U12427 (N_12427,N_12291,N_12127);
xnor U12428 (N_12428,N_12229,N_12122);
or U12429 (N_12429,N_12244,N_12056);
xnor U12430 (N_12430,N_12080,N_12288);
nor U12431 (N_12431,N_12218,N_12099);
and U12432 (N_12432,N_12048,N_12128);
nor U12433 (N_12433,N_12148,N_12009);
or U12434 (N_12434,N_12098,N_12075);
xnor U12435 (N_12435,N_12256,N_12105);
nand U12436 (N_12436,N_12059,N_12100);
nor U12437 (N_12437,N_12136,N_12126);
and U12438 (N_12438,N_12209,N_12210);
nand U12439 (N_12439,N_12144,N_12047);
nand U12440 (N_12440,N_12202,N_12061);
and U12441 (N_12441,N_12212,N_12143);
or U12442 (N_12442,N_12235,N_12001);
nand U12443 (N_12443,N_12208,N_12106);
and U12444 (N_12444,N_12187,N_12186);
or U12445 (N_12445,N_12257,N_12068);
nand U12446 (N_12446,N_12282,N_12050);
nor U12447 (N_12447,N_12275,N_12270);
or U12448 (N_12448,N_12000,N_12184);
nand U12449 (N_12449,N_12003,N_12274);
and U12450 (N_12450,N_12288,N_12026);
xnor U12451 (N_12451,N_12291,N_12040);
and U12452 (N_12452,N_12140,N_12061);
nor U12453 (N_12453,N_12016,N_12178);
nor U12454 (N_12454,N_12062,N_12049);
xnor U12455 (N_12455,N_12236,N_12199);
and U12456 (N_12456,N_12053,N_12075);
or U12457 (N_12457,N_12022,N_12273);
xor U12458 (N_12458,N_12236,N_12256);
nand U12459 (N_12459,N_12150,N_12194);
nor U12460 (N_12460,N_12188,N_12239);
nor U12461 (N_12461,N_12042,N_12099);
xnor U12462 (N_12462,N_12043,N_12003);
xor U12463 (N_12463,N_12103,N_12241);
or U12464 (N_12464,N_12136,N_12272);
nand U12465 (N_12465,N_12253,N_12014);
xnor U12466 (N_12466,N_12042,N_12178);
nand U12467 (N_12467,N_12094,N_12133);
nor U12468 (N_12468,N_12150,N_12246);
nand U12469 (N_12469,N_12297,N_12288);
and U12470 (N_12470,N_12260,N_12081);
nor U12471 (N_12471,N_12039,N_12282);
xnor U12472 (N_12472,N_12106,N_12174);
nor U12473 (N_12473,N_12200,N_12081);
nand U12474 (N_12474,N_12178,N_12235);
xor U12475 (N_12475,N_12145,N_12129);
xnor U12476 (N_12476,N_12222,N_12050);
nand U12477 (N_12477,N_12212,N_12208);
nand U12478 (N_12478,N_12222,N_12254);
nand U12479 (N_12479,N_12273,N_12042);
nor U12480 (N_12480,N_12132,N_12259);
or U12481 (N_12481,N_12163,N_12046);
or U12482 (N_12482,N_12196,N_12282);
nand U12483 (N_12483,N_12027,N_12275);
nor U12484 (N_12484,N_12210,N_12046);
or U12485 (N_12485,N_12023,N_12115);
and U12486 (N_12486,N_12121,N_12044);
nor U12487 (N_12487,N_12019,N_12150);
and U12488 (N_12488,N_12236,N_12123);
nor U12489 (N_12489,N_12113,N_12283);
or U12490 (N_12490,N_12202,N_12257);
xnor U12491 (N_12491,N_12157,N_12257);
and U12492 (N_12492,N_12009,N_12192);
xor U12493 (N_12493,N_12214,N_12158);
xor U12494 (N_12494,N_12217,N_12271);
and U12495 (N_12495,N_12232,N_12089);
xnor U12496 (N_12496,N_12209,N_12026);
nand U12497 (N_12497,N_12048,N_12293);
nor U12498 (N_12498,N_12022,N_12054);
nand U12499 (N_12499,N_12063,N_12205);
nor U12500 (N_12500,N_12288,N_12293);
xnor U12501 (N_12501,N_12262,N_12031);
or U12502 (N_12502,N_12098,N_12274);
nand U12503 (N_12503,N_12053,N_12106);
or U12504 (N_12504,N_12265,N_12063);
or U12505 (N_12505,N_12201,N_12030);
nor U12506 (N_12506,N_12109,N_12241);
and U12507 (N_12507,N_12033,N_12023);
nand U12508 (N_12508,N_12041,N_12064);
or U12509 (N_12509,N_12118,N_12229);
or U12510 (N_12510,N_12282,N_12120);
and U12511 (N_12511,N_12016,N_12145);
nor U12512 (N_12512,N_12234,N_12079);
nand U12513 (N_12513,N_12054,N_12221);
xnor U12514 (N_12514,N_12249,N_12296);
nor U12515 (N_12515,N_12139,N_12170);
nor U12516 (N_12516,N_12141,N_12087);
xor U12517 (N_12517,N_12113,N_12257);
nor U12518 (N_12518,N_12041,N_12141);
nand U12519 (N_12519,N_12035,N_12131);
or U12520 (N_12520,N_12138,N_12284);
nand U12521 (N_12521,N_12213,N_12098);
and U12522 (N_12522,N_12109,N_12243);
xor U12523 (N_12523,N_12031,N_12205);
nand U12524 (N_12524,N_12156,N_12287);
or U12525 (N_12525,N_12161,N_12207);
nor U12526 (N_12526,N_12181,N_12037);
or U12527 (N_12527,N_12033,N_12295);
or U12528 (N_12528,N_12239,N_12148);
nand U12529 (N_12529,N_12191,N_12170);
nand U12530 (N_12530,N_12088,N_12199);
and U12531 (N_12531,N_12208,N_12080);
nor U12532 (N_12532,N_12261,N_12089);
nand U12533 (N_12533,N_12156,N_12159);
nor U12534 (N_12534,N_12161,N_12022);
and U12535 (N_12535,N_12162,N_12106);
nor U12536 (N_12536,N_12137,N_12104);
and U12537 (N_12537,N_12124,N_12241);
nor U12538 (N_12538,N_12009,N_12120);
xor U12539 (N_12539,N_12134,N_12054);
or U12540 (N_12540,N_12185,N_12260);
and U12541 (N_12541,N_12024,N_12004);
nor U12542 (N_12542,N_12024,N_12278);
and U12543 (N_12543,N_12225,N_12297);
and U12544 (N_12544,N_12273,N_12259);
xor U12545 (N_12545,N_12288,N_12198);
or U12546 (N_12546,N_12290,N_12231);
or U12547 (N_12547,N_12192,N_12141);
and U12548 (N_12548,N_12037,N_12198);
xor U12549 (N_12549,N_12080,N_12176);
nor U12550 (N_12550,N_12240,N_12011);
nand U12551 (N_12551,N_12135,N_12145);
and U12552 (N_12552,N_12195,N_12001);
xnor U12553 (N_12553,N_12073,N_12185);
nand U12554 (N_12554,N_12048,N_12256);
nor U12555 (N_12555,N_12258,N_12131);
xor U12556 (N_12556,N_12139,N_12127);
and U12557 (N_12557,N_12287,N_12033);
or U12558 (N_12558,N_12164,N_12203);
or U12559 (N_12559,N_12068,N_12275);
or U12560 (N_12560,N_12114,N_12264);
xnor U12561 (N_12561,N_12277,N_12072);
and U12562 (N_12562,N_12133,N_12042);
and U12563 (N_12563,N_12282,N_12030);
xnor U12564 (N_12564,N_12073,N_12255);
nand U12565 (N_12565,N_12019,N_12114);
nor U12566 (N_12566,N_12024,N_12254);
nand U12567 (N_12567,N_12138,N_12085);
nand U12568 (N_12568,N_12246,N_12235);
xnor U12569 (N_12569,N_12067,N_12041);
and U12570 (N_12570,N_12065,N_12099);
nand U12571 (N_12571,N_12033,N_12227);
or U12572 (N_12572,N_12236,N_12089);
or U12573 (N_12573,N_12103,N_12094);
and U12574 (N_12574,N_12009,N_12179);
nand U12575 (N_12575,N_12217,N_12016);
xnor U12576 (N_12576,N_12126,N_12175);
or U12577 (N_12577,N_12181,N_12290);
nor U12578 (N_12578,N_12108,N_12250);
nor U12579 (N_12579,N_12150,N_12026);
nand U12580 (N_12580,N_12254,N_12205);
nand U12581 (N_12581,N_12233,N_12169);
nand U12582 (N_12582,N_12169,N_12115);
nor U12583 (N_12583,N_12030,N_12195);
nand U12584 (N_12584,N_12163,N_12112);
xnor U12585 (N_12585,N_12076,N_12026);
nand U12586 (N_12586,N_12211,N_12166);
and U12587 (N_12587,N_12238,N_12148);
nand U12588 (N_12588,N_12104,N_12080);
nand U12589 (N_12589,N_12041,N_12209);
xor U12590 (N_12590,N_12219,N_12088);
xor U12591 (N_12591,N_12254,N_12080);
nand U12592 (N_12592,N_12007,N_12235);
or U12593 (N_12593,N_12006,N_12015);
and U12594 (N_12594,N_12003,N_12170);
xor U12595 (N_12595,N_12184,N_12177);
and U12596 (N_12596,N_12039,N_12162);
and U12597 (N_12597,N_12191,N_12213);
nand U12598 (N_12598,N_12101,N_12153);
and U12599 (N_12599,N_12282,N_12299);
nand U12600 (N_12600,N_12446,N_12427);
and U12601 (N_12601,N_12323,N_12346);
or U12602 (N_12602,N_12553,N_12362);
and U12603 (N_12603,N_12337,N_12322);
nand U12604 (N_12604,N_12375,N_12502);
or U12605 (N_12605,N_12458,N_12503);
and U12606 (N_12606,N_12352,N_12542);
and U12607 (N_12607,N_12565,N_12329);
nor U12608 (N_12608,N_12302,N_12435);
and U12609 (N_12609,N_12440,N_12593);
or U12610 (N_12610,N_12585,N_12580);
or U12611 (N_12611,N_12527,N_12442);
nor U12612 (N_12612,N_12336,N_12415);
and U12613 (N_12613,N_12573,N_12439);
or U12614 (N_12614,N_12391,N_12596);
nand U12615 (N_12615,N_12549,N_12398);
or U12616 (N_12616,N_12547,N_12574);
nor U12617 (N_12617,N_12570,N_12463);
xnor U12618 (N_12618,N_12557,N_12489);
or U12619 (N_12619,N_12353,N_12450);
and U12620 (N_12620,N_12347,N_12470);
nor U12621 (N_12621,N_12444,N_12515);
or U12622 (N_12622,N_12524,N_12312);
nor U12623 (N_12623,N_12348,N_12507);
and U12624 (N_12624,N_12571,N_12340);
xnor U12625 (N_12625,N_12445,N_12392);
nand U12626 (N_12626,N_12330,N_12568);
and U12627 (N_12627,N_12599,N_12388);
nor U12628 (N_12628,N_12321,N_12447);
nand U12629 (N_12629,N_12484,N_12555);
or U12630 (N_12630,N_12384,N_12394);
nand U12631 (N_12631,N_12335,N_12460);
nand U12632 (N_12632,N_12522,N_12532);
nor U12633 (N_12633,N_12588,N_12455);
nand U12634 (N_12634,N_12584,N_12491);
nor U12635 (N_12635,N_12472,N_12512);
xor U12636 (N_12636,N_12310,N_12399);
nor U12637 (N_12637,N_12357,N_12495);
xor U12638 (N_12638,N_12591,N_12426);
nand U12639 (N_12639,N_12509,N_12514);
nor U12640 (N_12640,N_12339,N_12309);
nand U12641 (N_12641,N_12490,N_12566);
nor U12642 (N_12642,N_12389,N_12479);
nor U12643 (N_12643,N_12378,N_12342);
or U12644 (N_12644,N_12420,N_12303);
and U12645 (N_12645,N_12405,N_12341);
nand U12646 (N_12646,N_12385,N_12561);
xor U12647 (N_12647,N_12480,N_12437);
and U12648 (N_12648,N_12314,N_12453);
xnor U12649 (N_12649,N_12459,N_12334);
and U12650 (N_12650,N_12523,N_12595);
or U12651 (N_12651,N_12386,N_12350);
or U12652 (N_12652,N_12505,N_12421);
nor U12653 (N_12653,N_12543,N_12559);
nand U12654 (N_12654,N_12587,N_12477);
xor U12655 (N_12655,N_12454,N_12541);
nand U12656 (N_12656,N_12544,N_12349);
nor U12657 (N_12657,N_12583,N_12423);
and U12658 (N_12658,N_12493,N_12556);
and U12659 (N_12659,N_12418,N_12368);
nand U12660 (N_12660,N_12538,N_12483);
xnor U12661 (N_12661,N_12438,N_12464);
or U12662 (N_12662,N_12448,N_12598);
nor U12663 (N_12663,N_12590,N_12400);
xor U12664 (N_12664,N_12513,N_12521);
and U12665 (N_12665,N_12533,N_12371);
xnor U12666 (N_12666,N_12520,N_12494);
or U12667 (N_12667,N_12501,N_12551);
and U12668 (N_12668,N_12525,N_12387);
nor U12669 (N_12669,N_12572,N_12361);
nand U12670 (N_12670,N_12372,N_12311);
nor U12671 (N_12671,N_12554,N_12403);
and U12672 (N_12672,N_12518,N_12481);
and U12673 (N_12673,N_12488,N_12428);
or U12674 (N_12674,N_12408,N_12578);
xor U12675 (N_12675,N_12457,N_12496);
or U12676 (N_12676,N_12531,N_12563);
or U12677 (N_12677,N_12345,N_12316);
nand U12678 (N_12678,N_12377,N_12540);
nor U12679 (N_12679,N_12318,N_12517);
xnor U12680 (N_12680,N_12526,N_12456);
nand U12681 (N_12681,N_12468,N_12376);
nor U12682 (N_12682,N_12308,N_12550);
xnor U12683 (N_12683,N_12324,N_12304);
nor U12684 (N_12684,N_12510,N_12382);
nand U12685 (N_12685,N_12485,N_12402);
or U12686 (N_12686,N_12497,N_12597);
nor U12687 (N_12687,N_12373,N_12325);
nor U12688 (N_12688,N_12451,N_12344);
nor U12689 (N_12689,N_12492,N_12473);
nor U12690 (N_12690,N_12576,N_12409);
and U12691 (N_12691,N_12461,N_12511);
nand U12692 (N_12692,N_12545,N_12343);
and U12693 (N_12693,N_12410,N_12366);
xnor U12694 (N_12694,N_12412,N_12516);
xor U12695 (N_12695,N_12552,N_12370);
or U12696 (N_12696,N_12414,N_12536);
nand U12697 (N_12697,N_12327,N_12575);
xor U12698 (N_12698,N_12356,N_12567);
and U12699 (N_12699,N_12395,N_12535);
nand U12700 (N_12700,N_12582,N_12379);
or U12701 (N_12701,N_12300,N_12354);
nor U12702 (N_12702,N_12360,N_12534);
or U12703 (N_12703,N_12449,N_12365);
nand U12704 (N_12704,N_12326,N_12333);
and U12705 (N_12705,N_12407,N_12305);
nor U12706 (N_12706,N_12380,N_12562);
xnor U12707 (N_12707,N_12430,N_12564);
xor U12708 (N_12708,N_12539,N_12560);
nand U12709 (N_12709,N_12363,N_12528);
nand U12710 (N_12710,N_12441,N_12471);
or U12711 (N_12711,N_12529,N_12338);
nand U12712 (N_12712,N_12317,N_12579);
or U12713 (N_12713,N_12504,N_12537);
nor U12714 (N_12714,N_12315,N_12328);
nor U12715 (N_12715,N_12594,N_12436);
nand U12716 (N_12716,N_12301,N_12397);
or U12717 (N_12717,N_12433,N_12381);
or U12718 (N_12718,N_12467,N_12508);
xor U12719 (N_12719,N_12469,N_12307);
or U12720 (N_12720,N_12569,N_12351);
xnor U12721 (N_12721,N_12359,N_12364);
nor U12722 (N_12722,N_12424,N_12519);
xor U12723 (N_12723,N_12411,N_12500);
and U12724 (N_12724,N_12462,N_12369);
xor U12725 (N_12725,N_12474,N_12499);
nor U12726 (N_12726,N_12367,N_12452);
xnor U12727 (N_12727,N_12487,N_12425);
nand U12728 (N_12728,N_12406,N_12417);
and U12729 (N_12729,N_12443,N_12404);
and U12730 (N_12730,N_12313,N_12431);
nand U12731 (N_12731,N_12306,N_12413);
xor U12732 (N_12732,N_12498,N_12383);
or U12733 (N_12733,N_12592,N_12355);
nor U12734 (N_12734,N_12478,N_12581);
nand U12735 (N_12735,N_12419,N_12358);
nor U12736 (N_12736,N_12396,N_12530);
or U12737 (N_12737,N_12374,N_12475);
nand U12738 (N_12738,N_12401,N_12466);
nand U12739 (N_12739,N_12434,N_12422);
nand U12740 (N_12740,N_12319,N_12558);
nor U12741 (N_12741,N_12577,N_12482);
xnor U12742 (N_12742,N_12589,N_12390);
xor U12743 (N_12743,N_12332,N_12465);
or U12744 (N_12744,N_12586,N_12548);
nand U12745 (N_12745,N_12393,N_12429);
xnor U12746 (N_12746,N_12331,N_12320);
and U12747 (N_12747,N_12506,N_12432);
and U12748 (N_12748,N_12486,N_12416);
nand U12749 (N_12749,N_12546,N_12476);
nand U12750 (N_12750,N_12537,N_12511);
nor U12751 (N_12751,N_12442,N_12479);
xnor U12752 (N_12752,N_12423,N_12573);
and U12753 (N_12753,N_12518,N_12339);
and U12754 (N_12754,N_12458,N_12393);
xnor U12755 (N_12755,N_12496,N_12402);
nand U12756 (N_12756,N_12319,N_12564);
or U12757 (N_12757,N_12304,N_12342);
nor U12758 (N_12758,N_12370,N_12470);
nand U12759 (N_12759,N_12367,N_12521);
nand U12760 (N_12760,N_12576,N_12544);
or U12761 (N_12761,N_12441,N_12575);
xor U12762 (N_12762,N_12393,N_12462);
xnor U12763 (N_12763,N_12366,N_12587);
xnor U12764 (N_12764,N_12339,N_12456);
nand U12765 (N_12765,N_12515,N_12388);
and U12766 (N_12766,N_12490,N_12436);
and U12767 (N_12767,N_12592,N_12366);
xnor U12768 (N_12768,N_12500,N_12374);
xnor U12769 (N_12769,N_12530,N_12576);
or U12770 (N_12770,N_12596,N_12496);
nand U12771 (N_12771,N_12475,N_12571);
nor U12772 (N_12772,N_12572,N_12501);
xor U12773 (N_12773,N_12365,N_12445);
xnor U12774 (N_12774,N_12305,N_12319);
nand U12775 (N_12775,N_12421,N_12368);
and U12776 (N_12776,N_12592,N_12446);
or U12777 (N_12777,N_12469,N_12419);
xnor U12778 (N_12778,N_12364,N_12569);
xnor U12779 (N_12779,N_12334,N_12305);
nand U12780 (N_12780,N_12378,N_12395);
and U12781 (N_12781,N_12468,N_12529);
or U12782 (N_12782,N_12309,N_12402);
and U12783 (N_12783,N_12381,N_12559);
xor U12784 (N_12784,N_12494,N_12598);
or U12785 (N_12785,N_12436,N_12338);
xnor U12786 (N_12786,N_12301,N_12380);
nor U12787 (N_12787,N_12568,N_12408);
or U12788 (N_12788,N_12322,N_12547);
nor U12789 (N_12789,N_12479,N_12473);
and U12790 (N_12790,N_12467,N_12558);
xnor U12791 (N_12791,N_12477,N_12316);
nand U12792 (N_12792,N_12386,N_12468);
and U12793 (N_12793,N_12587,N_12344);
or U12794 (N_12794,N_12545,N_12468);
xnor U12795 (N_12795,N_12389,N_12456);
xnor U12796 (N_12796,N_12549,N_12546);
or U12797 (N_12797,N_12506,N_12515);
nor U12798 (N_12798,N_12449,N_12523);
xnor U12799 (N_12799,N_12458,N_12469);
or U12800 (N_12800,N_12501,N_12590);
xor U12801 (N_12801,N_12463,N_12512);
nand U12802 (N_12802,N_12399,N_12598);
nor U12803 (N_12803,N_12559,N_12480);
or U12804 (N_12804,N_12430,N_12362);
nor U12805 (N_12805,N_12591,N_12395);
nor U12806 (N_12806,N_12525,N_12329);
and U12807 (N_12807,N_12490,N_12397);
nor U12808 (N_12808,N_12398,N_12441);
xor U12809 (N_12809,N_12438,N_12485);
and U12810 (N_12810,N_12402,N_12599);
nand U12811 (N_12811,N_12393,N_12428);
or U12812 (N_12812,N_12420,N_12424);
and U12813 (N_12813,N_12413,N_12488);
xnor U12814 (N_12814,N_12374,N_12381);
nor U12815 (N_12815,N_12357,N_12349);
or U12816 (N_12816,N_12460,N_12530);
or U12817 (N_12817,N_12547,N_12385);
xor U12818 (N_12818,N_12565,N_12534);
nor U12819 (N_12819,N_12557,N_12597);
nand U12820 (N_12820,N_12465,N_12533);
xor U12821 (N_12821,N_12396,N_12550);
nor U12822 (N_12822,N_12581,N_12369);
nor U12823 (N_12823,N_12498,N_12524);
and U12824 (N_12824,N_12445,N_12339);
or U12825 (N_12825,N_12314,N_12564);
nand U12826 (N_12826,N_12553,N_12547);
xor U12827 (N_12827,N_12324,N_12477);
xnor U12828 (N_12828,N_12463,N_12388);
nor U12829 (N_12829,N_12345,N_12364);
xnor U12830 (N_12830,N_12538,N_12597);
or U12831 (N_12831,N_12424,N_12372);
or U12832 (N_12832,N_12435,N_12525);
nor U12833 (N_12833,N_12396,N_12470);
and U12834 (N_12834,N_12351,N_12318);
nand U12835 (N_12835,N_12302,N_12339);
or U12836 (N_12836,N_12387,N_12556);
nand U12837 (N_12837,N_12333,N_12374);
nor U12838 (N_12838,N_12326,N_12597);
xor U12839 (N_12839,N_12456,N_12383);
and U12840 (N_12840,N_12445,N_12594);
nand U12841 (N_12841,N_12361,N_12409);
or U12842 (N_12842,N_12438,N_12421);
or U12843 (N_12843,N_12389,N_12399);
nand U12844 (N_12844,N_12338,N_12592);
nor U12845 (N_12845,N_12587,N_12345);
xnor U12846 (N_12846,N_12496,N_12394);
or U12847 (N_12847,N_12433,N_12448);
nor U12848 (N_12848,N_12408,N_12302);
nand U12849 (N_12849,N_12388,N_12500);
xor U12850 (N_12850,N_12405,N_12419);
nand U12851 (N_12851,N_12430,N_12312);
or U12852 (N_12852,N_12330,N_12540);
or U12853 (N_12853,N_12560,N_12304);
and U12854 (N_12854,N_12573,N_12458);
or U12855 (N_12855,N_12425,N_12343);
nor U12856 (N_12856,N_12345,N_12520);
and U12857 (N_12857,N_12341,N_12541);
or U12858 (N_12858,N_12454,N_12428);
nor U12859 (N_12859,N_12549,N_12344);
nand U12860 (N_12860,N_12427,N_12345);
or U12861 (N_12861,N_12558,N_12476);
xnor U12862 (N_12862,N_12569,N_12554);
and U12863 (N_12863,N_12580,N_12486);
nand U12864 (N_12864,N_12361,N_12342);
or U12865 (N_12865,N_12448,N_12309);
xor U12866 (N_12866,N_12333,N_12477);
or U12867 (N_12867,N_12526,N_12451);
xor U12868 (N_12868,N_12449,N_12390);
nor U12869 (N_12869,N_12345,N_12596);
and U12870 (N_12870,N_12307,N_12313);
nand U12871 (N_12871,N_12415,N_12340);
or U12872 (N_12872,N_12543,N_12546);
or U12873 (N_12873,N_12377,N_12457);
or U12874 (N_12874,N_12515,N_12363);
xor U12875 (N_12875,N_12584,N_12442);
nor U12876 (N_12876,N_12338,N_12476);
or U12877 (N_12877,N_12419,N_12519);
nand U12878 (N_12878,N_12434,N_12409);
nand U12879 (N_12879,N_12374,N_12519);
xor U12880 (N_12880,N_12346,N_12381);
and U12881 (N_12881,N_12301,N_12483);
nand U12882 (N_12882,N_12503,N_12455);
nand U12883 (N_12883,N_12483,N_12532);
and U12884 (N_12884,N_12334,N_12469);
xnor U12885 (N_12885,N_12372,N_12552);
nand U12886 (N_12886,N_12371,N_12577);
or U12887 (N_12887,N_12365,N_12492);
and U12888 (N_12888,N_12388,N_12365);
nand U12889 (N_12889,N_12330,N_12326);
or U12890 (N_12890,N_12547,N_12423);
nand U12891 (N_12891,N_12462,N_12366);
nand U12892 (N_12892,N_12411,N_12359);
or U12893 (N_12893,N_12437,N_12498);
nand U12894 (N_12894,N_12485,N_12350);
and U12895 (N_12895,N_12593,N_12365);
nor U12896 (N_12896,N_12391,N_12520);
nor U12897 (N_12897,N_12417,N_12440);
or U12898 (N_12898,N_12408,N_12567);
nand U12899 (N_12899,N_12411,N_12429);
or U12900 (N_12900,N_12771,N_12860);
nand U12901 (N_12901,N_12739,N_12743);
nand U12902 (N_12902,N_12656,N_12622);
xor U12903 (N_12903,N_12630,N_12772);
xor U12904 (N_12904,N_12751,N_12632);
or U12905 (N_12905,N_12741,N_12847);
or U12906 (N_12906,N_12608,N_12726);
and U12907 (N_12907,N_12817,N_12840);
or U12908 (N_12908,N_12681,N_12648);
nand U12909 (N_12909,N_12807,N_12742);
nor U12910 (N_12910,N_12798,N_12809);
nand U12911 (N_12911,N_12799,N_12725);
nor U12912 (N_12912,N_12891,N_12781);
or U12913 (N_12913,N_12796,N_12615);
xor U12914 (N_12914,N_12680,N_12861);
nand U12915 (N_12915,N_12665,N_12869);
nor U12916 (N_12916,N_12894,N_12709);
xor U12917 (N_12917,N_12858,N_12835);
and U12918 (N_12918,N_12713,N_12821);
nor U12919 (N_12919,N_12694,N_12673);
nand U12920 (N_12920,N_12760,N_12856);
or U12921 (N_12921,N_12857,N_12810);
xor U12922 (N_12922,N_12634,N_12754);
xnor U12923 (N_12923,N_12750,N_12778);
and U12924 (N_12924,N_12877,N_12682);
or U12925 (N_12925,N_12818,N_12733);
xnor U12926 (N_12926,N_12710,N_12649);
nor U12927 (N_12927,N_12624,N_12606);
nand U12928 (N_12928,N_12604,N_12723);
or U12929 (N_12929,N_12613,N_12612);
nor U12930 (N_12930,N_12720,N_12805);
nand U12931 (N_12931,N_12832,N_12792);
nand U12932 (N_12932,N_12631,N_12688);
nand U12933 (N_12933,N_12859,N_12602);
xnor U12934 (N_12934,N_12672,N_12868);
xnor U12935 (N_12935,N_12645,N_12700);
or U12936 (N_12936,N_12647,N_12621);
and U12937 (N_12937,N_12697,N_12892);
or U12938 (N_12938,N_12875,N_12716);
and U12939 (N_12939,N_12603,N_12834);
or U12940 (N_12940,N_12676,N_12782);
nor U12941 (N_12941,N_12813,N_12837);
or U12942 (N_12942,N_12728,N_12619);
nor U12943 (N_12943,N_12666,N_12887);
or U12944 (N_12944,N_12628,N_12825);
xnor U12945 (N_12945,N_12671,N_12789);
and U12946 (N_12946,N_12836,N_12611);
and U12947 (N_12947,N_12661,N_12849);
and U12948 (N_12948,N_12788,N_12879);
or U12949 (N_12949,N_12629,N_12839);
xnor U12950 (N_12950,N_12740,N_12765);
and U12951 (N_12951,N_12679,N_12862);
xor U12952 (N_12952,N_12668,N_12812);
and U12953 (N_12953,N_12800,N_12761);
nand U12954 (N_12954,N_12643,N_12841);
xor U12955 (N_12955,N_12642,N_12797);
nor U12956 (N_12956,N_12639,N_12724);
xor U12957 (N_12957,N_12747,N_12829);
xnor U12958 (N_12958,N_12823,N_12816);
or U12959 (N_12959,N_12690,N_12752);
or U12960 (N_12960,N_12824,N_12678);
or U12961 (N_12961,N_12732,N_12734);
and U12962 (N_12962,N_12691,N_12769);
xnor U12963 (N_12963,N_12784,N_12696);
or U12964 (N_12964,N_12746,N_12828);
or U12965 (N_12965,N_12625,N_12702);
and U12966 (N_12966,N_12623,N_12731);
nor U12967 (N_12967,N_12863,N_12779);
and U12968 (N_12968,N_12852,N_12706);
nand U12969 (N_12969,N_12795,N_12756);
and U12970 (N_12970,N_12773,N_12766);
xnor U12971 (N_12971,N_12614,N_12684);
nand U12972 (N_12972,N_12701,N_12777);
or U12973 (N_12973,N_12801,N_12659);
xor U12974 (N_12974,N_12827,N_12893);
and U12975 (N_12975,N_12895,N_12844);
or U12976 (N_12976,N_12610,N_12637);
nor U12977 (N_12977,N_12870,N_12708);
or U12978 (N_12978,N_12670,N_12833);
nor U12979 (N_12979,N_12685,N_12808);
nor U12980 (N_12980,N_12652,N_12881);
nor U12981 (N_12981,N_12683,N_12729);
nand U12982 (N_12982,N_12896,N_12794);
nor U12983 (N_12983,N_12699,N_12646);
xor U12984 (N_12984,N_12884,N_12770);
and U12985 (N_12985,N_12826,N_12635);
nand U12986 (N_12986,N_12638,N_12871);
or U12987 (N_12987,N_12758,N_12698);
nand U12988 (N_12988,N_12851,N_12722);
nand U12989 (N_12989,N_12793,N_12889);
nand U12990 (N_12990,N_12867,N_12855);
nor U12991 (N_12991,N_12848,N_12650);
xor U12992 (N_12992,N_12675,N_12744);
nor U12993 (N_12993,N_12669,N_12662);
or U12994 (N_12994,N_12790,N_12830);
or U12995 (N_12995,N_12759,N_12618);
nor U12996 (N_12996,N_12719,N_12674);
nand U12997 (N_12997,N_12717,N_12876);
xnor U12998 (N_12998,N_12854,N_12787);
nor U12999 (N_12999,N_12695,N_12890);
nor U13000 (N_13000,N_12711,N_12601);
and U13001 (N_13001,N_12735,N_12667);
nor U13002 (N_13002,N_12644,N_12850);
and U13003 (N_13003,N_12768,N_12609);
nor U13004 (N_13004,N_12687,N_12745);
xor U13005 (N_13005,N_12802,N_12885);
or U13006 (N_13006,N_12806,N_12880);
nand U13007 (N_13007,N_12791,N_12627);
xnor U13008 (N_13008,N_12873,N_12874);
or U13009 (N_13009,N_12705,N_12714);
or U13010 (N_13010,N_12677,N_12882);
or U13011 (N_13011,N_12822,N_12866);
or U13012 (N_13012,N_12814,N_12712);
or U13013 (N_13013,N_12727,N_12783);
nor U13014 (N_13014,N_12626,N_12686);
nand U13015 (N_13015,N_12605,N_12755);
or U13016 (N_13016,N_12774,N_12641);
and U13017 (N_13017,N_12831,N_12721);
nand U13018 (N_13018,N_12704,N_12693);
or U13019 (N_13019,N_12707,N_12636);
or U13020 (N_13020,N_12872,N_12757);
or U13021 (N_13021,N_12703,N_12660);
nand U13022 (N_13022,N_12617,N_12657);
xnor U13023 (N_13023,N_12838,N_12842);
xor U13024 (N_13024,N_12748,N_12763);
xnor U13025 (N_13025,N_12762,N_12715);
xnor U13026 (N_13026,N_12776,N_12815);
and U13027 (N_13027,N_12845,N_12730);
and U13028 (N_13028,N_12653,N_12883);
nand U13029 (N_13029,N_12736,N_12897);
nand U13030 (N_13030,N_12620,N_12864);
and U13031 (N_13031,N_12786,N_12767);
nor U13032 (N_13032,N_12753,N_12654);
nor U13033 (N_13033,N_12737,N_12689);
or U13034 (N_13034,N_12898,N_12600);
nand U13035 (N_13035,N_12775,N_12785);
xnor U13036 (N_13036,N_12607,N_12651);
nor U13037 (N_13037,N_12764,N_12853);
nor U13038 (N_13038,N_12692,N_12616);
nor U13039 (N_13039,N_12811,N_12718);
and U13040 (N_13040,N_12738,N_12804);
xor U13041 (N_13041,N_12640,N_12886);
nand U13042 (N_13042,N_12865,N_12820);
xnor U13043 (N_13043,N_12878,N_12843);
xor U13044 (N_13044,N_12749,N_12658);
or U13045 (N_13045,N_12655,N_12803);
xnor U13046 (N_13046,N_12899,N_12819);
and U13047 (N_13047,N_12888,N_12664);
nor U13048 (N_13048,N_12633,N_12780);
xnor U13049 (N_13049,N_12846,N_12663);
nand U13050 (N_13050,N_12877,N_12883);
nand U13051 (N_13051,N_12702,N_12637);
xor U13052 (N_13052,N_12785,N_12886);
nand U13053 (N_13053,N_12830,N_12651);
and U13054 (N_13054,N_12636,N_12885);
xor U13055 (N_13055,N_12642,N_12773);
and U13056 (N_13056,N_12673,N_12659);
and U13057 (N_13057,N_12872,N_12644);
nor U13058 (N_13058,N_12668,N_12895);
xor U13059 (N_13059,N_12747,N_12816);
or U13060 (N_13060,N_12646,N_12711);
nor U13061 (N_13061,N_12895,N_12791);
nand U13062 (N_13062,N_12749,N_12789);
nand U13063 (N_13063,N_12677,N_12829);
nand U13064 (N_13064,N_12806,N_12794);
and U13065 (N_13065,N_12657,N_12782);
nor U13066 (N_13066,N_12803,N_12786);
or U13067 (N_13067,N_12807,N_12857);
nand U13068 (N_13068,N_12660,N_12729);
and U13069 (N_13069,N_12892,N_12634);
nand U13070 (N_13070,N_12826,N_12802);
nor U13071 (N_13071,N_12715,N_12748);
xor U13072 (N_13072,N_12831,N_12634);
xnor U13073 (N_13073,N_12889,N_12875);
nor U13074 (N_13074,N_12849,N_12844);
nand U13075 (N_13075,N_12618,N_12796);
and U13076 (N_13076,N_12859,N_12757);
and U13077 (N_13077,N_12899,N_12710);
or U13078 (N_13078,N_12643,N_12784);
and U13079 (N_13079,N_12882,N_12660);
and U13080 (N_13080,N_12696,N_12754);
or U13081 (N_13081,N_12692,N_12868);
nand U13082 (N_13082,N_12623,N_12654);
or U13083 (N_13083,N_12682,N_12837);
nand U13084 (N_13084,N_12822,N_12834);
and U13085 (N_13085,N_12716,N_12866);
nand U13086 (N_13086,N_12725,N_12625);
and U13087 (N_13087,N_12762,N_12600);
nor U13088 (N_13088,N_12681,N_12852);
nand U13089 (N_13089,N_12616,N_12704);
xnor U13090 (N_13090,N_12856,N_12822);
and U13091 (N_13091,N_12615,N_12620);
nand U13092 (N_13092,N_12631,N_12829);
xor U13093 (N_13093,N_12644,N_12756);
xnor U13094 (N_13094,N_12609,N_12832);
xor U13095 (N_13095,N_12858,N_12654);
xnor U13096 (N_13096,N_12825,N_12654);
and U13097 (N_13097,N_12855,N_12645);
and U13098 (N_13098,N_12820,N_12790);
nand U13099 (N_13099,N_12613,N_12663);
xnor U13100 (N_13100,N_12838,N_12757);
and U13101 (N_13101,N_12772,N_12655);
xnor U13102 (N_13102,N_12773,N_12847);
xor U13103 (N_13103,N_12825,N_12606);
nand U13104 (N_13104,N_12673,N_12858);
nand U13105 (N_13105,N_12787,N_12712);
or U13106 (N_13106,N_12702,N_12742);
and U13107 (N_13107,N_12715,N_12757);
xor U13108 (N_13108,N_12743,N_12736);
and U13109 (N_13109,N_12705,N_12760);
xnor U13110 (N_13110,N_12682,N_12849);
or U13111 (N_13111,N_12853,N_12803);
and U13112 (N_13112,N_12874,N_12861);
nor U13113 (N_13113,N_12818,N_12706);
xnor U13114 (N_13114,N_12609,N_12662);
and U13115 (N_13115,N_12679,N_12820);
or U13116 (N_13116,N_12894,N_12658);
and U13117 (N_13117,N_12810,N_12651);
xnor U13118 (N_13118,N_12876,N_12683);
xor U13119 (N_13119,N_12769,N_12774);
and U13120 (N_13120,N_12620,N_12654);
or U13121 (N_13121,N_12625,N_12846);
and U13122 (N_13122,N_12693,N_12681);
and U13123 (N_13123,N_12629,N_12898);
and U13124 (N_13124,N_12712,N_12755);
nor U13125 (N_13125,N_12824,N_12702);
xor U13126 (N_13126,N_12778,N_12854);
or U13127 (N_13127,N_12671,N_12878);
and U13128 (N_13128,N_12733,N_12776);
and U13129 (N_13129,N_12644,N_12810);
nor U13130 (N_13130,N_12722,N_12627);
nor U13131 (N_13131,N_12738,N_12764);
nand U13132 (N_13132,N_12659,N_12885);
nand U13133 (N_13133,N_12831,N_12751);
and U13134 (N_13134,N_12608,N_12770);
xnor U13135 (N_13135,N_12769,N_12756);
and U13136 (N_13136,N_12815,N_12810);
or U13137 (N_13137,N_12789,N_12792);
and U13138 (N_13138,N_12839,N_12784);
nor U13139 (N_13139,N_12722,N_12799);
and U13140 (N_13140,N_12713,N_12637);
nand U13141 (N_13141,N_12818,N_12890);
and U13142 (N_13142,N_12619,N_12813);
and U13143 (N_13143,N_12818,N_12773);
nand U13144 (N_13144,N_12722,N_12619);
xor U13145 (N_13145,N_12639,N_12858);
xor U13146 (N_13146,N_12710,N_12860);
or U13147 (N_13147,N_12885,N_12669);
nand U13148 (N_13148,N_12653,N_12821);
xnor U13149 (N_13149,N_12707,N_12659);
xor U13150 (N_13150,N_12814,N_12836);
xor U13151 (N_13151,N_12840,N_12803);
xor U13152 (N_13152,N_12601,N_12726);
nand U13153 (N_13153,N_12886,N_12749);
nand U13154 (N_13154,N_12668,N_12695);
nor U13155 (N_13155,N_12844,N_12812);
nor U13156 (N_13156,N_12875,N_12655);
or U13157 (N_13157,N_12635,N_12816);
nand U13158 (N_13158,N_12642,N_12699);
xor U13159 (N_13159,N_12758,N_12629);
nor U13160 (N_13160,N_12742,N_12725);
nor U13161 (N_13161,N_12820,N_12729);
and U13162 (N_13162,N_12615,N_12712);
xor U13163 (N_13163,N_12632,N_12899);
and U13164 (N_13164,N_12799,N_12816);
nand U13165 (N_13165,N_12771,N_12839);
xor U13166 (N_13166,N_12627,N_12810);
nand U13167 (N_13167,N_12894,N_12752);
nor U13168 (N_13168,N_12787,N_12823);
nor U13169 (N_13169,N_12864,N_12626);
nor U13170 (N_13170,N_12685,N_12749);
nand U13171 (N_13171,N_12641,N_12850);
and U13172 (N_13172,N_12737,N_12749);
nor U13173 (N_13173,N_12791,N_12613);
nand U13174 (N_13174,N_12669,N_12603);
nor U13175 (N_13175,N_12683,N_12635);
or U13176 (N_13176,N_12811,N_12883);
xnor U13177 (N_13177,N_12811,N_12664);
nor U13178 (N_13178,N_12773,N_12646);
or U13179 (N_13179,N_12697,N_12668);
nor U13180 (N_13180,N_12653,N_12648);
or U13181 (N_13181,N_12683,N_12721);
nand U13182 (N_13182,N_12755,N_12879);
nor U13183 (N_13183,N_12772,N_12615);
xor U13184 (N_13184,N_12617,N_12618);
nor U13185 (N_13185,N_12788,N_12672);
nand U13186 (N_13186,N_12706,N_12814);
or U13187 (N_13187,N_12898,N_12841);
and U13188 (N_13188,N_12772,N_12868);
nor U13189 (N_13189,N_12633,N_12728);
nor U13190 (N_13190,N_12840,N_12893);
nor U13191 (N_13191,N_12773,N_12822);
nand U13192 (N_13192,N_12753,N_12797);
or U13193 (N_13193,N_12663,N_12636);
nor U13194 (N_13194,N_12790,N_12827);
xor U13195 (N_13195,N_12887,N_12693);
xnor U13196 (N_13196,N_12823,N_12753);
and U13197 (N_13197,N_12839,N_12640);
and U13198 (N_13198,N_12767,N_12863);
xnor U13199 (N_13199,N_12688,N_12707);
nor U13200 (N_13200,N_13074,N_13016);
xnor U13201 (N_13201,N_13003,N_13006);
xnor U13202 (N_13202,N_12929,N_12981);
and U13203 (N_13203,N_12909,N_13154);
or U13204 (N_13204,N_13099,N_13014);
and U13205 (N_13205,N_12924,N_12991);
and U13206 (N_13206,N_13095,N_13189);
xnor U13207 (N_13207,N_13166,N_13011);
and U13208 (N_13208,N_13057,N_13182);
nand U13209 (N_13209,N_13158,N_12978);
nand U13210 (N_13210,N_13104,N_13174);
xnor U13211 (N_13211,N_13021,N_13114);
nand U13212 (N_13212,N_13181,N_13025);
xnor U13213 (N_13213,N_12999,N_13098);
and U13214 (N_13214,N_12920,N_13130);
or U13215 (N_13215,N_13116,N_13086);
or U13216 (N_13216,N_13050,N_13176);
nand U13217 (N_13217,N_13037,N_12917);
and U13218 (N_13218,N_12911,N_13190);
or U13219 (N_13219,N_12919,N_13083);
nor U13220 (N_13220,N_13162,N_13091);
xnor U13221 (N_13221,N_13070,N_13022);
xnor U13222 (N_13222,N_13069,N_13043);
or U13223 (N_13223,N_13065,N_13005);
xnor U13224 (N_13224,N_12961,N_13122);
or U13225 (N_13225,N_12923,N_12957);
and U13226 (N_13226,N_13113,N_13072);
nand U13227 (N_13227,N_13044,N_13109);
xor U13228 (N_13228,N_13096,N_13080);
nor U13229 (N_13229,N_13101,N_13157);
and U13230 (N_13230,N_13046,N_12966);
nand U13231 (N_13231,N_13103,N_12944);
and U13232 (N_13232,N_13150,N_12943);
xnor U13233 (N_13233,N_13068,N_13035);
nand U13234 (N_13234,N_13172,N_12928);
nand U13235 (N_13235,N_12922,N_12954);
nor U13236 (N_13236,N_13085,N_13087);
or U13237 (N_13237,N_13020,N_13160);
xnor U13238 (N_13238,N_13115,N_13028);
and U13239 (N_13239,N_13144,N_13141);
xnor U13240 (N_13240,N_13032,N_12962);
nor U13241 (N_13241,N_13030,N_13052);
or U13242 (N_13242,N_12987,N_13049);
and U13243 (N_13243,N_13169,N_13064);
xnor U13244 (N_13244,N_13004,N_12939);
or U13245 (N_13245,N_13017,N_12903);
nor U13246 (N_13246,N_12964,N_13075);
nand U13247 (N_13247,N_12960,N_12912);
nand U13248 (N_13248,N_13105,N_12998);
nand U13249 (N_13249,N_12951,N_13156);
xor U13250 (N_13250,N_12977,N_13077);
nand U13251 (N_13251,N_13094,N_13051);
nor U13252 (N_13252,N_13009,N_13082);
nor U13253 (N_13253,N_12915,N_13053);
xor U13254 (N_13254,N_12933,N_13121);
nor U13255 (N_13255,N_12916,N_13131);
or U13256 (N_13256,N_13000,N_13055);
or U13257 (N_13257,N_12972,N_12948);
or U13258 (N_13258,N_13112,N_13071);
and U13259 (N_13259,N_13159,N_13183);
and U13260 (N_13260,N_13041,N_12973);
or U13261 (N_13261,N_12988,N_12935);
or U13262 (N_13262,N_13061,N_12996);
and U13263 (N_13263,N_13117,N_12979);
nand U13264 (N_13264,N_12905,N_13171);
nor U13265 (N_13265,N_13067,N_13127);
nor U13266 (N_13266,N_12983,N_13018);
xor U13267 (N_13267,N_13066,N_12985);
xor U13268 (N_13268,N_12900,N_13140);
nand U13269 (N_13269,N_13111,N_13180);
nor U13270 (N_13270,N_12997,N_13084);
nor U13271 (N_13271,N_13060,N_13164);
nor U13272 (N_13272,N_13059,N_12982);
xor U13273 (N_13273,N_12971,N_13142);
or U13274 (N_13274,N_13048,N_13007);
and U13275 (N_13275,N_12927,N_13123);
and U13276 (N_13276,N_13073,N_13036);
nor U13277 (N_13277,N_13147,N_13078);
xnor U13278 (N_13278,N_13196,N_13042);
nor U13279 (N_13279,N_13175,N_13034);
nand U13280 (N_13280,N_13145,N_13155);
xnor U13281 (N_13281,N_13188,N_13143);
nor U13282 (N_13282,N_13081,N_13015);
nand U13283 (N_13283,N_13107,N_13139);
nor U13284 (N_13284,N_12934,N_12952);
nand U13285 (N_13285,N_13001,N_12993);
or U13286 (N_13286,N_12989,N_13187);
nor U13287 (N_13287,N_13199,N_12975);
or U13288 (N_13288,N_13178,N_12907);
and U13289 (N_13289,N_13118,N_13177);
nor U13290 (N_13290,N_13038,N_13108);
nand U13291 (N_13291,N_13152,N_13076);
or U13292 (N_13292,N_12930,N_13100);
nand U13293 (N_13293,N_12955,N_13029);
or U13294 (N_13294,N_13056,N_12970);
nand U13295 (N_13295,N_13023,N_12994);
and U13296 (N_13296,N_13184,N_12990);
xor U13297 (N_13297,N_12965,N_12901);
xnor U13298 (N_13298,N_13161,N_13024);
xor U13299 (N_13299,N_12913,N_13137);
or U13300 (N_13300,N_13008,N_12940);
nor U13301 (N_13301,N_13198,N_13179);
nor U13302 (N_13302,N_13165,N_13129);
or U13303 (N_13303,N_12968,N_13125);
nor U13304 (N_13304,N_12918,N_12932);
or U13305 (N_13305,N_13193,N_13092);
and U13306 (N_13306,N_12969,N_13058);
and U13307 (N_13307,N_13089,N_13136);
xnor U13308 (N_13308,N_13132,N_12984);
and U13309 (N_13309,N_13191,N_13135);
or U13310 (N_13310,N_13047,N_13192);
and U13311 (N_13311,N_13063,N_13170);
and U13312 (N_13312,N_12986,N_13149);
nand U13313 (N_13313,N_13033,N_13013);
xnor U13314 (N_13314,N_12945,N_13045);
or U13315 (N_13315,N_12906,N_13102);
and U13316 (N_13316,N_13133,N_13012);
xnor U13317 (N_13317,N_12910,N_13054);
xnor U13318 (N_13318,N_13138,N_13163);
nand U13319 (N_13319,N_13167,N_12995);
and U13320 (N_13320,N_13194,N_12980);
and U13321 (N_13321,N_13088,N_13090);
or U13322 (N_13322,N_12908,N_13195);
nand U13323 (N_13323,N_13134,N_12967);
xor U13324 (N_13324,N_13173,N_12921);
nor U13325 (N_13325,N_13126,N_13151);
and U13326 (N_13326,N_13039,N_12963);
nand U13327 (N_13327,N_12941,N_12925);
xor U13328 (N_13328,N_12953,N_12938);
nor U13329 (N_13329,N_12992,N_12942);
xnor U13330 (N_13330,N_13119,N_13019);
nand U13331 (N_13331,N_12958,N_12937);
and U13332 (N_13332,N_13106,N_13079);
nand U13333 (N_13333,N_13146,N_12950);
nor U13334 (N_13334,N_13062,N_12974);
and U13335 (N_13335,N_13027,N_12902);
or U13336 (N_13336,N_13186,N_12947);
nand U13337 (N_13337,N_13110,N_13097);
nor U13338 (N_13338,N_13197,N_13002);
xnor U13339 (N_13339,N_13040,N_12959);
nor U13340 (N_13340,N_13128,N_13168);
nand U13341 (N_13341,N_12914,N_13093);
nand U13342 (N_13342,N_12946,N_13148);
xor U13343 (N_13343,N_13153,N_13010);
and U13344 (N_13344,N_13124,N_12936);
and U13345 (N_13345,N_13026,N_12956);
nor U13346 (N_13346,N_12931,N_12904);
nor U13347 (N_13347,N_12949,N_12926);
xor U13348 (N_13348,N_13031,N_12976);
or U13349 (N_13349,N_13120,N_13185);
nand U13350 (N_13350,N_13086,N_13144);
or U13351 (N_13351,N_13164,N_12999);
xor U13352 (N_13352,N_12991,N_12973);
and U13353 (N_13353,N_12972,N_12924);
or U13354 (N_13354,N_13187,N_13009);
and U13355 (N_13355,N_12930,N_12949);
or U13356 (N_13356,N_13119,N_12986);
nand U13357 (N_13357,N_12927,N_13042);
and U13358 (N_13358,N_12992,N_13091);
and U13359 (N_13359,N_13053,N_13164);
nor U13360 (N_13360,N_12912,N_13098);
nand U13361 (N_13361,N_12946,N_12905);
or U13362 (N_13362,N_12972,N_13101);
nor U13363 (N_13363,N_13048,N_13016);
nand U13364 (N_13364,N_13160,N_13151);
or U13365 (N_13365,N_12905,N_13061);
nand U13366 (N_13366,N_13118,N_12919);
and U13367 (N_13367,N_12968,N_13091);
and U13368 (N_13368,N_13170,N_13002);
nand U13369 (N_13369,N_13038,N_13091);
and U13370 (N_13370,N_13174,N_13141);
nor U13371 (N_13371,N_13094,N_12953);
nand U13372 (N_13372,N_13056,N_12911);
or U13373 (N_13373,N_13156,N_13093);
and U13374 (N_13374,N_12968,N_12956);
nand U13375 (N_13375,N_13176,N_13083);
nor U13376 (N_13376,N_13030,N_12904);
nand U13377 (N_13377,N_13003,N_13122);
or U13378 (N_13378,N_12958,N_13040);
or U13379 (N_13379,N_12944,N_13024);
nor U13380 (N_13380,N_13061,N_13187);
xnor U13381 (N_13381,N_12973,N_12979);
xor U13382 (N_13382,N_13035,N_13171);
or U13383 (N_13383,N_12999,N_13149);
xor U13384 (N_13384,N_13099,N_12944);
nand U13385 (N_13385,N_12925,N_12912);
nand U13386 (N_13386,N_13196,N_12908);
xnor U13387 (N_13387,N_12984,N_13041);
or U13388 (N_13388,N_13144,N_13149);
xor U13389 (N_13389,N_13028,N_12916);
or U13390 (N_13390,N_12941,N_12981);
nand U13391 (N_13391,N_13166,N_12911);
and U13392 (N_13392,N_12963,N_13071);
xnor U13393 (N_13393,N_13006,N_13137);
xor U13394 (N_13394,N_12915,N_13196);
nor U13395 (N_13395,N_12905,N_12954);
nor U13396 (N_13396,N_12986,N_13136);
nand U13397 (N_13397,N_13116,N_13046);
xor U13398 (N_13398,N_13130,N_13162);
xnor U13399 (N_13399,N_12974,N_13110);
nand U13400 (N_13400,N_13125,N_13118);
xnor U13401 (N_13401,N_12974,N_12926);
and U13402 (N_13402,N_13074,N_13094);
nand U13403 (N_13403,N_12980,N_12915);
or U13404 (N_13404,N_13123,N_12923);
and U13405 (N_13405,N_13197,N_13037);
or U13406 (N_13406,N_12924,N_13083);
and U13407 (N_13407,N_13141,N_13138);
or U13408 (N_13408,N_13015,N_12905);
or U13409 (N_13409,N_13187,N_12999);
or U13410 (N_13410,N_13189,N_13153);
xor U13411 (N_13411,N_12906,N_13059);
xnor U13412 (N_13412,N_13112,N_13026);
or U13413 (N_13413,N_13193,N_13056);
and U13414 (N_13414,N_12918,N_13122);
and U13415 (N_13415,N_12941,N_12931);
or U13416 (N_13416,N_12944,N_12918);
and U13417 (N_13417,N_12958,N_13111);
and U13418 (N_13418,N_12922,N_13121);
nor U13419 (N_13419,N_12944,N_13187);
nand U13420 (N_13420,N_13011,N_13155);
and U13421 (N_13421,N_12980,N_13085);
nand U13422 (N_13422,N_13156,N_13166);
nor U13423 (N_13423,N_13162,N_13045);
and U13424 (N_13424,N_12956,N_12912);
xor U13425 (N_13425,N_13015,N_13108);
and U13426 (N_13426,N_13172,N_12918);
or U13427 (N_13427,N_13022,N_12991);
xnor U13428 (N_13428,N_13030,N_13062);
or U13429 (N_13429,N_13040,N_13060);
xor U13430 (N_13430,N_12953,N_13023);
nor U13431 (N_13431,N_13080,N_13139);
nand U13432 (N_13432,N_12910,N_13137);
nand U13433 (N_13433,N_13074,N_12994);
nor U13434 (N_13434,N_12904,N_13086);
or U13435 (N_13435,N_12989,N_13047);
nor U13436 (N_13436,N_12964,N_12974);
nor U13437 (N_13437,N_12992,N_12931);
or U13438 (N_13438,N_12992,N_13001);
nor U13439 (N_13439,N_13153,N_13191);
and U13440 (N_13440,N_12928,N_13060);
xnor U13441 (N_13441,N_13129,N_13195);
nand U13442 (N_13442,N_13042,N_12913);
and U13443 (N_13443,N_12946,N_13025);
nand U13444 (N_13444,N_12981,N_13119);
and U13445 (N_13445,N_13199,N_13144);
and U13446 (N_13446,N_13118,N_13023);
or U13447 (N_13447,N_12997,N_13077);
and U13448 (N_13448,N_13189,N_12949);
nor U13449 (N_13449,N_13058,N_13195);
xor U13450 (N_13450,N_12982,N_12917);
or U13451 (N_13451,N_13111,N_13106);
and U13452 (N_13452,N_13047,N_12949);
or U13453 (N_13453,N_13127,N_13179);
nor U13454 (N_13454,N_13088,N_13018);
xnor U13455 (N_13455,N_12998,N_13070);
nor U13456 (N_13456,N_12938,N_13171);
nor U13457 (N_13457,N_12914,N_12974);
nor U13458 (N_13458,N_12940,N_12984);
and U13459 (N_13459,N_13012,N_13044);
or U13460 (N_13460,N_13015,N_13045);
or U13461 (N_13461,N_13181,N_12905);
and U13462 (N_13462,N_12963,N_13022);
nor U13463 (N_13463,N_12929,N_13124);
xnor U13464 (N_13464,N_13067,N_13003);
xor U13465 (N_13465,N_13067,N_13042);
or U13466 (N_13466,N_12971,N_13037);
xor U13467 (N_13467,N_13077,N_13022);
nand U13468 (N_13468,N_13162,N_12903);
or U13469 (N_13469,N_13018,N_12904);
xor U13470 (N_13470,N_13131,N_12991);
nor U13471 (N_13471,N_12914,N_12934);
nand U13472 (N_13472,N_12995,N_13013);
nor U13473 (N_13473,N_13142,N_12909);
xor U13474 (N_13474,N_13053,N_13152);
or U13475 (N_13475,N_13141,N_13038);
nand U13476 (N_13476,N_13134,N_12954);
and U13477 (N_13477,N_12995,N_13182);
xnor U13478 (N_13478,N_12903,N_12948);
or U13479 (N_13479,N_13102,N_13161);
xnor U13480 (N_13480,N_12932,N_13014);
nand U13481 (N_13481,N_13074,N_13045);
xor U13482 (N_13482,N_12901,N_12908);
or U13483 (N_13483,N_13148,N_13049);
and U13484 (N_13484,N_13103,N_13087);
nor U13485 (N_13485,N_13160,N_13054);
xnor U13486 (N_13486,N_13009,N_13116);
or U13487 (N_13487,N_13119,N_13104);
or U13488 (N_13488,N_12985,N_12926);
nor U13489 (N_13489,N_12911,N_13194);
and U13490 (N_13490,N_12993,N_13123);
and U13491 (N_13491,N_13129,N_13105);
nor U13492 (N_13492,N_12957,N_13128);
nor U13493 (N_13493,N_13163,N_12949);
or U13494 (N_13494,N_13187,N_13091);
or U13495 (N_13495,N_13025,N_13104);
nor U13496 (N_13496,N_12933,N_13193);
or U13497 (N_13497,N_13083,N_12929);
or U13498 (N_13498,N_13166,N_13115);
and U13499 (N_13499,N_12952,N_13084);
xor U13500 (N_13500,N_13335,N_13364);
nand U13501 (N_13501,N_13458,N_13366);
nand U13502 (N_13502,N_13444,N_13322);
or U13503 (N_13503,N_13202,N_13467);
nor U13504 (N_13504,N_13445,N_13496);
nor U13505 (N_13505,N_13280,N_13422);
xor U13506 (N_13506,N_13240,N_13242);
and U13507 (N_13507,N_13468,N_13227);
or U13508 (N_13508,N_13442,N_13420);
and U13509 (N_13509,N_13218,N_13469);
and U13510 (N_13510,N_13315,N_13248);
xor U13511 (N_13511,N_13474,N_13452);
or U13512 (N_13512,N_13303,N_13299);
or U13513 (N_13513,N_13284,N_13257);
or U13514 (N_13514,N_13300,N_13493);
and U13515 (N_13515,N_13358,N_13217);
nor U13516 (N_13516,N_13352,N_13282);
or U13517 (N_13517,N_13237,N_13373);
and U13518 (N_13518,N_13292,N_13250);
xor U13519 (N_13519,N_13255,N_13367);
or U13520 (N_13520,N_13409,N_13351);
xor U13521 (N_13521,N_13285,N_13392);
nor U13522 (N_13522,N_13453,N_13421);
nor U13523 (N_13523,N_13375,N_13414);
nand U13524 (N_13524,N_13370,N_13490);
nor U13525 (N_13525,N_13349,N_13447);
or U13526 (N_13526,N_13321,N_13244);
xnor U13527 (N_13527,N_13419,N_13354);
and U13528 (N_13528,N_13434,N_13332);
and U13529 (N_13529,N_13397,N_13441);
xor U13530 (N_13530,N_13439,N_13215);
nor U13531 (N_13531,N_13395,N_13462);
nand U13532 (N_13532,N_13219,N_13473);
nor U13533 (N_13533,N_13340,N_13334);
nand U13534 (N_13534,N_13376,N_13211);
and U13535 (N_13535,N_13466,N_13247);
or U13536 (N_13536,N_13446,N_13231);
or U13537 (N_13537,N_13311,N_13221);
nand U13538 (N_13538,N_13296,N_13293);
or U13539 (N_13539,N_13341,N_13314);
nand U13540 (N_13540,N_13382,N_13239);
and U13541 (N_13541,N_13460,N_13309);
or U13542 (N_13542,N_13384,N_13472);
or U13543 (N_13543,N_13200,N_13302);
xnor U13544 (N_13544,N_13436,N_13264);
nand U13545 (N_13545,N_13383,N_13417);
and U13546 (N_13546,N_13222,N_13353);
nor U13547 (N_13547,N_13440,N_13203);
nor U13548 (N_13548,N_13254,N_13438);
and U13549 (N_13549,N_13249,N_13450);
nor U13550 (N_13550,N_13325,N_13412);
xnor U13551 (N_13551,N_13330,N_13386);
or U13552 (N_13552,N_13430,N_13301);
nand U13553 (N_13553,N_13324,N_13443);
and U13554 (N_13554,N_13210,N_13258);
nand U13555 (N_13555,N_13333,N_13475);
or U13556 (N_13556,N_13357,N_13269);
or U13557 (N_13557,N_13253,N_13377);
and U13558 (N_13558,N_13424,N_13429);
nand U13559 (N_13559,N_13489,N_13274);
xor U13560 (N_13560,N_13278,N_13359);
or U13561 (N_13561,N_13497,N_13437);
and U13562 (N_13562,N_13213,N_13481);
nor U13563 (N_13563,N_13262,N_13245);
nor U13564 (N_13564,N_13279,N_13336);
and U13565 (N_13565,N_13480,N_13476);
or U13566 (N_13566,N_13317,N_13337);
or U13567 (N_13567,N_13344,N_13312);
nand U13568 (N_13568,N_13319,N_13362);
nand U13569 (N_13569,N_13294,N_13291);
or U13570 (N_13570,N_13298,N_13492);
and U13571 (N_13571,N_13243,N_13426);
nor U13572 (N_13572,N_13451,N_13459);
nand U13573 (N_13573,N_13410,N_13204);
nand U13574 (N_13574,N_13347,N_13295);
nand U13575 (N_13575,N_13498,N_13246);
nor U13576 (N_13576,N_13477,N_13380);
nor U13577 (N_13577,N_13495,N_13224);
nand U13578 (N_13578,N_13394,N_13273);
xnor U13579 (N_13579,N_13270,N_13307);
and U13580 (N_13580,N_13398,N_13406);
or U13581 (N_13581,N_13327,N_13401);
and U13582 (N_13582,N_13281,N_13234);
nor U13583 (N_13583,N_13431,N_13252);
or U13584 (N_13584,N_13400,N_13486);
and U13585 (N_13585,N_13407,N_13471);
nand U13586 (N_13586,N_13360,N_13350);
nand U13587 (N_13587,N_13220,N_13287);
nand U13588 (N_13588,N_13416,N_13484);
nor U13589 (N_13589,N_13404,N_13478);
nor U13590 (N_13590,N_13232,N_13365);
and U13591 (N_13591,N_13313,N_13433);
and U13592 (N_13592,N_13355,N_13361);
or U13593 (N_13593,N_13356,N_13374);
nor U13594 (N_13594,N_13263,N_13228);
and U13595 (N_13595,N_13230,N_13449);
xor U13596 (N_13596,N_13212,N_13372);
or U13597 (N_13597,N_13241,N_13205);
nand U13598 (N_13598,N_13229,N_13448);
and U13599 (N_13599,N_13415,N_13368);
and U13600 (N_13600,N_13271,N_13316);
or U13601 (N_13601,N_13482,N_13206);
xnor U13602 (N_13602,N_13487,N_13290);
or U13603 (N_13603,N_13207,N_13331);
nand U13604 (N_13604,N_13251,N_13209);
or U13605 (N_13605,N_13223,N_13308);
nor U13606 (N_13606,N_13260,N_13304);
and U13607 (N_13607,N_13328,N_13310);
nand U13608 (N_13608,N_13432,N_13379);
and U13609 (N_13609,N_13286,N_13268);
nor U13610 (N_13610,N_13236,N_13387);
xnor U13611 (N_13611,N_13411,N_13413);
nand U13612 (N_13612,N_13235,N_13369);
nor U13613 (N_13613,N_13454,N_13485);
and U13614 (N_13614,N_13435,N_13388);
or U13615 (N_13615,N_13266,N_13348);
and U13616 (N_13616,N_13423,N_13339);
or U13617 (N_13617,N_13425,N_13233);
xor U13618 (N_13618,N_13488,N_13399);
and U13619 (N_13619,N_13297,N_13214);
xor U13620 (N_13620,N_13216,N_13342);
xnor U13621 (N_13621,N_13455,N_13201);
nor U13622 (N_13622,N_13463,N_13346);
or U13623 (N_13623,N_13385,N_13343);
and U13624 (N_13624,N_13403,N_13378);
or U13625 (N_13625,N_13329,N_13272);
and U13626 (N_13626,N_13289,N_13326);
or U13627 (N_13627,N_13256,N_13418);
nand U13628 (N_13628,N_13499,N_13470);
or U13629 (N_13629,N_13491,N_13371);
nor U13630 (N_13630,N_13265,N_13226);
xnor U13631 (N_13631,N_13456,N_13277);
or U13632 (N_13632,N_13338,N_13428);
or U13633 (N_13633,N_13276,N_13461);
nor U13634 (N_13634,N_13318,N_13381);
nor U13635 (N_13635,N_13391,N_13267);
nand U13636 (N_13636,N_13320,N_13389);
nor U13637 (N_13637,N_13283,N_13494);
or U13638 (N_13638,N_13457,N_13479);
or U13639 (N_13639,N_13261,N_13405);
or U13640 (N_13640,N_13225,N_13427);
nor U13641 (N_13641,N_13305,N_13464);
and U13642 (N_13642,N_13465,N_13402);
and U13643 (N_13643,N_13208,N_13306);
or U13644 (N_13644,N_13238,N_13393);
nand U13645 (N_13645,N_13483,N_13363);
xnor U13646 (N_13646,N_13408,N_13345);
nor U13647 (N_13647,N_13259,N_13275);
or U13648 (N_13648,N_13288,N_13396);
or U13649 (N_13649,N_13323,N_13390);
nor U13650 (N_13650,N_13320,N_13273);
nand U13651 (N_13651,N_13424,N_13482);
or U13652 (N_13652,N_13450,N_13357);
and U13653 (N_13653,N_13343,N_13369);
and U13654 (N_13654,N_13493,N_13263);
nor U13655 (N_13655,N_13299,N_13210);
xnor U13656 (N_13656,N_13469,N_13247);
or U13657 (N_13657,N_13333,N_13451);
or U13658 (N_13658,N_13387,N_13370);
xnor U13659 (N_13659,N_13423,N_13231);
nand U13660 (N_13660,N_13209,N_13328);
nor U13661 (N_13661,N_13396,N_13321);
or U13662 (N_13662,N_13449,N_13469);
and U13663 (N_13663,N_13283,N_13437);
xor U13664 (N_13664,N_13469,N_13261);
nand U13665 (N_13665,N_13401,N_13355);
nor U13666 (N_13666,N_13370,N_13427);
nor U13667 (N_13667,N_13317,N_13476);
and U13668 (N_13668,N_13410,N_13400);
and U13669 (N_13669,N_13495,N_13382);
xor U13670 (N_13670,N_13454,N_13443);
xor U13671 (N_13671,N_13327,N_13431);
xor U13672 (N_13672,N_13333,N_13452);
nand U13673 (N_13673,N_13379,N_13241);
nand U13674 (N_13674,N_13388,N_13331);
xor U13675 (N_13675,N_13347,N_13466);
nor U13676 (N_13676,N_13434,N_13338);
nor U13677 (N_13677,N_13246,N_13273);
and U13678 (N_13678,N_13462,N_13322);
xnor U13679 (N_13679,N_13360,N_13486);
and U13680 (N_13680,N_13423,N_13259);
nand U13681 (N_13681,N_13456,N_13474);
and U13682 (N_13682,N_13284,N_13245);
and U13683 (N_13683,N_13260,N_13317);
or U13684 (N_13684,N_13357,N_13367);
and U13685 (N_13685,N_13255,N_13478);
xnor U13686 (N_13686,N_13251,N_13287);
nand U13687 (N_13687,N_13394,N_13475);
xnor U13688 (N_13688,N_13336,N_13385);
nand U13689 (N_13689,N_13232,N_13450);
xor U13690 (N_13690,N_13415,N_13251);
or U13691 (N_13691,N_13318,N_13271);
nand U13692 (N_13692,N_13306,N_13238);
or U13693 (N_13693,N_13479,N_13476);
nand U13694 (N_13694,N_13272,N_13289);
nand U13695 (N_13695,N_13380,N_13413);
or U13696 (N_13696,N_13430,N_13265);
or U13697 (N_13697,N_13211,N_13416);
xor U13698 (N_13698,N_13435,N_13398);
nor U13699 (N_13699,N_13231,N_13311);
nor U13700 (N_13700,N_13397,N_13458);
and U13701 (N_13701,N_13396,N_13443);
nand U13702 (N_13702,N_13356,N_13264);
and U13703 (N_13703,N_13329,N_13347);
xor U13704 (N_13704,N_13282,N_13476);
or U13705 (N_13705,N_13489,N_13223);
and U13706 (N_13706,N_13240,N_13224);
xor U13707 (N_13707,N_13315,N_13450);
nor U13708 (N_13708,N_13405,N_13226);
nand U13709 (N_13709,N_13298,N_13417);
or U13710 (N_13710,N_13257,N_13288);
xor U13711 (N_13711,N_13481,N_13398);
xor U13712 (N_13712,N_13218,N_13306);
xnor U13713 (N_13713,N_13211,N_13241);
and U13714 (N_13714,N_13396,N_13417);
xor U13715 (N_13715,N_13392,N_13485);
and U13716 (N_13716,N_13350,N_13364);
or U13717 (N_13717,N_13441,N_13475);
nor U13718 (N_13718,N_13287,N_13349);
nand U13719 (N_13719,N_13279,N_13376);
or U13720 (N_13720,N_13261,N_13262);
nor U13721 (N_13721,N_13373,N_13301);
nor U13722 (N_13722,N_13321,N_13217);
nor U13723 (N_13723,N_13474,N_13298);
or U13724 (N_13724,N_13470,N_13383);
xor U13725 (N_13725,N_13367,N_13340);
and U13726 (N_13726,N_13324,N_13407);
or U13727 (N_13727,N_13307,N_13321);
or U13728 (N_13728,N_13415,N_13494);
and U13729 (N_13729,N_13350,N_13493);
and U13730 (N_13730,N_13277,N_13304);
xor U13731 (N_13731,N_13301,N_13329);
xnor U13732 (N_13732,N_13334,N_13420);
and U13733 (N_13733,N_13313,N_13237);
nor U13734 (N_13734,N_13204,N_13340);
and U13735 (N_13735,N_13313,N_13406);
nor U13736 (N_13736,N_13488,N_13299);
xor U13737 (N_13737,N_13238,N_13421);
nand U13738 (N_13738,N_13270,N_13370);
nand U13739 (N_13739,N_13267,N_13335);
or U13740 (N_13740,N_13219,N_13484);
or U13741 (N_13741,N_13475,N_13380);
and U13742 (N_13742,N_13299,N_13219);
nor U13743 (N_13743,N_13394,N_13485);
and U13744 (N_13744,N_13348,N_13201);
and U13745 (N_13745,N_13351,N_13244);
xor U13746 (N_13746,N_13286,N_13302);
nor U13747 (N_13747,N_13486,N_13461);
and U13748 (N_13748,N_13229,N_13458);
or U13749 (N_13749,N_13363,N_13463);
or U13750 (N_13750,N_13498,N_13226);
or U13751 (N_13751,N_13377,N_13331);
or U13752 (N_13752,N_13351,N_13369);
nor U13753 (N_13753,N_13324,N_13498);
or U13754 (N_13754,N_13451,N_13296);
and U13755 (N_13755,N_13286,N_13252);
nor U13756 (N_13756,N_13219,N_13400);
or U13757 (N_13757,N_13277,N_13426);
nor U13758 (N_13758,N_13333,N_13484);
nor U13759 (N_13759,N_13398,N_13420);
and U13760 (N_13760,N_13350,N_13321);
or U13761 (N_13761,N_13386,N_13249);
nor U13762 (N_13762,N_13307,N_13214);
xor U13763 (N_13763,N_13451,N_13367);
nand U13764 (N_13764,N_13341,N_13220);
nor U13765 (N_13765,N_13436,N_13393);
nand U13766 (N_13766,N_13251,N_13283);
or U13767 (N_13767,N_13486,N_13369);
and U13768 (N_13768,N_13251,N_13311);
and U13769 (N_13769,N_13491,N_13219);
nand U13770 (N_13770,N_13250,N_13333);
nand U13771 (N_13771,N_13482,N_13488);
nor U13772 (N_13772,N_13381,N_13330);
and U13773 (N_13773,N_13484,N_13413);
nand U13774 (N_13774,N_13463,N_13273);
nor U13775 (N_13775,N_13490,N_13329);
nand U13776 (N_13776,N_13235,N_13347);
xor U13777 (N_13777,N_13286,N_13210);
nand U13778 (N_13778,N_13459,N_13209);
and U13779 (N_13779,N_13259,N_13415);
and U13780 (N_13780,N_13455,N_13301);
or U13781 (N_13781,N_13241,N_13346);
nor U13782 (N_13782,N_13243,N_13325);
nand U13783 (N_13783,N_13442,N_13497);
or U13784 (N_13784,N_13467,N_13409);
nor U13785 (N_13785,N_13328,N_13408);
xor U13786 (N_13786,N_13485,N_13311);
nand U13787 (N_13787,N_13427,N_13463);
nor U13788 (N_13788,N_13310,N_13245);
nor U13789 (N_13789,N_13295,N_13289);
and U13790 (N_13790,N_13210,N_13352);
and U13791 (N_13791,N_13373,N_13452);
nor U13792 (N_13792,N_13342,N_13255);
or U13793 (N_13793,N_13277,N_13309);
and U13794 (N_13794,N_13429,N_13334);
nor U13795 (N_13795,N_13475,N_13495);
nor U13796 (N_13796,N_13343,N_13498);
xor U13797 (N_13797,N_13480,N_13479);
nand U13798 (N_13798,N_13374,N_13361);
xnor U13799 (N_13799,N_13433,N_13346);
nand U13800 (N_13800,N_13744,N_13613);
nor U13801 (N_13801,N_13611,N_13711);
and U13802 (N_13802,N_13630,N_13547);
xnor U13803 (N_13803,N_13799,N_13761);
or U13804 (N_13804,N_13790,N_13747);
nor U13805 (N_13805,N_13581,N_13692);
nand U13806 (N_13806,N_13776,N_13794);
and U13807 (N_13807,N_13762,N_13585);
or U13808 (N_13808,N_13737,N_13636);
nor U13809 (N_13809,N_13663,N_13622);
or U13810 (N_13810,N_13798,N_13774);
xnor U13811 (N_13811,N_13796,N_13669);
or U13812 (N_13812,N_13781,N_13722);
xor U13813 (N_13813,N_13589,N_13536);
nand U13814 (N_13814,N_13600,N_13787);
nand U13815 (N_13815,N_13683,N_13700);
and U13816 (N_13816,N_13518,N_13727);
nand U13817 (N_13817,N_13690,N_13642);
xnor U13818 (N_13818,N_13718,N_13745);
nor U13819 (N_13819,N_13563,N_13608);
or U13820 (N_13820,N_13684,N_13785);
nor U13821 (N_13821,N_13521,N_13674);
and U13822 (N_13822,N_13623,N_13549);
nand U13823 (N_13823,N_13621,N_13609);
and U13824 (N_13824,N_13569,N_13716);
nand U13825 (N_13825,N_13616,N_13657);
or U13826 (N_13826,N_13558,N_13707);
and U13827 (N_13827,N_13784,N_13594);
nand U13828 (N_13828,N_13542,N_13702);
and U13829 (N_13829,N_13713,N_13618);
and U13830 (N_13830,N_13695,N_13668);
or U13831 (N_13831,N_13714,N_13527);
xor U13832 (N_13832,N_13640,N_13502);
xnor U13833 (N_13833,N_13561,N_13773);
nand U13834 (N_13834,N_13780,N_13541);
nand U13835 (N_13835,N_13634,N_13679);
nand U13836 (N_13836,N_13673,N_13649);
xnor U13837 (N_13837,N_13658,N_13544);
nor U13838 (N_13838,N_13672,N_13633);
and U13839 (N_13839,N_13639,N_13537);
xnor U13840 (N_13840,N_13705,N_13763);
nand U13841 (N_13841,N_13726,N_13554);
xor U13842 (N_13842,N_13660,N_13550);
and U13843 (N_13843,N_13789,N_13689);
or U13844 (N_13844,N_13530,N_13520);
xnor U13845 (N_13845,N_13746,N_13641);
and U13846 (N_13846,N_13645,N_13715);
nand U13847 (N_13847,N_13562,N_13666);
or U13848 (N_13848,N_13506,N_13548);
and U13849 (N_13849,N_13756,N_13771);
nand U13850 (N_13850,N_13595,N_13748);
or U13851 (N_13851,N_13768,N_13652);
and U13852 (N_13852,N_13680,N_13632);
nor U13853 (N_13853,N_13535,N_13731);
or U13854 (N_13854,N_13571,N_13532);
or U13855 (N_13855,N_13741,N_13597);
xnor U13856 (N_13856,N_13511,N_13583);
or U13857 (N_13857,N_13661,N_13693);
and U13858 (N_13858,N_13650,N_13709);
xor U13859 (N_13859,N_13753,N_13625);
xor U13860 (N_13860,N_13552,N_13540);
xor U13861 (N_13861,N_13729,N_13777);
nand U13862 (N_13862,N_13531,N_13512);
or U13863 (N_13863,N_13566,N_13792);
xnor U13864 (N_13864,N_13703,N_13628);
xor U13865 (N_13865,N_13637,N_13783);
nand U13866 (N_13866,N_13648,N_13617);
nor U13867 (N_13867,N_13720,N_13681);
or U13868 (N_13868,N_13643,N_13578);
nor U13869 (N_13869,N_13769,N_13685);
nand U13870 (N_13870,N_13739,N_13651);
nor U13871 (N_13871,N_13507,N_13534);
or U13872 (N_13872,N_13717,N_13691);
xnor U13873 (N_13873,N_13513,N_13508);
nor U13874 (N_13874,N_13570,N_13568);
xnor U13875 (N_13875,N_13665,N_13515);
or U13876 (N_13876,N_13797,N_13754);
and U13877 (N_13877,N_13580,N_13559);
nand U13878 (N_13878,N_13606,N_13565);
nor U13879 (N_13879,N_13601,N_13553);
nand U13880 (N_13880,N_13503,N_13505);
xnor U13881 (N_13881,N_13675,N_13593);
xor U13882 (N_13882,N_13765,N_13587);
nor U13883 (N_13883,N_13759,N_13500);
nand U13884 (N_13884,N_13750,N_13701);
xor U13885 (N_13885,N_13529,N_13599);
xnor U13886 (N_13886,N_13574,N_13626);
or U13887 (N_13887,N_13667,N_13671);
or U13888 (N_13888,N_13696,N_13670);
xor U13889 (N_13889,N_13539,N_13560);
nor U13890 (N_13890,N_13749,N_13743);
or U13891 (N_13891,N_13712,N_13575);
nor U13892 (N_13892,N_13579,N_13688);
nand U13893 (N_13893,N_13708,N_13545);
or U13894 (N_13894,N_13786,N_13721);
xor U13895 (N_13895,N_13591,N_13504);
xnor U13896 (N_13896,N_13778,N_13653);
nand U13897 (N_13897,N_13704,N_13576);
xnor U13898 (N_13898,N_13620,N_13733);
or U13899 (N_13899,N_13751,N_13772);
xor U13900 (N_13900,N_13647,N_13619);
xor U13901 (N_13901,N_13742,N_13728);
or U13902 (N_13902,N_13723,N_13629);
nor U13903 (N_13903,N_13698,N_13584);
xnor U13904 (N_13904,N_13551,N_13662);
nand U13905 (N_13905,N_13755,N_13725);
nor U13906 (N_13906,N_13795,N_13596);
and U13907 (N_13907,N_13546,N_13706);
or U13908 (N_13908,N_13510,N_13555);
and U13909 (N_13909,N_13735,N_13697);
or U13910 (N_13910,N_13738,N_13627);
and U13911 (N_13911,N_13614,N_13710);
or U13912 (N_13912,N_13770,N_13528);
nor U13913 (N_13913,N_13590,N_13564);
xnor U13914 (N_13914,N_13501,N_13644);
xnor U13915 (N_13915,N_13730,N_13538);
and U13916 (N_13916,N_13752,N_13682);
nand U13917 (N_13917,N_13582,N_13516);
nand U13918 (N_13918,N_13646,N_13740);
or U13919 (N_13919,N_13519,N_13655);
and U13920 (N_13920,N_13719,N_13677);
nor U13921 (N_13921,N_13602,N_13514);
and U13922 (N_13922,N_13557,N_13615);
nor U13923 (N_13923,N_13543,N_13631);
nand U13924 (N_13924,N_13699,N_13654);
or U13925 (N_13925,N_13760,N_13577);
and U13926 (N_13926,N_13757,N_13694);
xor U13927 (N_13927,N_13604,N_13605);
or U13928 (N_13928,N_13509,N_13767);
nor U13929 (N_13929,N_13573,N_13524);
or U13930 (N_13930,N_13775,N_13624);
nand U13931 (N_13931,N_13724,N_13676);
or U13932 (N_13932,N_13758,N_13793);
nor U13933 (N_13933,N_13686,N_13687);
or U13934 (N_13934,N_13607,N_13782);
nor U13935 (N_13935,N_13664,N_13526);
or U13936 (N_13936,N_13659,N_13791);
nor U13937 (N_13937,N_13567,N_13764);
nand U13938 (N_13938,N_13588,N_13788);
and U13939 (N_13939,N_13635,N_13525);
and U13940 (N_13940,N_13638,N_13517);
and U13941 (N_13941,N_13592,N_13523);
nand U13942 (N_13942,N_13603,N_13556);
and U13943 (N_13943,N_13610,N_13736);
xor U13944 (N_13944,N_13586,N_13522);
nor U13945 (N_13945,N_13572,N_13656);
or U13946 (N_13946,N_13533,N_13598);
nand U13947 (N_13947,N_13766,N_13732);
and U13948 (N_13948,N_13779,N_13678);
and U13949 (N_13949,N_13612,N_13734);
or U13950 (N_13950,N_13796,N_13682);
or U13951 (N_13951,N_13711,N_13510);
nor U13952 (N_13952,N_13690,N_13623);
xor U13953 (N_13953,N_13616,N_13547);
and U13954 (N_13954,N_13666,N_13786);
nor U13955 (N_13955,N_13618,N_13752);
xor U13956 (N_13956,N_13610,N_13524);
and U13957 (N_13957,N_13672,N_13623);
or U13958 (N_13958,N_13583,N_13549);
xnor U13959 (N_13959,N_13504,N_13520);
and U13960 (N_13960,N_13656,N_13559);
nand U13961 (N_13961,N_13653,N_13777);
and U13962 (N_13962,N_13744,N_13544);
or U13963 (N_13963,N_13587,N_13609);
xnor U13964 (N_13964,N_13607,N_13784);
or U13965 (N_13965,N_13576,N_13593);
xor U13966 (N_13966,N_13731,N_13693);
and U13967 (N_13967,N_13533,N_13512);
xor U13968 (N_13968,N_13653,N_13631);
nand U13969 (N_13969,N_13698,N_13781);
nor U13970 (N_13970,N_13552,N_13658);
nor U13971 (N_13971,N_13794,N_13738);
xor U13972 (N_13972,N_13553,N_13659);
and U13973 (N_13973,N_13555,N_13704);
nor U13974 (N_13974,N_13603,N_13682);
and U13975 (N_13975,N_13635,N_13733);
xnor U13976 (N_13976,N_13573,N_13793);
or U13977 (N_13977,N_13709,N_13517);
nand U13978 (N_13978,N_13717,N_13536);
or U13979 (N_13979,N_13593,N_13670);
and U13980 (N_13980,N_13621,N_13553);
or U13981 (N_13981,N_13766,N_13638);
nand U13982 (N_13982,N_13723,N_13587);
or U13983 (N_13983,N_13630,N_13738);
nor U13984 (N_13984,N_13684,N_13612);
and U13985 (N_13985,N_13638,N_13589);
nor U13986 (N_13986,N_13631,N_13652);
and U13987 (N_13987,N_13519,N_13551);
or U13988 (N_13988,N_13714,N_13698);
xnor U13989 (N_13989,N_13721,N_13517);
and U13990 (N_13990,N_13606,N_13513);
nand U13991 (N_13991,N_13526,N_13716);
nor U13992 (N_13992,N_13588,N_13577);
xnor U13993 (N_13993,N_13595,N_13710);
and U13994 (N_13994,N_13704,N_13655);
nor U13995 (N_13995,N_13672,N_13543);
nand U13996 (N_13996,N_13613,N_13784);
nor U13997 (N_13997,N_13721,N_13574);
or U13998 (N_13998,N_13689,N_13614);
nand U13999 (N_13999,N_13656,N_13590);
or U14000 (N_14000,N_13799,N_13576);
or U14001 (N_14001,N_13640,N_13660);
or U14002 (N_14002,N_13737,N_13685);
xor U14003 (N_14003,N_13616,N_13775);
nor U14004 (N_14004,N_13734,N_13560);
xor U14005 (N_14005,N_13799,N_13534);
nand U14006 (N_14006,N_13540,N_13521);
and U14007 (N_14007,N_13772,N_13749);
or U14008 (N_14008,N_13727,N_13593);
nand U14009 (N_14009,N_13783,N_13773);
nor U14010 (N_14010,N_13755,N_13658);
xor U14011 (N_14011,N_13771,N_13733);
nor U14012 (N_14012,N_13744,N_13558);
or U14013 (N_14013,N_13775,N_13517);
nor U14014 (N_14014,N_13655,N_13611);
nor U14015 (N_14015,N_13739,N_13503);
nor U14016 (N_14016,N_13760,N_13580);
and U14017 (N_14017,N_13727,N_13764);
nand U14018 (N_14018,N_13776,N_13730);
or U14019 (N_14019,N_13736,N_13735);
and U14020 (N_14020,N_13708,N_13565);
nor U14021 (N_14021,N_13699,N_13718);
nor U14022 (N_14022,N_13710,N_13659);
and U14023 (N_14023,N_13740,N_13722);
xnor U14024 (N_14024,N_13534,N_13728);
nor U14025 (N_14025,N_13525,N_13790);
nor U14026 (N_14026,N_13620,N_13510);
nand U14027 (N_14027,N_13623,N_13573);
and U14028 (N_14028,N_13505,N_13756);
or U14029 (N_14029,N_13504,N_13585);
nand U14030 (N_14030,N_13768,N_13534);
and U14031 (N_14031,N_13507,N_13787);
xnor U14032 (N_14032,N_13552,N_13614);
or U14033 (N_14033,N_13622,N_13510);
or U14034 (N_14034,N_13748,N_13787);
nor U14035 (N_14035,N_13533,N_13544);
xor U14036 (N_14036,N_13761,N_13520);
and U14037 (N_14037,N_13586,N_13594);
nor U14038 (N_14038,N_13649,N_13683);
nand U14039 (N_14039,N_13653,N_13537);
xnor U14040 (N_14040,N_13669,N_13599);
nor U14041 (N_14041,N_13577,N_13604);
nand U14042 (N_14042,N_13720,N_13766);
or U14043 (N_14043,N_13726,N_13580);
nand U14044 (N_14044,N_13721,N_13615);
nor U14045 (N_14045,N_13704,N_13551);
or U14046 (N_14046,N_13586,N_13596);
and U14047 (N_14047,N_13615,N_13730);
and U14048 (N_14048,N_13734,N_13752);
xor U14049 (N_14049,N_13615,N_13631);
xnor U14050 (N_14050,N_13710,N_13739);
and U14051 (N_14051,N_13653,N_13740);
nor U14052 (N_14052,N_13557,N_13629);
nor U14053 (N_14053,N_13733,N_13688);
or U14054 (N_14054,N_13749,N_13549);
or U14055 (N_14055,N_13506,N_13514);
or U14056 (N_14056,N_13663,N_13648);
nand U14057 (N_14057,N_13567,N_13672);
xnor U14058 (N_14058,N_13791,N_13502);
or U14059 (N_14059,N_13793,N_13790);
or U14060 (N_14060,N_13609,N_13748);
or U14061 (N_14061,N_13508,N_13717);
xnor U14062 (N_14062,N_13535,N_13581);
xor U14063 (N_14063,N_13765,N_13656);
nor U14064 (N_14064,N_13774,N_13640);
nand U14065 (N_14065,N_13621,N_13683);
nand U14066 (N_14066,N_13553,N_13629);
nand U14067 (N_14067,N_13720,N_13693);
and U14068 (N_14068,N_13614,N_13747);
nand U14069 (N_14069,N_13621,N_13543);
nor U14070 (N_14070,N_13688,N_13552);
or U14071 (N_14071,N_13797,N_13761);
or U14072 (N_14072,N_13563,N_13609);
and U14073 (N_14073,N_13600,N_13655);
and U14074 (N_14074,N_13744,N_13576);
nand U14075 (N_14075,N_13692,N_13641);
and U14076 (N_14076,N_13639,N_13791);
or U14077 (N_14077,N_13522,N_13717);
nor U14078 (N_14078,N_13734,N_13783);
or U14079 (N_14079,N_13746,N_13795);
xnor U14080 (N_14080,N_13569,N_13516);
xnor U14081 (N_14081,N_13739,N_13571);
xor U14082 (N_14082,N_13580,N_13754);
xnor U14083 (N_14083,N_13509,N_13608);
nand U14084 (N_14084,N_13701,N_13552);
nand U14085 (N_14085,N_13678,N_13572);
or U14086 (N_14086,N_13643,N_13517);
nor U14087 (N_14087,N_13566,N_13578);
and U14088 (N_14088,N_13789,N_13655);
or U14089 (N_14089,N_13592,N_13719);
and U14090 (N_14090,N_13561,N_13786);
or U14091 (N_14091,N_13713,N_13613);
nor U14092 (N_14092,N_13598,N_13671);
nor U14093 (N_14093,N_13793,N_13690);
and U14094 (N_14094,N_13528,N_13706);
xnor U14095 (N_14095,N_13592,N_13549);
xor U14096 (N_14096,N_13731,N_13625);
and U14097 (N_14097,N_13662,N_13710);
xor U14098 (N_14098,N_13544,N_13768);
nand U14099 (N_14099,N_13641,N_13675);
xnor U14100 (N_14100,N_13991,N_13936);
xnor U14101 (N_14101,N_14020,N_13962);
nand U14102 (N_14102,N_13801,N_13860);
or U14103 (N_14103,N_13859,N_13820);
nand U14104 (N_14104,N_14029,N_14076);
nand U14105 (N_14105,N_13893,N_13949);
and U14106 (N_14106,N_13881,N_13823);
or U14107 (N_14107,N_13954,N_14062);
nor U14108 (N_14108,N_14084,N_14060);
nand U14109 (N_14109,N_13910,N_14061);
xnor U14110 (N_14110,N_14093,N_13919);
nand U14111 (N_14111,N_13886,N_13869);
nand U14112 (N_14112,N_13916,N_13953);
and U14113 (N_14113,N_13846,N_14000);
xor U14114 (N_14114,N_14053,N_13883);
nor U14115 (N_14115,N_14049,N_13840);
or U14116 (N_14116,N_13818,N_13926);
and U14117 (N_14117,N_13826,N_13845);
and U14118 (N_14118,N_13987,N_14044);
and U14119 (N_14119,N_13838,N_13969);
nor U14120 (N_14120,N_13872,N_14006);
or U14121 (N_14121,N_13849,N_14099);
xor U14122 (N_14122,N_13973,N_13951);
nor U14123 (N_14123,N_13810,N_13937);
nor U14124 (N_14124,N_13829,N_14041);
and U14125 (N_14125,N_13842,N_14040);
xor U14126 (N_14126,N_14046,N_13929);
nor U14127 (N_14127,N_13993,N_13855);
nor U14128 (N_14128,N_13986,N_13992);
nor U14129 (N_14129,N_14032,N_13806);
nand U14130 (N_14130,N_13912,N_14086);
nand U14131 (N_14131,N_14072,N_13945);
xor U14132 (N_14132,N_14048,N_13894);
nand U14133 (N_14133,N_13964,N_13915);
or U14134 (N_14134,N_13958,N_14083);
and U14135 (N_14135,N_14024,N_13983);
nor U14136 (N_14136,N_13808,N_13807);
or U14137 (N_14137,N_13999,N_14003);
or U14138 (N_14138,N_14092,N_13815);
or U14139 (N_14139,N_13866,N_13988);
and U14140 (N_14140,N_13946,N_14097);
or U14141 (N_14141,N_13914,N_13952);
nor U14142 (N_14142,N_14052,N_13997);
nand U14143 (N_14143,N_13880,N_14069);
nand U14144 (N_14144,N_14002,N_14026);
nand U14145 (N_14145,N_13856,N_13963);
nand U14146 (N_14146,N_14057,N_13800);
nand U14147 (N_14147,N_14047,N_13994);
nand U14148 (N_14148,N_14085,N_13904);
xor U14149 (N_14149,N_13955,N_13871);
xor U14150 (N_14150,N_13874,N_13802);
xor U14151 (N_14151,N_13911,N_13972);
xnor U14152 (N_14152,N_13876,N_14038);
or U14153 (N_14153,N_14095,N_14028);
xor U14154 (N_14154,N_13947,N_13821);
nand U14155 (N_14155,N_13966,N_14001);
or U14156 (N_14156,N_14054,N_14096);
and U14157 (N_14157,N_13903,N_14017);
and U14158 (N_14158,N_13899,N_13998);
nor U14159 (N_14159,N_13822,N_13933);
xor U14160 (N_14160,N_13882,N_14005);
nand U14161 (N_14161,N_14025,N_13907);
or U14162 (N_14162,N_13948,N_13878);
nand U14163 (N_14163,N_14063,N_14070);
or U14164 (N_14164,N_14066,N_13943);
nor U14165 (N_14165,N_13819,N_14014);
or U14166 (N_14166,N_13934,N_13835);
nor U14167 (N_14167,N_14012,N_13978);
and U14168 (N_14168,N_13853,N_13956);
xor U14169 (N_14169,N_13844,N_14064);
xnor U14170 (N_14170,N_14015,N_14090);
and U14171 (N_14171,N_14058,N_13901);
or U14172 (N_14172,N_13909,N_13982);
and U14173 (N_14173,N_13913,N_13864);
nand U14174 (N_14174,N_14027,N_13977);
nor U14175 (N_14175,N_13809,N_14088);
nor U14176 (N_14176,N_14087,N_13885);
nor U14177 (N_14177,N_14075,N_13989);
nor U14178 (N_14178,N_14078,N_13925);
nand U14179 (N_14179,N_14091,N_13839);
xor U14180 (N_14180,N_14094,N_13879);
nor U14181 (N_14181,N_13967,N_13961);
or U14182 (N_14182,N_13873,N_13990);
xnor U14183 (N_14183,N_13892,N_14050);
xor U14184 (N_14184,N_14008,N_13939);
xor U14185 (N_14185,N_13862,N_13980);
nor U14186 (N_14186,N_14013,N_13870);
nor U14187 (N_14187,N_13922,N_13889);
xnor U14188 (N_14188,N_14059,N_13817);
xor U14189 (N_14189,N_13906,N_14071);
or U14190 (N_14190,N_13924,N_13935);
nor U14191 (N_14191,N_14089,N_13971);
nand U14192 (N_14192,N_13902,N_13861);
nor U14193 (N_14193,N_14010,N_13804);
nand U14194 (N_14194,N_13996,N_14004);
and U14195 (N_14195,N_14022,N_13985);
and U14196 (N_14196,N_13831,N_13975);
nor U14197 (N_14197,N_14098,N_13965);
and U14198 (N_14198,N_13865,N_14081);
nand U14199 (N_14199,N_13841,N_13921);
nor U14200 (N_14200,N_14051,N_13928);
nand U14201 (N_14201,N_13931,N_13984);
and U14202 (N_14202,N_13938,N_14042);
nand U14203 (N_14203,N_14080,N_13968);
xnor U14204 (N_14204,N_14019,N_13898);
nor U14205 (N_14205,N_14016,N_13863);
nand U14206 (N_14206,N_13868,N_13854);
xnor U14207 (N_14207,N_14067,N_13976);
xnor U14208 (N_14208,N_14045,N_13888);
and U14209 (N_14209,N_13867,N_14018);
xnor U14210 (N_14210,N_13837,N_13917);
nand U14211 (N_14211,N_13814,N_13850);
xor U14212 (N_14212,N_13828,N_14021);
and U14213 (N_14213,N_13852,N_14055);
and U14214 (N_14214,N_13995,N_13896);
nand U14215 (N_14215,N_13825,N_13930);
or U14216 (N_14216,N_14030,N_13858);
or U14217 (N_14217,N_13805,N_13900);
and U14218 (N_14218,N_13918,N_13942);
xnor U14219 (N_14219,N_13957,N_13891);
and U14220 (N_14220,N_13960,N_13847);
nor U14221 (N_14221,N_13836,N_13824);
nor U14222 (N_14222,N_14009,N_13884);
nand U14223 (N_14223,N_14074,N_14034);
xor U14224 (N_14224,N_13897,N_13908);
or U14225 (N_14225,N_13923,N_13927);
xnor U14226 (N_14226,N_13944,N_13890);
or U14227 (N_14227,N_14056,N_13981);
nor U14228 (N_14228,N_14068,N_14082);
or U14229 (N_14229,N_13857,N_13848);
or U14230 (N_14230,N_14035,N_14073);
and U14231 (N_14231,N_13950,N_13877);
and U14232 (N_14232,N_14007,N_14037);
or U14233 (N_14233,N_13827,N_13803);
nor U14234 (N_14234,N_13812,N_14065);
nor U14235 (N_14235,N_13970,N_13830);
xor U14236 (N_14236,N_14077,N_13851);
xor U14237 (N_14237,N_14031,N_13875);
or U14238 (N_14238,N_13941,N_13895);
nand U14239 (N_14239,N_14043,N_14023);
and U14240 (N_14240,N_13887,N_13932);
nor U14241 (N_14241,N_13832,N_13905);
and U14242 (N_14242,N_14033,N_13940);
nand U14243 (N_14243,N_14011,N_13979);
and U14244 (N_14244,N_13811,N_13833);
nand U14245 (N_14245,N_13816,N_13843);
nor U14246 (N_14246,N_14039,N_13813);
xnor U14247 (N_14247,N_13834,N_13920);
nand U14248 (N_14248,N_13959,N_14079);
nand U14249 (N_14249,N_13974,N_14036);
xnor U14250 (N_14250,N_13933,N_14045);
xor U14251 (N_14251,N_13979,N_14081);
xnor U14252 (N_14252,N_13852,N_14067);
xnor U14253 (N_14253,N_14070,N_13880);
nor U14254 (N_14254,N_14043,N_13880);
nand U14255 (N_14255,N_13904,N_14024);
and U14256 (N_14256,N_13866,N_14026);
nand U14257 (N_14257,N_14020,N_14083);
nand U14258 (N_14258,N_14018,N_13894);
xnor U14259 (N_14259,N_14035,N_13949);
xnor U14260 (N_14260,N_14027,N_13957);
nor U14261 (N_14261,N_14062,N_13902);
nor U14262 (N_14262,N_14017,N_13957);
xor U14263 (N_14263,N_14022,N_14065);
or U14264 (N_14264,N_13972,N_14042);
xnor U14265 (N_14265,N_13974,N_13840);
nand U14266 (N_14266,N_13942,N_13971);
nand U14267 (N_14267,N_14019,N_14044);
and U14268 (N_14268,N_13824,N_13914);
nand U14269 (N_14269,N_14084,N_13967);
xor U14270 (N_14270,N_13863,N_13894);
nand U14271 (N_14271,N_14048,N_14009);
or U14272 (N_14272,N_13955,N_14080);
nand U14273 (N_14273,N_14033,N_14028);
xor U14274 (N_14274,N_14047,N_13913);
nor U14275 (N_14275,N_14082,N_13809);
and U14276 (N_14276,N_13934,N_13829);
nand U14277 (N_14277,N_13940,N_13805);
or U14278 (N_14278,N_13920,N_13971);
or U14279 (N_14279,N_13853,N_13883);
nand U14280 (N_14280,N_13997,N_14049);
nor U14281 (N_14281,N_13964,N_13803);
xor U14282 (N_14282,N_14067,N_13906);
and U14283 (N_14283,N_13925,N_14015);
or U14284 (N_14284,N_14011,N_13984);
and U14285 (N_14285,N_13891,N_13936);
or U14286 (N_14286,N_13876,N_13804);
or U14287 (N_14287,N_13974,N_13893);
xor U14288 (N_14288,N_13850,N_13985);
xor U14289 (N_14289,N_14083,N_13889);
and U14290 (N_14290,N_13814,N_13887);
or U14291 (N_14291,N_13922,N_13958);
and U14292 (N_14292,N_13906,N_13827);
or U14293 (N_14293,N_14053,N_13917);
nor U14294 (N_14294,N_14022,N_14060);
xnor U14295 (N_14295,N_14017,N_14039);
or U14296 (N_14296,N_14003,N_13888);
xnor U14297 (N_14297,N_13999,N_13934);
and U14298 (N_14298,N_13956,N_13965);
nand U14299 (N_14299,N_14006,N_14021);
xor U14300 (N_14300,N_13816,N_13859);
and U14301 (N_14301,N_13923,N_13989);
or U14302 (N_14302,N_13911,N_14032);
nand U14303 (N_14303,N_13977,N_13937);
xor U14304 (N_14304,N_13945,N_13946);
xor U14305 (N_14305,N_13804,N_13991);
or U14306 (N_14306,N_14087,N_13868);
and U14307 (N_14307,N_13953,N_13982);
xor U14308 (N_14308,N_14068,N_14022);
or U14309 (N_14309,N_14016,N_14063);
nand U14310 (N_14310,N_13802,N_13867);
nor U14311 (N_14311,N_13911,N_14004);
nor U14312 (N_14312,N_13870,N_13955);
nor U14313 (N_14313,N_13973,N_13959);
or U14314 (N_14314,N_13911,N_13956);
and U14315 (N_14315,N_13961,N_13807);
xor U14316 (N_14316,N_13973,N_13820);
xnor U14317 (N_14317,N_14034,N_14095);
or U14318 (N_14318,N_13956,N_14040);
nor U14319 (N_14319,N_13883,N_13919);
or U14320 (N_14320,N_13861,N_14096);
nor U14321 (N_14321,N_14077,N_13852);
or U14322 (N_14322,N_13812,N_13920);
xor U14323 (N_14323,N_14009,N_13949);
or U14324 (N_14324,N_13825,N_14016);
xor U14325 (N_14325,N_14010,N_13881);
or U14326 (N_14326,N_13915,N_13978);
nor U14327 (N_14327,N_13888,N_14052);
or U14328 (N_14328,N_14067,N_14039);
and U14329 (N_14329,N_13800,N_13814);
and U14330 (N_14330,N_14073,N_13870);
xor U14331 (N_14331,N_13973,N_14094);
nor U14332 (N_14332,N_13836,N_13850);
nor U14333 (N_14333,N_13810,N_13872);
and U14334 (N_14334,N_13951,N_14061);
or U14335 (N_14335,N_14035,N_13804);
nor U14336 (N_14336,N_13818,N_14013);
nand U14337 (N_14337,N_14048,N_13924);
xor U14338 (N_14338,N_13903,N_14000);
and U14339 (N_14339,N_13891,N_13805);
nor U14340 (N_14340,N_14026,N_13872);
xnor U14341 (N_14341,N_14044,N_13946);
and U14342 (N_14342,N_14018,N_13980);
and U14343 (N_14343,N_13896,N_14019);
xor U14344 (N_14344,N_14064,N_14001);
nand U14345 (N_14345,N_13846,N_14049);
or U14346 (N_14346,N_14091,N_13984);
xor U14347 (N_14347,N_14065,N_13865);
nand U14348 (N_14348,N_13811,N_13810);
or U14349 (N_14349,N_13960,N_13908);
or U14350 (N_14350,N_13934,N_13961);
or U14351 (N_14351,N_13951,N_13946);
xor U14352 (N_14352,N_14033,N_13907);
nand U14353 (N_14353,N_13836,N_14066);
nand U14354 (N_14354,N_14006,N_13888);
and U14355 (N_14355,N_13830,N_13925);
xnor U14356 (N_14356,N_14096,N_14022);
xnor U14357 (N_14357,N_14076,N_14001);
nor U14358 (N_14358,N_13869,N_13966);
or U14359 (N_14359,N_14056,N_13912);
xor U14360 (N_14360,N_13803,N_13885);
or U14361 (N_14361,N_13881,N_13811);
or U14362 (N_14362,N_13828,N_13908);
or U14363 (N_14363,N_14091,N_13953);
and U14364 (N_14364,N_14058,N_14085);
and U14365 (N_14365,N_14018,N_13897);
nand U14366 (N_14366,N_13838,N_13896);
nand U14367 (N_14367,N_13905,N_13857);
xor U14368 (N_14368,N_13943,N_13824);
nand U14369 (N_14369,N_13937,N_13813);
and U14370 (N_14370,N_14040,N_13979);
or U14371 (N_14371,N_13811,N_14090);
or U14372 (N_14372,N_13950,N_14012);
and U14373 (N_14373,N_13909,N_13942);
nor U14374 (N_14374,N_14027,N_14016);
and U14375 (N_14375,N_13840,N_14025);
or U14376 (N_14376,N_13832,N_14008);
and U14377 (N_14377,N_13932,N_13916);
nand U14378 (N_14378,N_13863,N_13856);
or U14379 (N_14379,N_13849,N_13940);
nor U14380 (N_14380,N_14080,N_13823);
xnor U14381 (N_14381,N_13962,N_14089);
nor U14382 (N_14382,N_14065,N_13982);
nor U14383 (N_14383,N_13978,N_14082);
or U14384 (N_14384,N_14048,N_13931);
and U14385 (N_14385,N_13989,N_14085);
or U14386 (N_14386,N_13979,N_13801);
nand U14387 (N_14387,N_13960,N_13993);
xor U14388 (N_14388,N_13918,N_14082);
nor U14389 (N_14389,N_13968,N_14072);
or U14390 (N_14390,N_14059,N_13810);
xnor U14391 (N_14391,N_14032,N_14019);
nand U14392 (N_14392,N_14052,N_14026);
nor U14393 (N_14393,N_14057,N_13815);
xnor U14394 (N_14394,N_14084,N_13878);
xor U14395 (N_14395,N_13828,N_13974);
xnor U14396 (N_14396,N_14045,N_14086);
nand U14397 (N_14397,N_13926,N_13905);
xor U14398 (N_14398,N_13859,N_13956);
nand U14399 (N_14399,N_13936,N_13931);
or U14400 (N_14400,N_14321,N_14129);
xnor U14401 (N_14401,N_14396,N_14273);
nand U14402 (N_14402,N_14278,N_14209);
or U14403 (N_14403,N_14234,N_14322);
and U14404 (N_14404,N_14242,N_14153);
nand U14405 (N_14405,N_14225,N_14120);
nand U14406 (N_14406,N_14115,N_14187);
xor U14407 (N_14407,N_14305,N_14260);
xor U14408 (N_14408,N_14372,N_14375);
xor U14409 (N_14409,N_14335,N_14292);
and U14410 (N_14410,N_14371,N_14175);
or U14411 (N_14411,N_14337,N_14384);
nand U14412 (N_14412,N_14320,N_14295);
xor U14413 (N_14413,N_14154,N_14307);
or U14414 (N_14414,N_14394,N_14301);
nor U14415 (N_14415,N_14171,N_14395);
nand U14416 (N_14416,N_14147,N_14308);
nand U14417 (N_14417,N_14298,N_14205);
nand U14418 (N_14418,N_14208,N_14282);
and U14419 (N_14419,N_14252,N_14228);
nor U14420 (N_14420,N_14102,N_14286);
nand U14421 (N_14421,N_14233,N_14219);
xor U14422 (N_14422,N_14347,N_14204);
and U14423 (N_14423,N_14101,N_14151);
xnor U14424 (N_14424,N_14336,N_14266);
nor U14425 (N_14425,N_14203,N_14217);
xnor U14426 (N_14426,N_14330,N_14210);
xor U14427 (N_14427,N_14181,N_14196);
or U14428 (N_14428,N_14363,N_14393);
and U14429 (N_14429,N_14170,N_14274);
xnor U14430 (N_14430,N_14141,N_14190);
nor U14431 (N_14431,N_14133,N_14345);
nor U14432 (N_14432,N_14327,N_14328);
xnor U14433 (N_14433,N_14213,N_14119);
nand U14434 (N_14434,N_14155,N_14388);
or U14435 (N_14435,N_14382,N_14379);
or U14436 (N_14436,N_14332,N_14279);
xnor U14437 (N_14437,N_14265,N_14366);
nand U14438 (N_14438,N_14331,N_14104);
and U14439 (N_14439,N_14106,N_14240);
and U14440 (N_14440,N_14317,N_14387);
nor U14441 (N_14441,N_14362,N_14270);
xor U14442 (N_14442,N_14296,N_14177);
xnor U14443 (N_14443,N_14199,N_14244);
xor U14444 (N_14444,N_14168,N_14235);
nor U14445 (N_14445,N_14340,N_14229);
xor U14446 (N_14446,N_14289,N_14367);
nand U14447 (N_14447,N_14140,N_14276);
or U14448 (N_14448,N_14113,N_14223);
or U14449 (N_14449,N_14294,N_14360);
xnor U14450 (N_14450,N_14125,N_14248);
xnor U14451 (N_14451,N_14373,N_14356);
nor U14452 (N_14452,N_14221,N_14185);
nand U14453 (N_14453,N_14231,N_14202);
nand U14454 (N_14454,N_14156,N_14145);
xnor U14455 (N_14455,N_14198,N_14355);
nor U14456 (N_14456,N_14297,N_14112);
and U14457 (N_14457,N_14211,N_14136);
and U14458 (N_14458,N_14287,N_14293);
or U14459 (N_14459,N_14267,N_14315);
nand U14460 (N_14460,N_14348,N_14251);
xnor U14461 (N_14461,N_14368,N_14126);
xnor U14462 (N_14462,N_14281,N_14299);
or U14463 (N_14463,N_14342,N_14232);
xnor U14464 (N_14464,N_14364,N_14132);
and U14465 (N_14465,N_14280,N_14316);
or U14466 (N_14466,N_14338,N_14121);
xnor U14467 (N_14467,N_14300,N_14116);
or U14468 (N_14468,N_14161,N_14146);
and U14469 (N_14469,N_14117,N_14285);
nor U14470 (N_14470,N_14344,N_14257);
nor U14471 (N_14471,N_14169,N_14165);
xor U14472 (N_14472,N_14263,N_14374);
nor U14473 (N_14473,N_14166,N_14172);
nor U14474 (N_14474,N_14207,N_14230);
nand U14475 (N_14475,N_14167,N_14152);
nor U14476 (N_14476,N_14107,N_14139);
and U14477 (N_14477,N_14343,N_14313);
nand U14478 (N_14478,N_14160,N_14188);
and U14479 (N_14479,N_14222,N_14191);
xnor U14480 (N_14480,N_14100,N_14163);
and U14481 (N_14481,N_14365,N_14186);
or U14482 (N_14482,N_14318,N_14159);
nor U14483 (N_14483,N_14310,N_14246);
and U14484 (N_14484,N_14179,N_14227);
or U14485 (N_14485,N_14253,N_14245);
and U14486 (N_14486,N_14150,N_14114);
nand U14487 (N_14487,N_14135,N_14250);
or U14488 (N_14488,N_14369,N_14137);
or U14489 (N_14489,N_14224,N_14323);
xnor U14490 (N_14490,N_14324,N_14398);
and U14491 (N_14491,N_14241,N_14123);
xnor U14492 (N_14492,N_14383,N_14206);
nor U14493 (N_14493,N_14226,N_14130);
and U14494 (N_14494,N_14329,N_14128);
xnor U14495 (N_14495,N_14385,N_14268);
nor U14496 (N_14496,N_14359,N_14214);
and U14497 (N_14497,N_14258,N_14264);
nand U14498 (N_14498,N_14108,N_14131);
xor U14499 (N_14499,N_14390,N_14326);
or U14500 (N_14500,N_14184,N_14124);
xor U14501 (N_14501,N_14256,N_14197);
xnor U14502 (N_14502,N_14148,N_14358);
nand U14503 (N_14503,N_14122,N_14290);
nand U14504 (N_14504,N_14110,N_14239);
xnor U14505 (N_14505,N_14157,N_14397);
nor U14506 (N_14506,N_14283,N_14312);
xor U14507 (N_14507,N_14192,N_14311);
and U14508 (N_14508,N_14386,N_14237);
nor U14509 (N_14509,N_14339,N_14194);
nor U14510 (N_14510,N_14346,N_14218);
or U14511 (N_14511,N_14334,N_14118);
nor U14512 (N_14512,N_14333,N_14183);
and U14513 (N_14513,N_14220,N_14353);
nand U14514 (N_14514,N_14288,N_14351);
and U14515 (N_14515,N_14275,N_14189);
nand U14516 (N_14516,N_14349,N_14303);
xor U14517 (N_14517,N_14105,N_14378);
nor U14518 (N_14518,N_14291,N_14103);
or U14519 (N_14519,N_14255,N_14361);
nand U14520 (N_14520,N_14238,N_14284);
nand U14521 (N_14521,N_14142,N_14277);
nand U14522 (N_14522,N_14261,N_14243);
and U14523 (N_14523,N_14182,N_14164);
nor U14524 (N_14524,N_14352,N_14306);
xor U14525 (N_14525,N_14109,N_14381);
or U14526 (N_14526,N_14271,N_14269);
nor U14527 (N_14527,N_14138,N_14134);
or U14528 (N_14528,N_14309,N_14180);
or U14529 (N_14529,N_14357,N_14389);
and U14530 (N_14530,N_14247,N_14236);
and U14531 (N_14531,N_14215,N_14127);
nand U14532 (N_14532,N_14376,N_14319);
xnor U14533 (N_14533,N_14149,N_14201);
xor U14534 (N_14534,N_14178,N_14314);
and U14535 (N_14535,N_14304,N_14262);
and U14536 (N_14536,N_14249,N_14212);
xor U14537 (N_14537,N_14143,N_14302);
nor U14538 (N_14538,N_14195,N_14216);
xnor U14539 (N_14539,N_14370,N_14377);
or U14540 (N_14540,N_14325,N_14158);
or U14541 (N_14541,N_14272,N_14162);
xor U14542 (N_14542,N_14176,N_14354);
or U14543 (N_14543,N_14399,N_14200);
or U14544 (N_14544,N_14254,N_14341);
xor U14545 (N_14545,N_14111,N_14174);
nor U14546 (N_14546,N_14380,N_14193);
or U14547 (N_14547,N_14350,N_14259);
nand U14548 (N_14548,N_14392,N_14391);
and U14549 (N_14549,N_14173,N_14144);
nand U14550 (N_14550,N_14245,N_14133);
and U14551 (N_14551,N_14106,N_14251);
nand U14552 (N_14552,N_14106,N_14333);
xnor U14553 (N_14553,N_14362,N_14259);
or U14554 (N_14554,N_14236,N_14164);
and U14555 (N_14555,N_14275,N_14397);
nor U14556 (N_14556,N_14292,N_14252);
nand U14557 (N_14557,N_14366,N_14216);
xnor U14558 (N_14558,N_14282,N_14358);
xnor U14559 (N_14559,N_14331,N_14119);
nor U14560 (N_14560,N_14392,N_14323);
or U14561 (N_14561,N_14390,N_14360);
and U14562 (N_14562,N_14330,N_14347);
nor U14563 (N_14563,N_14299,N_14397);
nand U14564 (N_14564,N_14123,N_14112);
nand U14565 (N_14565,N_14226,N_14302);
xnor U14566 (N_14566,N_14198,N_14177);
nand U14567 (N_14567,N_14135,N_14144);
or U14568 (N_14568,N_14238,N_14301);
or U14569 (N_14569,N_14174,N_14107);
or U14570 (N_14570,N_14206,N_14248);
and U14571 (N_14571,N_14101,N_14265);
or U14572 (N_14572,N_14308,N_14393);
and U14573 (N_14573,N_14140,N_14261);
and U14574 (N_14574,N_14266,N_14254);
and U14575 (N_14575,N_14108,N_14191);
or U14576 (N_14576,N_14294,N_14266);
and U14577 (N_14577,N_14388,N_14242);
xnor U14578 (N_14578,N_14256,N_14181);
and U14579 (N_14579,N_14149,N_14219);
xor U14580 (N_14580,N_14190,N_14148);
and U14581 (N_14581,N_14191,N_14337);
nand U14582 (N_14582,N_14393,N_14206);
and U14583 (N_14583,N_14163,N_14155);
or U14584 (N_14584,N_14331,N_14181);
and U14585 (N_14585,N_14185,N_14182);
nor U14586 (N_14586,N_14253,N_14291);
nand U14587 (N_14587,N_14166,N_14117);
and U14588 (N_14588,N_14133,N_14328);
or U14589 (N_14589,N_14157,N_14311);
nor U14590 (N_14590,N_14395,N_14311);
nor U14591 (N_14591,N_14298,N_14101);
nor U14592 (N_14592,N_14241,N_14331);
xnor U14593 (N_14593,N_14266,N_14233);
or U14594 (N_14594,N_14282,N_14243);
xor U14595 (N_14595,N_14286,N_14355);
nor U14596 (N_14596,N_14333,N_14250);
or U14597 (N_14597,N_14123,N_14166);
nand U14598 (N_14598,N_14341,N_14375);
or U14599 (N_14599,N_14143,N_14132);
or U14600 (N_14600,N_14132,N_14346);
or U14601 (N_14601,N_14240,N_14366);
or U14602 (N_14602,N_14322,N_14379);
or U14603 (N_14603,N_14179,N_14316);
nor U14604 (N_14604,N_14315,N_14277);
and U14605 (N_14605,N_14110,N_14215);
or U14606 (N_14606,N_14265,N_14123);
nor U14607 (N_14607,N_14309,N_14307);
nand U14608 (N_14608,N_14214,N_14114);
xnor U14609 (N_14609,N_14280,N_14108);
xnor U14610 (N_14610,N_14153,N_14305);
xnor U14611 (N_14611,N_14268,N_14187);
nand U14612 (N_14612,N_14228,N_14197);
nand U14613 (N_14613,N_14186,N_14319);
and U14614 (N_14614,N_14348,N_14387);
nor U14615 (N_14615,N_14236,N_14153);
xnor U14616 (N_14616,N_14180,N_14386);
nor U14617 (N_14617,N_14158,N_14310);
or U14618 (N_14618,N_14248,N_14258);
or U14619 (N_14619,N_14346,N_14237);
nand U14620 (N_14620,N_14247,N_14397);
or U14621 (N_14621,N_14336,N_14208);
xor U14622 (N_14622,N_14295,N_14147);
or U14623 (N_14623,N_14335,N_14144);
or U14624 (N_14624,N_14383,N_14238);
or U14625 (N_14625,N_14213,N_14357);
or U14626 (N_14626,N_14379,N_14151);
xnor U14627 (N_14627,N_14384,N_14339);
xnor U14628 (N_14628,N_14192,N_14211);
or U14629 (N_14629,N_14113,N_14263);
xor U14630 (N_14630,N_14266,N_14102);
nor U14631 (N_14631,N_14224,N_14350);
xnor U14632 (N_14632,N_14261,N_14238);
nor U14633 (N_14633,N_14304,N_14139);
nand U14634 (N_14634,N_14323,N_14123);
xor U14635 (N_14635,N_14257,N_14119);
xor U14636 (N_14636,N_14203,N_14334);
nand U14637 (N_14637,N_14191,N_14129);
xnor U14638 (N_14638,N_14179,N_14231);
xor U14639 (N_14639,N_14188,N_14303);
and U14640 (N_14640,N_14267,N_14113);
or U14641 (N_14641,N_14230,N_14312);
and U14642 (N_14642,N_14181,N_14253);
nand U14643 (N_14643,N_14137,N_14278);
and U14644 (N_14644,N_14204,N_14274);
or U14645 (N_14645,N_14144,N_14236);
nand U14646 (N_14646,N_14310,N_14186);
or U14647 (N_14647,N_14316,N_14360);
or U14648 (N_14648,N_14266,N_14166);
nand U14649 (N_14649,N_14351,N_14125);
nand U14650 (N_14650,N_14227,N_14218);
xor U14651 (N_14651,N_14288,N_14114);
and U14652 (N_14652,N_14260,N_14252);
and U14653 (N_14653,N_14115,N_14199);
xor U14654 (N_14654,N_14205,N_14227);
and U14655 (N_14655,N_14253,N_14377);
nor U14656 (N_14656,N_14265,N_14357);
xnor U14657 (N_14657,N_14253,N_14236);
and U14658 (N_14658,N_14348,N_14276);
and U14659 (N_14659,N_14104,N_14207);
xor U14660 (N_14660,N_14259,N_14280);
xor U14661 (N_14661,N_14262,N_14300);
xor U14662 (N_14662,N_14283,N_14202);
and U14663 (N_14663,N_14149,N_14228);
and U14664 (N_14664,N_14179,N_14124);
and U14665 (N_14665,N_14349,N_14235);
nand U14666 (N_14666,N_14216,N_14318);
nor U14667 (N_14667,N_14384,N_14312);
nor U14668 (N_14668,N_14250,N_14387);
and U14669 (N_14669,N_14375,N_14271);
nand U14670 (N_14670,N_14219,N_14354);
and U14671 (N_14671,N_14238,N_14283);
nand U14672 (N_14672,N_14197,N_14276);
or U14673 (N_14673,N_14266,N_14385);
or U14674 (N_14674,N_14134,N_14137);
or U14675 (N_14675,N_14152,N_14397);
nand U14676 (N_14676,N_14175,N_14149);
nor U14677 (N_14677,N_14276,N_14258);
nor U14678 (N_14678,N_14286,N_14235);
nand U14679 (N_14679,N_14170,N_14396);
xnor U14680 (N_14680,N_14336,N_14163);
and U14681 (N_14681,N_14103,N_14355);
nor U14682 (N_14682,N_14277,N_14242);
xor U14683 (N_14683,N_14385,N_14348);
or U14684 (N_14684,N_14282,N_14372);
or U14685 (N_14685,N_14393,N_14333);
nor U14686 (N_14686,N_14193,N_14138);
xor U14687 (N_14687,N_14329,N_14280);
nor U14688 (N_14688,N_14260,N_14234);
xor U14689 (N_14689,N_14120,N_14179);
xnor U14690 (N_14690,N_14312,N_14363);
or U14691 (N_14691,N_14278,N_14396);
or U14692 (N_14692,N_14159,N_14176);
xor U14693 (N_14693,N_14178,N_14395);
and U14694 (N_14694,N_14354,N_14389);
or U14695 (N_14695,N_14318,N_14373);
and U14696 (N_14696,N_14206,N_14236);
and U14697 (N_14697,N_14194,N_14159);
nor U14698 (N_14698,N_14197,N_14223);
and U14699 (N_14699,N_14203,N_14166);
or U14700 (N_14700,N_14401,N_14543);
xor U14701 (N_14701,N_14672,N_14520);
and U14702 (N_14702,N_14587,N_14421);
nand U14703 (N_14703,N_14552,N_14661);
nor U14704 (N_14704,N_14585,N_14618);
and U14705 (N_14705,N_14446,N_14603);
and U14706 (N_14706,N_14505,N_14696);
xor U14707 (N_14707,N_14665,N_14464);
and U14708 (N_14708,N_14581,N_14481);
nor U14709 (N_14709,N_14572,N_14644);
nand U14710 (N_14710,N_14594,N_14676);
nand U14711 (N_14711,N_14402,N_14638);
and U14712 (N_14712,N_14438,N_14443);
or U14713 (N_14713,N_14441,N_14525);
nand U14714 (N_14714,N_14573,N_14569);
nor U14715 (N_14715,N_14452,N_14433);
nand U14716 (N_14716,N_14560,N_14537);
nand U14717 (N_14717,N_14612,N_14629);
nor U14718 (N_14718,N_14406,N_14664);
and U14719 (N_14719,N_14440,N_14496);
and U14720 (N_14720,N_14574,N_14506);
nor U14721 (N_14721,N_14508,N_14545);
and U14722 (N_14722,N_14654,N_14474);
nand U14723 (N_14723,N_14436,N_14691);
or U14724 (N_14724,N_14586,N_14655);
nor U14725 (N_14725,N_14453,N_14686);
nor U14726 (N_14726,N_14681,N_14634);
or U14727 (N_14727,N_14487,N_14549);
and U14728 (N_14728,N_14529,N_14411);
nand U14729 (N_14729,N_14559,N_14582);
and U14730 (N_14730,N_14454,N_14404);
xor U14731 (N_14731,N_14652,N_14610);
or U14732 (N_14732,N_14486,N_14554);
nand U14733 (N_14733,N_14504,N_14413);
nor U14734 (N_14734,N_14418,N_14456);
nand U14735 (N_14735,N_14533,N_14432);
and U14736 (N_14736,N_14512,N_14689);
nand U14737 (N_14737,N_14547,N_14579);
or U14738 (N_14738,N_14675,N_14470);
nor U14739 (N_14739,N_14499,N_14492);
xor U14740 (N_14740,N_14476,N_14528);
nor U14741 (N_14741,N_14518,N_14658);
and U14742 (N_14742,N_14494,N_14480);
xnor U14743 (N_14743,N_14576,N_14534);
or U14744 (N_14744,N_14444,N_14601);
or U14745 (N_14745,N_14604,N_14422);
and U14746 (N_14746,N_14619,N_14426);
xnor U14747 (N_14747,N_14465,N_14489);
nor U14748 (N_14748,N_14437,N_14683);
or U14749 (N_14749,N_14690,N_14613);
or U14750 (N_14750,N_14427,N_14469);
xnor U14751 (N_14751,N_14632,N_14620);
or U14752 (N_14752,N_14420,N_14478);
xor U14753 (N_14753,N_14449,N_14414);
or U14754 (N_14754,N_14530,N_14460);
nand U14755 (N_14755,N_14684,N_14692);
nand U14756 (N_14756,N_14685,N_14498);
nand U14757 (N_14757,N_14516,N_14532);
or U14758 (N_14758,N_14631,N_14615);
and U14759 (N_14759,N_14561,N_14477);
nand U14760 (N_14760,N_14577,N_14571);
xnor U14761 (N_14761,N_14442,N_14542);
or U14762 (N_14762,N_14531,N_14588);
and U14763 (N_14763,N_14502,N_14641);
xnor U14764 (N_14764,N_14431,N_14558);
nor U14765 (N_14765,N_14417,N_14666);
or U14766 (N_14766,N_14595,N_14483);
xor U14767 (N_14767,N_14546,N_14584);
or U14768 (N_14768,N_14600,N_14607);
nand U14769 (N_14769,N_14415,N_14482);
nor U14770 (N_14770,N_14566,N_14628);
xnor U14771 (N_14771,N_14682,N_14621);
or U14772 (N_14772,N_14503,N_14524);
or U14773 (N_14773,N_14510,N_14539);
xnor U14774 (N_14774,N_14650,N_14695);
or U14775 (N_14775,N_14567,N_14556);
and U14776 (N_14776,N_14425,N_14562);
xor U14777 (N_14777,N_14403,N_14495);
nor U14778 (N_14778,N_14564,N_14687);
nor U14779 (N_14779,N_14697,N_14541);
or U14780 (N_14780,N_14630,N_14522);
or U14781 (N_14781,N_14535,N_14428);
and U14782 (N_14782,N_14694,N_14647);
nor U14783 (N_14783,N_14674,N_14670);
and U14784 (N_14784,N_14511,N_14471);
nor U14785 (N_14785,N_14430,N_14490);
xnor U14786 (N_14786,N_14626,N_14445);
and U14787 (N_14787,N_14678,N_14563);
and U14788 (N_14788,N_14636,N_14536);
and U14789 (N_14789,N_14459,N_14521);
and U14790 (N_14790,N_14515,N_14698);
and U14791 (N_14791,N_14640,N_14590);
nand U14792 (N_14792,N_14497,N_14458);
and U14793 (N_14793,N_14693,N_14578);
nand U14794 (N_14794,N_14592,N_14448);
or U14795 (N_14795,N_14596,N_14468);
nand U14796 (N_14796,N_14523,N_14625);
or U14797 (N_14797,N_14667,N_14527);
xnor U14798 (N_14798,N_14659,N_14648);
xnor U14799 (N_14799,N_14699,N_14643);
nor U14800 (N_14800,N_14540,N_14423);
and U14801 (N_14801,N_14624,N_14407);
or U14802 (N_14802,N_14606,N_14416);
or U14803 (N_14803,N_14656,N_14660);
xor U14804 (N_14804,N_14410,N_14688);
and U14805 (N_14805,N_14509,N_14472);
nor U14806 (N_14806,N_14663,N_14617);
nand U14807 (N_14807,N_14405,N_14461);
xnor U14808 (N_14808,N_14517,N_14668);
or U14809 (N_14809,N_14642,N_14565);
and U14810 (N_14810,N_14639,N_14623);
or U14811 (N_14811,N_14673,N_14580);
xor U14812 (N_14812,N_14519,N_14645);
and U14813 (N_14813,N_14570,N_14679);
nor U14814 (N_14814,N_14627,N_14611);
nand U14815 (N_14815,N_14671,N_14575);
and U14816 (N_14816,N_14553,N_14500);
nand U14817 (N_14817,N_14466,N_14488);
and U14818 (N_14818,N_14616,N_14457);
nor U14819 (N_14819,N_14637,N_14653);
or U14820 (N_14820,N_14646,N_14633);
or U14821 (N_14821,N_14635,N_14669);
and U14822 (N_14822,N_14408,N_14491);
nand U14823 (N_14823,N_14614,N_14593);
and U14824 (N_14824,N_14591,N_14485);
nand U14825 (N_14825,N_14484,N_14493);
and U14826 (N_14826,N_14429,N_14450);
or U14827 (N_14827,N_14568,N_14662);
xnor U14828 (N_14828,N_14501,N_14434);
and U14829 (N_14829,N_14447,N_14473);
xor U14830 (N_14830,N_14555,N_14424);
and U14831 (N_14831,N_14439,N_14557);
nand U14832 (N_14832,N_14538,N_14677);
xnor U14833 (N_14833,N_14589,N_14548);
xor U14834 (N_14834,N_14455,N_14680);
xnor U14835 (N_14835,N_14657,N_14598);
nor U14836 (N_14836,N_14514,N_14599);
nor U14837 (N_14837,N_14609,N_14479);
xnor U14838 (N_14838,N_14435,N_14649);
or U14839 (N_14839,N_14463,N_14507);
nand U14840 (N_14840,N_14475,N_14451);
xnor U14841 (N_14841,N_14412,N_14622);
xor U14842 (N_14842,N_14462,N_14550);
and U14843 (N_14843,N_14544,N_14409);
nor U14844 (N_14844,N_14551,N_14526);
and U14845 (N_14845,N_14400,N_14513);
xnor U14846 (N_14846,N_14651,N_14602);
nand U14847 (N_14847,N_14597,N_14605);
nand U14848 (N_14848,N_14583,N_14608);
or U14849 (N_14849,N_14419,N_14467);
or U14850 (N_14850,N_14573,N_14663);
or U14851 (N_14851,N_14425,N_14592);
nand U14852 (N_14852,N_14447,N_14405);
xor U14853 (N_14853,N_14561,N_14486);
nand U14854 (N_14854,N_14499,N_14577);
xnor U14855 (N_14855,N_14614,N_14568);
xnor U14856 (N_14856,N_14541,N_14404);
nand U14857 (N_14857,N_14686,N_14484);
and U14858 (N_14858,N_14431,N_14596);
nor U14859 (N_14859,N_14546,N_14635);
and U14860 (N_14860,N_14500,N_14677);
or U14861 (N_14861,N_14698,N_14572);
or U14862 (N_14862,N_14413,N_14662);
xnor U14863 (N_14863,N_14648,N_14491);
nor U14864 (N_14864,N_14554,N_14404);
or U14865 (N_14865,N_14594,N_14433);
and U14866 (N_14866,N_14557,N_14618);
xnor U14867 (N_14867,N_14651,N_14492);
nor U14868 (N_14868,N_14598,N_14653);
and U14869 (N_14869,N_14445,N_14467);
nand U14870 (N_14870,N_14670,N_14690);
nand U14871 (N_14871,N_14569,N_14428);
and U14872 (N_14872,N_14507,N_14542);
and U14873 (N_14873,N_14510,N_14416);
or U14874 (N_14874,N_14682,N_14556);
xnor U14875 (N_14875,N_14447,N_14692);
xor U14876 (N_14876,N_14674,N_14667);
and U14877 (N_14877,N_14479,N_14662);
and U14878 (N_14878,N_14482,N_14554);
and U14879 (N_14879,N_14594,N_14563);
nor U14880 (N_14880,N_14580,N_14667);
xor U14881 (N_14881,N_14663,N_14541);
and U14882 (N_14882,N_14497,N_14507);
and U14883 (N_14883,N_14594,N_14665);
and U14884 (N_14884,N_14660,N_14478);
or U14885 (N_14885,N_14615,N_14543);
nor U14886 (N_14886,N_14526,N_14644);
nor U14887 (N_14887,N_14574,N_14697);
xnor U14888 (N_14888,N_14462,N_14609);
nor U14889 (N_14889,N_14411,N_14455);
xnor U14890 (N_14890,N_14582,N_14677);
and U14891 (N_14891,N_14693,N_14423);
xor U14892 (N_14892,N_14407,N_14444);
nor U14893 (N_14893,N_14584,N_14623);
or U14894 (N_14894,N_14406,N_14656);
nand U14895 (N_14895,N_14580,N_14475);
xnor U14896 (N_14896,N_14408,N_14483);
or U14897 (N_14897,N_14537,N_14443);
xor U14898 (N_14898,N_14693,N_14518);
and U14899 (N_14899,N_14433,N_14412);
nor U14900 (N_14900,N_14577,N_14470);
and U14901 (N_14901,N_14508,N_14460);
nand U14902 (N_14902,N_14433,N_14517);
xnor U14903 (N_14903,N_14493,N_14430);
nor U14904 (N_14904,N_14428,N_14418);
or U14905 (N_14905,N_14500,N_14422);
or U14906 (N_14906,N_14436,N_14611);
nand U14907 (N_14907,N_14611,N_14507);
nor U14908 (N_14908,N_14593,N_14620);
and U14909 (N_14909,N_14578,N_14698);
nor U14910 (N_14910,N_14421,N_14622);
nand U14911 (N_14911,N_14469,N_14548);
or U14912 (N_14912,N_14686,N_14692);
and U14913 (N_14913,N_14571,N_14439);
or U14914 (N_14914,N_14521,N_14579);
nand U14915 (N_14915,N_14417,N_14640);
xor U14916 (N_14916,N_14641,N_14550);
nand U14917 (N_14917,N_14514,N_14447);
xnor U14918 (N_14918,N_14534,N_14545);
and U14919 (N_14919,N_14594,N_14480);
and U14920 (N_14920,N_14638,N_14543);
nor U14921 (N_14921,N_14582,N_14667);
nor U14922 (N_14922,N_14410,N_14697);
xnor U14923 (N_14923,N_14603,N_14636);
and U14924 (N_14924,N_14548,N_14543);
nand U14925 (N_14925,N_14573,N_14612);
and U14926 (N_14926,N_14429,N_14536);
nand U14927 (N_14927,N_14560,N_14491);
and U14928 (N_14928,N_14599,N_14586);
or U14929 (N_14929,N_14693,N_14555);
nand U14930 (N_14930,N_14654,N_14505);
nand U14931 (N_14931,N_14572,N_14442);
nand U14932 (N_14932,N_14426,N_14403);
xor U14933 (N_14933,N_14454,N_14444);
or U14934 (N_14934,N_14578,N_14569);
nor U14935 (N_14935,N_14486,N_14645);
nand U14936 (N_14936,N_14508,N_14433);
or U14937 (N_14937,N_14691,N_14470);
xnor U14938 (N_14938,N_14482,N_14583);
and U14939 (N_14939,N_14613,N_14616);
nor U14940 (N_14940,N_14695,N_14544);
or U14941 (N_14941,N_14457,N_14424);
or U14942 (N_14942,N_14446,N_14520);
or U14943 (N_14943,N_14696,N_14411);
xor U14944 (N_14944,N_14400,N_14451);
nand U14945 (N_14945,N_14501,N_14545);
and U14946 (N_14946,N_14456,N_14682);
and U14947 (N_14947,N_14406,N_14500);
nand U14948 (N_14948,N_14469,N_14461);
or U14949 (N_14949,N_14571,N_14419);
and U14950 (N_14950,N_14506,N_14480);
and U14951 (N_14951,N_14661,N_14534);
xor U14952 (N_14952,N_14440,N_14471);
nor U14953 (N_14953,N_14463,N_14423);
or U14954 (N_14954,N_14652,N_14544);
nor U14955 (N_14955,N_14588,N_14500);
nor U14956 (N_14956,N_14660,N_14488);
or U14957 (N_14957,N_14568,N_14466);
xor U14958 (N_14958,N_14637,N_14568);
nor U14959 (N_14959,N_14467,N_14556);
nor U14960 (N_14960,N_14553,N_14654);
nand U14961 (N_14961,N_14541,N_14591);
nor U14962 (N_14962,N_14435,N_14487);
and U14963 (N_14963,N_14679,N_14469);
or U14964 (N_14964,N_14616,N_14566);
and U14965 (N_14965,N_14414,N_14555);
or U14966 (N_14966,N_14675,N_14666);
and U14967 (N_14967,N_14666,N_14460);
xor U14968 (N_14968,N_14598,N_14507);
nand U14969 (N_14969,N_14430,N_14457);
nor U14970 (N_14970,N_14696,N_14694);
nor U14971 (N_14971,N_14614,N_14554);
nor U14972 (N_14972,N_14496,N_14604);
xnor U14973 (N_14973,N_14473,N_14555);
nor U14974 (N_14974,N_14480,N_14584);
and U14975 (N_14975,N_14447,N_14456);
nor U14976 (N_14976,N_14635,N_14499);
xnor U14977 (N_14977,N_14630,N_14510);
nor U14978 (N_14978,N_14403,N_14458);
nor U14979 (N_14979,N_14499,N_14474);
or U14980 (N_14980,N_14612,N_14518);
nand U14981 (N_14981,N_14643,N_14497);
nand U14982 (N_14982,N_14547,N_14616);
and U14983 (N_14983,N_14460,N_14558);
nor U14984 (N_14984,N_14470,N_14674);
and U14985 (N_14985,N_14666,N_14663);
nor U14986 (N_14986,N_14444,N_14590);
nand U14987 (N_14987,N_14648,N_14443);
xnor U14988 (N_14988,N_14577,N_14536);
and U14989 (N_14989,N_14582,N_14496);
and U14990 (N_14990,N_14473,N_14649);
or U14991 (N_14991,N_14683,N_14673);
or U14992 (N_14992,N_14620,N_14679);
xor U14993 (N_14993,N_14414,N_14525);
and U14994 (N_14994,N_14611,N_14654);
and U14995 (N_14995,N_14587,N_14612);
nor U14996 (N_14996,N_14627,N_14401);
nor U14997 (N_14997,N_14421,N_14605);
xor U14998 (N_14998,N_14572,N_14605);
and U14999 (N_14999,N_14493,N_14667);
or U15000 (N_15000,N_14996,N_14817);
nor U15001 (N_15001,N_14871,N_14720);
nand U15002 (N_15002,N_14910,N_14751);
xor U15003 (N_15003,N_14744,N_14734);
nor U15004 (N_15004,N_14754,N_14867);
or U15005 (N_15005,N_14998,N_14761);
and U15006 (N_15006,N_14798,N_14799);
nand U15007 (N_15007,N_14913,N_14932);
xor U15008 (N_15008,N_14718,N_14764);
nand U15009 (N_15009,N_14872,N_14947);
xor U15010 (N_15010,N_14784,N_14729);
or U15011 (N_15011,N_14879,N_14722);
and U15012 (N_15012,N_14735,N_14836);
or U15013 (N_15013,N_14916,N_14738);
xor U15014 (N_15014,N_14939,N_14736);
nor U15015 (N_15015,N_14746,N_14762);
xor U15016 (N_15016,N_14948,N_14753);
and U15017 (N_15017,N_14815,N_14887);
nand U15018 (N_15018,N_14975,N_14908);
xor U15019 (N_15019,N_14968,N_14859);
nor U15020 (N_15020,N_14919,N_14864);
and U15021 (N_15021,N_14776,N_14701);
or U15022 (N_15022,N_14758,N_14844);
nor U15023 (N_15023,N_14726,N_14828);
xor U15024 (N_15024,N_14770,N_14896);
or U15025 (N_15025,N_14955,N_14849);
nand U15026 (N_15026,N_14774,N_14834);
xor U15027 (N_15027,N_14742,N_14991);
or U15028 (N_15028,N_14831,N_14856);
or U15029 (N_15029,N_14760,N_14780);
nor U15030 (N_15030,N_14768,N_14940);
nand U15031 (N_15031,N_14731,N_14778);
nand U15032 (N_15032,N_14902,N_14728);
and U15033 (N_15033,N_14763,N_14714);
nand U15034 (N_15034,N_14988,N_14709);
xor U15035 (N_15035,N_14737,N_14878);
and U15036 (N_15036,N_14961,N_14886);
and U15037 (N_15037,N_14857,N_14851);
xor U15038 (N_15038,N_14806,N_14813);
nor U15039 (N_15039,N_14953,N_14786);
xor U15040 (N_15040,N_14860,N_14765);
xor U15041 (N_15041,N_14712,N_14927);
xor U15042 (N_15042,N_14824,N_14790);
xor U15043 (N_15043,N_14981,N_14755);
or U15044 (N_15044,N_14873,N_14829);
or U15045 (N_15045,N_14924,N_14854);
or U15046 (N_15046,N_14861,N_14715);
nor U15047 (N_15047,N_14875,N_14915);
or U15048 (N_15048,N_14952,N_14766);
nor U15049 (N_15049,N_14819,N_14997);
nand U15050 (N_15050,N_14822,N_14992);
and U15051 (N_15051,N_14787,N_14852);
xor U15052 (N_15052,N_14983,N_14750);
xnor U15053 (N_15053,N_14733,N_14892);
and U15054 (N_15054,N_14876,N_14959);
and U15055 (N_15055,N_14779,N_14757);
nor U15056 (N_15056,N_14781,N_14707);
xor U15057 (N_15057,N_14724,N_14802);
nand U15058 (N_15058,N_14835,N_14727);
or U15059 (N_15059,N_14805,N_14882);
and U15060 (N_15060,N_14803,N_14783);
and U15061 (N_15061,N_14772,N_14796);
xor U15062 (N_15062,N_14777,N_14956);
or U15063 (N_15063,N_14708,N_14972);
nor U15064 (N_15064,N_14946,N_14999);
xnor U15065 (N_15065,N_14848,N_14889);
xnor U15066 (N_15066,N_14740,N_14967);
or U15067 (N_15067,N_14745,N_14801);
and U15068 (N_15068,N_14880,N_14909);
nand U15069 (N_15069,N_14903,N_14853);
nand U15070 (N_15070,N_14782,N_14730);
nand U15071 (N_15071,N_14769,N_14989);
xnor U15072 (N_15072,N_14840,N_14905);
and U15073 (N_15073,N_14984,N_14929);
and U15074 (N_15074,N_14870,N_14716);
xnor U15075 (N_15075,N_14756,N_14969);
nand U15076 (N_15076,N_14973,N_14914);
and U15077 (N_15077,N_14904,N_14721);
xnor U15078 (N_15078,N_14850,N_14960);
xnor U15079 (N_15079,N_14890,N_14845);
or U15080 (N_15080,N_14966,N_14926);
or U15081 (N_15081,N_14943,N_14936);
or U15082 (N_15082,N_14931,N_14881);
xnor U15083 (N_15083,N_14884,N_14888);
and U15084 (N_15084,N_14855,N_14771);
nand U15085 (N_15085,N_14814,N_14944);
nor U15086 (N_15086,N_14862,N_14797);
and U15087 (N_15087,N_14812,N_14723);
or U15088 (N_15088,N_14832,N_14901);
or U15089 (N_15089,N_14893,N_14816);
and U15090 (N_15090,N_14789,N_14962);
nand U15091 (N_15091,N_14842,N_14739);
nor U15092 (N_15092,N_14917,N_14963);
nor U15093 (N_15093,N_14868,N_14704);
and U15094 (N_15094,N_14841,N_14964);
nand U15095 (N_15095,N_14976,N_14820);
nand U15096 (N_15096,N_14930,N_14847);
xor U15097 (N_15097,N_14928,N_14748);
xor U15098 (N_15098,N_14874,N_14711);
nor U15099 (N_15099,N_14818,N_14885);
or U15100 (N_15100,N_14970,N_14839);
nand U15101 (N_15101,N_14826,N_14749);
or U15102 (N_15102,N_14994,N_14920);
nor U15103 (N_15103,N_14858,N_14794);
or U15104 (N_15104,N_14922,N_14958);
and U15105 (N_15105,N_14921,N_14971);
xnor U15106 (N_15106,N_14775,N_14894);
nand U15107 (N_15107,N_14865,N_14907);
and U15108 (N_15108,N_14937,N_14950);
or U15109 (N_15109,N_14793,N_14705);
nand U15110 (N_15110,N_14838,N_14900);
or U15111 (N_15111,N_14978,N_14911);
xnor U15112 (N_15112,N_14743,N_14942);
nand U15113 (N_15113,N_14897,N_14759);
nand U15114 (N_15114,N_14846,N_14895);
xnor U15115 (N_15115,N_14767,N_14833);
xnor U15116 (N_15116,N_14933,N_14837);
and U15117 (N_15117,N_14823,N_14883);
nand U15118 (N_15118,N_14843,N_14791);
xnor U15119 (N_15119,N_14700,N_14891);
nor U15120 (N_15120,N_14987,N_14993);
xnor U15121 (N_15121,N_14732,N_14788);
nand U15122 (N_15122,N_14703,N_14785);
xnor U15123 (N_15123,N_14923,N_14741);
and U15124 (N_15124,N_14811,N_14935);
or U15125 (N_15125,N_14710,N_14980);
or U15126 (N_15126,N_14830,N_14906);
xor U15127 (N_15127,N_14934,N_14706);
nand U15128 (N_15128,N_14957,N_14899);
or U15129 (N_15129,N_14713,N_14747);
nor U15130 (N_15130,N_14800,N_14949);
nor U15131 (N_15131,N_14965,N_14717);
nand U15132 (N_15132,N_14804,N_14941);
nand U15133 (N_15133,N_14945,N_14809);
xor U15134 (N_15134,N_14827,N_14810);
or U15135 (N_15135,N_14985,N_14808);
and U15136 (N_15136,N_14877,N_14821);
or U15137 (N_15137,N_14938,N_14912);
and U15138 (N_15138,N_14954,N_14979);
nand U15139 (N_15139,N_14773,N_14807);
or U15140 (N_15140,N_14995,N_14792);
xor U15141 (N_15141,N_14898,N_14795);
nand U15142 (N_15142,N_14825,N_14719);
nand U15143 (N_15143,N_14752,N_14863);
nand U15144 (N_15144,N_14866,N_14974);
nor U15145 (N_15145,N_14725,N_14925);
and U15146 (N_15146,N_14702,N_14982);
or U15147 (N_15147,N_14977,N_14869);
and U15148 (N_15148,N_14986,N_14918);
xor U15149 (N_15149,N_14951,N_14990);
nand U15150 (N_15150,N_14803,N_14915);
and U15151 (N_15151,N_14842,N_14716);
and U15152 (N_15152,N_14973,N_14803);
xor U15153 (N_15153,N_14753,N_14985);
or U15154 (N_15154,N_14908,N_14830);
or U15155 (N_15155,N_14834,N_14844);
xor U15156 (N_15156,N_14993,N_14738);
xor U15157 (N_15157,N_14771,N_14709);
xor U15158 (N_15158,N_14938,N_14773);
nor U15159 (N_15159,N_14849,N_14857);
or U15160 (N_15160,N_14994,N_14911);
xor U15161 (N_15161,N_14743,N_14870);
xor U15162 (N_15162,N_14718,N_14754);
nor U15163 (N_15163,N_14829,N_14897);
xor U15164 (N_15164,N_14891,N_14898);
nor U15165 (N_15165,N_14878,N_14923);
xnor U15166 (N_15166,N_14757,N_14727);
nor U15167 (N_15167,N_14900,N_14711);
nor U15168 (N_15168,N_14876,N_14990);
xnor U15169 (N_15169,N_14942,N_14953);
and U15170 (N_15170,N_14874,N_14954);
and U15171 (N_15171,N_14816,N_14922);
and U15172 (N_15172,N_14978,N_14831);
nor U15173 (N_15173,N_14702,N_14827);
nand U15174 (N_15174,N_14849,N_14967);
nand U15175 (N_15175,N_14762,N_14818);
nand U15176 (N_15176,N_14780,N_14959);
nand U15177 (N_15177,N_14998,N_14736);
nand U15178 (N_15178,N_14883,N_14972);
xor U15179 (N_15179,N_14919,N_14946);
and U15180 (N_15180,N_14904,N_14704);
or U15181 (N_15181,N_14877,N_14999);
and U15182 (N_15182,N_14742,N_14856);
and U15183 (N_15183,N_14865,N_14835);
or U15184 (N_15184,N_14948,N_14872);
nor U15185 (N_15185,N_14711,N_14708);
or U15186 (N_15186,N_14858,N_14773);
nand U15187 (N_15187,N_14881,N_14755);
nor U15188 (N_15188,N_14858,N_14733);
xor U15189 (N_15189,N_14937,N_14834);
and U15190 (N_15190,N_14806,N_14907);
or U15191 (N_15191,N_14713,N_14841);
nor U15192 (N_15192,N_14774,N_14854);
or U15193 (N_15193,N_14760,N_14982);
or U15194 (N_15194,N_14980,N_14828);
xnor U15195 (N_15195,N_14879,N_14714);
nand U15196 (N_15196,N_14885,N_14948);
nand U15197 (N_15197,N_14887,N_14851);
nor U15198 (N_15198,N_14888,N_14873);
and U15199 (N_15199,N_14967,N_14906);
xnor U15200 (N_15200,N_14819,N_14709);
nand U15201 (N_15201,N_14875,N_14834);
nand U15202 (N_15202,N_14701,N_14774);
or U15203 (N_15203,N_14973,N_14784);
nor U15204 (N_15204,N_14715,N_14743);
nand U15205 (N_15205,N_14929,N_14845);
nor U15206 (N_15206,N_14745,N_14946);
nand U15207 (N_15207,N_14719,N_14717);
and U15208 (N_15208,N_14722,N_14976);
nor U15209 (N_15209,N_14988,N_14766);
nor U15210 (N_15210,N_14732,N_14875);
or U15211 (N_15211,N_14988,N_14765);
or U15212 (N_15212,N_14900,N_14725);
xor U15213 (N_15213,N_14745,N_14819);
nor U15214 (N_15214,N_14839,N_14902);
or U15215 (N_15215,N_14925,N_14862);
xor U15216 (N_15216,N_14875,N_14879);
nand U15217 (N_15217,N_14797,N_14972);
nor U15218 (N_15218,N_14876,N_14781);
xor U15219 (N_15219,N_14758,N_14969);
nor U15220 (N_15220,N_14908,N_14902);
and U15221 (N_15221,N_14915,N_14703);
nor U15222 (N_15222,N_14762,N_14873);
and U15223 (N_15223,N_14868,N_14702);
or U15224 (N_15224,N_14987,N_14767);
nand U15225 (N_15225,N_14751,N_14842);
xnor U15226 (N_15226,N_14842,N_14964);
xor U15227 (N_15227,N_14995,N_14999);
nor U15228 (N_15228,N_14825,N_14931);
nand U15229 (N_15229,N_14846,N_14884);
or U15230 (N_15230,N_14701,N_14946);
nor U15231 (N_15231,N_14910,N_14844);
xnor U15232 (N_15232,N_14985,N_14872);
or U15233 (N_15233,N_14993,N_14885);
and U15234 (N_15234,N_14781,N_14989);
or U15235 (N_15235,N_14746,N_14753);
nand U15236 (N_15236,N_14819,N_14951);
nor U15237 (N_15237,N_14721,N_14871);
nand U15238 (N_15238,N_14889,N_14855);
and U15239 (N_15239,N_14753,N_14742);
or U15240 (N_15240,N_14921,N_14861);
xnor U15241 (N_15241,N_14710,N_14867);
and U15242 (N_15242,N_14800,N_14918);
or U15243 (N_15243,N_14881,N_14779);
or U15244 (N_15244,N_14751,N_14797);
xor U15245 (N_15245,N_14916,N_14701);
or U15246 (N_15246,N_14751,N_14961);
or U15247 (N_15247,N_14832,N_14993);
xor U15248 (N_15248,N_14778,N_14994);
or U15249 (N_15249,N_14761,N_14866);
nor U15250 (N_15250,N_14871,N_14855);
nor U15251 (N_15251,N_14937,N_14794);
nor U15252 (N_15252,N_14951,N_14860);
xnor U15253 (N_15253,N_14703,N_14904);
nor U15254 (N_15254,N_14895,N_14999);
nor U15255 (N_15255,N_14866,N_14853);
nand U15256 (N_15256,N_14901,N_14979);
or U15257 (N_15257,N_14716,N_14912);
nand U15258 (N_15258,N_14944,N_14851);
and U15259 (N_15259,N_14782,N_14834);
nand U15260 (N_15260,N_14752,N_14942);
and U15261 (N_15261,N_14818,N_14775);
or U15262 (N_15262,N_14976,N_14886);
nand U15263 (N_15263,N_14979,N_14806);
xor U15264 (N_15264,N_14865,N_14754);
nor U15265 (N_15265,N_14974,N_14944);
or U15266 (N_15266,N_14922,N_14751);
or U15267 (N_15267,N_14834,N_14702);
nand U15268 (N_15268,N_14719,N_14908);
and U15269 (N_15269,N_14987,N_14812);
nor U15270 (N_15270,N_14957,N_14930);
and U15271 (N_15271,N_14969,N_14836);
and U15272 (N_15272,N_14774,N_14930);
or U15273 (N_15273,N_14721,N_14977);
and U15274 (N_15274,N_14739,N_14847);
or U15275 (N_15275,N_14786,N_14764);
xor U15276 (N_15276,N_14792,N_14891);
nor U15277 (N_15277,N_14783,N_14786);
or U15278 (N_15278,N_14834,N_14942);
xnor U15279 (N_15279,N_14928,N_14996);
or U15280 (N_15280,N_14978,N_14841);
and U15281 (N_15281,N_14838,N_14929);
and U15282 (N_15282,N_14714,N_14770);
nand U15283 (N_15283,N_14993,N_14888);
xnor U15284 (N_15284,N_14773,N_14748);
xnor U15285 (N_15285,N_14741,N_14879);
or U15286 (N_15286,N_14771,N_14796);
and U15287 (N_15287,N_14847,N_14959);
or U15288 (N_15288,N_14831,N_14983);
and U15289 (N_15289,N_14930,N_14978);
xor U15290 (N_15290,N_14780,N_14869);
or U15291 (N_15291,N_14877,N_14726);
or U15292 (N_15292,N_14727,N_14813);
nor U15293 (N_15293,N_14851,N_14795);
nor U15294 (N_15294,N_14815,N_14980);
nor U15295 (N_15295,N_14998,N_14808);
or U15296 (N_15296,N_14810,N_14826);
or U15297 (N_15297,N_14812,N_14809);
nand U15298 (N_15298,N_14787,N_14945);
or U15299 (N_15299,N_14912,N_14898);
or U15300 (N_15300,N_15178,N_15236);
nor U15301 (N_15301,N_15261,N_15093);
or U15302 (N_15302,N_15248,N_15255);
and U15303 (N_15303,N_15085,N_15217);
xnor U15304 (N_15304,N_15260,N_15029);
or U15305 (N_15305,N_15100,N_15212);
nand U15306 (N_15306,N_15058,N_15210);
and U15307 (N_15307,N_15017,N_15252);
nor U15308 (N_15308,N_15195,N_15191);
nor U15309 (N_15309,N_15071,N_15069);
nor U15310 (N_15310,N_15298,N_15243);
nand U15311 (N_15311,N_15270,N_15180);
and U15312 (N_15312,N_15202,N_15228);
nand U15313 (N_15313,N_15133,N_15173);
nor U15314 (N_15314,N_15204,N_15274);
or U15315 (N_15315,N_15157,N_15175);
xor U15316 (N_15316,N_15235,N_15049);
nand U15317 (N_15317,N_15283,N_15139);
and U15318 (N_15318,N_15165,N_15281);
xnor U15319 (N_15319,N_15084,N_15155);
nor U15320 (N_15320,N_15192,N_15138);
xor U15321 (N_15321,N_15159,N_15064);
or U15322 (N_15322,N_15036,N_15096);
xnor U15323 (N_15323,N_15123,N_15237);
and U15324 (N_15324,N_15201,N_15014);
and U15325 (N_15325,N_15249,N_15272);
and U15326 (N_15326,N_15023,N_15055);
xor U15327 (N_15327,N_15004,N_15080);
xnor U15328 (N_15328,N_15024,N_15140);
xor U15329 (N_15329,N_15063,N_15122);
and U15330 (N_15330,N_15208,N_15297);
nor U15331 (N_15331,N_15168,N_15259);
and U15332 (N_15332,N_15182,N_15124);
and U15333 (N_15333,N_15184,N_15137);
and U15334 (N_15334,N_15041,N_15246);
and U15335 (N_15335,N_15289,N_15282);
or U15336 (N_15336,N_15188,N_15291);
or U15337 (N_15337,N_15083,N_15089);
nand U15338 (N_15338,N_15244,N_15053);
and U15339 (N_15339,N_15211,N_15117);
xnor U15340 (N_15340,N_15129,N_15194);
or U15341 (N_15341,N_15148,N_15088);
or U15342 (N_15342,N_15003,N_15278);
nand U15343 (N_15343,N_15242,N_15144);
xnor U15344 (N_15344,N_15240,N_15176);
nor U15345 (N_15345,N_15108,N_15189);
xor U15346 (N_15346,N_15146,N_15214);
nand U15347 (N_15347,N_15038,N_15264);
and U15348 (N_15348,N_15154,N_15010);
and U15349 (N_15349,N_15200,N_15054);
or U15350 (N_15350,N_15197,N_15040);
nor U15351 (N_15351,N_15126,N_15187);
nand U15352 (N_15352,N_15193,N_15179);
nor U15353 (N_15353,N_15273,N_15121);
and U15354 (N_15354,N_15229,N_15099);
nand U15355 (N_15355,N_15152,N_15031);
nor U15356 (N_15356,N_15044,N_15062);
or U15357 (N_15357,N_15151,N_15143);
xor U15358 (N_15358,N_15042,N_15112);
nor U15359 (N_15359,N_15156,N_15160);
nand U15360 (N_15360,N_15196,N_15141);
nor U15361 (N_15361,N_15039,N_15056);
or U15362 (N_15362,N_15022,N_15256);
or U15363 (N_15363,N_15276,N_15005);
xnor U15364 (N_15364,N_15111,N_15215);
xor U15365 (N_15365,N_15070,N_15269);
or U15366 (N_15366,N_15043,N_15206);
or U15367 (N_15367,N_15292,N_15057);
and U15368 (N_15368,N_15263,N_15115);
nand U15369 (N_15369,N_15241,N_15199);
or U15370 (N_15370,N_15198,N_15275);
or U15371 (N_15371,N_15268,N_15072);
xor U15372 (N_15372,N_15086,N_15052);
nor U15373 (N_15373,N_15186,N_15142);
nand U15374 (N_15374,N_15149,N_15073);
nand U15375 (N_15375,N_15113,N_15081);
or U15376 (N_15376,N_15098,N_15225);
nor U15377 (N_15377,N_15231,N_15277);
xnor U15378 (N_15378,N_15279,N_15094);
xor U15379 (N_15379,N_15035,N_15163);
nor U15380 (N_15380,N_15245,N_15131);
and U15381 (N_15381,N_15000,N_15147);
nor U15382 (N_15382,N_15128,N_15021);
nor U15383 (N_15383,N_15103,N_15107);
nor U15384 (N_15384,N_15018,N_15266);
nor U15385 (N_15385,N_15234,N_15092);
or U15386 (N_15386,N_15271,N_15284);
nor U15387 (N_15387,N_15183,N_15015);
nor U15388 (N_15388,N_15177,N_15078);
nor U15389 (N_15389,N_15050,N_15068);
nand U15390 (N_15390,N_15087,N_15104);
and U15391 (N_15391,N_15046,N_15207);
and U15392 (N_15392,N_15290,N_15170);
or U15393 (N_15393,N_15221,N_15267);
nor U15394 (N_15394,N_15145,N_15265);
or U15395 (N_15395,N_15065,N_15226);
and U15396 (N_15396,N_15101,N_15153);
nor U15397 (N_15397,N_15213,N_15167);
xor U15398 (N_15398,N_15033,N_15075);
and U15399 (N_15399,N_15219,N_15037);
nor U15400 (N_15400,N_15060,N_15171);
or U15401 (N_15401,N_15016,N_15006);
and U15402 (N_15402,N_15119,N_15090);
or U15403 (N_15403,N_15285,N_15007);
or U15404 (N_15404,N_15251,N_15066);
or U15405 (N_15405,N_15253,N_15220);
and U15406 (N_15406,N_15106,N_15095);
nand U15407 (N_15407,N_15216,N_15002);
xor U15408 (N_15408,N_15091,N_15025);
and U15409 (N_15409,N_15132,N_15059);
or U15410 (N_15410,N_15114,N_15079);
nor U15411 (N_15411,N_15120,N_15295);
or U15412 (N_15412,N_15209,N_15190);
or U15413 (N_15413,N_15028,N_15164);
and U15414 (N_15414,N_15247,N_15116);
xnor U15415 (N_15415,N_15181,N_15230);
and U15416 (N_15416,N_15250,N_15258);
nand U15417 (N_15417,N_15013,N_15222);
nor U15418 (N_15418,N_15118,N_15136);
and U15419 (N_15419,N_15223,N_15218);
nor U15420 (N_15420,N_15232,N_15011);
xor U15421 (N_15421,N_15296,N_15262);
nand U15422 (N_15422,N_15130,N_15001);
nand U15423 (N_15423,N_15082,N_15097);
and U15424 (N_15424,N_15280,N_15047);
nor U15425 (N_15425,N_15224,N_15299);
xor U15426 (N_15426,N_15020,N_15287);
xor U15427 (N_15427,N_15019,N_15161);
xnor U15428 (N_15428,N_15286,N_15125);
or U15429 (N_15429,N_15150,N_15203);
xnor U15430 (N_15430,N_15166,N_15110);
or U15431 (N_15431,N_15032,N_15134);
xnor U15432 (N_15432,N_15238,N_15048);
or U15433 (N_15433,N_15077,N_15067);
nand U15434 (N_15434,N_15027,N_15294);
nand U15435 (N_15435,N_15185,N_15169);
nor U15436 (N_15436,N_15030,N_15174);
or U15437 (N_15437,N_15293,N_15008);
nand U15438 (N_15438,N_15257,N_15102);
xnor U15439 (N_15439,N_15135,N_15009);
xor U15440 (N_15440,N_15172,N_15162);
or U15441 (N_15441,N_15254,N_15127);
and U15442 (N_15442,N_15105,N_15233);
and U15443 (N_15443,N_15061,N_15227);
or U15444 (N_15444,N_15051,N_15158);
xor U15445 (N_15445,N_15012,N_15205);
and U15446 (N_15446,N_15074,N_15045);
or U15447 (N_15447,N_15026,N_15288);
and U15448 (N_15448,N_15076,N_15034);
or U15449 (N_15449,N_15109,N_15239);
and U15450 (N_15450,N_15152,N_15206);
or U15451 (N_15451,N_15257,N_15043);
xnor U15452 (N_15452,N_15296,N_15194);
and U15453 (N_15453,N_15229,N_15244);
xnor U15454 (N_15454,N_15158,N_15152);
and U15455 (N_15455,N_15269,N_15058);
nor U15456 (N_15456,N_15266,N_15030);
or U15457 (N_15457,N_15049,N_15104);
xnor U15458 (N_15458,N_15108,N_15047);
nor U15459 (N_15459,N_15213,N_15214);
and U15460 (N_15460,N_15237,N_15291);
or U15461 (N_15461,N_15057,N_15138);
and U15462 (N_15462,N_15118,N_15014);
nand U15463 (N_15463,N_15145,N_15047);
and U15464 (N_15464,N_15179,N_15108);
xnor U15465 (N_15465,N_15293,N_15192);
nor U15466 (N_15466,N_15226,N_15111);
nand U15467 (N_15467,N_15036,N_15063);
or U15468 (N_15468,N_15156,N_15090);
or U15469 (N_15469,N_15013,N_15069);
and U15470 (N_15470,N_15225,N_15276);
and U15471 (N_15471,N_15208,N_15147);
or U15472 (N_15472,N_15195,N_15222);
xnor U15473 (N_15473,N_15239,N_15287);
nand U15474 (N_15474,N_15052,N_15274);
nand U15475 (N_15475,N_15103,N_15190);
nor U15476 (N_15476,N_15081,N_15133);
nor U15477 (N_15477,N_15293,N_15159);
nand U15478 (N_15478,N_15035,N_15294);
or U15479 (N_15479,N_15101,N_15134);
nor U15480 (N_15480,N_15081,N_15099);
xor U15481 (N_15481,N_15096,N_15105);
or U15482 (N_15482,N_15137,N_15104);
nor U15483 (N_15483,N_15274,N_15266);
or U15484 (N_15484,N_15018,N_15038);
or U15485 (N_15485,N_15104,N_15008);
nand U15486 (N_15486,N_15242,N_15052);
and U15487 (N_15487,N_15266,N_15290);
or U15488 (N_15488,N_15045,N_15267);
nand U15489 (N_15489,N_15091,N_15112);
and U15490 (N_15490,N_15121,N_15275);
and U15491 (N_15491,N_15228,N_15223);
nand U15492 (N_15492,N_15269,N_15215);
or U15493 (N_15493,N_15132,N_15229);
nand U15494 (N_15494,N_15127,N_15048);
and U15495 (N_15495,N_15017,N_15184);
or U15496 (N_15496,N_15057,N_15135);
nor U15497 (N_15497,N_15231,N_15000);
nor U15498 (N_15498,N_15083,N_15055);
nand U15499 (N_15499,N_15027,N_15251);
or U15500 (N_15500,N_15040,N_15298);
and U15501 (N_15501,N_15272,N_15172);
and U15502 (N_15502,N_15089,N_15113);
nand U15503 (N_15503,N_15193,N_15140);
or U15504 (N_15504,N_15298,N_15122);
and U15505 (N_15505,N_15109,N_15102);
and U15506 (N_15506,N_15262,N_15223);
or U15507 (N_15507,N_15053,N_15184);
or U15508 (N_15508,N_15195,N_15298);
nor U15509 (N_15509,N_15107,N_15088);
xor U15510 (N_15510,N_15186,N_15016);
and U15511 (N_15511,N_15051,N_15043);
xnor U15512 (N_15512,N_15186,N_15036);
xor U15513 (N_15513,N_15260,N_15182);
and U15514 (N_15514,N_15100,N_15146);
or U15515 (N_15515,N_15298,N_15100);
nor U15516 (N_15516,N_15049,N_15190);
and U15517 (N_15517,N_15002,N_15093);
or U15518 (N_15518,N_15240,N_15278);
nand U15519 (N_15519,N_15217,N_15155);
or U15520 (N_15520,N_15229,N_15283);
or U15521 (N_15521,N_15106,N_15221);
xor U15522 (N_15522,N_15288,N_15296);
nor U15523 (N_15523,N_15192,N_15003);
nor U15524 (N_15524,N_15053,N_15242);
nor U15525 (N_15525,N_15154,N_15250);
nand U15526 (N_15526,N_15120,N_15078);
or U15527 (N_15527,N_15047,N_15000);
xnor U15528 (N_15528,N_15148,N_15165);
or U15529 (N_15529,N_15140,N_15085);
nor U15530 (N_15530,N_15153,N_15064);
or U15531 (N_15531,N_15162,N_15023);
nand U15532 (N_15532,N_15180,N_15025);
nand U15533 (N_15533,N_15108,N_15130);
and U15534 (N_15534,N_15009,N_15112);
and U15535 (N_15535,N_15163,N_15055);
nor U15536 (N_15536,N_15198,N_15238);
or U15537 (N_15537,N_15130,N_15016);
nor U15538 (N_15538,N_15029,N_15051);
xor U15539 (N_15539,N_15031,N_15032);
nand U15540 (N_15540,N_15110,N_15136);
nand U15541 (N_15541,N_15038,N_15128);
nand U15542 (N_15542,N_15290,N_15124);
xor U15543 (N_15543,N_15183,N_15042);
and U15544 (N_15544,N_15235,N_15217);
xnor U15545 (N_15545,N_15107,N_15032);
xnor U15546 (N_15546,N_15123,N_15170);
nor U15547 (N_15547,N_15228,N_15270);
nand U15548 (N_15548,N_15131,N_15107);
nand U15549 (N_15549,N_15226,N_15268);
or U15550 (N_15550,N_15099,N_15185);
nor U15551 (N_15551,N_15275,N_15288);
nor U15552 (N_15552,N_15249,N_15173);
nand U15553 (N_15553,N_15217,N_15248);
nor U15554 (N_15554,N_15236,N_15148);
or U15555 (N_15555,N_15204,N_15195);
nor U15556 (N_15556,N_15038,N_15120);
nand U15557 (N_15557,N_15014,N_15166);
and U15558 (N_15558,N_15126,N_15052);
and U15559 (N_15559,N_15162,N_15243);
and U15560 (N_15560,N_15207,N_15065);
nor U15561 (N_15561,N_15101,N_15089);
nor U15562 (N_15562,N_15043,N_15139);
nand U15563 (N_15563,N_15044,N_15231);
nand U15564 (N_15564,N_15171,N_15184);
nor U15565 (N_15565,N_15036,N_15085);
nor U15566 (N_15566,N_15160,N_15075);
xnor U15567 (N_15567,N_15026,N_15101);
nor U15568 (N_15568,N_15263,N_15167);
xnor U15569 (N_15569,N_15051,N_15090);
or U15570 (N_15570,N_15203,N_15102);
and U15571 (N_15571,N_15277,N_15284);
nand U15572 (N_15572,N_15275,N_15264);
nor U15573 (N_15573,N_15217,N_15141);
and U15574 (N_15574,N_15287,N_15011);
nor U15575 (N_15575,N_15235,N_15297);
and U15576 (N_15576,N_15211,N_15121);
or U15577 (N_15577,N_15192,N_15134);
or U15578 (N_15578,N_15241,N_15004);
or U15579 (N_15579,N_15143,N_15033);
or U15580 (N_15580,N_15086,N_15266);
and U15581 (N_15581,N_15025,N_15119);
nor U15582 (N_15582,N_15117,N_15286);
nand U15583 (N_15583,N_15112,N_15061);
nand U15584 (N_15584,N_15142,N_15146);
and U15585 (N_15585,N_15273,N_15021);
nor U15586 (N_15586,N_15210,N_15062);
nor U15587 (N_15587,N_15049,N_15240);
xnor U15588 (N_15588,N_15135,N_15213);
and U15589 (N_15589,N_15271,N_15105);
xor U15590 (N_15590,N_15289,N_15042);
or U15591 (N_15591,N_15294,N_15230);
nor U15592 (N_15592,N_15067,N_15217);
and U15593 (N_15593,N_15252,N_15041);
or U15594 (N_15594,N_15191,N_15057);
nand U15595 (N_15595,N_15216,N_15078);
or U15596 (N_15596,N_15194,N_15131);
xnor U15597 (N_15597,N_15151,N_15007);
or U15598 (N_15598,N_15074,N_15237);
nor U15599 (N_15599,N_15244,N_15045);
or U15600 (N_15600,N_15559,N_15357);
nor U15601 (N_15601,N_15430,N_15325);
nor U15602 (N_15602,N_15327,N_15411);
and U15603 (N_15603,N_15393,N_15491);
or U15604 (N_15604,N_15377,N_15317);
nand U15605 (N_15605,N_15319,N_15336);
and U15606 (N_15606,N_15314,N_15520);
nand U15607 (N_15607,N_15570,N_15361);
or U15608 (N_15608,N_15376,N_15577);
nand U15609 (N_15609,N_15534,N_15443);
nand U15610 (N_15610,N_15472,N_15363);
xor U15611 (N_15611,N_15300,N_15490);
nand U15612 (N_15612,N_15392,N_15598);
xnor U15613 (N_15613,N_15349,N_15350);
xnor U15614 (N_15614,N_15425,N_15398);
xor U15615 (N_15615,N_15503,N_15473);
nand U15616 (N_15616,N_15429,N_15501);
or U15617 (N_15617,N_15588,N_15388);
xor U15618 (N_15618,N_15365,N_15590);
and U15619 (N_15619,N_15482,N_15304);
xnor U15620 (N_15620,N_15551,N_15435);
or U15621 (N_15621,N_15511,N_15541);
nor U15622 (N_15622,N_15306,N_15455);
or U15623 (N_15623,N_15535,N_15409);
xor U15624 (N_15624,N_15316,N_15466);
and U15625 (N_15625,N_15468,N_15487);
nor U15626 (N_15626,N_15318,N_15563);
nor U15627 (N_15627,N_15369,N_15475);
nor U15628 (N_15628,N_15460,N_15539);
or U15629 (N_15629,N_15366,N_15574);
or U15630 (N_15630,N_15567,N_15390);
nand U15631 (N_15631,N_15315,N_15510);
or U15632 (N_15632,N_15575,N_15387);
nand U15633 (N_15633,N_15404,N_15421);
nand U15634 (N_15634,N_15334,N_15572);
xnor U15635 (N_15635,N_15498,N_15529);
nand U15636 (N_15636,N_15332,N_15562);
xor U15637 (N_15637,N_15513,N_15348);
xor U15638 (N_15638,N_15444,N_15449);
nor U15639 (N_15639,N_15508,N_15457);
and U15640 (N_15640,N_15335,N_15434);
and U15641 (N_15641,N_15507,N_15586);
nand U15642 (N_15642,N_15424,N_15523);
xor U15643 (N_15643,N_15420,N_15368);
or U15644 (N_15644,N_15599,N_15470);
xor U15645 (N_15645,N_15462,N_15354);
nand U15646 (N_15646,N_15439,N_15389);
nor U15647 (N_15647,N_15545,N_15313);
and U15648 (N_15648,N_15433,N_15403);
and U15649 (N_15649,N_15483,N_15423);
xnor U15650 (N_15650,N_15419,N_15564);
nor U15651 (N_15651,N_15589,N_15308);
nor U15652 (N_15652,N_15395,N_15372);
or U15653 (N_15653,N_15373,N_15383);
and U15654 (N_15654,N_15526,N_15499);
or U15655 (N_15655,N_15587,N_15518);
and U15656 (N_15656,N_15305,N_15394);
nor U15657 (N_15657,N_15346,N_15480);
nor U15658 (N_15658,N_15525,N_15431);
or U15659 (N_15659,N_15543,N_15374);
nand U15660 (N_15660,N_15464,N_15307);
nand U15661 (N_15661,N_15581,N_15320);
nand U15662 (N_15662,N_15597,N_15408);
or U15663 (N_15663,N_15532,N_15322);
and U15664 (N_15664,N_15362,N_15331);
or U15665 (N_15665,N_15445,N_15502);
or U15666 (N_15666,N_15509,N_15522);
or U15667 (N_15667,N_15592,N_15355);
xnor U15668 (N_15668,N_15427,N_15323);
xnor U15669 (N_15669,N_15301,N_15517);
and U15670 (N_15670,N_15370,N_15552);
xnor U15671 (N_15671,N_15358,N_15527);
or U15672 (N_15672,N_15340,N_15407);
nor U15673 (N_15673,N_15359,N_15573);
or U15674 (N_15674,N_15382,N_15437);
or U15675 (N_15675,N_15345,N_15414);
or U15676 (N_15676,N_15413,N_15302);
xnor U15677 (N_15677,N_15494,N_15440);
nor U15678 (N_15678,N_15533,N_15536);
or U15679 (N_15679,N_15337,N_15530);
nand U15680 (N_15680,N_15579,N_15479);
xnor U15681 (N_15681,N_15446,N_15519);
nor U15682 (N_15682,N_15339,N_15546);
and U15683 (N_15683,N_15516,N_15399);
xnor U15684 (N_15684,N_15585,N_15488);
nor U15685 (N_15685,N_15576,N_15338);
or U15686 (N_15686,N_15416,N_15594);
nand U15687 (N_15687,N_15512,N_15593);
or U15688 (N_15688,N_15578,N_15415);
xnor U15689 (N_15689,N_15451,N_15463);
or U15690 (N_15690,N_15310,N_15474);
nor U15691 (N_15691,N_15356,N_15381);
and U15692 (N_15692,N_15344,N_15458);
xor U15693 (N_15693,N_15418,N_15537);
xor U15694 (N_15694,N_15426,N_15412);
and U15695 (N_15695,N_15448,N_15540);
and U15696 (N_15696,N_15422,N_15561);
nand U15697 (N_15697,N_15506,N_15524);
nor U15698 (N_15698,N_15405,N_15486);
nor U15699 (N_15699,N_15595,N_15330);
or U15700 (N_15700,N_15584,N_15556);
nor U15701 (N_15701,N_15496,N_15568);
nand U15702 (N_15702,N_15401,N_15391);
xor U15703 (N_15703,N_15341,N_15542);
and U15704 (N_15704,N_15514,N_15452);
xor U15705 (N_15705,N_15554,N_15569);
or U15706 (N_15706,N_15428,N_15371);
or U15707 (N_15707,N_15493,N_15495);
nand U15708 (N_15708,N_15504,N_15347);
nand U15709 (N_15709,N_15438,N_15565);
or U15710 (N_15710,N_15549,N_15465);
xor U15711 (N_15711,N_15402,N_15453);
nor U15712 (N_15712,N_15571,N_15467);
and U15713 (N_15713,N_15410,N_15515);
xnor U15714 (N_15714,N_15384,N_15459);
nor U15715 (N_15715,N_15353,N_15312);
xnor U15716 (N_15716,N_15521,N_15454);
xnor U15717 (N_15717,N_15471,N_15591);
xor U15718 (N_15718,N_15528,N_15500);
and U15719 (N_15719,N_15324,N_15555);
xnor U15720 (N_15720,N_15580,N_15328);
xor U15721 (N_15721,N_15550,N_15560);
and U15722 (N_15722,N_15478,N_15558);
or U15723 (N_15723,N_15544,N_15477);
xor U15724 (N_15724,N_15385,N_15476);
or U15725 (N_15725,N_15436,N_15333);
nand U15726 (N_15726,N_15342,N_15492);
xnor U15727 (N_15727,N_15484,N_15380);
and U15728 (N_15728,N_15378,N_15469);
and U15729 (N_15729,N_15303,N_15351);
or U15730 (N_15730,N_15343,N_15406);
nand U15731 (N_15731,N_15326,N_15596);
nor U15732 (N_15732,N_15379,N_15538);
or U15733 (N_15733,N_15553,N_15386);
nor U15734 (N_15734,N_15364,N_15505);
nor U15735 (N_15735,N_15583,N_15450);
or U15736 (N_15736,N_15557,N_15447);
or U15737 (N_15737,N_15441,N_15329);
or U15738 (N_15738,N_15547,N_15432);
nand U15739 (N_15739,N_15531,N_15400);
and U15740 (N_15740,N_15396,N_15461);
xor U15741 (N_15741,N_15481,N_15582);
nor U15742 (N_15742,N_15397,N_15566);
nand U15743 (N_15743,N_15321,N_15456);
or U15744 (N_15744,N_15352,N_15311);
nor U15745 (N_15745,N_15442,N_15360);
and U15746 (N_15746,N_15548,N_15417);
nand U15747 (N_15747,N_15497,N_15367);
xnor U15748 (N_15748,N_15485,N_15309);
or U15749 (N_15749,N_15489,N_15375);
or U15750 (N_15750,N_15572,N_15403);
nor U15751 (N_15751,N_15532,N_15354);
nor U15752 (N_15752,N_15461,N_15360);
xnor U15753 (N_15753,N_15583,N_15368);
nor U15754 (N_15754,N_15342,N_15502);
and U15755 (N_15755,N_15373,N_15391);
nand U15756 (N_15756,N_15572,N_15465);
and U15757 (N_15757,N_15338,N_15431);
xnor U15758 (N_15758,N_15386,N_15402);
nor U15759 (N_15759,N_15542,N_15547);
nand U15760 (N_15760,N_15356,N_15376);
and U15761 (N_15761,N_15329,N_15313);
nor U15762 (N_15762,N_15361,N_15439);
xnor U15763 (N_15763,N_15439,N_15486);
and U15764 (N_15764,N_15501,N_15548);
nor U15765 (N_15765,N_15345,N_15560);
nand U15766 (N_15766,N_15436,N_15393);
xor U15767 (N_15767,N_15410,N_15482);
or U15768 (N_15768,N_15301,N_15320);
or U15769 (N_15769,N_15382,N_15306);
nor U15770 (N_15770,N_15378,N_15531);
nor U15771 (N_15771,N_15535,N_15483);
and U15772 (N_15772,N_15491,N_15441);
and U15773 (N_15773,N_15471,N_15334);
and U15774 (N_15774,N_15303,N_15342);
and U15775 (N_15775,N_15595,N_15421);
and U15776 (N_15776,N_15468,N_15443);
nor U15777 (N_15777,N_15340,N_15579);
or U15778 (N_15778,N_15548,N_15317);
or U15779 (N_15779,N_15333,N_15520);
xor U15780 (N_15780,N_15579,N_15416);
or U15781 (N_15781,N_15378,N_15367);
nor U15782 (N_15782,N_15430,N_15451);
or U15783 (N_15783,N_15368,N_15537);
and U15784 (N_15784,N_15569,N_15452);
xnor U15785 (N_15785,N_15489,N_15477);
nor U15786 (N_15786,N_15576,N_15579);
and U15787 (N_15787,N_15300,N_15432);
nor U15788 (N_15788,N_15419,N_15553);
or U15789 (N_15789,N_15469,N_15322);
or U15790 (N_15790,N_15445,N_15326);
or U15791 (N_15791,N_15495,N_15519);
nand U15792 (N_15792,N_15580,N_15406);
xnor U15793 (N_15793,N_15469,N_15548);
or U15794 (N_15794,N_15311,N_15449);
xnor U15795 (N_15795,N_15523,N_15393);
and U15796 (N_15796,N_15374,N_15352);
or U15797 (N_15797,N_15558,N_15590);
and U15798 (N_15798,N_15487,N_15561);
nor U15799 (N_15799,N_15553,N_15562);
nand U15800 (N_15800,N_15407,N_15424);
and U15801 (N_15801,N_15384,N_15403);
nand U15802 (N_15802,N_15364,N_15367);
or U15803 (N_15803,N_15363,N_15348);
or U15804 (N_15804,N_15562,N_15593);
nor U15805 (N_15805,N_15479,N_15310);
nor U15806 (N_15806,N_15592,N_15353);
and U15807 (N_15807,N_15587,N_15464);
or U15808 (N_15808,N_15502,N_15424);
xnor U15809 (N_15809,N_15312,N_15544);
nand U15810 (N_15810,N_15569,N_15326);
and U15811 (N_15811,N_15430,N_15332);
xnor U15812 (N_15812,N_15551,N_15591);
or U15813 (N_15813,N_15537,N_15487);
or U15814 (N_15814,N_15336,N_15422);
nor U15815 (N_15815,N_15557,N_15543);
or U15816 (N_15816,N_15554,N_15480);
and U15817 (N_15817,N_15523,N_15323);
nand U15818 (N_15818,N_15339,N_15421);
xnor U15819 (N_15819,N_15409,N_15568);
nor U15820 (N_15820,N_15432,N_15349);
nand U15821 (N_15821,N_15507,N_15497);
xnor U15822 (N_15822,N_15539,N_15486);
xor U15823 (N_15823,N_15329,N_15507);
nor U15824 (N_15824,N_15371,N_15336);
nor U15825 (N_15825,N_15493,N_15312);
xnor U15826 (N_15826,N_15342,N_15579);
or U15827 (N_15827,N_15422,N_15567);
or U15828 (N_15828,N_15376,N_15556);
xor U15829 (N_15829,N_15512,N_15546);
and U15830 (N_15830,N_15558,N_15556);
xor U15831 (N_15831,N_15425,N_15477);
and U15832 (N_15832,N_15373,N_15490);
xnor U15833 (N_15833,N_15589,N_15544);
or U15834 (N_15834,N_15500,N_15431);
or U15835 (N_15835,N_15345,N_15342);
or U15836 (N_15836,N_15478,N_15403);
nand U15837 (N_15837,N_15401,N_15362);
and U15838 (N_15838,N_15548,N_15459);
nand U15839 (N_15839,N_15491,N_15364);
and U15840 (N_15840,N_15450,N_15447);
or U15841 (N_15841,N_15473,N_15558);
or U15842 (N_15842,N_15307,N_15367);
or U15843 (N_15843,N_15357,N_15523);
nor U15844 (N_15844,N_15465,N_15426);
and U15845 (N_15845,N_15551,N_15303);
nor U15846 (N_15846,N_15474,N_15435);
xnor U15847 (N_15847,N_15514,N_15449);
nand U15848 (N_15848,N_15500,N_15478);
or U15849 (N_15849,N_15381,N_15410);
xnor U15850 (N_15850,N_15549,N_15306);
and U15851 (N_15851,N_15458,N_15483);
nand U15852 (N_15852,N_15330,N_15407);
and U15853 (N_15853,N_15468,N_15308);
or U15854 (N_15854,N_15315,N_15472);
and U15855 (N_15855,N_15393,N_15423);
nor U15856 (N_15856,N_15478,N_15490);
and U15857 (N_15857,N_15587,N_15450);
nor U15858 (N_15858,N_15347,N_15512);
xor U15859 (N_15859,N_15356,N_15523);
xor U15860 (N_15860,N_15411,N_15429);
and U15861 (N_15861,N_15378,N_15430);
xnor U15862 (N_15862,N_15522,N_15447);
nor U15863 (N_15863,N_15340,N_15491);
nand U15864 (N_15864,N_15545,N_15552);
xnor U15865 (N_15865,N_15534,N_15493);
nor U15866 (N_15866,N_15356,N_15565);
nand U15867 (N_15867,N_15467,N_15380);
nand U15868 (N_15868,N_15532,N_15530);
or U15869 (N_15869,N_15387,N_15430);
and U15870 (N_15870,N_15576,N_15449);
nand U15871 (N_15871,N_15352,N_15594);
nor U15872 (N_15872,N_15381,N_15334);
nand U15873 (N_15873,N_15382,N_15313);
nand U15874 (N_15874,N_15361,N_15336);
or U15875 (N_15875,N_15403,N_15416);
nor U15876 (N_15876,N_15403,N_15335);
or U15877 (N_15877,N_15480,N_15522);
nor U15878 (N_15878,N_15365,N_15426);
or U15879 (N_15879,N_15569,N_15447);
or U15880 (N_15880,N_15540,N_15452);
nor U15881 (N_15881,N_15497,N_15356);
and U15882 (N_15882,N_15565,N_15579);
xnor U15883 (N_15883,N_15399,N_15377);
or U15884 (N_15884,N_15540,N_15460);
and U15885 (N_15885,N_15519,N_15433);
xnor U15886 (N_15886,N_15415,N_15502);
and U15887 (N_15887,N_15507,N_15462);
xnor U15888 (N_15888,N_15419,N_15397);
nor U15889 (N_15889,N_15489,N_15320);
and U15890 (N_15890,N_15525,N_15395);
and U15891 (N_15891,N_15401,N_15412);
or U15892 (N_15892,N_15310,N_15594);
and U15893 (N_15893,N_15311,N_15340);
and U15894 (N_15894,N_15426,N_15356);
and U15895 (N_15895,N_15491,N_15543);
nor U15896 (N_15896,N_15402,N_15463);
nor U15897 (N_15897,N_15533,N_15306);
and U15898 (N_15898,N_15559,N_15367);
and U15899 (N_15899,N_15417,N_15523);
or U15900 (N_15900,N_15714,N_15831);
nand U15901 (N_15901,N_15671,N_15746);
nor U15902 (N_15902,N_15867,N_15793);
or U15903 (N_15903,N_15672,N_15639);
and U15904 (N_15904,N_15777,N_15760);
and U15905 (N_15905,N_15873,N_15801);
and U15906 (N_15906,N_15790,N_15641);
xnor U15907 (N_15907,N_15841,N_15897);
xor U15908 (N_15908,N_15886,N_15706);
xnor U15909 (N_15909,N_15617,N_15614);
xnor U15910 (N_15910,N_15788,N_15845);
and U15911 (N_15911,N_15705,N_15797);
and U15912 (N_15912,N_15895,N_15724);
xor U15913 (N_15913,N_15715,N_15835);
or U15914 (N_15914,N_15851,N_15602);
and U15915 (N_15915,N_15838,N_15635);
xnor U15916 (N_15916,N_15823,N_15761);
and U15917 (N_15917,N_15758,N_15811);
xnor U15918 (N_15918,N_15814,N_15670);
and U15919 (N_15919,N_15855,N_15794);
xnor U15920 (N_15920,N_15654,N_15698);
nor U15921 (N_15921,N_15629,N_15604);
nand U15922 (N_15922,N_15800,N_15843);
nand U15923 (N_15923,N_15829,N_15711);
nor U15924 (N_15924,N_15680,N_15870);
nor U15925 (N_15925,N_15741,N_15721);
nand U15926 (N_15926,N_15806,N_15893);
xnor U15927 (N_15927,N_15807,N_15858);
xor U15928 (N_15928,N_15815,N_15633);
nand U15929 (N_15929,N_15780,N_15749);
nand U15930 (N_15930,N_15837,N_15691);
nand U15931 (N_15931,N_15832,N_15609);
and U15932 (N_15932,N_15630,N_15877);
or U15933 (N_15933,N_15891,N_15669);
and U15934 (N_15934,N_15628,N_15701);
nand U15935 (N_15935,N_15673,N_15659);
nor U15936 (N_15936,N_15764,N_15735);
and U15937 (N_15937,N_15812,N_15871);
and U15938 (N_15938,N_15846,N_15729);
or U15939 (N_15939,N_15637,N_15658);
or U15940 (N_15940,N_15616,N_15830);
xor U15941 (N_15941,N_15876,N_15679);
xnor U15942 (N_15942,N_15852,N_15736);
or U15943 (N_15943,N_15767,N_15779);
nor U15944 (N_15944,N_15881,N_15896);
nor U15945 (N_15945,N_15888,N_15803);
or U15946 (N_15946,N_15697,N_15748);
and U15947 (N_15947,N_15847,N_15799);
and U15948 (N_15948,N_15603,N_15791);
or U15949 (N_15949,N_15763,N_15821);
nand U15950 (N_15950,N_15663,N_15681);
nand U15951 (N_15951,N_15668,N_15605);
or U15952 (N_15952,N_15720,N_15700);
and U15953 (N_15953,N_15693,N_15827);
xor U15954 (N_15954,N_15685,N_15770);
xor U15955 (N_15955,N_15613,N_15836);
xnor U15956 (N_15956,N_15684,N_15733);
and U15957 (N_15957,N_15833,N_15622);
or U15958 (N_15958,N_15734,N_15861);
and U15959 (N_15959,N_15784,N_15822);
nand U15960 (N_15960,N_15849,N_15810);
nor U15961 (N_15961,N_15772,N_15677);
nand U15962 (N_15962,N_15620,N_15786);
xnor U15963 (N_15963,N_15712,N_15728);
nor U15964 (N_15964,N_15774,N_15854);
or U15965 (N_15965,N_15675,N_15664);
or U15966 (N_15966,N_15828,N_15879);
or U15967 (N_15967,N_15740,N_15783);
or U15968 (N_15968,N_15642,N_15752);
or U15969 (N_15969,N_15632,N_15765);
or U15970 (N_15970,N_15696,N_15730);
xnor U15971 (N_15971,N_15826,N_15690);
nand U15972 (N_15972,N_15844,N_15762);
and U15973 (N_15973,N_15703,N_15688);
nand U15974 (N_15974,N_15636,N_15878);
and U15975 (N_15975,N_15816,N_15716);
xor U15976 (N_15976,N_15731,N_15775);
nand U15977 (N_15977,N_15709,N_15742);
or U15978 (N_15978,N_15808,N_15725);
nand U15979 (N_15979,N_15645,N_15638);
or U15980 (N_15980,N_15789,N_15651);
nand U15981 (N_15981,N_15623,N_15695);
or U15982 (N_15982,N_15899,N_15866);
nand U15983 (N_15983,N_15708,N_15750);
nand U15984 (N_15984,N_15853,N_15759);
nor U15985 (N_15985,N_15880,N_15850);
or U15986 (N_15986,N_15771,N_15648);
and U15987 (N_15987,N_15805,N_15656);
xnor U15988 (N_15988,N_15834,N_15683);
xor U15989 (N_15989,N_15615,N_15666);
nand U15990 (N_15990,N_15678,N_15610);
nand U15991 (N_15991,N_15719,N_15792);
and U15992 (N_15992,N_15824,N_15694);
nand U15993 (N_15993,N_15860,N_15722);
nand U15994 (N_15994,N_15732,N_15754);
nand U15995 (N_15995,N_15600,N_15862);
and U15996 (N_15996,N_15612,N_15773);
or U15997 (N_15997,N_15813,N_15650);
nor U15998 (N_15998,N_15753,N_15796);
nor U15999 (N_15999,N_15809,N_15781);
and U16000 (N_16000,N_15624,N_15874);
and U16001 (N_16001,N_15665,N_15872);
xnor U16002 (N_16002,N_15757,N_15782);
and U16003 (N_16003,N_15739,N_15787);
nand U16004 (N_16004,N_15898,N_15857);
or U16005 (N_16005,N_15768,N_15713);
xor U16006 (N_16006,N_15621,N_15820);
nand U16007 (N_16007,N_15848,N_15737);
nor U16008 (N_16008,N_15798,N_15869);
nor U16009 (N_16009,N_15755,N_15640);
and U16010 (N_16010,N_15692,N_15661);
and U16011 (N_16011,N_15892,N_15751);
and U16012 (N_16012,N_15887,N_15894);
xor U16013 (N_16013,N_15611,N_15747);
xnor U16014 (N_16014,N_15804,N_15743);
nor U16015 (N_16015,N_15723,N_15889);
nand U16016 (N_16016,N_15634,N_15864);
nand U16017 (N_16017,N_15819,N_15676);
and U16018 (N_16018,N_15704,N_15646);
or U16019 (N_16019,N_15601,N_15618);
nor U16020 (N_16020,N_15863,N_15776);
and U16021 (N_16021,N_15756,N_15882);
xnor U16022 (N_16022,N_15607,N_15608);
nor U16023 (N_16023,N_15842,N_15689);
xor U16024 (N_16024,N_15840,N_15859);
nor U16025 (N_16025,N_15643,N_15884);
xor U16026 (N_16026,N_15883,N_15868);
or U16027 (N_16027,N_15660,N_15745);
xor U16028 (N_16028,N_15686,N_15710);
and U16029 (N_16029,N_15653,N_15631);
nor U16030 (N_16030,N_15795,N_15785);
xor U16031 (N_16031,N_15699,N_15652);
nor U16032 (N_16032,N_15839,N_15718);
and U16033 (N_16033,N_15606,N_15744);
or U16034 (N_16034,N_15687,N_15657);
and U16035 (N_16035,N_15619,N_15682);
nor U16036 (N_16036,N_15626,N_15856);
nand U16037 (N_16037,N_15865,N_15717);
nand U16038 (N_16038,N_15802,N_15885);
xnor U16039 (N_16039,N_15738,N_15778);
and U16040 (N_16040,N_15707,N_15649);
nand U16041 (N_16041,N_15625,N_15766);
and U16042 (N_16042,N_15655,N_15667);
xnor U16043 (N_16043,N_15818,N_15817);
or U16044 (N_16044,N_15644,N_15726);
nor U16045 (N_16045,N_15702,N_15674);
or U16046 (N_16046,N_15727,N_15769);
nand U16047 (N_16047,N_15627,N_15825);
or U16048 (N_16048,N_15890,N_15662);
or U16049 (N_16049,N_15647,N_15875);
or U16050 (N_16050,N_15693,N_15897);
nand U16051 (N_16051,N_15710,N_15607);
nand U16052 (N_16052,N_15737,N_15633);
nor U16053 (N_16053,N_15619,N_15758);
or U16054 (N_16054,N_15871,N_15834);
xnor U16055 (N_16055,N_15624,N_15620);
nand U16056 (N_16056,N_15858,N_15673);
nor U16057 (N_16057,N_15762,N_15770);
xor U16058 (N_16058,N_15813,N_15876);
or U16059 (N_16059,N_15676,N_15698);
nand U16060 (N_16060,N_15880,N_15832);
xnor U16061 (N_16061,N_15630,N_15770);
or U16062 (N_16062,N_15705,N_15696);
xor U16063 (N_16063,N_15848,N_15638);
nor U16064 (N_16064,N_15686,N_15765);
xor U16065 (N_16065,N_15624,N_15666);
and U16066 (N_16066,N_15771,N_15721);
xor U16067 (N_16067,N_15804,N_15746);
nand U16068 (N_16068,N_15649,N_15683);
nand U16069 (N_16069,N_15767,N_15692);
or U16070 (N_16070,N_15713,N_15896);
and U16071 (N_16071,N_15737,N_15877);
nand U16072 (N_16072,N_15733,N_15840);
or U16073 (N_16073,N_15682,N_15741);
and U16074 (N_16074,N_15887,N_15802);
xnor U16075 (N_16075,N_15691,N_15886);
and U16076 (N_16076,N_15781,N_15628);
xor U16077 (N_16077,N_15857,N_15708);
xnor U16078 (N_16078,N_15751,N_15805);
xnor U16079 (N_16079,N_15610,N_15688);
nand U16080 (N_16080,N_15717,N_15707);
and U16081 (N_16081,N_15829,N_15787);
xnor U16082 (N_16082,N_15681,N_15651);
nor U16083 (N_16083,N_15616,N_15864);
nor U16084 (N_16084,N_15748,N_15852);
xor U16085 (N_16085,N_15738,N_15803);
nand U16086 (N_16086,N_15690,N_15844);
nand U16087 (N_16087,N_15844,N_15659);
xnor U16088 (N_16088,N_15773,N_15737);
nand U16089 (N_16089,N_15748,N_15678);
and U16090 (N_16090,N_15752,N_15678);
nor U16091 (N_16091,N_15879,N_15679);
xor U16092 (N_16092,N_15675,N_15744);
and U16093 (N_16093,N_15676,N_15710);
nor U16094 (N_16094,N_15634,N_15631);
xor U16095 (N_16095,N_15640,N_15673);
and U16096 (N_16096,N_15633,N_15784);
or U16097 (N_16097,N_15872,N_15804);
or U16098 (N_16098,N_15880,N_15728);
nand U16099 (N_16099,N_15730,N_15660);
or U16100 (N_16100,N_15817,N_15873);
nand U16101 (N_16101,N_15776,N_15724);
xor U16102 (N_16102,N_15685,N_15710);
or U16103 (N_16103,N_15739,N_15775);
nand U16104 (N_16104,N_15618,N_15605);
xor U16105 (N_16105,N_15624,N_15767);
nor U16106 (N_16106,N_15635,N_15825);
xnor U16107 (N_16107,N_15794,N_15703);
and U16108 (N_16108,N_15891,N_15803);
or U16109 (N_16109,N_15641,N_15635);
xor U16110 (N_16110,N_15785,N_15606);
nor U16111 (N_16111,N_15792,N_15784);
nand U16112 (N_16112,N_15791,N_15737);
nand U16113 (N_16113,N_15802,N_15867);
xor U16114 (N_16114,N_15689,N_15851);
xnor U16115 (N_16115,N_15623,N_15762);
and U16116 (N_16116,N_15673,N_15619);
xor U16117 (N_16117,N_15837,N_15710);
nor U16118 (N_16118,N_15780,N_15793);
or U16119 (N_16119,N_15890,N_15786);
or U16120 (N_16120,N_15698,N_15786);
nand U16121 (N_16121,N_15707,N_15806);
xnor U16122 (N_16122,N_15824,N_15665);
and U16123 (N_16123,N_15793,N_15826);
or U16124 (N_16124,N_15669,N_15800);
xor U16125 (N_16125,N_15742,N_15692);
nand U16126 (N_16126,N_15875,N_15610);
xor U16127 (N_16127,N_15854,N_15787);
and U16128 (N_16128,N_15736,N_15744);
xnor U16129 (N_16129,N_15759,N_15672);
or U16130 (N_16130,N_15838,N_15639);
nor U16131 (N_16131,N_15756,N_15671);
nand U16132 (N_16132,N_15766,N_15795);
xor U16133 (N_16133,N_15789,N_15613);
or U16134 (N_16134,N_15628,N_15846);
xnor U16135 (N_16135,N_15629,N_15642);
and U16136 (N_16136,N_15762,N_15811);
nand U16137 (N_16137,N_15856,N_15777);
and U16138 (N_16138,N_15617,N_15804);
xnor U16139 (N_16139,N_15765,N_15806);
or U16140 (N_16140,N_15812,N_15771);
nor U16141 (N_16141,N_15725,N_15603);
and U16142 (N_16142,N_15613,N_15723);
nand U16143 (N_16143,N_15840,N_15804);
nor U16144 (N_16144,N_15717,N_15676);
nor U16145 (N_16145,N_15781,N_15785);
or U16146 (N_16146,N_15722,N_15727);
and U16147 (N_16147,N_15887,N_15610);
xnor U16148 (N_16148,N_15619,N_15739);
xnor U16149 (N_16149,N_15825,N_15762);
nor U16150 (N_16150,N_15796,N_15807);
nor U16151 (N_16151,N_15801,N_15695);
xnor U16152 (N_16152,N_15763,N_15812);
or U16153 (N_16153,N_15634,N_15622);
xor U16154 (N_16154,N_15677,N_15600);
nor U16155 (N_16155,N_15840,N_15686);
nor U16156 (N_16156,N_15701,N_15820);
nand U16157 (N_16157,N_15630,N_15647);
and U16158 (N_16158,N_15676,N_15650);
or U16159 (N_16159,N_15814,N_15610);
nor U16160 (N_16160,N_15671,N_15751);
nor U16161 (N_16161,N_15681,N_15886);
or U16162 (N_16162,N_15614,N_15625);
nand U16163 (N_16163,N_15897,N_15691);
nor U16164 (N_16164,N_15699,N_15761);
xnor U16165 (N_16165,N_15846,N_15860);
nand U16166 (N_16166,N_15643,N_15602);
and U16167 (N_16167,N_15786,N_15892);
and U16168 (N_16168,N_15693,N_15882);
nor U16169 (N_16169,N_15867,N_15758);
or U16170 (N_16170,N_15823,N_15774);
and U16171 (N_16171,N_15790,N_15733);
or U16172 (N_16172,N_15833,N_15788);
nor U16173 (N_16173,N_15627,N_15640);
nor U16174 (N_16174,N_15731,N_15740);
xor U16175 (N_16175,N_15610,N_15659);
and U16176 (N_16176,N_15683,N_15867);
xor U16177 (N_16177,N_15889,N_15665);
or U16178 (N_16178,N_15793,N_15766);
or U16179 (N_16179,N_15671,N_15742);
xnor U16180 (N_16180,N_15888,N_15841);
nand U16181 (N_16181,N_15836,N_15897);
nor U16182 (N_16182,N_15604,N_15616);
nand U16183 (N_16183,N_15642,N_15616);
nor U16184 (N_16184,N_15660,N_15651);
nand U16185 (N_16185,N_15615,N_15620);
and U16186 (N_16186,N_15639,N_15704);
xnor U16187 (N_16187,N_15696,N_15672);
xor U16188 (N_16188,N_15807,N_15827);
nor U16189 (N_16189,N_15714,N_15712);
nand U16190 (N_16190,N_15829,N_15660);
or U16191 (N_16191,N_15887,N_15826);
nor U16192 (N_16192,N_15797,N_15846);
xor U16193 (N_16193,N_15695,N_15813);
nor U16194 (N_16194,N_15791,N_15727);
nor U16195 (N_16195,N_15774,N_15760);
nand U16196 (N_16196,N_15729,N_15735);
nand U16197 (N_16197,N_15718,N_15649);
or U16198 (N_16198,N_15801,N_15898);
nor U16199 (N_16199,N_15723,N_15800);
xor U16200 (N_16200,N_15923,N_16130);
nor U16201 (N_16201,N_15944,N_15995);
and U16202 (N_16202,N_16195,N_16158);
xor U16203 (N_16203,N_15912,N_16100);
nor U16204 (N_16204,N_15918,N_16095);
nand U16205 (N_16205,N_16099,N_16044);
nand U16206 (N_16206,N_15903,N_15971);
nor U16207 (N_16207,N_16010,N_16058);
and U16208 (N_16208,N_16017,N_15951);
nor U16209 (N_16209,N_16114,N_15902);
and U16210 (N_16210,N_16021,N_16077);
and U16211 (N_16211,N_16034,N_16137);
and U16212 (N_16212,N_16084,N_16080);
nand U16213 (N_16213,N_16116,N_16008);
nor U16214 (N_16214,N_16161,N_16167);
xor U16215 (N_16215,N_16157,N_16170);
or U16216 (N_16216,N_15982,N_16165);
nand U16217 (N_16217,N_15927,N_16073);
and U16218 (N_16218,N_16122,N_15970);
xor U16219 (N_16219,N_16191,N_15996);
nor U16220 (N_16220,N_15973,N_16036);
or U16221 (N_16221,N_16139,N_16138);
nor U16222 (N_16222,N_16169,N_15922);
nor U16223 (N_16223,N_16088,N_16063);
xor U16224 (N_16224,N_16107,N_16082);
xor U16225 (N_16225,N_16031,N_15985);
xor U16226 (N_16226,N_16052,N_15939);
nand U16227 (N_16227,N_16192,N_15924);
and U16228 (N_16228,N_15954,N_15901);
nand U16229 (N_16229,N_15916,N_16019);
and U16230 (N_16230,N_16150,N_15919);
xnor U16231 (N_16231,N_16164,N_15943);
xnor U16232 (N_16232,N_16042,N_16096);
or U16233 (N_16233,N_16018,N_16033);
nand U16234 (N_16234,N_16127,N_16079);
xnor U16235 (N_16235,N_15921,N_15959);
nor U16236 (N_16236,N_16009,N_16133);
or U16237 (N_16237,N_15917,N_16120);
xor U16238 (N_16238,N_15932,N_16119);
xor U16239 (N_16239,N_15975,N_16196);
xnor U16240 (N_16240,N_16135,N_16003);
nand U16241 (N_16241,N_16145,N_15962);
xnor U16242 (N_16242,N_15910,N_16179);
xnor U16243 (N_16243,N_16012,N_15987);
or U16244 (N_16244,N_16043,N_16154);
or U16245 (N_16245,N_15976,N_16051);
xor U16246 (N_16246,N_15984,N_15994);
xnor U16247 (N_16247,N_16013,N_16155);
nor U16248 (N_16248,N_15960,N_15993);
and U16249 (N_16249,N_16027,N_15964);
or U16250 (N_16250,N_16014,N_16144);
nor U16251 (N_16251,N_16109,N_16177);
and U16252 (N_16252,N_16175,N_16186);
or U16253 (N_16253,N_16152,N_16029);
or U16254 (N_16254,N_16199,N_15940);
or U16255 (N_16255,N_16092,N_16136);
nor U16256 (N_16256,N_16190,N_15999);
xor U16257 (N_16257,N_16141,N_16129);
and U16258 (N_16258,N_16056,N_16184);
xnor U16259 (N_16259,N_16030,N_16185);
nand U16260 (N_16260,N_15988,N_16097);
nand U16261 (N_16261,N_15956,N_16053);
nor U16262 (N_16262,N_16041,N_16047);
nand U16263 (N_16263,N_15926,N_16070);
nor U16264 (N_16264,N_16168,N_16124);
nand U16265 (N_16265,N_16037,N_16083);
xnor U16266 (N_16266,N_16151,N_16061);
or U16267 (N_16267,N_16085,N_15908);
and U16268 (N_16268,N_16148,N_15950);
and U16269 (N_16269,N_16194,N_15935);
and U16270 (N_16270,N_15915,N_16032);
xor U16271 (N_16271,N_16011,N_16005);
nand U16272 (N_16272,N_15933,N_16121);
nand U16273 (N_16273,N_16147,N_16113);
or U16274 (N_16274,N_16086,N_16140);
nor U16275 (N_16275,N_15930,N_15969);
or U16276 (N_16276,N_16112,N_16125);
or U16277 (N_16277,N_16038,N_15997);
xnor U16278 (N_16278,N_16143,N_16183);
or U16279 (N_16279,N_15913,N_16171);
nand U16280 (N_16280,N_15909,N_16098);
nand U16281 (N_16281,N_16103,N_15946);
or U16282 (N_16282,N_16166,N_16162);
and U16283 (N_16283,N_15977,N_16015);
or U16284 (N_16284,N_16105,N_16134);
nor U16285 (N_16285,N_16068,N_16176);
nor U16286 (N_16286,N_15907,N_15952);
xor U16287 (N_16287,N_15953,N_16101);
nand U16288 (N_16288,N_16146,N_16123);
and U16289 (N_16289,N_16142,N_15928);
nor U16290 (N_16290,N_15947,N_16132);
or U16291 (N_16291,N_16126,N_15948);
and U16292 (N_16292,N_15938,N_15972);
nor U16293 (N_16293,N_16023,N_15961);
or U16294 (N_16294,N_16000,N_15941);
or U16295 (N_16295,N_16045,N_16057);
nand U16296 (N_16296,N_15931,N_15966);
or U16297 (N_16297,N_15942,N_16048);
nor U16298 (N_16298,N_16102,N_16002);
nand U16299 (N_16299,N_16060,N_16090);
and U16300 (N_16300,N_16024,N_16160);
nand U16301 (N_16301,N_16078,N_15968);
or U16302 (N_16302,N_16035,N_16159);
or U16303 (N_16303,N_15929,N_16091);
nor U16304 (N_16304,N_15989,N_16075);
and U16305 (N_16305,N_16128,N_16016);
and U16306 (N_16306,N_15983,N_16111);
nand U16307 (N_16307,N_16094,N_15958);
or U16308 (N_16308,N_16004,N_15900);
xor U16309 (N_16309,N_16153,N_16087);
nand U16310 (N_16310,N_16180,N_16055);
nor U16311 (N_16311,N_16059,N_15992);
or U16312 (N_16312,N_16039,N_16065);
or U16313 (N_16313,N_15914,N_15986);
or U16314 (N_16314,N_16028,N_15967);
xor U16315 (N_16315,N_16174,N_16001);
xnor U16316 (N_16316,N_16049,N_16007);
nand U16317 (N_16317,N_16093,N_16072);
or U16318 (N_16318,N_16081,N_16110);
xnor U16319 (N_16319,N_15998,N_15904);
or U16320 (N_16320,N_16178,N_15963);
nand U16321 (N_16321,N_15925,N_16067);
xnor U16322 (N_16322,N_16117,N_16163);
nor U16323 (N_16323,N_16198,N_15978);
nor U16324 (N_16324,N_16173,N_16187);
and U16325 (N_16325,N_16089,N_16046);
nor U16326 (N_16326,N_16156,N_15936);
and U16327 (N_16327,N_16074,N_16149);
nand U16328 (N_16328,N_16106,N_16115);
or U16329 (N_16329,N_16182,N_16069);
nand U16330 (N_16330,N_16104,N_16189);
or U16331 (N_16331,N_15979,N_16108);
nor U16332 (N_16332,N_16022,N_16131);
nor U16333 (N_16333,N_16006,N_15981);
xor U16334 (N_16334,N_16064,N_16062);
and U16335 (N_16335,N_16040,N_15957);
and U16336 (N_16336,N_15965,N_16076);
nand U16337 (N_16337,N_15906,N_15990);
nand U16338 (N_16338,N_15920,N_16197);
or U16339 (N_16339,N_15937,N_15949);
and U16340 (N_16340,N_15991,N_16188);
or U16341 (N_16341,N_16054,N_16025);
or U16342 (N_16342,N_16066,N_16181);
or U16343 (N_16343,N_15945,N_15974);
nand U16344 (N_16344,N_15955,N_15905);
nor U16345 (N_16345,N_16026,N_16172);
nand U16346 (N_16346,N_15911,N_15934);
or U16347 (N_16347,N_16118,N_16193);
and U16348 (N_16348,N_16020,N_16050);
nand U16349 (N_16349,N_16071,N_15980);
nor U16350 (N_16350,N_15982,N_16020);
and U16351 (N_16351,N_16171,N_15981);
and U16352 (N_16352,N_15964,N_16174);
or U16353 (N_16353,N_15998,N_16027);
nand U16354 (N_16354,N_16122,N_16019);
nand U16355 (N_16355,N_15994,N_16061);
xor U16356 (N_16356,N_16001,N_16158);
nand U16357 (N_16357,N_16164,N_16015);
nand U16358 (N_16358,N_16083,N_16068);
nor U16359 (N_16359,N_16070,N_15969);
nand U16360 (N_16360,N_16058,N_16085);
nor U16361 (N_16361,N_15919,N_16197);
xnor U16362 (N_16362,N_15998,N_16048);
nor U16363 (N_16363,N_16027,N_15996);
nor U16364 (N_16364,N_16163,N_16074);
nand U16365 (N_16365,N_15907,N_15973);
nor U16366 (N_16366,N_15966,N_16192);
nor U16367 (N_16367,N_16136,N_16036);
xor U16368 (N_16368,N_16061,N_16114);
xnor U16369 (N_16369,N_16018,N_16190);
nand U16370 (N_16370,N_16127,N_16055);
nand U16371 (N_16371,N_16170,N_16018);
xnor U16372 (N_16372,N_16011,N_16035);
xnor U16373 (N_16373,N_15950,N_15914);
xor U16374 (N_16374,N_15943,N_16194);
nand U16375 (N_16375,N_16010,N_15942);
nor U16376 (N_16376,N_16015,N_16030);
xor U16377 (N_16377,N_16050,N_16135);
nand U16378 (N_16378,N_16033,N_16025);
nor U16379 (N_16379,N_16043,N_16119);
and U16380 (N_16380,N_16095,N_16153);
or U16381 (N_16381,N_16012,N_16029);
nor U16382 (N_16382,N_16072,N_16145);
or U16383 (N_16383,N_16089,N_16018);
xor U16384 (N_16384,N_15943,N_16122);
or U16385 (N_16385,N_16050,N_16171);
and U16386 (N_16386,N_16081,N_16163);
and U16387 (N_16387,N_16027,N_15966);
nor U16388 (N_16388,N_15932,N_15933);
nand U16389 (N_16389,N_16014,N_16147);
nand U16390 (N_16390,N_16096,N_16073);
and U16391 (N_16391,N_16034,N_15989);
or U16392 (N_16392,N_15984,N_16054);
nand U16393 (N_16393,N_16188,N_16081);
or U16394 (N_16394,N_15939,N_16116);
nor U16395 (N_16395,N_15960,N_16010);
nand U16396 (N_16396,N_16104,N_16096);
and U16397 (N_16397,N_16184,N_16195);
or U16398 (N_16398,N_16140,N_16115);
nor U16399 (N_16399,N_16131,N_15961);
xnor U16400 (N_16400,N_16194,N_16061);
nor U16401 (N_16401,N_16185,N_16162);
xor U16402 (N_16402,N_16190,N_15980);
and U16403 (N_16403,N_15977,N_15972);
xor U16404 (N_16404,N_16134,N_16085);
nand U16405 (N_16405,N_15964,N_15953);
nor U16406 (N_16406,N_15992,N_15922);
nand U16407 (N_16407,N_16010,N_16057);
nor U16408 (N_16408,N_16134,N_16068);
and U16409 (N_16409,N_15927,N_16090);
xnor U16410 (N_16410,N_15985,N_16069);
nor U16411 (N_16411,N_15934,N_16111);
or U16412 (N_16412,N_16118,N_16141);
and U16413 (N_16413,N_16153,N_16180);
nand U16414 (N_16414,N_15901,N_16142);
nand U16415 (N_16415,N_16179,N_16105);
and U16416 (N_16416,N_16142,N_16116);
nand U16417 (N_16417,N_15978,N_16121);
and U16418 (N_16418,N_16178,N_16126);
or U16419 (N_16419,N_16100,N_15961);
xor U16420 (N_16420,N_15966,N_16038);
or U16421 (N_16421,N_15938,N_16005);
or U16422 (N_16422,N_16189,N_15959);
and U16423 (N_16423,N_15908,N_16198);
nor U16424 (N_16424,N_16130,N_16145);
nand U16425 (N_16425,N_15988,N_16099);
xor U16426 (N_16426,N_15929,N_15930);
nor U16427 (N_16427,N_16190,N_15938);
nand U16428 (N_16428,N_16010,N_16054);
nor U16429 (N_16429,N_16162,N_16157);
and U16430 (N_16430,N_16024,N_16094);
nor U16431 (N_16431,N_16150,N_15942);
and U16432 (N_16432,N_16095,N_15982);
xnor U16433 (N_16433,N_16106,N_16147);
nor U16434 (N_16434,N_15993,N_16062);
xnor U16435 (N_16435,N_15983,N_16174);
xor U16436 (N_16436,N_16005,N_16101);
or U16437 (N_16437,N_16102,N_16044);
xor U16438 (N_16438,N_15919,N_16104);
nand U16439 (N_16439,N_16163,N_16156);
and U16440 (N_16440,N_15954,N_16052);
nor U16441 (N_16441,N_16187,N_15952);
xor U16442 (N_16442,N_16160,N_15925);
and U16443 (N_16443,N_16073,N_16106);
and U16444 (N_16444,N_16087,N_16092);
nand U16445 (N_16445,N_16145,N_16112);
and U16446 (N_16446,N_15962,N_15972);
xnor U16447 (N_16447,N_15967,N_16026);
or U16448 (N_16448,N_15947,N_16185);
xnor U16449 (N_16449,N_16156,N_15906);
nand U16450 (N_16450,N_16185,N_15988);
or U16451 (N_16451,N_16151,N_16164);
and U16452 (N_16452,N_16097,N_16134);
and U16453 (N_16453,N_16145,N_16062);
xor U16454 (N_16454,N_16100,N_16114);
and U16455 (N_16455,N_16043,N_16175);
or U16456 (N_16456,N_16108,N_16128);
xnor U16457 (N_16457,N_16149,N_16104);
nor U16458 (N_16458,N_16197,N_15934);
nand U16459 (N_16459,N_16191,N_15914);
or U16460 (N_16460,N_15957,N_16070);
and U16461 (N_16461,N_16175,N_16161);
xor U16462 (N_16462,N_15984,N_15955);
nand U16463 (N_16463,N_16153,N_15995);
nor U16464 (N_16464,N_16037,N_16190);
and U16465 (N_16465,N_16111,N_15941);
xnor U16466 (N_16466,N_16054,N_16027);
or U16467 (N_16467,N_15985,N_16198);
and U16468 (N_16468,N_16028,N_15947);
nor U16469 (N_16469,N_15995,N_16048);
xor U16470 (N_16470,N_16061,N_15973);
xor U16471 (N_16471,N_16050,N_16048);
and U16472 (N_16472,N_16138,N_16110);
and U16473 (N_16473,N_16014,N_16043);
or U16474 (N_16474,N_16152,N_16192);
and U16475 (N_16475,N_16048,N_16022);
xnor U16476 (N_16476,N_16163,N_16183);
or U16477 (N_16477,N_16070,N_16199);
and U16478 (N_16478,N_16172,N_15914);
xor U16479 (N_16479,N_16072,N_16127);
xor U16480 (N_16480,N_16025,N_16022);
or U16481 (N_16481,N_16078,N_15908);
nand U16482 (N_16482,N_16079,N_15905);
and U16483 (N_16483,N_16152,N_16093);
nor U16484 (N_16484,N_16035,N_15972);
nor U16485 (N_16485,N_16006,N_16179);
xnor U16486 (N_16486,N_16085,N_16154);
and U16487 (N_16487,N_16043,N_15965);
xor U16488 (N_16488,N_16032,N_15903);
and U16489 (N_16489,N_16171,N_16001);
xnor U16490 (N_16490,N_16038,N_16152);
nor U16491 (N_16491,N_16191,N_16046);
or U16492 (N_16492,N_15962,N_16038);
and U16493 (N_16493,N_16055,N_16131);
nand U16494 (N_16494,N_15922,N_16183);
nor U16495 (N_16495,N_16158,N_15905);
nor U16496 (N_16496,N_15939,N_16115);
nand U16497 (N_16497,N_16119,N_16065);
and U16498 (N_16498,N_16059,N_16130);
nor U16499 (N_16499,N_16119,N_16134);
or U16500 (N_16500,N_16383,N_16251);
nor U16501 (N_16501,N_16283,N_16200);
xnor U16502 (N_16502,N_16417,N_16370);
nand U16503 (N_16503,N_16221,N_16236);
nand U16504 (N_16504,N_16422,N_16474);
and U16505 (N_16505,N_16354,N_16272);
xnor U16506 (N_16506,N_16223,N_16477);
nor U16507 (N_16507,N_16374,N_16202);
and U16508 (N_16508,N_16489,N_16387);
nor U16509 (N_16509,N_16267,N_16364);
nor U16510 (N_16510,N_16382,N_16280);
nor U16511 (N_16511,N_16259,N_16427);
nor U16512 (N_16512,N_16342,N_16429);
nor U16513 (N_16513,N_16344,N_16301);
xor U16514 (N_16514,N_16219,N_16490);
nand U16515 (N_16515,N_16320,N_16210);
and U16516 (N_16516,N_16303,N_16234);
and U16517 (N_16517,N_16231,N_16350);
nand U16518 (N_16518,N_16266,N_16414);
nor U16519 (N_16519,N_16304,N_16415);
or U16520 (N_16520,N_16478,N_16472);
nand U16521 (N_16521,N_16392,N_16444);
nand U16522 (N_16522,N_16361,N_16248);
xnor U16523 (N_16523,N_16449,N_16465);
xor U16524 (N_16524,N_16341,N_16306);
and U16525 (N_16525,N_16201,N_16212);
nand U16526 (N_16526,N_16277,N_16235);
xor U16527 (N_16527,N_16228,N_16243);
and U16528 (N_16528,N_16335,N_16327);
nand U16529 (N_16529,N_16332,N_16416);
nor U16530 (N_16530,N_16365,N_16456);
nand U16531 (N_16531,N_16268,N_16360);
or U16532 (N_16532,N_16488,N_16239);
or U16533 (N_16533,N_16476,N_16255);
xnor U16534 (N_16534,N_16211,N_16264);
xor U16535 (N_16535,N_16443,N_16278);
and U16536 (N_16536,N_16400,N_16351);
or U16537 (N_16537,N_16486,N_16302);
xnor U16538 (N_16538,N_16402,N_16294);
nor U16539 (N_16539,N_16419,N_16492);
and U16540 (N_16540,N_16324,N_16406);
nor U16541 (N_16541,N_16300,N_16205);
and U16542 (N_16542,N_16436,N_16377);
nand U16543 (N_16543,N_16273,N_16222);
or U16544 (N_16544,N_16495,N_16282);
xor U16545 (N_16545,N_16390,N_16346);
and U16546 (N_16546,N_16440,N_16404);
or U16547 (N_16547,N_16394,N_16225);
nand U16548 (N_16548,N_16467,N_16314);
nand U16549 (N_16549,N_16286,N_16224);
and U16550 (N_16550,N_16322,N_16499);
xnor U16551 (N_16551,N_16213,N_16330);
and U16552 (N_16552,N_16216,N_16423);
or U16553 (N_16553,N_16497,N_16431);
and U16554 (N_16554,N_16362,N_16437);
and U16555 (N_16555,N_16295,N_16418);
xnor U16556 (N_16556,N_16408,N_16289);
xnor U16557 (N_16557,N_16353,N_16333);
nor U16558 (N_16558,N_16454,N_16307);
or U16559 (N_16559,N_16349,N_16291);
nor U16560 (N_16560,N_16494,N_16411);
or U16561 (N_16561,N_16359,N_16217);
and U16562 (N_16562,N_16451,N_16410);
nor U16563 (N_16563,N_16479,N_16458);
nand U16564 (N_16564,N_16275,N_16297);
nand U16565 (N_16565,N_16457,N_16373);
and U16566 (N_16566,N_16347,N_16218);
and U16567 (N_16567,N_16355,N_16241);
and U16568 (N_16568,N_16203,N_16331);
or U16569 (N_16569,N_16305,N_16397);
nor U16570 (N_16570,N_16401,N_16396);
and U16571 (N_16571,N_16317,N_16460);
nand U16572 (N_16572,N_16384,N_16263);
xnor U16573 (N_16573,N_16484,N_16475);
or U16574 (N_16574,N_16238,N_16348);
nor U16575 (N_16575,N_16336,N_16244);
nor U16576 (N_16576,N_16481,N_16215);
nor U16577 (N_16577,N_16376,N_16292);
xnor U16578 (N_16578,N_16230,N_16247);
xnor U16579 (N_16579,N_16473,N_16375);
and U16580 (N_16580,N_16385,N_16206);
xnor U16581 (N_16581,N_16453,N_16338);
and U16582 (N_16582,N_16452,N_16455);
and U16583 (N_16583,N_16480,N_16381);
xor U16584 (N_16584,N_16288,N_16405);
xnor U16585 (N_16585,N_16391,N_16312);
and U16586 (N_16586,N_16464,N_16233);
or U16587 (N_16587,N_16246,N_16352);
and U16588 (N_16588,N_16372,N_16293);
and U16589 (N_16589,N_16462,N_16493);
nand U16590 (N_16590,N_16432,N_16363);
nand U16591 (N_16591,N_16298,N_16471);
nand U16592 (N_16592,N_16389,N_16334);
xor U16593 (N_16593,N_16463,N_16340);
xor U16594 (N_16594,N_16237,N_16380);
and U16595 (N_16595,N_16459,N_16445);
and U16596 (N_16596,N_16254,N_16367);
nor U16597 (N_16597,N_16369,N_16496);
nand U16598 (N_16598,N_16240,N_16220);
nor U16599 (N_16599,N_16366,N_16214);
xor U16600 (N_16600,N_16242,N_16262);
nand U16601 (N_16601,N_16326,N_16227);
and U16602 (N_16602,N_16448,N_16426);
or U16603 (N_16603,N_16466,N_16442);
nand U16604 (N_16604,N_16276,N_16207);
nor U16605 (N_16605,N_16325,N_16424);
or U16606 (N_16606,N_16296,N_16357);
xnor U16607 (N_16607,N_16321,N_16439);
xor U16608 (N_16608,N_16487,N_16409);
xor U16609 (N_16609,N_16270,N_16345);
xor U16610 (N_16610,N_16469,N_16485);
and U16611 (N_16611,N_16269,N_16433);
nand U16612 (N_16612,N_16287,N_16461);
nand U16613 (N_16613,N_16328,N_16318);
nor U16614 (N_16614,N_16249,N_16450);
xor U16615 (N_16615,N_16395,N_16308);
nand U16616 (N_16616,N_16204,N_16285);
or U16617 (N_16617,N_16398,N_16271);
nor U16618 (N_16618,N_16470,N_16393);
nor U16619 (N_16619,N_16343,N_16313);
xor U16620 (N_16620,N_16430,N_16319);
xnor U16621 (N_16621,N_16252,N_16209);
and U16622 (N_16622,N_16329,N_16309);
xnor U16623 (N_16623,N_16281,N_16229);
and U16624 (N_16624,N_16379,N_16434);
xor U16625 (N_16625,N_16378,N_16446);
nor U16626 (N_16626,N_16356,N_16428);
nor U16627 (N_16627,N_16388,N_16257);
nor U16628 (N_16628,N_16290,N_16368);
xor U16629 (N_16629,N_16258,N_16311);
xor U16630 (N_16630,N_16323,N_16425);
and U16631 (N_16631,N_16399,N_16253);
xor U16632 (N_16632,N_16284,N_16310);
and U16633 (N_16633,N_16265,N_16208);
nor U16634 (N_16634,N_16420,N_16412);
nor U16635 (N_16635,N_16299,N_16407);
nor U16636 (N_16636,N_16421,N_16250);
nand U16637 (N_16637,N_16358,N_16261);
xnor U16638 (N_16638,N_16245,N_16482);
and U16639 (N_16639,N_16483,N_16260);
xnor U16640 (N_16640,N_16274,N_16435);
xnor U16641 (N_16641,N_16279,N_16468);
nor U16642 (N_16642,N_16386,N_16256);
or U16643 (N_16643,N_16232,N_16315);
or U16644 (N_16644,N_16403,N_16438);
xor U16645 (N_16645,N_16339,N_16371);
or U16646 (N_16646,N_16491,N_16441);
xor U16647 (N_16647,N_16337,N_16498);
nor U16648 (N_16648,N_16447,N_16316);
nor U16649 (N_16649,N_16226,N_16413);
nor U16650 (N_16650,N_16362,N_16404);
nor U16651 (N_16651,N_16482,N_16219);
xnor U16652 (N_16652,N_16338,N_16279);
and U16653 (N_16653,N_16333,N_16464);
nand U16654 (N_16654,N_16410,N_16356);
xor U16655 (N_16655,N_16471,N_16433);
nand U16656 (N_16656,N_16366,N_16410);
nand U16657 (N_16657,N_16208,N_16409);
and U16658 (N_16658,N_16242,N_16218);
nor U16659 (N_16659,N_16369,N_16329);
nand U16660 (N_16660,N_16330,N_16313);
and U16661 (N_16661,N_16363,N_16382);
and U16662 (N_16662,N_16272,N_16361);
and U16663 (N_16663,N_16426,N_16374);
nand U16664 (N_16664,N_16207,N_16450);
or U16665 (N_16665,N_16445,N_16448);
and U16666 (N_16666,N_16267,N_16284);
xor U16667 (N_16667,N_16219,N_16363);
xor U16668 (N_16668,N_16494,N_16366);
nand U16669 (N_16669,N_16291,N_16216);
xnor U16670 (N_16670,N_16415,N_16456);
or U16671 (N_16671,N_16242,N_16477);
xnor U16672 (N_16672,N_16394,N_16370);
nand U16673 (N_16673,N_16245,N_16420);
or U16674 (N_16674,N_16323,N_16381);
nor U16675 (N_16675,N_16352,N_16476);
and U16676 (N_16676,N_16354,N_16393);
xnor U16677 (N_16677,N_16316,N_16439);
and U16678 (N_16678,N_16382,N_16481);
xnor U16679 (N_16679,N_16495,N_16489);
or U16680 (N_16680,N_16232,N_16422);
nor U16681 (N_16681,N_16338,N_16269);
nor U16682 (N_16682,N_16420,N_16342);
nor U16683 (N_16683,N_16499,N_16262);
nand U16684 (N_16684,N_16378,N_16457);
and U16685 (N_16685,N_16289,N_16399);
xnor U16686 (N_16686,N_16214,N_16277);
xor U16687 (N_16687,N_16412,N_16436);
or U16688 (N_16688,N_16478,N_16460);
xnor U16689 (N_16689,N_16272,N_16423);
or U16690 (N_16690,N_16230,N_16276);
xor U16691 (N_16691,N_16220,N_16295);
nor U16692 (N_16692,N_16336,N_16243);
and U16693 (N_16693,N_16224,N_16321);
or U16694 (N_16694,N_16320,N_16361);
nand U16695 (N_16695,N_16286,N_16237);
or U16696 (N_16696,N_16254,N_16286);
or U16697 (N_16697,N_16436,N_16271);
or U16698 (N_16698,N_16340,N_16333);
nor U16699 (N_16699,N_16461,N_16294);
and U16700 (N_16700,N_16477,N_16469);
or U16701 (N_16701,N_16287,N_16204);
and U16702 (N_16702,N_16220,N_16419);
nor U16703 (N_16703,N_16430,N_16318);
or U16704 (N_16704,N_16382,N_16294);
nand U16705 (N_16705,N_16300,N_16302);
xor U16706 (N_16706,N_16235,N_16256);
or U16707 (N_16707,N_16380,N_16460);
or U16708 (N_16708,N_16418,N_16225);
or U16709 (N_16709,N_16456,N_16313);
and U16710 (N_16710,N_16273,N_16373);
nor U16711 (N_16711,N_16392,N_16499);
or U16712 (N_16712,N_16308,N_16489);
xnor U16713 (N_16713,N_16291,N_16223);
and U16714 (N_16714,N_16387,N_16375);
or U16715 (N_16715,N_16251,N_16359);
xor U16716 (N_16716,N_16230,N_16304);
xor U16717 (N_16717,N_16309,N_16245);
nor U16718 (N_16718,N_16261,N_16399);
or U16719 (N_16719,N_16285,N_16261);
xnor U16720 (N_16720,N_16405,N_16237);
nand U16721 (N_16721,N_16312,N_16456);
and U16722 (N_16722,N_16389,N_16456);
and U16723 (N_16723,N_16276,N_16376);
nor U16724 (N_16724,N_16287,N_16479);
nor U16725 (N_16725,N_16243,N_16366);
nor U16726 (N_16726,N_16333,N_16359);
or U16727 (N_16727,N_16417,N_16273);
nor U16728 (N_16728,N_16242,N_16430);
and U16729 (N_16729,N_16225,N_16337);
or U16730 (N_16730,N_16348,N_16364);
and U16731 (N_16731,N_16216,N_16270);
or U16732 (N_16732,N_16238,N_16438);
and U16733 (N_16733,N_16305,N_16395);
nand U16734 (N_16734,N_16470,N_16385);
xnor U16735 (N_16735,N_16392,N_16334);
nand U16736 (N_16736,N_16484,N_16450);
and U16737 (N_16737,N_16471,N_16241);
or U16738 (N_16738,N_16265,N_16446);
nand U16739 (N_16739,N_16330,N_16363);
or U16740 (N_16740,N_16416,N_16329);
and U16741 (N_16741,N_16419,N_16493);
nor U16742 (N_16742,N_16360,N_16453);
and U16743 (N_16743,N_16299,N_16450);
nand U16744 (N_16744,N_16458,N_16330);
nor U16745 (N_16745,N_16453,N_16282);
or U16746 (N_16746,N_16427,N_16207);
xnor U16747 (N_16747,N_16336,N_16317);
xnor U16748 (N_16748,N_16439,N_16270);
nand U16749 (N_16749,N_16338,N_16200);
xnor U16750 (N_16750,N_16472,N_16492);
nor U16751 (N_16751,N_16495,N_16260);
xor U16752 (N_16752,N_16308,N_16408);
nor U16753 (N_16753,N_16364,N_16269);
or U16754 (N_16754,N_16282,N_16206);
nor U16755 (N_16755,N_16348,N_16404);
nand U16756 (N_16756,N_16487,N_16415);
nand U16757 (N_16757,N_16329,N_16235);
or U16758 (N_16758,N_16321,N_16370);
and U16759 (N_16759,N_16481,N_16433);
nor U16760 (N_16760,N_16491,N_16361);
nand U16761 (N_16761,N_16292,N_16341);
and U16762 (N_16762,N_16271,N_16372);
and U16763 (N_16763,N_16450,N_16419);
nand U16764 (N_16764,N_16331,N_16368);
or U16765 (N_16765,N_16293,N_16329);
and U16766 (N_16766,N_16456,N_16261);
nor U16767 (N_16767,N_16385,N_16201);
and U16768 (N_16768,N_16410,N_16316);
nor U16769 (N_16769,N_16240,N_16270);
nor U16770 (N_16770,N_16292,N_16470);
nand U16771 (N_16771,N_16318,N_16206);
and U16772 (N_16772,N_16300,N_16266);
nand U16773 (N_16773,N_16404,N_16430);
xnor U16774 (N_16774,N_16268,N_16263);
nand U16775 (N_16775,N_16379,N_16219);
and U16776 (N_16776,N_16312,N_16477);
nor U16777 (N_16777,N_16416,N_16290);
xor U16778 (N_16778,N_16273,N_16227);
and U16779 (N_16779,N_16254,N_16375);
xnor U16780 (N_16780,N_16337,N_16445);
or U16781 (N_16781,N_16469,N_16364);
nor U16782 (N_16782,N_16483,N_16208);
xor U16783 (N_16783,N_16405,N_16481);
nand U16784 (N_16784,N_16290,N_16264);
or U16785 (N_16785,N_16257,N_16326);
or U16786 (N_16786,N_16313,N_16364);
nor U16787 (N_16787,N_16484,N_16406);
or U16788 (N_16788,N_16416,N_16486);
nor U16789 (N_16789,N_16315,N_16299);
and U16790 (N_16790,N_16331,N_16403);
xor U16791 (N_16791,N_16307,N_16391);
and U16792 (N_16792,N_16236,N_16345);
xor U16793 (N_16793,N_16498,N_16358);
nand U16794 (N_16794,N_16277,N_16484);
and U16795 (N_16795,N_16298,N_16445);
and U16796 (N_16796,N_16400,N_16349);
or U16797 (N_16797,N_16311,N_16251);
xor U16798 (N_16798,N_16267,N_16328);
xor U16799 (N_16799,N_16484,N_16457);
xnor U16800 (N_16800,N_16548,N_16622);
and U16801 (N_16801,N_16647,N_16641);
or U16802 (N_16802,N_16660,N_16670);
xor U16803 (N_16803,N_16781,N_16631);
nand U16804 (N_16804,N_16630,N_16603);
nor U16805 (N_16805,N_16634,N_16519);
nand U16806 (N_16806,N_16503,N_16510);
or U16807 (N_16807,N_16564,N_16539);
xnor U16808 (N_16808,N_16667,N_16763);
and U16809 (N_16809,N_16502,N_16579);
or U16810 (N_16810,N_16595,N_16535);
xor U16811 (N_16811,N_16512,N_16669);
nand U16812 (N_16812,N_16786,N_16668);
nand U16813 (N_16813,N_16727,N_16561);
nor U16814 (N_16814,N_16626,N_16590);
or U16815 (N_16815,N_16697,N_16618);
and U16816 (N_16816,N_16505,N_16770);
nand U16817 (N_16817,N_16704,N_16735);
and U16818 (N_16818,N_16774,N_16683);
or U16819 (N_16819,N_16756,N_16625);
xnor U16820 (N_16820,N_16555,N_16705);
or U16821 (N_16821,N_16734,N_16644);
nor U16822 (N_16822,N_16788,N_16674);
nor U16823 (N_16823,N_16723,N_16717);
nor U16824 (N_16824,N_16587,N_16521);
nor U16825 (N_16825,N_16524,N_16602);
nand U16826 (N_16826,N_16643,N_16558);
nand U16827 (N_16827,N_16580,N_16741);
or U16828 (N_16828,N_16703,N_16550);
nand U16829 (N_16829,N_16720,N_16699);
nand U16830 (N_16830,N_16517,N_16591);
nand U16831 (N_16831,N_16744,N_16769);
nor U16832 (N_16832,N_16573,N_16716);
nand U16833 (N_16833,N_16585,N_16650);
nand U16834 (N_16834,N_16693,N_16515);
or U16835 (N_16835,N_16766,N_16633);
nor U16836 (N_16836,N_16533,N_16662);
nand U16837 (N_16837,N_16568,N_16549);
nand U16838 (N_16838,N_16627,N_16765);
or U16839 (N_16839,N_16612,N_16557);
xor U16840 (N_16840,N_16746,N_16728);
or U16841 (N_16841,N_16513,N_16552);
and U16842 (N_16842,N_16624,N_16500);
or U16843 (N_16843,N_16575,N_16787);
nand U16844 (N_16844,N_16676,N_16509);
nor U16845 (N_16845,N_16702,N_16684);
or U16846 (N_16846,N_16791,N_16785);
xor U16847 (N_16847,N_16732,N_16594);
xor U16848 (N_16848,N_16598,N_16520);
nand U16849 (N_16849,N_16758,N_16721);
xor U16850 (N_16850,N_16745,N_16589);
and U16851 (N_16851,N_16711,N_16501);
nand U16852 (N_16852,N_16678,N_16530);
or U16853 (N_16853,N_16572,N_16783);
and U16854 (N_16854,N_16547,N_16688);
and U16855 (N_16855,N_16712,N_16692);
and U16856 (N_16856,N_16563,N_16709);
nor U16857 (N_16857,N_16581,N_16751);
or U16858 (N_16858,N_16556,N_16784);
xnor U16859 (N_16859,N_16689,N_16682);
xor U16860 (N_16860,N_16742,N_16796);
xnor U16861 (N_16861,N_16691,N_16588);
or U16862 (N_16862,N_16687,N_16708);
nand U16863 (N_16863,N_16738,N_16753);
xor U16864 (N_16864,N_16652,N_16780);
nor U16865 (N_16865,N_16752,N_16772);
nor U16866 (N_16866,N_16729,N_16565);
xor U16867 (N_16867,N_16764,N_16518);
nor U16868 (N_16868,N_16777,N_16790);
or U16869 (N_16869,N_16761,N_16794);
and U16870 (N_16870,N_16760,N_16642);
or U16871 (N_16871,N_16648,N_16645);
nor U16872 (N_16872,N_16577,N_16560);
nor U16873 (N_16873,N_16640,N_16593);
nand U16874 (N_16874,N_16508,N_16722);
xor U16875 (N_16875,N_16606,N_16661);
and U16876 (N_16876,N_16628,N_16554);
xnor U16877 (N_16877,N_16506,N_16797);
nand U16878 (N_16878,N_16750,N_16511);
nand U16879 (N_16879,N_16617,N_16657);
nand U16880 (N_16880,N_16775,N_16616);
nor U16881 (N_16881,N_16599,N_16671);
and U16882 (N_16882,N_16672,N_16675);
xnor U16883 (N_16883,N_16686,N_16632);
nand U16884 (N_16884,N_16586,N_16619);
nand U16885 (N_16885,N_16799,N_16559);
or U16886 (N_16886,N_16733,N_16719);
nand U16887 (N_16887,N_16639,N_16659);
xor U16888 (N_16888,N_16714,N_16706);
xor U16889 (N_16889,N_16516,N_16528);
xnor U16890 (N_16890,N_16677,N_16656);
and U16891 (N_16891,N_16615,N_16649);
nand U16892 (N_16892,N_16701,N_16740);
xor U16893 (N_16893,N_16507,N_16608);
nand U16894 (N_16894,N_16743,N_16798);
and U16895 (N_16895,N_16578,N_16654);
xor U16896 (N_16896,N_16685,N_16597);
xor U16897 (N_16897,N_16663,N_16567);
nor U16898 (N_16898,N_16646,N_16596);
and U16899 (N_16899,N_16638,N_16601);
or U16900 (N_16900,N_16525,N_16782);
nand U16901 (N_16901,N_16605,N_16522);
nor U16902 (N_16902,N_16610,N_16757);
xor U16903 (N_16903,N_16540,N_16607);
and U16904 (N_16904,N_16523,N_16747);
or U16905 (N_16905,N_16600,N_16504);
or U16906 (N_16906,N_16623,N_16541);
nor U16907 (N_16907,N_16749,N_16582);
and U16908 (N_16908,N_16576,N_16710);
xor U16909 (N_16909,N_16695,N_16566);
or U16910 (N_16910,N_16621,N_16551);
or U16911 (N_16911,N_16653,N_16694);
or U16912 (N_16912,N_16537,N_16536);
and U16913 (N_16913,N_16793,N_16574);
xor U16914 (N_16914,N_16544,N_16731);
nand U16915 (N_16915,N_16529,N_16754);
xor U16916 (N_16916,N_16637,N_16609);
nor U16917 (N_16917,N_16666,N_16680);
xor U16918 (N_16918,N_16771,N_16707);
nor U16919 (N_16919,N_16718,N_16534);
nand U16920 (N_16920,N_16759,N_16789);
or U16921 (N_16921,N_16543,N_16737);
xnor U16922 (N_16922,N_16553,N_16584);
or U16923 (N_16923,N_16532,N_16636);
and U16924 (N_16924,N_16773,N_16514);
xnor U16925 (N_16925,N_16604,N_16542);
nor U16926 (N_16926,N_16762,N_16778);
or U16927 (N_16927,N_16776,N_16739);
and U16928 (N_16928,N_16715,N_16779);
or U16929 (N_16929,N_16526,N_16571);
or U16930 (N_16930,N_16768,N_16613);
and U16931 (N_16931,N_16665,N_16726);
and U16932 (N_16932,N_16629,N_16673);
or U16933 (N_16933,N_16725,N_16748);
and U16934 (N_16934,N_16736,N_16583);
nand U16935 (N_16935,N_16679,N_16713);
and U16936 (N_16936,N_16545,N_16527);
or U16937 (N_16937,N_16655,N_16651);
xnor U16938 (N_16938,N_16611,N_16658);
or U16939 (N_16939,N_16755,N_16614);
nand U16940 (N_16940,N_16698,N_16620);
nand U16941 (N_16941,N_16538,N_16635);
and U16942 (N_16942,N_16696,N_16569);
nand U16943 (N_16943,N_16681,N_16795);
xor U16944 (N_16944,N_16690,N_16570);
or U16945 (N_16945,N_16664,N_16531);
nor U16946 (N_16946,N_16792,N_16730);
and U16947 (N_16947,N_16592,N_16562);
nor U16948 (N_16948,N_16724,N_16700);
or U16949 (N_16949,N_16767,N_16546);
xnor U16950 (N_16950,N_16752,N_16737);
nand U16951 (N_16951,N_16737,N_16666);
nand U16952 (N_16952,N_16718,N_16708);
nand U16953 (N_16953,N_16660,N_16549);
nor U16954 (N_16954,N_16639,N_16584);
nand U16955 (N_16955,N_16794,N_16518);
and U16956 (N_16956,N_16644,N_16695);
or U16957 (N_16957,N_16668,N_16572);
nand U16958 (N_16958,N_16545,N_16703);
xor U16959 (N_16959,N_16715,N_16602);
nor U16960 (N_16960,N_16564,N_16752);
xor U16961 (N_16961,N_16581,N_16580);
or U16962 (N_16962,N_16797,N_16551);
and U16963 (N_16963,N_16604,N_16543);
xnor U16964 (N_16964,N_16620,N_16539);
nor U16965 (N_16965,N_16667,N_16504);
xnor U16966 (N_16966,N_16720,N_16676);
nand U16967 (N_16967,N_16643,N_16517);
xnor U16968 (N_16968,N_16783,N_16562);
xor U16969 (N_16969,N_16657,N_16622);
or U16970 (N_16970,N_16547,N_16797);
or U16971 (N_16971,N_16677,N_16662);
and U16972 (N_16972,N_16553,N_16564);
and U16973 (N_16973,N_16780,N_16770);
xnor U16974 (N_16974,N_16637,N_16770);
and U16975 (N_16975,N_16643,N_16689);
or U16976 (N_16976,N_16717,N_16728);
nor U16977 (N_16977,N_16733,N_16789);
or U16978 (N_16978,N_16558,N_16759);
nand U16979 (N_16979,N_16566,N_16569);
nor U16980 (N_16980,N_16796,N_16726);
nor U16981 (N_16981,N_16624,N_16777);
and U16982 (N_16982,N_16681,N_16533);
xnor U16983 (N_16983,N_16577,N_16633);
nand U16984 (N_16984,N_16799,N_16664);
nor U16985 (N_16985,N_16708,N_16503);
xor U16986 (N_16986,N_16709,N_16692);
or U16987 (N_16987,N_16607,N_16600);
and U16988 (N_16988,N_16529,N_16602);
nor U16989 (N_16989,N_16626,N_16665);
xor U16990 (N_16990,N_16749,N_16612);
nor U16991 (N_16991,N_16734,N_16588);
nand U16992 (N_16992,N_16625,N_16723);
nor U16993 (N_16993,N_16689,N_16757);
nor U16994 (N_16994,N_16661,N_16543);
nor U16995 (N_16995,N_16787,N_16662);
or U16996 (N_16996,N_16506,N_16737);
xnor U16997 (N_16997,N_16753,N_16682);
nand U16998 (N_16998,N_16682,N_16561);
xnor U16999 (N_16999,N_16739,N_16794);
and U17000 (N_17000,N_16662,N_16768);
nor U17001 (N_17001,N_16588,N_16650);
or U17002 (N_17002,N_16660,N_16770);
nor U17003 (N_17003,N_16641,N_16519);
nor U17004 (N_17004,N_16762,N_16637);
xnor U17005 (N_17005,N_16777,N_16567);
xnor U17006 (N_17006,N_16782,N_16510);
nand U17007 (N_17007,N_16555,N_16579);
nand U17008 (N_17008,N_16613,N_16690);
or U17009 (N_17009,N_16520,N_16737);
nor U17010 (N_17010,N_16518,N_16684);
or U17011 (N_17011,N_16728,N_16500);
or U17012 (N_17012,N_16581,N_16539);
xor U17013 (N_17013,N_16796,N_16762);
nor U17014 (N_17014,N_16702,N_16701);
nand U17015 (N_17015,N_16749,N_16679);
xor U17016 (N_17016,N_16544,N_16539);
nand U17017 (N_17017,N_16798,N_16562);
or U17018 (N_17018,N_16759,N_16682);
nor U17019 (N_17019,N_16698,N_16546);
and U17020 (N_17020,N_16564,N_16547);
nor U17021 (N_17021,N_16795,N_16759);
and U17022 (N_17022,N_16664,N_16503);
xnor U17023 (N_17023,N_16772,N_16606);
nand U17024 (N_17024,N_16722,N_16783);
and U17025 (N_17025,N_16573,N_16734);
xor U17026 (N_17026,N_16772,N_16513);
and U17027 (N_17027,N_16693,N_16637);
nor U17028 (N_17028,N_16634,N_16550);
nand U17029 (N_17029,N_16775,N_16707);
xnor U17030 (N_17030,N_16565,N_16648);
nand U17031 (N_17031,N_16542,N_16619);
xnor U17032 (N_17032,N_16522,N_16534);
xnor U17033 (N_17033,N_16501,N_16523);
and U17034 (N_17034,N_16798,N_16555);
or U17035 (N_17035,N_16663,N_16699);
and U17036 (N_17036,N_16508,N_16561);
or U17037 (N_17037,N_16531,N_16563);
nor U17038 (N_17038,N_16736,N_16625);
and U17039 (N_17039,N_16555,N_16564);
xor U17040 (N_17040,N_16664,N_16759);
nor U17041 (N_17041,N_16607,N_16764);
nand U17042 (N_17042,N_16574,N_16797);
and U17043 (N_17043,N_16550,N_16704);
nand U17044 (N_17044,N_16628,N_16540);
xnor U17045 (N_17045,N_16748,N_16720);
or U17046 (N_17046,N_16724,N_16707);
or U17047 (N_17047,N_16791,N_16746);
nand U17048 (N_17048,N_16706,N_16713);
xor U17049 (N_17049,N_16714,N_16694);
xnor U17050 (N_17050,N_16724,N_16543);
nand U17051 (N_17051,N_16676,N_16675);
or U17052 (N_17052,N_16721,N_16794);
or U17053 (N_17053,N_16773,N_16709);
and U17054 (N_17054,N_16575,N_16737);
nor U17055 (N_17055,N_16648,N_16524);
nand U17056 (N_17056,N_16580,N_16592);
or U17057 (N_17057,N_16595,N_16747);
nand U17058 (N_17058,N_16776,N_16549);
or U17059 (N_17059,N_16785,N_16704);
or U17060 (N_17060,N_16713,N_16715);
and U17061 (N_17061,N_16638,N_16526);
nand U17062 (N_17062,N_16651,N_16795);
nand U17063 (N_17063,N_16721,N_16646);
or U17064 (N_17064,N_16554,N_16635);
and U17065 (N_17065,N_16764,N_16656);
and U17066 (N_17066,N_16793,N_16581);
nor U17067 (N_17067,N_16559,N_16690);
xnor U17068 (N_17068,N_16529,N_16715);
nand U17069 (N_17069,N_16753,N_16691);
nand U17070 (N_17070,N_16735,N_16796);
xnor U17071 (N_17071,N_16628,N_16702);
nand U17072 (N_17072,N_16603,N_16674);
nor U17073 (N_17073,N_16542,N_16556);
and U17074 (N_17074,N_16761,N_16618);
or U17075 (N_17075,N_16560,N_16722);
and U17076 (N_17076,N_16542,N_16514);
nand U17077 (N_17077,N_16611,N_16693);
nand U17078 (N_17078,N_16787,N_16643);
or U17079 (N_17079,N_16545,N_16764);
nor U17080 (N_17080,N_16587,N_16511);
nand U17081 (N_17081,N_16586,N_16653);
nor U17082 (N_17082,N_16762,N_16634);
xnor U17083 (N_17083,N_16625,N_16630);
xor U17084 (N_17084,N_16694,N_16785);
xnor U17085 (N_17085,N_16571,N_16713);
and U17086 (N_17086,N_16536,N_16725);
nand U17087 (N_17087,N_16541,N_16770);
and U17088 (N_17088,N_16685,N_16674);
or U17089 (N_17089,N_16772,N_16567);
nor U17090 (N_17090,N_16759,N_16564);
and U17091 (N_17091,N_16527,N_16730);
nand U17092 (N_17092,N_16745,N_16664);
and U17093 (N_17093,N_16785,N_16729);
nor U17094 (N_17094,N_16729,N_16745);
xor U17095 (N_17095,N_16590,N_16549);
or U17096 (N_17096,N_16664,N_16601);
and U17097 (N_17097,N_16651,N_16797);
nor U17098 (N_17098,N_16623,N_16659);
xnor U17099 (N_17099,N_16547,N_16672);
xor U17100 (N_17100,N_16929,N_16916);
nor U17101 (N_17101,N_16823,N_16953);
or U17102 (N_17102,N_17070,N_16944);
or U17103 (N_17103,N_16937,N_16907);
and U17104 (N_17104,N_17065,N_16868);
nand U17105 (N_17105,N_16933,N_17080);
or U17106 (N_17106,N_16906,N_16915);
nand U17107 (N_17107,N_16967,N_16959);
nor U17108 (N_17108,N_17063,N_16973);
nor U17109 (N_17109,N_16840,N_16845);
nand U17110 (N_17110,N_17040,N_17067);
and U17111 (N_17111,N_16971,N_16816);
and U17112 (N_17112,N_16930,N_17034);
nand U17113 (N_17113,N_16895,N_16851);
xnor U17114 (N_17114,N_17026,N_16897);
nor U17115 (N_17115,N_16888,N_16969);
and U17116 (N_17116,N_17058,N_17086);
and U17117 (N_17117,N_16963,N_16908);
nor U17118 (N_17118,N_17093,N_17015);
or U17119 (N_17119,N_16941,N_16873);
nor U17120 (N_17120,N_17077,N_17002);
and U17121 (N_17121,N_17068,N_16945);
xor U17122 (N_17122,N_17021,N_17051);
nor U17123 (N_17123,N_16936,N_16875);
or U17124 (N_17124,N_17087,N_16882);
nor U17125 (N_17125,N_16821,N_17017);
and U17126 (N_17126,N_16866,N_16859);
nand U17127 (N_17127,N_16842,N_16827);
and U17128 (N_17128,N_16808,N_16849);
nor U17129 (N_17129,N_16834,N_17011);
nand U17130 (N_17130,N_16939,N_17033);
nand U17131 (N_17131,N_16976,N_16863);
or U17132 (N_17132,N_16870,N_16826);
nor U17133 (N_17133,N_16817,N_16932);
xnor U17134 (N_17134,N_17006,N_16996);
or U17135 (N_17135,N_17031,N_16865);
or U17136 (N_17136,N_16979,N_16946);
or U17137 (N_17137,N_16975,N_17007);
nand U17138 (N_17138,N_16954,N_16843);
nor U17139 (N_17139,N_17055,N_16950);
nand U17140 (N_17140,N_16813,N_16890);
nor U17141 (N_17141,N_16854,N_17013);
or U17142 (N_17142,N_16923,N_16948);
nand U17143 (N_17143,N_16958,N_16919);
and U17144 (N_17144,N_16861,N_17035);
and U17145 (N_17145,N_16892,N_17062);
nor U17146 (N_17146,N_16925,N_16984);
xnor U17147 (N_17147,N_16893,N_17053);
or U17148 (N_17148,N_16912,N_16980);
xor U17149 (N_17149,N_17092,N_16855);
nand U17150 (N_17150,N_16911,N_16998);
and U17151 (N_17151,N_16942,N_16844);
nor U17152 (N_17152,N_17066,N_17010);
xor U17153 (N_17153,N_17064,N_16830);
and U17154 (N_17154,N_16981,N_16904);
nand U17155 (N_17155,N_17044,N_16928);
xor U17156 (N_17156,N_17001,N_17003);
xnor U17157 (N_17157,N_16957,N_17050);
and U17158 (N_17158,N_16978,N_17041);
nand U17159 (N_17159,N_16860,N_16920);
or U17160 (N_17160,N_16815,N_16898);
and U17161 (N_17161,N_16804,N_16803);
or U17162 (N_17162,N_17060,N_17098);
nor U17163 (N_17163,N_16924,N_16814);
or U17164 (N_17164,N_17019,N_16972);
nand U17165 (N_17165,N_16955,N_16931);
nand U17166 (N_17166,N_16820,N_16995);
xnor U17167 (N_17167,N_16993,N_17042);
or U17168 (N_17168,N_16988,N_16856);
or U17169 (N_17169,N_16974,N_16951);
xnor U17170 (N_17170,N_16881,N_16837);
and U17171 (N_17171,N_16864,N_17032);
nor U17172 (N_17172,N_16968,N_16848);
nand U17173 (N_17173,N_16934,N_16901);
and U17174 (N_17174,N_16990,N_17012);
and U17175 (N_17175,N_16889,N_16852);
nor U17176 (N_17176,N_16987,N_16879);
or U17177 (N_17177,N_17048,N_16811);
and U17178 (N_17178,N_16836,N_16961);
xnor U17179 (N_17179,N_17029,N_16994);
nand U17180 (N_17180,N_16805,N_17038);
nor U17181 (N_17181,N_16902,N_16956);
xnor U17182 (N_17182,N_16986,N_16943);
or U17183 (N_17183,N_17085,N_17099);
and U17184 (N_17184,N_16867,N_17084);
or U17185 (N_17185,N_16896,N_16921);
or U17186 (N_17186,N_16846,N_17024);
or U17187 (N_17187,N_17046,N_17005);
or U17188 (N_17188,N_16997,N_16831);
xnor U17189 (N_17189,N_16985,N_16964);
and U17190 (N_17190,N_16802,N_16887);
nand U17191 (N_17191,N_16914,N_16886);
xor U17192 (N_17192,N_17081,N_16913);
and U17193 (N_17193,N_17061,N_17047);
nor U17194 (N_17194,N_16917,N_17057);
nor U17195 (N_17195,N_16960,N_17014);
xor U17196 (N_17196,N_16853,N_16922);
and U17197 (N_17197,N_16819,N_16927);
xnor U17198 (N_17198,N_17089,N_17071);
and U17199 (N_17199,N_17083,N_17095);
nor U17200 (N_17200,N_16926,N_16812);
and U17201 (N_17201,N_16839,N_16938);
nor U17202 (N_17202,N_16806,N_16878);
or U17203 (N_17203,N_16983,N_16874);
and U17204 (N_17204,N_16900,N_17079);
xor U17205 (N_17205,N_17056,N_17096);
or U17206 (N_17206,N_16807,N_16977);
and U17207 (N_17207,N_16838,N_17088);
nor U17208 (N_17208,N_16999,N_16810);
or U17209 (N_17209,N_17039,N_17027);
and U17210 (N_17210,N_16847,N_17052);
xor U17211 (N_17211,N_16884,N_16850);
nor U17212 (N_17212,N_16876,N_16872);
nor U17213 (N_17213,N_16891,N_17000);
or U17214 (N_17214,N_16862,N_16899);
or U17215 (N_17215,N_16952,N_17028);
nand U17216 (N_17216,N_16857,N_17022);
nand U17217 (N_17217,N_16828,N_17043);
and U17218 (N_17218,N_16841,N_16935);
and U17219 (N_17219,N_17075,N_16949);
nand U17220 (N_17220,N_16910,N_16880);
and U17221 (N_17221,N_16829,N_17049);
xor U17222 (N_17222,N_16918,N_17030);
nand U17223 (N_17223,N_17078,N_17023);
nor U17224 (N_17224,N_16962,N_16883);
and U17225 (N_17225,N_16801,N_16905);
or U17226 (N_17226,N_17037,N_17045);
nor U17227 (N_17227,N_16903,N_17016);
and U17228 (N_17228,N_16822,N_17059);
nand U17229 (N_17229,N_17020,N_16982);
nor U17230 (N_17230,N_17091,N_16858);
and U17231 (N_17231,N_17073,N_17072);
nor U17232 (N_17232,N_16869,N_16947);
xor U17233 (N_17233,N_17074,N_17097);
nand U17234 (N_17234,N_16885,N_16894);
nor U17235 (N_17235,N_16970,N_17036);
nor U17236 (N_17236,N_17009,N_16965);
or U17237 (N_17237,N_16833,N_16809);
nor U17238 (N_17238,N_16940,N_17076);
or U17239 (N_17239,N_16909,N_17069);
xor U17240 (N_17240,N_16824,N_17090);
and U17241 (N_17241,N_16877,N_17004);
nand U17242 (N_17242,N_16871,N_16992);
and U17243 (N_17243,N_16800,N_16818);
nand U17244 (N_17244,N_16989,N_17094);
nand U17245 (N_17245,N_17025,N_17082);
nor U17246 (N_17246,N_16825,N_16832);
nand U17247 (N_17247,N_16966,N_16991);
and U17248 (N_17248,N_17008,N_17018);
and U17249 (N_17249,N_17054,N_16835);
and U17250 (N_17250,N_17064,N_16897);
or U17251 (N_17251,N_16890,N_17094);
nand U17252 (N_17252,N_17088,N_17022);
or U17253 (N_17253,N_16990,N_16867);
or U17254 (N_17254,N_16911,N_16872);
nand U17255 (N_17255,N_17013,N_16943);
nor U17256 (N_17256,N_17028,N_17095);
nand U17257 (N_17257,N_16977,N_16953);
nand U17258 (N_17258,N_17078,N_17065);
nor U17259 (N_17259,N_16823,N_16937);
nor U17260 (N_17260,N_16928,N_16970);
nand U17261 (N_17261,N_17027,N_17046);
nor U17262 (N_17262,N_16916,N_16911);
nor U17263 (N_17263,N_16916,N_17085);
nand U17264 (N_17264,N_16875,N_16953);
or U17265 (N_17265,N_17023,N_16845);
nor U17266 (N_17266,N_16970,N_16923);
and U17267 (N_17267,N_16955,N_16923);
and U17268 (N_17268,N_17016,N_17026);
nor U17269 (N_17269,N_17063,N_16970);
nand U17270 (N_17270,N_16846,N_16927);
nand U17271 (N_17271,N_17095,N_16810);
xnor U17272 (N_17272,N_16894,N_17075);
or U17273 (N_17273,N_16935,N_16834);
nand U17274 (N_17274,N_17079,N_17028);
or U17275 (N_17275,N_16950,N_16922);
and U17276 (N_17276,N_16829,N_16846);
or U17277 (N_17277,N_17034,N_16959);
or U17278 (N_17278,N_16991,N_16891);
and U17279 (N_17279,N_16829,N_16848);
and U17280 (N_17280,N_16974,N_16801);
and U17281 (N_17281,N_16942,N_16900);
nand U17282 (N_17282,N_16994,N_16969);
nor U17283 (N_17283,N_16965,N_17038);
or U17284 (N_17284,N_17013,N_17009);
xor U17285 (N_17285,N_17049,N_16883);
or U17286 (N_17286,N_17034,N_17018);
xor U17287 (N_17287,N_16910,N_16931);
nand U17288 (N_17288,N_16957,N_17091);
or U17289 (N_17289,N_16971,N_16848);
and U17290 (N_17290,N_16918,N_16855);
or U17291 (N_17291,N_16912,N_16981);
nand U17292 (N_17292,N_17059,N_16991);
nor U17293 (N_17293,N_16859,N_17035);
or U17294 (N_17294,N_17086,N_17049);
xor U17295 (N_17295,N_17097,N_17086);
and U17296 (N_17296,N_16956,N_17004);
or U17297 (N_17297,N_17064,N_17003);
xnor U17298 (N_17298,N_16911,N_16980);
and U17299 (N_17299,N_16863,N_16937);
or U17300 (N_17300,N_17036,N_16835);
or U17301 (N_17301,N_17020,N_17058);
nand U17302 (N_17302,N_17029,N_16855);
nor U17303 (N_17303,N_16833,N_16937);
nor U17304 (N_17304,N_16997,N_16939);
xor U17305 (N_17305,N_16920,N_17055);
nor U17306 (N_17306,N_17044,N_17089);
or U17307 (N_17307,N_17006,N_16982);
or U17308 (N_17308,N_16809,N_16900);
nor U17309 (N_17309,N_16819,N_16877);
and U17310 (N_17310,N_17018,N_17022);
or U17311 (N_17311,N_17057,N_16946);
and U17312 (N_17312,N_16858,N_17071);
xnor U17313 (N_17313,N_16955,N_16932);
and U17314 (N_17314,N_17070,N_16942);
nor U17315 (N_17315,N_16966,N_16913);
and U17316 (N_17316,N_16965,N_17083);
xnor U17317 (N_17317,N_16837,N_16935);
nor U17318 (N_17318,N_16966,N_17001);
nor U17319 (N_17319,N_17014,N_17046);
and U17320 (N_17320,N_16973,N_17092);
nand U17321 (N_17321,N_16854,N_16879);
or U17322 (N_17322,N_16860,N_16807);
nand U17323 (N_17323,N_17079,N_16998);
or U17324 (N_17324,N_16841,N_17009);
nor U17325 (N_17325,N_16975,N_16950);
xnor U17326 (N_17326,N_17082,N_16967);
xnor U17327 (N_17327,N_17046,N_17019);
and U17328 (N_17328,N_16862,N_17089);
nand U17329 (N_17329,N_16876,N_16937);
xnor U17330 (N_17330,N_17002,N_16866);
xor U17331 (N_17331,N_17052,N_16852);
nor U17332 (N_17332,N_17087,N_17036);
nor U17333 (N_17333,N_16923,N_16817);
and U17334 (N_17334,N_17043,N_17087);
nor U17335 (N_17335,N_16841,N_16840);
nand U17336 (N_17336,N_17009,N_16901);
xor U17337 (N_17337,N_16801,N_16899);
or U17338 (N_17338,N_17019,N_17040);
nor U17339 (N_17339,N_17008,N_17074);
xnor U17340 (N_17340,N_17042,N_16879);
nor U17341 (N_17341,N_16975,N_16944);
nand U17342 (N_17342,N_17016,N_16978);
or U17343 (N_17343,N_16976,N_16804);
nor U17344 (N_17344,N_16936,N_17090);
xnor U17345 (N_17345,N_17058,N_17055);
or U17346 (N_17346,N_16933,N_16880);
nand U17347 (N_17347,N_17009,N_16999);
nor U17348 (N_17348,N_16960,N_16827);
xnor U17349 (N_17349,N_16976,N_16942);
nor U17350 (N_17350,N_17009,N_16859);
or U17351 (N_17351,N_16814,N_16847);
xor U17352 (N_17352,N_17022,N_16861);
xor U17353 (N_17353,N_17038,N_16852);
xnor U17354 (N_17354,N_16929,N_17022);
and U17355 (N_17355,N_16962,N_16948);
xor U17356 (N_17356,N_16953,N_16962);
or U17357 (N_17357,N_16870,N_17077);
nand U17358 (N_17358,N_17022,N_16997);
nand U17359 (N_17359,N_16817,N_17018);
nand U17360 (N_17360,N_16966,N_17046);
nor U17361 (N_17361,N_16935,N_16813);
nor U17362 (N_17362,N_17049,N_16868);
and U17363 (N_17363,N_16918,N_16967);
nand U17364 (N_17364,N_16986,N_16913);
nand U17365 (N_17365,N_16912,N_17005);
nor U17366 (N_17366,N_16911,N_16975);
nand U17367 (N_17367,N_16979,N_17092);
or U17368 (N_17368,N_16844,N_16971);
and U17369 (N_17369,N_16903,N_16896);
or U17370 (N_17370,N_16860,N_16824);
or U17371 (N_17371,N_17051,N_17007);
and U17372 (N_17372,N_17075,N_17059);
or U17373 (N_17373,N_16839,N_16999);
and U17374 (N_17374,N_17009,N_16982);
or U17375 (N_17375,N_17080,N_17009);
xor U17376 (N_17376,N_17030,N_17065);
and U17377 (N_17377,N_16849,N_16824);
or U17378 (N_17378,N_16891,N_17003);
or U17379 (N_17379,N_16840,N_16848);
or U17380 (N_17380,N_16841,N_17066);
nand U17381 (N_17381,N_16926,N_16935);
and U17382 (N_17382,N_17020,N_16887);
nor U17383 (N_17383,N_16998,N_17025);
nor U17384 (N_17384,N_17068,N_16847);
nor U17385 (N_17385,N_17088,N_16974);
nand U17386 (N_17386,N_17090,N_16918);
nor U17387 (N_17387,N_16845,N_16810);
and U17388 (N_17388,N_17054,N_16888);
nor U17389 (N_17389,N_16841,N_16878);
xnor U17390 (N_17390,N_16824,N_16900);
nand U17391 (N_17391,N_17003,N_17033);
xor U17392 (N_17392,N_17062,N_17092);
nor U17393 (N_17393,N_16800,N_17076);
xnor U17394 (N_17394,N_16861,N_16871);
or U17395 (N_17395,N_17004,N_16833);
nor U17396 (N_17396,N_16901,N_17069);
nor U17397 (N_17397,N_17010,N_17070);
nor U17398 (N_17398,N_16979,N_16857);
xnor U17399 (N_17399,N_16989,N_17019);
nor U17400 (N_17400,N_17274,N_17169);
nor U17401 (N_17401,N_17133,N_17152);
nand U17402 (N_17402,N_17389,N_17178);
xnor U17403 (N_17403,N_17354,N_17368);
or U17404 (N_17404,N_17172,N_17342);
nor U17405 (N_17405,N_17211,N_17275);
and U17406 (N_17406,N_17159,N_17300);
nor U17407 (N_17407,N_17331,N_17106);
nand U17408 (N_17408,N_17265,N_17201);
nor U17409 (N_17409,N_17132,N_17388);
or U17410 (N_17410,N_17234,N_17120);
nor U17411 (N_17411,N_17358,N_17341);
nor U17412 (N_17412,N_17261,N_17314);
nor U17413 (N_17413,N_17279,N_17239);
xnor U17414 (N_17414,N_17303,N_17123);
nor U17415 (N_17415,N_17107,N_17394);
nand U17416 (N_17416,N_17363,N_17174);
xnor U17417 (N_17417,N_17210,N_17127);
and U17418 (N_17418,N_17164,N_17311);
or U17419 (N_17419,N_17166,N_17278);
and U17420 (N_17420,N_17369,N_17187);
nand U17421 (N_17421,N_17301,N_17286);
nor U17422 (N_17422,N_17167,N_17284);
and U17423 (N_17423,N_17141,N_17204);
and U17424 (N_17424,N_17395,N_17380);
or U17425 (N_17425,N_17397,N_17293);
and U17426 (N_17426,N_17245,N_17296);
nand U17427 (N_17427,N_17244,N_17111);
nor U17428 (N_17428,N_17105,N_17387);
and U17429 (N_17429,N_17119,N_17207);
or U17430 (N_17430,N_17113,N_17365);
xnor U17431 (N_17431,N_17154,N_17145);
and U17432 (N_17432,N_17230,N_17103);
xor U17433 (N_17433,N_17128,N_17375);
and U17434 (N_17434,N_17294,N_17143);
nand U17435 (N_17435,N_17112,N_17247);
or U17436 (N_17436,N_17327,N_17243);
or U17437 (N_17437,N_17183,N_17162);
or U17438 (N_17438,N_17147,N_17376);
nand U17439 (N_17439,N_17309,N_17306);
nand U17440 (N_17440,N_17100,N_17281);
xor U17441 (N_17441,N_17260,N_17194);
and U17442 (N_17442,N_17336,N_17248);
nand U17443 (N_17443,N_17351,N_17224);
xor U17444 (N_17444,N_17176,N_17258);
xor U17445 (N_17445,N_17292,N_17372);
or U17446 (N_17446,N_17102,N_17222);
nor U17447 (N_17447,N_17269,N_17209);
and U17448 (N_17448,N_17377,N_17242);
or U17449 (N_17449,N_17285,N_17264);
nand U17450 (N_17450,N_17362,N_17216);
nand U17451 (N_17451,N_17237,N_17116);
nor U17452 (N_17452,N_17257,N_17254);
and U17453 (N_17453,N_17349,N_17228);
nand U17454 (N_17454,N_17195,N_17208);
and U17455 (N_17455,N_17364,N_17339);
and U17456 (N_17456,N_17227,N_17333);
or U17457 (N_17457,N_17393,N_17241);
xnor U17458 (N_17458,N_17280,N_17318);
xnor U17459 (N_17459,N_17315,N_17262);
xor U17460 (N_17460,N_17206,N_17215);
xnor U17461 (N_17461,N_17268,N_17263);
xor U17462 (N_17462,N_17399,N_17348);
nand U17463 (N_17463,N_17151,N_17190);
and U17464 (N_17464,N_17108,N_17383);
or U17465 (N_17465,N_17277,N_17332);
and U17466 (N_17466,N_17193,N_17236);
nor U17467 (N_17467,N_17214,N_17273);
nand U17468 (N_17468,N_17182,N_17197);
nand U17469 (N_17469,N_17140,N_17173);
and U17470 (N_17470,N_17240,N_17334);
xnor U17471 (N_17471,N_17310,N_17370);
and U17472 (N_17472,N_17114,N_17101);
nand U17473 (N_17473,N_17386,N_17287);
or U17474 (N_17474,N_17288,N_17168);
xnor U17475 (N_17475,N_17109,N_17373);
or U17476 (N_17476,N_17199,N_17177);
xor U17477 (N_17477,N_17213,N_17316);
nand U17478 (N_17478,N_17136,N_17171);
and U17479 (N_17479,N_17129,N_17124);
and U17480 (N_17480,N_17104,N_17252);
xor U17481 (N_17481,N_17352,N_17226);
xnor U17482 (N_17482,N_17165,N_17329);
nand U17483 (N_17483,N_17361,N_17320);
nand U17484 (N_17484,N_17192,N_17360);
or U17485 (N_17485,N_17250,N_17188);
nand U17486 (N_17486,N_17139,N_17157);
and U17487 (N_17487,N_17379,N_17312);
nand U17488 (N_17488,N_17282,N_17142);
nor U17489 (N_17489,N_17321,N_17337);
xnor U17490 (N_17490,N_17371,N_17322);
nand U17491 (N_17491,N_17344,N_17367);
or U17492 (N_17492,N_17202,N_17121);
nor U17493 (N_17493,N_17117,N_17200);
nor U17494 (N_17494,N_17153,N_17205);
nand U17495 (N_17495,N_17155,N_17137);
and U17496 (N_17496,N_17156,N_17225);
nand U17497 (N_17497,N_17345,N_17356);
nand U17498 (N_17498,N_17355,N_17196);
and U17499 (N_17499,N_17325,N_17175);
and U17500 (N_17500,N_17125,N_17290);
nand U17501 (N_17501,N_17381,N_17343);
or U17502 (N_17502,N_17346,N_17347);
nor U17503 (N_17503,N_17185,N_17267);
nand U17504 (N_17504,N_17229,N_17272);
and U17505 (N_17505,N_17353,N_17218);
or U17506 (N_17506,N_17256,N_17249);
xnor U17507 (N_17507,N_17251,N_17297);
nand U17508 (N_17508,N_17110,N_17134);
nor U17509 (N_17509,N_17253,N_17259);
xor U17510 (N_17510,N_17289,N_17283);
or U17511 (N_17511,N_17135,N_17323);
xor U17512 (N_17512,N_17305,N_17122);
and U17513 (N_17513,N_17126,N_17392);
nor U17514 (N_17514,N_17130,N_17295);
nand U17515 (N_17515,N_17366,N_17291);
nor U17516 (N_17516,N_17179,N_17181);
xnor U17517 (N_17517,N_17115,N_17138);
xnor U17518 (N_17518,N_17340,N_17160);
or U17519 (N_17519,N_17382,N_17335);
or U17520 (N_17520,N_17231,N_17385);
and U17521 (N_17521,N_17235,N_17203);
nor U17522 (N_17522,N_17299,N_17131);
or U17523 (N_17523,N_17313,N_17238);
xor U17524 (N_17524,N_17170,N_17326);
xnor U17525 (N_17525,N_17118,N_17255);
or U17526 (N_17526,N_17350,N_17357);
nor U17527 (N_17527,N_17319,N_17390);
and U17528 (N_17528,N_17276,N_17223);
or U17529 (N_17529,N_17324,N_17374);
nand U17530 (N_17530,N_17246,N_17271);
xnor U17531 (N_17531,N_17163,N_17391);
xnor U17532 (N_17532,N_17233,N_17219);
xnor U17533 (N_17533,N_17148,N_17270);
nand U17534 (N_17534,N_17317,N_17330);
or U17535 (N_17535,N_17302,N_17180);
nor U17536 (N_17536,N_17232,N_17184);
nor U17537 (N_17537,N_17338,N_17212);
nand U17538 (N_17538,N_17398,N_17359);
xor U17539 (N_17539,N_17396,N_17220);
and U17540 (N_17540,N_17189,N_17221);
and U17541 (N_17541,N_17144,N_17161);
nand U17542 (N_17542,N_17307,N_17191);
or U17543 (N_17543,N_17308,N_17378);
or U17544 (N_17544,N_17304,N_17217);
nor U17545 (N_17545,N_17266,N_17158);
and U17546 (N_17546,N_17149,N_17186);
and U17547 (N_17547,N_17298,N_17146);
and U17548 (N_17548,N_17198,N_17150);
nand U17549 (N_17549,N_17328,N_17384);
xnor U17550 (N_17550,N_17127,N_17204);
nand U17551 (N_17551,N_17101,N_17354);
nand U17552 (N_17552,N_17367,N_17112);
nor U17553 (N_17553,N_17263,N_17134);
xor U17554 (N_17554,N_17114,N_17263);
and U17555 (N_17555,N_17352,N_17277);
and U17556 (N_17556,N_17237,N_17101);
or U17557 (N_17557,N_17373,N_17179);
xor U17558 (N_17558,N_17177,N_17352);
or U17559 (N_17559,N_17259,N_17111);
nand U17560 (N_17560,N_17303,N_17105);
xnor U17561 (N_17561,N_17275,N_17138);
xor U17562 (N_17562,N_17310,N_17329);
xor U17563 (N_17563,N_17117,N_17268);
nand U17564 (N_17564,N_17258,N_17326);
nor U17565 (N_17565,N_17364,N_17159);
or U17566 (N_17566,N_17202,N_17287);
nand U17567 (N_17567,N_17122,N_17338);
or U17568 (N_17568,N_17159,N_17202);
or U17569 (N_17569,N_17159,N_17253);
or U17570 (N_17570,N_17216,N_17285);
and U17571 (N_17571,N_17279,N_17309);
xnor U17572 (N_17572,N_17138,N_17312);
xnor U17573 (N_17573,N_17144,N_17167);
xnor U17574 (N_17574,N_17312,N_17339);
or U17575 (N_17575,N_17376,N_17371);
nand U17576 (N_17576,N_17346,N_17232);
or U17577 (N_17577,N_17295,N_17241);
nor U17578 (N_17578,N_17246,N_17229);
nor U17579 (N_17579,N_17220,N_17279);
and U17580 (N_17580,N_17126,N_17156);
nand U17581 (N_17581,N_17310,N_17224);
xnor U17582 (N_17582,N_17318,N_17334);
or U17583 (N_17583,N_17154,N_17211);
nor U17584 (N_17584,N_17223,N_17194);
nor U17585 (N_17585,N_17308,N_17328);
and U17586 (N_17586,N_17215,N_17130);
and U17587 (N_17587,N_17396,N_17336);
and U17588 (N_17588,N_17103,N_17232);
or U17589 (N_17589,N_17294,N_17108);
xor U17590 (N_17590,N_17110,N_17189);
xor U17591 (N_17591,N_17361,N_17231);
nand U17592 (N_17592,N_17216,N_17106);
nor U17593 (N_17593,N_17135,N_17363);
and U17594 (N_17594,N_17350,N_17150);
and U17595 (N_17595,N_17195,N_17328);
and U17596 (N_17596,N_17165,N_17310);
and U17597 (N_17597,N_17131,N_17204);
or U17598 (N_17598,N_17133,N_17219);
xnor U17599 (N_17599,N_17232,N_17144);
and U17600 (N_17600,N_17126,N_17258);
nand U17601 (N_17601,N_17261,N_17226);
xor U17602 (N_17602,N_17187,N_17118);
nand U17603 (N_17603,N_17315,N_17251);
nand U17604 (N_17604,N_17345,N_17177);
or U17605 (N_17605,N_17310,N_17207);
xor U17606 (N_17606,N_17140,N_17151);
or U17607 (N_17607,N_17218,N_17269);
xnor U17608 (N_17608,N_17343,N_17160);
xor U17609 (N_17609,N_17101,N_17398);
and U17610 (N_17610,N_17187,N_17167);
or U17611 (N_17611,N_17179,N_17272);
xor U17612 (N_17612,N_17332,N_17214);
or U17613 (N_17613,N_17272,N_17386);
nor U17614 (N_17614,N_17348,N_17305);
nor U17615 (N_17615,N_17233,N_17190);
and U17616 (N_17616,N_17328,N_17137);
or U17617 (N_17617,N_17103,N_17130);
and U17618 (N_17618,N_17396,N_17353);
and U17619 (N_17619,N_17274,N_17269);
nand U17620 (N_17620,N_17357,N_17185);
nor U17621 (N_17621,N_17258,N_17321);
and U17622 (N_17622,N_17382,N_17101);
nand U17623 (N_17623,N_17396,N_17182);
and U17624 (N_17624,N_17115,N_17156);
or U17625 (N_17625,N_17395,N_17154);
xor U17626 (N_17626,N_17351,N_17398);
or U17627 (N_17627,N_17174,N_17116);
and U17628 (N_17628,N_17393,N_17262);
xor U17629 (N_17629,N_17350,N_17339);
or U17630 (N_17630,N_17115,N_17232);
and U17631 (N_17631,N_17307,N_17326);
and U17632 (N_17632,N_17214,N_17235);
nor U17633 (N_17633,N_17108,N_17381);
nand U17634 (N_17634,N_17200,N_17266);
xnor U17635 (N_17635,N_17240,N_17241);
and U17636 (N_17636,N_17344,N_17349);
nor U17637 (N_17637,N_17382,N_17354);
or U17638 (N_17638,N_17396,N_17211);
nor U17639 (N_17639,N_17366,N_17386);
xor U17640 (N_17640,N_17317,N_17134);
xnor U17641 (N_17641,N_17372,N_17221);
or U17642 (N_17642,N_17202,N_17171);
nand U17643 (N_17643,N_17255,N_17377);
or U17644 (N_17644,N_17279,N_17194);
nor U17645 (N_17645,N_17292,N_17117);
or U17646 (N_17646,N_17206,N_17273);
xnor U17647 (N_17647,N_17312,N_17223);
or U17648 (N_17648,N_17134,N_17173);
nor U17649 (N_17649,N_17254,N_17386);
xnor U17650 (N_17650,N_17355,N_17103);
and U17651 (N_17651,N_17265,N_17231);
or U17652 (N_17652,N_17248,N_17341);
or U17653 (N_17653,N_17138,N_17186);
xnor U17654 (N_17654,N_17350,N_17157);
or U17655 (N_17655,N_17110,N_17204);
and U17656 (N_17656,N_17361,N_17296);
or U17657 (N_17657,N_17192,N_17322);
and U17658 (N_17658,N_17199,N_17354);
and U17659 (N_17659,N_17332,N_17387);
xnor U17660 (N_17660,N_17392,N_17303);
and U17661 (N_17661,N_17152,N_17149);
nor U17662 (N_17662,N_17250,N_17129);
or U17663 (N_17663,N_17210,N_17172);
or U17664 (N_17664,N_17286,N_17250);
nor U17665 (N_17665,N_17212,N_17330);
nor U17666 (N_17666,N_17390,N_17266);
or U17667 (N_17667,N_17262,N_17399);
nand U17668 (N_17668,N_17334,N_17161);
or U17669 (N_17669,N_17317,N_17357);
and U17670 (N_17670,N_17124,N_17173);
or U17671 (N_17671,N_17238,N_17109);
or U17672 (N_17672,N_17334,N_17226);
xor U17673 (N_17673,N_17370,N_17302);
xor U17674 (N_17674,N_17257,N_17363);
nor U17675 (N_17675,N_17232,N_17215);
xnor U17676 (N_17676,N_17190,N_17166);
nand U17677 (N_17677,N_17209,N_17156);
xor U17678 (N_17678,N_17277,N_17191);
nor U17679 (N_17679,N_17371,N_17140);
nand U17680 (N_17680,N_17174,N_17118);
xnor U17681 (N_17681,N_17166,N_17154);
nor U17682 (N_17682,N_17328,N_17389);
or U17683 (N_17683,N_17256,N_17197);
or U17684 (N_17684,N_17280,N_17388);
and U17685 (N_17685,N_17120,N_17250);
nand U17686 (N_17686,N_17275,N_17288);
and U17687 (N_17687,N_17324,N_17107);
or U17688 (N_17688,N_17291,N_17138);
or U17689 (N_17689,N_17379,N_17157);
nor U17690 (N_17690,N_17168,N_17368);
nand U17691 (N_17691,N_17102,N_17290);
and U17692 (N_17692,N_17302,N_17208);
xnor U17693 (N_17693,N_17200,N_17178);
or U17694 (N_17694,N_17197,N_17360);
xnor U17695 (N_17695,N_17290,N_17208);
xor U17696 (N_17696,N_17394,N_17175);
nand U17697 (N_17697,N_17176,N_17365);
or U17698 (N_17698,N_17176,N_17186);
and U17699 (N_17699,N_17220,N_17298);
nand U17700 (N_17700,N_17637,N_17684);
and U17701 (N_17701,N_17518,N_17657);
or U17702 (N_17702,N_17506,N_17692);
or U17703 (N_17703,N_17580,N_17442);
and U17704 (N_17704,N_17698,N_17455);
and U17705 (N_17705,N_17560,N_17691);
nand U17706 (N_17706,N_17421,N_17630);
nand U17707 (N_17707,N_17429,N_17443);
nand U17708 (N_17708,N_17505,N_17614);
nor U17709 (N_17709,N_17495,N_17496);
and U17710 (N_17710,N_17603,N_17482);
nor U17711 (N_17711,N_17504,N_17563);
and U17712 (N_17712,N_17418,N_17659);
xnor U17713 (N_17713,N_17581,N_17405);
nand U17714 (N_17714,N_17594,N_17669);
xor U17715 (N_17715,N_17400,N_17683);
nor U17716 (N_17716,N_17693,N_17524);
xnor U17717 (N_17717,N_17570,N_17523);
nand U17718 (N_17718,N_17578,N_17522);
nand U17719 (N_17719,N_17648,N_17542);
xor U17720 (N_17720,N_17546,N_17468);
xnor U17721 (N_17721,N_17419,N_17699);
and U17722 (N_17722,N_17626,N_17508);
nor U17723 (N_17723,N_17551,N_17612);
and U17724 (N_17724,N_17574,N_17601);
nand U17725 (N_17725,N_17447,N_17557);
nand U17726 (N_17726,N_17485,N_17410);
and U17727 (N_17727,N_17475,N_17620);
or U17728 (N_17728,N_17463,N_17573);
nor U17729 (N_17729,N_17527,N_17680);
xor U17730 (N_17730,N_17655,N_17685);
or U17731 (N_17731,N_17510,N_17513);
or U17732 (N_17732,N_17634,N_17619);
and U17733 (N_17733,N_17528,N_17424);
nor U17734 (N_17734,N_17583,N_17498);
nor U17735 (N_17735,N_17640,N_17596);
nand U17736 (N_17736,N_17434,N_17458);
and U17737 (N_17737,N_17534,N_17431);
nor U17738 (N_17738,N_17456,N_17571);
nand U17739 (N_17739,N_17449,N_17526);
or U17740 (N_17740,N_17440,N_17582);
and U17741 (N_17741,N_17439,N_17493);
nand U17742 (N_17742,N_17589,N_17519);
xor U17743 (N_17743,N_17535,N_17644);
or U17744 (N_17744,N_17480,N_17432);
and U17745 (N_17745,N_17695,N_17413);
or U17746 (N_17746,N_17552,N_17629);
nand U17747 (N_17747,N_17569,N_17411);
nor U17748 (N_17748,N_17512,N_17478);
nand U17749 (N_17749,N_17517,N_17547);
nand U17750 (N_17750,N_17689,N_17661);
or U17751 (N_17751,N_17651,N_17562);
and U17752 (N_17752,N_17558,N_17672);
nor U17753 (N_17753,N_17445,N_17404);
or U17754 (N_17754,N_17696,N_17401);
xor U17755 (N_17755,N_17617,N_17556);
xor U17756 (N_17756,N_17566,N_17605);
or U17757 (N_17757,N_17467,N_17406);
nor U17758 (N_17758,N_17511,N_17460);
nand U17759 (N_17759,N_17540,N_17476);
and U17760 (N_17760,N_17652,N_17676);
nand U17761 (N_17761,N_17417,N_17464);
xnor U17762 (N_17762,N_17427,N_17670);
nand U17763 (N_17763,N_17587,N_17553);
nor U17764 (N_17764,N_17638,N_17600);
xor U17765 (N_17765,N_17567,N_17687);
nand U17766 (N_17766,N_17621,N_17479);
nor U17767 (N_17767,N_17592,N_17608);
or U17768 (N_17768,N_17470,N_17425);
nand U17769 (N_17769,N_17665,N_17416);
nor U17770 (N_17770,N_17444,N_17446);
nand U17771 (N_17771,N_17533,N_17613);
or U17772 (N_17772,N_17494,N_17525);
nand U17773 (N_17773,N_17541,N_17507);
or U17774 (N_17774,N_17585,N_17466);
nor U17775 (N_17775,N_17635,N_17678);
xor U17776 (N_17776,N_17611,N_17489);
or U17777 (N_17777,N_17453,N_17545);
or U17778 (N_17778,N_17609,N_17591);
xnor U17779 (N_17779,N_17641,N_17666);
nand U17780 (N_17780,N_17572,N_17686);
or U17781 (N_17781,N_17544,N_17515);
and U17782 (N_17782,N_17514,N_17491);
or U17783 (N_17783,N_17653,N_17536);
and U17784 (N_17784,N_17675,N_17658);
and U17785 (N_17785,N_17593,N_17503);
nand U17786 (N_17786,N_17679,N_17428);
nand U17787 (N_17787,N_17462,N_17577);
or U17788 (N_17788,N_17586,N_17632);
xnor U17789 (N_17789,N_17588,N_17697);
nand U17790 (N_17790,N_17636,N_17500);
xnor U17791 (N_17791,N_17615,N_17403);
xnor U17792 (N_17792,N_17576,N_17579);
or U17793 (N_17793,N_17673,N_17465);
xor U17794 (N_17794,N_17667,N_17543);
or U17795 (N_17795,N_17568,N_17663);
nor U17796 (N_17796,N_17477,N_17437);
or U17797 (N_17797,N_17529,N_17471);
and U17798 (N_17798,N_17597,N_17602);
nor U17799 (N_17799,N_17499,N_17627);
nand U17800 (N_17800,N_17438,N_17488);
xnor U17801 (N_17801,N_17481,N_17497);
nor U17802 (N_17802,N_17564,N_17422);
and U17803 (N_17803,N_17414,N_17423);
nor U17804 (N_17804,N_17646,N_17407);
nor U17805 (N_17805,N_17677,N_17625);
and U17806 (N_17806,N_17565,N_17473);
nor U17807 (N_17807,N_17590,N_17509);
or U17808 (N_17808,N_17454,N_17415);
or U17809 (N_17809,N_17457,N_17520);
or U17810 (N_17810,N_17532,N_17674);
nor U17811 (N_17811,N_17610,N_17654);
nand U17812 (N_17812,N_17642,N_17559);
or U17813 (N_17813,N_17486,N_17668);
nand U17814 (N_17814,N_17530,N_17616);
nand U17815 (N_17815,N_17660,N_17452);
and U17816 (N_17816,N_17426,N_17521);
xor U17817 (N_17817,N_17502,N_17549);
nand U17818 (N_17818,N_17682,N_17538);
or U17819 (N_17819,N_17694,N_17474);
xor U17820 (N_17820,N_17555,N_17450);
and U17821 (N_17821,N_17501,N_17575);
or U17822 (N_17822,N_17622,N_17599);
and U17823 (N_17823,N_17435,N_17516);
nor U17824 (N_17824,N_17484,N_17631);
or U17825 (N_17825,N_17671,N_17647);
nand U17826 (N_17826,N_17688,N_17628);
nand U17827 (N_17827,N_17664,N_17490);
or U17828 (N_17828,N_17408,N_17584);
nor U17829 (N_17829,N_17430,N_17420);
nand U17830 (N_17830,N_17409,N_17539);
nor U17831 (N_17831,N_17604,N_17433);
nor U17832 (N_17832,N_17402,N_17607);
and U17833 (N_17833,N_17595,N_17441);
xor U17834 (N_17834,N_17690,N_17487);
or U17835 (N_17835,N_17550,N_17448);
nand U17836 (N_17836,N_17492,N_17461);
and U17837 (N_17837,N_17561,N_17436);
and U17838 (N_17838,N_17412,N_17681);
xnor U17839 (N_17839,N_17606,N_17624);
nand U17840 (N_17840,N_17472,N_17656);
nand U17841 (N_17841,N_17554,N_17531);
or U17842 (N_17842,N_17662,N_17618);
nor U17843 (N_17843,N_17650,N_17643);
xnor U17844 (N_17844,N_17598,N_17649);
nand U17845 (N_17845,N_17639,N_17537);
nor U17846 (N_17846,N_17633,N_17469);
or U17847 (N_17847,N_17623,N_17548);
and U17848 (N_17848,N_17483,N_17451);
or U17849 (N_17849,N_17645,N_17459);
or U17850 (N_17850,N_17438,N_17622);
xor U17851 (N_17851,N_17405,N_17473);
xor U17852 (N_17852,N_17496,N_17693);
nor U17853 (N_17853,N_17634,N_17633);
and U17854 (N_17854,N_17508,N_17660);
and U17855 (N_17855,N_17466,N_17442);
nand U17856 (N_17856,N_17694,N_17578);
xor U17857 (N_17857,N_17483,N_17644);
nor U17858 (N_17858,N_17500,N_17493);
nand U17859 (N_17859,N_17593,N_17636);
and U17860 (N_17860,N_17447,N_17432);
nand U17861 (N_17861,N_17587,N_17684);
and U17862 (N_17862,N_17527,N_17493);
xnor U17863 (N_17863,N_17407,N_17552);
xor U17864 (N_17864,N_17438,N_17672);
nand U17865 (N_17865,N_17667,N_17629);
nor U17866 (N_17866,N_17508,N_17493);
xor U17867 (N_17867,N_17527,N_17448);
or U17868 (N_17868,N_17682,N_17519);
and U17869 (N_17869,N_17423,N_17668);
nor U17870 (N_17870,N_17483,N_17690);
and U17871 (N_17871,N_17697,N_17651);
nand U17872 (N_17872,N_17582,N_17532);
xnor U17873 (N_17873,N_17590,N_17462);
and U17874 (N_17874,N_17577,N_17412);
xor U17875 (N_17875,N_17570,N_17502);
nand U17876 (N_17876,N_17427,N_17402);
xor U17877 (N_17877,N_17677,N_17485);
or U17878 (N_17878,N_17689,N_17496);
nor U17879 (N_17879,N_17582,N_17697);
nor U17880 (N_17880,N_17533,N_17598);
nor U17881 (N_17881,N_17477,N_17440);
xnor U17882 (N_17882,N_17424,N_17697);
nor U17883 (N_17883,N_17425,N_17448);
nor U17884 (N_17884,N_17420,N_17656);
and U17885 (N_17885,N_17601,N_17469);
nor U17886 (N_17886,N_17467,N_17468);
nand U17887 (N_17887,N_17628,N_17695);
nand U17888 (N_17888,N_17464,N_17497);
xnor U17889 (N_17889,N_17514,N_17678);
xor U17890 (N_17890,N_17472,N_17534);
and U17891 (N_17891,N_17642,N_17681);
or U17892 (N_17892,N_17519,N_17529);
nor U17893 (N_17893,N_17457,N_17628);
nor U17894 (N_17894,N_17515,N_17652);
xnor U17895 (N_17895,N_17565,N_17606);
and U17896 (N_17896,N_17685,N_17543);
xnor U17897 (N_17897,N_17652,N_17436);
xor U17898 (N_17898,N_17431,N_17679);
or U17899 (N_17899,N_17644,N_17573);
xor U17900 (N_17900,N_17577,N_17578);
nor U17901 (N_17901,N_17409,N_17541);
xnor U17902 (N_17902,N_17478,N_17614);
nor U17903 (N_17903,N_17631,N_17656);
xor U17904 (N_17904,N_17482,N_17651);
xor U17905 (N_17905,N_17440,N_17590);
and U17906 (N_17906,N_17459,N_17594);
nand U17907 (N_17907,N_17538,N_17582);
and U17908 (N_17908,N_17583,N_17644);
nor U17909 (N_17909,N_17432,N_17426);
nand U17910 (N_17910,N_17504,N_17449);
and U17911 (N_17911,N_17686,N_17600);
nand U17912 (N_17912,N_17543,N_17453);
nor U17913 (N_17913,N_17699,N_17412);
nand U17914 (N_17914,N_17518,N_17532);
nor U17915 (N_17915,N_17513,N_17678);
nor U17916 (N_17916,N_17600,N_17681);
and U17917 (N_17917,N_17521,N_17461);
nor U17918 (N_17918,N_17641,N_17450);
xor U17919 (N_17919,N_17625,N_17429);
or U17920 (N_17920,N_17623,N_17448);
xnor U17921 (N_17921,N_17528,N_17608);
nand U17922 (N_17922,N_17628,N_17654);
xor U17923 (N_17923,N_17684,N_17688);
or U17924 (N_17924,N_17461,N_17454);
nand U17925 (N_17925,N_17480,N_17579);
xor U17926 (N_17926,N_17692,N_17495);
xnor U17927 (N_17927,N_17573,N_17544);
and U17928 (N_17928,N_17495,N_17569);
or U17929 (N_17929,N_17448,N_17502);
or U17930 (N_17930,N_17507,N_17486);
xnor U17931 (N_17931,N_17675,N_17553);
xnor U17932 (N_17932,N_17509,N_17663);
nand U17933 (N_17933,N_17687,N_17621);
nor U17934 (N_17934,N_17509,N_17487);
xnor U17935 (N_17935,N_17553,N_17543);
nor U17936 (N_17936,N_17618,N_17508);
or U17937 (N_17937,N_17626,N_17615);
or U17938 (N_17938,N_17644,N_17410);
or U17939 (N_17939,N_17409,N_17672);
xnor U17940 (N_17940,N_17608,N_17461);
and U17941 (N_17941,N_17524,N_17587);
nand U17942 (N_17942,N_17419,N_17400);
xnor U17943 (N_17943,N_17450,N_17454);
xor U17944 (N_17944,N_17491,N_17455);
and U17945 (N_17945,N_17404,N_17561);
or U17946 (N_17946,N_17670,N_17654);
nor U17947 (N_17947,N_17459,N_17452);
and U17948 (N_17948,N_17425,N_17517);
xor U17949 (N_17949,N_17571,N_17559);
or U17950 (N_17950,N_17607,N_17625);
or U17951 (N_17951,N_17661,N_17698);
xnor U17952 (N_17952,N_17487,N_17637);
and U17953 (N_17953,N_17498,N_17615);
nand U17954 (N_17954,N_17544,N_17448);
and U17955 (N_17955,N_17692,N_17695);
nor U17956 (N_17956,N_17558,N_17444);
and U17957 (N_17957,N_17561,N_17506);
and U17958 (N_17958,N_17482,N_17496);
or U17959 (N_17959,N_17560,N_17505);
xor U17960 (N_17960,N_17573,N_17653);
and U17961 (N_17961,N_17623,N_17699);
xor U17962 (N_17962,N_17496,N_17560);
nor U17963 (N_17963,N_17637,N_17582);
nor U17964 (N_17964,N_17695,N_17503);
or U17965 (N_17965,N_17529,N_17420);
xor U17966 (N_17966,N_17435,N_17642);
and U17967 (N_17967,N_17408,N_17519);
nand U17968 (N_17968,N_17518,N_17604);
xor U17969 (N_17969,N_17633,N_17589);
nand U17970 (N_17970,N_17532,N_17596);
nand U17971 (N_17971,N_17496,N_17471);
nand U17972 (N_17972,N_17697,N_17405);
nand U17973 (N_17973,N_17686,N_17461);
and U17974 (N_17974,N_17610,N_17665);
or U17975 (N_17975,N_17449,N_17673);
nand U17976 (N_17976,N_17602,N_17587);
nand U17977 (N_17977,N_17599,N_17623);
or U17978 (N_17978,N_17511,N_17619);
and U17979 (N_17979,N_17563,N_17465);
or U17980 (N_17980,N_17507,N_17418);
nand U17981 (N_17981,N_17611,N_17533);
xor U17982 (N_17982,N_17403,N_17420);
or U17983 (N_17983,N_17612,N_17555);
or U17984 (N_17984,N_17558,N_17496);
xnor U17985 (N_17985,N_17568,N_17620);
xor U17986 (N_17986,N_17690,N_17671);
nor U17987 (N_17987,N_17517,N_17482);
nor U17988 (N_17988,N_17463,N_17680);
nand U17989 (N_17989,N_17671,N_17499);
nand U17990 (N_17990,N_17633,N_17465);
and U17991 (N_17991,N_17640,N_17409);
and U17992 (N_17992,N_17429,N_17664);
xnor U17993 (N_17993,N_17574,N_17694);
xor U17994 (N_17994,N_17567,N_17575);
nand U17995 (N_17995,N_17417,N_17472);
xor U17996 (N_17996,N_17512,N_17554);
nor U17997 (N_17997,N_17686,N_17513);
nand U17998 (N_17998,N_17633,N_17694);
or U17999 (N_17999,N_17674,N_17609);
and U18000 (N_18000,N_17998,N_17817);
and U18001 (N_18001,N_17831,N_17830);
nand U18002 (N_18002,N_17852,N_17885);
nor U18003 (N_18003,N_17864,N_17874);
xnor U18004 (N_18004,N_17750,N_17819);
xnor U18005 (N_18005,N_17937,N_17707);
or U18006 (N_18006,N_17753,N_17919);
and U18007 (N_18007,N_17785,N_17995);
nand U18008 (N_18008,N_17717,N_17867);
nor U18009 (N_18009,N_17912,N_17795);
nor U18010 (N_18010,N_17964,N_17842);
or U18011 (N_18011,N_17906,N_17732);
or U18012 (N_18012,N_17947,N_17776);
and U18013 (N_18013,N_17837,N_17748);
and U18014 (N_18014,N_17909,N_17975);
nand U18015 (N_18015,N_17738,N_17803);
nor U18016 (N_18016,N_17742,N_17950);
nand U18017 (N_18017,N_17807,N_17915);
nor U18018 (N_18018,N_17706,N_17938);
and U18019 (N_18019,N_17914,N_17815);
nand U18020 (N_18020,N_17703,N_17982);
and U18021 (N_18021,N_17722,N_17930);
xnor U18022 (N_18022,N_17929,N_17812);
nor U18023 (N_18023,N_17756,N_17939);
xnor U18024 (N_18024,N_17701,N_17734);
and U18025 (N_18025,N_17754,N_17956);
xor U18026 (N_18026,N_17926,N_17936);
nand U18027 (N_18027,N_17820,N_17927);
and U18028 (N_18028,N_17871,N_17992);
xor U18029 (N_18029,N_17916,N_17784);
nor U18030 (N_18030,N_17805,N_17743);
or U18031 (N_18031,N_17869,N_17720);
or U18032 (N_18032,N_17882,N_17973);
and U18033 (N_18033,N_17715,N_17994);
xnor U18034 (N_18034,N_17856,N_17941);
or U18035 (N_18035,N_17987,N_17757);
nand U18036 (N_18036,N_17779,N_17758);
or U18037 (N_18037,N_17848,N_17846);
nor U18038 (N_18038,N_17782,N_17902);
or U18039 (N_18039,N_17990,N_17900);
nor U18040 (N_18040,N_17976,N_17872);
or U18041 (N_18041,N_17928,N_17963);
xnor U18042 (N_18042,N_17777,N_17759);
nor U18043 (N_18043,N_17708,N_17770);
nand U18044 (N_18044,N_17955,N_17923);
or U18045 (N_18045,N_17878,N_17739);
nand U18046 (N_18046,N_17797,N_17932);
or U18047 (N_18047,N_17881,N_17769);
or U18048 (N_18048,N_17765,N_17858);
xnor U18049 (N_18049,N_17783,N_17951);
nand U18050 (N_18050,N_17755,N_17724);
or U18051 (N_18051,N_17713,N_17814);
nand U18052 (N_18052,N_17786,N_17723);
and U18053 (N_18053,N_17761,N_17727);
xnor U18054 (N_18054,N_17851,N_17980);
nor U18055 (N_18055,N_17983,N_17752);
and U18056 (N_18056,N_17835,N_17959);
and U18057 (N_18057,N_17935,N_17892);
nand U18058 (N_18058,N_17845,N_17793);
or U18059 (N_18059,N_17823,N_17735);
or U18060 (N_18060,N_17897,N_17711);
nand U18061 (N_18061,N_17808,N_17908);
and U18062 (N_18062,N_17746,N_17799);
nor U18063 (N_18063,N_17953,N_17876);
xnor U18064 (N_18064,N_17904,N_17767);
nor U18065 (N_18065,N_17890,N_17921);
nor U18066 (N_18066,N_17873,N_17850);
xnor U18067 (N_18067,N_17899,N_17917);
nand U18068 (N_18068,N_17824,N_17792);
or U18069 (N_18069,N_17968,N_17828);
and U18070 (N_18070,N_17991,N_17733);
nand U18071 (N_18071,N_17944,N_17967);
nand U18072 (N_18072,N_17969,N_17903);
or U18073 (N_18073,N_17719,N_17996);
nor U18074 (N_18074,N_17868,N_17925);
nand U18075 (N_18075,N_17979,N_17961);
or U18076 (N_18076,N_17787,N_17965);
and U18077 (N_18077,N_17911,N_17714);
nor U18078 (N_18078,N_17788,N_17934);
nand U18079 (N_18079,N_17857,N_17763);
nor U18080 (N_18080,N_17700,N_17918);
nand U18081 (N_18081,N_17806,N_17863);
xor U18082 (N_18082,N_17843,N_17774);
nand U18083 (N_18083,N_17778,N_17811);
or U18084 (N_18084,N_17804,N_17838);
or U18085 (N_18085,N_17762,N_17726);
or U18086 (N_18086,N_17725,N_17833);
and U18087 (N_18087,N_17933,N_17883);
xor U18088 (N_18088,N_17862,N_17839);
nand U18089 (N_18089,N_17721,N_17920);
nand U18090 (N_18090,N_17896,N_17791);
xnor U18091 (N_18091,N_17747,N_17737);
xnor U18092 (N_18092,N_17768,N_17773);
or U18093 (N_18093,N_17854,N_17986);
nor U18094 (N_18094,N_17802,N_17999);
or U18095 (N_18095,N_17859,N_17702);
or U18096 (N_18096,N_17772,N_17977);
nor U18097 (N_18097,N_17891,N_17974);
and U18098 (N_18098,N_17981,N_17741);
or U18099 (N_18099,N_17993,N_17877);
and U18100 (N_18100,N_17905,N_17894);
or U18101 (N_18101,N_17736,N_17841);
nor U18102 (N_18102,N_17948,N_17822);
or U18103 (N_18103,N_17818,N_17718);
nand U18104 (N_18104,N_17710,N_17813);
nor U18105 (N_18105,N_17886,N_17826);
or U18106 (N_18106,N_17730,N_17840);
xor U18107 (N_18107,N_17884,N_17985);
and U18108 (N_18108,N_17960,N_17972);
and U18109 (N_18109,N_17931,N_17962);
nand U18110 (N_18110,N_17870,N_17922);
xor U18111 (N_18111,N_17945,N_17875);
nor U18112 (N_18112,N_17913,N_17866);
nor U18113 (N_18113,N_17888,N_17853);
nor U18114 (N_18114,N_17880,N_17709);
nand U18115 (N_18115,N_17704,N_17834);
or U18116 (N_18116,N_17901,N_17958);
nand U18117 (N_18117,N_17907,N_17957);
or U18118 (N_18118,N_17829,N_17949);
and U18119 (N_18119,N_17832,N_17809);
nor U18120 (N_18120,N_17744,N_17766);
nor U18121 (N_18121,N_17728,N_17849);
nor U18122 (N_18122,N_17895,N_17887);
xnor U18123 (N_18123,N_17751,N_17971);
nor U18124 (N_18124,N_17954,N_17943);
and U18125 (N_18125,N_17889,N_17865);
nor U18126 (N_18126,N_17790,N_17771);
xnor U18127 (N_18127,N_17893,N_17789);
nor U18128 (N_18128,N_17827,N_17940);
nand U18129 (N_18129,N_17796,N_17712);
or U18130 (N_18130,N_17780,N_17910);
nor U18131 (N_18131,N_17924,N_17988);
xnor U18132 (N_18132,N_17800,N_17860);
and U18133 (N_18133,N_17740,N_17821);
xor U18134 (N_18134,N_17997,N_17942);
or U18135 (N_18135,N_17861,N_17952);
nand U18136 (N_18136,N_17855,N_17794);
nand U18137 (N_18137,N_17970,N_17825);
nand U18138 (N_18138,N_17729,N_17984);
nand U18139 (N_18139,N_17946,N_17798);
xnor U18140 (N_18140,N_17716,N_17705);
nor U18141 (N_18141,N_17978,N_17745);
xnor U18142 (N_18142,N_17816,N_17898);
or U18143 (N_18143,N_17879,N_17781);
xnor U18144 (N_18144,N_17966,N_17989);
or U18145 (N_18145,N_17836,N_17749);
xor U18146 (N_18146,N_17801,N_17810);
nand U18147 (N_18147,N_17844,N_17764);
nor U18148 (N_18148,N_17760,N_17775);
nand U18149 (N_18149,N_17731,N_17847);
or U18150 (N_18150,N_17850,N_17735);
nor U18151 (N_18151,N_17853,N_17772);
nor U18152 (N_18152,N_17721,N_17781);
or U18153 (N_18153,N_17855,N_17905);
and U18154 (N_18154,N_17830,N_17727);
xnor U18155 (N_18155,N_17749,N_17854);
or U18156 (N_18156,N_17892,N_17761);
xnor U18157 (N_18157,N_17892,N_17772);
xnor U18158 (N_18158,N_17804,N_17830);
and U18159 (N_18159,N_17799,N_17999);
xnor U18160 (N_18160,N_17733,N_17823);
xnor U18161 (N_18161,N_17854,N_17998);
and U18162 (N_18162,N_17706,N_17928);
or U18163 (N_18163,N_17993,N_17720);
or U18164 (N_18164,N_17723,N_17847);
nand U18165 (N_18165,N_17945,N_17845);
nor U18166 (N_18166,N_17787,N_17953);
xnor U18167 (N_18167,N_17831,N_17750);
and U18168 (N_18168,N_17780,N_17967);
nor U18169 (N_18169,N_17872,N_17705);
and U18170 (N_18170,N_17716,N_17801);
and U18171 (N_18171,N_17894,N_17897);
nand U18172 (N_18172,N_17752,N_17841);
nor U18173 (N_18173,N_17717,N_17902);
and U18174 (N_18174,N_17748,N_17801);
or U18175 (N_18175,N_17753,N_17897);
nand U18176 (N_18176,N_17780,N_17950);
nor U18177 (N_18177,N_17986,N_17727);
or U18178 (N_18178,N_17762,N_17801);
nand U18179 (N_18179,N_17926,N_17835);
nand U18180 (N_18180,N_17786,N_17826);
nand U18181 (N_18181,N_17915,N_17926);
xor U18182 (N_18182,N_17817,N_17787);
or U18183 (N_18183,N_17829,N_17936);
xnor U18184 (N_18184,N_17738,N_17886);
nand U18185 (N_18185,N_17978,N_17739);
or U18186 (N_18186,N_17845,N_17740);
and U18187 (N_18187,N_17870,N_17756);
nor U18188 (N_18188,N_17836,N_17741);
nand U18189 (N_18189,N_17966,N_17918);
and U18190 (N_18190,N_17742,N_17935);
nor U18191 (N_18191,N_17999,N_17727);
xnor U18192 (N_18192,N_17906,N_17809);
nor U18193 (N_18193,N_17838,N_17851);
nor U18194 (N_18194,N_17960,N_17869);
or U18195 (N_18195,N_17801,N_17807);
xnor U18196 (N_18196,N_17963,N_17736);
nor U18197 (N_18197,N_17973,N_17907);
or U18198 (N_18198,N_17921,N_17749);
nand U18199 (N_18199,N_17809,N_17956);
or U18200 (N_18200,N_17993,N_17830);
nand U18201 (N_18201,N_17731,N_17911);
and U18202 (N_18202,N_17792,N_17829);
nor U18203 (N_18203,N_17889,N_17809);
xnor U18204 (N_18204,N_17871,N_17776);
nor U18205 (N_18205,N_17732,N_17841);
or U18206 (N_18206,N_17827,N_17713);
nor U18207 (N_18207,N_17774,N_17946);
or U18208 (N_18208,N_17745,N_17755);
nand U18209 (N_18209,N_17994,N_17938);
or U18210 (N_18210,N_17737,N_17918);
xor U18211 (N_18211,N_17770,N_17847);
and U18212 (N_18212,N_17742,N_17786);
or U18213 (N_18213,N_17837,N_17869);
and U18214 (N_18214,N_17873,N_17762);
nand U18215 (N_18215,N_17956,N_17846);
or U18216 (N_18216,N_17703,N_17797);
nor U18217 (N_18217,N_17744,N_17990);
xor U18218 (N_18218,N_17700,N_17811);
xor U18219 (N_18219,N_17796,N_17763);
nor U18220 (N_18220,N_17756,N_17925);
xor U18221 (N_18221,N_17777,N_17942);
nand U18222 (N_18222,N_17785,N_17812);
nand U18223 (N_18223,N_17701,N_17852);
xnor U18224 (N_18224,N_17828,N_17982);
or U18225 (N_18225,N_17960,N_17734);
nor U18226 (N_18226,N_17988,N_17771);
or U18227 (N_18227,N_17726,N_17801);
or U18228 (N_18228,N_17974,N_17748);
xnor U18229 (N_18229,N_17732,N_17954);
nand U18230 (N_18230,N_17736,N_17749);
nor U18231 (N_18231,N_17919,N_17788);
and U18232 (N_18232,N_17774,N_17898);
nand U18233 (N_18233,N_17806,N_17773);
nor U18234 (N_18234,N_17911,N_17989);
nor U18235 (N_18235,N_17786,N_17801);
nor U18236 (N_18236,N_17857,N_17815);
xnor U18237 (N_18237,N_17723,N_17716);
or U18238 (N_18238,N_17777,N_17733);
and U18239 (N_18239,N_17738,N_17855);
and U18240 (N_18240,N_17960,N_17861);
nor U18241 (N_18241,N_17906,N_17902);
nand U18242 (N_18242,N_17764,N_17751);
nor U18243 (N_18243,N_17717,N_17971);
and U18244 (N_18244,N_17844,N_17707);
and U18245 (N_18245,N_17984,N_17925);
nand U18246 (N_18246,N_17996,N_17709);
nor U18247 (N_18247,N_17837,N_17889);
xnor U18248 (N_18248,N_17903,N_17701);
and U18249 (N_18249,N_17905,N_17997);
xor U18250 (N_18250,N_17721,N_17728);
nand U18251 (N_18251,N_17894,N_17920);
xor U18252 (N_18252,N_17731,N_17908);
or U18253 (N_18253,N_17750,N_17927);
nand U18254 (N_18254,N_17702,N_17891);
xor U18255 (N_18255,N_17993,N_17824);
xnor U18256 (N_18256,N_17921,N_17978);
nand U18257 (N_18257,N_17714,N_17778);
nor U18258 (N_18258,N_17823,N_17700);
and U18259 (N_18259,N_17856,N_17909);
and U18260 (N_18260,N_17897,N_17966);
nor U18261 (N_18261,N_17937,N_17757);
or U18262 (N_18262,N_17781,N_17842);
nor U18263 (N_18263,N_17996,N_17842);
nand U18264 (N_18264,N_17743,N_17781);
and U18265 (N_18265,N_17726,N_17832);
or U18266 (N_18266,N_17729,N_17767);
nor U18267 (N_18267,N_17944,N_17745);
xor U18268 (N_18268,N_17870,N_17960);
nor U18269 (N_18269,N_17956,N_17968);
xor U18270 (N_18270,N_17919,N_17756);
nand U18271 (N_18271,N_17854,N_17924);
nor U18272 (N_18272,N_17715,N_17852);
or U18273 (N_18273,N_17852,N_17955);
or U18274 (N_18274,N_17795,N_17719);
nand U18275 (N_18275,N_17846,N_17843);
nor U18276 (N_18276,N_17980,N_17928);
and U18277 (N_18277,N_17739,N_17897);
or U18278 (N_18278,N_17729,N_17960);
or U18279 (N_18279,N_17905,N_17794);
or U18280 (N_18280,N_17951,N_17772);
or U18281 (N_18281,N_17989,N_17932);
nand U18282 (N_18282,N_17700,N_17991);
nand U18283 (N_18283,N_17986,N_17748);
xnor U18284 (N_18284,N_17937,N_17702);
or U18285 (N_18285,N_17988,N_17734);
nand U18286 (N_18286,N_17794,N_17723);
nor U18287 (N_18287,N_17917,N_17811);
nor U18288 (N_18288,N_17703,N_17823);
nor U18289 (N_18289,N_17898,N_17966);
nor U18290 (N_18290,N_17899,N_17823);
and U18291 (N_18291,N_17955,N_17918);
and U18292 (N_18292,N_17811,N_17786);
or U18293 (N_18293,N_17799,N_17900);
nand U18294 (N_18294,N_17816,N_17741);
nor U18295 (N_18295,N_17912,N_17777);
or U18296 (N_18296,N_17761,N_17869);
or U18297 (N_18297,N_17898,N_17974);
and U18298 (N_18298,N_17879,N_17822);
xnor U18299 (N_18299,N_17830,N_17750);
xnor U18300 (N_18300,N_18269,N_18204);
and U18301 (N_18301,N_18015,N_18068);
nand U18302 (N_18302,N_18261,N_18194);
nand U18303 (N_18303,N_18124,N_18232);
or U18304 (N_18304,N_18205,N_18207);
or U18305 (N_18305,N_18043,N_18198);
xor U18306 (N_18306,N_18127,N_18132);
and U18307 (N_18307,N_18169,N_18137);
nand U18308 (N_18308,N_18123,N_18187);
nor U18309 (N_18309,N_18150,N_18184);
xnor U18310 (N_18310,N_18144,N_18138);
or U18311 (N_18311,N_18271,N_18297);
and U18312 (N_18312,N_18176,N_18029);
xor U18313 (N_18313,N_18088,N_18109);
nand U18314 (N_18314,N_18134,N_18173);
and U18315 (N_18315,N_18285,N_18246);
and U18316 (N_18316,N_18274,N_18027);
xnor U18317 (N_18317,N_18142,N_18094);
nor U18318 (N_18318,N_18133,N_18023);
nand U18319 (N_18319,N_18037,N_18089);
and U18320 (N_18320,N_18103,N_18003);
or U18321 (N_18321,N_18292,N_18146);
or U18322 (N_18322,N_18051,N_18175);
and U18323 (N_18323,N_18046,N_18069);
nor U18324 (N_18324,N_18291,N_18014);
or U18325 (N_18325,N_18226,N_18259);
or U18326 (N_18326,N_18071,N_18136);
and U18327 (N_18327,N_18026,N_18171);
xor U18328 (N_18328,N_18262,N_18155);
and U18329 (N_18329,N_18206,N_18091);
or U18330 (N_18330,N_18202,N_18077);
or U18331 (N_18331,N_18217,N_18076);
or U18332 (N_18332,N_18005,N_18244);
and U18333 (N_18333,N_18122,N_18061);
or U18334 (N_18334,N_18019,N_18036);
or U18335 (N_18335,N_18099,N_18113);
nor U18336 (N_18336,N_18097,N_18240);
xor U18337 (N_18337,N_18209,N_18152);
xnor U18338 (N_18338,N_18108,N_18073);
and U18339 (N_18339,N_18065,N_18273);
or U18340 (N_18340,N_18030,N_18154);
or U18341 (N_18341,N_18256,N_18254);
xor U18342 (N_18342,N_18038,N_18048);
or U18343 (N_18343,N_18060,N_18100);
or U18344 (N_18344,N_18128,N_18252);
nand U18345 (N_18345,N_18234,N_18296);
nor U18346 (N_18346,N_18191,N_18129);
nand U18347 (N_18347,N_18268,N_18018);
and U18348 (N_18348,N_18177,N_18236);
or U18349 (N_18349,N_18057,N_18188);
xor U18350 (N_18350,N_18126,N_18264);
and U18351 (N_18351,N_18238,N_18181);
xnor U18352 (N_18352,N_18096,N_18275);
nor U18353 (N_18353,N_18199,N_18004);
nor U18354 (N_18354,N_18024,N_18280);
or U18355 (N_18355,N_18193,N_18201);
or U18356 (N_18356,N_18286,N_18172);
or U18357 (N_18357,N_18047,N_18075);
nand U18358 (N_18358,N_18016,N_18101);
xor U18359 (N_18359,N_18197,N_18008);
or U18360 (N_18360,N_18167,N_18163);
nand U18361 (N_18361,N_18053,N_18298);
xor U18362 (N_18362,N_18220,N_18118);
xnor U18363 (N_18363,N_18112,N_18162);
xor U18364 (N_18364,N_18074,N_18082);
xnor U18365 (N_18365,N_18230,N_18241);
and U18366 (N_18366,N_18164,N_18042);
xor U18367 (N_18367,N_18165,N_18039);
and U18368 (N_18368,N_18001,N_18010);
nand U18369 (N_18369,N_18151,N_18294);
xnor U18370 (N_18370,N_18235,N_18102);
or U18371 (N_18371,N_18270,N_18145);
nand U18372 (N_18372,N_18125,N_18214);
or U18373 (N_18373,N_18290,N_18179);
nor U18374 (N_18374,N_18227,N_18195);
xnor U18375 (N_18375,N_18277,N_18218);
and U18376 (N_18376,N_18282,N_18224);
nand U18377 (N_18377,N_18260,N_18156);
and U18378 (N_18378,N_18021,N_18272);
nor U18379 (N_18379,N_18006,N_18114);
and U18380 (N_18380,N_18249,N_18013);
nand U18381 (N_18381,N_18295,N_18034);
and U18382 (N_18382,N_18288,N_18093);
or U18383 (N_18383,N_18032,N_18233);
or U18384 (N_18384,N_18095,N_18098);
and U18385 (N_18385,N_18284,N_18157);
nor U18386 (N_18386,N_18067,N_18063);
or U18387 (N_18387,N_18266,N_18168);
and U18388 (N_18388,N_18219,N_18161);
nand U18389 (N_18389,N_18212,N_18033);
xnor U18390 (N_18390,N_18243,N_18178);
nor U18391 (N_18391,N_18009,N_18121);
nor U18392 (N_18392,N_18158,N_18222);
nor U18393 (N_18393,N_18000,N_18225);
and U18394 (N_18394,N_18106,N_18007);
or U18395 (N_18395,N_18017,N_18044);
or U18396 (N_18396,N_18265,N_18031);
xor U18397 (N_18397,N_18041,N_18058);
xor U18398 (N_18398,N_18090,N_18064);
or U18399 (N_18399,N_18131,N_18221);
and U18400 (N_18400,N_18247,N_18054);
xnor U18401 (N_18401,N_18231,N_18130);
nand U18402 (N_18402,N_18159,N_18183);
or U18403 (N_18403,N_18045,N_18251);
or U18404 (N_18404,N_18255,N_18174);
nor U18405 (N_18405,N_18020,N_18080);
xor U18406 (N_18406,N_18012,N_18299);
nand U18407 (N_18407,N_18160,N_18149);
or U18408 (N_18408,N_18115,N_18056);
or U18409 (N_18409,N_18028,N_18186);
xor U18410 (N_18410,N_18283,N_18104);
nand U18411 (N_18411,N_18248,N_18084);
xor U18412 (N_18412,N_18208,N_18229);
nor U18413 (N_18413,N_18223,N_18279);
nand U18414 (N_18414,N_18120,N_18213);
and U18415 (N_18415,N_18141,N_18166);
nand U18416 (N_18416,N_18210,N_18025);
and U18417 (N_18417,N_18135,N_18050);
and U18418 (N_18418,N_18035,N_18228);
nand U18419 (N_18419,N_18140,N_18083);
and U18420 (N_18420,N_18287,N_18148);
xor U18421 (N_18421,N_18022,N_18066);
or U18422 (N_18422,N_18072,N_18062);
or U18423 (N_18423,N_18216,N_18079);
nor U18424 (N_18424,N_18263,N_18002);
nand U18425 (N_18425,N_18293,N_18257);
xnor U18426 (N_18426,N_18147,N_18211);
and U18427 (N_18427,N_18086,N_18107);
and U18428 (N_18428,N_18087,N_18258);
xnor U18429 (N_18429,N_18250,N_18081);
nand U18430 (N_18430,N_18203,N_18052);
nand U18431 (N_18431,N_18105,N_18281);
and U18432 (N_18432,N_18111,N_18215);
nor U18433 (N_18433,N_18117,N_18055);
and U18434 (N_18434,N_18040,N_18170);
or U18435 (N_18435,N_18110,N_18180);
or U18436 (N_18436,N_18182,N_18276);
and U18437 (N_18437,N_18011,N_18245);
or U18438 (N_18438,N_18242,N_18185);
xnor U18439 (N_18439,N_18070,N_18192);
and U18440 (N_18440,N_18289,N_18059);
nor U18441 (N_18441,N_18049,N_18139);
nand U18442 (N_18442,N_18196,N_18092);
or U18443 (N_18443,N_18119,N_18189);
xnor U18444 (N_18444,N_18267,N_18078);
or U18445 (N_18445,N_18278,N_18153);
and U18446 (N_18446,N_18116,N_18085);
or U18447 (N_18447,N_18253,N_18200);
nor U18448 (N_18448,N_18237,N_18190);
nor U18449 (N_18449,N_18239,N_18143);
and U18450 (N_18450,N_18274,N_18128);
nand U18451 (N_18451,N_18024,N_18238);
nand U18452 (N_18452,N_18188,N_18103);
nor U18453 (N_18453,N_18290,N_18004);
or U18454 (N_18454,N_18107,N_18061);
nor U18455 (N_18455,N_18250,N_18267);
nand U18456 (N_18456,N_18102,N_18144);
nand U18457 (N_18457,N_18188,N_18005);
nand U18458 (N_18458,N_18114,N_18293);
xnor U18459 (N_18459,N_18279,N_18298);
nor U18460 (N_18460,N_18115,N_18002);
xor U18461 (N_18461,N_18071,N_18082);
nor U18462 (N_18462,N_18205,N_18021);
and U18463 (N_18463,N_18188,N_18208);
or U18464 (N_18464,N_18194,N_18057);
or U18465 (N_18465,N_18182,N_18237);
nand U18466 (N_18466,N_18093,N_18205);
nor U18467 (N_18467,N_18228,N_18233);
nand U18468 (N_18468,N_18140,N_18018);
nand U18469 (N_18469,N_18143,N_18211);
nand U18470 (N_18470,N_18288,N_18047);
and U18471 (N_18471,N_18141,N_18084);
xnor U18472 (N_18472,N_18087,N_18221);
or U18473 (N_18473,N_18199,N_18105);
and U18474 (N_18474,N_18194,N_18254);
nor U18475 (N_18475,N_18268,N_18170);
xnor U18476 (N_18476,N_18035,N_18291);
and U18477 (N_18477,N_18126,N_18072);
nor U18478 (N_18478,N_18046,N_18210);
nor U18479 (N_18479,N_18139,N_18056);
or U18480 (N_18480,N_18101,N_18172);
nand U18481 (N_18481,N_18199,N_18158);
or U18482 (N_18482,N_18072,N_18152);
nor U18483 (N_18483,N_18241,N_18076);
xor U18484 (N_18484,N_18223,N_18104);
and U18485 (N_18485,N_18106,N_18063);
or U18486 (N_18486,N_18115,N_18193);
nor U18487 (N_18487,N_18283,N_18235);
and U18488 (N_18488,N_18269,N_18008);
and U18489 (N_18489,N_18285,N_18284);
xor U18490 (N_18490,N_18035,N_18169);
or U18491 (N_18491,N_18290,N_18082);
and U18492 (N_18492,N_18074,N_18015);
xor U18493 (N_18493,N_18115,N_18205);
or U18494 (N_18494,N_18117,N_18041);
nand U18495 (N_18495,N_18130,N_18228);
and U18496 (N_18496,N_18116,N_18104);
xor U18497 (N_18497,N_18025,N_18176);
and U18498 (N_18498,N_18276,N_18263);
or U18499 (N_18499,N_18154,N_18189);
or U18500 (N_18500,N_18047,N_18042);
and U18501 (N_18501,N_18059,N_18077);
nand U18502 (N_18502,N_18180,N_18084);
and U18503 (N_18503,N_18007,N_18031);
nor U18504 (N_18504,N_18025,N_18203);
nor U18505 (N_18505,N_18036,N_18262);
xor U18506 (N_18506,N_18285,N_18086);
xnor U18507 (N_18507,N_18003,N_18228);
xor U18508 (N_18508,N_18022,N_18176);
xnor U18509 (N_18509,N_18173,N_18113);
nand U18510 (N_18510,N_18133,N_18019);
nand U18511 (N_18511,N_18101,N_18157);
xnor U18512 (N_18512,N_18022,N_18144);
nor U18513 (N_18513,N_18257,N_18264);
xnor U18514 (N_18514,N_18290,N_18170);
nand U18515 (N_18515,N_18116,N_18160);
nand U18516 (N_18516,N_18123,N_18261);
and U18517 (N_18517,N_18209,N_18166);
nor U18518 (N_18518,N_18230,N_18029);
and U18519 (N_18519,N_18028,N_18083);
and U18520 (N_18520,N_18275,N_18117);
xnor U18521 (N_18521,N_18172,N_18173);
or U18522 (N_18522,N_18065,N_18252);
nor U18523 (N_18523,N_18106,N_18273);
nand U18524 (N_18524,N_18267,N_18097);
nor U18525 (N_18525,N_18226,N_18040);
nand U18526 (N_18526,N_18046,N_18127);
xor U18527 (N_18527,N_18010,N_18220);
and U18528 (N_18528,N_18235,N_18154);
nand U18529 (N_18529,N_18232,N_18186);
and U18530 (N_18530,N_18028,N_18007);
xnor U18531 (N_18531,N_18050,N_18231);
and U18532 (N_18532,N_18047,N_18084);
nor U18533 (N_18533,N_18045,N_18283);
or U18534 (N_18534,N_18294,N_18129);
nand U18535 (N_18535,N_18146,N_18256);
nand U18536 (N_18536,N_18210,N_18231);
or U18537 (N_18537,N_18000,N_18102);
or U18538 (N_18538,N_18255,N_18142);
xnor U18539 (N_18539,N_18049,N_18288);
or U18540 (N_18540,N_18245,N_18292);
nor U18541 (N_18541,N_18071,N_18219);
nor U18542 (N_18542,N_18150,N_18073);
nand U18543 (N_18543,N_18223,N_18033);
and U18544 (N_18544,N_18213,N_18270);
nand U18545 (N_18545,N_18070,N_18034);
or U18546 (N_18546,N_18285,N_18054);
xnor U18547 (N_18547,N_18170,N_18258);
nor U18548 (N_18548,N_18294,N_18099);
and U18549 (N_18549,N_18239,N_18226);
or U18550 (N_18550,N_18229,N_18127);
nor U18551 (N_18551,N_18032,N_18227);
nand U18552 (N_18552,N_18297,N_18228);
or U18553 (N_18553,N_18125,N_18160);
xor U18554 (N_18554,N_18059,N_18256);
nor U18555 (N_18555,N_18024,N_18063);
xnor U18556 (N_18556,N_18019,N_18042);
nor U18557 (N_18557,N_18013,N_18151);
nor U18558 (N_18558,N_18211,N_18085);
xor U18559 (N_18559,N_18279,N_18274);
xor U18560 (N_18560,N_18036,N_18218);
xor U18561 (N_18561,N_18061,N_18111);
nor U18562 (N_18562,N_18208,N_18009);
or U18563 (N_18563,N_18081,N_18075);
or U18564 (N_18564,N_18227,N_18237);
xnor U18565 (N_18565,N_18048,N_18220);
nand U18566 (N_18566,N_18284,N_18238);
and U18567 (N_18567,N_18159,N_18223);
nor U18568 (N_18568,N_18265,N_18055);
nor U18569 (N_18569,N_18073,N_18088);
xnor U18570 (N_18570,N_18054,N_18204);
nor U18571 (N_18571,N_18289,N_18096);
xor U18572 (N_18572,N_18103,N_18058);
xor U18573 (N_18573,N_18221,N_18229);
xor U18574 (N_18574,N_18080,N_18134);
nand U18575 (N_18575,N_18250,N_18070);
xor U18576 (N_18576,N_18165,N_18177);
xnor U18577 (N_18577,N_18189,N_18244);
or U18578 (N_18578,N_18048,N_18244);
nand U18579 (N_18579,N_18253,N_18223);
and U18580 (N_18580,N_18172,N_18071);
or U18581 (N_18581,N_18150,N_18291);
or U18582 (N_18582,N_18086,N_18201);
and U18583 (N_18583,N_18148,N_18216);
nand U18584 (N_18584,N_18243,N_18189);
and U18585 (N_18585,N_18019,N_18050);
nand U18586 (N_18586,N_18151,N_18267);
nand U18587 (N_18587,N_18005,N_18017);
nand U18588 (N_18588,N_18255,N_18251);
nor U18589 (N_18589,N_18229,N_18291);
and U18590 (N_18590,N_18197,N_18086);
xor U18591 (N_18591,N_18132,N_18041);
nand U18592 (N_18592,N_18292,N_18004);
or U18593 (N_18593,N_18010,N_18265);
nand U18594 (N_18594,N_18208,N_18070);
nand U18595 (N_18595,N_18236,N_18287);
and U18596 (N_18596,N_18135,N_18182);
or U18597 (N_18597,N_18173,N_18208);
nand U18598 (N_18598,N_18103,N_18294);
nand U18599 (N_18599,N_18125,N_18275);
nor U18600 (N_18600,N_18378,N_18484);
nor U18601 (N_18601,N_18511,N_18341);
and U18602 (N_18602,N_18317,N_18590);
xnor U18603 (N_18603,N_18561,N_18486);
or U18604 (N_18604,N_18455,N_18438);
xor U18605 (N_18605,N_18475,N_18539);
or U18606 (N_18606,N_18565,N_18540);
xor U18607 (N_18607,N_18366,N_18570);
or U18608 (N_18608,N_18593,N_18535);
xnor U18609 (N_18609,N_18333,N_18300);
nor U18610 (N_18610,N_18571,N_18458);
and U18611 (N_18611,N_18301,N_18356);
nand U18612 (N_18612,N_18547,N_18493);
nor U18613 (N_18613,N_18360,N_18574);
or U18614 (N_18614,N_18367,N_18418);
and U18615 (N_18615,N_18572,N_18477);
and U18616 (N_18616,N_18435,N_18414);
and U18617 (N_18617,N_18334,N_18454);
nor U18618 (N_18618,N_18501,N_18421);
and U18619 (N_18619,N_18448,N_18498);
and U18620 (N_18620,N_18546,N_18329);
and U18621 (N_18621,N_18401,N_18453);
xor U18622 (N_18622,N_18528,N_18372);
or U18623 (N_18623,N_18507,N_18550);
xnor U18624 (N_18624,N_18504,N_18588);
xnor U18625 (N_18625,N_18568,N_18405);
or U18626 (N_18626,N_18383,N_18524);
and U18627 (N_18627,N_18361,N_18464);
xnor U18628 (N_18628,N_18312,N_18375);
nand U18629 (N_18629,N_18388,N_18362);
or U18630 (N_18630,N_18575,N_18434);
nor U18631 (N_18631,N_18488,N_18577);
nand U18632 (N_18632,N_18440,N_18363);
nand U18633 (N_18633,N_18496,N_18479);
nand U18634 (N_18634,N_18542,N_18393);
nor U18635 (N_18635,N_18328,N_18397);
or U18636 (N_18636,N_18323,N_18324);
xnor U18637 (N_18637,N_18558,N_18519);
nor U18638 (N_18638,N_18555,N_18514);
or U18639 (N_18639,N_18553,N_18599);
nor U18640 (N_18640,N_18340,N_18306);
xnor U18641 (N_18641,N_18441,N_18564);
nand U18642 (N_18642,N_18410,N_18580);
xor U18643 (N_18643,N_18344,N_18512);
or U18644 (N_18644,N_18469,N_18552);
and U18645 (N_18645,N_18569,N_18303);
and U18646 (N_18646,N_18487,N_18389);
xor U18647 (N_18647,N_18497,N_18338);
nand U18648 (N_18648,N_18499,N_18374);
and U18649 (N_18649,N_18373,N_18357);
nor U18650 (N_18650,N_18415,N_18359);
xnor U18651 (N_18651,N_18473,N_18581);
xnor U18652 (N_18652,N_18330,N_18355);
nor U18653 (N_18653,N_18520,N_18460);
or U18654 (N_18654,N_18489,N_18591);
nor U18655 (N_18655,N_18308,N_18320);
nand U18656 (N_18656,N_18457,N_18508);
or U18657 (N_18657,N_18480,N_18560);
and U18658 (N_18658,N_18326,N_18380);
xnor U18659 (N_18659,N_18398,N_18534);
or U18660 (N_18660,N_18381,N_18402);
or U18661 (N_18661,N_18428,N_18382);
nor U18662 (N_18662,N_18545,N_18567);
nor U18663 (N_18663,N_18364,N_18439);
and U18664 (N_18664,N_18468,N_18331);
nand U18665 (N_18665,N_18379,N_18307);
or U18666 (N_18666,N_18387,N_18302);
or U18667 (N_18667,N_18327,N_18465);
or U18668 (N_18668,N_18598,N_18490);
nand U18669 (N_18669,N_18530,N_18304);
and U18670 (N_18670,N_18482,N_18597);
xnor U18671 (N_18671,N_18573,N_18370);
and U18672 (N_18672,N_18502,N_18579);
and U18673 (N_18673,N_18583,N_18335);
and U18674 (N_18674,N_18517,N_18495);
or U18675 (N_18675,N_18523,N_18400);
or U18676 (N_18676,N_18436,N_18551);
and U18677 (N_18677,N_18423,N_18339);
xor U18678 (N_18678,N_18509,N_18314);
nor U18679 (N_18679,N_18549,N_18424);
and U18680 (N_18680,N_18527,N_18466);
nand U18681 (N_18681,N_18399,N_18521);
and U18682 (N_18682,N_18538,N_18369);
nor U18683 (N_18683,N_18596,N_18316);
xnor U18684 (N_18684,N_18510,N_18322);
nand U18685 (N_18685,N_18492,N_18313);
nand U18686 (N_18686,N_18345,N_18406);
xor U18687 (N_18687,N_18557,N_18472);
or U18688 (N_18688,N_18420,N_18587);
nand U18689 (N_18689,N_18430,N_18595);
nor U18690 (N_18690,N_18503,N_18445);
and U18691 (N_18691,N_18544,N_18347);
nand U18692 (N_18692,N_18404,N_18315);
nor U18693 (N_18693,N_18516,N_18525);
or U18694 (N_18694,N_18478,N_18522);
xor U18695 (N_18695,N_18485,N_18442);
or U18696 (N_18696,N_18470,N_18491);
nor U18697 (N_18697,N_18319,N_18461);
or U18698 (N_18698,N_18385,N_18513);
nand U18699 (N_18699,N_18377,N_18518);
nor U18700 (N_18700,N_18505,N_18589);
xor U18701 (N_18701,N_18433,N_18395);
nor U18702 (N_18702,N_18417,N_18529);
and U18703 (N_18703,N_18451,N_18346);
xor U18704 (N_18704,N_18443,N_18407);
nor U18705 (N_18705,N_18576,N_18321);
or U18706 (N_18706,N_18358,N_18427);
and U18707 (N_18707,N_18337,N_18390);
or U18708 (N_18708,N_18408,N_18449);
xnor U18709 (N_18709,N_18419,N_18531);
or U18710 (N_18710,N_18467,N_18586);
and U18711 (N_18711,N_18559,N_18350);
and U18712 (N_18712,N_18474,N_18594);
and U18713 (N_18713,N_18309,N_18409);
xor U18714 (N_18714,N_18376,N_18543);
or U18715 (N_18715,N_18343,N_18500);
nand U18716 (N_18716,N_18578,N_18584);
and U18717 (N_18717,N_18450,N_18463);
nand U18718 (N_18718,N_18471,N_18348);
and U18719 (N_18719,N_18332,N_18452);
or U18720 (N_18720,N_18305,N_18310);
and U18721 (N_18721,N_18533,N_18563);
xnor U18722 (N_18722,N_18566,N_18476);
and U18723 (N_18723,N_18368,N_18365);
nor U18724 (N_18724,N_18392,N_18311);
or U18725 (N_18725,N_18352,N_18429);
and U18726 (N_18726,N_18411,N_18462);
nand U18727 (N_18727,N_18384,N_18532);
nor U18728 (N_18728,N_18554,N_18426);
or U18729 (N_18729,N_18562,N_18592);
and U18730 (N_18730,N_18351,N_18541);
xor U18731 (N_18731,N_18481,N_18342);
and U18732 (N_18732,N_18459,N_18354);
nand U18733 (N_18733,N_18396,N_18536);
nand U18734 (N_18734,N_18391,N_18548);
or U18735 (N_18735,N_18371,N_18437);
nand U18736 (N_18736,N_18412,N_18494);
xor U18737 (N_18737,N_18353,N_18444);
nand U18738 (N_18738,N_18556,N_18336);
nor U18739 (N_18739,N_18422,N_18537);
or U18740 (N_18740,N_18582,N_18506);
xor U18741 (N_18741,N_18349,N_18403);
xnor U18742 (N_18742,N_18432,N_18585);
nor U18743 (N_18743,N_18425,N_18526);
nor U18744 (N_18744,N_18325,N_18386);
nand U18745 (N_18745,N_18394,N_18416);
or U18746 (N_18746,N_18446,N_18447);
nor U18747 (N_18747,N_18483,N_18431);
nand U18748 (N_18748,N_18515,N_18413);
or U18749 (N_18749,N_18456,N_18318);
and U18750 (N_18750,N_18561,N_18492);
or U18751 (N_18751,N_18515,N_18571);
or U18752 (N_18752,N_18586,N_18583);
or U18753 (N_18753,N_18426,N_18301);
or U18754 (N_18754,N_18551,N_18529);
xnor U18755 (N_18755,N_18565,N_18490);
or U18756 (N_18756,N_18337,N_18459);
nor U18757 (N_18757,N_18420,N_18348);
and U18758 (N_18758,N_18452,N_18438);
xor U18759 (N_18759,N_18552,N_18324);
or U18760 (N_18760,N_18311,N_18424);
or U18761 (N_18761,N_18338,N_18431);
nor U18762 (N_18762,N_18590,N_18356);
or U18763 (N_18763,N_18514,N_18534);
xnor U18764 (N_18764,N_18433,N_18467);
nor U18765 (N_18765,N_18535,N_18492);
xor U18766 (N_18766,N_18335,N_18300);
and U18767 (N_18767,N_18331,N_18462);
xnor U18768 (N_18768,N_18582,N_18451);
nand U18769 (N_18769,N_18408,N_18454);
xnor U18770 (N_18770,N_18524,N_18512);
or U18771 (N_18771,N_18499,N_18300);
nor U18772 (N_18772,N_18373,N_18516);
xor U18773 (N_18773,N_18493,N_18361);
or U18774 (N_18774,N_18383,N_18432);
and U18775 (N_18775,N_18429,N_18551);
and U18776 (N_18776,N_18455,N_18433);
nor U18777 (N_18777,N_18519,N_18561);
nor U18778 (N_18778,N_18553,N_18393);
nor U18779 (N_18779,N_18566,N_18407);
or U18780 (N_18780,N_18582,N_18349);
nor U18781 (N_18781,N_18377,N_18559);
and U18782 (N_18782,N_18330,N_18417);
nand U18783 (N_18783,N_18444,N_18489);
and U18784 (N_18784,N_18501,N_18458);
nor U18785 (N_18785,N_18460,N_18519);
xor U18786 (N_18786,N_18501,N_18452);
and U18787 (N_18787,N_18529,N_18304);
nor U18788 (N_18788,N_18370,N_18533);
nor U18789 (N_18789,N_18447,N_18436);
and U18790 (N_18790,N_18515,N_18421);
xnor U18791 (N_18791,N_18343,N_18318);
or U18792 (N_18792,N_18430,N_18411);
nand U18793 (N_18793,N_18356,N_18326);
nor U18794 (N_18794,N_18477,N_18504);
nor U18795 (N_18795,N_18510,N_18501);
nor U18796 (N_18796,N_18596,N_18405);
xor U18797 (N_18797,N_18576,N_18324);
nor U18798 (N_18798,N_18385,N_18330);
xor U18799 (N_18799,N_18513,N_18444);
nand U18800 (N_18800,N_18354,N_18557);
and U18801 (N_18801,N_18403,N_18504);
and U18802 (N_18802,N_18314,N_18466);
xor U18803 (N_18803,N_18595,N_18526);
nor U18804 (N_18804,N_18452,N_18399);
nand U18805 (N_18805,N_18309,N_18575);
nor U18806 (N_18806,N_18551,N_18307);
and U18807 (N_18807,N_18379,N_18301);
or U18808 (N_18808,N_18351,N_18374);
or U18809 (N_18809,N_18467,N_18360);
or U18810 (N_18810,N_18428,N_18345);
and U18811 (N_18811,N_18353,N_18336);
xor U18812 (N_18812,N_18477,N_18525);
xor U18813 (N_18813,N_18321,N_18375);
nor U18814 (N_18814,N_18349,N_18307);
nand U18815 (N_18815,N_18422,N_18404);
xor U18816 (N_18816,N_18493,N_18442);
and U18817 (N_18817,N_18550,N_18383);
xnor U18818 (N_18818,N_18586,N_18354);
nor U18819 (N_18819,N_18331,N_18378);
nor U18820 (N_18820,N_18445,N_18556);
nand U18821 (N_18821,N_18326,N_18344);
and U18822 (N_18822,N_18595,N_18498);
and U18823 (N_18823,N_18594,N_18385);
nor U18824 (N_18824,N_18322,N_18508);
and U18825 (N_18825,N_18599,N_18350);
and U18826 (N_18826,N_18495,N_18313);
nor U18827 (N_18827,N_18575,N_18501);
nor U18828 (N_18828,N_18454,N_18592);
and U18829 (N_18829,N_18389,N_18441);
nand U18830 (N_18830,N_18434,N_18527);
nand U18831 (N_18831,N_18487,N_18403);
xor U18832 (N_18832,N_18378,N_18489);
nor U18833 (N_18833,N_18442,N_18465);
xnor U18834 (N_18834,N_18345,N_18366);
xor U18835 (N_18835,N_18511,N_18571);
xnor U18836 (N_18836,N_18319,N_18514);
or U18837 (N_18837,N_18562,N_18437);
xnor U18838 (N_18838,N_18406,N_18487);
and U18839 (N_18839,N_18508,N_18516);
or U18840 (N_18840,N_18516,N_18560);
nor U18841 (N_18841,N_18504,N_18414);
nor U18842 (N_18842,N_18596,N_18573);
nor U18843 (N_18843,N_18504,N_18502);
xnor U18844 (N_18844,N_18350,N_18375);
or U18845 (N_18845,N_18306,N_18454);
xnor U18846 (N_18846,N_18448,N_18575);
nand U18847 (N_18847,N_18440,N_18391);
and U18848 (N_18848,N_18336,N_18528);
nand U18849 (N_18849,N_18469,N_18324);
and U18850 (N_18850,N_18481,N_18376);
or U18851 (N_18851,N_18525,N_18424);
nand U18852 (N_18852,N_18500,N_18572);
nor U18853 (N_18853,N_18511,N_18574);
xor U18854 (N_18854,N_18596,N_18400);
xor U18855 (N_18855,N_18592,N_18468);
nand U18856 (N_18856,N_18485,N_18511);
or U18857 (N_18857,N_18534,N_18319);
xor U18858 (N_18858,N_18531,N_18597);
or U18859 (N_18859,N_18337,N_18345);
nand U18860 (N_18860,N_18502,N_18328);
or U18861 (N_18861,N_18359,N_18469);
or U18862 (N_18862,N_18362,N_18453);
and U18863 (N_18863,N_18445,N_18447);
nor U18864 (N_18864,N_18435,N_18407);
or U18865 (N_18865,N_18568,N_18366);
nor U18866 (N_18866,N_18451,N_18385);
nor U18867 (N_18867,N_18517,N_18573);
nor U18868 (N_18868,N_18395,N_18451);
nor U18869 (N_18869,N_18454,N_18431);
nand U18870 (N_18870,N_18305,N_18491);
or U18871 (N_18871,N_18446,N_18373);
and U18872 (N_18872,N_18479,N_18527);
nand U18873 (N_18873,N_18394,N_18510);
and U18874 (N_18874,N_18356,N_18462);
nor U18875 (N_18875,N_18589,N_18330);
or U18876 (N_18876,N_18469,N_18319);
xnor U18877 (N_18877,N_18352,N_18459);
nand U18878 (N_18878,N_18474,N_18331);
and U18879 (N_18879,N_18557,N_18318);
and U18880 (N_18880,N_18586,N_18571);
nor U18881 (N_18881,N_18306,N_18553);
and U18882 (N_18882,N_18531,N_18495);
nand U18883 (N_18883,N_18446,N_18559);
and U18884 (N_18884,N_18478,N_18414);
and U18885 (N_18885,N_18475,N_18471);
and U18886 (N_18886,N_18482,N_18365);
or U18887 (N_18887,N_18542,N_18312);
xnor U18888 (N_18888,N_18351,N_18334);
nand U18889 (N_18889,N_18482,N_18321);
nor U18890 (N_18890,N_18389,N_18556);
and U18891 (N_18891,N_18572,N_18479);
and U18892 (N_18892,N_18584,N_18376);
xnor U18893 (N_18893,N_18310,N_18560);
nor U18894 (N_18894,N_18325,N_18558);
xnor U18895 (N_18895,N_18447,N_18334);
and U18896 (N_18896,N_18458,N_18536);
nor U18897 (N_18897,N_18463,N_18401);
or U18898 (N_18898,N_18569,N_18513);
or U18899 (N_18899,N_18524,N_18531);
and U18900 (N_18900,N_18806,N_18851);
nand U18901 (N_18901,N_18721,N_18757);
nand U18902 (N_18902,N_18655,N_18882);
nor U18903 (N_18903,N_18801,N_18672);
nor U18904 (N_18904,N_18862,N_18724);
nor U18905 (N_18905,N_18636,N_18787);
xor U18906 (N_18906,N_18855,N_18758);
xnor U18907 (N_18907,N_18684,N_18830);
nor U18908 (N_18908,N_18641,N_18698);
nand U18909 (N_18909,N_18844,N_18867);
xor U18910 (N_18910,N_18891,N_18837);
nand U18911 (N_18911,N_18709,N_18642);
nor U18912 (N_18912,N_18826,N_18768);
nand U18913 (N_18913,N_18663,N_18648);
and U18914 (N_18914,N_18870,N_18835);
and U18915 (N_18915,N_18649,N_18689);
or U18916 (N_18916,N_18853,N_18734);
or U18917 (N_18917,N_18866,N_18736);
nand U18918 (N_18918,N_18739,N_18679);
xor U18919 (N_18919,N_18833,N_18859);
nand U18920 (N_18920,N_18681,N_18693);
nor U18921 (N_18921,N_18717,N_18883);
nor U18922 (N_18922,N_18817,N_18659);
nand U18923 (N_18923,N_18700,N_18623);
nor U18924 (N_18924,N_18701,N_18605);
nand U18925 (N_18925,N_18857,N_18720);
nand U18926 (N_18926,N_18621,N_18687);
nor U18927 (N_18927,N_18827,N_18874);
or U18928 (N_18928,N_18766,N_18619);
nor U18929 (N_18929,N_18873,N_18706);
xnor U18930 (N_18930,N_18751,N_18645);
or U18931 (N_18931,N_18775,N_18601);
nand U18932 (N_18932,N_18617,N_18776);
and U18933 (N_18933,N_18748,N_18676);
or U18934 (N_18934,N_18887,N_18694);
and U18935 (N_18935,N_18633,N_18761);
nor U18936 (N_18936,N_18695,N_18781);
xor U18937 (N_18937,N_18732,N_18777);
nor U18938 (N_18938,N_18746,N_18860);
or U18939 (N_18939,N_18772,N_18750);
or U18940 (N_18940,N_18666,N_18795);
or U18941 (N_18941,N_18635,N_18865);
nor U18942 (N_18942,N_18823,N_18712);
xor U18943 (N_18943,N_18728,N_18760);
nand U18944 (N_18944,N_18847,N_18697);
xor U18945 (N_18945,N_18869,N_18639);
and U18946 (N_18946,N_18618,N_18799);
nor U18947 (N_18947,N_18626,N_18685);
nor U18948 (N_18948,N_18754,N_18767);
and U18949 (N_18949,N_18638,N_18811);
or U18950 (N_18950,N_18771,N_18843);
nor U18951 (N_18951,N_18731,N_18778);
nor U18952 (N_18952,N_18877,N_18825);
and U18953 (N_18953,N_18670,N_18674);
and U18954 (N_18954,N_18861,N_18890);
and U18955 (N_18955,N_18699,N_18790);
nor U18956 (N_18956,N_18752,N_18682);
nand U18957 (N_18957,N_18840,N_18856);
and U18958 (N_18958,N_18664,N_18667);
xor U18959 (N_18959,N_18640,N_18714);
nand U18960 (N_18960,N_18646,N_18722);
nor U18961 (N_18961,N_18846,N_18774);
or U18962 (N_18962,N_18675,N_18730);
xnor U18963 (N_18963,N_18669,N_18763);
nor U18964 (N_18964,N_18749,N_18885);
nand U18965 (N_18965,N_18602,N_18872);
nor U18966 (N_18966,N_18807,N_18785);
and U18967 (N_18967,N_18654,N_18610);
nor U18968 (N_18968,N_18686,N_18688);
nor U18969 (N_18969,N_18824,N_18741);
xnor U18970 (N_18970,N_18719,N_18813);
and U18971 (N_18971,N_18707,N_18634);
and U18972 (N_18972,N_18651,N_18703);
or U18973 (N_18973,N_18899,N_18660);
or U18974 (N_18974,N_18880,N_18747);
or U18975 (N_18975,N_18845,N_18756);
or U18976 (N_18976,N_18783,N_18611);
nor U18977 (N_18977,N_18710,N_18737);
nand U18978 (N_18978,N_18692,N_18662);
xnor U18979 (N_18979,N_18656,N_18759);
or U18980 (N_18980,N_18897,N_18627);
or U18981 (N_18981,N_18613,N_18744);
and U18982 (N_18982,N_18755,N_18793);
nand U18983 (N_18983,N_18852,N_18839);
and U18984 (N_18984,N_18821,N_18604);
or U18985 (N_18985,N_18632,N_18650);
and U18986 (N_18986,N_18735,N_18643);
nor U18987 (N_18987,N_18784,N_18624);
nor U18988 (N_18988,N_18832,N_18849);
xor U18989 (N_18989,N_18716,N_18644);
xor U18990 (N_18990,N_18796,N_18616);
xnor U18991 (N_18991,N_18657,N_18665);
xor U18992 (N_18992,N_18765,N_18745);
or U18993 (N_18993,N_18671,N_18858);
or U18994 (N_18994,N_18863,N_18895);
nand U18995 (N_18995,N_18727,N_18678);
xor U18996 (N_18996,N_18898,N_18854);
or U18997 (N_18997,N_18888,N_18808);
nor U18998 (N_18998,N_18889,N_18810);
or U18999 (N_18999,N_18612,N_18805);
nor U19000 (N_19000,N_18705,N_18600);
nand U19001 (N_19001,N_18875,N_18715);
or U19002 (N_19002,N_18892,N_18871);
and U19003 (N_19003,N_18628,N_18708);
nand U19004 (N_19004,N_18631,N_18615);
nand U19005 (N_19005,N_18668,N_18803);
xnor U19006 (N_19006,N_18637,N_18658);
or U19007 (N_19007,N_18702,N_18723);
xnor U19008 (N_19008,N_18828,N_18896);
nor U19009 (N_19009,N_18680,N_18725);
nor U19010 (N_19010,N_18886,N_18786);
and U19011 (N_19011,N_18809,N_18622);
and U19012 (N_19012,N_18794,N_18652);
xnor U19013 (N_19013,N_18677,N_18729);
nor U19014 (N_19014,N_18738,N_18743);
xor U19015 (N_19015,N_18673,N_18822);
and U19016 (N_19016,N_18893,N_18726);
or U19017 (N_19017,N_18630,N_18881);
or U19018 (N_19018,N_18647,N_18802);
nor U19019 (N_19019,N_18780,N_18798);
and U19020 (N_19020,N_18829,N_18620);
nand U19021 (N_19021,N_18814,N_18789);
nand U19022 (N_19022,N_18764,N_18713);
xor U19023 (N_19023,N_18608,N_18762);
and U19024 (N_19024,N_18603,N_18607);
or U19025 (N_19025,N_18683,N_18816);
nand U19026 (N_19026,N_18812,N_18797);
and U19027 (N_19027,N_18614,N_18606);
nand U19028 (N_19028,N_18791,N_18848);
nand U19029 (N_19029,N_18773,N_18879);
nor U19030 (N_19030,N_18850,N_18769);
nor U19031 (N_19031,N_18696,N_18704);
or U19032 (N_19032,N_18629,N_18834);
xor U19033 (N_19033,N_18718,N_18876);
or U19034 (N_19034,N_18884,N_18878);
nand U19035 (N_19035,N_18818,N_18804);
or U19036 (N_19036,N_18820,N_18864);
or U19037 (N_19037,N_18661,N_18841);
and U19038 (N_19038,N_18711,N_18753);
nor U19039 (N_19039,N_18625,N_18831);
or U19040 (N_19040,N_18838,N_18782);
xor U19041 (N_19041,N_18690,N_18609);
or U19042 (N_19042,N_18894,N_18800);
nor U19043 (N_19043,N_18788,N_18733);
nand U19044 (N_19044,N_18691,N_18815);
nor U19045 (N_19045,N_18792,N_18842);
or U19046 (N_19046,N_18740,N_18770);
nor U19047 (N_19047,N_18819,N_18742);
or U19048 (N_19048,N_18779,N_18653);
nand U19049 (N_19049,N_18836,N_18868);
nand U19050 (N_19050,N_18671,N_18794);
nor U19051 (N_19051,N_18702,N_18747);
or U19052 (N_19052,N_18648,N_18608);
nor U19053 (N_19053,N_18726,N_18688);
xnor U19054 (N_19054,N_18653,N_18752);
nand U19055 (N_19055,N_18803,N_18881);
or U19056 (N_19056,N_18643,N_18881);
and U19057 (N_19057,N_18868,N_18837);
and U19058 (N_19058,N_18877,N_18726);
and U19059 (N_19059,N_18666,N_18713);
nand U19060 (N_19060,N_18651,N_18699);
nor U19061 (N_19061,N_18623,N_18874);
or U19062 (N_19062,N_18836,N_18630);
nand U19063 (N_19063,N_18619,N_18716);
nor U19064 (N_19064,N_18878,N_18773);
and U19065 (N_19065,N_18756,N_18795);
xor U19066 (N_19066,N_18862,N_18647);
xnor U19067 (N_19067,N_18827,N_18772);
or U19068 (N_19068,N_18826,N_18712);
xnor U19069 (N_19069,N_18801,N_18688);
or U19070 (N_19070,N_18678,N_18664);
nand U19071 (N_19071,N_18681,N_18804);
or U19072 (N_19072,N_18602,N_18863);
nor U19073 (N_19073,N_18833,N_18719);
or U19074 (N_19074,N_18620,N_18826);
or U19075 (N_19075,N_18893,N_18809);
xor U19076 (N_19076,N_18605,N_18792);
and U19077 (N_19077,N_18801,N_18765);
or U19078 (N_19078,N_18846,N_18887);
or U19079 (N_19079,N_18660,N_18736);
or U19080 (N_19080,N_18816,N_18768);
nand U19081 (N_19081,N_18848,N_18637);
xor U19082 (N_19082,N_18693,N_18855);
nor U19083 (N_19083,N_18657,N_18808);
xor U19084 (N_19084,N_18770,N_18676);
nand U19085 (N_19085,N_18684,N_18743);
xor U19086 (N_19086,N_18736,N_18877);
or U19087 (N_19087,N_18851,N_18875);
nand U19088 (N_19088,N_18784,N_18678);
and U19089 (N_19089,N_18784,N_18862);
xor U19090 (N_19090,N_18674,N_18878);
or U19091 (N_19091,N_18707,N_18855);
or U19092 (N_19092,N_18704,N_18660);
or U19093 (N_19093,N_18741,N_18757);
or U19094 (N_19094,N_18624,N_18701);
xnor U19095 (N_19095,N_18846,N_18603);
xnor U19096 (N_19096,N_18713,N_18812);
or U19097 (N_19097,N_18833,N_18722);
and U19098 (N_19098,N_18711,N_18787);
xor U19099 (N_19099,N_18736,N_18672);
nor U19100 (N_19100,N_18793,N_18640);
nor U19101 (N_19101,N_18671,N_18646);
nand U19102 (N_19102,N_18785,N_18637);
and U19103 (N_19103,N_18825,N_18657);
xnor U19104 (N_19104,N_18625,N_18644);
and U19105 (N_19105,N_18621,N_18872);
and U19106 (N_19106,N_18619,N_18715);
nor U19107 (N_19107,N_18842,N_18835);
nor U19108 (N_19108,N_18635,N_18604);
xor U19109 (N_19109,N_18732,N_18803);
xor U19110 (N_19110,N_18774,N_18811);
nand U19111 (N_19111,N_18781,N_18849);
nand U19112 (N_19112,N_18807,N_18782);
xor U19113 (N_19113,N_18813,N_18686);
xor U19114 (N_19114,N_18612,N_18701);
nand U19115 (N_19115,N_18798,N_18819);
nor U19116 (N_19116,N_18625,N_18712);
nor U19117 (N_19117,N_18640,N_18858);
xor U19118 (N_19118,N_18632,N_18881);
or U19119 (N_19119,N_18660,N_18871);
or U19120 (N_19120,N_18694,N_18899);
xnor U19121 (N_19121,N_18676,N_18695);
nand U19122 (N_19122,N_18696,N_18885);
nor U19123 (N_19123,N_18896,N_18745);
or U19124 (N_19124,N_18661,N_18894);
nor U19125 (N_19125,N_18667,N_18722);
nor U19126 (N_19126,N_18800,N_18832);
xor U19127 (N_19127,N_18782,N_18661);
and U19128 (N_19128,N_18712,N_18650);
nor U19129 (N_19129,N_18727,N_18890);
nand U19130 (N_19130,N_18729,N_18892);
or U19131 (N_19131,N_18655,N_18699);
and U19132 (N_19132,N_18810,N_18801);
or U19133 (N_19133,N_18618,N_18829);
xor U19134 (N_19134,N_18893,N_18706);
nand U19135 (N_19135,N_18688,N_18689);
nor U19136 (N_19136,N_18738,N_18679);
or U19137 (N_19137,N_18827,N_18830);
or U19138 (N_19138,N_18878,N_18756);
xor U19139 (N_19139,N_18738,N_18889);
and U19140 (N_19140,N_18847,N_18727);
nand U19141 (N_19141,N_18652,N_18838);
and U19142 (N_19142,N_18616,N_18691);
or U19143 (N_19143,N_18843,N_18783);
nor U19144 (N_19144,N_18812,N_18897);
nand U19145 (N_19145,N_18761,N_18863);
and U19146 (N_19146,N_18804,N_18796);
and U19147 (N_19147,N_18682,N_18828);
xor U19148 (N_19148,N_18629,N_18784);
xor U19149 (N_19149,N_18693,N_18609);
and U19150 (N_19150,N_18680,N_18889);
xnor U19151 (N_19151,N_18794,N_18795);
nor U19152 (N_19152,N_18893,N_18627);
and U19153 (N_19153,N_18828,N_18808);
nand U19154 (N_19154,N_18847,N_18859);
and U19155 (N_19155,N_18670,N_18876);
or U19156 (N_19156,N_18646,N_18811);
xnor U19157 (N_19157,N_18813,N_18601);
nand U19158 (N_19158,N_18884,N_18835);
xnor U19159 (N_19159,N_18614,N_18748);
or U19160 (N_19160,N_18647,N_18651);
xnor U19161 (N_19161,N_18611,N_18839);
nand U19162 (N_19162,N_18693,N_18722);
or U19163 (N_19163,N_18801,N_18745);
nor U19164 (N_19164,N_18728,N_18813);
nand U19165 (N_19165,N_18619,N_18791);
xor U19166 (N_19166,N_18812,N_18772);
nor U19167 (N_19167,N_18602,N_18603);
or U19168 (N_19168,N_18610,N_18765);
xor U19169 (N_19169,N_18683,N_18715);
nand U19170 (N_19170,N_18666,N_18851);
nor U19171 (N_19171,N_18672,N_18601);
nand U19172 (N_19172,N_18744,N_18716);
or U19173 (N_19173,N_18748,N_18864);
or U19174 (N_19174,N_18628,N_18779);
nor U19175 (N_19175,N_18692,N_18808);
nand U19176 (N_19176,N_18886,N_18896);
or U19177 (N_19177,N_18648,N_18873);
and U19178 (N_19178,N_18877,N_18849);
nor U19179 (N_19179,N_18844,N_18655);
xor U19180 (N_19180,N_18800,N_18699);
or U19181 (N_19181,N_18688,N_18802);
or U19182 (N_19182,N_18675,N_18770);
and U19183 (N_19183,N_18650,N_18772);
or U19184 (N_19184,N_18707,N_18731);
and U19185 (N_19185,N_18877,N_18632);
xnor U19186 (N_19186,N_18785,N_18672);
nor U19187 (N_19187,N_18730,N_18852);
nand U19188 (N_19188,N_18826,N_18854);
nor U19189 (N_19189,N_18678,N_18680);
or U19190 (N_19190,N_18694,N_18772);
and U19191 (N_19191,N_18730,N_18842);
nand U19192 (N_19192,N_18629,N_18799);
nor U19193 (N_19193,N_18730,N_18869);
nor U19194 (N_19194,N_18816,N_18896);
nor U19195 (N_19195,N_18677,N_18775);
or U19196 (N_19196,N_18680,N_18687);
nor U19197 (N_19197,N_18688,N_18644);
and U19198 (N_19198,N_18884,N_18662);
and U19199 (N_19199,N_18785,N_18643);
xor U19200 (N_19200,N_19146,N_19162);
nand U19201 (N_19201,N_19054,N_18995);
and U19202 (N_19202,N_19108,N_18976);
nand U19203 (N_19203,N_19104,N_19190);
xnor U19204 (N_19204,N_18913,N_19094);
xor U19205 (N_19205,N_19121,N_19082);
nor U19206 (N_19206,N_19112,N_19167);
nand U19207 (N_19207,N_19182,N_19010);
xnor U19208 (N_19208,N_19083,N_19175);
nor U19209 (N_19209,N_19067,N_18960);
or U19210 (N_19210,N_18981,N_19140);
and U19211 (N_19211,N_18907,N_18967);
nand U19212 (N_19212,N_19030,N_18991);
nor U19213 (N_19213,N_18997,N_19169);
nand U19214 (N_19214,N_19038,N_18935);
or U19215 (N_19215,N_18923,N_18987);
and U19216 (N_19216,N_19195,N_18980);
or U19217 (N_19217,N_19143,N_18944);
nor U19218 (N_19218,N_19034,N_19022);
xnor U19219 (N_19219,N_19168,N_19124);
or U19220 (N_19220,N_19062,N_19046);
and U19221 (N_19221,N_19047,N_19078);
or U19222 (N_19222,N_19120,N_18945);
nor U19223 (N_19223,N_18956,N_19107);
nand U19224 (N_19224,N_19081,N_19187);
nand U19225 (N_19225,N_19127,N_19123);
or U19226 (N_19226,N_18916,N_18977);
and U19227 (N_19227,N_19184,N_19070);
or U19228 (N_19228,N_19171,N_19088);
or U19229 (N_19229,N_18912,N_18921);
xnor U19230 (N_19230,N_19045,N_19065);
xnor U19231 (N_19231,N_19024,N_18920);
nand U19232 (N_19232,N_19136,N_18958);
nor U19233 (N_19233,N_19141,N_18904);
or U19234 (N_19234,N_19178,N_19037);
nor U19235 (N_19235,N_18950,N_18910);
and U19236 (N_19236,N_18905,N_19019);
or U19237 (N_19237,N_19007,N_19192);
or U19238 (N_19238,N_18983,N_19051);
nor U19239 (N_19239,N_18943,N_18900);
and U19240 (N_19240,N_18909,N_19059);
nor U19241 (N_19241,N_19170,N_19092);
nand U19242 (N_19242,N_19036,N_18911);
or U19243 (N_19243,N_18954,N_19027);
and U19244 (N_19244,N_19134,N_19096);
xnor U19245 (N_19245,N_18924,N_19110);
nand U19246 (N_19246,N_18988,N_19157);
and U19247 (N_19247,N_19023,N_18902);
or U19248 (N_19248,N_19125,N_19117);
and U19249 (N_19249,N_19011,N_19166);
nand U19250 (N_19250,N_18928,N_18964);
or U19251 (N_19251,N_19183,N_19197);
and U19252 (N_19252,N_19016,N_19032);
or U19253 (N_19253,N_19149,N_18972);
nand U19254 (N_19254,N_19164,N_19105);
nor U19255 (N_19255,N_19189,N_19041);
or U19256 (N_19256,N_18970,N_19111);
nor U19257 (N_19257,N_18949,N_18940);
and U19258 (N_19258,N_19151,N_19172);
and U19259 (N_19259,N_19133,N_19100);
and U19260 (N_19260,N_19020,N_19072);
nor U19261 (N_19261,N_19028,N_19147);
nor U19262 (N_19262,N_18927,N_18971);
nand U19263 (N_19263,N_18986,N_19040);
nand U19264 (N_19264,N_18925,N_19014);
or U19265 (N_19265,N_19013,N_18975);
nand U19266 (N_19266,N_18959,N_19050);
nor U19267 (N_19267,N_19057,N_19017);
nand U19268 (N_19268,N_18951,N_19074);
and U19269 (N_19269,N_19031,N_18998);
nand U19270 (N_19270,N_18941,N_19130);
or U19271 (N_19271,N_19185,N_19090);
nand U19272 (N_19272,N_19077,N_19179);
and U19273 (N_19273,N_18989,N_18901);
nor U19274 (N_19274,N_19139,N_19085);
nor U19275 (N_19275,N_19132,N_19152);
nand U19276 (N_19276,N_19091,N_19015);
xor U19277 (N_19277,N_19196,N_19122);
xor U19278 (N_19278,N_18952,N_18965);
xnor U19279 (N_19279,N_18906,N_18938);
and U19280 (N_19280,N_19076,N_19048);
and U19281 (N_19281,N_19115,N_19001);
nor U19282 (N_19282,N_19069,N_18985);
or U19283 (N_19283,N_18946,N_18919);
nor U19284 (N_19284,N_18937,N_19089);
nand U19285 (N_19285,N_18966,N_19003);
nor U19286 (N_19286,N_19118,N_19116);
nand U19287 (N_19287,N_19060,N_19165);
nand U19288 (N_19288,N_19005,N_19018);
nand U19289 (N_19289,N_19021,N_19042);
xor U19290 (N_19290,N_19066,N_19061);
nor U19291 (N_19291,N_19075,N_19145);
and U19292 (N_19292,N_19012,N_19154);
xor U19293 (N_19293,N_18973,N_19153);
nand U19294 (N_19294,N_19039,N_18918);
nor U19295 (N_19295,N_19173,N_19064);
or U19296 (N_19296,N_19102,N_19002);
or U19297 (N_19297,N_19073,N_18930);
nand U19298 (N_19298,N_19155,N_18982);
nand U19299 (N_19299,N_19071,N_18974);
or U19300 (N_19300,N_18926,N_19160);
nor U19301 (N_19301,N_18969,N_19159);
and U19302 (N_19302,N_19161,N_19079);
xor U19303 (N_19303,N_19137,N_18994);
or U19304 (N_19304,N_19158,N_19186);
or U19305 (N_19305,N_19063,N_18934);
nor U19306 (N_19306,N_19029,N_18963);
or U19307 (N_19307,N_19087,N_19098);
nor U19308 (N_19308,N_18903,N_19177);
or U19309 (N_19309,N_18915,N_19000);
xor U19310 (N_19310,N_19086,N_19114);
nand U19311 (N_19311,N_18984,N_19058);
or U19312 (N_19312,N_18957,N_19056);
and U19313 (N_19313,N_18996,N_19095);
nor U19314 (N_19314,N_19055,N_19135);
xor U19315 (N_19315,N_19199,N_19053);
nand U19316 (N_19316,N_18999,N_18968);
xnor U19317 (N_19317,N_19043,N_19128);
nor U19318 (N_19318,N_19138,N_19101);
and U19319 (N_19319,N_19193,N_18979);
and U19320 (N_19320,N_18936,N_19148);
or U19321 (N_19321,N_19049,N_18955);
nor U19322 (N_19322,N_18939,N_19093);
nor U19323 (N_19323,N_19194,N_18931);
and U19324 (N_19324,N_19176,N_19119);
xor U19325 (N_19325,N_19142,N_18992);
nand U19326 (N_19326,N_19033,N_19180);
nand U19327 (N_19327,N_19188,N_18990);
nand U19328 (N_19328,N_19191,N_19084);
nor U19329 (N_19329,N_19126,N_18932);
nor U19330 (N_19330,N_19174,N_19044);
and U19331 (N_19331,N_18922,N_18953);
and U19332 (N_19332,N_18947,N_19144);
xnor U19333 (N_19333,N_19035,N_19103);
and U19334 (N_19334,N_19106,N_18933);
nand U19335 (N_19335,N_19131,N_19129);
xor U19336 (N_19336,N_18962,N_19068);
nor U19337 (N_19337,N_19026,N_19163);
or U19338 (N_19338,N_18978,N_19006);
or U19339 (N_19339,N_19004,N_18942);
nand U19340 (N_19340,N_18908,N_18929);
xor U19341 (N_19341,N_18961,N_19109);
nor U19342 (N_19342,N_19080,N_19025);
and U19343 (N_19343,N_19008,N_18948);
nand U19344 (N_19344,N_19181,N_19099);
nor U19345 (N_19345,N_19097,N_19113);
nor U19346 (N_19346,N_18917,N_19198);
nor U19347 (N_19347,N_19150,N_19009);
nor U19348 (N_19348,N_19156,N_18993);
nand U19349 (N_19349,N_18914,N_19052);
nor U19350 (N_19350,N_19162,N_18987);
nand U19351 (N_19351,N_19077,N_19094);
xor U19352 (N_19352,N_19174,N_19154);
and U19353 (N_19353,N_19008,N_19023);
xnor U19354 (N_19354,N_18905,N_19041);
and U19355 (N_19355,N_18992,N_19168);
and U19356 (N_19356,N_19031,N_19071);
nand U19357 (N_19357,N_19142,N_18951);
xor U19358 (N_19358,N_19065,N_19086);
nand U19359 (N_19359,N_19010,N_19026);
nor U19360 (N_19360,N_18926,N_18931);
xor U19361 (N_19361,N_19185,N_19101);
or U19362 (N_19362,N_19043,N_19172);
xor U19363 (N_19363,N_18940,N_18992);
nor U19364 (N_19364,N_19118,N_19124);
nand U19365 (N_19365,N_18910,N_18956);
xor U19366 (N_19366,N_19136,N_18922);
nand U19367 (N_19367,N_18989,N_19018);
xnor U19368 (N_19368,N_18928,N_19009);
xnor U19369 (N_19369,N_19129,N_19134);
nand U19370 (N_19370,N_19048,N_19033);
nand U19371 (N_19371,N_18976,N_18986);
nor U19372 (N_19372,N_19125,N_19162);
nor U19373 (N_19373,N_18928,N_19005);
xor U19374 (N_19374,N_19119,N_19033);
xnor U19375 (N_19375,N_19027,N_18999);
xnor U19376 (N_19376,N_19075,N_19036);
nor U19377 (N_19377,N_19169,N_19050);
nand U19378 (N_19378,N_19106,N_19037);
nand U19379 (N_19379,N_18970,N_19166);
nor U19380 (N_19380,N_19197,N_18989);
xnor U19381 (N_19381,N_19170,N_18907);
or U19382 (N_19382,N_19109,N_19045);
or U19383 (N_19383,N_19020,N_19130);
nand U19384 (N_19384,N_19086,N_19121);
nor U19385 (N_19385,N_19143,N_19018);
nand U19386 (N_19386,N_19180,N_19058);
xor U19387 (N_19387,N_19194,N_19154);
nand U19388 (N_19388,N_19019,N_19027);
nand U19389 (N_19389,N_19023,N_18970);
and U19390 (N_19390,N_19038,N_18977);
nand U19391 (N_19391,N_18965,N_19099);
nand U19392 (N_19392,N_19104,N_18906);
nand U19393 (N_19393,N_18916,N_19074);
nand U19394 (N_19394,N_19000,N_18912);
nand U19395 (N_19395,N_19102,N_18901);
nor U19396 (N_19396,N_19102,N_18919);
xnor U19397 (N_19397,N_18905,N_18955);
or U19398 (N_19398,N_19130,N_18987);
or U19399 (N_19399,N_18942,N_19018);
xnor U19400 (N_19400,N_18912,N_19140);
nor U19401 (N_19401,N_18909,N_19075);
and U19402 (N_19402,N_19158,N_18984);
xnor U19403 (N_19403,N_18973,N_19173);
nor U19404 (N_19404,N_19078,N_19137);
nor U19405 (N_19405,N_18952,N_19101);
nor U19406 (N_19406,N_19063,N_19107);
nor U19407 (N_19407,N_19186,N_19141);
xor U19408 (N_19408,N_19089,N_19017);
nand U19409 (N_19409,N_18919,N_19156);
xnor U19410 (N_19410,N_18922,N_19032);
xor U19411 (N_19411,N_19196,N_19043);
and U19412 (N_19412,N_18968,N_19079);
nor U19413 (N_19413,N_19066,N_19058);
nand U19414 (N_19414,N_19060,N_19063);
nor U19415 (N_19415,N_18903,N_18912);
xnor U19416 (N_19416,N_19035,N_19126);
xor U19417 (N_19417,N_19008,N_19162);
nand U19418 (N_19418,N_19124,N_19161);
xnor U19419 (N_19419,N_18966,N_19052);
and U19420 (N_19420,N_19137,N_18972);
nor U19421 (N_19421,N_18901,N_19014);
nand U19422 (N_19422,N_19041,N_19090);
xnor U19423 (N_19423,N_18901,N_19099);
nor U19424 (N_19424,N_19076,N_19077);
nand U19425 (N_19425,N_19091,N_19038);
or U19426 (N_19426,N_19092,N_19166);
nand U19427 (N_19427,N_19001,N_19162);
or U19428 (N_19428,N_19137,N_19101);
and U19429 (N_19429,N_19171,N_18981);
or U19430 (N_19430,N_19149,N_18933);
or U19431 (N_19431,N_19169,N_19018);
and U19432 (N_19432,N_19170,N_19175);
or U19433 (N_19433,N_19151,N_18901);
and U19434 (N_19434,N_19104,N_18910);
or U19435 (N_19435,N_19011,N_18994);
nand U19436 (N_19436,N_19175,N_18987);
and U19437 (N_19437,N_19153,N_18992);
nor U19438 (N_19438,N_19179,N_19096);
and U19439 (N_19439,N_19157,N_18972);
or U19440 (N_19440,N_19030,N_19005);
nand U19441 (N_19441,N_19088,N_19110);
nand U19442 (N_19442,N_19135,N_18952);
nor U19443 (N_19443,N_18974,N_19111);
nor U19444 (N_19444,N_18902,N_18905);
xnor U19445 (N_19445,N_19011,N_19147);
and U19446 (N_19446,N_19140,N_18968);
or U19447 (N_19447,N_18985,N_19014);
or U19448 (N_19448,N_19110,N_18915);
nor U19449 (N_19449,N_18950,N_19043);
nand U19450 (N_19450,N_18969,N_19172);
xor U19451 (N_19451,N_19012,N_19004);
nand U19452 (N_19452,N_19047,N_18922);
nand U19453 (N_19453,N_19068,N_19143);
nor U19454 (N_19454,N_19103,N_18945);
nand U19455 (N_19455,N_19163,N_19043);
nand U19456 (N_19456,N_19171,N_19192);
or U19457 (N_19457,N_19048,N_19113);
and U19458 (N_19458,N_19127,N_19065);
xnor U19459 (N_19459,N_19076,N_19173);
nor U19460 (N_19460,N_18974,N_19018);
or U19461 (N_19461,N_19079,N_18982);
nor U19462 (N_19462,N_19146,N_18966);
or U19463 (N_19463,N_18994,N_19189);
xnor U19464 (N_19464,N_19041,N_18999);
xor U19465 (N_19465,N_18922,N_19008);
nor U19466 (N_19466,N_19034,N_19054);
nor U19467 (N_19467,N_19048,N_18926);
nand U19468 (N_19468,N_19081,N_18941);
xnor U19469 (N_19469,N_19089,N_18912);
nor U19470 (N_19470,N_18935,N_18927);
or U19471 (N_19471,N_19047,N_19019);
or U19472 (N_19472,N_19095,N_18990);
nor U19473 (N_19473,N_19005,N_19171);
nor U19474 (N_19474,N_19086,N_19081);
or U19475 (N_19475,N_19095,N_18963);
xnor U19476 (N_19476,N_19135,N_19117);
and U19477 (N_19477,N_19174,N_19034);
xor U19478 (N_19478,N_19032,N_18956);
nor U19479 (N_19479,N_19122,N_19092);
nand U19480 (N_19480,N_19000,N_19080);
or U19481 (N_19481,N_18943,N_18930);
and U19482 (N_19482,N_18961,N_19042);
and U19483 (N_19483,N_19199,N_18987);
nor U19484 (N_19484,N_18961,N_19169);
nor U19485 (N_19485,N_18955,N_19038);
nor U19486 (N_19486,N_19012,N_19108);
nand U19487 (N_19487,N_19172,N_18976);
and U19488 (N_19488,N_18918,N_19137);
and U19489 (N_19489,N_19035,N_19045);
nand U19490 (N_19490,N_19137,N_19017);
xnor U19491 (N_19491,N_19170,N_18936);
or U19492 (N_19492,N_18974,N_18986);
nand U19493 (N_19493,N_19189,N_19015);
or U19494 (N_19494,N_18918,N_19070);
nand U19495 (N_19495,N_19175,N_18939);
or U19496 (N_19496,N_19009,N_19191);
xor U19497 (N_19497,N_19018,N_19183);
xor U19498 (N_19498,N_18966,N_19030);
nand U19499 (N_19499,N_18989,N_18931);
and U19500 (N_19500,N_19488,N_19279);
nor U19501 (N_19501,N_19366,N_19411);
nand U19502 (N_19502,N_19478,N_19328);
and U19503 (N_19503,N_19445,N_19368);
and U19504 (N_19504,N_19305,N_19281);
and U19505 (N_19505,N_19342,N_19285);
or U19506 (N_19506,N_19341,N_19270);
nand U19507 (N_19507,N_19431,N_19485);
nand U19508 (N_19508,N_19472,N_19425);
nor U19509 (N_19509,N_19336,N_19467);
or U19510 (N_19510,N_19493,N_19477);
or U19511 (N_19511,N_19350,N_19400);
xor U19512 (N_19512,N_19399,N_19294);
and U19513 (N_19513,N_19422,N_19345);
xnor U19514 (N_19514,N_19450,N_19359);
nor U19515 (N_19515,N_19401,N_19297);
nor U19516 (N_19516,N_19409,N_19358);
nand U19517 (N_19517,N_19417,N_19239);
xor U19518 (N_19518,N_19241,N_19206);
or U19519 (N_19519,N_19267,N_19248);
or U19520 (N_19520,N_19448,N_19339);
xor U19521 (N_19521,N_19338,N_19288);
nand U19522 (N_19522,N_19362,N_19455);
xnor U19523 (N_19523,N_19429,N_19262);
xnor U19524 (N_19524,N_19250,N_19302);
or U19525 (N_19525,N_19233,N_19352);
nor U19526 (N_19526,N_19218,N_19363);
xnor U19527 (N_19527,N_19325,N_19443);
or U19528 (N_19528,N_19230,N_19377);
nand U19529 (N_19529,N_19433,N_19404);
nor U19530 (N_19530,N_19437,N_19249);
nor U19531 (N_19531,N_19292,N_19231);
nor U19532 (N_19532,N_19474,N_19462);
nand U19533 (N_19533,N_19286,N_19290);
and U19534 (N_19534,N_19298,N_19200);
and U19535 (N_19535,N_19313,N_19322);
xor U19536 (N_19536,N_19211,N_19309);
and U19537 (N_19537,N_19390,N_19441);
nand U19538 (N_19538,N_19215,N_19349);
xor U19539 (N_19539,N_19255,N_19293);
nand U19540 (N_19540,N_19329,N_19348);
xnor U19541 (N_19541,N_19266,N_19224);
xnor U19542 (N_19542,N_19291,N_19436);
nand U19543 (N_19543,N_19439,N_19407);
or U19544 (N_19544,N_19387,N_19303);
or U19545 (N_19545,N_19227,N_19376);
xor U19546 (N_19546,N_19383,N_19419);
nor U19547 (N_19547,N_19269,N_19463);
or U19548 (N_19548,N_19316,N_19415);
or U19549 (N_19549,N_19259,N_19347);
or U19550 (N_19550,N_19207,N_19274);
nor U19551 (N_19551,N_19413,N_19337);
or U19552 (N_19552,N_19476,N_19395);
xnor U19553 (N_19553,N_19213,N_19382);
or U19554 (N_19554,N_19310,N_19226);
nor U19555 (N_19555,N_19311,N_19278);
nor U19556 (N_19556,N_19331,N_19289);
nand U19557 (N_19557,N_19217,N_19205);
xor U19558 (N_19558,N_19497,N_19396);
xor U19559 (N_19559,N_19287,N_19466);
or U19560 (N_19560,N_19464,N_19410);
and U19561 (N_19561,N_19457,N_19388);
and U19562 (N_19562,N_19458,N_19499);
or U19563 (N_19563,N_19452,N_19245);
xnor U19564 (N_19564,N_19364,N_19204);
nand U19565 (N_19565,N_19451,N_19494);
and U19566 (N_19566,N_19475,N_19263);
and U19567 (N_19567,N_19228,N_19386);
or U19568 (N_19568,N_19375,N_19384);
or U19569 (N_19569,N_19210,N_19496);
xnor U19570 (N_19570,N_19421,N_19324);
nand U19571 (N_19571,N_19299,N_19238);
or U19572 (N_19572,N_19470,N_19276);
or U19573 (N_19573,N_19481,N_19357);
nand U19574 (N_19574,N_19371,N_19402);
or U19575 (N_19575,N_19237,N_19435);
nand U19576 (N_19576,N_19355,N_19317);
or U19577 (N_19577,N_19381,N_19315);
xnor U19578 (N_19578,N_19498,N_19418);
and U19579 (N_19579,N_19356,N_19326);
or U19580 (N_19580,N_19244,N_19469);
xor U19581 (N_19581,N_19361,N_19374);
xor U19582 (N_19582,N_19414,N_19403);
nand U19583 (N_19583,N_19365,N_19440);
and U19584 (N_19584,N_19487,N_19434);
xnor U19585 (N_19585,N_19379,N_19453);
nor U19586 (N_19586,N_19296,N_19420);
and U19587 (N_19587,N_19327,N_19335);
and U19588 (N_19588,N_19408,N_19214);
xor U19589 (N_19589,N_19430,N_19254);
or U19590 (N_19590,N_19235,N_19412);
and U19591 (N_19591,N_19427,N_19219);
or U19592 (N_19592,N_19438,N_19260);
nor U19593 (N_19593,N_19209,N_19392);
nor U19594 (N_19594,N_19491,N_19490);
and U19595 (N_19595,N_19265,N_19312);
and U19596 (N_19596,N_19301,N_19372);
xnor U19597 (N_19597,N_19221,N_19268);
and U19598 (N_19598,N_19232,N_19203);
or U19599 (N_19599,N_19405,N_19489);
nor U19600 (N_19600,N_19480,N_19447);
nor U19601 (N_19601,N_19449,N_19252);
nor U19602 (N_19602,N_19277,N_19460);
or U19603 (N_19603,N_19484,N_19321);
nand U19604 (N_19604,N_19246,N_19343);
or U19605 (N_19605,N_19240,N_19353);
nand U19606 (N_19606,N_19202,N_19222);
nor U19607 (N_19607,N_19243,N_19212);
or U19608 (N_19608,N_19334,N_19471);
nand U19609 (N_19609,N_19479,N_19229);
nor U19610 (N_19610,N_19495,N_19378);
nand U19611 (N_19611,N_19406,N_19323);
or U19612 (N_19612,N_19423,N_19247);
and U19613 (N_19613,N_19370,N_19454);
nand U19614 (N_19614,N_19424,N_19275);
xnor U19615 (N_19615,N_19393,N_19236);
xor U19616 (N_19616,N_19242,N_19461);
nor U19617 (N_19617,N_19442,N_19483);
or U19618 (N_19618,N_19320,N_19426);
nor U19619 (N_19619,N_19223,N_19280);
nor U19620 (N_19620,N_19253,N_19330);
xor U19621 (N_19621,N_19373,N_19354);
nor U19622 (N_19622,N_19284,N_19308);
nor U19623 (N_19623,N_19306,N_19258);
xor U19624 (N_19624,N_19264,N_19360);
nor U19625 (N_19625,N_19389,N_19256);
xor U19626 (N_19626,N_19307,N_19333);
nand U19627 (N_19627,N_19304,N_19398);
nand U19628 (N_19628,N_19482,N_19319);
and U19629 (N_19629,N_19391,N_19394);
nand U19630 (N_19630,N_19444,N_19257);
and U19631 (N_19631,N_19428,N_19346);
or U19632 (N_19632,N_19272,N_19456);
nand U19633 (N_19633,N_19273,N_19397);
and U19634 (N_19634,N_19282,N_19251);
xnor U19635 (N_19635,N_19314,N_19459);
and U19636 (N_19636,N_19201,N_19261);
and U19637 (N_19637,N_19271,N_19369);
nor U19638 (N_19638,N_19225,N_19220);
nor U19639 (N_19639,N_19344,N_19318);
xnor U19640 (N_19640,N_19380,N_19300);
or U19641 (N_19641,N_19416,N_19486);
nand U19642 (N_19642,N_19468,N_19367);
and U19643 (N_19643,N_19473,N_19351);
nand U19644 (N_19644,N_19208,N_19446);
or U19645 (N_19645,N_19465,N_19295);
xnor U19646 (N_19646,N_19216,N_19332);
nor U19647 (N_19647,N_19340,N_19283);
or U19648 (N_19648,N_19492,N_19385);
nand U19649 (N_19649,N_19234,N_19432);
nor U19650 (N_19650,N_19428,N_19469);
nand U19651 (N_19651,N_19211,N_19413);
or U19652 (N_19652,N_19323,N_19359);
and U19653 (N_19653,N_19416,N_19433);
xor U19654 (N_19654,N_19203,N_19476);
xor U19655 (N_19655,N_19409,N_19231);
nor U19656 (N_19656,N_19224,N_19306);
xor U19657 (N_19657,N_19368,N_19420);
and U19658 (N_19658,N_19215,N_19212);
nor U19659 (N_19659,N_19363,N_19227);
xor U19660 (N_19660,N_19397,N_19337);
xor U19661 (N_19661,N_19253,N_19213);
nand U19662 (N_19662,N_19235,N_19465);
nand U19663 (N_19663,N_19240,N_19338);
nand U19664 (N_19664,N_19436,N_19260);
or U19665 (N_19665,N_19374,N_19286);
and U19666 (N_19666,N_19263,N_19221);
nand U19667 (N_19667,N_19219,N_19443);
nor U19668 (N_19668,N_19420,N_19253);
and U19669 (N_19669,N_19299,N_19289);
nand U19670 (N_19670,N_19284,N_19261);
nor U19671 (N_19671,N_19202,N_19352);
or U19672 (N_19672,N_19242,N_19494);
or U19673 (N_19673,N_19410,N_19298);
and U19674 (N_19674,N_19422,N_19348);
nor U19675 (N_19675,N_19419,N_19498);
xor U19676 (N_19676,N_19401,N_19222);
and U19677 (N_19677,N_19278,N_19319);
or U19678 (N_19678,N_19390,N_19346);
and U19679 (N_19679,N_19225,N_19389);
or U19680 (N_19680,N_19474,N_19231);
or U19681 (N_19681,N_19426,N_19356);
and U19682 (N_19682,N_19355,N_19486);
and U19683 (N_19683,N_19326,N_19477);
nor U19684 (N_19684,N_19338,N_19361);
or U19685 (N_19685,N_19245,N_19492);
nor U19686 (N_19686,N_19265,N_19477);
xor U19687 (N_19687,N_19316,N_19419);
xnor U19688 (N_19688,N_19496,N_19252);
xor U19689 (N_19689,N_19216,N_19234);
nand U19690 (N_19690,N_19223,N_19264);
nand U19691 (N_19691,N_19482,N_19371);
nor U19692 (N_19692,N_19348,N_19458);
or U19693 (N_19693,N_19495,N_19404);
xnor U19694 (N_19694,N_19231,N_19422);
nand U19695 (N_19695,N_19206,N_19462);
and U19696 (N_19696,N_19264,N_19464);
nor U19697 (N_19697,N_19321,N_19366);
nand U19698 (N_19698,N_19231,N_19254);
or U19699 (N_19699,N_19237,N_19252);
nor U19700 (N_19700,N_19333,N_19382);
nand U19701 (N_19701,N_19307,N_19270);
or U19702 (N_19702,N_19269,N_19341);
and U19703 (N_19703,N_19249,N_19476);
nor U19704 (N_19704,N_19230,N_19287);
nor U19705 (N_19705,N_19436,N_19344);
nand U19706 (N_19706,N_19363,N_19249);
nand U19707 (N_19707,N_19202,N_19309);
nand U19708 (N_19708,N_19294,N_19264);
or U19709 (N_19709,N_19389,N_19402);
or U19710 (N_19710,N_19391,N_19246);
or U19711 (N_19711,N_19271,N_19375);
xor U19712 (N_19712,N_19253,N_19244);
nand U19713 (N_19713,N_19330,N_19260);
nor U19714 (N_19714,N_19324,N_19425);
nor U19715 (N_19715,N_19393,N_19201);
nand U19716 (N_19716,N_19497,N_19445);
or U19717 (N_19717,N_19355,N_19322);
nand U19718 (N_19718,N_19473,N_19201);
and U19719 (N_19719,N_19372,N_19298);
xor U19720 (N_19720,N_19433,N_19217);
or U19721 (N_19721,N_19258,N_19288);
nand U19722 (N_19722,N_19260,N_19468);
xnor U19723 (N_19723,N_19205,N_19261);
and U19724 (N_19724,N_19408,N_19432);
nor U19725 (N_19725,N_19303,N_19483);
nor U19726 (N_19726,N_19285,N_19497);
or U19727 (N_19727,N_19297,N_19405);
nor U19728 (N_19728,N_19415,N_19383);
nand U19729 (N_19729,N_19393,N_19360);
or U19730 (N_19730,N_19284,N_19459);
and U19731 (N_19731,N_19304,N_19341);
xnor U19732 (N_19732,N_19255,N_19316);
xor U19733 (N_19733,N_19391,N_19363);
nand U19734 (N_19734,N_19252,N_19466);
xor U19735 (N_19735,N_19465,N_19281);
nor U19736 (N_19736,N_19485,N_19397);
and U19737 (N_19737,N_19220,N_19463);
or U19738 (N_19738,N_19289,N_19484);
or U19739 (N_19739,N_19427,N_19346);
nand U19740 (N_19740,N_19412,N_19278);
nor U19741 (N_19741,N_19373,N_19318);
nor U19742 (N_19742,N_19438,N_19467);
and U19743 (N_19743,N_19259,N_19311);
and U19744 (N_19744,N_19302,N_19205);
and U19745 (N_19745,N_19430,N_19308);
and U19746 (N_19746,N_19382,N_19205);
nand U19747 (N_19747,N_19406,N_19332);
nor U19748 (N_19748,N_19338,N_19386);
or U19749 (N_19749,N_19296,N_19417);
or U19750 (N_19750,N_19297,N_19266);
or U19751 (N_19751,N_19472,N_19290);
and U19752 (N_19752,N_19430,N_19460);
nand U19753 (N_19753,N_19425,N_19240);
and U19754 (N_19754,N_19346,N_19373);
nand U19755 (N_19755,N_19294,N_19246);
nor U19756 (N_19756,N_19417,N_19360);
xor U19757 (N_19757,N_19472,N_19211);
or U19758 (N_19758,N_19403,N_19418);
and U19759 (N_19759,N_19223,N_19438);
or U19760 (N_19760,N_19276,N_19361);
xnor U19761 (N_19761,N_19324,N_19222);
or U19762 (N_19762,N_19279,N_19262);
and U19763 (N_19763,N_19366,N_19334);
nor U19764 (N_19764,N_19412,N_19228);
or U19765 (N_19765,N_19363,N_19487);
nor U19766 (N_19766,N_19271,N_19432);
nand U19767 (N_19767,N_19450,N_19314);
nand U19768 (N_19768,N_19417,N_19427);
nand U19769 (N_19769,N_19234,N_19427);
nor U19770 (N_19770,N_19318,N_19269);
xor U19771 (N_19771,N_19498,N_19294);
or U19772 (N_19772,N_19364,N_19362);
xnor U19773 (N_19773,N_19323,N_19258);
and U19774 (N_19774,N_19200,N_19256);
and U19775 (N_19775,N_19400,N_19379);
nor U19776 (N_19776,N_19447,N_19345);
nand U19777 (N_19777,N_19477,N_19372);
xor U19778 (N_19778,N_19356,N_19408);
nor U19779 (N_19779,N_19381,N_19482);
or U19780 (N_19780,N_19219,N_19288);
nor U19781 (N_19781,N_19465,N_19455);
nand U19782 (N_19782,N_19297,N_19212);
nand U19783 (N_19783,N_19242,N_19301);
nor U19784 (N_19784,N_19499,N_19309);
nor U19785 (N_19785,N_19496,N_19243);
and U19786 (N_19786,N_19301,N_19244);
nand U19787 (N_19787,N_19208,N_19336);
xor U19788 (N_19788,N_19329,N_19291);
xor U19789 (N_19789,N_19371,N_19413);
and U19790 (N_19790,N_19378,N_19346);
or U19791 (N_19791,N_19343,N_19353);
nor U19792 (N_19792,N_19385,N_19334);
and U19793 (N_19793,N_19472,N_19220);
nor U19794 (N_19794,N_19227,N_19257);
nor U19795 (N_19795,N_19235,N_19322);
and U19796 (N_19796,N_19313,N_19335);
nand U19797 (N_19797,N_19306,N_19215);
nand U19798 (N_19798,N_19343,N_19383);
or U19799 (N_19799,N_19263,N_19355);
xnor U19800 (N_19800,N_19760,N_19537);
xor U19801 (N_19801,N_19622,N_19595);
or U19802 (N_19802,N_19665,N_19511);
or U19803 (N_19803,N_19777,N_19520);
or U19804 (N_19804,N_19653,N_19671);
xor U19805 (N_19805,N_19798,N_19580);
and U19806 (N_19806,N_19536,N_19692);
and U19807 (N_19807,N_19594,N_19654);
xnor U19808 (N_19808,N_19574,N_19538);
nand U19809 (N_19809,N_19601,N_19613);
nor U19810 (N_19810,N_19540,N_19640);
nand U19811 (N_19811,N_19651,N_19605);
and U19812 (N_19812,N_19576,N_19614);
xnor U19813 (N_19813,N_19592,N_19701);
nor U19814 (N_19814,N_19512,N_19784);
xnor U19815 (N_19815,N_19697,N_19603);
or U19816 (N_19816,N_19578,N_19523);
and U19817 (N_19817,N_19567,N_19694);
xnor U19818 (N_19818,N_19772,N_19588);
xnor U19819 (N_19819,N_19747,N_19794);
and U19820 (N_19820,N_19677,N_19650);
and U19821 (N_19821,N_19531,N_19624);
and U19822 (N_19822,N_19673,N_19717);
nor U19823 (N_19823,N_19733,N_19725);
or U19824 (N_19824,N_19556,N_19795);
and U19825 (N_19825,N_19663,N_19690);
nor U19826 (N_19826,N_19749,N_19658);
xor U19827 (N_19827,N_19593,N_19771);
xnor U19828 (N_19828,N_19645,N_19604);
xor U19829 (N_19829,N_19708,N_19790);
or U19830 (N_19830,N_19590,N_19646);
and U19831 (N_19831,N_19517,N_19786);
nor U19832 (N_19832,N_19639,N_19530);
nand U19833 (N_19833,N_19674,N_19695);
and U19834 (N_19834,N_19579,N_19791);
nor U19835 (N_19835,N_19630,N_19670);
and U19836 (N_19836,N_19687,N_19766);
nand U19837 (N_19837,N_19596,N_19737);
and U19838 (N_19838,N_19734,N_19738);
xor U19839 (N_19839,N_19775,N_19634);
xor U19840 (N_19840,N_19551,N_19713);
or U19841 (N_19841,N_19657,N_19757);
nor U19842 (N_19842,N_19507,N_19621);
nor U19843 (N_19843,N_19788,N_19689);
xor U19844 (N_19844,N_19608,N_19669);
nor U19845 (N_19845,N_19611,N_19545);
nand U19846 (N_19846,N_19575,N_19732);
xnor U19847 (N_19847,N_19615,N_19504);
and U19848 (N_19848,N_19526,N_19680);
nor U19849 (N_19849,N_19529,N_19704);
xor U19850 (N_19850,N_19516,N_19660);
nand U19851 (N_19851,N_19702,N_19513);
and U19852 (N_19852,N_19623,N_19503);
nor U19853 (N_19853,N_19719,N_19607);
nand U19854 (N_19854,N_19612,N_19550);
and U19855 (N_19855,N_19779,N_19635);
or U19856 (N_19856,N_19632,N_19548);
and U19857 (N_19857,N_19647,N_19561);
xor U19858 (N_19858,N_19500,N_19618);
and U19859 (N_19859,N_19714,N_19649);
and U19860 (N_19860,N_19533,N_19711);
or U19861 (N_19861,N_19644,N_19678);
xnor U19862 (N_19862,N_19557,N_19724);
and U19863 (N_19863,N_19797,N_19706);
nand U19864 (N_19864,N_19570,N_19569);
and U19865 (N_19865,N_19782,N_19528);
xor U19866 (N_19866,N_19721,N_19666);
or U19867 (N_19867,N_19787,N_19633);
nand U19868 (N_19868,N_19769,N_19506);
nand U19869 (N_19869,N_19655,N_19744);
and U19870 (N_19870,N_19763,N_19643);
nor U19871 (N_19871,N_19573,N_19552);
nand U19872 (N_19872,N_19761,N_19686);
nand U19873 (N_19873,N_19542,N_19586);
xor U19874 (N_19874,N_19572,N_19683);
nand U19875 (N_19875,N_19781,N_19659);
and U19876 (N_19876,N_19793,N_19652);
nor U19877 (N_19877,N_19774,N_19524);
or U19878 (N_19878,N_19532,N_19637);
nor U19879 (N_19879,N_19543,N_19606);
nand U19880 (N_19880,N_19541,N_19510);
or U19881 (N_19881,N_19589,N_19508);
and U19882 (N_19882,N_19765,N_19558);
nand U19883 (N_19883,N_19672,N_19745);
nor U19884 (N_19884,N_19581,N_19656);
nand U19885 (N_19885,N_19722,N_19696);
or U19886 (N_19886,N_19554,N_19707);
xnor U19887 (N_19887,N_19591,N_19549);
nor U19888 (N_19888,N_19667,N_19699);
nor U19889 (N_19889,N_19705,N_19560);
and U19890 (N_19890,N_19514,N_19584);
xnor U19891 (N_19891,N_19662,N_19741);
and U19892 (N_19892,N_19585,N_19746);
and U19893 (N_19893,N_19735,N_19522);
xor U19894 (N_19894,N_19712,N_19750);
and U19895 (N_19895,N_19789,N_19703);
nor U19896 (N_19896,N_19502,N_19521);
nor U19897 (N_19897,N_19571,N_19748);
or U19898 (N_19898,N_19559,N_19739);
xor U19899 (N_19899,N_19783,N_19676);
nor U19900 (N_19900,N_19636,N_19715);
or U19901 (N_19901,N_19627,N_19718);
and U19902 (N_19902,N_19698,N_19756);
and U19903 (N_19903,N_19726,N_19778);
or U19904 (N_19904,N_19641,N_19742);
and U19905 (N_19905,N_19723,N_19727);
nand U19906 (N_19906,N_19664,N_19693);
nor U19907 (N_19907,N_19768,N_19610);
xor U19908 (N_19908,N_19598,N_19505);
xor U19909 (N_19909,N_19720,N_19616);
or U19910 (N_19910,N_19562,N_19602);
and U19911 (N_19911,N_19518,N_19759);
nand U19912 (N_19912,N_19752,N_19762);
and U19913 (N_19913,N_19758,N_19780);
and U19914 (N_19914,N_19675,N_19688);
xor U19915 (N_19915,N_19620,N_19736);
or U19916 (N_19916,N_19565,N_19619);
xnor U19917 (N_19917,N_19740,N_19583);
xnor U19918 (N_19918,N_19582,N_19638);
or U19919 (N_19919,N_19519,N_19764);
xor U19920 (N_19920,N_19773,N_19642);
xor U19921 (N_19921,N_19710,N_19568);
or U19922 (N_19922,N_19700,N_19527);
nand U19923 (N_19923,N_19755,N_19709);
nor U19924 (N_19924,N_19515,N_19626);
nor U19925 (N_19925,N_19587,N_19679);
and U19926 (N_19926,N_19563,N_19600);
xor U19927 (N_19927,N_19730,N_19754);
and U19928 (N_19928,N_19685,N_19785);
xor U19929 (N_19929,N_19544,N_19731);
xnor U19930 (N_19930,N_19597,N_19564);
and U19931 (N_19931,N_19792,N_19770);
or U19932 (N_19932,N_19566,N_19525);
nand U19933 (N_19933,N_19625,N_19553);
or U19934 (N_19934,N_19796,N_19729);
nand U19935 (N_19935,N_19599,N_19535);
and U19936 (N_19936,N_19629,N_19539);
xor U19937 (N_19937,N_19753,N_19509);
nand U19938 (N_19938,N_19728,N_19577);
or U19939 (N_19939,N_19609,N_19716);
nor U19940 (N_19940,N_19547,N_19617);
nor U19941 (N_19941,N_19546,N_19767);
nand U19942 (N_19942,N_19684,N_19534);
nor U19943 (N_19943,N_19751,N_19628);
nand U19944 (N_19944,N_19799,N_19661);
xnor U19945 (N_19945,N_19776,N_19648);
or U19946 (N_19946,N_19682,N_19681);
xnor U19947 (N_19947,N_19555,N_19501);
nor U19948 (N_19948,N_19631,N_19668);
nand U19949 (N_19949,N_19691,N_19743);
nand U19950 (N_19950,N_19679,N_19616);
and U19951 (N_19951,N_19552,N_19641);
nand U19952 (N_19952,N_19601,N_19747);
xor U19953 (N_19953,N_19741,N_19760);
and U19954 (N_19954,N_19638,N_19775);
or U19955 (N_19955,N_19746,N_19783);
or U19956 (N_19956,N_19711,N_19529);
or U19957 (N_19957,N_19535,N_19506);
xnor U19958 (N_19958,N_19601,N_19528);
nand U19959 (N_19959,N_19711,N_19634);
nor U19960 (N_19960,N_19791,N_19664);
or U19961 (N_19961,N_19782,N_19739);
or U19962 (N_19962,N_19652,N_19795);
or U19963 (N_19963,N_19710,N_19671);
and U19964 (N_19964,N_19517,N_19688);
xor U19965 (N_19965,N_19506,N_19601);
xnor U19966 (N_19966,N_19728,N_19663);
and U19967 (N_19967,N_19597,N_19614);
nand U19968 (N_19968,N_19716,N_19677);
or U19969 (N_19969,N_19526,N_19734);
nor U19970 (N_19970,N_19590,N_19602);
xnor U19971 (N_19971,N_19513,N_19714);
nor U19972 (N_19972,N_19596,N_19767);
nor U19973 (N_19973,N_19770,N_19618);
and U19974 (N_19974,N_19793,N_19692);
nand U19975 (N_19975,N_19518,N_19520);
nor U19976 (N_19976,N_19556,N_19791);
or U19977 (N_19977,N_19669,N_19651);
nand U19978 (N_19978,N_19550,N_19788);
or U19979 (N_19979,N_19744,N_19746);
and U19980 (N_19980,N_19686,N_19792);
nor U19981 (N_19981,N_19607,N_19750);
nand U19982 (N_19982,N_19504,N_19777);
xnor U19983 (N_19983,N_19512,N_19578);
nor U19984 (N_19984,N_19606,N_19623);
or U19985 (N_19985,N_19592,N_19507);
nor U19986 (N_19986,N_19618,N_19672);
or U19987 (N_19987,N_19682,N_19716);
xor U19988 (N_19988,N_19780,N_19744);
xor U19989 (N_19989,N_19681,N_19524);
nor U19990 (N_19990,N_19585,N_19622);
or U19991 (N_19991,N_19757,N_19670);
and U19992 (N_19992,N_19783,N_19736);
xor U19993 (N_19993,N_19683,N_19705);
and U19994 (N_19994,N_19557,N_19746);
or U19995 (N_19995,N_19568,N_19758);
or U19996 (N_19996,N_19600,N_19755);
or U19997 (N_19997,N_19547,N_19756);
and U19998 (N_19998,N_19615,N_19666);
nand U19999 (N_19999,N_19569,N_19708);
nor U20000 (N_20000,N_19767,N_19725);
or U20001 (N_20001,N_19526,N_19631);
xnor U20002 (N_20002,N_19558,N_19734);
or U20003 (N_20003,N_19775,N_19628);
nor U20004 (N_20004,N_19637,N_19615);
xnor U20005 (N_20005,N_19520,N_19661);
nand U20006 (N_20006,N_19638,N_19640);
and U20007 (N_20007,N_19545,N_19796);
and U20008 (N_20008,N_19580,N_19533);
and U20009 (N_20009,N_19759,N_19723);
nor U20010 (N_20010,N_19542,N_19784);
or U20011 (N_20011,N_19781,N_19793);
and U20012 (N_20012,N_19574,N_19549);
nor U20013 (N_20013,N_19605,N_19671);
or U20014 (N_20014,N_19705,N_19503);
and U20015 (N_20015,N_19548,N_19710);
and U20016 (N_20016,N_19652,N_19783);
and U20017 (N_20017,N_19700,N_19684);
or U20018 (N_20018,N_19564,N_19568);
or U20019 (N_20019,N_19510,N_19687);
xor U20020 (N_20020,N_19640,N_19669);
or U20021 (N_20021,N_19524,N_19682);
nand U20022 (N_20022,N_19697,N_19713);
nand U20023 (N_20023,N_19601,N_19609);
xnor U20024 (N_20024,N_19548,N_19620);
xnor U20025 (N_20025,N_19519,N_19602);
or U20026 (N_20026,N_19513,N_19532);
nand U20027 (N_20027,N_19559,N_19636);
nor U20028 (N_20028,N_19549,N_19656);
and U20029 (N_20029,N_19545,N_19522);
nor U20030 (N_20030,N_19508,N_19575);
or U20031 (N_20031,N_19700,N_19729);
or U20032 (N_20032,N_19606,N_19685);
nor U20033 (N_20033,N_19664,N_19601);
nor U20034 (N_20034,N_19549,N_19530);
xnor U20035 (N_20035,N_19500,N_19545);
or U20036 (N_20036,N_19621,N_19573);
and U20037 (N_20037,N_19690,N_19572);
xor U20038 (N_20038,N_19777,N_19665);
xnor U20039 (N_20039,N_19538,N_19743);
nand U20040 (N_20040,N_19582,N_19564);
and U20041 (N_20041,N_19703,N_19662);
nand U20042 (N_20042,N_19793,N_19601);
and U20043 (N_20043,N_19539,N_19711);
nor U20044 (N_20044,N_19608,N_19683);
nor U20045 (N_20045,N_19562,N_19516);
or U20046 (N_20046,N_19709,N_19745);
nand U20047 (N_20047,N_19574,N_19592);
or U20048 (N_20048,N_19680,N_19675);
nand U20049 (N_20049,N_19651,N_19773);
or U20050 (N_20050,N_19740,N_19778);
nor U20051 (N_20051,N_19674,N_19523);
or U20052 (N_20052,N_19517,N_19782);
xor U20053 (N_20053,N_19579,N_19641);
nand U20054 (N_20054,N_19642,N_19788);
nor U20055 (N_20055,N_19792,N_19782);
nor U20056 (N_20056,N_19534,N_19696);
nor U20057 (N_20057,N_19516,N_19577);
nand U20058 (N_20058,N_19791,N_19691);
and U20059 (N_20059,N_19668,N_19719);
or U20060 (N_20060,N_19773,N_19541);
nor U20061 (N_20061,N_19508,N_19695);
and U20062 (N_20062,N_19781,N_19586);
nor U20063 (N_20063,N_19654,N_19513);
nand U20064 (N_20064,N_19540,N_19680);
and U20065 (N_20065,N_19631,N_19751);
or U20066 (N_20066,N_19524,N_19749);
or U20067 (N_20067,N_19577,N_19778);
and U20068 (N_20068,N_19772,N_19516);
nor U20069 (N_20069,N_19712,N_19613);
or U20070 (N_20070,N_19533,N_19733);
or U20071 (N_20071,N_19746,N_19533);
or U20072 (N_20072,N_19585,N_19630);
nor U20073 (N_20073,N_19526,N_19607);
nor U20074 (N_20074,N_19696,N_19524);
nand U20075 (N_20075,N_19618,N_19659);
xor U20076 (N_20076,N_19693,N_19697);
xor U20077 (N_20077,N_19661,N_19720);
xnor U20078 (N_20078,N_19659,N_19784);
nand U20079 (N_20079,N_19691,N_19765);
nor U20080 (N_20080,N_19604,N_19771);
and U20081 (N_20081,N_19582,N_19536);
or U20082 (N_20082,N_19738,N_19652);
nand U20083 (N_20083,N_19504,N_19545);
nand U20084 (N_20084,N_19748,N_19682);
xor U20085 (N_20085,N_19635,N_19624);
nand U20086 (N_20086,N_19797,N_19512);
nand U20087 (N_20087,N_19747,N_19511);
xor U20088 (N_20088,N_19584,N_19735);
nand U20089 (N_20089,N_19798,N_19691);
and U20090 (N_20090,N_19503,N_19591);
nor U20091 (N_20091,N_19577,N_19736);
nor U20092 (N_20092,N_19756,N_19624);
or U20093 (N_20093,N_19635,N_19536);
or U20094 (N_20094,N_19582,N_19672);
xnor U20095 (N_20095,N_19581,N_19785);
or U20096 (N_20096,N_19640,N_19520);
and U20097 (N_20097,N_19587,N_19536);
and U20098 (N_20098,N_19622,N_19647);
nand U20099 (N_20099,N_19730,N_19587);
and U20100 (N_20100,N_19808,N_19910);
xnor U20101 (N_20101,N_19852,N_19956);
xor U20102 (N_20102,N_19893,N_19960);
xor U20103 (N_20103,N_19881,N_19961);
nor U20104 (N_20104,N_20052,N_20077);
nor U20105 (N_20105,N_19928,N_20057);
nand U20106 (N_20106,N_19877,N_19965);
nand U20107 (N_20107,N_19952,N_19879);
or U20108 (N_20108,N_20092,N_20041);
xor U20109 (N_20109,N_20055,N_19812);
and U20110 (N_20110,N_19837,N_19942);
and U20111 (N_20111,N_20087,N_20083);
xor U20112 (N_20112,N_19828,N_20014);
xor U20113 (N_20113,N_20051,N_19823);
nand U20114 (N_20114,N_19935,N_19996);
xnor U20115 (N_20115,N_19885,N_19816);
xor U20116 (N_20116,N_19941,N_19826);
nor U20117 (N_20117,N_19882,N_19806);
nand U20118 (N_20118,N_19983,N_20089);
or U20119 (N_20119,N_20029,N_19886);
or U20120 (N_20120,N_19814,N_19957);
or U20121 (N_20121,N_19921,N_19979);
nor U20122 (N_20122,N_20062,N_20048);
and U20123 (N_20123,N_19973,N_19829);
nor U20124 (N_20124,N_20037,N_19844);
and U20125 (N_20125,N_19800,N_19834);
xnor U20126 (N_20126,N_20069,N_20064);
and U20127 (N_20127,N_20043,N_20028);
nor U20128 (N_20128,N_20073,N_19891);
nor U20129 (N_20129,N_20007,N_19999);
xor U20130 (N_20130,N_20090,N_19909);
nand U20131 (N_20131,N_19905,N_19997);
nand U20132 (N_20132,N_19987,N_19975);
xor U20133 (N_20133,N_19914,N_20006);
nand U20134 (N_20134,N_19873,N_19818);
nor U20135 (N_20135,N_19995,N_19802);
or U20136 (N_20136,N_20097,N_19892);
nor U20137 (N_20137,N_20024,N_19867);
nand U20138 (N_20138,N_20049,N_19878);
or U20139 (N_20139,N_20032,N_19856);
nand U20140 (N_20140,N_19863,N_19858);
and U20141 (N_20141,N_19930,N_20063);
xnor U20142 (N_20142,N_19972,N_19809);
and U20143 (N_20143,N_20082,N_20017);
xnor U20144 (N_20144,N_20046,N_19984);
xor U20145 (N_20145,N_20076,N_19865);
nor U20146 (N_20146,N_19980,N_20096);
nor U20147 (N_20147,N_19929,N_20036);
or U20148 (N_20148,N_19846,N_19845);
nor U20149 (N_20149,N_19925,N_19832);
nand U20150 (N_20150,N_20065,N_20093);
nand U20151 (N_20151,N_20027,N_20053);
xnor U20152 (N_20152,N_20058,N_19861);
nor U20153 (N_20153,N_20059,N_19815);
xor U20154 (N_20154,N_20066,N_19974);
xnor U20155 (N_20155,N_19945,N_19920);
xnor U20156 (N_20156,N_19934,N_20005);
or U20157 (N_20157,N_20009,N_20068);
and U20158 (N_20158,N_20050,N_19847);
and U20159 (N_20159,N_19841,N_19944);
nor U20160 (N_20160,N_20084,N_19962);
and U20161 (N_20161,N_19913,N_19978);
nor U20162 (N_20162,N_20056,N_19854);
nand U20163 (N_20163,N_19989,N_19949);
nor U20164 (N_20164,N_19831,N_19968);
or U20165 (N_20165,N_20020,N_19880);
and U20166 (N_20166,N_20086,N_19947);
or U20167 (N_20167,N_19993,N_19966);
nand U20168 (N_20168,N_19981,N_19932);
nand U20169 (N_20169,N_19872,N_20095);
nor U20170 (N_20170,N_19883,N_19839);
and U20171 (N_20171,N_20085,N_19931);
or U20172 (N_20172,N_19906,N_19959);
nor U20173 (N_20173,N_19933,N_20088);
nand U20174 (N_20174,N_19948,N_20026);
and U20175 (N_20175,N_20039,N_19970);
or U20176 (N_20176,N_20022,N_19884);
xnor U20177 (N_20177,N_19803,N_20003);
nand U20178 (N_20178,N_19898,N_19915);
nand U20179 (N_20179,N_19991,N_19821);
nand U20180 (N_20180,N_19801,N_19848);
nor U20181 (N_20181,N_19866,N_19967);
and U20182 (N_20182,N_19922,N_19977);
and U20183 (N_20183,N_19890,N_19969);
and U20184 (N_20184,N_19864,N_20025);
and U20185 (N_20185,N_19860,N_19888);
xnor U20186 (N_20186,N_19874,N_19849);
nand U20187 (N_20187,N_19958,N_19908);
or U20188 (N_20188,N_19838,N_19868);
nand U20189 (N_20189,N_19807,N_20030);
nor U20190 (N_20190,N_19889,N_19937);
nand U20191 (N_20191,N_19982,N_20015);
or U20192 (N_20192,N_19902,N_19918);
or U20193 (N_20193,N_19871,N_20094);
xnor U20194 (N_20194,N_19911,N_19859);
or U20195 (N_20195,N_19819,N_19899);
nor U20196 (N_20196,N_20047,N_20067);
nand U20197 (N_20197,N_20012,N_19901);
nand U20198 (N_20198,N_20099,N_20045);
xnor U20199 (N_20199,N_19938,N_19950);
nor U20200 (N_20200,N_19875,N_19805);
nand U20201 (N_20201,N_20072,N_19855);
nor U20202 (N_20202,N_20018,N_20091);
xor U20203 (N_20203,N_19923,N_19912);
and U20204 (N_20204,N_19924,N_20004);
and U20205 (N_20205,N_20021,N_20019);
xor U20206 (N_20206,N_19927,N_19940);
nand U20207 (N_20207,N_19954,N_19951);
xor U20208 (N_20208,N_19810,N_19862);
nand U20209 (N_20209,N_20035,N_19843);
nor U20210 (N_20210,N_19853,N_20042);
and U20211 (N_20211,N_19963,N_20001);
and U20212 (N_20212,N_19904,N_19971);
nor U20213 (N_20213,N_19851,N_20075);
xor U20214 (N_20214,N_19990,N_19964);
nor U20215 (N_20215,N_19985,N_19998);
nor U20216 (N_20216,N_20010,N_19896);
and U20217 (N_20217,N_19804,N_19988);
or U20218 (N_20218,N_19835,N_19926);
nor U20219 (N_20219,N_20002,N_20074);
nor U20220 (N_20220,N_20079,N_19817);
or U20221 (N_20221,N_19903,N_19994);
nand U20222 (N_20222,N_20008,N_19992);
nand U20223 (N_20223,N_19917,N_20070);
xnor U20224 (N_20224,N_19876,N_20054);
xnor U20225 (N_20225,N_19953,N_19986);
or U20226 (N_20226,N_19887,N_19813);
or U20227 (N_20227,N_20078,N_19936);
nand U20228 (N_20228,N_20016,N_19919);
nor U20229 (N_20229,N_19894,N_20031);
or U20230 (N_20230,N_19830,N_19939);
nand U20231 (N_20231,N_19822,N_20098);
or U20232 (N_20232,N_19857,N_20011);
and U20233 (N_20233,N_20071,N_20061);
and U20234 (N_20234,N_20034,N_19869);
and U20235 (N_20235,N_20033,N_19820);
and U20236 (N_20236,N_19811,N_19946);
nand U20237 (N_20237,N_20044,N_19842);
or U20238 (N_20238,N_20000,N_20080);
nor U20239 (N_20239,N_19870,N_19900);
and U20240 (N_20240,N_19833,N_20060);
nand U20241 (N_20241,N_19850,N_19836);
nor U20242 (N_20242,N_19943,N_20013);
nor U20243 (N_20243,N_19955,N_20038);
or U20244 (N_20244,N_20040,N_20081);
and U20245 (N_20245,N_19895,N_19827);
or U20246 (N_20246,N_20023,N_19916);
nor U20247 (N_20247,N_19824,N_19907);
and U20248 (N_20248,N_19840,N_19976);
xor U20249 (N_20249,N_19825,N_19897);
nor U20250 (N_20250,N_19822,N_20032);
nor U20251 (N_20251,N_19836,N_19985);
nor U20252 (N_20252,N_20078,N_19946);
or U20253 (N_20253,N_19818,N_19896);
nor U20254 (N_20254,N_20079,N_19897);
xnor U20255 (N_20255,N_19869,N_19908);
nor U20256 (N_20256,N_19867,N_20085);
nor U20257 (N_20257,N_19856,N_20058);
nand U20258 (N_20258,N_19966,N_20044);
nor U20259 (N_20259,N_20083,N_19985);
and U20260 (N_20260,N_20023,N_19947);
xnor U20261 (N_20261,N_20029,N_19968);
nor U20262 (N_20262,N_19834,N_20034);
or U20263 (N_20263,N_20027,N_20084);
nor U20264 (N_20264,N_19894,N_20036);
and U20265 (N_20265,N_19802,N_20039);
and U20266 (N_20266,N_20052,N_19857);
and U20267 (N_20267,N_19908,N_20014);
nor U20268 (N_20268,N_19953,N_20020);
nor U20269 (N_20269,N_19942,N_20023);
nand U20270 (N_20270,N_20091,N_19864);
or U20271 (N_20271,N_20017,N_19958);
nand U20272 (N_20272,N_20086,N_20002);
nand U20273 (N_20273,N_20035,N_19897);
nand U20274 (N_20274,N_19891,N_19947);
xnor U20275 (N_20275,N_19839,N_19886);
xor U20276 (N_20276,N_19907,N_19885);
or U20277 (N_20277,N_19997,N_19915);
or U20278 (N_20278,N_19931,N_20055);
nor U20279 (N_20279,N_20022,N_20039);
and U20280 (N_20280,N_19940,N_19807);
or U20281 (N_20281,N_20018,N_20046);
nor U20282 (N_20282,N_20081,N_19848);
or U20283 (N_20283,N_19995,N_19834);
nand U20284 (N_20284,N_20097,N_19911);
xnor U20285 (N_20285,N_20019,N_19806);
nor U20286 (N_20286,N_19897,N_20049);
xnor U20287 (N_20287,N_19990,N_19865);
and U20288 (N_20288,N_19972,N_19842);
xnor U20289 (N_20289,N_19961,N_20073);
or U20290 (N_20290,N_19853,N_19810);
nor U20291 (N_20291,N_19980,N_19932);
xor U20292 (N_20292,N_19993,N_19905);
nand U20293 (N_20293,N_19903,N_19877);
nor U20294 (N_20294,N_19961,N_19995);
or U20295 (N_20295,N_19859,N_19838);
xnor U20296 (N_20296,N_19921,N_20071);
and U20297 (N_20297,N_19805,N_20047);
nand U20298 (N_20298,N_19903,N_20017);
and U20299 (N_20299,N_19832,N_19814);
xnor U20300 (N_20300,N_20088,N_20024);
or U20301 (N_20301,N_19882,N_20084);
xnor U20302 (N_20302,N_20015,N_19931);
nand U20303 (N_20303,N_19874,N_20030);
nor U20304 (N_20304,N_19913,N_20073);
nand U20305 (N_20305,N_19872,N_20046);
nor U20306 (N_20306,N_19804,N_19961);
or U20307 (N_20307,N_19998,N_20089);
and U20308 (N_20308,N_19934,N_19977);
or U20309 (N_20309,N_20094,N_20019);
nor U20310 (N_20310,N_19950,N_19819);
and U20311 (N_20311,N_19901,N_19885);
nor U20312 (N_20312,N_19978,N_19801);
and U20313 (N_20313,N_19827,N_19965);
and U20314 (N_20314,N_19814,N_20030);
and U20315 (N_20315,N_19836,N_19956);
nor U20316 (N_20316,N_20040,N_19966);
nor U20317 (N_20317,N_19912,N_19802);
xnor U20318 (N_20318,N_20028,N_19947);
or U20319 (N_20319,N_19904,N_19888);
or U20320 (N_20320,N_20059,N_19888);
or U20321 (N_20321,N_20051,N_20068);
xor U20322 (N_20322,N_19911,N_20085);
nor U20323 (N_20323,N_19891,N_20037);
xnor U20324 (N_20324,N_19984,N_19912);
nor U20325 (N_20325,N_19881,N_19988);
and U20326 (N_20326,N_19930,N_19814);
and U20327 (N_20327,N_19861,N_19983);
or U20328 (N_20328,N_20087,N_19998);
and U20329 (N_20329,N_20012,N_19879);
nand U20330 (N_20330,N_19846,N_19830);
nor U20331 (N_20331,N_20006,N_19934);
and U20332 (N_20332,N_20087,N_19831);
nand U20333 (N_20333,N_19996,N_19879);
xor U20334 (N_20334,N_19828,N_19877);
and U20335 (N_20335,N_20079,N_19996);
nor U20336 (N_20336,N_19889,N_19936);
or U20337 (N_20337,N_20045,N_19895);
nor U20338 (N_20338,N_19892,N_19877);
xnor U20339 (N_20339,N_19956,N_19962);
nor U20340 (N_20340,N_19907,N_20075);
nand U20341 (N_20341,N_20081,N_20068);
nand U20342 (N_20342,N_19810,N_20059);
nor U20343 (N_20343,N_19806,N_20074);
xnor U20344 (N_20344,N_19829,N_20084);
nor U20345 (N_20345,N_19994,N_19975);
or U20346 (N_20346,N_20099,N_19832);
and U20347 (N_20347,N_19872,N_20072);
and U20348 (N_20348,N_20037,N_19819);
nor U20349 (N_20349,N_19809,N_19862);
xnor U20350 (N_20350,N_20046,N_20016);
nor U20351 (N_20351,N_20011,N_19924);
and U20352 (N_20352,N_19936,N_19949);
and U20353 (N_20353,N_19901,N_20094);
nand U20354 (N_20354,N_19937,N_19968);
and U20355 (N_20355,N_20057,N_19817);
nor U20356 (N_20356,N_20071,N_19888);
and U20357 (N_20357,N_19917,N_19875);
nor U20358 (N_20358,N_20066,N_19952);
or U20359 (N_20359,N_19915,N_19828);
nor U20360 (N_20360,N_20007,N_20028);
xnor U20361 (N_20361,N_19913,N_19998);
xor U20362 (N_20362,N_19928,N_19843);
nor U20363 (N_20363,N_20022,N_20088);
nor U20364 (N_20364,N_19855,N_20002);
nand U20365 (N_20365,N_20033,N_20092);
or U20366 (N_20366,N_19954,N_19923);
xnor U20367 (N_20367,N_19857,N_19973);
nor U20368 (N_20368,N_19818,N_19996);
nand U20369 (N_20369,N_20050,N_19902);
and U20370 (N_20370,N_19963,N_20016);
or U20371 (N_20371,N_19844,N_20068);
nor U20372 (N_20372,N_19848,N_20026);
or U20373 (N_20373,N_20038,N_20007);
or U20374 (N_20374,N_19935,N_20087);
or U20375 (N_20375,N_20032,N_19998);
nor U20376 (N_20376,N_20093,N_19928);
or U20377 (N_20377,N_19811,N_20021);
or U20378 (N_20378,N_19851,N_20032);
xnor U20379 (N_20379,N_19921,N_19865);
nand U20380 (N_20380,N_19916,N_19877);
or U20381 (N_20381,N_19836,N_20042);
xor U20382 (N_20382,N_19977,N_19870);
xor U20383 (N_20383,N_20088,N_19820);
nor U20384 (N_20384,N_19883,N_19948);
xor U20385 (N_20385,N_20062,N_19890);
xor U20386 (N_20386,N_19896,N_20036);
nand U20387 (N_20387,N_20075,N_19815);
nand U20388 (N_20388,N_19834,N_20079);
nand U20389 (N_20389,N_19817,N_19948);
nand U20390 (N_20390,N_20054,N_20010);
nand U20391 (N_20391,N_19819,N_19957);
or U20392 (N_20392,N_19970,N_19814);
and U20393 (N_20393,N_19856,N_20040);
nand U20394 (N_20394,N_19835,N_19921);
nor U20395 (N_20395,N_20075,N_19841);
nand U20396 (N_20396,N_19835,N_19837);
and U20397 (N_20397,N_19946,N_20042);
and U20398 (N_20398,N_19813,N_20067);
nand U20399 (N_20399,N_19835,N_19865);
nand U20400 (N_20400,N_20126,N_20144);
nor U20401 (N_20401,N_20357,N_20231);
nor U20402 (N_20402,N_20109,N_20377);
nand U20403 (N_20403,N_20224,N_20110);
or U20404 (N_20404,N_20367,N_20286);
or U20405 (N_20405,N_20235,N_20351);
nor U20406 (N_20406,N_20196,N_20240);
nor U20407 (N_20407,N_20354,N_20300);
xor U20408 (N_20408,N_20362,N_20128);
nand U20409 (N_20409,N_20147,N_20160);
nand U20410 (N_20410,N_20325,N_20385);
xnor U20411 (N_20411,N_20330,N_20179);
and U20412 (N_20412,N_20275,N_20309);
or U20413 (N_20413,N_20138,N_20168);
nand U20414 (N_20414,N_20242,N_20305);
nor U20415 (N_20415,N_20254,N_20181);
or U20416 (N_20416,N_20302,N_20184);
xnor U20417 (N_20417,N_20101,N_20156);
nor U20418 (N_20418,N_20393,N_20399);
nor U20419 (N_20419,N_20256,N_20328);
nand U20420 (N_20420,N_20392,N_20382);
and U20421 (N_20421,N_20165,N_20200);
and U20422 (N_20422,N_20182,N_20365);
nor U20423 (N_20423,N_20271,N_20143);
and U20424 (N_20424,N_20215,N_20263);
or U20425 (N_20425,N_20121,N_20206);
xor U20426 (N_20426,N_20232,N_20250);
nand U20427 (N_20427,N_20313,N_20304);
xnor U20428 (N_20428,N_20148,N_20282);
nor U20429 (N_20429,N_20386,N_20288);
nor U20430 (N_20430,N_20387,N_20380);
and U20431 (N_20431,N_20149,N_20205);
nor U20432 (N_20432,N_20381,N_20376);
and U20433 (N_20433,N_20237,N_20145);
nor U20434 (N_20434,N_20295,N_20344);
nand U20435 (N_20435,N_20312,N_20326);
nand U20436 (N_20436,N_20100,N_20293);
nor U20437 (N_20437,N_20290,N_20236);
nor U20438 (N_20438,N_20324,N_20241);
nor U20439 (N_20439,N_20177,N_20199);
nor U20440 (N_20440,N_20105,N_20135);
and U20441 (N_20441,N_20310,N_20142);
or U20442 (N_20442,N_20358,N_20187);
or U20443 (N_20443,N_20146,N_20227);
and U20444 (N_20444,N_20244,N_20315);
nor U20445 (N_20445,N_20183,N_20391);
and U20446 (N_20446,N_20174,N_20139);
nand U20447 (N_20447,N_20347,N_20269);
or U20448 (N_20448,N_20397,N_20363);
and U20449 (N_20449,N_20189,N_20141);
nand U20450 (N_20450,N_20249,N_20117);
or U20451 (N_20451,N_20172,N_20252);
or U20452 (N_20452,N_20297,N_20259);
or U20453 (N_20453,N_20116,N_20319);
nand U20454 (N_20454,N_20229,N_20216);
or U20455 (N_20455,N_20296,N_20372);
or U20456 (N_20456,N_20337,N_20151);
nand U20457 (N_20457,N_20191,N_20276);
nor U20458 (N_20458,N_20374,N_20281);
nand U20459 (N_20459,N_20343,N_20140);
and U20460 (N_20460,N_20278,N_20308);
xor U20461 (N_20461,N_20348,N_20118);
xor U20462 (N_20462,N_20336,N_20209);
or U20463 (N_20463,N_20122,N_20211);
xnor U20464 (N_20464,N_20217,N_20112);
nand U20465 (N_20465,N_20125,N_20132);
nor U20466 (N_20466,N_20341,N_20280);
nor U20467 (N_20467,N_20192,N_20257);
xor U20468 (N_20468,N_20219,N_20245);
and U20469 (N_20469,N_20131,N_20154);
nor U20470 (N_20470,N_20329,N_20306);
or U20471 (N_20471,N_20208,N_20111);
xor U20472 (N_20472,N_20133,N_20207);
nand U20473 (N_20473,N_20137,N_20195);
or U20474 (N_20474,N_20180,N_20338);
and U20475 (N_20475,N_20332,N_20314);
xnor U20476 (N_20476,N_20167,N_20394);
xnor U20477 (N_20477,N_20178,N_20103);
nor U20478 (N_20478,N_20123,N_20353);
and U20479 (N_20479,N_20210,N_20292);
nand U20480 (N_20480,N_20369,N_20262);
nand U20481 (N_20481,N_20194,N_20106);
nor U20482 (N_20482,N_20359,N_20352);
and U20483 (N_20483,N_20294,N_20222);
nand U20484 (N_20484,N_20113,N_20258);
nor U20485 (N_20485,N_20284,N_20220);
xnor U20486 (N_20486,N_20102,N_20120);
and U20487 (N_20487,N_20150,N_20361);
and U20488 (N_20488,N_20193,N_20339);
nand U20489 (N_20489,N_20134,N_20318);
or U20490 (N_20490,N_20230,N_20107);
nand U20491 (N_20491,N_20289,N_20171);
nand U20492 (N_20492,N_20238,N_20157);
and U20493 (N_20493,N_20114,N_20153);
nand U20494 (N_20494,N_20162,N_20248);
or U20495 (N_20495,N_20158,N_20264);
xor U20496 (N_20496,N_20340,N_20270);
nor U20497 (N_20497,N_20127,N_20228);
or U20498 (N_20498,N_20169,N_20175);
and U20499 (N_20499,N_20342,N_20108);
and U20500 (N_20500,N_20287,N_20334);
nor U20501 (N_20501,N_20185,N_20322);
nand U20502 (N_20502,N_20360,N_20299);
and U20503 (N_20503,N_20366,N_20214);
nand U20504 (N_20504,N_20331,N_20246);
nand U20505 (N_20505,N_20203,N_20190);
and U20506 (N_20506,N_20223,N_20272);
nand U20507 (N_20507,N_20159,N_20204);
nor U20508 (N_20508,N_20115,N_20291);
nor U20509 (N_20509,N_20186,N_20323);
and U20510 (N_20510,N_20213,N_20375);
xnor U20511 (N_20511,N_20283,N_20368);
xor U20512 (N_20512,N_20349,N_20298);
xor U20513 (N_20513,N_20124,N_20234);
xor U20514 (N_20514,N_20389,N_20333);
nand U20515 (N_20515,N_20233,N_20379);
xor U20516 (N_20516,N_20201,N_20350);
xor U20517 (N_20517,N_20396,N_20188);
xor U20518 (N_20518,N_20218,N_20267);
nor U20519 (N_20519,N_20212,N_20370);
nor U20520 (N_20520,N_20265,N_20260);
nor U20521 (N_20521,N_20335,N_20225);
nand U20522 (N_20522,N_20384,N_20176);
xnor U20523 (N_20523,N_20317,N_20345);
nand U20524 (N_20524,N_20129,N_20301);
xor U20525 (N_20525,N_20198,N_20261);
or U20526 (N_20526,N_20255,N_20320);
or U20527 (N_20527,N_20164,N_20371);
nor U20528 (N_20528,N_20356,N_20163);
xnor U20529 (N_20529,N_20197,N_20398);
or U20530 (N_20530,N_20239,N_20266);
or U20531 (N_20531,N_20253,N_20136);
nand U20532 (N_20532,N_20247,N_20321);
and U20533 (N_20533,N_20173,N_20243);
nand U20534 (N_20534,N_20170,N_20355);
and U20535 (N_20535,N_20166,N_20285);
nand U20536 (N_20536,N_20395,N_20130);
nor U20537 (N_20537,N_20268,N_20155);
xnor U20538 (N_20538,N_20273,N_20307);
nor U20539 (N_20539,N_20383,N_20303);
nor U20540 (N_20540,N_20316,N_20119);
nand U20541 (N_20541,N_20152,N_20221);
and U20542 (N_20542,N_20279,N_20390);
nor U20543 (N_20543,N_20277,N_20274);
nand U20544 (N_20544,N_20104,N_20202);
nand U20545 (N_20545,N_20327,N_20388);
and U20546 (N_20546,N_20226,N_20373);
nand U20547 (N_20547,N_20251,N_20311);
or U20548 (N_20548,N_20364,N_20378);
nor U20549 (N_20549,N_20346,N_20161);
and U20550 (N_20550,N_20197,N_20248);
or U20551 (N_20551,N_20235,N_20122);
nor U20552 (N_20552,N_20196,N_20221);
nor U20553 (N_20553,N_20396,N_20364);
nor U20554 (N_20554,N_20285,N_20301);
or U20555 (N_20555,N_20236,N_20192);
or U20556 (N_20556,N_20196,N_20365);
and U20557 (N_20557,N_20358,N_20285);
xor U20558 (N_20558,N_20379,N_20319);
and U20559 (N_20559,N_20234,N_20242);
nor U20560 (N_20560,N_20339,N_20207);
nor U20561 (N_20561,N_20181,N_20158);
or U20562 (N_20562,N_20397,N_20364);
or U20563 (N_20563,N_20299,N_20300);
nand U20564 (N_20564,N_20162,N_20304);
xnor U20565 (N_20565,N_20190,N_20132);
xnor U20566 (N_20566,N_20168,N_20201);
xor U20567 (N_20567,N_20149,N_20115);
nand U20568 (N_20568,N_20251,N_20270);
xor U20569 (N_20569,N_20207,N_20130);
or U20570 (N_20570,N_20387,N_20278);
xor U20571 (N_20571,N_20210,N_20113);
nor U20572 (N_20572,N_20229,N_20113);
and U20573 (N_20573,N_20385,N_20176);
nor U20574 (N_20574,N_20142,N_20139);
and U20575 (N_20575,N_20137,N_20133);
and U20576 (N_20576,N_20334,N_20145);
xor U20577 (N_20577,N_20119,N_20145);
nand U20578 (N_20578,N_20240,N_20163);
and U20579 (N_20579,N_20150,N_20161);
or U20580 (N_20580,N_20324,N_20132);
or U20581 (N_20581,N_20282,N_20193);
nor U20582 (N_20582,N_20100,N_20345);
or U20583 (N_20583,N_20273,N_20136);
and U20584 (N_20584,N_20219,N_20294);
and U20585 (N_20585,N_20303,N_20231);
nor U20586 (N_20586,N_20187,N_20337);
nand U20587 (N_20587,N_20152,N_20272);
and U20588 (N_20588,N_20256,N_20305);
or U20589 (N_20589,N_20246,N_20188);
and U20590 (N_20590,N_20328,N_20284);
nand U20591 (N_20591,N_20158,N_20363);
and U20592 (N_20592,N_20281,N_20394);
and U20593 (N_20593,N_20384,N_20197);
and U20594 (N_20594,N_20111,N_20181);
nor U20595 (N_20595,N_20255,N_20151);
or U20596 (N_20596,N_20260,N_20369);
xnor U20597 (N_20597,N_20385,N_20371);
nand U20598 (N_20598,N_20184,N_20392);
xor U20599 (N_20599,N_20355,N_20360);
and U20600 (N_20600,N_20253,N_20126);
and U20601 (N_20601,N_20126,N_20234);
and U20602 (N_20602,N_20284,N_20152);
xor U20603 (N_20603,N_20276,N_20251);
or U20604 (N_20604,N_20191,N_20281);
nor U20605 (N_20605,N_20241,N_20226);
and U20606 (N_20606,N_20219,N_20153);
or U20607 (N_20607,N_20209,N_20206);
or U20608 (N_20608,N_20262,N_20296);
nor U20609 (N_20609,N_20269,N_20310);
xor U20610 (N_20610,N_20184,N_20270);
and U20611 (N_20611,N_20152,N_20222);
and U20612 (N_20612,N_20225,N_20357);
or U20613 (N_20613,N_20315,N_20161);
nand U20614 (N_20614,N_20324,N_20303);
and U20615 (N_20615,N_20125,N_20239);
and U20616 (N_20616,N_20163,N_20138);
nor U20617 (N_20617,N_20382,N_20154);
and U20618 (N_20618,N_20275,N_20297);
nor U20619 (N_20619,N_20221,N_20388);
or U20620 (N_20620,N_20389,N_20151);
and U20621 (N_20621,N_20123,N_20223);
and U20622 (N_20622,N_20100,N_20391);
or U20623 (N_20623,N_20102,N_20210);
or U20624 (N_20624,N_20167,N_20340);
xnor U20625 (N_20625,N_20389,N_20266);
nor U20626 (N_20626,N_20167,N_20118);
or U20627 (N_20627,N_20318,N_20316);
and U20628 (N_20628,N_20372,N_20263);
and U20629 (N_20629,N_20227,N_20287);
nor U20630 (N_20630,N_20173,N_20338);
nor U20631 (N_20631,N_20376,N_20345);
nor U20632 (N_20632,N_20134,N_20155);
or U20633 (N_20633,N_20199,N_20106);
nor U20634 (N_20634,N_20381,N_20343);
nor U20635 (N_20635,N_20162,N_20389);
or U20636 (N_20636,N_20215,N_20214);
nor U20637 (N_20637,N_20152,N_20228);
nor U20638 (N_20638,N_20352,N_20189);
nor U20639 (N_20639,N_20385,N_20244);
nand U20640 (N_20640,N_20371,N_20156);
nand U20641 (N_20641,N_20154,N_20359);
and U20642 (N_20642,N_20343,N_20399);
or U20643 (N_20643,N_20300,N_20123);
or U20644 (N_20644,N_20295,N_20215);
xnor U20645 (N_20645,N_20271,N_20118);
xnor U20646 (N_20646,N_20246,N_20185);
or U20647 (N_20647,N_20132,N_20329);
nor U20648 (N_20648,N_20212,N_20371);
nand U20649 (N_20649,N_20366,N_20161);
nor U20650 (N_20650,N_20344,N_20308);
xnor U20651 (N_20651,N_20306,N_20301);
and U20652 (N_20652,N_20186,N_20292);
nand U20653 (N_20653,N_20275,N_20303);
and U20654 (N_20654,N_20269,N_20121);
nor U20655 (N_20655,N_20286,N_20202);
nand U20656 (N_20656,N_20321,N_20285);
nand U20657 (N_20657,N_20310,N_20194);
xnor U20658 (N_20658,N_20389,N_20357);
or U20659 (N_20659,N_20252,N_20129);
nand U20660 (N_20660,N_20285,N_20179);
nor U20661 (N_20661,N_20399,N_20166);
and U20662 (N_20662,N_20307,N_20369);
nor U20663 (N_20663,N_20289,N_20396);
or U20664 (N_20664,N_20153,N_20254);
xor U20665 (N_20665,N_20345,N_20342);
and U20666 (N_20666,N_20275,N_20185);
and U20667 (N_20667,N_20207,N_20248);
xnor U20668 (N_20668,N_20222,N_20119);
nor U20669 (N_20669,N_20105,N_20177);
and U20670 (N_20670,N_20291,N_20249);
nor U20671 (N_20671,N_20298,N_20361);
nand U20672 (N_20672,N_20142,N_20193);
xnor U20673 (N_20673,N_20215,N_20349);
or U20674 (N_20674,N_20162,N_20374);
and U20675 (N_20675,N_20299,N_20272);
and U20676 (N_20676,N_20163,N_20321);
xor U20677 (N_20677,N_20383,N_20145);
or U20678 (N_20678,N_20182,N_20187);
nor U20679 (N_20679,N_20266,N_20247);
nand U20680 (N_20680,N_20140,N_20210);
and U20681 (N_20681,N_20310,N_20299);
or U20682 (N_20682,N_20278,N_20380);
or U20683 (N_20683,N_20312,N_20371);
xnor U20684 (N_20684,N_20347,N_20184);
and U20685 (N_20685,N_20305,N_20316);
xnor U20686 (N_20686,N_20398,N_20355);
nor U20687 (N_20687,N_20116,N_20284);
xnor U20688 (N_20688,N_20165,N_20148);
nand U20689 (N_20689,N_20283,N_20388);
nor U20690 (N_20690,N_20290,N_20333);
and U20691 (N_20691,N_20214,N_20176);
or U20692 (N_20692,N_20111,N_20202);
or U20693 (N_20693,N_20239,N_20385);
nand U20694 (N_20694,N_20210,N_20112);
xnor U20695 (N_20695,N_20214,N_20282);
and U20696 (N_20696,N_20211,N_20372);
nand U20697 (N_20697,N_20166,N_20345);
and U20698 (N_20698,N_20230,N_20197);
nor U20699 (N_20699,N_20295,N_20294);
and U20700 (N_20700,N_20595,N_20488);
nor U20701 (N_20701,N_20640,N_20635);
nor U20702 (N_20702,N_20517,N_20431);
and U20703 (N_20703,N_20423,N_20599);
xor U20704 (N_20704,N_20427,N_20471);
xnor U20705 (N_20705,N_20612,N_20472);
or U20706 (N_20706,N_20619,N_20668);
xnor U20707 (N_20707,N_20490,N_20665);
nand U20708 (N_20708,N_20422,N_20634);
nor U20709 (N_20709,N_20499,N_20456);
or U20710 (N_20710,N_20501,N_20560);
nand U20711 (N_20711,N_20406,N_20544);
xnor U20712 (N_20712,N_20643,N_20615);
and U20713 (N_20713,N_20584,N_20420);
or U20714 (N_20714,N_20486,N_20687);
nor U20715 (N_20715,N_20401,N_20575);
nor U20716 (N_20716,N_20625,N_20419);
or U20717 (N_20717,N_20463,N_20551);
nand U20718 (N_20718,N_20411,N_20506);
and U20719 (N_20719,N_20491,N_20571);
and U20720 (N_20720,N_20441,N_20547);
or U20721 (N_20721,N_20636,N_20404);
or U20722 (N_20722,N_20458,N_20695);
nand U20723 (N_20723,N_20641,N_20620);
or U20724 (N_20724,N_20631,N_20493);
nand U20725 (N_20725,N_20526,N_20610);
nand U20726 (N_20726,N_20416,N_20429);
xor U20727 (N_20727,N_20541,N_20597);
nand U20728 (N_20728,N_20662,N_20462);
xnor U20729 (N_20729,N_20459,N_20601);
nor U20730 (N_20730,N_20698,N_20538);
nor U20731 (N_20731,N_20494,N_20572);
or U20732 (N_20732,N_20677,N_20503);
and U20733 (N_20733,N_20696,N_20521);
or U20734 (N_20734,N_20505,N_20661);
nand U20735 (N_20735,N_20626,N_20651);
xor U20736 (N_20736,N_20623,N_20482);
nand U20737 (N_20737,N_20632,N_20469);
xnor U20738 (N_20738,N_20415,N_20583);
and U20739 (N_20739,N_20679,N_20443);
or U20740 (N_20740,N_20699,N_20522);
xor U20741 (N_20741,N_20574,N_20414);
nand U20742 (N_20742,N_20581,N_20566);
nor U20743 (N_20743,N_20524,N_20417);
and U20744 (N_20744,N_20489,N_20559);
or U20745 (N_20745,N_20444,N_20563);
xnor U20746 (N_20746,N_20539,N_20585);
and U20747 (N_20747,N_20564,N_20592);
nor U20748 (N_20748,N_20495,N_20487);
xnor U20749 (N_20749,N_20658,N_20473);
nand U20750 (N_20750,N_20536,N_20629);
or U20751 (N_20751,N_20600,N_20450);
nand U20752 (N_20752,N_20504,N_20447);
or U20753 (N_20753,N_20475,N_20525);
nand U20754 (N_20754,N_20673,N_20652);
and U20755 (N_20755,N_20480,N_20681);
nor U20756 (N_20756,N_20511,N_20680);
nand U20757 (N_20757,N_20694,N_20688);
or U20758 (N_20758,N_20424,N_20582);
nor U20759 (N_20759,N_20693,N_20616);
xor U20760 (N_20760,N_20573,N_20611);
or U20761 (N_20761,N_20607,N_20510);
and U20762 (N_20762,N_20557,N_20622);
and U20763 (N_20763,N_20650,N_20543);
nor U20764 (N_20764,N_20664,N_20654);
or U20765 (N_20765,N_20527,N_20497);
and U20766 (N_20766,N_20613,N_20697);
and U20767 (N_20767,N_20682,N_20466);
xor U20768 (N_20768,N_20580,N_20430);
nand U20769 (N_20769,N_20534,N_20666);
nand U20770 (N_20770,N_20591,N_20418);
or U20771 (N_20771,N_20545,N_20402);
or U20772 (N_20772,N_20644,N_20484);
or U20773 (N_20773,N_20425,N_20530);
nor U20774 (N_20774,N_20608,N_20514);
nor U20775 (N_20775,N_20577,N_20671);
nand U20776 (N_20776,N_20405,N_20535);
xnor U20777 (N_20777,N_20452,N_20553);
and U20778 (N_20778,N_20637,N_20435);
nand U20779 (N_20779,N_20589,N_20542);
or U20780 (N_20780,N_20576,N_20434);
nand U20781 (N_20781,N_20438,N_20691);
xnor U20782 (N_20782,N_20627,N_20642);
xnor U20783 (N_20783,N_20528,N_20529);
or U20784 (N_20784,N_20432,N_20492);
nor U20785 (N_20785,N_20532,N_20579);
or U20786 (N_20786,N_20686,N_20421);
and U20787 (N_20787,N_20485,N_20478);
or U20788 (N_20788,N_20516,N_20467);
nand U20789 (N_20789,N_20437,N_20587);
and U20790 (N_20790,N_20647,N_20550);
nor U20791 (N_20791,N_20606,N_20655);
nand U20792 (N_20792,N_20523,N_20555);
nand U20793 (N_20793,N_20552,N_20477);
or U20794 (N_20794,N_20451,N_20474);
nor U20795 (N_20795,N_20483,N_20609);
or U20796 (N_20796,N_20496,N_20628);
nand U20797 (N_20797,N_20548,N_20624);
nand U20798 (N_20798,N_20412,N_20509);
and U20799 (N_20799,N_20457,N_20449);
nand U20800 (N_20800,N_20596,N_20618);
nor U20801 (N_20801,N_20657,N_20403);
nand U20802 (N_20802,N_20678,N_20461);
and U20803 (N_20803,N_20672,N_20436);
nor U20804 (N_20804,N_20446,N_20659);
and U20805 (N_20805,N_20598,N_20502);
and U20806 (N_20806,N_20500,N_20603);
xor U20807 (N_20807,N_20645,N_20540);
nand U20808 (N_20808,N_20407,N_20633);
xnor U20809 (N_20809,N_20578,N_20683);
or U20810 (N_20810,N_20690,N_20533);
nor U20811 (N_20811,N_20413,N_20605);
xor U20812 (N_20812,N_20685,N_20684);
nor U20813 (N_20813,N_20400,N_20433);
and U20814 (N_20814,N_20586,N_20507);
nand U20815 (N_20815,N_20537,N_20676);
nor U20816 (N_20816,N_20439,N_20428);
nand U20817 (N_20817,N_20565,N_20630);
nor U20818 (N_20818,N_20508,N_20692);
xor U20819 (N_20819,N_20570,N_20519);
nand U20820 (N_20820,N_20465,N_20674);
xor U20821 (N_20821,N_20588,N_20410);
xnor U20822 (N_20822,N_20476,N_20454);
or U20823 (N_20823,N_20667,N_20669);
nor U20824 (N_20824,N_20518,N_20554);
xor U20825 (N_20825,N_20513,N_20442);
nand U20826 (N_20826,N_20653,N_20408);
nor U20827 (N_20827,N_20512,N_20549);
or U20828 (N_20828,N_20621,N_20569);
nor U20829 (N_20829,N_20594,N_20498);
nand U20830 (N_20830,N_20479,N_20481);
xor U20831 (N_20831,N_20663,N_20648);
xnor U20832 (N_20832,N_20593,N_20660);
and U20833 (N_20833,N_20445,N_20590);
or U20834 (N_20834,N_20520,N_20460);
nor U20835 (N_20835,N_20675,N_20638);
or U20836 (N_20836,N_20440,N_20426);
nor U20837 (N_20837,N_20561,N_20567);
nand U20838 (N_20838,N_20453,N_20470);
nand U20839 (N_20839,N_20646,N_20604);
and U20840 (N_20840,N_20531,N_20562);
nor U20841 (N_20841,N_20556,N_20448);
or U20842 (N_20842,N_20649,N_20614);
nand U20843 (N_20843,N_20568,N_20468);
xor U20844 (N_20844,N_20656,N_20515);
and U20845 (N_20845,N_20455,N_20464);
and U20846 (N_20846,N_20409,N_20617);
nor U20847 (N_20847,N_20546,N_20558);
xnor U20848 (N_20848,N_20639,N_20689);
or U20849 (N_20849,N_20670,N_20602);
nand U20850 (N_20850,N_20546,N_20468);
nand U20851 (N_20851,N_20631,N_20562);
or U20852 (N_20852,N_20525,N_20485);
nand U20853 (N_20853,N_20484,N_20686);
and U20854 (N_20854,N_20604,N_20632);
xor U20855 (N_20855,N_20607,N_20605);
nand U20856 (N_20856,N_20497,N_20565);
nor U20857 (N_20857,N_20449,N_20614);
or U20858 (N_20858,N_20408,N_20691);
nand U20859 (N_20859,N_20612,N_20609);
nand U20860 (N_20860,N_20412,N_20630);
nor U20861 (N_20861,N_20569,N_20600);
nand U20862 (N_20862,N_20681,N_20485);
nor U20863 (N_20863,N_20652,N_20578);
or U20864 (N_20864,N_20633,N_20667);
nor U20865 (N_20865,N_20460,N_20420);
nand U20866 (N_20866,N_20554,N_20405);
nor U20867 (N_20867,N_20415,N_20616);
nor U20868 (N_20868,N_20536,N_20617);
nor U20869 (N_20869,N_20599,N_20539);
nor U20870 (N_20870,N_20496,N_20528);
and U20871 (N_20871,N_20460,N_20596);
nor U20872 (N_20872,N_20408,N_20554);
nand U20873 (N_20873,N_20421,N_20427);
and U20874 (N_20874,N_20661,N_20556);
xnor U20875 (N_20875,N_20543,N_20596);
xnor U20876 (N_20876,N_20467,N_20532);
nand U20877 (N_20877,N_20665,N_20466);
or U20878 (N_20878,N_20437,N_20639);
xor U20879 (N_20879,N_20448,N_20650);
nand U20880 (N_20880,N_20450,N_20653);
nand U20881 (N_20881,N_20647,N_20678);
xor U20882 (N_20882,N_20565,N_20599);
nand U20883 (N_20883,N_20545,N_20430);
or U20884 (N_20884,N_20660,N_20457);
nor U20885 (N_20885,N_20659,N_20419);
nand U20886 (N_20886,N_20648,N_20530);
and U20887 (N_20887,N_20465,N_20683);
or U20888 (N_20888,N_20514,N_20560);
and U20889 (N_20889,N_20580,N_20491);
nand U20890 (N_20890,N_20440,N_20526);
or U20891 (N_20891,N_20514,N_20481);
nand U20892 (N_20892,N_20483,N_20560);
nor U20893 (N_20893,N_20513,N_20506);
nor U20894 (N_20894,N_20404,N_20475);
nand U20895 (N_20895,N_20422,N_20596);
and U20896 (N_20896,N_20649,N_20543);
nor U20897 (N_20897,N_20637,N_20413);
nand U20898 (N_20898,N_20402,N_20490);
nor U20899 (N_20899,N_20592,N_20683);
nor U20900 (N_20900,N_20657,N_20410);
and U20901 (N_20901,N_20557,N_20554);
nor U20902 (N_20902,N_20524,N_20648);
or U20903 (N_20903,N_20434,N_20647);
nor U20904 (N_20904,N_20436,N_20491);
and U20905 (N_20905,N_20423,N_20403);
xnor U20906 (N_20906,N_20414,N_20502);
or U20907 (N_20907,N_20448,N_20590);
nand U20908 (N_20908,N_20460,N_20685);
or U20909 (N_20909,N_20501,N_20547);
xor U20910 (N_20910,N_20668,N_20591);
nand U20911 (N_20911,N_20447,N_20561);
xor U20912 (N_20912,N_20616,N_20528);
xor U20913 (N_20913,N_20501,N_20520);
nand U20914 (N_20914,N_20517,N_20661);
or U20915 (N_20915,N_20537,N_20446);
or U20916 (N_20916,N_20621,N_20518);
and U20917 (N_20917,N_20588,N_20523);
and U20918 (N_20918,N_20572,N_20655);
xor U20919 (N_20919,N_20421,N_20586);
or U20920 (N_20920,N_20554,N_20534);
and U20921 (N_20921,N_20570,N_20422);
xnor U20922 (N_20922,N_20523,N_20455);
nor U20923 (N_20923,N_20507,N_20640);
and U20924 (N_20924,N_20438,N_20453);
and U20925 (N_20925,N_20588,N_20486);
nor U20926 (N_20926,N_20568,N_20555);
nor U20927 (N_20927,N_20504,N_20457);
nor U20928 (N_20928,N_20420,N_20637);
and U20929 (N_20929,N_20533,N_20511);
xnor U20930 (N_20930,N_20532,N_20517);
xnor U20931 (N_20931,N_20601,N_20524);
nor U20932 (N_20932,N_20565,N_20427);
nor U20933 (N_20933,N_20675,N_20699);
nor U20934 (N_20934,N_20674,N_20435);
and U20935 (N_20935,N_20409,N_20436);
and U20936 (N_20936,N_20431,N_20672);
nor U20937 (N_20937,N_20466,N_20609);
xnor U20938 (N_20938,N_20649,N_20528);
xnor U20939 (N_20939,N_20477,N_20436);
nor U20940 (N_20940,N_20568,N_20556);
or U20941 (N_20941,N_20467,N_20459);
or U20942 (N_20942,N_20445,N_20638);
xor U20943 (N_20943,N_20632,N_20520);
and U20944 (N_20944,N_20573,N_20566);
and U20945 (N_20945,N_20646,N_20638);
or U20946 (N_20946,N_20675,N_20687);
nor U20947 (N_20947,N_20436,N_20503);
nand U20948 (N_20948,N_20636,N_20444);
and U20949 (N_20949,N_20475,N_20527);
xnor U20950 (N_20950,N_20693,N_20634);
nor U20951 (N_20951,N_20593,N_20616);
xnor U20952 (N_20952,N_20453,N_20660);
or U20953 (N_20953,N_20463,N_20565);
or U20954 (N_20954,N_20668,N_20464);
nor U20955 (N_20955,N_20630,N_20498);
xor U20956 (N_20956,N_20676,N_20446);
xnor U20957 (N_20957,N_20511,N_20653);
xnor U20958 (N_20958,N_20654,N_20686);
or U20959 (N_20959,N_20638,N_20579);
or U20960 (N_20960,N_20616,N_20648);
and U20961 (N_20961,N_20657,N_20502);
and U20962 (N_20962,N_20503,N_20431);
xor U20963 (N_20963,N_20618,N_20585);
and U20964 (N_20964,N_20490,N_20554);
nor U20965 (N_20965,N_20510,N_20495);
or U20966 (N_20966,N_20523,N_20412);
and U20967 (N_20967,N_20541,N_20693);
nand U20968 (N_20968,N_20590,N_20637);
nand U20969 (N_20969,N_20410,N_20531);
and U20970 (N_20970,N_20664,N_20554);
nor U20971 (N_20971,N_20518,N_20609);
and U20972 (N_20972,N_20577,N_20698);
and U20973 (N_20973,N_20426,N_20626);
xnor U20974 (N_20974,N_20645,N_20631);
and U20975 (N_20975,N_20545,N_20502);
nand U20976 (N_20976,N_20600,N_20445);
xor U20977 (N_20977,N_20437,N_20455);
and U20978 (N_20978,N_20601,N_20547);
or U20979 (N_20979,N_20442,N_20426);
xnor U20980 (N_20980,N_20633,N_20430);
or U20981 (N_20981,N_20596,N_20457);
xor U20982 (N_20982,N_20564,N_20565);
xor U20983 (N_20983,N_20521,N_20506);
xor U20984 (N_20984,N_20435,N_20503);
nor U20985 (N_20985,N_20568,N_20506);
and U20986 (N_20986,N_20610,N_20405);
nand U20987 (N_20987,N_20649,N_20616);
or U20988 (N_20988,N_20415,N_20479);
or U20989 (N_20989,N_20697,N_20696);
nor U20990 (N_20990,N_20534,N_20636);
xor U20991 (N_20991,N_20618,N_20530);
or U20992 (N_20992,N_20682,N_20608);
and U20993 (N_20993,N_20570,N_20432);
nand U20994 (N_20994,N_20686,N_20540);
or U20995 (N_20995,N_20664,N_20665);
nor U20996 (N_20996,N_20536,N_20596);
or U20997 (N_20997,N_20571,N_20527);
nor U20998 (N_20998,N_20418,N_20590);
nand U20999 (N_20999,N_20695,N_20537);
nor U21000 (N_21000,N_20973,N_20870);
or U21001 (N_21001,N_20865,N_20788);
nand U21002 (N_21002,N_20827,N_20730);
and U21003 (N_21003,N_20928,N_20960);
or U21004 (N_21004,N_20842,N_20716);
and U21005 (N_21005,N_20706,N_20725);
or U21006 (N_21006,N_20976,N_20805);
nand U21007 (N_21007,N_20894,N_20999);
and U21008 (N_21008,N_20708,N_20944);
nor U21009 (N_21009,N_20906,N_20850);
nor U21010 (N_21010,N_20834,N_20811);
and U21011 (N_21011,N_20790,N_20801);
nor U21012 (N_21012,N_20829,N_20777);
nor U21013 (N_21013,N_20797,N_20998);
nand U21014 (N_21014,N_20779,N_20830);
or U21015 (N_21015,N_20980,N_20953);
or U21016 (N_21016,N_20733,N_20896);
nor U21017 (N_21017,N_20971,N_20886);
nor U21018 (N_21018,N_20993,N_20796);
xor U21019 (N_21019,N_20852,N_20726);
nor U21020 (N_21020,N_20970,N_20756);
nor U21021 (N_21021,N_20914,N_20718);
nand U21022 (N_21022,N_20774,N_20964);
nand U21023 (N_21023,N_20957,N_20715);
xor U21024 (N_21024,N_20893,N_20904);
and U21025 (N_21025,N_20739,N_20736);
xnor U21026 (N_21026,N_20924,N_20901);
and U21027 (N_21027,N_20895,N_20758);
and U21028 (N_21028,N_20798,N_20744);
and U21029 (N_21029,N_20804,N_20968);
or U21030 (N_21030,N_20961,N_20866);
xnor U21031 (N_21031,N_20782,N_20878);
nor U21032 (N_21032,N_20907,N_20818);
xor U21033 (N_21033,N_20781,N_20713);
nand U21034 (N_21034,N_20859,N_20823);
and U21035 (N_21035,N_20753,N_20707);
and U21036 (N_21036,N_20986,N_20768);
and U21037 (N_21037,N_20737,N_20995);
and U21038 (N_21038,N_20919,N_20989);
xnor U21039 (N_21039,N_20812,N_20892);
xnor U21040 (N_21040,N_20845,N_20831);
xnor U21041 (N_21041,N_20888,N_20792);
nor U21042 (N_21042,N_20764,N_20701);
xnor U21043 (N_21043,N_20824,N_20742);
and U21044 (N_21044,N_20871,N_20860);
or U21045 (N_21045,N_20856,N_20988);
xnor U21046 (N_21046,N_20990,N_20916);
nor U21047 (N_21047,N_20900,N_20817);
and U21048 (N_21048,N_20826,N_20727);
nand U21049 (N_21049,N_20939,N_20837);
or U21050 (N_21050,N_20729,N_20816);
and U21051 (N_21051,N_20740,N_20940);
and U21052 (N_21052,N_20984,N_20841);
nor U21053 (N_21053,N_20748,N_20926);
or U21054 (N_21054,N_20853,N_20931);
nor U21055 (N_21055,N_20905,N_20952);
and U21056 (N_21056,N_20757,N_20825);
nor U21057 (N_21057,N_20815,N_20941);
xnor U21058 (N_21058,N_20942,N_20963);
xnor U21059 (N_21059,N_20955,N_20806);
nand U21060 (N_21060,N_20854,N_20884);
nor U21061 (N_21061,N_20843,N_20759);
nor U21062 (N_21062,N_20734,N_20975);
nor U21063 (N_21063,N_20923,N_20938);
nand U21064 (N_21064,N_20720,N_20956);
or U21065 (N_21065,N_20863,N_20991);
xnor U21066 (N_21066,N_20763,N_20920);
xnor U21067 (N_21067,N_20762,N_20838);
and U21068 (N_21068,N_20839,N_20754);
nand U21069 (N_21069,N_20891,N_20722);
or U21070 (N_21070,N_20765,N_20703);
nor U21071 (N_21071,N_20848,N_20925);
nor U21072 (N_21072,N_20723,N_20962);
and U21073 (N_21073,N_20709,N_20783);
or U21074 (N_21074,N_20704,N_20819);
xor U21075 (N_21075,N_20844,N_20857);
nand U21076 (N_21076,N_20885,N_20799);
and U21077 (N_21077,N_20800,N_20840);
nor U21078 (N_21078,N_20882,N_20743);
and U21079 (N_21079,N_20977,N_20933);
and U21080 (N_21080,N_20712,N_20769);
and U21081 (N_21081,N_20867,N_20809);
nand U21082 (N_21082,N_20847,N_20864);
and U21083 (N_21083,N_20773,N_20994);
or U21084 (N_21084,N_20717,N_20802);
and U21085 (N_21085,N_20710,N_20992);
nand U21086 (N_21086,N_20851,N_20948);
nand U21087 (N_21087,N_20858,N_20947);
nand U21088 (N_21088,N_20965,N_20775);
nand U21089 (N_21089,N_20833,N_20776);
or U21090 (N_21090,N_20982,N_20897);
xnor U21091 (N_21091,N_20814,N_20903);
xor U21092 (N_21092,N_20930,N_20922);
xor U21093 (N_21093,N_20705,N_20789);
xor U21094 (N_21094,N_20969,N_20978);
nor U21095 (N_21095,N_20784,N_20700);
xnor U21096 (N_21096,N_20750,N_20937);
or U21097 (N_21097,N_20849,N_20836);
and U21098 (N_21098,N_20902,N_20951);
nand U21099 (N_21099,N_20735,N_20927);
nor U21100 (N_21100,N_20945,N_20910);
and U21101 (N_21101,N_20741,N_20912);
and U21102 (N_21102,N_20771,N_20972);
or U21103 (N_21103,N_20996,N_20898);
and U21104 (N_21104,N_20890,N_20909);
nand U21105 (N_21105,N_20760,N_20881);
xnor U21106 (N_21106,N_20887,N_20810);
nor U21107 (N_21107,N_20807,N_20950);
and U21108 (N_21108,N_20997,N_20936);
nand U21109 (N_21109,N_20832,N_20767);
nand U21110 (N_21110,N_20808,N_20728);
and U21111 (N_21111,N_20846,N_20946);
and U21112 (N_21112,N_20943,N_20778);
nor U21113 (N_21113,N_20772,N_20855);
and U21114 (N_21114,N_20822,N_20949);
and U21115 (N_21115,N_20985,N_20835);
xnor U21116 (N_21116,N_20869,N_20731);
nor U21117 (N_21117,N_20958,N_20934);
xnor U21118 (N_21118,N_20921,N_20821);
or U21119 (N_21119,N_20981,N_20791);
nand U21120 (N_21120,N_20786,N_20861);
or U21121 (N_21121,N_20794,N_20785);
nor U21122 (N_21122,N_20966,N_20702);
or U21123 (N_21123,N_20787,N_20880);
nor U21124 (N_21124,N_20908,N_20766);
xor U21125 (N_21125,N_20987,N_20780);
or U21126 (N_21126,N_20724,N_20974);
nand U21127 (N_21127,N_20913,N_20876);
and U21128 (N_21128,N_20874,N_20917);
nor U21129 (N_21129,N_20747,N_20803);
and U21130 (N_21130,N_20746,N_20918);
and U21131 (N_21131,N_20883,N_20983);
and U21132 (N_21132,N_20751,N_20929);
xor U21133 (N_21133,N_20879,N_20979);
nand U21134 (N_21134,N_20732,N_20795);
nand U21135 (N_21135,N_20862,N_20872);
nand U21136 (N_21136,N_20813,N_20935);
nand U21137 (N_21137,N_20967,N_20954);
nor U21138 (N_21138,N_20820,N_20752);
or U21139 (N_21139,N_20745,N_20711);
nor U21140 (N_21140,N_20738,N_20714);
xnor U21141 (N_21141,N_20877,N_20755);
nand U21142 (N_21142,N_20899,N_20932);
nand U21143 (N_21143,N_20761,N_20828);
xnor U21144 (N_21144,N_20749,N_20873);
and U21145 (N_21145,N_20875,N_20793);
nand U21146 (N_21146,N_20911,N_20770);
nor U21147 (N_21147,N_20915,N_20719);
xnor U21148 (N_21148,N_20721,N_20889);
and U21149 (N_21149,N_20959,N_20868);
or U21150 (N_21150,N_20811,N_20764);
or U21151 (N_21151,N_20978,N_20902);
nand U21152 (N_21152,N_20927,N_20738);
nor U21153 (N_21153,N_20884,N_20754);
nor U21154 (N_21154,N_20815,N_20887);
xnor U21155 (N_21155,N_20875,N_20775);
xor U21156 (N_21156,N_20801,N_20775);
or U21157 (N_21157,N_20901,N_20820);
and U21158 (N_21158,N_20871,N_20836);
or U21159 (N_21159,N_20761,N_20977);
nand U21160 (N_21160,N_20979,N_20787);
and U21161 (N_21161,N_20798,N_20725);
or U21162 (N_21162,N_20891,N_20831);
and U21163 (N_21163,N_20724,N_20922);
or U21164 (N_21164,N_20863,N_20821);
nor U21165 (N_21165,N_20875,N_20761);
nor U21166 (N_21166,N_20817,N_20757);
xor U21167 (N_21167,N_20963,N_20904);
nand U21168 (N_21168,N_20945,N_20840);
or U21169 (N_21169,N_20847,N_20708);
nand U21170 (N_21170,N_20994,N_20898);
xnor U21171 (N_21171,N_20710,N_20967);
and U21172 (N_21172,N_20802,N_20781);
or U21173 (N_21173,N_20700,N_20980);
xnor U21174 (N_21174,N_20911,N_20947);
or U21175 (N_21175,N_20920,N_20970);
or U21176 (N_21176,N_20966,N_20796);
and U21177 (N_21177,N_20936,N_20750);
nor U21178 (N_21178,N_20767,N_20799);
nor U21179 (N_21179,N_20818,N_20796);
xnor U21180 (N_21180,N_20781,N_20721);
xor U21181 (N_21181,N_20971,N_20727);
or U21182 (N_21182,N_20948,N_20791);
or U21183 (N_21183,N_20716,N_20992);
nor U21184 (N_21184,N_20942,N_20923);
nor U21185 (N_21185,N_20809,N_20709);
nor U21186 (N_21186,N_20765,N_20894);
nor U21187 (N_21187,N_20924,N_20902);
and U21188 (N_21188,N_20836,N_20893);
nand U21189 (N_21189,N_20932,N_20884);
xnor U21190 (N_21190,N_20816,N_20960);
nand U21191 (N_21191,N_20721,N_20958);
xnor U21192 (N_21192,N_20869,N_20799);
xor U21193 (N_21193,N_20863,N_20792);
or U21194 (N_21194,N_20788,N_20939);
nor U21195 (N_21195,N_20710,N_20960);
xnor U21196 (N_21196,N_20702,N_20775);
nor U21197 (N_21197,N_20738,N_20719);
nand U21198 (N_21198,N_20989,N_20731);
nor U21199 (N_21199,N_20981,N_20704);
nor U21200 (N_21200,N_20893,N_20809);
nor U21201 (N_21201,N_20856,N_20835);
nand U21202 (N_21202,N_20702,N_20718);
nand U21203 (N_21203,N_20884,N_20938);
or U21204 (N_21204,N_20961,N_20998);
xnor U21205 (N_21205,N_20881,N_20947);
and U21206 (N_21206,N_20847,N_20929);
xnor U21207 (N_21207,N_20931,N_20718);
and U21208 (N_21208,N_20790,N_20864);
or U21209 (N_21209,N_20937,N_20781);
or U21210 (N_21210,N_20970,N_20738);
and U21211 (N_21211,N_20980,N_20718);
or U21212 (N_21212,N_20935,N_20870);
xnor U21213 (N_21213,N_20836,N_20837);
xor U21214 (N_21214,N_20993,N_20727);
or U21215 (N_21215,N_20920,N_20792);
xor U21216 (N_21216,N_20997,N_20896);
nor U21217 (N_21217,N_20801,N_20896);
nand U21218 (N_21218,N_20735,N_20775);
or U21219 (N_21219,N_20741,N_20864);
xnor U21220 (N_21220,N_20734,N_20959);
xor U21221 (N_21221,N_20810,N_20958);
or U21222 (N_21222,N_20722,N_20958);
nand U21223 (N_21223,N_20910,N_20922);
or U21224 (N_21224,N_20882,N_20899);
xor U21225 (N_21225,N_20934,N_20769);
or U21226 (N_21226,N_20856,N_20916);
xor U21227 (N_21227,N_20703,N_20825);
and U21228 (N_21228,N_20919,N_20750);
xor U21229 (N_21229,N_20944,N_20870);
xor U21230 (N_21230,N_20850,N_20920);
nor U21231 (N_21231,N_20918,N_20927);
and U21232 (N_21232,N_20809,N_20965);
and U21233 (N_21233,N_20998,N_20906);
xnor U21234 (N_21234,N_20807,N_20949);
and U21235 (N_21235,N_20772,N_20846);
and U21236 (N_21236,N_20980,N_20829);
or U21237 (N_21237,N_20948,N_20970);
and U21238 (N_21238,N_20866,N_20734);
nor U21239 (N_21239,N_20940,N_20764);
or U21240 (N_21240,N_20759,N_20707);
or U21241 (N_21241,N_20808,N_20719);
or U21242 (N_21242,N_20945,N_20744);
and U21243 (N_21243,N_20768,N_20932);
nor U21244 (N_21244,N_20787,N_20804);
nor U21245 (N_21245,N_20817,N_20761);
nor U21246 (N_21246,N_20834,N_20857);
or U21247 (N_21247,N_20850,N_20710);
or U21248 (N_21248,N_20889,N_20700);
or U21249 (N_21249,N_20789,N_20715);
nand U21250 (N_21250,N_20735,N_20828);
and U21251 (N_21251,N_20925,N_20868);
nor U21252 (N_21252,N_20999,N_20958);
nor U21253 (N_21253,N_20879,N_20720);
nand U21254 (N_21254,N_20851,N_20879);
nand U21255 (N_21255,N_20983,N_20822);
nor U21256 (N_21256,N_20904,N_20715);
and U21257 (N_21257,N_20805,N_20821);
nor U21258 (N_21258,N_20732,N_20817);
or U21259 (N_21259,N_20895,N_20897);
nand U21260 (N_21260,N_20841,N_20825);
and U21261 (N_21261,N_20704,N_20886);
xor U21262 (N_21262,N_20714,N_20769);
nor U21263 (N_21263,N_20804,N_20986);
nor U21264 (N_21264,N_20837,N_20774);
nor U21265 (N_21265,N_20706,N_20714);
and U21266 (N_21266,N_20758,N_20714);
nor U21267 (N_21267,N_20932,N_20784);
or U21268 (N_21268,N_20782,N_20930);
xnor U21269 (N_21269,N_20888,N_20879);
and U21270 (N_21270,N_20804,N_20752);
and U21271 (N_21271,N_20878,N_20785);
and U21272 (N_21272,N_20982,N_20779);
xnor U21273 (N_21273,N_20807,N_20831);
nand U21274 (N_21274,N_20812,N_20700);
xor U21275 (N_21275,N_20799,N_20946);
xor U21276 (N_21276,N_20874,N_20745);
nand U21277 (N_21277,N_20782,N_20953);
nor U21278 (N_21278,N_20776,N_20904);
xnor U21279 (N_21279,N_20758,N_20820);
nor U21280 (N_21280,N_20743,N_20860);
or U21281 (N_21281,N_20809,N_20795);
xor U21282 (N_21282,N_20837,N_20846);
or U21283 (N_21283,N_20788,N_20922);
xnor U21284 (N_21284,N_20802,N_20996);
nand U21285 (N_21285,N_20846,N_20955);
nor U21286 (N_21286,N_20960,N_20856);
or U21287 (N_21287,N_20825,N_20820);
or U21288 (N_21288,N_20946,N_20908);
or U21289 (N_21289,N_20782,N_20859);
nand U21290 (N_21290,N_20762,N_20940);
xor U21291 (N_21291,N_20760,N_20780);
nor U21292 (N_21292,N_20900,N_20743);
xor U21293 (N_21293,N_20799,N_20822);
nand U21294 (N_21294,N_20937,N_20832);
nand U21295 (N_21295,N_20909,N_20901);
nand U21296 (N_21296,N_20970,N_20741);
or U21297 (N_21297,N_20978,N_20859);
nand U21298 (N_21298,N_20882,N_20980);
nand U21299 (N_21299,N_20864,N_20950);
xnor U21300 (N_21300,N_21126,N_21251);
and U21301 (N_21301,N_21068,N_21023);
and U21302 (N_21302,N_21152,N_21008);
or U21303 (N_21303,N_21276,N_21039);
and U21304 (N_21304,N_21018,N_21278);
xor U21305 (N_21305,N_21121,N_21195);
and U21306 (N_21306,N_21258,N_21167);
xor U21307 (N_21307,N_21200,N_21024);
or U21308 (N_21308,N_21299,N_21004);
xnor U21309 (N_21309,N_21135,N_21203);
and U21310 (N_21310,N_21230,N_21030);
xor U21311 (N_21311,N_21185,N_21127);
nand U21312 (N_21312,N_21026,N_21058);
nor U21313 (N_21313,N_21071,N_21160);
and U21314 (N_21314,N_21297,N_21257);
xor U21315 (N_21315,N_21218,N_21273);
or U21316 (N_21316,N_21138,N_21074);
and U21317 (N_21317,N_21097,N_21099);
xor U21318 (N_21318,N_21022,N_21002);
nand U21319 (N_21319,N_21104,N_21182);
nor U21320 (N_21320,N_21073,N_21249);
nor U21321 (N_21321,N_21226,N_21267);
or U21322 (N_21322,N_21107,N_21217);
and U21323 (N_21323,N_21063,N_21198);
xnor U21324 (N_21324,N_21268,N_21043);
nand U21325 (N_21325,N_21188,N_21298);
and U21326 (N_21326,N_21046,N_21227);
xnor U21327 (N_21327,N_21211,N_21283);
or U21328 (N_21328,N_21146,N_21184);
nand U21329 (N_21329,N_21165,N_21037);
nand U21330 (N_21330,N_21168,N_21262);
or U21331 (N_21331,N_21001,N_21095);
or U21332 (N_21332,N_21212,N_21153);
xor U21333 (N_21333,N_21052,N_21154);
xnor U21334 (N_21334,N_21035,N_21114);
and U21335 (N_21335,N_21285,N_21162);
xor U21336 (N_21336,N_21089,N_21000);
nand U21337 (N_21337,N_21072,N_21122);
nor U21338 (N_21338,N_21124,N_21157);
nor U21339 (N_21339,N_21156,N_21096);
nand U21340 (N_21340,N_21291,N_21134);
xor U21341 (N_21341,N_21028,N_21295);
or U21342 (N_21342,N_21236,N_21274);
xor U21343 (N_21343,N_21256,N_21192);
xnor U21344 (N_21344,N_21080,N_21110);
nor U21345 (N_21345,N_21202,N_21091);
nand U21346 (N_21346,N_21150,N_21141);
and U21347 (N_21347,N_21147,N_21120);
nor U21348 (N_21348,N_21244,N_21151);
xor U21349 (N_21349,N_21207,N_21209);
and U21350 (N_21350,N_21014,N_21036);
and U21351 (N_21351,N_21243,N_21288);
nand U21352 (N_21352,N_21102,N_21189);
or U21353 (N_21353,N_21015,N_21136);
nand U21354 (N_21354,N_21021,N_21266);
or U21355 (N_21355,N_21197,N_21186);
or U21356 (N_21356,N_21050,N_21245);
nor U21357 (N_21357,N_21223,N_21016);
nand U21358 (N_21358,N_21264,N_21215);
or U21359 (N_21359,N_21289,N_21020);
nor U21360 (N_21360,N_21060,N_21142);
and U21361 (N_21361,N_21204,N_21077);
and U21362 (N_21362,N_21092,N_21235);
or U21363 (N_21363,N_21086,N_21287);
nand U21364 (N_21364,N_21233,N_21131);
nand U21365 (N_21365,N_21144,N_21048);
or U21366 (N_21366,N_21201,N_21280);
nor U21367 (N_21367,N_21208,N_21100);
xnor U21368 (N_21368,N_21234,N_21017);
xnor U21369 (N_21369,N_21025,N_21158);
xor U21370 (N_21370,N_21159,N_21232);
nand U21371 (N_21371,N_21224,N_21190);
nor U21372 (N_21372,N_21255,N_21260);
xnor U21373 (N_21373,N_21065,N_21140);
and U21374 (N_21374,N_21270,N_21205);
nand U21375 (N_21375,N_21132,N_21051);
or U21376 (N_21376,N_21139,N_21174);
or U21377 (N_21377,N_21179,N_21148);
xor U21378 (N_21378,N_21061,N_21076);
xnor U21379 (N_21379,N_21173,N_21161);
xnor U21380 (N_21380,N_21237,N_21279);
and U21381 (N_21381,N_21054,N_21041);
or U21382 (N_21382,N_21254,N_21253);
or U21383 (N_21383,N_21067,N_21115);
nor U21384 (N_21384,N_21199,N_21293);
and U21385 (N_21385,N_21261,N_21166);
and U21386 (N_21386,N_21281,N_21118);
nand U21387 (N_21387,N_21130,N_21032);
xor U21388 (N_21388,N_21292,N_21013);
or U21389 (N_21389,N_21175,N_21210);
nor U21390 (N_21390,N_21010,N_21047);
or U21391 (N_21391,N_21213,N_21216);
nand U21392 (N_21392,N_21128,N_21040);
nand U21393 (N_21393,N_21178,N_21033);
and U21394 (N_21394,N_21087,N_21075);
xor U21395 (N_21395,N_21084,N_21059);
and U21396 (N_21396,N_21214,N_21064);
or U21397 (N_21397,N_21206,N_21240);
and U21398 (N_21398,N_21006,N_21094);
or U21399 (N_21399,N_21108,N_21106);
and U21400 (N_21400,N_21225,N_21252);
or U21401 (N_21401,N_21183,N_21241);
nor U21402 (N_21402,N_21117,N_21238);
xnor U21403 (N_21403,N_21133,N_21042);
xor U21404 (N_21404,N_21066,N_21123);
and U21405 (N_21405,N_21078,N_21044);
and U21406 (N_21406,N_21088,N_21027);
or U21407 (N_21407,N_21019,N_21222);
or U21408 (N_21408,N_21221,N_21247);
or U21409 (N_21409,N_21070,N_21105);
and U21410 (N_21410,N_21263,N_21176);
nor U21411 (N_21411,N_21231,N_21220);
and U21412 (N_21412,N_21271,N_21145);
nor U21413 (N_21413,N_21265,N_21053);
xnor U21414 (N_21414,N_21103,N_21143);
nand U21415 (N_21415,N_21284,N_21093);
or U21416 (N_21416,N_21194,N_21045);
nand U21417 (N_21417,N_21034,N_21009);
nor U21418 (N_21418,N_21219,N_21031);
or U21419 (N_21419,N_21277,N_21187);
nor U21420 (N_21420,N_21116,N_21125);
nor U21421 (N_21421,N_21294,N_21012);
xnor U21422 (N_21422,N_21079,N_21113);
nor U21423 (N_21423,N_21193,N_21191);
or U21424 (N_21424,N_21164,N_21282);
and U21425 (N_21425,N_21081,N_21228);
or U21426 (N_21426,N_21239,N_21011);
xor U21427 (N_21427,N_21119,N_21038);
and U21428 (N_21428,N_21163,N_21109);
nand U21429 (N_21429,N_21171,N_21055);
nand U21430 (N_21430,N_21246,N_21180);
and U21431 (N_21431,N_21137,N_21098);
xnor U21432 (N_21432,N_21111,N_21062);
xnor U21433 (N_21433,N_21069,N_21275);
xnor U21434 (N_21434,N_21286,N_21085);
or U21435 (N_21435,N_21296,N_21029);
nor U21436 (N_21436,N_21242,N_21248);
and U21437 (N_21437,N_21005,N_21181);
nor U21438 (N_21438,N_21083,N_21090);
xnor U21439 (N_21439,N_21155,N_21229);
or U21440 (N_21440,N_21196,N_21250);
nand U21441 (N_21441,N_21177,N_21112);
xor U21442 (N_21442,N_21272,N_21149);
xor U21443 (N_21443,N_21056,N_21170);
nor U21444 (N_21444,N_21259,N_21172);
or U21445 (N_21445,N_21169,N_21290);
nand U21446 (N_21446,N_21129,N_21057);
nor U21447 (N_21447,N_21049,N_21082);
or U21448 (N_21448,N_21003,N_21101);
xnor U21449 (N_21449,N_21269,N_21007);
or U21450 (N_21450,N_21099,N_21140);
nand U21451 (N_21451,N_21099,N_21142);
xor U21452 (N_21452,N_21239,N_21105);
and U21453 (N_21453,N_21027,N_21107);
or U21454 (N_21454,N_21266,N_21023);
xnor U21455 (N_21455,N_21022,N_21161);
or U21456 (N_21456,N_21165,N_21049);
or U21457 (N_21457,N_21297,N_21265);
or U21458 (N_21458,N_21263,N_21175);
or U21459 (N_21459,N_21096,N_21018);
xnor U21460 (N_21460,N_21277,N_21152);
nor U21461 (N_21461,N_21214,N_21021);
and U21462 (N_21462,N_21295,N_21206);
nor U21463 (N_21463,N_21041,N_21033);
nor U21464 (N_21464,N_21260,N_21158);
nor U21465 (N_21465,N_21147,N_21183);
and U21466 (N_21466,N_21136,N_21250);
and U21467 (N_21467,N_21188,N_21235);
xnor U21468 (N_21468,N_21004,N_21016);
xnor U21469 (N_21469,N_21266,N_21055);
nor U21470 (N_21470,N_21212,N_21074);
and U21471 (N_21471,N_21205,N_21029);
and U21472 (N_21472,N_21116,N_21207);
nand U21473 (N_21473,N_21024,N_21030);
nand U21474 (N_21474,N_21182,N_21096);
and U21475 (N_21475,N_21129,N_21109);
nor U21476 (N_21476,N_21255,N_21169);
or U21477 (N_21477,N_21104,N_21166);
nand U21478 (N_21478,N_21006,N_21069);
and U21479 (N_21479,N_21113,N_21168);
xor U21480 (N_21480,N_21103,N_21141);
nand U21481 (N_21481,N_21047,N_21112);
or U21482 (N_21482,N_21127,N_21086);
nand U21483 (N_21483,N_21063,N_21263);
xnor U21484 (N_21484,N_21211,N_21073);
nand U21485 (N_21485,N_21181,N_21147);
xnor U21486 (N_21486,N_21283,N_21117);
nor U21487 (N_21487,N_21271,N_21134);
nor U21488 (N_21488,N_21148,N_21213);
xor U21489 (N_21489,N_21109,N_21050);
xnor U21490 (N_21490,N_21266,N_21270);
xor U21491 (N_21491,N_21181,N_21261);
or U21492 (N_21492,N_21066,N_21235);
nand U21493 (N_21493,N_21053,N_21064);
nor U21494 (N_21494,N_21202,N_21266);
or U21495 (N_21495,N_21247,N_21069);
and U21496 (N_21496,N_21175,N_21289);
nand U21497 (N_21497,N_21111,N_21122);
nand U21498 (N_21498,N_21102,N_21103);
xor U21499 (N_21499,N_21176,N_21225);
and U21500 (N_21500,N_21064,N_21245);
and U21501 (N_21501,N_21168,N_21086);
xor U21502 (N_21502,N_21028,N_21161);
and U21503 (N_21503,N_21246,N_21131);
or U21504 (N_21504,N_21254,N_21143);
and U21505 (N_21505,N_21055,N_21192);
or U21506 (N_21506,N_21096,N_21174);
and U21507 (N_21507,N_21222,N_21146);
xnor U21508 (N_21508,N_21176,N_21295);
xor U21509 (N_21509,N_21158,N_21135);
nand U21510 (N_21510,N_21066,N_21216);
nand U21511 (N_21511,N_21116,N_21006);
xnor U21512 (N_21512,N_21215,N_21107);
xor U21513 (N_21513,N_21212,N_21024);
xor U21514 (N_21514,N_21049,N_21123);
or U21515 (N_21515,N_21007,N_21250);
and U21516 (N_21516,N_21095,N_21253);
and U21517 (N_21517,N_21271,N_21006);
nand U21518 (N_21518,N_21176,N_21006);
xor U21519 (N_21519,N_21090,N_21160);
xnor U21520 (N_21520,N_21224,N_21275);
xor U21521 (N_21521,N_21241,N_21261);
or U21522 (N_21522,N_21112,N_21227);
nor U21523 (N_21523,N_21259,N_21142);
nand U21524 (N_21524,N_21019,N_21146);
nor U21525 (N_21525,N_21143,N_21127);
and U21526 (N_21526,N_21149,N_21178);
nor U21527 (N_21527,N_21059,N_21095);
and U21528 (N_21528,N_21216,N_21110);
xor U21529 (N_21529,N_21168,N_21026);
and U21530 (N_21530,N_21205,N_21299);
xnor U21531 (N_21531,N_21051,N_21060);
nand U21532 (N_21532,N_21114,N_21057);
nand U21533 (N_21533,N_21226,N_21017);
or U21534 (N_21534,N_21273,N_21264);
or U21535 (N_21535,N_21184,N_21121);
nor U21536 (N_21536,N_21198,N_21219);
nand U21537 (N_21537,N_21237,N_21238);
xor U21538 (N_21538,N_21230,N_21023);
nor U21539 (N_21539,N_21177,N_21131);
nand U21540 (N_21540,N_21222,N_21135);
or U21541 (N_21541,N_21026,N_21255);
xor U21542 (N_21542,N_21073,N_21285);
nor U21543 (N_21543,N_21062,N_21034);
nand U21544 (N_21544,N_21252,N_21118);
and U21545 (N_21545,N_21025,N_21069);
xor U21546 (N_21546,N_21030,N_21096);
nor U21547 (N_21547,N_21299,N_21170);
nor U21548 (N_21548,N_21140,N_21166);
nand U21549 (N_21549,N_21291,N_21175);
nor U21550 (N_21550,N_21039,N_21140);
or U21551 (N_21551,N_21132,N_21136);
nor U21552 (N_21552,N_21048,N_21165);
and U21553 (N_21553,N_21006,N_21220);
or U21554 (N_21554,N_21076,N_21091);
nand U21555 (N_21555,N_21074,N_21089);
and U21556 (N_21556,N_21024,N_21120);
or U21557 (N_21557,N_21126,N_21136);
xor U21558 (N_21558,N_21162,N_21000);
nor U21559 (N_21559,N_21147,N_21220);
or U21560 (N_21560,N_21198,N_21006);
and U21561 (N_21561,N_21200,N_21239);
and U21562 (N_21562,N_21149,N_21228);
nor U21563 (N_21563,N_21134,N_21290);
nand U21564 (N_21564,N_21212,N_21072);
xor U21565 (N_21565,N_21255,N_21204);
and U21566 (N_21566,N_21216,N_21012);
nor U21567 (N_21567,N_21261,N_21010);
nor U21568 (N_21568,N_21016,N_21024);
and U21569 (N_21569,N_21147,N_21001);
and U21570 (N_21570,N_21294,N_21141);
nor U21571 (N_21571,N_21200,N_21026);
and U21572 (N_21572,N_21003,N_21295);
or U21573 (N_21573,N_21142,N_21007);
and U21574 (N_21574,N_21234,N_21005);
or U21575 (N_21575,N_21132,N_21281);
and U21576 (N_21576,N_21025,N_21257);
xnor U21577 (N_21577,N_21085,N_21098);
and U21578 (N_21578,N_21136,N_21049);
nand U21579 (N_21579,N_21202,N_21126);
nand U21580 (N_21580,N_21197,N_21064);
and U21581 (N_21581,N_21055,N_21177);
nor U21582 (N_21582,N_21253,N_21272);
nand U21583 (N_21583,N_21053,N_21272);
nand U21584 (N_21584,N_21167,N_21295);
and U21585 (N_21585,N_21298,N_21282);
or U21586 (N_21586,N_21046,N_21201);
xnor U21587 (N_21587,N_21130,N_21276);
xnor U21588 (N_21588,N_21012,N_21264);
nor U21589 (N_21589,N_21055,N_21045);
or U21590 (N_21590,N_21277,N_21091);
or U21591 (N_21591,N_21099,N_21082);
xor U21592 (N_21592,N_21198,N_21189);
nand U21593 (N_21593,N_21209,N_21230);
xnor U21594 (N_21594,N_21295,N_21163);
nor U21595 (N_21595,N_21116,N_21039);
xnor U21596 (N_21596,N_21299,N_21186);
or U21597 (N_21597,N_21078,N_21185);
nand U21598 (N_21598,N_21172,N_21280);
or U21599 (N_21599,N_21139,N_21121);
nand U21600 (N_21600,N_21554,N_21544);
or U21601 (N_21601,N_21514,N_21459);
nor U21602 (N_21602,N_21522,N_21548);
or U21603 (N_21603,N_21582,N_21537);
or U21604 (N_21604,N_21507,N_21335);
and U21605 (N_21605,N_21431,N_21306);
nor U21606 (N_21606,N_21447,N_21468);
nor U21607 (N_21607,N_21323,N_21474);
nand U21608 (N_21608,N_21588,N_21477);
nand U21609 (N_21609,N_21325,N_21592);
nand U21610 (N_21610,N_21317,N_21495);
nor U21611 (N_21611,N_21476,N_21432);
and U21612 (N_21612,N_21412,N_21585);
or U21613 (N_21613,N_21384,N_21307);
nor U21614 (N_21614,N_21524,N_21430);
nand U21615 (N_21615,N_21442,N_21342);
nor U21616 (N_21616,N_21419,N_21408);
nand U21617 (N_21617,N_21300,N_21454);
nand U21618 (N_21618,N_21395,N_21471);
xor U21619 (N_21619,N_21556,N_21318);
and U21620 (N_21620,N_21547,N_21532);
and U21621 (N_21621,N_21399,N_21493);
or U21622 (N_21622,N_21349,N_21390);
nand U21623 (N_21623,N_21566,N_21309);
nand U21624 (N_21624,N_21561,N_21340);
nor U21625 (N_21625,N_21387,N_21483);
nor U21626 (N_21626,N_21543,N_21310);
xnor U21627 (N_21627,N_21385,N_21417);
or U21628 (N_21628,N_21329,N_21456);
or U21629 (N_21629,N_21478,N_21389);
and U21630 (N_21630,N_21303,N_21527);
or U21631 (N_21631,N_21565,N_21348);
or U21632 (N_21632,N_21350,N_21392);
and U21633 (N_21633,N_21552,N_21518);
or U21634 (N_21634,N_21433,N_21455);
or U21635 (N_21635,N_21555,N_21376);
nand U21636 (N_21636,N_21511,N_21510);
nand U21637 (N_21637,N_21405,N_21579);
xor U21638 (N_21638,N_21311,N_21458);
xor U21639 (N_21639,N_21439,N_21469);
or U21640 (N_21640,N_21595,N_21407);
or U21641 (N_21641,N_21370,N_21573);
or U21642 (N_21642,N_21328,N_21429);
nand U21643 (N_21643,N_21400,N_21330);
xnor U21644 (N_21644,N_21396,N_21457);
or U21645 (N_21645,N_21393,N_21418);
or U21646 (N_21646,N_21529,N_21533);
nor U21647 (N_21647,N_21558,N_21485);
xor U21648 (N_21648,N_21539,N_21578);
or U21649 (N_21649,N_21386,N_21319);
nor U21650 (N_21650,N_21308,N_21502);
nand U21651 (N_21651,N_21375,N_21540);
nor U21652 (N_21652,N_21353,N_21314);
and U21653 (N_21653,N_21491,N_21321);
or U21654 (N_21654,N_21327,N_21336);
nor U21655 (N_21655,N_21538,N_21568);
and U21656 (N_21656,N_21461,N_21591);
nor U21657 (N_21657,N_21362,N_21427);
nand U21658 (N_21658,N_21453,N_21531);
and U21659 (N_21659,N_21535,N_21480);
or U21660 (N_21660,N_21356,N_21346);
and U21661 (N_21661,N_21519,N_21574);
or U21662 (N_21662,N_21363,N_21504);
and U21663 (N_21663,N_21545,N_21445);
xnor U21664 (N_21664,N_21435,N_21572);
nor U21665 (N_21665,N_21551,N_21377);
xnor U21666 (N_21666,N_21489,N_21517);
or U21667 (N_21667,N_21557,N_21438);
nor U21668 (N_21668,N_21422,N_21313);
and U21669 (N_21669,N_21357,N_21406);
xnor U21670 (N_21670,N_21496,N_21379);
xnor U21671 (N_21671,N_21351,N_21304);
xnor U21672 (N_21672,N_21508,N_21589);
nand U21673 (N_21673,N_21382,N_21497);
xor U21674 (N_21674,N_21449,N_21580);
and U21675 (N_21675,N_21597,N_21562);
nor U21676 (N_21676,N_21423,N_21549);
xor U21677 (N_21677,N_21426,N_21398);
and U21678 (N_21678,N_21437,N_21440);
nand U21679 (N_21679,N_21479,N_21443);
or U21680 (N_21680,N_21486,N_21421);
and U21681 (N_21681,N_21420,N_21584);
xnor U21682 (N_21682,N_21409,N_21371);
nor U21683 (N_21683,N_21467,N_21364);
nand U21684 (N_21684,N_21465,N_21506);
nor U21685 (N_21685,N_21301,N_21345);
nor U21686 (N_21686,N_21475,N_21521);
nor U21687 (N_21687,N_21594,N_21470);
and U21688 (N_21688,N_21305,N_21494);
nand U21689 (N_21689,N_21450,N_21596);
or U21690 (N_21690,N_21586,N_21359);
or U21691 (N_21691,N_21500,N_21394);
xnor U21692 (N_21692,N_21541,N_21397);
and U21693 (N_21693,N_21593,N_21341);
or U21694 (N_21694,N_21373,N_21368);
nand U21695 (N_21695,N_21516,N_21515);
or U21696 (N_21696,N_21320,N_21571);
nor U21697 (N_21697,N_21583,N_21372);
or U21698 (N_21698,N_21490,N_21367);
xnor U21699 (N_21699,N_21365,N_21331);
nand U21700 (N_21700,N_21425,N_21481);
or U21701 (N_21701,N_21347,N_21404);
and U21702 (N_21702,N_21416,N_21316);
or U21703 (N_21703,N_21463,N_21599);
xnor U21704 (N_21704,N_21570,N_21513);
and U21705 (N_21705,N_21472,N_21360);
xor U21706 (N_21706,N_21464,N_21403);
or U21707 (N_21707,N_21520,N_21302);
nor U21708 (N_21708,N_21546,N_21492);
or U21709 (N_21709,N_21523,N_21473);
or U21710 (N_21710,N_21460,N_21381);
and U21711 (N_21711,N_21452,N_21569);
and U21712 (N_21712,N_21576,N_21354);
xor U21713 (N_21713,N_21448,N_21441);
nand U21714 (N_21714,N_21512,N_21388);
nand U21715 (N_21715,N_21499,N_21401);
xnor U21716 (N_21716,N_21509,N_21322);
xnor U21717 (N_21717,N_21414,N_21451);
xor U21718 (N_21718,N_21369,N_21366);
and U21719 (N_21719,N_21587,N_21488);
and U21720 (N_21720,N_21567,N_21324);
xnor U21721 (N_21721,N_21575,N_21530);
nand U21722 (N_21722,N_21487,N_21410);
and U21723 (N_21723,N_21374,N_21553);
or U21724 (N_21724,N_21528,N_21332);
nor U21725 (N_21725,N_21315,N_21436);
xnor U21726 (N_21726,N_21355,N_21581);
and U21727 (N_21727,N_21484,N_21337);
and U21728 (N_21728,N_21590,N_21413);
nor U21729 (N_21729,N_21501,N_21526);
nor U21730 (N_21730,N_21334,N_21505);
nand U21731 (N_21731,N_21434,N_21358);
and U21732 (N_21732,N_21391,N_21444);
xnor U21733 (N_21733,N_21577,N_21339);
and U21734 (N_21734,N_21498,N_21482);
xor U21735 (N_21735,N_21312,N_21383);
nor U21736 (N_21736,N_21338,N_21415);
nand U21737 (N_21737,N_21428,N_21361);
nor U21738 (N_21738,N_21559,N_21563);
xnor U21739 (N_21739,N_21550,N_21326);
xnor U21740 (N_21740,N_21564,N_21411);
and U21741 (N_21741,N_21378,N_21462);
and U21742 (N_21742,N_21333,N_21534);
nor U21743 (N_21743,N_21525,N_21343);
nand U21744 (N_21744,N_21560,N_21380);
or U21745 (N_21745,N_21466,N_21344);
and U21746 (N_21746,N_21446,N_21542);
nand U21747 (N_21747,N_21424,N_21402);
or U21748 (N_21748,N_21536,N_21598);
nand U21749 (N_21749,N_21352,N_21503);
xor U21750 (N_21750,N_21572,N_21396);
and U21751 (N_21751,N_21399,N_21396);
or U21752 (N_21752,N_21509,N_21347);
xnor U21753 (N_21753,N_21476,N_21438);
nor U21754 (N_21754,N_21506,N_21595);
nand U21755 (N_21755,N_21336,N_21325);
or U21756 (N_21756,N_21593,N_21442);
and U21757 (N_21757,N_21535,N_21356);
and U21758 (N_21758,N_21458,N_21484);
or U21759 (N_21759,N_21538,N_21363);
xnor U21760 (N_21760,N_21543,N_21394);
or U21761 (N_21761,N_21314,N_21316);
xor U21762 (N_21762,N_21397,N_21510);
nor U21763 (N_21763,N_21480,N_21572);
or U21764 (N_21764,N_21379,N_21543);
nor U21765 (N_21765,N_21446,N_21519);
nor U21766 (N_21766,N_21318,N_21471);
nand U21767 (N_21767,N_21405,N_21483);
nand U21768 (N_21768,N_21424,N_21422);
nor U21769 (N_21769,N_21460,N_21302);
nand U21770 (N_21770,N_21503,N_21312);
xnor U21771 (N_21771,N_21376,N_21465);
or U21772 (N_21772,N_21556,N_21451);
nand U21773 (N_21773,N_21560,N_21572);
xnor U21774 (N_21774,N_21571,N_21598);
and U21775 (N_21775,N_21510,N_21381);
and U21776 (N_21776,N_21348,N_21528);
nor U21777 (N_21777,N_21547,N_21589);
or U21778 (N_21778,N_21365,N_21426);
xor U21779 (N_21779,N_21370,N_21381);
nand U21780 (N_21780,N_21500,N_21573);
nand U21781 (N_21781,N_21494,N_21398);
and U21782 (N_21782,N_21384,N_21460);
xnor U21783 (N_21783,N_21586,N_21349);
xor U21784 (N_21784,N_21418,N_21324);
or U21785 (N_21785,N_21512,N_21410);
nor U21786 (N_21786,N_21556,N_21417);
nor U21787 (N_21787,N_21392,N_21414);
nor U21788 (N_21788,N_21555,N_21364);
xor U21789 (N_21789,N_21368,N_21354);
and U21790 (N_21790,N_21459,N_21482);
xor U21791 (N_21791,N_21438,N_21317);
nor U21792 (N_21792,N_21346,N_21427);
nor U21793 (N_21793,N_21394,N_21383);
nor U21794 (N_21794,N_21581,N_21548);
xnor U21795 (N_21795,N_21476,N_21389);
nor U21796 (N_21796,N_21322,N_21531);
xnor U21797 (N_21797,N_21319,N_21324);
xor U21798 (N_21798,N_21376,N_21455);
nand U21799 (N_21799,N_21553,N_21570);
xor U21800 (N_21800,N_21334,N_21585);
and U21801 (N_21801,N_21459,N_21369);
and U21802 (N_21802,N_21379,N_21310);
and U21803 (N_21803,N_21567,N_21424);
nor U21804 (N_21804,N_21469,N_21496);
xnor U21805 (N_21805,N_21497,N_21324);
and U21806 (N_21806,N_21551,N_21354);
nand U21807 (N_21807,N_21529,N_21462);
and U21808 (N_21808,N_21323,N_21427);
nor U21809 (N_21809,N_21302,N_21310);
nand U21810 (N_21810,N_21478,N_21308);
nand U21811 (N_21811,N_21440,N_21359);
and U21812 (N_21812,N_21450,N_21474);
and U21813 (N_21813,N_21474,N_21391);
and U21814 (N_21814,N_21479,N_21410);
xor U21815 (N_21815,N_21414,N_21535);
nor U21816 (N_21816,N_21472,N_21481);
xnor U21817 (N_21817,N_21329,N_21581);
xor U21818 (N_21818,N_21564,N_21469);
or U21819 (N_21819,N_21405,N_21446);
xnor U21820 (N_21820,N_21510,N_21484);
nand U21821 (N_21821,N_21408,N_21431);
nor U21822 (N_21822,N_21462,N_21568);
and U21823 (N_21823,N_21504,N_21539);
or U21824 (N_21824,N_21438,N_21571);
and U21825 (N_21825,N_21411,N_21433);
nand U21826 (N_21826,N_21521,N_21326);
nand U21827 (N_21827,N_21320,N_21452);
nor U21828 (N_21828,N_21500,N_21537);
or U21829 (N_21829,N_21494,N_21548);
nand U21830 (N_21830,N_21496,N_21425);
or U21831 (N_21831,N_21542,N_21511);
xor U21832 (N_21832,N_21598,N_21531);
nor U21833 (N_21833,N_21599,N_21532);
or U21834 (N_21834,N_21307,N_21548);
xor U21835 (N_21835,N_21581,N_21549);
nand U21836 (N_21836,N_21344,N_21567);
nor U21837 (N_21837,N_21436,N_21373);
xor U21838 (N_21838,N_21348,N_21452);
xnor U21839 (N_21839,N_21491,N_21536);
and U21840 (N_21840,N_21411,N_21418);
or U21841 (N_21841,N_21321,N_21303);
xor U21842 (N_21842,N_21566,N_21473);
or U21843 (N_21843,N_21581,N_21518);
nor U21844 (N_21844,N_21590,N_21544);
and U21845 (N_21845,N_21390,N_21388);
and U21846 (N_21846,N_21427,N_21438);
and U21847 (N_21847,N_21508,N_21435);
or U21848 (N_21848,N_21487,N_21400);
and U21849 (N_21849,N_21495,N_21470);
and U21850 (N_21850,N_21544,N_21579);
or U21851 (N_21851,N_21468,N_21366);
xor U21852 (N_21852,N_21598,N_21568);
and U21853 (N_21853,N_21322,N_21583);
and U21854 (N_21854,N_21467,N_21537);
xnor U21855 (N_21855,N_21368,N_21465);
nand U21856 (N_21856,N_21458,N_21410);
or U21857 (N_21857,N_21493,N_21488);
or U21858 (N_21858,N_21461,N_21379);
xnor U21859 (N_21859,N_21589,N_21393);
xor U21860 (N_21860,N_21573,N_21319);
nor U21861 (N_21861,N_21377,N_21533);
and U21862 (N_21862,N_21395,N_21428);
nand U21863 (N_21863,N_21571,N_21398);
or U21864 (N_21864,N_21494,N_21556);
nor U21865 (N_21865,N_21461,N_21467);
and U21866 (N_21866,N_21535,N_21347);
nand U21867 (N_21867,N_21459,N_21351);
or U21868 (N_21868,N_21507,N_21535);
and U21869 (N_21869,N_21518,N_21565);
xor U21870 (N_21870,N_21313,N_21490);
nand U21871 (N_21871,N_21566,N_21347);
and U21872 (N_21872,N_21327,N_21437);
xnor U21873 (N_21873,N_21465,N_21585);
nand U21874 (N_21874,N_21311,N_21420);
nor U21875 (N_21875,N_21359,N_21544);
xnor U21876 (N_21876,N_21419,N_21411);
xor U21877 (N_21877,N_21583,N_21566);
and U21878 (N_21878,N_21353,N_21330);
nor U21879 (N_21879,N_21315,N_21362);
and U21880 (N_21880,N_21516,N_21372);
nor U21881 (N_21881,N_21545,N_21500);
nand U21882 (N_21882,N_21443,N_21346);
or U21883 (N_21883,N_21426,N_21409);
nand U21884 (N_21884,N_21417,N_21390);
nor U21885 (N_21885,N_21478,N_21589);
or U21886 (N_21886,N_21569,N_21300);
nor U21887 (N_21887,N_21542,N_21419);
and U21888 (N_21888,N_21520,N_21560);
nor U21889 (N_21889,N_21591,N_21431);
or U21890 (N_21890,N_21320,N_21433);
or U21891 (N_21891,N_21455,N_21425);
or U21892 (N_21892,N_21326,N_21463);
nor U21893 (N_21893,N_21399,N_21358);
xnor U21894 (N_21894,N_21431,N_21378);
and U21895 (N_21895,N_21394,N_21421);
nor U21896 (N_21896,N_21556,N_21335);
or U21897 (N_21897,N_21352,N_21499);
nand U21898 (N_21898,N_21486,N_21303);
nor U21899 (N_21899,N_21585,N_21318);
or U21900 (N_21900,N_21656,N_21696);
and U21901 (N_21901,N_21894,N_21637);
nor U21902 (N_21902,N_21748,N_21796);
nand U21903 (N_21903,N_21784,N_21850);
and U21904 (N_21904,N_21604,N_21650);
or U21905 (N_21905,N_21742,N_21855);
nand U21906 (N_21906,N_21833,N_21835);
xor U21907 (N_21907,N_21633,N_21773);
and U21908 (N_21908,N_21752,N_21876);
and U21909 (N_21909,N_21660,N_21783);
and U21910 (N_21910,N_21781,N_21654);
nand U21911 (N_21911,N_21628,N_21821);
xor U21912 (N_21912,N_21763,N_21780);
nand U21913 (N_21913,N_21775,N_21615);
or U21914 (N_21914,N_21738,N_21778);
xnor U21915 (N_21915,N_21756,N_21725);
nor U21916 (N_21916,N_21834,N_21768);
and U21917 (N_21917,N_21639,N_21795);
nor U21918 (N_21918,N_21886,N_21652);
xor U21919 (N_21919,N_21716,N_21769);
xor U21920 (N_21920,N_21772,N_21644);
and U21921 (N_21921,N_21642,N_21811);
or U21922 (N_21922,N_21718,N_21865);
or U21923 (N_21923,N_21840,N_21706);
nor U21924 (N_21924,N_21852,N_21793);
or U21925 (N_21925,N_21826,N_21856);
and U21926 (N_21926,N_21627,N_21875);
nor U21927 (N_21927,N_21661,N_21609);
or U21928 (N_21928,N_21662,N_21740);
nor U21929 (N_21929,N_21729,N_21683);
nand U21930 (N_21930,N_21694,N_21761);
xnor U21931 (N_21931,N_21798,N_21843);
or U21932 (N_21932,N_21680,N_21638);
xor U21933 (N_21933,N_21805,N_21734);
and U21934 (N_21934,N_21816,N_21676);
nand U21935 (N_21935,N_21817,N_21787);
or U21936 (N_21936,N_21732,N_21704);
or U21937 (N_21937,N_21657,N_21606);
xor U21938 (N_21938,N_21744,N_21836);
or U21939 (N_21939,N_21668,N_21622);
nand U21940 (N_21940,N_21818,N_21803);
and U21941 (N_21941,N_21667,N_21617);
nor U21942 (N_21942,N_21646,N_21714);
xnor U21943 (N_21943,N_21736,N_21831);
xor U21944 (N_21944,N_21789,N_21653);
nor U21945 (N_21945,N_21669,N_21874);
and U21946 (N_21946,N_21708,N_21681);
and U21947 (N_21947,N_21621,N_21619);
xor U21948 (N_21948,N_21624,N_21685);
nor U21949 (N_21949,N_21695,N_21705);
and U21950 (N_21950,N_21765,N_21655);
or U21951 (N_21951,N_21790,N_21877);
nand U21952 (N_21952,N_21895,N_21693);
and U21953 (N_21953,N_21869,N_21632);
nor U21954 (N_21954,N_21883,N_21777);
nand U21955 (N_21955,N_21814,N_21794);
nand U21956 (N_21956,N_21849,N_21829);
or U21957 (N_21957,N_21675,N_21717);
xnor U21958 (N_21958,N_21827,N_21864);
nor U21959 (N_21959,N_21888,N_21866);
or U21960 (N_21960,N_21641,N_21601);
and U21961 (N_21961,N_21824,N_21616);
or U21962 (N_21962,N_21688,N_21678);
nand U21963 (N_21963,N_21643,N_21801);
xnor U21964 (N_21964,N_21698,N_21721);
nor U21965 (N_21965,N_21853,N_21719);
nand U21966 (N_21966,N_21699,N_21697);
or U21967 (N_21967,N_21726,N_21844);
xor U21968 (N_21968,N_21722,N_21700);
and U21969 (N_21969,N_21792,N_21707);
and U21970 (N_21970,N_21647,N_21770);
and U21971 (N_21971,N_21860,N_21879);
or U21972 (N_21972,N_21749,N_21898);
nor U21973 (N_21973,N_21602,N_21762);
xnor U21974 (N_21974,N_21750,N_21851);
nand U21975 (N_21975,N_21753,N_21614);
nor U21976 (N_21976,N_21679,N_21723);
or U21977 (N_21977,N_21603,N_21782);
nand U21978 (N_21978,N_21797,N_21873);
nor U21979 (N_21979,N_21806,N_21820);
nor U21980 (N_21980,N_21737,N_21684);
xnor U21981 (N_21981,N_21871,N_21702);
and U21982 (N_21982,N_21823,N_21649);
and U21983 (N_21983,N_21691,N_21677);
or U21984 (N_21984,N_21881,N_21857);
and U21985 (N_21985,N_21659,N_21880);
xor U21986 (N_21986,N_21832,N_21727);
xor U21987 (N_21987,N_21760,N_21893);
and U21988 (N_21988,N_21735,N_21837);
or U21989 (N_21989,N_21776,N_21728);
xor U21990 (N_21990,N_21636,N_21730);
and U21991 (N_21991,N_21897,N_21613);
nand U21992 (N_21992,N_21799,N_21870);
or U21993 (N_21993,N_21672,N_21743);
xor U21994 (N_21994,N_21774,N_21758);
and U21995 (N_21995,N_21611,N_21885);
xnor U21996 (N_21996,N_21810,N_21623);
or U21997 (N_21997,N_21846,N_21896);
nand U21998 (N_21998,N_21626,N_21682);
nor U21999 (N_21999,N_21755,N_21884);
nor U22000 (N_22000,N_21890,N_21607);
xor U22001 (N_22001,N_21779,N_21634);
xnor U22002 (N_22002,N_21629,N_21800);
xnor U22003 (N_22003,N_21701,N_21709);
xor U22004 (N_22004,N_21712,N_21862);
xor U22005 (N_22005,N_21664,N_21686);
nand U22006 (N_22006,N_21731,N_21631);
xnor U22007 (N_22007,N_21670,N_21635);
or U22008 (N_22008,N_21747,N_21625);
xnor U22009 (N_22009,N_21618,N_21600);
nand U22010 (N_22010,N_21889,N_21665);
xnor U22011 (N_22011,N_21812,N_21751);
or U22012 (N_22012,N_21809,N_21651);
nor U22013 (N_22013,N_21839,N_21802);
nor U22014 (N_22014,N_21845,N_21741);
xor U22015 (N_22015,N_21746,N_21733);
nor U22016 (N_22016,N_21620,N_21767);
nand U22017 (N_22017,N_21674,N_21892);
or U22018 (N_22018,N_21658,N_21819);
and U22019 (N_22019,N_21703,N_21858);
and U22020 (N_22020,N_21608,N_21757);
or U22021 (N_22021,N_21724,N_21745);
or U22022 (N_22022,N_21671,N_21891);
or U22023 (N_22023,N_21822,N_21715);
and U22024 (N_22024,N_21610,N_21785);
nand U22025 (N_22025,N_21807,N_21791);
xor U22026 (N_22026,N_21766,N_21838);
nor U22027 (N_22027,N_21663,N_21689);
or U22028 (N_22028,N_21804,N_21648);
xnor U22029 (N_22029,N_21815,N_21605);
xnor U22030 (N_22030,N_21666,N_21687);
xnor U22031 (N_22031,N_21720,N_21630);
nor U22032 (N_22032,N_21711,N_21788);
and U22033 (N_22033,N_21771,N_21878);
nor U22034 (N_22034,N_21612,N_21673);
nand U22035 (N_22035,N_21813,N_21830);
xor U22036 (N_22036,N_21713,N_21841);
nor U22037 (N_22037,N_21640,N_21882);
xnor U22038 (N_22038,N_21868,N_21692);
and U22039 (N_22039,N_21825,N_21887);
xor U22040 (N_22040,N_21872,N_21786);
xor U22041 (N_22041,N_21645,N_21690);
or U22042 (N_22042,N_21828,N_21764);
xor U22043 (N_22043,N_21710,N_21848);
nor U22044 (N_22044,N_21854,N_21859);
and U22045 (N_22045,N_21739,N_21754);
or U22046 (N_22046,N_21863,N_21899);
nand U22047 (N_22047,N_21759,N_21808);
xnor U22048 (N_22048,N_21842,N_21847);
or U22049 (N_22049,N_21867,N_21861);
xor U22050 (N_22050,N_21680,N_21633);
and U22051 (N_22051,N_21657,N_21811);
xor U22052 (N_22052,N_21790,N_21727);
xor U22053 (N_22053,N_21771,N_21844);
and U22054 (N_22054,N_21714,N_21842);
or U22055 (N_22055,N_21742,N_21646);
or U22056 (N_22056,N_21862,N_21819);
and U22057 (N_22057,N_21698,N_21810);
or U22058 (N_22058,N_21732,N_21702);
xor U22059 (N_22059,N_21769,N_21863);
or U22060 (N_22060,N_21845,N_21816);
and U22061 (N_22061,N_21686,N_21681);
nand U22062 (N_22062,N_21685,N_21808);
and U22063 (N_22063,N_21732,N_21640);
nand U22064 (N_22064,N_21824,N_21621);
nand U22065 (N_22065,N_21733,N_21763);
or U22066 (N_22066,N_21772,N_21656);
and U22067 (N_22067,N_21705,N_21742);
nand U22068 (N_22068,N_21716,N_21643);
and U22069 (N_22069,N_21787,N_21767);
nor U22070 (N_22070,N_21711,N_21755);
xor U22071 (N_22071,N_21682,N_21820);
and U22072 (N_22072,N_21604,N_21624);
nor U22073 (N_22073,N_21673,N_21625);
nor U22074 (N_22074,N_21775,N_21837);
or U22075 (N_22075,N_21673,N_21834);
xnor U22076 (N_22076,N_21881,N_21823);
and U22077 (N_22077,N_21674,N_21607);
nor U22078 (N_22078,N_21790,N_21859);
nand U22079 (N_22079,N_21767,N_21881);
and U22080 (N_22080,N_21701,N_21645);
and U22081 (N_22081,N_21634,N_21601);
or U22082 (N_22082,N_21655,N_21822);
or U22083 (N_22083,N_21714,N_21783);
nor U22084 (N_22084,N_21677,N_21636);
nor U22085 (N_22085,N_21828,N_21833);
and U22086 (N_22086,N_21735,N_21602);
xor U22087 (N_22087,N_21693,N_21867);
xor U22088 (N_22088,N_21802,N_21757);
nand U22089 (N_22089,N_21725,N_21846);
nand U22090 (N_22090,N_21693,N_21847);
and U22091 (N_22091,N_21743,N_21742);
nor U22092 (N_22092,N_21836,N_21615);
nor U22093 (N_22093,N_21662,N_21681);
or U22094 (N_22094,N_21738,N_21874);
nor U22095 (N_22095,N_21879,N_21883);
and U22096 (N_22096,N_21795,N_21783);
nor U22097 (N_22097,N_21830,N_21705);
nor U22098 (N_22098,N_21726,N_21645);
nor U22099 (N_22099,N_21625,N_21670);
or U22100 (N_22100,N_21699,N_21634);
and U22101 (N_22101,N_21810,N_21691);
and U22102 (N_22102,N_21754,N_21729);
xnor U22103 (N_22103,N_21667,N_21643);
nand U22104 (N_22104,N_21879,N_21880);
and U22105 (N_22105,N_21801,N_21719);
xor U22106 (N_22106,N_21835,N_21825);
and U22107 (N_22107,N_21882,N_21616);
or U22108 (N_22108,N_21878,N_21813);
or U22109 (N_22109,N_21601,N_21646);
nor U22110 (N_22110,N_21703,N_21805);
nor U22111 (N_22111,N_21605,N_21868);
nor U22112 (N_22112,N_21811,N_21660);
and U22113 (N_22113,N_21614,N_21745);
nor U22114 (N_22114,N_21618,N_21655);
and U22115 (N_22115,N_21649,N_21623);
and U22116 (N_22116,N_21751,N_21629);
nand U22117 (N_22117,N_21883,N_21607);
or U22118 (N_22118,N_21831,N_21795);
xnor U22119 (N_22119,N_21831,N_21698);
or U22120 (N_22120,N_21659,N_21621);
and U22121 (N_22121,N_21683,N_21815);
xor U22122 (N_22122,N_21811,N_21607);
and U22123 (N_22123,N_21639,N_21804);
nor U22124 (N_22124,N_21843,N_21861);
nand U22125 (N_22125,N_21764,N_21811);
or U22126 (N_22126,N_21766,N_21687);
xnor U22127 (N_22127,N_21899,N_21859);
or U22128 (N_22128,N_21891,N_21604);
nand U22129 (N_22129,N_21858,N_21691);
or U22130 (N_22130,N_21704,N_21686);
nand U22131 (N_22131,N_21732,N_21711);
xor U22132 (N_22132,N_21616,N_21800);
and U22133 (N_22133,N_21772,N_21894);
nor U22134 (N_22134,N_21836,N_21729);
xor U22135 (N_22135,N_21702,N_21685);
nand U22136 (N_22136,N_21758,N_21721);
xor U22137 (N_22137,N_21777,N_21668);
or U22138 (N_22138,N_21760,N_21731);
xnor U22139 (N_22139,N_21801,N_21871);
xnor U22140 (N_22140,N_21631,N_21753);
nand U22141 (N_22141,N_21679,N_21712);
nor U22142 (N_22142,N_21609,N_21765);
xnor U22143 (N_22143,N_21817,N_21685);
nor U22144 (N_22144,N_21889,N_21856);
and U22145 (N_22145,N_21706,N_21861);
xnor U22146 (N_22146,N_21826,N_21879);
xnor U22147 (N_22147,N_21852,N_21652);
nand U22148 (N_22148,N_21650,N_21715);
nand U22149 (N_22149,N_21699,N_21720);
or U22150 (N_22150,N_21898,N_21667);
nand U22151 (N_22151,N_21756,N_21613);
nand U22152 (N_22152,N_21616,N_21776);
nor U22153 (N_22153,N_21844,N_21884);
or U22154 (N_22154,N_21899,N_21687);
nand U22155 (N_22155,N_21854,N_21841);
nor U22156 (N_22156,N_21676,N_21863);
xor U22157 (N_22157,N_21679,N_21672);
xor U22158 (N_22158,N_21803,N_21767);
xor U22159 (N_22159,N_21822,N_21737);
xnor U22160 (N_22160,N_21705,N_21680);
or U22161 (N_22161,N_21811,N_21785);
and U22162 (N_22162,N_21683,N_21862);
or U22163 (N_22163,N_21691,N_21655);
and U22164 (N_22164,N_21606,N_21760);
nand U22165 (N_22165,N_21775,N_21751);
or U22166 (N_22166,N_21817,N_21613);
or U22167 (N_22167,N_21799,N_21605);
or U22168 (N_22168,N_21858,N_21646);
nand U22169 (N_22169,N_21708,N_21677);
nor U22170 (N_22170,N_21709,N_21840);
nand U22171 (N_22171,N_21773,N_21719);
or U22172 (N_22172,N_21717,N_21788);
xor U22173 (N_22173,N_21818,N_21611);
and U22174 (N_22174,N_21822,N_21859);
or U22175 (N_22175,N_21788,N_21780);
and U22176 (N_22176,N_21732,N_21804);
xnor U22177 (N_22177,N_21808,N_21749);
xnor U22178 (N_22178,N_21710,N_21871);
nor U22179 (N_22179,N_21729,N_21840);
or U22180 (N_22180,N_21631,N_21699);
and U22181 (N_22181,N_21745,N_21898);
nor U22182 (N_22182,N_21630,N_21761);
nor U22183 (N_22183,N_21612,N_21876);
or U22184 (N_22184,N_21650,N_21646);
nor U22185 (N_22185,N_21715,N_21630);
nor U22186 (N_22186,N_21676,N_21795);
xnor U22187 (N_22187,N_21846,N_21705);
or U22188 (N_22188,N_21758,N_21695);
nor U22189 (N_22189,N_21848,N_21754);
xnor U22190 (N_22190,N_21862,N_21836);
nor U22191 (N_22191,N_21690,N_21822);
or U22192 (N_22192,N_21887,N_21620);
and U22193 (N_22193,N_21610,N_21671);
nand U22194 (N_22194,N_21652,N_21759);
nand U22195 (N_22195,N_21855,N_21845);
nor U22196 (N_22196,N_21783,N_21621);
xnor U22197 (N_22197,N_21885,N_21871);
xnor U22198 (N_22198,N_21714,N_21889);
and U22199 (N_22199,N_21814,N_21629);
and U22200 (N_22200,N_22177,N_21933);
nor U22201 (N_22201,N_22173,N_22061);
nand U22202 (N_22202,N_21907,N_21915);
xnor U22203 (N_22203,N_22165,N_22190);
or U22204 (N_22204,N_22099,N_21997);
nor U22205 (N_22205,N_22192,N_22068);
or U22206 (N_22206,N_22182,N_21917);
nand U22207 (N_22207,N_22101,N_22112);
or U22208 (N_22208,N_22123,N_22087);
nand U22209 (N_22209,N_22086,N_22089);
nand U22210 (N_22210,N_22075,N_22138);
or U22211 (N_22211,N_21920,N_22062);
nor U22212 (N_22212,N_22161,N_21991);
and U22213 (N_22213,N_22030,N_22103);
and U22214 (N_22214,N_21996,N_22104);
nor U22215 (N_22215,N_22047,N_22186);
nand U22216 (N_22216,N_22094,N_22096);
nor U22217 (N_22217,N_21938,N_22126);
nor U22218 (N_22218,N_22070,N_22083);
nor U22219 (N_22219,N_22105,N_22010);
or U22220 (N_22220,N_21926,N_22155);
xnor U22221 (N_22221,N_21990,N_22129);
and U22222 (N_22222,N_22137,N_22116);
nor U22223 (N_22223,N_22156,N_22102);
xnor U22224 (N_22224,N_21992,N_22072);
and U22225 (N_22225,N_22012,N_22019);
nor U22226 (N_22226,N_22179,N_22121);
nor U22227 (N_22227,N_22097,N_22014);
xor U22228 (N_22228,N_22154,N_22198);
or U22229 (N_22229,N_21930,N_22084);
and U22230 (N_22230,N_22039,N_21982);
nor U22231 (N_22231,N_22051,N_21989);
nor U22232 (N_22232,N_22018,N_22088);
nand U22233 (N_22233,N_22191,N_22195);
or U22234 (N_22234,N_22033,N_22076);
nand U22235 (N_22235,N_22036,N_21931);
nand U22236 (N_22236,N_22187,N_22042);
nand U22237 (N_22237,N_22170,N_22034);
and U22238 (N_22238,N_22189,N_22145);
or U22239 (N_22239,N_21932,N_21948);
and U22240 (N_22240,N_21949,N_21909);
xnor U22241 (N_22241,N_21954,N_21994);
nor U22242 (N_22242,N_22193,N_22082);
nor U22243 (N_22243,N_22168,N_22074);
or U22244 (N_22244,N_22060,N_22149);
nor U22245 (N_22245,N_21985,N_21934);
and U22246 (N_22246,N_21939,N_21906);
nor U22247 (N_22247,N_22150,N_22120);
nand U22248 (N_22248,N_22091,N_22058);
or U22249 (N_22249,N_22045,N_21945);
or U22250 (N_22250,N_21927,N_22079);
nor U22251 (N_22251,N_21973,N_22148);
nand U22252 (N_22252,N_22199,N_22057);
nand U22253 (N_22253,N_22122,N_21903);
and U22254 (N_22254,N_22171,N_22055);
xnor U22255 (N_22255,N_22181,N_22001);
nand U22256 (N_22256,N_22040,N_21957);
nand U22257 (N_22257,N_22002,N_22000);
and U22258 (N_22258,N_22024,N_21911);
xnor U22259 (N_22259,N_22081,N_22100);
and U22260 (N_22260,N_22174,N_21967);
and U22261 (N_22261,N_22038,N_21904);
nor U22262 (N_22262,N_21935,N_21966);
and U22263 (N_22263,N_22052,N_22020);
and U22264 (N_22264,N_21964,N_22163);
nand U22265 (N_22265,N_22064,N_21944);
or U22266 (N_22266,N_21942,N_21960);
xnor U22267 (N_22267,N_22118,N_22041);
xor U22268 (N_22268,N_22111,N_21914);
xnor U22269 (N_22269,N_21961,N_22085);
xnor U22270 (N_22270,N_21999,N_21955);
nor U22271 (N_22271,N_22028,N_21986);
or U22272 (N_22272,N_22140,N_21972);
nor U22273 (N_22273,N_22007,N_21987);
or U22274 (N_22274,N_22167,N_22152);
xnor U22275 (N_22275,N_22043,N_22166);
nor U22276 (N_22276,N_22108,N_22054);
or U22277 (N_22277,N_22106,N_21953);
nand U22278 (N_22278,N_22185,N_22157);
or U22279 (N_22279,N_22063,N_22127);
nor U22280 (N_22280,N_22027,N_22109);
or U22281 (N_22281,N_22169,N_21941);
nand U22282 (N_22282,N_22056,N_21965);
xnor U22283 (N_22283,N_22130,N_22004);
xnor U22284 (N_22284,N_22180,N_22069);
nor U22285 (N_22285,N_22066,N_22141);
or U22286 (N_22286,N_21902,N_22005);
nor U22287 (N_22287,N_22023,N_21922);
and U22288 (N_22288,N_22113,N_21988);
nand U22289 (N_22289,N_21910,N_22029);
nor U22290 (N_22290,N_21900,N_21950);
or U22291 (N_22291,N_21971,N_21976);
or U22292 (N_22292,N_21980,N_22151);
or U22293 (N_22293,N_21925,N_21977);
nor U22294 (N_22294,N_22124,N_21981);
nand U22295 (N_22295,N_21908,N_22176);
and U22296 (N_22296,N_21978,N_22065);
or U22297 (N_22297,N_21946,N_22194);
nand U22298 (N_22298,N_21952,N_22139);
nand U22299 (N_22299,N_21983,N_22071);
nor U22300 (N_22300,N_21947,N_22008);
or U22301 (N_22301,N_22172,N_22049);
nand U22302 (N_22302,N_21928,N_22134);
or U22303 (N_22303,N_21943,N_22184);
nand U22304 (N_22304,N_21998,N_21918);
nor U22305 (N_22305,N_22073,N_22053);
nand U22306 (N_22306,N_22114,N_22128);
nor U22307 (N_22307,N_21936,N_22025);
or U22308 (N_22308,N_21979,N_22110);
or U22309 (N_22309,N_22050,N_22133);
nand U22310 (N_22310,N_22136,N_22146);
nor U22311 (N_22311,N_21921,N_22006);
nand U22312 (N_22312,N_22021,N_22144);
or U22313 (N_22313,N_22044,N_22153);
and U22314 (N_22314,N_22078,N_22135);
and U22315 (N_22315,N_22048,N_22032);
nor U22316 (N_22316,N_21975,N_22026);
nor U22317 (N_22317,N_22017,N_21993);
xor U22318 (N_22318,N_22132,N_22093);
or U22319 (N_22319,N_22115,N_22175);
nand U22320 (N_22320,N_22117,N_22098);
or U22321 (N_22321,N_22125,N_22164);
nor U22322 (N_22322,N_22196,N_22162);
and U22323 (N_22323,N_22188,N_22090);
or U22324 (N_22324,N_22119,N_22037);
nand U22325 (N_22325,N_21912,N_21901);
nand U22326 (N_22326,N_22046,N_21919);
nor U22327 (N_22327,N_21962,N_21956);
nand U22328 (N_22328,N_22011,N_22022);
nand U22329 (N_22329,N_21913,N_22092);
nor U22330 (N_22330,N_21958,N_22178);
nand U22331 (N_22331,N_21916,N_22147);
or U22332 (N_22332,N_22031,N_22013);
xnor U22333 (N_22333,N_22143,N_21937);
nor U22334 (N_22334,N_21924,N_21951);
xor U22335 (N_22335,N_22009,N_22197);
or U22336 (N_22336,N_21974,N_22015);
nand U22337 (N_22337,N_21940,N_22159);
xor U22338 (N_22338,N_22131,N_22077);
and U22339 (N_22339,N_21969,N_21984);
nor U22340 (N_22340,N_21923,N_21905);
and U22341 (N_22341,N_21995,N_22160);
nor U22342 (N_22342,N_21963,N_21929);
and U22343 (N_22343,N_22095,N_22003);
xor U22344 (N_22344,N_21959,N_22035);
nor U22345 (N_22345,N_22107,N_21970);
or U22346 (N_22346,N_22016,N_22059);
nand U22347 (N_22347,N_22080,N_22067);
xor U22348 (N_22348,N_21968,N_22183);
xnor U22349 (N_22349,N_22158,N_22142);
xnor U22350 (N_22350,N_21931,N_22092);
and U22351 (N_22351,N_22160,N_22189);
xnor U22352 (N_22352,N_22136,N_22115);
nand U22353 (N_22353,N_22037,N_22132);
or U22354 (N_22354,N_22185,N_22153);
or U22355 (N_22355,N_22191,N_22074);
xor U22356 (N_22356,N_22054,N_22093);
nand U22357 (N_22357,N_22127,N_22132);
nand U22358 (N_22358,N_22024,N_21995);
nor U22359 (N_22359,N_21902,N_22073);
nor U22360 (N_22360,N_21959,N_22175);
and U22361 (N_22361,N_21921,N_22168);
or U22362 (N_22362,N_21981,N_21946);
or U22363 (N_22363,N_22173,N_22044);
xnor U22364 (N_22364,N_21928,N_22148);
and U22365 (N_22365,N_22063,N_21968);
nor U22366 (N_22366,N_22084,N_22122);
nand U22367 (N_22367,N_22177,N_22082);
xor U22368 (N_22368,N_22168,N_22115);
nor U22369 (N_22369,N_22011,N_22170);
or U22370 (N_22370,N_21976,N_22003);
nor U22371 (N_22371,N_22150,N_22027);
nor U22372 (N_22372,N_22012,N_22145);
nand U22373 (N_22373,N_21953,N_22152);
nand U22374 (N_22374,N_22086,N_21909);
xnor U22375 (N_22375,N_22177,N_22156);
nor U22376 (N_22376,N_22020,N_22186);
and U22377 (N_22377,N_22196,N_22193);
nand U22378 (N_22378,N_22176,N_21966);
and U22379 (N_22379,N_22022,N_22152);
nor U22380 (N_22380,N_21911,N_22155);
and U22381 (N_22381,N_21997,N_22081);
xnor U22382 (N_22382,N_22065,N_22076);
nor U22383 (N_22383,N_22094,N_21908);
and U22384 (N_22384,N_22135,N_22121);
nor U22385 (N_22385,N_21959,N_22032);
nand U22386 (N_22386,N_22111,N_21991);
xnor U22387 (N_22387,N_22009,N_21904);
nor U22388 (N_22388,N_22102,N_22076);
or U22389 (N_22389,N_22110,N_21920);
xor U22390 (N_22390,N_22164,N_22094);
or U22391 (N_22391,N_21993,N_22105);
xnor U22392 (N_22392,N_22197,N_22189);
xor U22393 (N_22393,N_22013,N_21978);
xnor U22394 (N_22394,N_22018,N_22015);
nor U22395 (N_22395,N_22182,N_22162);
nor U22396 (N_22396,N_22138,N_21947);
nand U22397 (N_22397,N_22067,N_22042);
and U22398 (N_22398,N_22055,N_22161);
nand U22399 (N_22399,N_22132,N_21949);
and U22400 (N_22400,N_22095,N_22027);
nand U22401 (N_22401,N_22026,N_22175);
or U22402 (N_22402,N_22135,N_22101);
or U22403 (N_22403,N_22054,N_22026);
or U22404 (N_22404,N_22148,N_21938);
nor U22405 (N_22405,N_22195,N_21999);
xor U22406 (N_22406,N_22157,N_21920);
or U22407 (N_22407,N_22190,N_22055);
or U22408 (N_22408,N_21947,N_21924);
and U22409 (N_22409,N_21981,N_22048);
and U22410 (N_22410,N_21931,N_22080);
nand U22411 (N_22411,N_22184,N_22024);
xnor U22412 (N_22412,N_21945,N_21992);
or U22413 (N_22413,N_22094,N_22035);
nand U22414 (N_22414,N_22045,N_22123);
nand U22415 (N_22415,N_21993,N_21992);
and U22416 (N_22416,N_22065,N_22178);
nand U22417 (N_22417,N_22152,N_22010);
xnor U22418 (N_22418,N_22028,N_21968);
nor U22419 (N_22419,N_21942,N_21914);
and U22420 (N_22420,N_22143,N_22183);
nor U22421 (N_22421,N_22156,N_21937);
or U22422 (N_22422,N_22010,N_21969);
nand U22423 (N_22423,N_21975,N_22137);
nor U22424 (N_22424,N_22035,N_22024);
nor U22425 (N_22425,N_22062,N_22139);
and U22426 (N_22426,N_22165,N_22083);
nor U22427 (N_22427,N_22048,N_21948);
and U22428 (N_22428,N_22131,N_21999);
nand U22429 (N_22429,N_22069,N_22086);
nand U22430 (N_22430,N_21945,N_21960);
or U22431 (N_22431,N_22179,N_22169);
xnor U22432 (N_22432,N_22112,N_21995);
xnor U22433 (N_22433,N_22112,N_22186);
nor U22434 (N_22434,N_22059,N_22024);
and U22435 (N_22435,N_22078,N_21998);
nor U22436 (N_22436,N_22135,N_22125);
nand U22437 (N_22437,N_22176,N_21950);
nor U22438 (N_22438,N_21993,N_22175);
nand U22439 (N_22439,N_22114,N_21905);
nand U22440 (N_22440,N_22169,N_22184);
xor U22441 (N_22441,N_22196,N_22035);
and U22442 (N_22442,N_21926,N_22024);
or U22443 (N_22443,N_21917,N_21900);
xnor U22444 (N_22444,N_21995,N_22080);
nor U22445 (N_22445,N_21919,N_21913);
xnor U22446 (N_22446,N_22144,N_22198);
and U22447 (N_22447,N_22119,N_21937);
nor U22448 (N_22448,N_22148,N_22195);
or U22449 (N_22449,N_22130,N_21966);
and U22450 (N_22450,N_22048,N_22091);
nand U22451 (N_22451,N_22120,N_22113);
nor U22452 (N_22452,N_21938,N_22125);
xnor U22453 (N_22453,N_22030,N_21994);
nand U22454 (N_22454,N_22062,N_22006);
nand U22455 (N_22455,N_22065,N_22075);
nand U22456 (N_22456,N_21925,N_22133);
xnor U22457 (N_22457,N_22089,N_22045);
xnor U22458 (N_22458,N_21955,N_22191);
and U22459 (N_22459,N_22107,N_21960);
or U22460 (N_22460,N_22072,N_22164);
xor U22461 (N_22461,N_21970,N_21922);
nand U22462 (N_22462,N_22165,N_21971);
and U22463 (N_22463,N_22129,N_22198);
or U22464 (N_22464,N_21962,N_22079);
nand U22465 (N_22465,N_21993,N_21958);
xor U22466 (N_22466,N_21994,N_22106);
xnor U22467 (N_22467,N_21958,N_22073);
nor U22468 (N_22468,N_21984,N_21915);
nor U22469 (N_22469,N_22189,N_22066);
nand U22470 (N_22470,N_22066,N_22002);
or U22471 (N_22471,N_21901,N_21925);
and U22472 (N_22472,N_21983,N_21975);
or U22473 (N_22473,N_22062,N_22073);
or U22474 (N_22474,N_21959,N_22081);
nor U22475 (N_22475,N_21972,N_21935);
and U22476 (N_22476,N_22026,N_22185);
xor U22477 (N_22477,N_22133,N_22135);
nand U22478 (N_22478,N_21979,N_22151);
and U22479 (N_22479,N_22102,N_21980);
and U22480 (N_22480,N_22048,N_22085);
nor U22481 (N_22481,N_21934,N_22189);
and U22482 (N_22482,N_21982,N_21970);
or U22483 (N_22483,N_21963,N_21971);
nor U22484 (N_22484,N_21979,N_22152);
nor U22485 (N_22485,N_22158,N_21904);
nand U22486 (N_22486,N_21971,N_22046);
xor U22487 (N_22487,N_21968,N_22082);
nand U22488 (N_22488,N_22056,N_22023);
and U22489 (N_22489,N_22111,N_22063);
xnor U22490 (N_22490,N_21939,N_22097);
nor U22491 (N_22491,N_21921,N_21929);
nand U22492 (N_22492,N_22103,N_22036);
nand U22493 (N_22493,N_22094,N_22075);
nor U22494 (N_22494,N_22022,N_21998);
xnor U22495 (N_22495,N_22065,N_21916);
nand U22496 (N_22496,N_21961,N_22081);
xnor U22497 (N_22497,N_22046,N_22039);
nor U22498 (N_22498,N_22099,N_21950);
nand U22499 (N_22499,N_22131,N_22003);
and U22500 (N_22500,N_22283,N_22412);
nand U22501 (N_22501,N_22256,N_22437);
or U22502 (N_22502,N_22278,N_22456);
or U22503 (N_22503,N_22353,N_22221);
nor U22504 (N_22504,N_22424,N_22428);
xor U22505 (N_22505,N_22472,N_22374);
or U22506 (N_22506,N_22457,N_22240);
nor U22507 (N_22507,N_22210,N_22388);
nand U22508 (N_22508,N_22406,N_22433);
or U22509 (N_22509,N_22325,N_22316);
and U22510 (N_22510,N_22274,N_22265);
nor U22511 (N_22511,N_22298,N_22461);
xnor U22512 (N_22512,N_22452,N_22273);
and U22513 (N_22513,N_22332,N_22211);
xnor U22514 (N_22514,N_22365,N_22276);
nor U22515 (N_22515,N_22259,N_22431);
or U22516 (N_22516,N_22225,N_22370);
nor U22517 (N_22517,N_22207,N_22439);
xor U22518 (N_22518,N_22268,N_22345);
and U22519 (N_22519,N_22277,N_22434);
xor U22520 (N_22520,N_22432,N_22214);
xor U22521 (N_22521,N_22385,N_22460);
or U22522 (N_22522,N_22299,N_22441);
or U22523 (N_22523,N_22425,N_22344);
xnor U22524 (N_22524,N_22422,N_22377);
nor U22525 (N_22525,N_22336,N_22464);
xnor U22526 (N_22526,N_22258,N_22414);
xnor U22527 (N_22527,N_22486,N_22279);
and U22528 (N_22528,N_22389,N_22384);
and U22529 (N_22529,N_22416,N_22409);
xnor U22530 (N_22530,N_22242,N_22339);
xor U22531 (N_22531,N_22322,N_22481);
or U22532 (N_22532,N_22371,N_22338);
nand U22533 (N_22533,N_22307,N_22466);
nor U22534 (N_22534,N_22482,N_22397);
or U22535 (N_22535,N_22287,N_22218);
nor U22536 (N_22536,N_22394,N_22266);
xor U22537 (N_22537,N_22204,N_22443);
and U22538 (N_22538,N_22224,N_22487);
xnor U22539 (N_22539,N_22491,N_22228);
nand U22540 (N_22540,N_22205,N_22324);
nor U22541 (N_22541,N_22230,N_22444);
xnor U22542 (N_22542,N_22311,N_22251);
xnor U22543 (N_22543,N_22216,N_22270);
xnor U22544 (N_22544,N_22372,N_22390);
and U22545 (N_22545,N_22420,N_22304);
or U22546 (N_22546,N_22354,N_22286);
nand U22547 (N_22547,N_22262,N_22368);
or U22548 (N_22548,N_22290,N_22227);
and U22549 (N_22549,N_22355,N_22260);
nand U22550 (N_22550,N_22296,N_22285);
and U22551 (N_22551,N_22471,N_22474);
and U22552 (N_22552,N_22253,N_22342);
xnor U22553 (N_22553,N_22319,N_22326);
xnor U22554 (N_22554,N_22217,N_22320);
nor U22555 (N_22555,N_22349,N_22475);
xnor U22556 (N_22556,N_22300,N_22301);
or U22557 (N_22557,N_22328,N_22498);
nand U22558 (N_22558,N_22243,N_22436);
xnor U22559 (N_22559,N_22423,N_22426);
xor U22560 (N_22560,N_22238,N_22239);
nand U22561 (N_22561,N_22459,N_22312);
and U22562 (N_22562,N_22293,N_22490);
xnor U22563 (N_22563,N_22333,N_22493);
nand U22564 (N_22564,N_22415,N_22295);
nand U22565 (N_22565,N_22418,N_22245);
nor U22566 (N_22566,N_22231,N_22201);
nor U22567 (N_22567,N_22376,N_22302);
or U22568 (N_22568,N_22395,N_22446);
xor U22569 (N_22569,N_22383,N_22366);
or U22570 (N_22570,N_22494,N_22484);
and U22571 (N_22571,N_22408,N_22367);
nor U22572 (N_22572,N_22246,N_22308);
nand U22573 (N_22573,N_22476,N_22249);
nand U22574 (N_22574,N_22363,N_22232);
nor U22575 (N_22575,N_22369,N_22313);
or U22576 (N_22576,N_22226,N_22241);
nand U22577 (N_22577,N_22222,N_22335);
or U22578 (N_22578,N_22417,N_22236);
nor U22579 (N_22579,N_22361,N_22254);
or U22580 (N_22580,N_22407,N_22220);
xor U22581 (N_22581,N_22250,N_22386);
nand U22582 (N_22582,N_22378,N_22359);
nand U22583 (N_22583,N_22483,N_22318);
nor U22584 (N_22584,N_22234,N_22309);
nor U22585 (N_22585,N_22334,N_22310);
and U22586 (N_22586,N_22393,N_22435);
xor U22587 (N_22587,N_22450,N_22429);
and U22588 (N_22588,N_22213,N_22496);
or U22589 (N_22589,N_22467,N_22282);
and U22590 (N_22590,N_22297,N_22479);
nand U22591 (N_22591,N_22458,N_22215);
xnor U22592 (N_22592,N_22305,N_22404);
xor U22593 (N_22593,N_22392,N_22350);
xor U22594 (N_22594,N_22317,N_22263);
or U22595 (N_22595,N_22375,N_22315);
or U22596 (N_22596,N_22454,N_22488);
nor U22597 (N_22597,N_22244,N_22427);
nor U22598 (N_22598,N_22288,N_22212);
or U22599 (N_22599,N_22399,N_22379);
xnor U22600 (N_22600,N_22411,N_22272);
xnor U22601 (N_22601,N_22391,N_22264);
nor U22602 (N_22602,N_22237,N_22247);
nor U22603 (N_22603,N_22352,N_22473);
xor U22604 (N_22604,N_22327,N_22348);
and U22605 (N_22605,N_22430,N_22403);
nand U22606 (N_22606,N_22248,N_22480);
nand U22607 (N_22607,N_22200,N_22440);
xnor U22608 (N_22608,N_22402,N_22303);
nor U22609 (N_22609,N_22485,N_22492);
xnor U22610 (N_22610,N_22356,N_22323);
nand U22611 (N_22611,N_22292,N_22499);
xnor U22612 (N_22612,N_22497,N_22209);
nand U22613 (N_22613,N_22387,N_22438);
nand U22614 (N_22614,N_22410,N_22235);
and U22615 (N_22615,N_22291,N_22453);
xor U22616 (N_22616,N_22362,N_22255);
nor U22617 (N_22617,N_22252,N_22229);
nor U22618 (N_22618,N_22271,N_22208);
or U22619 (N_22619,N_22489,N_22449);
nor U22620 (N_22620,N_22495,N_22381);
nor U22621 (N_22621,N_22223,N_22445);
xnor U22622 (N_22622,N_22347,N_22364);
or U22623 (N_22623,N_22343,N_22346);
or U22624 (N_22624,N_22373,N_22463);
xnor U22625 (N_22625,N_22289,N_22267);
or U22626 (N_22626,N_22401,N_22470);
and U22627 (N_22627,N_22448,N_22398);
xnor U22628 (N_22628,N_22351,N_22447);
or U22629 (N_22629,N_22451,N_22203);
and U22630 (N_22630,N_22468,N_22321);
and U22631 (N_22631,N_22337,N_22284);
or U22632 (N_22632,N_22419,N_22357);
and U22633 (N_22633,N_22478,N_22413);
nor U22634 (N_22634,N_22465,N_22294);
or U22635 (N_22635,N_22455,N_22382);
xor U22636 (N_22636,N_22306,N_22400);
xor U22637 (N_22637,N_22261,N_22219);
or U22638 (N_22638,N_22442,N_22462);
or U22639 (N_22639,N_22421,N_22280);
and U22640 (N_22640,N_22396,N_22331);
or U22641 (N_22641,N_22269,N_22275);
nor U22642 (N_22642,N_22233,N_22360);
nor U22643 (N_22643,N_22329,N_22469);
nand U22644 (N_22644,N_22405,N_22281);
or U22645 (N_22645,N_22477,N_22314);
xor U22646 (N_22646,N_22257,N_22340);
or U22647 (N_22647,N_22206,N_22380);
and U22648 (N_22648,N_22341,N_22358);
nand U22649 (N_22649,N_22330,N_22202);
nor U22650 (N_22650,N_22332,N_22402);
nand U22651 (N_22651,N_22390,N_22373);
or U22652 (N_22652,N_22495,N_22418);
nor U22653 (N_22653,N_22407,N_22489);
or U22654 (N_22654,N_22291,N_22369);
nand U22655 (N_22655,N_22377,N_22240);
xor U22656 (N_22656,N_22209,N_22284);
or U22657 (N_22657,N_22354,N_22392);
or U22658 (N_22658,N_22462,N_22394);
nor U22659 (N_22659,N_22261,N_22386);
and U22660 (N_22660,N_22378,N_22412);
or U22661 (N_22661,N_22385,N_22277);
and U22662 (N_22662,N_22297,N_22354);
and U22663 (N_22663,N_22309,N_22279);
xnor U22664 (N_22664,N_22294,N_22239);
or U22665 (N_22665,N_22315,N_22330);
or U22666 (N_22666,N_22309,N_22275);
or U22667 (N_22667,N_22349,N_22414);
and U22668 (N_22668,N_22464,N_22234);
nor U22669 (N_22669,N_22238,N_22202);
nand U22670 (N_22670,N_22431,N_22234);
and U22671 (N_22671,N_22271,N_22277);
nand U22672 (N_22672,N_22399,N_22473);
xor U22673 (N_22673,N_22247,N_22418);
or U22674 (N_22674,N_22388,N_22249);
nor U22675 (N_22675,N_22343,N_22202);
xor U22676 (N_22676,N_22433,N_22393);
nor U22677 (N_22677,N_22493,N_22325);
or U22678 (N_22678,N_22412,N_22495);
and U22679 (N_22679,N_22321,N_22294);
xnor U22680 (N_22680,N_22377,N_22393);
or U22681 (N_22681,N_22479,N_22243);
nand U22682 (N_22682,N_22289,N_22318);
nand U22683 (N_22683,N_22499,N_22482);
or U22684 (N_22684,N_22207,N_22297);
xor U22685 (N_22685,N_22498,N_22284);
nor U22686 (N_22686,N_22217,N_22444);
xnor U22687 (N_22687,N_22402,N_22421);
nor U22688 (N_22688,N_22458,N_22267);
nor U22689 (N_22689,N_22475,N_22292);
nor U22690 (N_22690,N_22230,N_22388);
nand U22691 (N_22691,N_22490,N_22376);
or U22692 (N_22692,N_22435,N_22437);
and U22693 (N_22693,N_22488,N_22450);
xor U22694 (N_22694,N_22289,N_22334);
xnor U22695 (N_22695,N_22393,N_22329);
and U22696 (N_22696,N_22405,N_22383);
nand U22697 (N_22697,N_22366,N_22395);
nand U22698 (N_22698,N_22451,N_22253);
nand U22699 (N_22699,N_22293,N_22223);
xnor U22700 (N_22700,N_22410,N_22319);
xor U22701 (N_22701,N_22354,N_22350);
nand U22702 (N_22702,N_22357,N_22262);
xnor U22703 (N_22703,N_22335,N_22279);
and U22704 (N_22704,N_22342,N_22493);
and U22705 (N_22705,N_22344,N_22249);
and U22706 (N_22706,N_22487,N_22348);
and U22707 (N_22707,N_22270,N_22340);
xnor U22708 (N_22708,N_22428,N_22449);
xor U22709 (N_22709,N_22490,N_22406);
and U22710 (N_22710,N_22270,N_22413);
nand U22711 (N_22711,N_22434,N_22359);
and U22712 (N_22712,N_22478,N_22397);
and U22713 (N_22713,N_22417,N_22200);
nor U22714 (N_22714,N_22251,N_22427);
nor U22715 (N_22715,N_22288,N_22466);
and U22716 (N_22716,N_22319,N_22214);
or U22717 (N_22717,N_22286,N_22236);
xnor U22718 (N_22718,N_22220,N_22362);
nor U22719 (N_22719,N_22368,N_22271);
xor U22720 (N_22720,N_22338,N_22346);
nand U22721 (N_22721,N_22480,N_22435);
nand U22722 (N_22722,N_22415,N_22240);
or U22723 (N_22723,N_22469,N_22338);
nand U22724 (N_22724,N_22247,N_22367);
or U22725 (N_22725,N_22248,N_22484);
and U22726 (N_22726,N_22291,N_22305);
nor U22727 (N_22727,N_22477,N_22270);
xnor U22728 (N_22728,N_22413,N_22297);
nand U22729 (N_22729,N_22339,N_22463);
xnor U22730 (N_22730,N_22400,N_22357);
and U22731 (N_22731,N_22374,N_22489);
xor U22732 (N_22732,N_22283,N_22353);
xnor U22733 (N_22733,N_22213,N_22454);
nand U22734 (N_22734,N_22219,N_22273);
or U22735 (N_22735,N_22231,N_22432);
nor U22736 (N_22736,N_22366,N_22465);
and U22737 (N_22737,N_22362,N_22277);
or U22738 (N_22738,N_22458,N_22391);
nor U22739 (N_22739,N_22226,N_22355);
and U22740 (N_22740,N_22246,N_22344);
or U22741 (N_22741,N_22282,N_22367);
or U22742 (N_22742,N_22303,N_22232);
or U22743 (N_22743,N_22328,N_22281);
xnor U22744 (N_22744,N_22449,N_22283);
xor U22745 (N_22745,N_22249,N_22240);
or U22746 (N_22746,N_22271,N_22492);
nand U22747 (N_22747,N_22433,N_22499);
and U22748 (N_22748,N_22428,N_22252);
or U22749 (N_22749,N_22273,N_22233);
nor U22750 (N_22750,N_22356,N_22240);
and U22751 (N_22751,N_22452,N_22265);
nor U22752 (N_22752,N_22415,N_22201);
xnor U22753 (N_22753,N_22313,N_22406);
and U22754 (N_22754,N_22439,N_22429);
nand U22755 (N_22755,N_22397,N_22299);
and U22756 (N_22756,N_22410,N_22467);
xnor U22757 (N_22757,N_22290,N_22374);
nand U22758 (N_22758,N_22250,N_22315);
xor U22759 (N_22759,N_22362,N_22453);
nor U22760 (N_22760,N_22264,N_22378);
nor U22761 (N_22761,N_22456,N_22372);
and U22762 (N_22762,N_22466,N_22204);
xor U22763 (N_22763,N_22339,N_22392);
nand U22764 (N_22764,N_22359,N_22446);
nand U22765 (N_22765,N_22343,N_22347);
xnor U22766 (N_22766,N_22275,N_22314);
nand U22767 (N_22767,N_22258,N_22381);
nand U22768 (N_22768,N_22212,N_22255);
and U22769 (N_22769,N_22492,N_22207);
and U22770 (N_22770,N_22392,N_22415);
or U22771 (N_22771,N_22449,N_22463);
nor U22772 (N_22772,N_22331,N_22478);
xor U22773 (N_22773,N_22447,N_22368);
or U22774 (N_22774,N_22266,N_22268);
nand U22775 (N_22775,N_22365,N_22462);
nor U22776 (N_22776,N_22254,N_22230);
or U22777 (N_22777,N_22393,N_22313);
and U22778 (N_22778,N_22302,N_22243);
or U22779 (N_22779,N_22319,N_22341);
nor U22780 (N_22780,N_22460,N_22352);
or U22781 (N_22781,N_22202,N_22368);
and U22782 (N_22782,N_22320,N_22256);
xor U22783 (N_22783,N_22239,N_22430);
nor U22784 (N_22784,N_22463,N_22270);
nand U22785 (N_22785,N_22227,N_22215);
and U22786 (N_22786,N_22385,N_22226);
nand U22787 (N_22787,N_22322,N_22228);
nor U22788 (N_22788,N_22318,N_22377);
nand U22789 (N_22789,N_22289,N_22386);
xnor U22790 (N_22790,N_22432,N_22475);
nand U22791 (N_22791,N_22444,N_22475);
nor U22792 (N_22792,N_22314,N_22435);
and U22793 (N_22793,N_22230,N_22252);
and U22794 (N_22794,N_22206,N_22403);
or U22795 (N_22795,N_22355,N_22455);
nand U22796 (N_22796,N_22299,N_22496);
nand U22797 (N_22797,N_22221,N_22286);
xnor U22798 (N_22798,N_22290,N_22318);
and U22799 (N_22799,N_22402,N_22344);
nor U22800 (N_22800,N_22763,N_22617);
xor U22801 (N_22801,N_22706,N_22574);
and U22802 (N_22802,N_22682,N_22510);
nand U22803 (N_22803,N_22699,N_22753);
nand U22804 (N_22804,N_22633,N_22775);
or U22805 (N_22805,N_22568,N_22500);
or U22806 (N_22806,N_22618,N_22695);
nand U22807 (N_22807,N_22790,N_22709);
nand U22808 (N_22808,N_22680,N_22615);
nand U22809 (N_22809,N_22592,N_22530);
and U22810 (N_22810,N_22623,N_22602);
or U22811 (N_22811,N_22789,N_22793);
nor U22812 (N_22812,N_22647,N_22521);
nand U22813 (N_22813,N_22750,N_22678);
and U22814 (N_22814,N_22721,N_22547);
xnor U22815 (N_22815,N_22628,N_22591);
and U22816 (N_22816,N_22771,N_22539);
xnor U22817 (N_22817,N_22584,N_22570);
nor U22818 (N_22818,N_22717,N_22794);
and U22819 (N_22819,N_22668,N_22774);
nor U22820 (N_22820,N_22579,N_22601);
and U22821 (N_22821,N_22693,N_22779);
xor U22822 (N_22822,N_22726,N_22754);
nor U22823 (N_22823,N_22517,N_22738);
and U22824 (N_22824,N_22590,N_22522);
nand U22825 (N_22825,N_22548,N_22605);
or U22826 (N_22826,N_22756,N_22519);
xor U22827 (N_22827,N_22666,N_22675);
or U22828 (N_22828,N_22515,N_22531);
nor U22829 (N_22829,N_22655,N_22652);
nor U22830 (N_22830,N_22528,N_22712);
xnor U22831 (N_22831,N_22550,N_22546);
xnor U22832 (N_22832,N_22578,N_22650);
nand U22833 (N_22833,N_22622,N_22659);
xor U22834 (N_22834,N_22799,N_22676);
nor U22835 (N_22835,N_22609,N_22733);
xnor U22836 (N_22836,N_22573,N_22506);
xnor U22837 (N_22837,N_22735,N_22569);
xnor U22838 (N_22838,N_22748,N_22757);
nand U22839 (N_22839,N_22543,N_22669);
nor U22840 (N_22840,N_22788,N_22671);
and U22841 (N_22841,N_22536,N_22729);
nor U22842 (N_22842,N_22612,N_22603);
nand U22843 (N_22843,N_22630,N_22684);
nand U22844 (N_22844,N_22713,N_22795);
nor U22845 (N_22845,N_22649,N_22632);
or U22846 (N_22846,N_22604,N_22782);
xnor U22847 (N_22847,N_22736,N_22556);
nand U22848 (N_22848,N_22672,N_22516);
nor U22849 (N_22849,N_22727,N_22777);
xor U22850 (N_22850,N_22724,N_22624);
nor U22851 (N_22851,N_22610,N_22532);
xnor U22852 (N_22852,N_22665,N_22648);
or U22853 (N_22853,N_22643,N_22714);
nand U22854 (N_22854,N_22744,N_22742);
nor U22855 (N_22855,N_22557,N_22765);
and U22856 (N_22856,N_22607,N_22747);
or U22857 (N_22857,N_22740,N_22577);
or U22858 (N_22858,N_22653,N_22798);
nor U22859 (N_22859,N_22527,N_22505);
nor U22860 (N_22860,N_22769,N_22581);
and U22861 (N_22861,N_22594,N_22638);
or U22862 (N_22862,N_22501,N_22762);
nand U22863 (N_22863,N_22778,N_22561);
nor U22864 (N_22864,N_22759,N_22772);
nor U22865 (N_22865,N_22502,N_22658);
and U22866 (N_22866,N_22707,N_22722);
nor U22867 (N_22867,N_22644,N_22796);
nand U22868 (N_22868,N_22585,N_22667);
xor U22869 (N_22869,N_22786,N_22723);
and U22870 (N_22870,N_22694,N_22639);
nor U22871 (N_22871,N_22525,N_22549);
nor U22872 (N_22872,N_22687,N_22711);
nor U22873 (N_22873,N_22563,N_22697);
nand U22874 (N_22874,N_22620,N_22529);
xnor U22875 (N_22875,N_22677,N_22596);
nand U22876 (N_22876,N_22634,N_22636);
nand U22877 (N_22877,N_22743,N_22673);
and U22878 (N_22878,N_22766,N_22567);
and U22879 (N_22879,N_22627,N_22719);
and U22880 (N_22880,N_22509,N_22507);
or U22881 (N_22881,N_22745,N_22580);
xnor U22882 (N_22882,N_22508,N_22692);
nand U22883 (N_22883,N_22646,N_22535);
nand U22884 (N_22884,N_22797,N_22732);
and U22885 (N_22885,N_22571,N_22552);
and U22886 (N_22886,N_22656,N_22688);
nand U22887 (N_22887,N_22651,N_22554);
or U22888 (N_22888,N_22503,N_22730);
xnor U22889 (N_22889,N_22504,N_22523);
or U22890 (N_22890,N_22588,N_22770);
nand U22891 (N_22891,N_22661,N_22597);
and U22892 (N_22892,N_22518,N_22690);
and U22893 (N_22893,N_22631,N_22749);
or U22894 (N_22894,N_22741,N_22701);
and U22895 (N_22895,N_22702,N_22514);
and U22896 (N_22896,N_22657,N_22737);
xor U22897 (N_22897,N_22582,N_22739);
nand U22898 (N_22898,N_22619,N_22511);
nand U22899 (N_22899,N_22758,N_22544);
xnor U22900 (N_22900,N_22642,N_22645);
nor U22901 (N_22901,N_22572,N_22686);
nand U22902 (N_22902,N_22513,N_22696);
or U22903 (N_22903,N_22613,N_22767);
or U22904 (N_22904,N_22553,N_22784);
or U22905 (N_22905,N_22512,N_22773);
xnor U22906 (N_22906,N_22614,N_22664);
or U22907 (N_22907,N_22559,N_22785);
xor U22908 (N_22908,N_22704,N_22595);
or U22909 (N_22909,N_22662,N_22761);
or U22910 (N_22910,N_22641,N_22755);
xnor U22911 (N_22911,N_22520,N_22708);
and U22912 (N_22912,N_22626,N_22608);
or U22913 (N_22913,N_22589,N_22599);
xor U22914 (N_22914,N_22751,N_22541);
nand U22915 (N_22915,N_22629,N_22685);
and U22916 (N_22916,N_22566,N_22560);
nor U22917 (N_22917,N_22640,N_22720);
and U22918 (N_22918,N_22526,N_22715);
xor U22919 (N_22919,N_22600,N_22681);
or U22920 (N_22920,N_22731,N_22674);
or U22921 (N_22921,N_22625,N_22524);
nor U22922 (N_22922,N_22576,N_22787);
nand U22923 (N_22923,N_22575,N_22781);
xnor U22924 (N_22924,N_22780,N_22545);
and U22925 (N_22925,N_22542,N_22586);
nor U22926 (N_22926,N_22562,N_22558);
nor U22927 (N_22927,N_22764,N_22768);
nor U22928 (N_22928,N_22654,N_22752);
or U22929 (N_22929,N_22564,N_22538);
nor U22930 (N_22930,N_22670,N_22663);
nand U22931 (N_22931,N_22616,N_22691);
and U22932 (N_22932,N_22587,N_22583);
nand U22933 (N_22933,N_22635,N_22660);
or U22934 (N_22934,N_22700,N_22791);
and U22935 (N_22935,N_22637,N_22593);
and U22936 (N_22936,N_22734,N_22621);
and U22937 (N_22937,N_22551,N_22728);
or U22938 (N_22938,N_22683,N_22703);
or U22939 (N_22939,N_22716,N_22606);
and U22940 (N_22940,N_22679,N_22698);
nand U22941 (N_22941,N_22760,N_22710);
or U22942 (N_22942,N_22565,N_22783);
and U22943 (N_22943,N_22792,N_22533);
xnor U22944 (N_22944,N_22598,N_22540);
nand U22945 (N_22945,N_22718,N_22725);
or U22946 (N_22946,N_22611,N_22705);
and U22947 (N_22947,N_22555,N_22689);
and U22948 (N_22948,N_22746,N_22534);
and U22949 (N_22949,N_22776,N_22537);
xnor U22950 (N_22950,N_22641,N_22625);
xor U22951 (N_22951,N_22748,N_22790);
xnor U22952 (N_22952,N_22660,N_22710);
and U22953 (N_22953,N_22518,N_22640);
or U22954 (N_22954,N_22718,N_22700);
nor U22955 (N_22955,N_22560,N_22773);
xnor U22956 (N_22956,N_22654,N_22785);
xor U22957 (N_22957,N_22607,N_22722);
nor U22958 (N_22958,N_22703,N_22515);
xor U22959 (N_22959,N_22621,N_22509);
nor U22960 (N_22960,N_22512,N_22578);
or U22961 (N_22961,N_22757,N_22552);
xnor U22962 (N_22962,N_22624,N_22604);
and U22963 (N_22963,N_22626,N_22629);
and U22964 (N_22964,N_22595,N_22749);
nand U22965 (N_22965,N_22565,N_22788);
nor U22966 (N_22966,N_22606,N_22523);
or U22967 (N_22967,N_22659,N_22794);
or U22968 (N_22968,N_22555,N_22663);
or U22969 (N_22969,N_22584,N_22631);
nor U22970 (N_22970,N_22518,N_22582);
xor U22971 (N_22971,N_22794,N_22602);
nand U22972 (N_22972,N_22612,N_22738);
and U22973 (N_22973,N_22510,N_22570);
nand U22974 (N_22974,N_22505,N_22780);
nand U22975 (N_22975,N_22571,N_22579);
nor U22976 (N_22976,N_22666,N_22517);
nand U22977 (N_22977,N_22530,N_22610);
and U22978 (N_22978,N_22690,N_22601);
xor U22979 (N_22979,N_22788,N_22662);
xnor U22980 (N_22980,N_22671,N_22654);
nand U22981 (N_22981,N_22645,N_22504);
nor U22982 (N_22982,N_22794,N_22771);
nand U22983 (N_22983,N_22527,N_22645);
xor U22984 (N_22984,N_22600,N_22602);
or U22985 (N_22985,N_22627,N_22516);
or U22986 (N_22986,N_22765,N_22692);
or U22987 (N_22987,N_22658,N_22693);
nor U22988 (N_22988,N_22687,N_22682);
or U22989 (N_22989,N_22693,N_22683);
and U22990 (N_22990,N_22759,N_22503);
xor U22991 (N_22991,N_22523,N_22710);
nand U22992 (N_22992,N_22680,N_22647);
and U22993 (N_22993,N_22623,N_22671);
and U22994 (N_22994,N_22767,N_22745);
nand U22995 (N_22995,N_22600,N_22664);
nand U22996 (N_22996,N_22765,N_22575);
xnor U22997 (N_22997,N_22732,N_22777);
nor U22998 (N_22998,N_22696,N_22522);
xnor U22999 (N_22999,N_22762,N_22720);
nor U23000 (N_23000,N_22657,N_22697);
or U23001 (N_23001,N_22669,N_22734);
nor U23002 (N_23002,N_22676,N_22679);
or U23003 (N_23003,N_22700,N_22659);
or U23004 (N_23004,N_22760,N_22667);
nor U23005 (N_23005,N_22751,N_22609);
or U23006 (N_23006,N_22743,N_22665);
or U23007 (N_23007,N_22595,N_22748);
or U23008 (N_23008,N_22525,N_22747);
xnor U23009 (N_23009,N_22703,N_22798);
nand U23010 (N_23010,N_22687,N_22616);
nand U23011 (N_23011,N_22628,N_22691);
or U23012 (N_23012,N_22693,N_22620);
xor U23013 (N_23013,N_22713,N_22630);
or U23014 (N_23014,N_22605,N_22791);
or U23015 (N_23015,N_22647,N_22539);
and U23016 (N_23016,N_22702,N_22599);
and U23017 (N_23017,N_22737,N_22515);
and U23018 (N_23018,N_22780,N_22563);
nor U23019 (N_23019,N_22716,N_22562);
or U23020 (N_23020,N_22770,N_22790);
xor U23021 (N_23021,N_22512,N_22743);
and U23022 (N_23022,N_22573,N_22640);
or U23023 (N_23023,N_22782,N_22687);
nor U23024 (N_23024,N_22554,N_22728);
xor U23025 (N_23025,N_22511,N_22527);
and U23026 (N_23026,N_22606,N_22613);
nand U23027 (N_23027,N_22721,N_22779);
nor U23028 (N_23028,N_22506,N_22536);
nand U23029 (N_23029,N_22612,N_22719);
xnor U23030 (N_23030,N_22799,N_22750);
nand U23031 (N_23031,N_22734,N_22739);
or U23032 (N_23032,N_22532,N_22501);
xor U23033 (N_23033,N_22749,N_22771);
and U23034 (N_23034,N_22661,N_22583);
or U23035 (N_23035,N_22745,N_22528);
or U23036 (N_23036,N_22594,N_22677);
xor U23037 (N_23037,N_22794,N_22721);
nand U23038 (N_23038,N_22612,N_22724);
or U23039 (N_23039,N_22778,N_22669);
nand U23040 (N_23040,N_22636,N_22725);
nand U23041 (N_23041,N_22675,N_22503);
xor U23042 (N_23042,N_22565,N_22634);
and U23043 (N_23043,N_22654,N_22726);
nand U23044 (N_23044,N_22709,N_22795);
or U23045 (N_23045,N_22669,N_22505);
xnor U23046 (N_23046,N_22599,N_22531);
nor U23047 (N_23047,N_22760,N_22749);
nand U23048 (N_23048,N_22711,N_22738);
and U23049 (N_23049,N_22518,N_22734);
nand U23050 (N_23050,N_22538,N_22590);
and U23051 (N_23051,N_22643,N_22571);
or U23052 (N_23052,N_22671,N_22520);
xor U23053 (N_23053,N_22727,N_22795);
nor U23054 (N_23054,N_22606,N_22746);
or U23055 (N_23055,N_22698,N_22570);
xnor U23056 (N_23056,N_22599,N_22796);
xnor U23057 (N_23057,N_22727,N_22735);
and U23058 (N_23058,N_22651,N_22569);
xor U23059 (N_23059,N_22726,N_22551);
and U23060 (N_23060,N_22660,N_22750);
or U23061 (N_23061,N_22558,N_22619);
and U23062 (N_23062,N_22654,N_22637);
nor U23063 (N_23063,N_22618,N_22622);
xnor U23064 (N_23064,N_22778,N_22638);
and U23065 (N_23065,N_22540,N_22758);
or U23066 (N_23066,N_22680,N_22748);
or U23067 (N_23067,N_22615,N_22685);
xor U23068 (N_23068,N_22683,N_22786);
or U23069 (N_23069,N_22771,N_22715);
nor U23070 (N_23070,N_22596,N_22604);
and U23071 (N_23071,N_22685,N_22581);
or U23072 (N_23072,N_22526,N_22696);
nor U23073 (N_23073,N_22640,N_22627);
and U23074 (N_23074,N_22621,N_22731);
nor U23075 (N_23075,N_22688,N_22613);
or U23076 (N_23076,N_22785,N_22703);
or U23077 (N_23077,N_22643,N_22671);
and U23078 (N_23078,N_22710,N_22714);
or U23079 (N_23079,N_22536,N_22606);
and U23080 (N_23080,N_22552,N_22768);
nor U23081 (N_23081,N_22571,N_22538);
xnor U23082 (N_23082,N_22606,N_22712);
or U23083 (N_23083,N_22710,N_22588);
nor U23084 (N_23084,N_22707,N_22748);
nand U23085 (N_23085,N_22765,N_22788);
nor U23086 (N_23086,N_22565,N_22556);
or U23087 (N_23087,N_22678,N_22779);
nand U23088 (N_23088,N_22706,N_22527);
and U23089 (N_23089,N_22786,N_22517);
or U23090 (N_23090,N_22730,N_22791);
nor U23091 (N_23091,N_22626,N_22685);
or U23092 (N_23092,N_22611,N_22672);
xnor U23093 (N_23093,N_22641,N_22511);
nand U23094 (N_23094,N_22689,N_22723);
and U23095 (N_23095,N_22502,N_22786);
xor U23096 (N_23096,N_22588,N_22627);
nor U23097 (N_23097,N_22771,N_22629);
nand U23098 (N_23098,N_22740,N_22766);
and U23099 (N_23099,N_22666,N_22553);
or U23100 (N_23100,N_22847,N_22886);
nand U23101 (N_23101,N_22864,N_23070);
nand U23102 (N_23102,N_23041,N_22943);
nand U23103 (N_23103,N_22889,N_23068);
nor U23104 (N_23104,N_22818,N_22994);
xnor U23105 (N_23105,N_22867,N_22995);
nor U23106 (N_23106,N_22916,N_22849);
or U23107 (N_23107,N_22858,N_22845);
xor U23108 (N_23108,N_22848,N_22925);
nor U23109 (N_23109,N_22972,N_22802);
xor U23110 (N_23110,N_22823,N_22969);
nand U23111 (N_23111,N_22963,N_22960);
nand U23112 (N_23112,N_22992,N_23037);
and U23113 (N_23113,N_22806,N_23001);
nand U23114 (N_23114,N_22839,N_22941);
or U23115 (N_23115,N_23042,N_22862);
nand U23116 (N_23116,N_22965,N_22819);
or U23117 (N_23117,N_23078,N_22974);
or U23118 (N_23118,N_22883,N_23036);
nand U23119 (N_23119,N_23004,N_23066);
nand U23120 (N_23120,N_22876,N_23019);
nor U23121 (N_23121,N_22826,N_22807);
nand U23122 (N_23122,N_22817,N_22966);
or U23123 (N_23123,N_22962,N_22846);
xor U23124 (N_23124,N_22815,N_23077);
nor U23125 (N_23125,N_23009,N_22860);
xnor U23126 (N_23126,N_22820,N_23047);
and U23127 (N_23127,N_23006,N_22953);
xnor U23128 (N_23128,N_22851,N_22875);
or U23129 (N_23129,N_23018,N_22959);
nor U23130 (N_23130,N_22859,N_22865);
and U23131 (N_23131,N_22927,N_23060);
or U23132 (N_23132,N_22948,N_22879);
nand U23133 (N_23133,N_23054,N_22863);
nand U23134 (N_23134,N_23026,N_22933);
or U23135 (N_23135,N_22811,N_23039);
or U23136 (N_23136,N_23000,N_22930);
and U23137 (N_23137,N_22982,N_23020);
and U23138 (N_23138,N_22829,N_22975);
nand U23139 (N_23139,N_23092,N_23096);
nor U23140 (N_23140,N_23098,N_23027);
nand U23141 (N_23141,N_23002,N_22989);
nor U23142 (N_23142,N_23012,N_23079);
xnor U23143 (N_23143,N_22956,N_22918);
nand U23144 (N_23144,N_22888,N_22996);
nand U23145 (N_23145,N_23014,N_22803);
or U23146 (N_23146,N_23071,N_23010);
and U23147 (N_23147,N_22840,N_22984);
or U23148 (N_23148,N_23062,N_22919);
and U23149 (N_23149,N_22850,N_22828);
xor U23150 (N_23150,N_22834,N_23017);
and U23151 (N_23151,N_22805,N_22800);
or U23152 (N_23152,N_23015,N_23011);
and U23153 (N_23153,N_22900,N_22866);
and U23154 (N_23154,N_22977,N_22999);
and U23155 (N_23155,N_22926,N_22801);
xor U23156 (N_23156,N_23072,N_22808);
nand U23157 (N_23157,N_23075,N_22920);
or U23158 (N_23158,N_22885,N_23097);
or U23159 (N_23159,N_23059,N_23055);
nand U23160 (N_23160,N_22874,N_23038);
and U23161 (N_23161,N_22830,N_22923);
xor U23162 (N_23162,N_22868,N_23034);
or U23163 (N_23163,N_22822,N_22946);
nor U23164 (N_23164,N_23046,N_22856);
nor U23165 (N_23165,N_23053,N_23030);
and U23166 (N_23166,N_22809,N_22968);
nand U23167 (N_23167,N_22832,N_22902);
and U23168 (N_23168,N_22877,N_22892);
and U23169 (N_23169,N_22951,N_22914);
or U23170 (N_23170,N_22852,N_23091);
and U23171 (N_23171,N_23048,N_22945);
nor U23172 (N_23172,N_22833,N_22928);
nor U23173 (N_23173,N_22993,N_22954);
xnor U23174 (N_23174,N_22821,N_23088);
nor U23175 (N_23175,N_22804,N_22952);
and U23176 (N_23176,N_22912,N_23067);
nor U23177 (N_23177,N_22841,N_22911);
and U23178 (N_23178,N_22986,N_22976);
xor U23179 (N_23179,N_22898,N_23090);
or U23180 (N_23180,N_23051,N_23087);
nor U23181 (N_23181,N_22981,N_23005);
or U23182 (N_23182,N_22907,N_22950);
or U23183 (N_23183,N_23099,N_22870);
nor U23184 (N_23184,N_22985,N_22831);
nor U23185 (N_23185,N_22924,N_22853);
nor U23186 (N_23186,N_22970,N_22838);
and U23187 (N_23187,N_22813,N_22882);
and U23188 (N_23188,N_22955,N_22979);
or U23189 (N_23189,N_22869,N_22964);
nand U23190 (N_23190,N_23095,N_22895);
xor U23191 (N_23191,N_22861,N_23003);
or U23192 (N_23192,N_23033,N_22987);
or U23193 (N_23193,N_23093,N_23094);
nor U23194 (N_23194,N_23013,N_23023);
and U23195 (N_23195,N_22922,N_22872);
and U23196 (N_23196,N_22896,N_22881);
nor U23197 (N_23197,N_22812,N_22947);
xor U23198 (N_23198,N_22936,N_22910);
or U23199 (N_23199,N_22942,N_22854);
xor U23200 (N_23200,N_23074,N_22871);
nor U23201 (N_23201,N_22837,N_22857);
or U23202 (N_23202,N_22901,N_22917);
xor U23203 (N_23203,N_22932,N_22938);
and U23204 (N_23204,N_22903,N_23025);
and U23205 (N_23205,N_23029,N_22988);
and U23206 (N_23206,N_22929,N_22921);
nor U23207 (N_23207,N_22961,N_23084);
nor U23208 (N_23208,N_22824,N_23050);
or U23209 (N_23209,N_22894,N_22997);
nor U23210 (N_23210,N_23021,N_23057);
nor U23211 (N_23211,N_23080,N_22810);
xnor U23212 (N_23212,N_23065,N_22887);
and U23213 (N_23213,N_22957,N_22880);
and U23214 (N_23214,N_23076,N_22873);
or U23215 (N_23215,N_22906,N_23016);
xor U23216 (N_23216,N_23056,N_23028);
and U23217 (N_23217,N_23043,N_22905);
xnor U23218 (N_23218,N_22884,N_22836);
or U23219 (N_23219,N_22971,N_23086);
xnor U23220 (N_23220,N_23089,N_22934);
xor U23221 (N_23221,N_22937,N_23031);
or U23222 (N_23222,N_22816,N_22958);
and U23223 (N_23223,N_23049,N_23052);
xor U23224 (N_23224,N_22915,N_23035);
xnor U23225 (N_23225,N_23064,N_22913);
xnor U23226 (N_23226,N_22931,N_23069);
and U23227 (N_23227,N_23007,N_22827);
xnor U23228 (N_23228,N_23008,N_22983);
xnor U23229 (N_23229,N_23032,N_22909);
and U23230 (N_23230,N_23024,N_22940);
nand U23231 (N_23231,N_22939,N_22897);
and U23232 (N_23232,N_22978,N_22967);
nand U23233 (N_23233,N_22980,N_23022);
xnor U23234 (N_23234,N_22814,N_23073);
nand U23235 (N_23235,N_23061,N_22949);
nand U23236 (N_23236,N_22973,N_22991);
or U23237 (N_23237,N_22843,N_22825);
and U23238 (N_23238,N_22844,N_22899);
xnor U23239 (N_23239,N_22998,N_22835);
nand U23240 (N_23240,N_23045,N_22904);
xnor U23241 (N_23241,N_23081,N_23083);
nand U23242 (N_23242,N_22990,N_22890);
or U23243 (N_23243,N_22842,N_23063);
nand U23244 (N_23244,N_23085,N_22855);
nor U23245 (N_23245,N_22908,N_22891);
nand U23246 (N_23246,N_22878,N_23058);
or U23247 (N_23247,N_22935,N_22893);
nand U23248 (N_23248,N_23082,N_23044);
or U23249 (N_23249,N_23040,N_22944);
nor U23250 (N_23250,N_23015,N_22967);
and U23251 (N_23251,N_22912,N_23095);
nor U23252 (N_23252,N_22810,N_22834);
nor U23253 (N_23253,N_22885,N_22822);
and U23254 (N_23254,N_23025,N_22954);
or U23255 (N_23255,N_22969,N_22915);
and U23256 (N_23256,N_22932,N_22984);
xnor U23257 (N_23257,N_22804,N_22812);
nor U23258 (N_23258,N_23007,N_23003);
or U23259 (N_23259,N_22980,N_23064);
and U23260 (N_23260,N_23062,N_22930);
nand U23261 (N_23261,N_22929,N_22920);
and U23262 (N_23262,N_22806,N_23004);
or U23263 (N_23263,N_23012,N_23058);
xor U23264 (N_23264,N_23028,N_23089);
or U23265 (N_23265,N_22974,N_22964);
or U23266 (N_23266,N_22973,N_23039);
or U23267 (N_23267,N_22810,N_22917);
or U23268 (N_23268,N_23000,N_22905);
or U23269 (N_23269,N_23025,N_22857);
nor U23270 (N_23270,N_22833,N_22990);
nand U23271 (N_23271,N_22864,N_22926);
nand U23272 (N_23272,N_22911,N_22927);
or U23273 (N_23273,N_22856,N_22920);
and U23274 (N_23274,N_22926,N_22997);
nor U23275 (N_23275,N_22933,N_22983);
or U23276 (N_23276,N_22897,N_22885);
nor U23277 (N_23277,N_22884,N_22859);
or U23278 (N_23278,N_22852,N_22907);
and U23279 (N_23279,N_23015,N_22907);
xor U23280 (N_23280,N_23041,N_23050);
nor U23281 (N_23281,N_22923,N_22846);
nor U23282 (N_23282,N_22930,N_22816);
xnor U23283 (N_23283,N_23087,N_22833);
xor U23284 (N_23284,N_22834,N_22906);
or U23285 (N_23285,N_22932,N_22887);
nand U23286 (N_23286,N_22813,N_22845);
nand U23287 (N_23287,N_23047,N_23043);
or U23288 (N_23288,N_22826,N_22966);
nand U23289 (N_23289,N_22814,N_22849);
or U23290 (N_23290,N_22962,N_22944);
nor U23291 (N_23291,N_23012,N_22948);
or U23292 (N_23292,N_23091,N_22918);
xor U23293 (N_23293,N_23065,N_22820);
xor U23294 (N_23294,N_23090,N_22997);
or U23295 (N_23295,N_22926,N_22986);
or U23296 (N_23296,N_22853,N_23054);
xor U23297 (N_23297,N_22926,N_22921);
nor U23298 (N_23298,N_22832,N_23078);
nor U23299 (N_23299,N_22837,N_22962);
or U23300 (N_23300,N_23092,N_22881);
or U23301 (N_23301,N_23065,N_22964);
nand U23302 (N_23302,N_22894,N_22943);
and U23303 (N_23303,N_22851,N_23028);
and U23304 (N_23304,N_23071,N_22967);
nor U23305 (N_23305,N_22975,N_22874);
and U23306 (N_23306,N_22956,N_22842);
nand U23307 (N_23307,N_22933,N_23027);
nand U23308 (N_23308,N_23098,N_23099);
nand U23309 (N_23309,N_22807,N_22874);
nor U23310 (N_23310,N_22873,N_23091);
xnor U23311 (N_23311,N_22965,N_22835);
nand U23312 (N_23312,N_23035,N_22846);
nor U23313 (N_23313,N_22967,N_22988);
xnor U23314 (N_23314,N_22944,N_22911);
nor U23315 (N_23315,N_22821,N_23085);
xor U23316 (N_23316,N_23051,N_23002);
or U23317 (N_23317,N_23024,N_22879);
or U23318 (N_23318,N_22922,N_22901);
or U23319 (N_23319,N_23012,N_22824);
and U23320 (N_23320,N_22934,N_22983);
and U23321 (N_23321,N_22860,N_22828);
xnor U23322 (N_23322,N_22838,N_23059);
or U23323 (N_23323,N_22917,N_22986);
and U23324 (N_23324,N_22968,N_23073);
nand U23325 (N_23325,N_22801,N_22871);
xnor U23326 (N_23326,N_22814,N_22974);
xnor U23327 (N_23327,N_22908,N_22942);
nor U23328 (N_23328,N_22872,N_23016);
xnor U23329 (N_23329,N_22972,N_23090);
xor U23330 (N_23330,N_22900,N_22804);
and U23331 (N_23331,N_23053,N_23046);
and U23332 (N_23332,N_23099,N_22999);
and U23333 (N_23333,N_23016,N_22831);
or U23334 (N_23334,N_23039,N_23076);
and U23335 (N_23335,N_22955,N_22943);
nor U23336 (N_23336,N_22853,N_22934);
or U23337 (N_23337,N_22969,N_22928);
and U23338 (N_23338,N_22947,N_23000);
nor U23339 (N_23339,N_22810,N_22909);
and U23340 (N_23340,N_22978,N_22973);
nor U23341 (N_23341,N_23023,N_22959);
or U23342 (N_23342,N_22916,N_22957);
nor U23343 (N_23343,N_22987,N_23004);
nand U23344 (N_23344,N_23006,N_22896);
or U23345 (N_23345,N_23031,N_23000);
xor U23346 (N_23346,N_23098,N_22989);
nor U23347 (N_23347,N_22901,N_23046);
nand U23348 (N_23348,N_22838,N_23025);
xnor U23349 (N_23349,N_23047,N_22860);
and U23350 (N_23350,N_23088,N_22979);
nand U23351 (N_23351,N_23080,N_23015);
xor U23352 (N_23352,N_22930,N_22946);
xor U23353 (N_23353,N_22872,N_22800);
nand U23354 (N_23354,N_22834,N_22812);
xnor U23355 (N_23355,N_23035,N_23050);
or U23356 (N_23356,N_23064,N_22952);
nor U23357 (N_23357,N_22839,N_22879);
and U23358 (N_23358,N_22927,N_22900);
and U23359 (N_23359,N_22821,N_23091);
xnor U23360 (N_23360,N_23011,N_23046);
or U23361 (N_23361,N_22842,N_22969);
and U23362 (N_23362,N_23043,N_23028);
or U23363 (N_23363,N_23054,N_23032);
xor U23364 (N_23364,N_22884,N_22844);
nand U23365 (N_23365,N_23034,N_22944);
nand U23366 (N_23366,N_23061,N_22919);
nor U23367 (N_23367,N_22930,N_23056);
or U23368 (N_23368,N_22904,N_22816);
xnor U23369 (N_23369,N_22973,N_22893);
nand U23370 (N_23370,N_22840,N_22897);
nand U23371 (N_23371,N_23089,N_22903);
or U23372 (N_23372,N_22813,N_22852);
xor U23373 (N_23373,N_22938,N_23007);
or U23374 (N_23374,N_22848,N_23032);
xor U23375 (N_23375,N_22949,N_22883);
nand U23376 (N_23376,N_23022,N_22842);
xnor U23377 (N_23377,N_23056,N_22873);
nor U23378 (N_23378,N_23068,N_23005);
or U23379 (N_23379,N_23086,N_22940);
xnor U23380 (N_23380,N_22901,N_22949);
nand U23381 (N_23381,N_22887,N_23046);
nor U23382 (N_23382,N_23090,N_22835);
nor U23383 (N_23383,N_22825,N_22957);
and U23384 (N_23384,N_22954,N_23061);
and U23385 (N_23385,N_22872,N_22975);
nand U23386 (N_23386,N_22851,N_23001);
and U23387 (N_23387,N_22970,N_22821);
nand U23388 (N_23388,N_23013,N_22866);
nor U23389 (N_23389,N_23022,N_22847);
nand U23390 (N_23390,N_23003,N_22927);
xnor U23391 (N_23391,N_22967,N_22806);
nor U23392 (N_23392,N_22822,N_22987);
nand U23393 (N_23393,N_22999,N_22896);
or U23394 (N_23394,N_22844,N_23071);
nor U23395 (N_23395,N_23083,N_22812);
xor U23396 (N_23396,N_23075,N_23032);
nand U23397 (N_23397,N_22805,N_22936);
nand U23398 (N_23398,N_23057,N_23035);
nor U23399 (N_23399,N_22951,N_23026);
and U23400 (N_23400,N_23202,N_23196);
or U23401 (N_23401,N_23132,N_23337);
or U23402 (N_23402,N_23248,N_23275);
nor U23403 (N_23403,N_23268,N_23242);
xor U23404 (N_23404,N_23367,N_23160);
and U23405 (N_23405,N_23375,N_23186);
nor U23406 (N_23406,N_23232,N_23321);
and U23407 (N_23407,N_23316,N_23287);
xor U23408 (N_23408,N_23201,N_23288);
xnor U23409 (N_23409,N_23263,N_23223);
or U23410 (N_23410,N_23168,N_23266);
nand U23411 (N_23411,N_23358,N_23347);
nand U23412 (N_23412,N_23306,N_23291);
or U23413 (N_23413,N_23159,N_23252);
xnor U23414 (N_23414,N_23125,N_23280);
and U23415 (N_23415,N_23397,N_23119);
and U23416 (N_23416,N_23224,N_23332);
and U23417 (N_23417,N_23244,N_23165);
xor U23418 (N_23418,N_23382,N_23378);
and U23419 (N_23419,N_23240,N_23210);
and U23420 (N_23420,N_23366,N_23187);
nor U23421 (N_23421,N_23258,N_23320);
xor U23422 (N_23422,N_23221,N_23310);
and U23423 (N_23423,N_23296,N_23117);
and U23424 (N_23424,N_23193,N_23178);
and U23425 (N_23425,N_23339,N_23345);
nor U23426 (N_23426,N_23396,N_23371);
nand U23427 (N_23427,N_23169,N_23365);
xor U23428 (N_23428,N_23215,N_23109);
nand U23429 (N_23429,N_23262,N_23220);
or U23430 (N_23430,N_23247,N_23254);
nor U23431 (N_23431,N_23318,N_23304);
nor U23432 (N_23432,N_23313,N_23189);
nor U23433 (N_23433,N_23317,N_23141);
nor U23434 (N_23434,N_23379,N_23206);
nor U23435 (N_23435,N_23342,N_23338);
or U23436 (N_23436,N_23239,N_23153);
nor U23437 (N_23437,N_23265,N_23108);
nor U23438 (N_23438,N_23324,N_23229);
nor U23439 (N_23439,N_23144,N_23302);
xnor U23440 (N_23440,N_23120,N_23185);
nor U23441 (N_23441,N_23179,N_23200);
xor U23442 (N_23442,N_23158,N_23286);
and U23443 (N_23443,N_23385,N_23162);
or U23444 (N_23444,N_23182,N_23100);
or U23445 (N_23445,N_23156,N_23173);
nand U23446 (N_23446,N_23194,N_23122);
or U23447 (N_23447,N_23389,N_23112);
and U23448 (N_23448,N_23136,N_23257);
nand U23449 (N_23449,N_23243,N_23138);
nor U23450 (N_23450,N_23219,N_23390);
nand U23451 (N_23451,N_23213,N_23103);
or U23452 (N_23452,N_23349,N_23155);
xnor U23453 (N_23453,N_23184,N_23361);
xnor U23454 (N_23454,N_23175,N_23134);
nor U23455 (N_23455,N_23340,N_23300);
xor U23456 (N_23456,N_23328,N_23373);
nor U23457 (N_23457,N_23163,N_23395);
or U23458 (N_23458,N_23391,N_23394);
and U23459 (N_23459,N_23250,N_23383);
nand U23460 (N_23460,N_23325,N_23272);
xor U23461 (N_23461,N_23102,N_23192);
xor U23462 (N_23462,N_23334,N_23131);
and U23463 (N_23463,N_23279,N_23166);
and U23464 (N_23464,N_23323,N_23350);
and U23465 (N_23465,N_23368,N_23128);
or U23466 (N_23466,N_23209,N_23249);
and U23467 (N_23467,N_23107,N_23148);
nand U23468 (N_23468,N_23298,N_23330);
nor U23469 (N_23469,N_23319,N_23203);
and U23470 (N_23470,N_23387,N_23113);
nor U23471 (N_23471,N_23135,N_23146);
nor U23472 (N_23472,N_23374,N_23301);
nand U23473 (N_23473,N_23253,N_23246);
and U23474 (N_23474,N_23157,N_23191);
nand U23475 (N_23475,N_23227,N_23237);
xnor U23476 (N_23476,N_23393,N_23362);
or U23477 (N_23477,N_23139,N_23376);
or U23478 (N_23478,N_23273,N_23151);
nand U23479 (N_23479,N_23147,N_23399);
and U23480 (N_23480,N_23176,N_23225);
or U23481 (N_23481,N_23177,N_23370);
nand U23482 (N_23482,N_23380,N_23284);
nand U23483 (N_23483,N_23343,N_23312);
or U23484 (N_23484,N_23212,N_23205);
xor U23485 (N_23485,N_23104,N_23398);
nand U23486 (N_23486,N_23110,N_23234);
nor U23487 (N_23487,N_23116,N_23384);
and U23488 (N_23488,N_23228,N_23336);
nor U23489 (N_23489,N_23233,N_23164);
nand U23490 (N_23490,N_23111,N_23124);
nor U23491 (N_23491,N_23211,N_23290);
nand U23492 (N_23492,N_23369,N_23230);
or U23493 (N_23493,N_23188,N_23129);
nor U23494 (N_23494,N_23303,N_23260);
xnor U23495 (N_23495,N_23207,N_23133);
xor U23496 (N_23496,N_23308,N_23142);
nand U23497 (N_23497,N_23359,N_23190);
and U23498 (N_23498,N_23314,N_23170);
nor U23499 (N_23499,N_23354,N_23217);
and U23500 (N_23500,N_23277,N_23335);
xnor U23501 (N_23501,N_23154,N_23114);
and U23502 (N_23502,N_23126,N_23259);
xnor U23503 (N_23503,N_23309,N_23241);
or U23504 (N_23504,N_23372,N_23145);
nor U23505 (N_23505,N_23333,N_23281);
xnor U23506 (N_23506,N_23305,N_23364);
or U23507 (N_23507,N_23115,N_23149);
nor U23508 (N_23508,N_23171,N_23236);
or U23509 (N_23509,N_23106,N_23282);
nor U23510 (N_23510,N_23222,N_23251);
or U23511 (N_23511,N_23167,N_23269);
or U23512 (N_23512,N_23355,N_23245);
or U23513 (N_23513,N_23276,N_23357);
and U23514 (N_23514,N_23181,N_23180);
nand U23515 (N_23515,N_23293,N_23255);
and U23516 (N_23516,N_23388,N_23331);
nand U23517 (N_23517,N_23392,N_23208);
or U23518 (N_23518,N_23183,N_23292);
or U23519 (N_23519,N_23121,N_23226);
xnor U23520 (N_23520,N_23214,N_23351);
or U23521 (N_23521,N_23197,N_23199);
and U23522 (N_23522,N_23307,N_23174);
nor U23523 (N_23523,N_23271,N_23381);
and U23524 (N_23524,N_23299,N_23315);
or U23525 (N_23525,N_23195,N_23137);
nor U23526 (N_23526,N_23274,N_23377);
or U23527 (N_23527,N_23295,N_23267);
nor U23528 (N_23528,N_23327,N_23285);
nor U23529 (N_23529,N_23261,N_23346);
nand U23530 (N_23530,N_23311,N_23152);
nor U23531 (N_23531,N_23353,N_23127);
nor U23532 (N_23532,N_23130,N_23231);
nand U23533 (N_23533,N_23204,N_23264);
or U23534 (N_23534,N_23278,N_23235);
nor U23535 (N_23535,N_23150,N_23386);
or U23536 (N_23536,N_23216,N_23289);
and U23537 (N_23537,N_23283,N_23198);
xor U23538 (N_23538,N_23297,N_23218);
nand U23539 (N_23539,N_23123,N_23352);
and U23540 (N_23540,N_23294,N_23238);
and U23541 (N_23541,N_23140,N_23322);
xor U23542 (N_23542,N_23326,N_23118);
or U23543 (N_23543,N_23105,N_23360);
xnor U23544 (N_23544,N_23256,N_23341);
nand U23545 (N_23545,N_23348,N_23356);
nand U23546 (N_23546,N_23363,N_23101);
nand U23547 (N_23547,N_23329,N_23161);
nor U23548 (N_23548,N_23172,N_23270);
nand U23549 (N_23549,N_23344,N_23143);
xor U23550 (N_23550,N_23235,N_23135);
and U23551 (N_23551,N_23221,N_23328);
nor U23552 (N_23552,N_23165,N_23108);
nand U23553 (N_23553,N_23246,N_23390);
or U23554 (N_23554,N_23379,N_23274);
nand U23555 (N_23555,N_23252,N_23371);
nand U23556 (N_23556,N_23123,N_23239);
and U23557 (N_23557,N_23229,N_23392);
nand U23558 (N_23558,N_23313,N_23326);
xnor U23559 (N_23559,N_23289,N_23297);
nand U23560 (N_23560,N_23387,N_23128);
or U23561 (N_23561,N_23169,N_23340);
and U23562 (N_23562,N_23204,N_23353);
and U23563 (N_23563,N_23193,N_23166);
and U23564 (N_23564,N_23195,N_23329);
and U23565 (N_23565,N_23108,N_23287);
or U23566 (N_23566,N_23298,N_23190);
nor U23567 (N_23567,N_23291,N_23166);
or U23568 (N_23568,N_23171,N_23125);
or U23569 (N_23569,N_23249,N_23215);
and U23570 (N_23570,N_23316,N_23175);
nand U23571 (N_23571,N_23327,N_23200);
nor U23572 (N_23572,N_23204,N_23133);
nor U23573 (N_23573,N_23197,N_23326);
nand U23574 (N_23574,N_23378,N_23155);
xor U23575 (N_23575,N_23395,N_23112);
nor U23576 (N_23576,N_23196,N_23285);
nand U23577 (N_23577,N_23114,N_23240);
xor U23578 (N_23578,N_23299,N_23158);
nand U23579 (N_23579,N_23291,N_23398);
or U23580 (N_23580,N_23215,N_23108);
nand U23581 (N_23581,N_23323,N_23235);
xnor U23582 (N_23582,N_23289,N_23363);
and U23583 (N_23583,N_23156,N_23116);
or U23584 (N_23584,N_23314,N_23348);
nor U23585 (N_23585,N_23115,N_23140);
nand U23586 (N_23586,N_23213,N_23381);
nor U23587 (N_23587,N_23178,N_23188);
xnor U23588 (N_23588,N_23336,N_23218);
nor U23589 (N_23589,N_23236,N_23138);
xnor U23590 (N_23590,N_23223,N_23335);
nor U23591 (N_23591,N_23205,N_23224);
xnor U23592 (N_23592,N_23300,N_23142);
xnor U23593 (N_23593,N_23238,N_23155);
or U23594 (N_23594,N_23129,N_23206);
and U23595 (N_23595,N_23329,N_23274);
nor U23596 (N_23596,N_23113,N_23209);
and U23597 (N_23597,N_23229,N_23108);
and U23598 (N_23598,N_23195,N_23239);
or U23599 (N_23599,N_23112,N_23349);
or U23600 (N_23600,N_23230,N_23158);
nand U23601 (N_23601,N_23384,N_23129);
or U23602 (N_23602,N_23197,N_23342);
nand U23603 (N_23603,N_23219,N_23398);
or U23604 (N_23604,N_23136,N_23316);
xor U23605 (N_23605,N_23356,N_23299);
nand U23606 (N_23606,N_23310,N_23363);
and U23607 (N_23607,N_23312,N_23246);
or U23608 (N_23608,N_23224,N_23335);
nor U23609 (N_23609,N_23167,N_23394);
xnor U23610 (N_23610,N_23338,N_23373);
nor U23611 (N_23611,N_23399,N_23384);
or U23612 (N_23612,N_23367,N_23195);
or U23613 (N_23613,N_23161,N_23189);
nand U23614 (N_23614,N_23227,N_23300);
nand U23615 (N_23615,N_23354,N_23231);
and U23616 (N_23616,N_23134,N_23207);
xnor U23617 (N_23617,N_23176,N_23312);
nor U23618 (N_23618,N_23389,N_23160);
nor U23619 (N_23619,N_23217,N_23345);
xor U23620 (N_23620,N_23349,N_23151);
nor U23621 (N_23621,N_23204,N_23335);
or U23622 (N_23622,N_23133,N_23300);
and U23623 (N_23623,N_23355,N_23200);
or U23624 (N_23624,N_23271,N_23322);
nor U23625 (N_23625,N_23271,N_23113);
nor U23626 (N_23626,N_23118,N_23198);
nor U23627 (N_23627,N_23266,N_23174);
xor U23628 (N_23628,N_23244,N_23121);
and U23629 (N_23629,N_23250,N_23207);
or U23630 (N_23630,N_23231,N_23163);
or U23631 (N_23631,N_23279,N_23324);
and U23632 (N_23632,N_23251,N_23366);
nand U23633 (N_23633,N_23324,N_23231);
nor U23634 (N_23634,N_23267,N_23135);
nor U23635 (N_23635,N_23287,N_23100);
nand U23636 (N_23636,N_23331,N_23189);
xnor U23637 (N_23637,N_23134,N_23310);
nand U23638 (N_23638,N_23342,N_23225);
and U23639 (N_23639,N_23182,N_23131);
or U23640 (N_23640,N_23323,N_23296);
and U23641 (N_23641,N_23168,N_23110);
or U23642 (N_23642,N_23253,N_23388);
or U23643 (N_23643,N_23266,N_23290);
xnor U23644 (N_23644,N_23237,N_23364);
nor U23645 (N_23645,N_23337,N_23103);
nand U23646 (N_23646,N_23173,N_23259);
nand U23647 (N_23647,N_23253,N_23118);
xor U23648 (N_23648,N_23375,N_23176);
nand U23649 (N_23649,N_23245,N_23318);
nand U23650 (N_23650,N_23282,N_23100);
xnor U23651 (N_23651,N_23324,N_23292);
nor U23652 (N_23652,N_23256,N_23361);
and U23653 (N_23653,N_23293,N_23397);
nor U23654 (N_23654,N_23148,N_23265);
xor U23655 (N_23655,N_23370,N_23112);
nand U23656 (N_23656,N_23221,N_23320);
or U23657 (N_23657,N_23127,N_23238);
nor U23658 (N_23658,N_23365,N_23100);
nand U23659 (N_23659,N_23334,N_23224);
or U23660 (N_23660,N_23172,N_23273);
xnor U23661 (N_23661,N_23302,N_23318);
xor U23662 (N_23662,N_23240,N_23353);
and U23663 (N_23663,N_23199,N_23203);
and U23664 (N_23664,N_23360,N_23285);
nor U23665 (N_23665,N_23347,N_23183);
xnor U23666 (N_23666,N_23193,N_23312);
xor U23667 (N_23667,N_23288,N_23244);
and U23668 (N_23668,N_23310,N_23255);
and U23669 (N_23669,N_23394,N_23105);
or U23670 (N_23670,N_23384,N_23350);
and U23671 (N_23671,N_23375,N_23136);
nor U23672 (N_23672,N_23312,N_23321);
or U23673 (N_23673,N_23372,N_23137);
nor U23674 (N_23674,N_23222,N_23206);
or U23675 (N_23675,N_23242,N_23320);
nor U23676 (N_23676,N_23249,N_23345);
and U23677 (N_23677,N_23298,N_23155);
nor U23678 (N_23678,N_23363,N_23141);
nor U23679 (N_23679,N_23322,N_23130);
xor U23680 (N_23680,N_23394,N_23182);
nand U23681 (N_23681,N_23197,N_23343);
and U23682 (N_23682,N_23255,N_23225);
or U23683 (N_23683,N_23357,N_23348);
xor U23684 (N_23684,N_23337,N_23106);
or U23685 (N_23685,N_23165,N_23304);
and U23686 (N_23686,N_23353,N_23211);
nor U23687 (N_23687,N_23228,N_23307);
or U23688 (N_23688,N_23348,N_23150);
nor U23689 (N_23689,N_23127,N_23150);
and U23690 (N_23690,N_23257,N_23224);
nor U23691 (N_23691,N_23154,N_23395);
or U23692 (N_23692,N_23112,N_23175);
and U23693 (N_23693,N_23349,N_23259);
or U23694 (N_23694,N_23154,N_23127);
nor U23695 (N_23695,N_23379,N_23398);
and U23696 (N_23696,N_23292,N_23172);
nor U23697 (N_23697,N_23272,N_23282);
nand U23698 (N_23698,N_23362,N_23213);
nor U23699 (N_23699,N_23154,N_23300);
nor U23700 (N_23700,N_23541,N_23611);
and U23701 (N_23701,N_23669,N_23489);
or U23702 (N_23702,N_23581,N_23675);
nand U23703 (N_23703,N_23658,N_23409);
xor U23704 (N_23704,N_23522,N_23661);
and U23705 (N_23705,N_23665,N_23504);
or U23706 (N_23706,N_23456,N_23556);
nand U23707 (N_23707,N_23627,N_23446);
xnor U23708 (N_23708,N_23411,N_23508);
and U23709 (N_23709,N_23485,N_23499);
and U23710 (N_23710,N_23653,N_23663);
nand U23711 (N_23711,N_23564,N_23625);
or U23712 (N_23712,N_23441,N_23496);
nand U23713 (N_23713,N_23563,N_23559);
nor U23714 (N_23714,N_23472,N_23596);
nor U23715 (N_23715,N_23694,N_23545);
xor U23716 (N_23716,N_23511,N_23547);
nor U23717 (N_23717,N_23652,N_23540);
and U23718 (N_23718,N_23461,N_23612);
nand U23719 (N_23719,N_23645,N_23530);
nand U23720 (N_23720,N_23413,N_23639);
xor U23721 (N_23721,N_23531,N_23647);
and U23722 (N_23722,N_23513,N_23417);
or U23723 (N_23723,N_23689,N_23697);
or U23724 (N_23724,N_23628,N_23475);
xor U23725 (N_23725,N_23687,N_23437);
nand U23726 (N_23726,N_23643,N_23699);
nand U23727 (N_23727,N_23660,N_23580);
nor U23728 (N_23728,N_23686,N_23400);
or U23729 (N_23729,N_23668,N_23671);
xor U23730 (N_23730,N_23442,N_23599);
or U23731 (N_23731,N_23623,N_23656);
or U23732 (N_23732,N_23664,N_23592);
or U23733 (N_23733,N_23458,N_23677);
nand U23734 (N_23734,N_23569,N_23479);
nand U23735 (N_23735,N_23698,N_23457);
nand U23736 (N_23736,N_23445,N_23609);
nor U23737 (N_23737,N_23488,N_23464);
and U23738 (N_23738,N_23607,N_23516);
nor U23739 (N_23739,N_23420,N_23512);
nor U23740 (N_23740,N_23659,N_23523);
and U23741 (N_23741,N_23492,N_23407);
xor U23742 (N_23742,N_23546,N_23598);
nand U23743 (N_23743,N_23486,N_23476);
xor U23744 (N_23744,N_23666,N_23493);
nor U23745 (N_23745,N_23535,N_23657);
xnor U23746 (N_23746,N_23520,N_23434);
or U23747 (N_23747,N_23593,N_23626);
nor U23748 (N_23748,N_23427,N_23480);
xnor U23749 (N_23749,N_23642,N_23415);
or U23750 (N_23750,N_23648,N_23405);
xor U23751 (N_23751,N_23690,N_23624);
nor U23752 (N_23752,N_23498,N_23528);
nor U23753 (N_23753,N_23662,N_23402);
xnor U23754 (N_23754,N_23575,N_23614);
nand U23755 (N_23755,N_23621,N_23558);
or U23756 (N_23756,N_23674,N_23544);
and U23757 (N_23757,N_23527,N_23421);
nand U23758 (N_23758,N_23565,N_23533);
nor U23759 (N_23759,N_23438,N_23510);
nand U23760 (N_23760,N_23422,N_23633);
or U23761 (N_23761,N_23622,N_23465);
xor U23762 (N_23762,N_23587,N_23601);
and U23763 (N_23763,N_23539,N_23574);
nor U23764 (N_23764,N_23518,N_23586);
xnor U23765 (N_23765,N_23495,N_23487);
xnor U23766 (N_23766,N_23632,N_23433);
and U23767 (N_23767,N_23497,N_23691);
or U23768 (N_23768,N_23631,N_23695);
nand U23769 (N_23769,N_23451,N_23406);
or U23770 (N_23770,N_23629,N_23473);
xnor U23771 (N_23771,N_23467,N_23655);
nor U23772 (N_23772,N_23579,N_23506);
xor U23773 (N_23773,N_23682,N_23517);
or U23774 (N_23774,N_23637,N_23505);
nor U23775 (N_23775,N_23426,N_23532);
xnor U23776 (N_23776,N_23432,N_23591);
xor U23777 (N_23777,N_23670,N_23572);
xor U23778 (N_23778,N_23678,N_23453);
xnor U23779 (N_23779,N_23685,N_23490);
nand U23780 (N_23780,N_23412,N_23447);
or U23781 (N_23781,N_23610,N_23693);
or U23782 (N_23782,N_23501,N_23606);
or U23783 (N_23783,N_23509,N_23435);
or U23784 (N_23784,N_23634,N_23424);
nand U23785 (N_23785,N_23401,N_23550);
xor U23786 (N_23786,N_23474,N_23482);
nand U23787 (N_23787,N_23617,N_23419);
and U23788 (N_23788,N_23640,N_23519);
xor U23789 (N_23789,N_23536,N_23650);
nand U23790 (N_23790,N_23568,N_23507);
xor U23791 (N_23791,N_23537,N_23462);
nor U23792 (N_23792,N_23679,N_23618);
and U23793 (N_23793,N_23654,N_23561);
or U23794 (N_23794,N_23673,N_23692);
or U23795 (N_23795,N_23429,N_23683);
and U23796 (N_23796,N_23455,N_23483);
or U23797 (N_23797,N_23410,N_23684);
or U23798 (N_23798,N_23478,N_23605);
xnor U23799 (N_23799,N_23408,N_23468);
or U23800 (N_23800,N_23676,N_23542);
or U23801 (N_23801,N_23484,N_23452);
xnor U23802 (N_23802,N_23651,N_23529);
xnor U23803 (N_23803,N_23557,N_23667);
xnor U23804 (N_23804,N_23641,N_23636);
nand U23805 (N_23805,N_23597,N_23589);
xnor U23806 (N_23806,N_23416,N_23672);
or U23807 (N_23807,N_23439,N_23463);
nor U23808 (N_23808,N_23595,N_23459);
xor U23809 (N_23809,N_23481,N_23584);
and U23810 (N_23810,N_23403,N_23428);
nand U23811 (N_23811,N_23514,N_23615);
nor U23812 (N_23812,N_23466,N_23649);
nor U23813 (N_23813,N_23551,N_23450);
nor U23814 (N_23814,N_23471,N_23552);
and U23815 (N_23815,N_23404,N_23616);
nor U23816 (N_23816,N_23454,N_23549);
xnor U23817 (N_23817,N_23414,N_23500);
nor U23818 (N_23818,N_23590,N_23583);
and U23819 (N_23819,N_23613,N_23494);
xnor U23820 (N_23820,N_23423,N_23608);
and U23821 (N_23821,N_23554,N_23562);
nor U23822 (N_23822,N_23515,N_23548);
and U23823 (N_23823,N_23630,N_23582);
or U23824 (N_23824,N_23578,N_23588);
and U23825 (N_23825,N_23570,N_23571);
or U23826 (N_23826,N_23555,N_23444);
and U23827 (N_23827,N_23567,N_23525);
and U23828 (N_23828,N_23449,N_23602);
and U23829 (N_23829,N_23440,N_23521);
and U23830 (N_23830,N_23696,N_23644);
and U23831 (N_23831,N_23681,N_23431);
nand U23832 (N_23832,N_23503,N_23585);
and U23833 (N_23833,N_23638,N_23560);
or U23834 (N_23834,N_23470,N_23620);
nand U23835 (N_23835,N_23436,N_23460);
xnor U23836 (N_23836,N_23680,N_23526);
nor U23837 (N_23837,N_23534,N_23576);
nand U23838 (N_23838,N_23635,N_23603);
or U23839 (N_23839,N_23577,N_23566);
nand U23840 (N_23840,N_23477,N_23553);
or U23841 (N_23841,N_23538,N_23418);
nor U23842 (N_23842,N_23619,N_23688);
and U23843 (N_23843,N_23573,N_23448);
and U23844 (N_23844,N_23425,N_23430);
and U23845 (N_23845,N_23524,N_23604);
nor U23846 (N_23846,N_23469,N_23443);
xnor U23847 (N_23847,N_23600,N_23502);
nand U23848 (N_23848,N_23491,N_23646);
nor U23849 (N_23849,N_23594,N_23543);
xnor U23850 (N_23850,N_23669,N_23510);
and U23851 (N_23851,N_23665,N_23678);
nor U23852 (N_23852,N_23610,N_23516);
nor U23853 (N_23853,N_23687,N_23415);
or U23854 (N_23854,N_23571,N_23622);
nor U23855 (N_23855,N_23572,N_23688);
and U23856 (N_23856,N_23518,N_23692);
nor U23857 (N_23857,N_23641,N_23629);
and U23858 (N_23858,N_23568,N_23574);
xor U23859 (N_23859,N_23665,N_23441);
xnor U23860 (N_23860,N_23558,N_23626);
or U23861 (N_23861,N_23414,N_23553);
or U23862 (N_23862,N_23683,N_23576);
xor U23863 (N_23863,N_23421,N_23529);
nor U23864 (N_23864,N_23683,N_23619);
xnor U23865 (N_23865,N_23635,N_23494);
xor U23866 (N_23866,N_23545,N_23517);
and U23867 (N_23867,N_23618,N_23649);
or U23868 (N_23868,N_23571,N_23482);
nor U23869 (N_23869,N_23548,N_23487);
nor U23870 (N_23870,N_23632,N_23687);
nand U23871 (N_23871,N_23469,N_23625);
xnor U23872 (N_23872,N_23421,N_23412);
nor U23873 (N_23873,N_23595,N_23587);
and U23874 (N_23874,N_23476,N_23490);
nand U23875 (N_23875,N_23695,N_23527);
or U23876 (N_23876,N_23415,N_23464);
and U23877 (N_23877,N_23501,N_23675);
and U23878 (N_23878,N_23676,N_23550);
xnor U23879 (N_23879,N_23517,N_23500);
or U23880 (N_23880,N_23506,N_23662);
xnor U23881 (N_23881,N_23616,N_23524);
nor U23882 (N_23882,N_23620,N_23409);
nand U23883 (N_23883,N_23483,N_23481);
and U23884 (N_23884,N_23472,N_23620);
xnor U23885 (N_23885,N_23647,N_23694);
and U23886 (N_23886,N_23650,N_23410);
nand U23887 (N_23887,N_23589,N_23529);
nand U23888 (N_23888,N_23455,N_23479);
nor U23889 (N_23889,N_23507,N_23496);
xor U23890 (N_23890,N_23446,N_23469);
and U23891 (N_23891,N_23523,N_23452);
and U23892 (N_23892,N_23557,N_23555);
and U23893 (N_23893,N_23637,N_23659);
or U23894 (N_23894,N_23484,N_23428);
or U23895 (N_23895,N_23563,N_23656);
xnor U23896 (N_23896,N_23429,N_23695);
nand U23897 (N_23897,N_23484,N_23582);
xor U23898 (N_23898,N_23522,N_23492);
xor U23899 (N_23899,N_23449,N_23442);
nand U23900 (N_23900,N_23514,N_23439);
xor U23901 (N_23901,N_23652,N_23445);
nand U23902 (N_23902,N_23670,N_23589);
xor U23903 (N_23903,N_23651,N_23693);
nand U23904 (N_23904,N_23408,N_23556);
nor U23905 (N_23905,N_23695,N_23520);
nand U23906 (N_23906,N_23436,N_23608);
nand U23907 (N_23907,N_23564,N_23618);
or U23908 (N_23908,N_23576,N_23626);
and U23909 (N_23909,N_23554,N_23465);
xnor U23910 (N_23910,N_23522,N_23484);
and U23911 (N_23911,N_23620,N_23418);
xnor U23912 (N_23912,N_23560,N_23429);
xnor U23913 (N_23913,N_23478,N_23416);
nor U23914 (N_23914,N_23640,N_23574);
xnor U23915 (N_23915,N_23559,N_23486);
nor U23916 (N_23916,N_23669,N_23591);
nand U23917 (N_23917,N_23582,N_23471);
nand U23918 (N_23918,N_23582,N_23460);
nor U23919 (N_23919,N_23688,N_23556);
and U23920 (N_23920,N_23619,N_23477);
and U23921 (N_23921,N_23645,N_23534);
nor U23922 (N_23922,N_23554,N_23462);
nor U23923 (N_23923,N_23670,N_23616);
or U23924 (N_23924,N_23580,N_23678);
xnor U23925 (N_23925,N_23653,N_23681);
nand U23926 (N_23926,N_23520,N_23550);
nand U23927 (N_23927,N_23560,N_23472);
nor U23928 (N_23928,N_23566,N_23475);
or U23929 (N_23929,N_23613,N_23473);
nand U23930 (N_23930,N_23562,N_23439);
or U23931 (N_23931,N_23626,N_23620);
nand U23932 (N_23932,N_23485,N_23513);
xnor U23933 (N_23933,N_23471,N_23571);
nand U23934 (N_23934,N_23575,N_23548);
nand U23935 (N_23935,N_23585,N_23574);
nor U23936 (N_23936,N_23579,N_23510);
or U23937 (N_23937,N_23610,N_23596);
xnor U23938 (N_23938,N_23524,N_23577);
nor U23939 (N_23939,N_23698,N_23663);
or U23940 (N_23940,N_23461,N_23664);
or U23941 (N_23941,N_23517,N_23597);
and U23942 (N_23942,N_23534,N_23697);
or U23943 (N_23943,N_23427,N_23440);
xor U23944 (N_23944,N_23521,N_23460);
nor U23945 (N_23945,N_23641,N_23597);
nand U23946 (N_23946,N_23477,N_23618);
nor U23947 (N_23947,N_23411,N_23584);
nand U23948 (N_23948,N_23525,N_23680);
nor U23949 (N_23949,N_23681,N_23437);
nand U23950 (N_23950,N_23425,N_23441);
nor U23951 (N_23951,N_23675,N_23536);
nand U23952 (N_23952,N_23659,N_23684);
nor U23953 (N_23953,N_23484,N_23488);
nand U23954 (N_23954,N_23477,N_23411);
nor U23955 (N_23955,N_23543,N_23642);
xnor U23956 (N_23956,N_23675,N_23453);
xnor U23957 (N_23957,N_23574,N_23686);
nor U23958 (N_23958,N_23548,N_23674);
or U23959 (N_23959,N_23519,N_23597);
xnor U23960 (N_23960,N_23560,N_23483);
or U23961 (N_23961,N_23452,N_23529);
or U23962 (N_23962,N_23682,N_23581);
xor U23963 (N_23963,N_23617,N_23548);
nand U23964 (N_23964,N_23506,N_23529);
or U23965 (N_23965,N_23436,N_23676);
nor U23966 (N_23966,N_23605,N_23655);
xnor U23967 (N_23967,N_23426,N_23638);
xnor U23968 (N_23968,N_23672,N_23555);
xnor U23969 (N_23969,N_23519,N_23560);
or U23970 (N_23970,N_23554,N_23524);
nand U23971 (N_23971,N_23443,N_23619);
nand U23972 (N_23972,N_23482,N_23699);
nor U23973 (N_23973,N_23636,N_23673);
or U23974 (N_23974,N_23511,N_23670);
and U23975 (N_23975,N_23569,N_23539);
xnor U23976 (N_23976,N_23499,N_23565);
nand U23977 (N_23977,N_23411,N_23550);
and U23978 (N_23978,N_23506,N_23695);
and U23979 (N_23979,N_23458,N_23596);
nand U23980 (N_23980,N_23446,N_23618);
and U23981 (N_23981,N_23588,N_23553);
or U23982 (N_23982,N_23570,N_23569);
xor U23983 (N_23983,N_23458,N_23649);
and U23984 (N_23984,N_23523,N_23521);
nor U23985 (N_23985,N_23497,N_23615);
nor U23986 (N_23986,N_23473,N_23447);
or U23987 (N_23987,N_23546,N_23414);
nand U23988 (N_23988,N_23405,N_23476);
xor U23989 (N_23989,N_23667,N_23692);
or U23990 (N_23990,N_23526,N_23539);
or U23991 (N_23991,N_23679,N_23581);
nor U23992 (N_23992,N_23637,N_23481);
nor U23993 (N_23993,N_23529,N_23616);
or U23994 (N_23994,N_23558,N_23484);
nand U23995 (N_23995,N_23675,N_23586);
nor U23996 (N_23996,N_23613,N_23475);
or U23997 (N_23997,N_23544,N_23611);
or U23998 (N_23998,N_23514,N_23481);
or U23999 (N_23999,N_23522,N_23670);
xnor U24000 (N_24000,N_23867,N_23737);
nor U24001 (N_24001,N_23870,N_23825);
nor U24002 (N_24002,N_23700,N_23952);
xnor U24003 (N_24003,N_23876,N_23794);
nand U24004 (N_24004,N_23832,N_23959);
nor U24005 (N_24005,N_23824,N_23845);
xor U24006 (N_24006,N_23759,N_23838);
xnor U24007 (N_24007,N_23793,N_23914);
and U24008 (N_24008,N_23815,N_23963);
xnor U24009 (N_24009,N_23816,N_23743);
nand U24010 (N_24010,N_23835,N_23813);
nand U24011 (N_24011,N_23976,N_23984);
nand U24012 (N_24012,N_23930,N_23970);
and U24013 (N_24013,N_23853,N_23884);
nor U24014 (N_24014,N_23846,N_23830);
or U24015 (N_24015,N_23782,N_23885);
nand U24016 (N_24016,N_23804,N_23950);
nand U24017 (N_24017,N_23858,N_23701);
xnor U24018 (N_24018,N_23968,N_23757);
xor U24019 (N_24019,N_23752,N_23738);
nor U24020 (N_24020,N_23863,N_23818);
and U24021 (N_24021,N_23716,N_23965);
or U24022 (N_24022,N_23948,N_23979);
or U24023 (N_24023,N_23719,N_23921);
and U24024 (N_24024,N_23896,N_23864);
nor U24025 (N_24025,N_23801,N_23826);
xnor U24026 (N_24026,N_23947,N_23722);
xnor U24027 (N_24027,N_23990,N_23988);
xnor U24028 (N_24028,N_23917,N_23809);
nor U24029 (N_24029,N_23873,N_23758);
xor U24030 (N_24030,N_23931,N_23842);
and U24031 (N_24031,N_23820,N_23903);
nand U24032 (N_24032,N_23945,N_23836);
and U24033 (N_24033,N_23895,N_23861);
xor U24034 (N_24034,N_23791,N_23848);
and U24035 (N_24035,N_23927,N_23956);
and U24036 (N_24036,N_23989,N_23953);
nor U24037 (N_24037,N_23754,N_23872);
xor U24038 (N_24038,N_23773,N_23975);
nor U24039 (N_24039,N_23933,N_23760);
nand U24040 (N_24040,N_23805,N_23742);
nor U24041 (N_24041,N_23783,N_23784);
and U24042 (N_24042,N_23750,N_23941);
or U24043 (N_24043,N_23899,N_23866);
and U24044 (N_24044,N_23960,N_23871);
nand U24045 (N_24045,N_23922,N_23943);
and U24046 (N_24046,N_23869,N_23912);
or U24047 (N_24047,N_23763,N_23995);
or U24048 (N_24048,N_23958,N_23734);
and U24049 (N_24049,N_23751,N_23781);
and U24050 (N_24050,N_23907,N_23799);
xnor U24051 (N_24051,N_23882,N_23982);
nand U24052 (N_24052,N_23854,N_23800);
and U24053 (N_24053,N_23755,N_23810);
nor U24054 (N_24054,N_23712,N_23926);
or U24055 (N_24055,N_23859,N_23807);
xor U24056 (N_24056,N_23875,N_23881);
nor U24057 (N_24057,N_23954,N_23851);
and U24058 (N_24058,N_23778,N_23776);
and U24059 (N_24059,N_23802,N_23906);
and U24060 (N_24060,N_23987,N_23844);
and U24061 (N_24061,N_23797,N_23822);
and U24062 (N_24062,N_23779,N_23736);
and U24063 (N_24063,N_23724,N_23991);
or U24064 (N_24064,N_23708,N_23983);
or U24065 (N_24065,N_23792,N_23957);
or U24066 (N_24066,N_23944,N_23973);
or U24067 (N_24067,N_23887,N_23936);
or U24068 (N_24068,N_23862,N_23946);
or U24069 (N_24069,N_23901,N_23744);
xor U24070 (N_24070,N_23980,N_23705);
nand U24071 (N_24071,N_23834,N_23811);
nand U24072 (N_24072,N_23741,N_23924);
nor U24073 (N_24073,N_23981,N_23932);
nand U24074 (N_24074,N_23715,N_23839);
and U24075 (N_24075,N_23874,N_23942);
or U24076 (N_24076,N_23790,N_23929);
nor U24077 (N_24077,N_23711,N_23729);
nand U24078 (N_24078,N_23771,N_23904);
nor U24079 (N_24079,N_23819,N_23774);
xnor U24080 (N_24080,N_23770,N_23923);
xnor U24081 (N_24081,N_23827,N_23749);
xor U24082 (N_24082,N_23764,N_23748);
xor U24083 (N_24083,N_23798,N_23812);
nor U24084 (N_24084,N_23786,N_23886);
or U24085 (N_24085,N_23706,N_23949);
nand U24086 (N_24086,N_23717,N_23919);
nand U24087 (N_24087,N_23891,N_23937);
and U24088 (N_24088,N_23785,N_23967);
xnor U24089 (N_24089,N_23803,N_23964);
xor U24090 (N_24090,N_23894,N_23787);
or U24091 (N_24091,N_23893,N_23928);
nand U24092 (N_24092,N_23994,N_23880);
or U24093 (N_24093,N_23777,N_23765);
or U24094 (N_24094,N_23993,N_23814);
and U24095 (N_24095,N_23726,N_23746);
xnor U24096 (N_24096,N_23780,N_23739);
or U24097 (N_24097,N_23828,N_23986);
nand U24098 (N_24098,N_23940,N_23732);
xor U24099 (N_24099,N_23740,N_23938);
or U24100 (N_24100,N_23902,N_23974);
xor U24101 (N_24101,N_23837,N_23865);
or U24102 (N_24102,N_23769,N_23951);
or U24103 (N_24103,N_23977,N_23728);
or U24104 (N_24104,N_23911,N_23788);
or U24105 (N_24105,N_23996,N_23998);
and U24106 (N_24106,N_23868,N_23879);
and U24107 (N_24107,N_23761,N_23731);
nand U24108 (N_24108,N_23910,N_23889);
or U24109 (N_24109,N_23892,N_23733);
or U24110 (N_24110,N_23898,N_23829);
and U24111 (N_24111,N_23841,N_23878);
nor U24112 (N_24112,N_23908,N_23969);
xnor U24113 (N_24113,N_23745,N_23897);
and U24114 (N_24114,N_23847,N_23999);
or U24115 (N_24115,N_23916,N_23720);
and U24116 (N_24116,N_23843,N_23756);
nand U24117 (N_24117,N_23714,N_23703);
xnor U24118 (N_24118,N_23935,N_23702);
nor U24119 (N_24119,N_23796,N_23730);
and U24120 (N_24120,N_23850,N_23962);
and U24121 (N_24121,N_23747,N_23831);
xnor U24122 (N_24122,N_23707,N_23849);
xnor U24123 (N_24123,N_23860,N_23789);
nor U24124 (N_24124,N_23900,N_23709);
or U24125 (N_24125,N_23909,N_23877);
nand U24126 (N_24126,N_23925,N_23762);
xnor U24127 (N_24127,N_23710,N_23767);
nand U24128 (N_24128,N_23883,N_23723);
nand U24129 (N_24129,N_23753,N_23735);
and U24130 (N_24130,N_23725,N_23972);
nor U24131 (N_24131,N_23817,N_23704);
nand U24132 (N_24132,N_23939,N_23718);
or U24133 (N_24133,N_23721,N_23833);
nand U24134 (N_24134,N_23775,N_23823);
nand U24135 (N_24135,N_23855,N_23985);
nand U24136 (N_24136,N_23992,N_23966);
or U24137 (N_24137,N_23971,N_23713);
nor U24138 (N_24138,N_23852,N_23913);
nand U24139 (N_24139,N_23888,N_23856);
nand U24140 (N_24140,N_23961,N_23905);
nand U24141 (N_24141,N_23955,N_23920);
nor U24142 (N_24142,N_23918,N_23795);
or U24143 (N_24143,N_23772,N_23890);
xor U24144 (N_24144,N_23978,N_23808);
and U24145 (N_24145,N_23934,N_23821);
nor U24146 (N_24146,N_23997,N_23915);
or U24147 (N_24147,N_23766,N_23857);
nor U24148 (N_24148,N_23727,N_23840);
or U24149 (N_24149,N_23806,N_23768);
nor U24150 (N_24150,N_23728,N_23793);
and U24151 (N_24151,N_23976,N_23893);
xnor U24152 (N_24152,N_23915,N_23861);
nand U24153 (N_24153,N_23836,N_23727);
xor U24154 (N_24154,N_23713,N_23756);
xnor U24155 (N_24155,N_23732,N_23969);
or U24156 (N_24156,N_23991,N_23855);
xor U24157 (N_24157,N_23747,N_23974);
xnor U24158 (N_24158,N_23744,N_23731);
and U24159 (N_24159,N_23899,N_23952);
xor U24160 (N_24160,N_23860,N_23839);
and U24161 (N_24161,N_23826,N_23961);
xor U24162 (N_24162,N_23713,N_23926);
and U24163 (N_24163,N_23730,N_23812);
and U24164 (N_24164,N_23903,N_23854);
and U24165 (N_24165,N_23800,N_23770);
or U24166 (N_24166,N_23753,N_23860);
and U24167 (N_24167,N_23925,N_23944);
and U24168 (N_24168,N_23807,N_23758);
nand U24169 (N_24169,N_23968,N_23822);
nand U24170 (N_24170,N_23842,N_23995);
xnor U24171 (N_24171,N_23958,N_23972);
xnor U24172 (N_24172,N_23976,N_23862);
nand U24173 (N_24173,N_23985,N_23718);
or U24174 (N_24174,N_23988,N_23931);
or U24175 (N_24175,N_23882,N_23714);
or U24176 (N_24176,N_23884,N_23922);
and U24177 (N_24177,N_23865,N_23948);
nand U24178 (N_24178,N_23876,N_23917);
xor U24179 (N_24179,N_23853,N_23721);
or U24180 (N_24180,N_23701,N_23714);
xnor U24181 (N_24181,N_23888,N_23769);
nand U24182 (N_24182,N_23735,N_23962);
nor U24183 (N_24183,N_23812,N_23959);
nor U24184 (N_24184,N_23729,N_23861);
xor U24185 (N_24185,N_23709,N_23933);
or U24186 (N_24186,N_23875,N_23786);
xnor U24187 (N_24187,N_23769,N_23918);
xnor U24188 (N_24188,N_23731,N_23953);
xnor U24189 (N_24189,N_23863,N_23839);
nand U24190 (N_24190,N_23923,N_23727);
nand U24191 (N_24191,N_23912,N_23722);
xnor U24192 (N_24192,N_23929,N_23878);
or U24193 (N_24193,N_23762,N_23719);
or U24194 (N_24194,N_23714,N_23888);
xor U24195 (N_24195,N_23944,N_23954);
xnor U24196 (N_24196,N_23883,N_23726);
nor U24197 (N_24197,N_23825,N_23700);
or U24198 (N_24198,N_23894,N_23760);
nor U24199 (N_24199,N_23973,N_23775);
or U24200 (N_24200,N_23987,N_23874);
nor U24201 (N_24201,N_23996,N_23815);
or U24202 (N_24202,N_23797,N_23868);
or U24203 (N_24203,N_23709,N_23772);
and U24204 (N_24204,N_23865,N_23955);
nand U24205 (N_24205,N_23985,N_23779);
or U24206 (N_24206,N_23739,N_23784);
and U24207 (N_24207,N_23806,N_23794);
xor U24208 (N_24208,N_23865,N_23780);
and U24209 (N_24209,N_23883,N_23914);
nand U24210 (N_24210,N_23994,N_23762);
xor U24211 (N_24211,N_23701,N_23976);
xor U24212 (N_24212,N_23941,N_23848);
xor U24213 (N_24213,N_23704,N_23766);
nand U24214 (N_24214,N_23828,N_23834);
nand U24215 (N_24215,N_23702,N_23776);
or U24216 (N_24216,N_23716,N_23911);
nor U24217 (N_24217,N_23914,N_23821);
nand U24218 (N_24218,N_23822,N_23912);
xnor U24219 (N_24219,N_23743,N_23944);
and U24220 (N_24220,N_23894,N_23972);
or U24221 (N_24221,N_23761,N_23790);
nand U24222 (N_24222,N_23752,N_23733);
xor U24223 (N_24223,N_23887,N_23992);
nand U24224 (N_24224,N_23855,N_23786);
and U24225 (N_24225,N_23706,N_23885);
or U24226 (N_24226,N_23719,N_23892);
or U24227 (N_24227,N_23810,N_23831);
and U24228 (N_24228,N_23952,N_23794);
and U24229 (N_24229,N_23755,N_23933);
or U24230 (N_24230,N_23823,N_23900);
nor U24231 (N_24231,N_23857,N_23939);
nand U24232 (N_24232,N_23838,N_23827);
nand U24233 (N_24233,N_23703,N_23796);
nor U24234 (N_24234,N_23769,N_23826);
nor U24235 (N_24235,N_23843,N_23812);
and U24236 (N_24236,N_23903,N_23763);
nor U24237 (N_24237,N_23762,N_23845);
xnor U24238 (N_24238,N_23867,N_23852);
and U24239 (N_24239,N_23926,N_23929);
and U24240 (N_24240,N_23797,N_23789);
nand U24241 (N_24241,N_23804,N_23853);
xor U24242 (N_24242,N_23795,N_23728);
and U24243 (N_24243,N_23758,N_23838);
and U24244 (N_24244,N_23926,N_23817);
and U24245 (N_24245,N_23854,N_23838);
or U24246 (N_24246,N_23981,N_23761);
nor U24247 (N_24247,N_23906,N_23726);
and U24248 (N_24248,N_23984,N_23804);
xor U24249 (N_24249,N_23810,N_23944);
and U24250 (N_24250,N_23921,N_23908);
and U24251 (N_24251,N_23779,N_23853);
xnor U24252 (N_24252,N_23918,N_23777);
and U24253 (N_24253,N_23722,N_23944);
and U24254 (N_24254,N_23929,N_23784);
or U24255 (N_24255,N_23798,N_23854);
nand U24256 (N_24256,N_23953,N_23794);
nor U24257 (N_24257,N_23743,N_23926);
or U24258 (N_24258,N_23828,N_23892);
nand U24259 (N_24259,N_23743,N_23714);
or U24260 (N_24260,N_23977,N_23881);
or U24261 (N_24261,N_23784,N_23838);
xnor U24262 (N_24262,N_23899,N_23712);
nor U24263 (N_24263,N_23767,N_23786);
nand U24264 (N_24264,N_23958,N_23967);
nor U24265 (N_24265,N_23813,N_23767);
or U24266 (N_24266,N_23788,N_23916);
nor U24267 (N_24267,N_23896,N_23984);
and U24268 (N_24268,N_23847,N_23712);
xnor U24269 (N_24269,N_23875,N_23972);
xnor U24270 (N_24270,N_23773,N_23861);
and U24271 (N_24271,N_23730,N_23928);
and U24272 (N_24272,N_23977,N_23763);
xnor U24273 (N_24273,N_23959,N_23728);
nor U24274 (N_24274,N_23993,N_23931);
nand U24275 (N_24275,N_23969,N_23859);
xnor U24276 (N_24276,N_23804,N_23813);
and U24277 (N_24277,N_23781,N_23808);
and U24278 (N_24278,N_23748,N_23869);
xnor U24279 (N_24279,N_23911,N_23754);
nand U24280 (N_24280,N_23903,N_23725);
xor U24281 (N_24281,N_23934,N_23719);
nor U24282 (N_24282,N_23776,N_23947);
nor U24283 (N_24283,N_23949,N_23998);
or U24284 (N_24284,N_23857,N_23762);
and U24285 (N_24285,N_23909,N_23707);
or U24286 (N_24286,N_23896,N_23791);
or U24287 (N_24287,N_23956,N_23971);
nand U24288 (N_24288,N_23941,N_23824);
and U24289 (N_24289,N_23959,N_23740);
or U24290 (N_24290,N_23935,N_23915);
nor U24291 (N_24291,N_23709,N_23813);
xor U24292 (N_24292,N_23755,N_23738);
xnor U24293 (N_24293,N_23735,N_23786);
or U24294 (N_24294,N_23815,N_23983);
and U24295 (N_24295,N_23768,N_23830);
or U24296 (N_24296,N_23715,N_23729);
nand U24297 (N_24297,N_23814,N_23706);
xor U24298 (N_24298,N_23759,N_23721);
nand U24299 (N_24299,N_23847,N_23813);
nand U24300 (N_24300,N_24178,N_24180);
nor U24301 (N_24301,N_24086,N_24185);
or U24302 (N_24302,N_24111,N_24192);
xnor U24303 (N_24303,N_24075,N_24044);
nor U24304 (N_24304,N_24288,N_24295);
nor U24305 (N_24305,N_24233,N_24214);
xor U24306 (N_24306,N_24070,N_24018);
or U24307 (N_24307,N_24121,N_24208);
and U24308 (N_24308,N_24087,N_24104);
or U24309 (N_24309,N_24110,N_24289);
nor U24310 (N_24310,N_24274,N_24097);
nand U24311 (N_24311,N_24265,N_24167);
or U24312 (N_24312,N_24098,N_24168);
nand U24313 (N_24313,N_24221,N_24241);
xor U24314 (N_24314,N_24029,N_24009);
nand U24315 (N_24315,N_24278,N_24023);
and U24316 (N_24316,N_24002,N_24232);
nor U24317 (N_24317,N_24024,N_24034);
nand U24318 (N_24318,N_24027,N_24131);
and U24319 (N_24319,N_24112,N_24188);
and U24320 (N_24320,N_24197,N_24299);
xnor U24321 (N_24321,N_24291,N_24127);
or U24322 (N_24322,N_24234,N_24176);
and U24323 (N_24323,N_24281,N_24043);
and U24324 (N_24324,N_24275,N_24133);
nand U24325 (N_24325,N_24063,N_24230);
nor U24326 (N_24326,N_24277,N_24280);
nand U24327 (N_24327,N_24038,N_24079);
and U24328 (N_24328,N_24139,N_24041);
xnor U24329 (N_24329,N_24003,N_24088);
nor U24330 (N_24330,N_24271,N_24285);
nor U24331 (N_24331,N_24227,N_24153);
nor U24332 (N_24332,N_24217,N_24200);
nor U24333 (N_24333,N_24261,N_24037);
and U24334 (N_24334,N_24036,N_24284);
nor U24335 (N_24335,N_24297,N_24251);
nand U24336 (N_24336,N_24219,N_24216);
or U24337 (N_24337,N_24117,N_24055);
nor U24338 (N_24338,N_24235,N_24160);
nand U24339 (N_24339,N_24021,N_24116);
xor U24340 (N_24340,N_24129,N_24262);
nor U24341 (N_24341,N_24165,N_24078);
or U24342 (N_24342,N_24052,N_24199);
and U24343 (N_24343,N_24132,N_24172);
or U24344 (N_24344,N_24174,N_24266);
xor U24345 (N_24345,N_24187,N_24193);
and U24346 (N_24346,N_24205,N_24220);
nor U24347 (N_24347,N_24267,N_24206);
or U24348 (N_24348,N_24015,N_24296);
and U24349 (N_24349,N_24294,N_24026);
nand U24350 (N_24350,N_24067,N_24103);
xnor U24351 (N_24351,N_24049,N_24290);
xor U24352 (N_24352,N_24010,N_24115);
or U24353 (N_24353,N_24231,N_24081);
or U24354 (N_24354,N_24091,N_24105);
and U24355 (N_24355,N_24239,N_24181);
or U24356 (N_24356,N_24244,N_24158);
or U24357 (N_24357,N_24102,N_24073);
xnor U24358 (N_24358,N_24173,N_24004);
and U24359 (N_24359,N_24286,N_24046);
or U24360 (N_24360,N_24171,N_24006);
or U24361 (N_24361,N_24005,N_24229);
xnor U24362 (N_24362,N_24000,N_24066);
and U24363 (N_24363,N_24106,N_24142);
or U24364 (N_24364,N_24039,N_24215);
or U24365 (N_24365,N_24226,N_24146);
or U24366 (N_24366,N_24014,N_24162);
xnor U24367 (N_24367,N_24134,N_24077);
nand U24368 (N_24368,N_24136,N_24090);
and U24369 (N_24369,N_24012,N_24202);
nand U24370 (N_24370,N_24019,N_24238);
nand U24371 (N_24371,N_24163,N_24076);
or U24372 (N_24372,N_24186,N_24025);
or U24373 (N_24373,N_24224,N_24258);
and U24374 (N_24374,N_24061,N_24085);
nor U24375 (N_24375,N_24054,N_24155);
and U24376 (N_24376,N_24152,N_24082);
nor U24377 (N_24377,N_24222,N_24028);
or U24378 (N_24378,N_24084,N_24175);
or U24379 (N_24379,N_24236,N_24184);
nor U24380 (N_24380,N_24279,N_24138);
nor U24381 (N_24381,N_24189,N_24298);
nand U24382 (N_24382,N_24096,N_24237);
and U24383 (N_24383,N_24196,N_24292);
or U24384 (N_24384,N_24264,N_24101);
or U24385 (N_24385,N_24245,N_24218);
or U24386 (N_24386,N_24100,N_24156);
xor U24387 (N_24387,N_24068,N_24246);
xor U24388 (N_24388,N_24157,N_24268);
xor U24389 (N_24389,N_24114,N_24151);
and U24390 (N_24390,N_24256,N_24001);
or U24391 (N_24391,N_24113,N_24056);
nor U24392 (N_24392,N_24249,N_24169);
and U24393 (N_24393,N_24161,N_24283);
nand U24394 (N_24394,N_24272,N_24276);
nand U24395 (N_24395,N_24240,N_24195);
nand U24396 (N_24396,N_24053,N_24016);
nor U24397 (N_24397,N_24017,N_24223);
nor U24398 (N_24398,N_24270,N_24047);
nand U24399 (N_24399,N_24108,N_24089);
xnor U24400 (N_24400,N_24095,N_24164);
xor U24401 (N_24401,N_24040,N_24145);
or U24402 (N_24402,N_24190,N_24159);
nor U24403 (N_24403,N_24191,N_24020);
xnor U24404 (N_24404,N_24254,N_24248);
nor U24405 (N_24405,N_24059,N_24042);
or U24406 (N_24406,N_24048,N_24069);
nand U24407 (N_24407,N_24045,N_24060);
or U24408 (N_24408,N_24260,N_24094);
or U24409 (N_24409,N_24148,N_24064);
xnor U24410 (N_24410,N_24282,N_24119);
and U24411 (N_24411,N_24140,N_24250);
nor U24412 (N_24412,N_24109,N_24032);
nand U24413 (N_24413,N_24050,N_24135);
nand U24414 (N_24414,N_24144,N_24074);
nand U24415 (N_24415,N_24255,N_24124);
and U24416 (N_24416,N_24072,N_24123);
nor U24417 (N_24417,N_24243,N_24125);
nand U24418 (N_24418,N_24213,N_24011);
nor U24419 (N_24419,N_24122,N_24263);
or U24420 (N_24420,N_24253,N_24259);
or U24421 (N_24421,N_24198,N_24225);
or U24422 (N_24422,N_24071,N_24211);
or U24423 (N_24423,N_24143,N_24033);
nor U24424 (N_24424,N_24183,N_24273);
or U24425 (N_24425,N_24008,N_24257);
and U24426 (N_24426,N_24154,N_24201);
and U24427 (N_24427,N_24062,N_24141);
xor U24428 (N_24428,N_24057,N_24099);
xor U24429 (N_24429,N_24182,N_24242);
or U24430 (N_24430,N_24126,N_24228);
and U24431 (N_24431,N_24287,N_24130);
nor U24432 (N_24432,N_24212,N_24210);
and U24433 (N_24433,N_24058,N_24107);
nand U24434 (N_24434,N_24149,N_24092);
and U24435 (N_24435,N_24166,N_24204);
nand U24436 (N_24436,N_24150,N_24120);
nand U24437 (N_24437,N_24209,N_24252);
xor U24438 (N_24438,N_24177,N_24203);
nor U24439 (N_24439,N_24147,N_24179);
or U24440 (N_24440,N_24293,N_24007);
xor U24441 (N_24441,N_24030,N_24093);
or U24442 (N_24442,N_24035,N_24022);
nor U24443 (N_24443,N_24194,N_24118);
or U24444 (N_24444,N_24128,N_24065);
nor U24445 (N_24445,N_24247,N_24269);
and U24446 (N_24446,N_24137,N_24083);
or U24447 (N_24447,N_24013,N_24051);
nor U24448 (N_24448,N_24080,N_24031);
and U24449 (N_24449,N_24207,N_24170);
nand U24450 (N_24450,N_24219,N_24169);
and U24451 (N_24451,N_24067,N_24064);
or U24452 (N_24452,N_24154,N_24012);
nor U24453 (N_24453,N_24027,N_24240);
nand U24454 (N_24454,N_24024,N_24014);
or U24455 (N_24455,N_24138,N_24129);
or U24456 (N_24456,N_24269,N_24237);
and U24457 (N_24457,N_24161,N_24041);
nor U24458 (N_24458,N_24232,N_24030);
and U24459 (N_24459,N_24052,N_24035);
nor U24460 (N_24460,N_24177,N_24205);
nor U24461 (N_24461,N_24028,N_24293);
and U24462 (N_24462,N_24249,N_24273);
nor U24463 (N_24463,N_24295,N_24057);
xor U24464 (N_24464,N_24025,N_24252);
nor U24465 (N_24465,N_24071,N_24015);
and U24466 (N_24466,N_24043,N_24271);
nor U24467 (N_24467,N_24206,N_24112);
or U24468 (N_24468,N_24209,N_24118);
nand U24469 (N_24469,N_24101,N_24141);
xnor U24470 (N_24470,N_24197,N_24151);
and U24471 (N_24471,N_24001,N_24061);
nor U24472 (N_24472,N_24131,N_24229);
nand U24473 (N_24473,N_24175,N_24249);
nand U24474 (N_24474,N_24187,N_24132);
xor U24475 (N_24475,N_24298,N_24185);
nor U24476 (N_24476,N_24292,N_24217);
nor U24477 (N_24477,N_24163,N_24121);
xor U24478 (N_24478,N_24239,N_24068);
or U24479 (N_24479,N_24176,N_24172);
xnor U24480 (N_24480,N_24292,N_24083);
and U24481 (N_24481,N_24151,N_24142);
xnor U24482 (N_24482,N_24286,N_24180);
nand U24483 (N_24483,N_24105,N_24063);
nor U24484 (N_24484,N_24143,N_24266);
or U24485 (N_24485,N_24184,N_24282);
nor U24486 (N_24486,N_24116,N_24260);
xnor U24487 (N_24487,N_24239,N_24238);
and U24488 (N_24488,N_24078,N_24143);
nor U24489 (N_24489,N_24269,N_24210);
nor U24490 (N_24490,N_24059,N_24095);
nor U24491 (N_24491,N_24105,N_24212);
and U24492 (N_24492,N_24146,N_24133);
and U24493 (N_24493,N_24151,N_24106);
nand U24494 (N_24494,N_24107,N_24096);
and U24495 (N_24495,N_24282,N_24209);
nor U24496 (N_24496,N_24094,N_24150);
and U24497 (N_24497,N_24275,N_24038);
nor U24498 (N_24498,N_24236,N_24125);
xnor U24499 (N_24499,N_24025,N_24271);
nand U24500 (N_24500,N_24231,N_24227);
or U24501 (N_24501,N_24128,N_24221);
xnor U24502 (N_24502,N_24162,N_24026);
nor U24503 (N_24503,N_24059,N_24050);
nand U24504 (N_24504,N_24294,N_24212);
or U24505 (N_24505,N_24174,N_24075);
nand U24506 (N_24506,N_24203,N_24236);
xnor U24507 (N_24507,N_24071,N_24218);
or U24508 (N_24508,N_24081,N_24176);
nor U24509 (N_24509,N_24109,N_24052);
or U24510 (N_24510,N_24146,N_24256);
or U24511 (N_24511,N_24193,N_24014);
nor U24512 (N_24512,N_24168,N_24075);
xnor U24513 (N_24513,N_24126,N_24205);
xnor U24514 (N_24514,N_24157,N_24174);
or U24515 (N_24515,N_24083,N_24222);
or U24516 (N_24516,N_24181,N_24229);
xnor U24517 (N_24517,N_24101,N_24134);
xor U24518 (N_24518,N_24056,N_24065);
xor U24519 (N_24519,N_24162,N_24077);
or U24520 (N_24520,N_24070,N_24003);
xor U24521 (N_24521,N_24059,N_24118);
nand U24522 (N_24522,N_24174,N_24245);
or U24523 (N_24523,N_24291,N_24281);
nor U24524 (N_24524,N_24101,N_24015);
nor U24525 (N_24525,N_24160,N_24209);
and U24526 (N_24526,N_24011,N_24025);
xnor U24527 (N_24527,N_24285,N_24127);
or U24528 (N_24528,N_24225,N_24073);
nand U24529 (N_24529,N_24064,N_24241);
nand U24530 (N_24530,N_24278,N_24254);
nand U24531 (N_24531,N_24166,N_24192);
nand U24532 (N_24532,N_24110,N_24023);
or U24533 (N_24533,N_24007,N_24150);
or U24534 (N_24534,N_24260,N_24075);
xnor U24535 (N_24535,N_24031,N_24211);
nor U24536 (N_24536,N_24239,N_24048);
or U24537 (N_24537,N_24183,N_24185);
nor U24538 (N_24538,N_24005,N_24079);
and U24539 (N_24539,N_24273,N_24112);
and U24540 (N_24540,N_24003,N_24006);
xor U24541 (N_24541,N_24262,N_24225);
xnor U24542 (N_24542,N_24242,N_24163);
xnor U24543 (N_24543,N_24164,N_24131);
xnor U24544 (N_24544,N_24281,N_24274);
and U24545 (N_24545,N_24254,N_24291);
xnor U24546 (N_24546,N_24140,N_24097);
and U24547 (N_24547,N_24292,N_24117);
or U24548 (N_24548,N_24215,N_24150);
xor U24549 (N_24549,N_24123,N_24288);
or U24550 (N_24550,N_24139,N_24018);
xnor U24551 (N_24551,N_24084,N_24174);
and U24552 (N_24552,N_24073,N_24190);
xnor U24553 (N_24553,N_24290,N_24285);
or U24554 (N_24554,N_24253,N_24146);
nand U24555 (N_24555,N_24230,N_24103);
nor U24556 (N_24556,N_24252,N_24243);
nor U24557 (N_24557,N_24011,N_24295);
or U24558 (N_24558,N_24269,N_24020);
and U24559 (N_24559,N_24193,N_24276);
nor U24560 (N_24560,N_24099,N_24116);
or U24561 (N_24561,N_24051,N_24187);
nand U24562 (N_24562,N_24081,N_24106);
nand U24563 (N_24563,N_24157,N_24262);
or U24564 (N_24564,N_24092,N_24103);
xor U24565 (N_24565,N_24143,N_24147);
xor U24566 (N_24566,N_24270,N_24026);
or U24567 (N_24567,N_24012,N_24257);
nor U24568 (N_24568,N_24251,N_24104);
nor U24569 (N_24569,N_24268,N_24164);
nor U24570 (N_24570,N_24146,N_24004);
or U24571 (N_24571,N_24051,N_24069);
xor U24572 (N_24572,N_24004,N_24253);
or U24573 (N_24573,N_24224,N_24277);
nor U24574 (N_24574,N_24050,N_24099);
nand U24575 (N_24575,N_24197,N_24252);
and U24576 (N_24576,N_24103,N_24277);
nor U24577 (N_24577,N_24129,N_24170);
nand U24578 (N_24578,N_24027,N_24014);
or U24579 (N_24579,N_24294,N_24151);
nand U24580 (N_24580,N_24193,N_24010);
nor U24581 (N_24581,N_24227,N_24230);
and U24582 (N_24582,N_24127,N_24071);
or U24583 (N_24583,N_24059,N_24200);
xor U24584 (N_24584,N_24196,N_24034);
nand U24585 (N_24585,N_24126,N_24196);
nor U24586 (N_24586,N_24292,N_24202);
nand U24587 (N_24587,N_24218,N_24296);
nor U24588 (N_24588,N_24281,N_24127);
and U24589 (N_24589,N_24034,N_24274);
nand U24590 (N_24590,N_24018,N_24122);
and U24591 (N_24591,N_24241,N_24172);
and U24592 (N_24592,N_24114,N_24147);
nand U24593 (N_24593,N_24081,N_24057);
or U24594 (N_24594,N_24008,N_24203);
nor U24595 (N_24595,N_24131,N_24279);
nand U24596 (N_24596,N_24234,N_24204);
nand U24597 (N_24597,N_24060,N_24262);
xnor U24598 (N_24598,N_24027,N_24116);
and U24599 (N_24599,N_24207,N_24199);
and U24600 (N_24600,N_24302,N_24357);
nor U24601 (N_24601,N_24443,N_24563);
and U24602 (N_24602,N_24548,N_24348);
and U24603 (N_24603,N_24324,N_24569);
and U24604 (N_24604,N_24577,N_24430);
or U24605 (N_24605,N_24365,N_24304);
xor U24606 (N_24606,N_24527,N_24415);
xnor U24607 (N_24607,N_24383,N_24439);
xnor U24608 (N_24608,N_24580,N_24401);
and U24609 (N_24609,N_24353,N_24586);
or U24610 (N_24610,N_24411,N_24350);
or U24611 (N_24611,N_24314,N_24378);
nand U24612 (N_24612,N_24472,N_24317);
and U24613 (N_24613,N_24478,N_24465);
nor U24614 (N_24614,N_24526,N_24456);
xor U24615 (N_24615,N_24554,N_24496);
and U24616 (N_24616,N_24504,N_24308);
xor U24617 (N_24617,N_24387,N_24520);
xnor U24618 (N_24618,N_24509,N_24538);
nor U24619 (N_24619,N_24547,N_24557);
and U24620 (N_24620,N_24523,N_24426);
or U24621 (N_24621,N_24433,N_24419);
xor U24622 (N_24622,N_24326,N_24346);
nand U24623 (N_24623,N_24593,N_24559);
nor U24624 (N_24624,N_24341,N_24518);
or U24625 (N_24625,N_24381,N_24438);
nand U24626 (N_24626,N_24400,N_24440);
xnor U24627 (N_24627,N_24335,N_24514);
nand U24628 (N_24628,N_24448,N_24442);
nand U24629 (N_24629,N_24423,N_24571);
or U24630 (N_24630,N_24510,N_24333);
and U24631 (N_24631,N_24587,N_24502);
and U24632 (N_24632,N_24345,N_24379);
and U24633 (N_24633,N_24582,N_24489);
and U24634 (N_24634,N_24390,N_24359);
nand U24635 (N_24635,N_24328,N_24477);
nor U24636 (N_24636,N_24543,N_24599);
xor U24637 (N_24637,N_24474,N_24590);
nor U24638 (N_24638,N_24408,N_24418);
nor U24639 (N_24639,N_24327,N_24434);
nand U24640 (N_24640,N_24573,N_24482);
nand U24641 (N_24641,N_24392,N_24597);
nand U24642 (N_24642,N_24393,N_24503);
and U24643 (N_24643,N_24432,N_24311);
nor U24644 (N_24644,N_24331,N_24453);
nand U24645 (N_24645,N_24508,N_24513);
nor U24646 (N_24646,N_24427,N_24519);
nor U24647 (N_24647,N_24402,N_24300);
and U24648 (N_24648,N_24583,N_24309);
nand U24649 (N_24649,N_24316,N_24531);
and U24650 (N_24650,N_24494,N_24512);
and U24651 (N_24651,N_24344,N_24539);
and U24652 (N_24652,N_24540,N_24460);
nand U24653 (N_24653,N_24407,N_24528);
nor U24654 (N_24654,N_24575,N_24319);
nand U24655 (N_24655,N_24332,N_24451);
or U24656 (N_24656,N_24564,N_24445);
nand U24657 (N_24657,N_24495,N_24342);
nor U24658 (N_24658,N_24458,N_24546);
and U24659 (N_24659,N_24459,N_24461);
and U24660 (N_24660,N_24579,N_24545);
and U24661 (N_24661,N_24487,N_24506);
nor U24662 (N_24662,N_24405,N_24467);
xnor U24663 (N_24663,N_24356,N_24553);
xor U24664 (N_24664,N_24585,N_24330);
xnor U24665 (N_24665,N_24367,N_24431);
or U24666 (N_24666,N_24534,N_24382);
or U24667 (N_24667,N_24444,N_24372);
nand U24668 (N_24668,N_24364,N_24437);
xnor U24669 (N_24669,N_24322,N_24533);
xnor U24670 (N_24670,N_24463,N_24421);
nor U24671 (N_24671,N_24476,N_24549);
nor U24672 (N_24672,N_24420,N_24325);
and U24673 (N_24673,N_24428,N_24521);
nand U24674 (N_24674,N_24354,N_24339);
nor U24675 (N_24675,N_24349,N_24578);
nand U24676 (N_24676,N_24429,N_24556);
and U24677 (N_24677,N_24446,N_24522);
and U24678 (N_24678,N_24391,N_24570);
and U24679 (N_24679,N_24370,N_24306);
nand U24680 (N_24680,N_24452,N_24491);
or U24681 (N_24681,N_24576,N_24532);
nor U24682 (N_24682,N_24529,N_24410);
xnor U24683 (N_24683,N_24473,N_24455);
nor U24684 (N_24684,N_24376,N_24323);
or U24685 (N_24685,N_24441,N_24413);
or U24686 (N_24686,N_24343,N_24484);
or U24687 (N_24687,N_24574,N_24493);
xor U24688 (N_24688,N_24307,N_24581);
xor U24689 (N_24689,N_24313,N_24388);
nor U24690 (N_24690,N_24436,N_24544);
nor U24691 (N_24691,N_24337,N_24374);
or U24692 (N_24692,N_24594,N_24396);
nor U24693 (N_24693,N_24369,N_24483);
nor U24694 (N_24694,N_24479,N_24565);
nor U24695 (N_24695,N_24366,N_24454);
and U24696 (N_24696,N_24501,N_24384);
nand U24697 (N_24697,N_24417,N_24377);
or U24698 (N_24698,N_24499,N_24475);
xnor U24699 (N_24699,N_24375,N_24368);
nand U24700 (N_24700,N_24470,N_24310);
nand U24701 (N_24701,N_24535,N_24488);
xor U24702 (N_24702,N_24598,N_24462);
xnor U24703 (N_24703,N_24498,N_24315);
nand U24704 (N_24704,N_24412,N_24386);
nor U24705 (N_24705,N_24525,N_24312);
and U24706 (N_24706,N_24567,N_24360);
nor U24707 (N_24707,N_24515,N_24449);
xor U24708 (N_24708,N_24380,N_24334);
and U24709 (N_24709,N_24481,N_24406);
or U24710 (N_24710,N_24394,N_24361);
and U24711 (N_24711,N_24457,N_24537);
nor U24712 (N_24712,N_24500,N_24592);
nor U24713 (N_24713,N_24351,N_24517);
or U24714 (N_24714,N_24568,N_24358);
or U24715 (N_24715,N_24589,N_24511);
xnor U24716 (N_24716,N_24447,N_24551);
nor U24717 (N_24717,N_24424,N_24566);
or U24718 (N_24718,N_24389,N_24562);
or U24719 (N_24719,N_24558,N_24422);
and U24720 (N_24720,N_24318,N_24507);
or U24721 (N_24721,N_24320,N_24404);
or U24722 (N_24722,N_24591,N_24505);
nor U24723 (N_24723,N_24414,N_24363);
and U24724 (N_24724,N_24338,N_24530);
nor U24725 (N_24725,N_24541,N_24468);
and U24726 (N_24726,N_24403,N_24595);
and U24727 (N_24727,N_24425,N_24409);
nor U24728 (N_24728,N_24397,N_24395);
nor U24729 (N_24729,N_24555,N_24542);
and U24730 (N_24730,N_24469,N_24584);
nand U24731 (N_24731,N_24471,N_24305);
nor U24732 (N_24732,N_24486,N_24560);
nor U24733 (N_24733,N_24524,N_24588);
nand U24734 (N_24734,N_24371,N_24399);
xnor U24735 (N_24735,N_24516,N_24347);
nor U24736 (N_24736,N_24466,N_24416);
and U24737 (N_24737,N_24485,N_24373);
nand U24738 (N_24738,N_24398,N_24301);
or U24739 (N_24739,N_24464,N_24352);
or U24740 (N_24740,N_24492,N_24303);
and U24741 (N_24741,N_24552,N_24536);
and U24742 (N_24742,N_24490,N_24385);
or U24743 (N_24743,N_24450,N_24572);
or U24744 (N_24744,N_24480,N_24497);
and U24745 (N_24745,N_24321,N_24336);
nor U24746 (N_24746,N_24550,N_24596);
nand U24747 (N_24747,N_24435,N_24329);
xor U24748 (N_24748,N_24355,N_24561);
xnor U24749 (N_24749,N_24362,N_24340);
or U24750 (N_24750,N_24424,N_24540);
xor U24751 (N_24751,N_24384,N_24453);
and U24752 (N_24752,N_24361,N_24404);
or U24753 (N_24753,N_24379,N_24522);
nand U24754 (N_24754,N_24337,N_24329);
or U24755 (N_24755,N_24541,N_24478);
and U24756 (N_24756,N_24522,N_24455);
and U24757 (N_24757,N_24317,N_24405);
xor U24758 (N_24758,N_24581,N_24324);
nor U24759 (N_24759,N_24494,N_24570);
nand U24760 (N_24760,N_24599,N_24447);
and U24761 (N_24761,N_24402,N_24492);
nand U24762 (N_24762,N_24362,N_24379);
xor U24763 (N_24763,N_24500,N_24480);
or U24764 (N_24764,N_24502,N_24395);
xor U24765 (N_24765,N_24438,N_24505);
nor U24766 (N_24766,N_24324,N_24453);
xnor U24767 (N_24767,N_24429,N_24526);
nand U24768 (N_24768,N_24556,N_24583);
nor U24769 (N_24769,N_24311,N_24510);
or U24770 (N_24770,N_24374,N_24409);
or U24771 (N_24771,N_24326,N_24515);
and U24772 (N_24772,N_24497,N_24437);
nor U24773 (N_24773,N_24327,N_24552);
nor U24774 (N_24774,N_24583,N_24519);
or U24775 (N_24775,N_24302,N_24438);
or U24776 (N_24776,N_24312,N_24539);
or U24777 (N_24777,N_24553,N_24489);
and U24778 (N_24778,N_24581,N_24395);
nand U24779 (N_24779,N_24517,N_24435);
nor U24780 (N_24780,N_24549,N_24437);
nand U24781 (N_24781,N_24318,N_24518);
nor U24782 (N_24782,N_24548,N_24530);
or U24783 (N_24783,N_24548,N_24560);
and U24784 (N_24784,N_24402,N_24351);
nand U24785 (N_24785,N_24381,N_24585);
xor U24786 (N_24786,N_24582,N_24475);
nand U24787 (N_24787,N_24461,N_24486);
or U24788 (N_24788,N_24548,N_24403);
nand U24789 (N_24789,N_24474,N_24307);
nor U24790 (N_24790,N_24587,N_24579);
nor U24791 (N_24791,N_24575,N_24474);
nand U24792 (N_24792,N_24594,N_24414);
and U24793 (N_24793,N_24458,N_24572);
nor U24794 (N_24794,N_24398,N_24510);
or U24795 (N_24795,N_24316,N_24390);
and U24796 (N_24796,N_24521,N_24540);
xor U24797 (N_24797,N_24372,N_24495);
and U24798 (N_24798,N_24412,N_24348);
nand U24799 (N_24799,N_24513,N_24445);
xnor U24800 (N_24800,N_24412,N_24486);
xnor U24801 (N_24801,N_24379,N_24431);
xor U24802 (N_24802,N_24417,N_24490);
nor U24803 (N_24803,N_24446,N_24509);
xnor U24804 (N_24804,N_24380,N_24505);
nor U24805 (N_24805,N_24455,N_24386);
nand U24806 (N_24806,N_24374,N_24573);
nand U24807 (N_24807,N_24444,N_24337);
and U24808 (N_24808,N_24433,N_24543);
or U24809 (N_24809,N_24333,N_24508);
nor U24810 (N_24810,N_24341,N_24568);
and U24811 (N_24811,N_24591,N_24319);
or U24812 (N_24812,N_24389,N_24301);
nor U24813 (N_24813,N_24531,N_24557);
nand U24814 (N_24814,N_24598,N_24591);
or U24815 (N_24815,N_24483,N_24449);
and U24816 (N_24816,N_24413,N_24404);
and U24817 (N_24817,N_24409,N_24523);
and U24818 (N_24818,N_24452,N_24587);
nor U24819 (N_24819,N_24510,N_24360);
and U24820 (N_24820,N_24396,N_24567);
nor U24821 (N_24821,N_24543,N_24558);
or U24822 (N_24822,N_24320,N_24434);
xor U24823 (N_24823,N_24454,N_24587);
and U24824 (N_24824,N_24314,N_24337);
xnor U24825 (N_24825,N_24333,N_24584);
nand U24826 (N_24826,N_24357,N_24544);
nor U24827 (N_24827,N_24478,N_24598);
nand U24828 (N_24828,N_24594,N_24491);
nor U24829 (N_24829,N_24550,N_24458);
nor U24830 (N_24830,N_24519,N_24411);
xnor U24831 (N_24831,N_24533,N_24304);
or U24832 (N_24832,N_24393,N_24552);
or U24833 (N_24833,N_24556,N_24460);
or U24834 (N_24834,N_24452,N_24337);
or U24835 (N_24835,N_24561,N_24577);
xnor U24836 (N_24836,N_24463,N_24399);
xor U24837 (N_24837,N_24313,N_24429);
xor U24838 (N_24838,N_24348,N_24533);
xnor U24839 (N_24839,N_24552,N_24518);
or U24840 (N_24840,N_24497,N_24567);
nor U24841 (N_24841,N_24549,N_24392);
or U24842 (N_24842,N_24395,N_24484);
and U24843 (N_24843,N_24413,N_24354);
or U24844 (N_24844,N_24512,N_24472);
xor U24845 (N_24845,N_24464,N_24554);
nand U24846 (N_24846,N_24386,N_24465);
xnor U24847 (N_24847,N_24385,N_24570);
xor U24848 (N_24848,N_24307,N_24358);
and U24849 (N_24849,N_24445,N_24317);
xnor U24850 (N_24850,N_24388,N_24302);
or U24851 (N_24851,N_24399,N_24340);
nor U24852 (N_24852,N_24458,N_24470);
nand U24853 (N_24853,N_24330,N_24310);
nor U24854 (N_24854,N_24456,N_24506);
or U24855 (N_24855,N_24303,N_24585);
or U24856 (N_24856,N_24354,N_24331);
and U24857 (N_24857,N_24515,N_24372);
xor U24858 (N_24858,N_24438,N_24553);
nand U24859 (N_24859,N_24549,N_24376);
nor U24860 (N_24860,N_24592,N_24437);
xor U24861 (N_24861,N_24324,N_24555);
or U24862 (N_24862,N_24496,N_24378);
xnor U24863 (N_24863,N_24312,N_24409);
nor U24864 (N_24864,N_24538,N_24340);
xnor U24865 (N_24865,N_24411,N_24433);
xor U24866 (N_24866,N_24312,N_24423);
nand U24867 (N_24867,N_24575,N_24302);
xor U24868 (N_24868,N_24582,N_24372);
and U24869 (N_24869,N_24354,N_24386);
and U24870 (N_24870,N_24454,N_24429);
nand U24871 (N_24871,N_24344,N_24453);
nand U24872 (N_24872,N_24459,N_24580);
and U24873 (N_24873,N_24529,N_24385);
and U24874 (N_24874,N_24461,N_24505);
nor U24875 (N_24875,N_24442,N_24544);
and U24876 (N_24876,N_24598,N_24443);
and U24877 (N_24877,N_24336,N_24498);
or U24878 (N_24878,N_24559,N_24415);
nand U24879 (N_24879,N_24558,N_24578);
xnor U24880 (N_24880,N_24373,N_24556);
nand U24881 (N_24881,N_24537,N_24510);
nor U24882 (N_24882,N_24390,N_24509);
nor U24883 (N_24883,N_24569,N_24524);
or U24884 (N_24884,N_24437,N_24486);
nand U24885 (N_24885,N_24369,N_24581);
xnor U24886 (N_24886,N_24447,N_24429);
nor U24887 (N_24887,N_24523,N_24459);
nand U24888 (N_24888,N_24434,N_24337);
nand U24889 (N_24889,N_24548,N_24421);
and U24890 (N_24890,N_24489,N_24445);
nor U24891 (N_24891,N_24536,N_24471);
nand U24892 (N_24892,N_24457,N_24544);
or U24893 (N_24893,N_24328,N_24535);
xor U24894 (N_24894,N_24456,N_24553);
or U24895 (N_24895,N_24347,N_24357);
nor U24896 (N_24896,N_24516,N_24375);
nor U24897 (N_24897,N_24488,N_24332);
and U24898 (N_24898,N_24440,N_24447);
nand U24899 (N_24899,N_24567,N_24425);
and U24900 (N_24900,N_24848,N_24878);
nor U24901 (N_24901,N_24866,N_24738);
and U24902 (N_24902,N_24623,N_24830);
and U24903 (N_24903,N_24638,N_24750);
nand U24904 (N_24904,N_24825,N_24645);
nand U24905 (N_24905,N_24677,N_24765);
xor U24906 (N_24906,N_24739,N_24846);
or U24907 (N_24907,N_24899,N_24736);
xor U24908 (N_24908,N_24618,N_24757);
nand U24909 (N_24909,N_24636,N_24662);
and U24910 (N_24910,N_24868,N_24772);
nand U24911 (N_24911,N_24760,N_24692);
or U24912 (N_24912,N_24798,N_24873);
and U24913 (N_24913,N_24656,N_24874);
and U24914 (N_24914,N_24784,N_24877);
nor U24915 (N_24915,N_24867,N_24713);
nor U24916 (N_24916,N_24891,N_24630);
nand U24917 (N_24917,N_24897,N_24801);
or U24918 (N_24918,N_24743,N_24763);
nor U24919 (N_24919,N_24755,N_24639);
nor U24920 (N_24920,N_24706,N_24882);
nand U24921 (N_24921,N_24614,N_24853);
or U24922 (N_24922,N_24894,N_24643);
nand U24923 (N_24923,N_24806,N_24740);
nand U24924 (N_24924,N_24881,N_24820);
xnor U24925 (N_24925,N_24754,N_24884);
nor U24926 (N_24926,N_24796,N_24734);
or U24927 (N_24927,N_24833,N_24729);
xor U24928 (N_24928,N_24604,N_24856);
and U24929 (N_24929,N_24646,N_24709);
nor U24930 (N_24930,N_24888,N_24603);
xnor U24931 (N_24931,N_24634,N_24702);
nand U24932 (N_24932,N_24691,N_24889);
or U24933 (N_24933,N_24762,N_24817);
xor U24934 (N_24934,N_24629,N_24771);
and U24935 (N_24935,N_24826,N_24625);
nand U24936 (N_24936,N_24628,N_24880);
nor U24937 (N_24937,N_24815,N_24758);
and U24938 (N_24938,N_24768,N_24697);
nor U24939 (N_24939,N_24865,N_24809);
and U24940 (N_24940,N_24847,N_24606);
xnor U24941 (N_24941,N_24816,N_24620);
and U24942 (N_24942,N_24745,N_24659);
nor U24943 (N_24943,N_24641,N_24624);
xor U24944 (N_24944,N_24876,N_24714);
nand U24945 (N_24945,N_24610,N_24631);
xor U24946 (N_24946,N_24663,N_24720);
nor U24947 (N_24947,N_24864,N_24658);
or U24948 (N_24948,N_24698,N_24753);
xnor U24949 (N_24949,N_24841,N_24674);
nand U24950 (N_24950,N_24651,N_24898);
nor U24951 (N_24951,N_24680,N_24794);
nand U24952 (N_24952,N_24759,N_24664);
and U24953 (N_24953,N_24727,N_24744);
xnor U24954 (N_24954,N_24642,N_24836);
or U24955 (N_24955,N_24667,N_24777);
xor U24956 (N_24956,N_24883,N_24653);
and U24957 (N_24957,N_24601,N_24886);
nor U24958 (N_24958,N_24723,N_24791);
and U24959 (N_24959,N_24704,N_24609);
nor U24960 (N_24960,N_24654,N_24752);
and U24961 (N_24961,N_24655,N_24756);
nor U24962 (N_24962,N_24751,N_24676);
xor U24963 (N_24963,N_24666,N_24797);
and U24964 (N_24964,N_24632,N_24838);
xnor U24965 (N_24965,N_24678,N_24657);
and U24966 (N_24966,N_24672,N_24887);
and U24967 (N_24967,N_24790,N_24776);
xor U24968 (N_24968,N_24792,N_24735);
nand U24969 (N_24969,N_24858,N_24681);
nand U24970 (N_24970,N_24863,N_24605);
nor U24971 (N_24971,N_24748,N_24679);
and U24972 (N_24972,N_24813,N_24840);
or U24973 (N_24973,N_24843,N_24731);
nand U24974 (N_24974,N_24842,N_24780);
and U24975 (N_24975,N_24694,N_24800);
nor U24976 (N_24976,N_24719,N_24885);
xor U24977 (N_24977,N_24823,N_24733);
or U24978 (N_24978,N_24795,N_24831);
and U24979 (N_24979,N_24724,N_24693);
xor U24980 (N_24980,N_24761,N_24728);
xnor U24981 (N_24981,N_24770,N_24730);
nand U24982 (N_24982,N_24608,N_24785);
xnor U24983 (N_24983,N_24712,N_24686);
nor U24984 (N_24984,N_24711,N_24786);
and U24985 (N_24985,N_24708,N_24721);
nand U24986 (N_24986,N_24774,N_24860);
nor U24987 (N_24987,N_24671,N_24742);
or U24988 (N_24988,N_24824,N_24879);
nor U24989 (N_24989,N_24890,N_24648);
xnor U24990 (N_24990,N_24635,N_24633);
or U24991 (N_24991,N_24640,N_24627);
or U24992 (N_24992,N_24644,N_24619);
and U24993 (N_24993,N_24819,N_24822);
nand U24994 (N_24994,N_24726,N_24715);
nand U24995 (N_24995,N_24696,N_24695);
nor U24996 (N_24996,N_24850,N_24861);
nor U24997 (N_24997,N_24647,N_24600);
nand U24998 (N_24998,N_24799,N_24732);
nand U24999 (N_24999,N_24849,N_24870);
nand U25000 (N_25000,N_24788,N_24773);
and U25001 (N_25001,N_24844,N_24805);
nor U25002 (N_25002,N_24893,N_24725);
nand U25003 (N_25003,N_24807,N_24649);
nor U25004 (N_25004,N_24829,N_24690);
xor U25005 (N_25005,N_24689,N_24789);
and U25006 (N_25006,N_24862,N_24812);
or U25007 (N_25007,N_24872,N_24718);
and U25008 (N_25008,N_24617,N_24675);
nor U25009 (N_25009,N_24746,N_24700);
xnor U25010 (N_25010,N_24749,N_24602);
nor U25011 (N_25011,N_24747,N_24717);
or U25012 (N_25012,N_24793,N_24787);
nand U25013 (N_25013,N_24811,N_24835);
xor U25014 (N_25014,N_24637,N_24783);
xnor U25015 (N_25015,N_24814,N_24802);
and U25016 (N_25016,N_24705,N_24661);
nor U25017 (N_25017,N_24626,N_24622);
or U25018 (N_25018,N_24703,N_24804);
and U25019 (N_25019,N_24699,N_24871);
or U25020 (N_25020,N_24845,N_24827);
nand U25021 (N_25021,N_24621,N_24611);
nor U25022 (N_25022,N_24779,N_24818);
or U25023 (N_25023,N_24716,N_24854);
nand U25024 (N_25024,N_24737,N_24767);
or U25025 (N_25025,N_24810,N_24828);
or U25026 (N_25026,N_24821,N_24688);
or U25027 (N_25027,N_24851,N_24684);
nand U25028 (N_25028,N_24685,N_24701);
or U25029 (N_25029,N_24741,N_24660);
or U25030 (N_25030,N_24710,N_24673);
nor U25031 (N_25031,N_24613,N_24669);
nand U25032 (N_25032,N_24896,N_24766);
and U25033 (N_25033,N_24612,N_24834);
nand U25034 (N_25034,N_24670,N_24895);
and U25035 (N_25035,N_24892,N_24832);
xor U25036 (N_25036,N_24859,N_24855);
and U25037 (N_25037,N_24687,N_24808);
or U25038 (N_25038,N_24837,N_24778);
xor U25039 (N_25039,N_24852,N_24707);
xnor U25040 (N_25040,N_24652,N_24683);
and U25041 (N_25041,N_24775,N_24665);
nand U25042 (N_25042,N_24875,N_24782);
and U25043 (N_25043,N_24607,N_24616);
and U25044 (N_25044,N_24839,N_24803);
nor U25045 (N_25045,N_24668,N_24650);
and U25046 (N_25046,N_24869,N_24769);
xor U25047 (N_25047,N_24682,N_24764);
nand U25048 (N_25048,N_24722,N_24857);
xnor U25049 (N_25049,N_24781,N_24615);
or U25050 (N_25050,N_24884,N_24894);
xor U25051 (N_25051,N_24668,N_24829);
xnor U25052 (N_25052,N_24785,N_24636);
nor U25053 (N_25053,N_24610,N_24873);
xor U25054 (N_25054,N_24839,N_24877);
nand U25055 (N_25055,N_24626,N_24892);
or U25056 (N_25056,N_24626,N_24742);
nor U25057 (N_25057,N_24892,N_24759);
nand U25058 (N_25058,N_24719,N_24790);
or U25059 (N_25059,N_24866,N_24777);
or U25060 (N_25060,N_24739,N_24799);
nor U25061 (N_25061,N_24763,N_24678);
and U25062 (N_25062,N_24692,N_24735);
nand U25063 (N_25063,N_24650,N_24789);
nor U25064 (N_25064,N_24605,N_24718);
nor U25065 (N_25065,N_24690,N_24804);
nand U25066 (N_25066,N_24787,N_24866);
nor U25067 (N_25067,N_24711,N_24698);
and U25068 (N_25068,N_24885,N_24748);
xnor U25069 (N_25069,N_24705,N_24644);
and U25070 (N_25070,N_24819,N_24636);
and U25071 (N_25071,N_24759,N_24662);
and U25072 (N_25072,N_24795,N_24640);
and U25073 (N_25073,N_24742,N_24835);
xnor U25074 (N_25074,N_24755,N_24673);
or U25075 (N_25075,N_24624,N_24857);
nor U25076 (N_25076,N_24891,N_24776);
or U25077 (N_25077,N_24668,N_24665);
xnor U25078 (N_25078,N_24745,N_24770);
nand U25079 (N_25079,N_24803,N_24681);
or U25080 (N_25080,N_24797,N_24644);
or U25081 (N_25081,N_24702,N_24787);
nor U25082 (N_25082,N_24707,N_24894);
nand U25083 (N_25083,N_24715,N_24616);
and U25084 (N_25084,N_24846,N_24876);
nor U25085 (N_25085,N_24633,N_24755);
nor U25086 (N_25086,N_24691,N_24704);
nand U25087 (N_25087,N_24783,N_24607);
nor U25088 (N_25088,N_24620,N_24664);
xor U25089 (N_25089,N_24885,N_24658);
and U25090 (N_25090,N_24822,N_24879);
and U25091 (N_25091,N_24773,N_24880);
nor U25092 (N_25092,N_24644,N_24860);
nor U25093 (N_25093,N_24659,N_24667);
and U25094 (N_25094,N_24722,N_24891);
and U25095 (N_25095,N_24827,N_24650);
or U25096 (N_25096,N_24809,N_24665);
and U25097 (N_25097,N_24752,N_24811);
xnor U25098 (N_25098,N_24694,N_24759);
nand U25099 (N_25099,N_24675,N_24747);
nand U25100 (N_25100,N_24729,N_24791);
nand U25101 (N_25101,N_24771,N_24665);
and U25102 (N_25102,N_24739,N_24669);
xnor U25103 (N_25103,N_24842,N_24747);
nand U25104 (N_25104,N_24837,N_24666);
or U25105 (N_25105,N_24802,N_24732);
nand U25106 (N_25106,N_24667,N_24757);
nand U25107 (N_25107,N_24674,N_24799);
nor U25108 (N_25108,N_24848,N_24756);
nor U25109 (N_25109,N_24734,N_24722);
nand U25110 (N_25110,N_24855,N_24621);
or U25111 (N_25111,N_24724,N_24801);
xor U25112 (N_25112,N_24741,N_24607);
xor U25113 (N_25113,N_24782,N_24799);
nor U25114 (N_25114,N_24723,N_24650);
nor U25115 (N_25115,N_24754,N_24649);
and U25116 (N_25116,N_24774,N_24735);
nor U25117 (N_25117,N_24783,N_24601);
or U25118 (N_25118,N_24625,N_24661);
nand U25119 (N_25119,N_24663,N_24624);
nand U25120 (N_25120,N_24662,N_24831);
nor U25121 (N_25121,N_24747,N_24694);
xnor U25122 (N_25122,N_24881,N_24607);
nor U25123 (N_25123,N_24863,N_24880);
nor U25124 (N_25124,N_24632,N_24767);
nand U25125 (N_25125,N_24686,N_24767);
and U25126 (N_25126,N_24734,N_24602);
or U25127 (N_25127,N_24693,N_24872);
and U25128 (N_25128,N_24833,N_24785);
xnor U25129 (N_25129,N_24796,N_24742);
nand U25130 (N_25130,N_24827,N_24683);
nand U25131 (N_25131,N_24666,N_24650);
nor U25132 (N_25132,N_24611,N_24828);
xnor U25133 (N_25133,N_24660,N_24632);
nor U25134 (N_25134,N_24687,N_24806);
nor U25135 (N_25135,N_24661,N_24893);
nand U25136 (N_25136,N_24689,N_24667);
and U25137 (N_25137,N_24700,N_24893);
and U25138 (N_25138,N_24777,N_24683);
nand U25139 (N_25139,N_24652,N_24792);
and U25140 (N_25140,N_24728,N_24811);
nor U25141 (N_25141,N_24841,N_24686);
xor U25142 (N_25142,N_24778,N_24824);
nor U25143 (N_25143,N_24852,N_24626);
nor U25144 (N_25144,N_24745,N_24850);
or U25145 (N_25145,N_24792,N_24801);
nor U25146 (N_25146,N_24816,N_24633);
and U25147 (N_25147,N_24615,N_24727);
and U25148 (N_25148,N_24630,N_24813);
and U25149 (N_25149,N_24784,N_24638);
xnor U25150 (N_25150,N_24652,N_24756);
nor U25151 (N_25151,N_24875,N_24702);
nand U25152 (N_25152,N_24891,N_24812);
or U25153 (N_25153,N_24804,N_24877);
nand U25154 (N_25154,N_24638,N_24861);
nor U25155 (N_25155,N_24818,N_24838);
and U25156 (N_25156,N_24796,N_24733);
xor U25157 (N_25157,N_24612,N_24656);
nand U25158 (N_25158,N_24757,N_24889);
or U25159 (N_25159,N_24731,N_24672);
xnor U25160 (N_25160,N_24893,N_24606);
or U25161 (N_25161,N_24856,N_24665);
xor U25162 (N_25162,N_24793,N_24797);
and U25163 (N_25163,N_24886,N_24724);
nand U25164 (N_25164,N_24771,N_24620);
and U25165 (N_25165,N_24867,N_24624);
or U25166 (N_25166,N_24828,N_24869);
and U25167 (N_25167,N_24899,N_24644);
xor U25168 (N_25168,N_24714,N_24745);
nand U25169 (N_25169,N_24891,N_24851);
nor U25170 (N_25170,N_24698,N_24848);
nor U25171 (N_25171,N_24805,N_24759);
xnor U25172 (N_25172,N_24854,N_24648);
and U25173 (N_25173,N_24647,N_24841);
and U25174 (N_25174,N_24795,N_24750);
and U25175 (N_25175,N_24815,N_24893);
xor U25176 (N_25176,N_24730,N_24758);
nor U25177 (N_25177,N_24731,N_24749);
nand U25178 (N_25178,N_24692,N_24736);
or U25179 (N_25179,N_24876,N_24661);
or U25180 (N_25180,N_24672,N_24774);
nand U25181 (N_25181,N_24818,N_24852);
or U25182 (N_25182,N_24812,N_24663);
and U25183 (N_25183,N_24615,N_24856);
and U25184 (N_25184,N_24671,N_24698);
nor U25185 (N_25185,N_24721,N_24719);
nand U25186 (N_25186,N_24877,N_24649);
nor U25187 (N_25187,N_24676,N_24647);
and U25188 (N_25188,N_24628,N_24699);
xor U25189 (N_25189,N_24624,N_24820);
or U25190 (N_25190,N_24662,N_24828);
or U25191 (N_25191,N_24622,N_24692);
or U25192 (N_25192,N_24767,N_24892);
nand U25193 (N_25193,N_24756,N_24648);
and U25194 (N_25194,N_24816,N_24824);
and U25195 (N_25195,N_24879,N_24765);
nand U25196 (N_25196,N_24729,N_24654);
and U25197 (N_25197,N_24673,N_24687);
xor U25198 (N_25198,N_24716,N_24783);
nand U25199 (N_25199,N_24865,N_24714);
nor U25200 (N_25200,N_24968,N_25071);
or U25201 (N_25201,N_25134,N_25157);
nand U25202 (N_25202,N_24975,N_24945);
nand U25203 (N_25203,N_25159,N_24942);
nor U25204 (N_25204,N_24982,N_25001);
nand U25205 (N_25205,N_25105,N_25058);
or U25206 (N_25206,N_25063,N_25016);
nor U25207 (N_25207,N_24907,N_25146);
and U25208 (N_25208,N_25083,N_24964);
nor U25209 (N_25209,N_24930,N_24997);
or U25210 (N_25210,N_25116,N_25149);
or U25211 (N_25211,N_25018,N_25052);
nor U25212 (N_25212,N_25190,N_25067);
and U25213 (N_25213,N_25039,N_24971);
and U25214 (N_25214,N_25129,N_25133);
or U25215 (N_25215,N_25174,N_25021);
xnor U25216 (N_25216,N_24969,N_24920);
or U25217 (N_25217,N_24958,N_25185);
and U25218 (N_25218,N_25101,N_25141);
xnor U25219 (N_25219,N_24913,N_24904);
xor U25220 (N_25220,N_25181,N_25050);
nor U25221 (N_25221,N_25119,N_25160);
or U25222 (N_25222,N_25009,N_25022);
xor U25223 (N_25223,N_25029,N_25010);
and U25224 (N_25224,N_25164,N_25162);
and U25225 (N_25225,N_25031,N_25128);
or U25226 (N_25226,N_24981,N_25121);
or U25227 (N_25227,N_25135,N_24993);
and U25228 (N_25228,N_25100,N_25172);
xnor U25229 (N_25229,N_25099,N_24980);
nor U25230 (N_25230,N_25048,N_24926);
or U25231 (N_25231,N_25056,N_25082);
or U25232 (N_25232,N_25095,N_24946);
or U25233 (N_25233,N_25012,N_25064);
and U25234 (N_25234,N_25168,N_24962);
or U25235 (N_25235,N_24972,N_25184);
nand U25236 (N_25236,N_25025,N_25166);
and U25237 (N_25237,N_24924,N_25109);
or U25238 (N_25238,N_25180,N_25078);
xor U25239 (N_25239,N_25177,N_25169);
and U25240 (N_25240,N_25062,N_25069);
nor U25241 (N_25241,N_24914,N_25028);
and U25242 (N_25242,N_25111,N_25192);
or U25243 (N_25243,N_25193,N_24955);
nor U25244 (N_25244,N_24952,N_25155);
nand U25245 (N_25245,N_25032,N_25175);
nor U25246 (N_25246,N_25096,N_25170);
and U25247 (N_25247,N_25092,N_25123);
or U25248 (N_25248,N_24929,N_24961);
or U25249 (N_25249,N_25167,N_25005);
and U25250 (N_25250,N_25183,N_25127);
xor U25251 (N_25251,N_25035,N_25026);
and U25252 (N_25252,N_25117,N_25088);
or U25253 (N_25253,N_25171,N_24934);
or U25254 (N_25254,N_25043,N_25036);
nor U25255 (N_25255,N_25107,N_24906);
nand U25256 (N_25256,N_24917,N_25076);
nand U25257 (N_25257,N_24918,N_25004);
or U25258 (N_25258,N_25103,N_25098);
nor U25259 (N_25259,N_25089,N_24931);
and U25260 (N_25260,N_24984,N_25113);
xnor U25261 (N_25261,N_25061,N_25131);
and U25262 (N_25262,N_24905,N_24996);
xnor U25263 (N_25263,N_25115,N_25199);
and U25264 (N_25264,N_24951,N_24992);
and U25265 (N_25265,N_25027,N_25173);
nand U25266 (N_25266,N_25077,N_24940);
nand U25267 (N_25267,N_25075,N_25042);
nor U25268 (N_25268,N_24999,N_24970);
xnor U25269 (N_25269,N_25030,N_24943);
nand U25270 (N_25270,N_24990,N_25110);
nor U25271 (N_25271,N_25065,N_25163);
nand U25272 (N_25272,N_25114,N_25142);
nor U25273 (N_25273,N_25084,N_25093);
nand U25274 (N_25274,N_25106,N_25102);
xnor U25275 (N_25275,N_25060,N_25156);
nor U25276 (N_25276,N_25158,N_25085);
nand U25277 (N_25277,N_25033,N_25140);
xnor U25278 (N_25278,N_25070,N_24973);
and U25279 (N_25279,N_24935,N_25047);
nand U25280 (N_25280,N_25148,N_25112);
or U25281 (N_25281,N_25057,N_24902);
or U25282 (N_25282,N_25153,N_24966);
nand U25283 (N_25283,N_24915,N_24938);
nor U25284 (N_25284,N_24919,N_24967);
or U25285 (N_25285,N_25037,N_25179);
xnor U25286 (N_25286,N_25197,N_25125);
xnor U25287 (N_25287,N_25013,N_25130);
nand U25288 (N_25288,N_25019,N_25139);
or U25289 (N_25289,N_24978,N_25194);
nand U25290 (N_25290,N_25132,N_24956);
xnor U25291 (N_25291,N_24909,N_25151);
nor U25292 (N_25292,N_24936,N_25154);
nor U25293 (N_25293,N_25104,N_25152);
xnor U25294 (N_25294,N_24985,N_25189);
and U25295 (N_25295,N_25161,N_25087);
xor U25296 (N_25296,N_24900,N_25002);
nand U25297 (N_25297,N_25147,N_24932);
nor U25298 (N_25298,N_24901,N_25079);
nor U25299 (N_25299,N_25003,N_25091);
nor U25300 (N_25300,N_24965,N_25086);
xor U25301 (N_25301,N_24954,N_25074);
or U25302 (N_25302,N_25007,N_25011);
or U25303 (N_25303,N_25186,N_24921);
or U25304 (N_25304,N_25040,N_24949);
nor U25305 (N_25305,N_25000,N_25024);
and U25306 (N_25306,N_25097,N_24994);
or U25307 (N_25307,N_24908,N_25138);
nor U25308 (N_25308,N_25195,N_24998);
and U25309 (N_25309,N_25046,N_24989);
xnor U25310 (N_25310,N_25108,N_24953);
or U25311 (N_25311,N_25122,N_25144);
nand U25312 (N_25312,N_24995,N_24977);
xnor U25313 (N_25313,N_24957,N_25118);
nor U25314 (N_25314,N_25196,N_24925);
nand U25315 (N_25315,N_24927,N_24939);
nand U25316 (N_25316,N_24944,N_25054);
and U25317 (N_25317,N_24947,N_25182);
nor U25318 (N_25318,N_25188,N_25198);
and U25319 (N_25319,N_25049,N_24991);
and U25320 (N_25320,N_25150,N_25051);
or U25321 (N_25321,N_25145,N_24922);
or U25322 (N_25322,N_25044,N_24941);
and U25323 (N_25323,N_25055,N_24923);
or U25324 (N_25324,N_25176,N_25072);
nand U25325 (N_25325,N_25073,N_25059);
or U25326 (N_25326,N_25126,N_25143);
or U25327 (N_25327,N_24976,N_25041);
or U25328 (N_25328,N_25017,N_24986);
nor U25329 (N_25329,N_24979,N_25053);
nor U25330 (N_25330,N_25178,N_25136);
xnor U25331 (N_25331,N_24983,N_25120);
nand U25332 (N_25332,N_25006,N_24911);
nand U25333 (N_25333,N_25081,N_24988);
and U25334 (N_25334,N_24974,N_24950);
or U25335 (N_25335,N_25124,N_24987);
or U25336 (N_25336,N_25008,N_24948);
or U25337 (N_25337,N_25066,N_24910);
xnor U25338 (N_25338,N_24963,N_24903);
or U25339 (N_25339,N_25165,N_24959);
and U25340 (N_25340,N_25090,N_25068);
nand U25341 (N_25341,N_24933,N_25014);
nor U25342 (N_25342,N_25015,N_25137);
nor U25343 (N_25343,N_25023,N_24916);
xnor U25344 (N_25344,N_25034,N_25080);
or U25345 (N_25345,N_25038,N_25094);
nand U25346 (N_25346,N_24912,N_25187);
or U25347 (N_25347,N_24928,N_24960);
or U25348 (N_25348,N_24937,N_25045);
or U25349 (N_25349,N_25191,N_25020);
or U25350 (N_25350,N_24941,N_24940);
xor U25351 (N_25351,N_24975,N_25156);
nand U25352 (N_25352,N_25103,N_24983);
or U25353 (N_25353,N_24974,N_25104);
and U25354 (N_25354,N_25183,N_24945);
xor U25355 (N_25355,N_24913,N_24903);
nor U25356 (N_25356,N_24965,N_25096);
nand U25357 (N_25357,N_24960,N_25113);
nor U25358 (N_25358,N_25056,N_24919);
or U25359 (N_25359,N_24973,N_24937);
nand U25360 (N_25360,N_25062,N_24965);
xnor U25361 (N_25361,N_24909,N_25120);
or U25362 (N_25362,N_24986,N_25087);
nor U25363 (N_25363,N_25047,N_24995);
xnor U25364 (N_25364,N_25001,N_25078);
and U25365 (N_25365,N_24985,N_24901);
or U25366 (N_25366,N_25191,N_25152);
xnor U25367 (N_25367,N_25011,N_25187);
or U25368 (N_25368,N_25078,N_24988);
xor U25369 (N_25369,N_25098,N_25174);
or U25370 (N_25370,N_25024,N_25152);
xor U25371 (N_25371,N_25156,N_24904);
nor U25372 (N_25372,N_24982,N_25043);
xnor U25373 (N_25373,N_25161,N_24998);
and U25374 (N_25374,N_25081,N_24934);
or U25375 (N_25375,N_25081,N_24955);
nand U25376 (N_25376,N_24919,N_25044);
nand U25377 (N_25377,N_24961,N_24921);
or U25378 (N_25378,N_25098,N_25151);
nand U25379 (N_25379,N_25154,N_25105);
and U25380 (N_25380,N_25115,N_25017);
or U25381 (N_25381,N_25026,N_25046);
and U25382 (N_25382,N_25160,N_24974);
or U25383 (N_25383,N_25186,N_25048);
nand U25384 (N_25384,N_24993,N_25157);
or U25385 (N_25385,N_25161,N_25034);
xnor U25386 (N_25386,N_25052,N_25108);
and U25387 (N_25387,N_24941,N_24904);
xor U25388 (N_25388,N_25025,N_24902);
or U25389 (N_25389,N_25159,N_24931);
or U25390 (N_25390,N_24963,N_24969);
nor U25391 (N_25391,N_25074,N_25012);
nand U25392 (N_25392,N_24939,N_25067);
nor U25393 (N_25393,N_25021,N_25045);
xnor U25394 (N_25394,N_25199,N_24916);
nor U25395 (N_25395,N_25180,N_25072);
nand U25396 (N_25396,N_25195,N_25015);
nand U25397 (N_25397,N_25112,N_25167);
and U25398 (N_25398,N_25111,N_25102);
xnor U25399 (N_25399,N_24975,N_24986);
and U25400 (N_25400,N_24967,N_25055);
xnor U25401 (N_25401,N_25011,N_25154);
nor U25402 (N_25402,N_25167,N_25001);
xor U25403 (N_25403,N_24945,N_25058);
nor U25404 (N_25404,N_24945,N_24921);
and U25405 (N_25405,N_25150,N_24980);
nor U25406 (N_25406,N_25179,N_25086);
xnor U25407 (N_25407,N_25180,N_24993);
or U25408 (N_25408,N_25138,N_24945);
nor U25409 (N_25409,N_25007,N_25153);
xor U25410 (N_25410,N_24990,N_25014);
nor U25411 (N_25411,N_25073,N_25139);
or U25412 (N_25412,N_24908,N_25128);
xor U25413 (N_25413,N_25038,N_25052);
and U25414 (N_25414,N_24986,N_24984);
and U25415 (N_25415,N_25123,N_25127);
and U25416 (N_25416,N_25070,N_25111);
and U25417 (N_25417,N_24923,N_25196);
and U25418 (N_25418,N_25117,N_24948);
or U25419 (N_25419,N_25160,N_25021);
or U25420 (N_25420,N_25164,N_25099);
and U25421 (N_25421,N_24997,N_25087);
or U25422 (N_25422,N_24930,N_24957);
xor U25423 (N_25423,N_24957,N_25077);
or U25424 (N_25424,N_24950,N_24957);
xor U25425 (N_25425,N_25134,N_25164);
nand U25426 (N_25426,N_25065,N_24996);
nor U25427 (N_25427,N_25154,N_25005);
nor U25428 (N_25428,N_24916,N_25104);
and U25429 (N_25429,N_24984,N_25160);
or U25430 (N_25430,N_24949,N_25084);
xnor U25431 (N_25431,N_25006,N_25183);
xnor U25432 (N_25432,N_25170,N_24967);
nand U25433 (N_25433,N_25132,N_25105);
nand U25434 (N_25434,N_25126,N_25009);
nand U25435 (N_25435,N_25061,N_25142);
xnor U25436 (N_25436,N_25095,N_24987);
or U25437 (N_25437,N_25011,N_24913);
and U25438 (N_25438,N_25171,N_25080);
xor U25439 (N_25439,N_24993,N_25177);
xor U25440 (N_25440,N_24901,N_24949);
xnor U25441 (N_25441,N_25197,N_25126);
nor U25442 (N_25442,N_24947,N_25194);
nand U25443 (N_25443,N_24971,N_25181);
xnor U25444 (N_25444,N_24911,N_25168);
nand U25445 (N_25445,N_25184,N_24973);
nor U25446 (N_25446,N_24963,N_25141);
nand U25447 (N_25447,N_25041,N_25098);
nor U25448 (N_25448,N_24909,N_25121);
xor U25449 (N_25449,N_25025,N_24955);
and U25450 (N_25450,N_25067,N_25059);
and U25451 (N_25451,N_25192,N_24999);
and U25452 (N_25452,N_24963,N_25140);
nor U25453 (N_25453,N_25190,N_25051);
nor U25454 (N_25454,N_24932,N_25191);
or U25455 (N_25455,N_24970,N_24931);
and U25456 (N_25456,N_25070,N_24920);
and U25457 (N_25457,N_24962,N_25167);
xor U25458 (N_25458,N_25147,N_25158);
xor U25459 (N_25459,N_25134,N_24949);
nor U25460 (N_25460,N_25061,N_25092);
and U25461 (N_25461,N_25186,N_24933);
xor U25462 (N_25462,N_25118,N_25173);
and U25463 (N_25463,N_25114,N_24900);
xnor U25464 (N_25464,N_25065,N_25054);
or U25465 (N_25465,N_25155,N_25082);
nand U25466 (N_25466,N_25135,N_25065);
xnor U25467 (N_25467,N_24904,N_25035);
nand U25468 (N_25468,N_24943,N_25171);
or U25469 (N_25469,N_25148,N_25175);
or U25470 (N_25470,N_25188,N_25008);
nor U25471 (N_25471,N_25010,N_25132);
xnor U25472 (N_25472,N_25156,N_25039);
nor U25473 (N_25473,N_25169,N_25141);
xor U25474 (N_25474,N_25034,N_25088);
nand U25475 (N_25475,N_24912,N_25066);
or U25476 (N_25476,N_25179,N_24929);
and U25477 (N_25477,N_25076,N_24942);
xor U25478 (N_25478,N_25021,N_25133);
nand U25479 (N_25479,N_24999,N_24950);
nor U25480 (N_25480,N_24927,N_25145);
xnor U25481 (N_25481,N_25076,N_25059);
nand U25482 (N_25482,N_24932,N_25113);
or U25483 (N_25483,N_25057,N_25012);
or U25484 (N_25484,N_25068,N_24920);
xnor U25485 (N_25485,N_25066,N_24909);
nor U25486 (N_25486,N_24979,N_25101);
nor U25487 (N_25487,N_24971,N_24925);
nor U25488 (N_25488,N_25025,N_24981);
nor U25489 (N_25489,N_24981,N_24923);
nor U25490 (N_25490,N_24957,N_25145);
or U25491 (N_25491,N_25115,N_25072);
xnor U25492 (N_25492,N_24991,N_24993);
or U25493 (N_25493,N_25058,N_25158);
or U25494 (N_25494,N_24947,N_25110);
nor U25495 (N_25495,N_25054,N_24920);
nand U25496 (N_25496,N_25005,N_25003);
nand U25497 (N_25497,N_25142,N_25144);
or U25498 (N_25498,N_25190,N_24912);
nor U25499 (N_25499,N_24934,N_24907);
nand U25500 (N_25500,N_25343,N_25425);
xor U25501 (N_25501,N_25332,N_25443);
or U25502 (N_25502,N_25255,N_25494);
and U25503 (N_25503,N_25473,N_25471);
nor U25504 (N_25504,N_25424,N_25366);
and U25505 (N_25505,N_25364,N_25479);
nor U25506 (N_25506,N_25340,N_25422);
nor U25507 (N_25507,N_25334,N_25347);
and U25508 (N_25508,N_25271,N_25220);
or U25509 (N_25509,N_25392,N_25469);
and U25510 (N_25510,N_25278,N_25468);
nand U25511 (N_25511,N_25326,N_25266);
or U25512 (N_25512,N_25493,N_25359);
xor U25513 (N_25513,N_25367,N_25263);
or U25514 (N_25514,N_25498,N_25476);
nand U25515 (N_25515,N_25400,N_25465);
nor U25516 (N_25516,N_25411,N_25451);
xnor U25517 (N_25517,N_25415,N_25279);
nand U25518 (N_25518,N_25224,N_25333);
nand U25519 (N_25519,N_25276,N_25368);
or U25520 (N_25520,N_25209,N_25416);
or U25521 (N_25521,N_25399,N_25251);
nor U25522 (N_25522,N_25254,N_25264);
nand U25523 (N_25523,N_25309,N_25310);
xnor U25524 (N_25524,N_25448,N_25337);
nand U25525 (N_25525,N_25436,N_25307);
nand U25526 (N_25526,N_25398,N_25496);
and U25527 (N_25527,N_25317,N_25236);
nand U25528 (N_25528,N_25238,N_25222);
or U25529 (N_25529,N_25201,N_25461);
xnor U25530 (N_25530,N_25256,N_25258);
xnor U25531 (N_25531,N_25381,N_25444);
nor U25532 (N_25532,N_25466,N_25235);
xnor U25533 (N_25533,N_25228,N_25316);
nor U25534 (N_25534,N_25455,N_25369);
and U25535 (N_25535,N_25357,N_25243);
nand U25536 (N_25536,N_25484,N_25402);
and U25537 (N_25537,N_25418,N_25295);
nand U25538 (N_25538,N_25352,N_25265);
or U25539 (N_25539,N_25430,N_25214);
nand U25540 (N_25540,N_25259,N_25312);
or U25541 (N_25541,N_25300,N_25252);
or U25542 (N_25542,N_25241,N_25495);
nand U25543 (N_25543,N_25287,N_25206);
nand U25544 (N_25544,N_25233,N_25290);
or U25545 (N_25545,N_25217,N_25377);
xnor U25546 (N_25546,N_25477,N_25480);
nand U25547 (N_25547,N_25410,N_25203);
nor U25548 (N_25548,N_25298,N_25325);
or U25549 (N_25549,N_25488,N_25296);
nand U25550 (N_25550,N_25239,N_25490);
and U25551 (N_25551,N_25302,N_25439);
xnor U25552 (N_25552,N_25331,N_25385);
xnor U25553 (N_25553,N_25285,N_25244);
nor U25554 (N_25554,N_25387,N_25375);
xor U25555 (N_25555,N_25210,N_25261);
xor U25556 (N_25556,N_25478,N_25237);
or U25557 (N_25557,N_25453,N_25274);
nand U25558 (N_25558,N_25486,N_25354);
nand U25559 (N_25559,N_25470,N_25240);
and U25560 (N_25560,N_25314,N_25351);
nand U25561 (N_25561,N_25219,N_25404);
nand U25562 (N_25562,N_25339,N_25345);
nor U25563 (N_25563,N_25463,N_25429);
xnor U25564 (N_25564,N_25313,N_25421);
nand U25565 (N_25565,N_25462,N_25474);
and U25566 (N_25566,N_25320,N_25389);
xnor U25567 (N_25567,N_25293,N_25407);
nand U25568 (N_25568,N_25268,N_25499);
or U25569 (N_25569,N_25412,N_25452);
nand U25570 (N_25570,N_25438,N_25289);
nor U25571 (N_25571,N_25207,N_25446);
and U25572 (N_25572,N_25353,N_25409);
nand U25573 (N_25573,N_25327,N_25342);
nand U25574 (N_25574,N_25401,N_25346);
nand U25575 (N_25575,N_25382,N_25384);
xor U25576 (N_25576,N_25344,N_25380);
nand U25577 (N_25577,N_25205,N_25202);
xnor U25578 (N_25578,N_25335,N_25482);
or U25579 (N_25579,N_25288,N_25456);
nor U25580 (N_25580,N_25489,N_25226);
xor U25581 (N_25581,N_25371,N_25286);
xnor U25582 (N_25582,N_25281,N_25267);
xor U25583 (N_25583,N_25437,N_25225);
and U25584 (N_25584,N_25397,N_25372);
and U25585 (N_25585,N_25200,N_25434);
and U25586 (N_25586,N_25291,N_25356);
or U25587 (N_25587,N_25294,N_25405);
and U25588 (N_25588,N_25472,N_25242);
and U25589 (N_25589,N_25458,N_25248);
or U25590 (N_25590,N_25445,N_25282);
nand U25591 (N_25591,N_25432,N_25403);
or U25592 (N_25592,N_25299,N_25379);
xor U25593 (N_25593,N_25459,N_25395);
and U25594 (N_25594,N_25460,N_25230);
nor U25595 (N_25595,N_25301,N_25360);
nand U25596 (N_25596,N_25249,N_25363);
xnor U25597 (N_25597,N_25348,N_25246);
and U25598 (N_25598,N_25336,N_25284);
nor U25599 (N_25599,N_25338,N_25441);
xor U25600 (N_25600,N_25215,N_25454);
xor U25601 (N_25601,N_25483,N_25341);
nand U25602 (N_25602,N_25303,N_25435);
nor U25603 (N_25603,N_25247,N_25370);
nor U25604 (N_25604,N_25250,N_25253);
nor U25605 (N_25605,N_25406,N_25277);
or U25606 (N_25606,N_25318,N_25433);
nor U25607 (N_25607,N_25417,N_25427);
nor U25608 (N_25608,N_25408,N_25213);
nand U25609 (N_25609,N_25362,N_25464);
xnor U25610 (N_25610,N_25485,N_25492);
xor U25611 (N_25611,N_25391,N_25328);
nor U25612 (N_25612,N_25204,N_25383);
nor U25613 (N_25613,N_25275,N_25229);
nor U25614 (N_25614,N_25283,N_25272);
xnor U25615 (N_25615,N_25423,N_25218);
nand U25616 (N_25616,N_25428,N_25390);
nand U25617 (N_25617,N_25450,N_25308);
nand U25618 (N_25618,N_25315,N_25413);
nor U25619 (N_25619,N_25440,N_25208);
and U25620 (N_25620,N_25306,N_25234);
or U25621 (N_25621,N_25467,N_25221);
nor U25622 (N_25622,N_25358,N_25324);
nand U25623 (N_25623,N_25420,N_25481);
nor U25624 (N_25624,N_25487,N_25319);
xnor U25625 (N_25625,N_25393,N_25475);
and U25626 (N_25626,N_25216,N_25223);
nor U25627 (N_25627,N_25311,N_25361);
and U25628 (N_25628,N_25442,N_25449);
and U25629 (N_25629,N_25227,N_25245);
and U25630 (N_25630,N_25373,N_25269);
or U25631 (N_25631,N_25376,N_25270);
nand U25632 (N_25632,N_25280,N_25447);
nor U25633 (N_25633,N_25232,N_25394);
xnor U25634 (N_25634,N_25330,N_25365);
or U25635 (N_25635,N_25304,N_25431);
nand U25636 (N_25636,N_25297,N_25497);
nand U25637 (N_25637,N_25260,N_25273);
xor U25638 (N_25638,N_25378,N_25419);
nor U25639 (N_25639,N_25349,N_25350);
and U25640 (N_25640,N_25329,N_25231);
xnor U25641 (N_25641,N_25388,N_25491);
or U25642 (N_25642,N_25322,N_25414);
or U25643 (N_25643,N_25211,N_25457);
or U25644 (N_25644,N_25262,N_25355);
xnor U25645 (N_25645,N_25257,N_25323);
nor U25646 (N_25646,N_25396,N_25292);
xor U25647 (N_25647,N_25374,N_25386);
nand U25648 (N_25648,N_25305,N_25212);
nand U25649 (N_25649,N_25321,N_25426);
nor U25650 (N_25650,N_25281,N_25373);
and U25651 (N_25651,N_25369,N_25249);
nor U25652 (N_25652,N_25370,N_25372);
and U25653 (N_25653,N_25332,N_25226);
nor U25654 (N_25654,N_25335,N_25441);
nand U25655 (N_25655,N_25394,N_25412);
xor U25656 (N_25656,N_25201,N_25200);
nor U25657 (N_25657,N_25251,N_25418);
or U25658 (N_25658,N_25271,N_25361);
nand U25659 (N_25659,N_25364,N_25254);
and U25660 (N_25660,N_25309,N_25218);
xnor U25661 (N_25661,N_25406,N_25440);
nand U25662 (N_25662,N_25348,N_25268);
or U25663 (N_25663,N_25220,N_25321);
xor U25664 (N_25664,N_25292,N_25331);
and U25665 (N_25665,N_25232,N_25219);
nor U25666 (N_25666,N_25217,N_25340);
and U25667 (N_25667,N_25498,N_25382);
and U25668 (N_25668,N_25229,N_25351);
xor U25669 (N_25669,N_25491,N_25422);
nand U25670 (N_25670,N_25272,N_25446);
xor U25671 (N_25671,N_25389,N_25327);
nor U25672 (N_25672,N_25381,N_25463);
and U25673 (N_25673,N_25219,N_25222);
nor U25674 (N_25674,N_25328,N_25413);
and U25675 (N_25675,N_25290,N_25454);
xor U25676 (N_25676,N_25306,N_25244);
and U25677 (N_25677,N_25449,N_25423);
nor U25678 (N_25678,N_25413,N_25201);
or U25679 (N_25679,N_25346,N_25440);
and U25680 (N_25680,N_25239,N_25284);
nor U25681 (N_25681,N_25250,N_25225);
nand U25682 (N_25682,N_25204,N_25393);
nand U25683 (N_25683,N_25400,N_25367);
or U25684 (N_25684,N_25339,N_25427);
nor U25685 (N_25685,N_25294,N_25357);
nand U25686 (N_25686,N_25360,N_25329);
and U25687 (N_25687,N_25213,N_25466);
or U25688 (N_25688,N_25245,N_25301);
or U25689 (N_25689,N_25337,N_25412);
nor U25690 (N_25690,N_25469,N_25210);
xor U25691 (N_25691,N_25247,N_25485);
and U25692 (N_25692,N_25200,N_25217);
xor U25693 (N_25693,N_25373,N_25200);
xor U25694 (N_25694,N_25249,N_25471);
and U25695 (N_25695,N_25328,N_25282);
and U25696 (N_25696,N_25327,N_25440);
nor U25697 (N_25697,N_25211,N_25330);
nor U25698 (N_25698,N_25427,N_25393);
or U25699 (N_25699,N_25302,N_25422);
or U25700 (N_25700,N_25402,N_25464);
nor U25701 (N_25701,N_25358,N_25308);
nor U25702 (N_25702,N_25432,N_25399);
or U25703 (N_25703,N_25427,N_25430);
and U25704 (N_25704,N_25292,N_25354);
nand U25705 (N_25705,N_25285,N_25368);
nor U25706 (N_25706,N_25319,N_25495);
nor U25707 (N_25707,N_25263,N_25438);
xor U25708 (N_25708,N_25232,N_25425);
nor U25709 (N_25709,N_25305,N_25488);
xnor U25710 (N_25710,N_25477,N_25448);
xor U25711 (N_25711,N_25472,N_25241);
nor U25712 (N_25712,N_25293,N_25435);
or U25713 (N_25713,N_25217,N_25416);
or U25714 (N_25714,N_25326,N_25353);
xnor U25715 (N_25715,N_25433,N_25361);
nor U25716 (N_25716,N_25477,N_25306);
or U25717 (N_25717,N_25323,N_25204);
or U25718 (N_25718,N_25243,N_25263);
nor U25719 (N_25719,N_25304,N_25345);
nor U25720 (N_25720,N_25387,N_25462);
or U25721 (N_25721,N_25491,N_25404);
and U25722 (N_25722,N_25472,N_25361);
or U25723 (N_25723,N_25412,N_25411);
and U25724 (N_25724,N_25251,N_25481);
nand U25725 (N_25725,N_25349,N_25348);
or U25726 (N_25726,N_25496,N_25392);
xnor U25727 (N_25727,N_25204,N_25316);
nor U25728 (N_25728,N_25292,N_25291);
nor U25729 (N_25729,N_25245,N_25232);
and U25730 (N_25730,N_25295,N_25270);
or U25731 (N_25731,N_25437,N_25235);
xor U25732 (N_25732,N_25346,N_25257);
and U25733 (N_25733,N_25248,N_25334);
or U25734 (N_25734,N_25408,N_25371);
nand U25735 (N_25735,N_25491,N_25395);
or U25736 (N_25736,N_25248,N_25333);
xor U25737 (N_25737,N_25343,N_25434);
and U25738 (N_25738,N_25227,N_25266);
xnor U25739 (N_25739,N_25450,N_25272);
xor U25740 (N_25740,N_25301,N_25330);
and U25741 (N_25741,N_25286,N_25455);
xor U25742 (N_25742,N_25356,N_25478);
and U25743 (N_25743,N_25447,N_25271);
or U25744 (N_25744,N_25492,N_25271);
xnor U25745 (N_25745,N_25224,N_25269);
xnor U25746 (N_25746,N_25358,N_25203);
and U25747 (N_25747,N_25405,N_25359);
nor U25748 (N_25748,N_25332,N_25273);
nor U25749 (N_25749,N_25386,N_25455);
xor U25750 (N_25750,N_25200,N_25311);
or U25751 (N_25751,N_25319,N_25359);
nor U25752 (N_25752,N_25497,N_25317);
xor U25753 (N_25753,N_25333,N_25211);
xor U25754 (N_25754,N_25350,N_25470);
nand U25755 (N_25755,N_25470,N_25265);
xor U25756 (N_25756,N_25413,N_25356);
xor U25757 (N_25757,N_25240,N_25328);
nand U25758 (N_25758,N_25401,N_25391);
xor U25759 (N_25759,N_25312,N_25341);
or U25760 (N_25760,N_25201,N_25253);
and U25761 (N_25761,N_25272,N_25441);
and U25762 (N_25762,N_25438,N_25357);
nor U25763 (N_25763,N_25385,N_25486);
and U25764 (N_25764,N_25390,N_25494);
and U25765 (N_25765,N_25334,N_25446);
nand U25766 (N_25766,N_25305,N_25277);
and U25767 (N_25767,N_25243,N_25286);
xnor U25768 (N_25768,N_25298,N_25453);
and U25769 (N_25769,N_25345,N_25474);
nand U25770 (N_25770,N_25331,N_25421);
or U25771 (N_25771,N_25220,N_25277);
or U25772 (N_25772,N_25375,N_25269);
nand U25773 (N_25773,N_25203,N_25460);
xnor U25774 (N_25774,N_25498,N_25259);
nor U25775 (N_25775,N_25321,N_25382);
and U25776 (N_25776,N_25368,N_25280);
xor U25777 (N_25777,N_25407,N_25367);
or U25778 (N_25778,N_25464,N_25267);
or U25779 (N_25779,N_25317,N_25361);
nor U25780 (N_25780,N_25225,N_25438);
xnor U25781 (N_25781,N_25400,N_25439);
and U25782 (N_25782,N_25445,N_25358);
nand U25783 (N_25783,N_25354,N_25207);
and U25784 (N_25784,N_25392,N_25464);
nor U25785 (N_25785,N_25202,N_25249);
nand U25786 (N_25786,N_25326,N_25294);
xor U25787 (N_25787,N_25456,N_25414);
xor U25788 (N_25788,N_25332,N_25401);
nor U25789 (N_25789,N_25316,N_25303);
or U25790 (N_25790,N_25406,N_25470);
and U25791 (N_25791,N_25207,N_25286);
nor U25792 (N_25792,N_25301,N_25318);
nand U25793 (N_25793,N_25460,N_25428);
nor U25794 (N_25794,N_25219,N_25427);
nand U25795 (N_25795,N_25395,N_25287);
nor U25796 (N_25796,N_25269,N_25365);
xnor U25797 (N_25797,N_25487,N_25498);
or U25798 (N_25798,N_25241,N_25218);
nor U25799 (N_25799,N_25208,N_25442);
nand U25800 (N_25800,N_25587,N_25700);
xor U25801 (N_25801,N_25754,N_25578);
or U25802 (N_25802,N_25728,N_25607);
and U25803 (N_25803,N_25570,N_25563);
xor U25804 (N_25804,N_25575,N_25509);
xnor U25805 (N_25805,N_25547,N_25651);
and U25806 (N_25806,N_25737,N_25784);
or U25807 (N_25807,N_25705,N_25565);
nand U25808 (N_25808,N_25715,N_25500);
xnor U25809 (N_25809,N_25615,N_25529);
nand U25810 (N_25810,N_25766,N_25709);
xor U25811 (N_25811,N_25600,N_25734);
xor U25812 (N_25812,N_25557,N_25512);
and U25813 (N_25813,N_25719,N_25538);
or U25814 (N_25814,N_25636,N_25762);
nand U25815 (N_25815,N_25723,N_25517);
or U25816 (N_25816,N_25535,N_25701);
nand U25817 (N_25817,N_25708,N_25748);
and U25818 (N_25818,N_25763,N_25634);
nand U25819 (N_25819,N_25664,N_25614);
nand U25820 (N_25820,N_25626,N_25716);
nor U25821 (N_25821,N_25585,N_25702);
or U25822 (N_25822,N_25528,N_25628);
and U25823 (N_25823,N_25774,N_25541);
nand U25824 (N_25824,N_25757,N_25554);
or U25825 (N_25825,N_25525,N_25521);
xor U25826 (N_25826,N_25610,N_25631);
and U25827 (N_25827,N_25520,N_25510);
nand U25828 (N_25828,N_25697,N_25682);
xor U25829 (N_25829,N_25523,N_25662);
xnor U25830 (N_25830,N_25759,N_25548);
nand U25831 (N_25831,N_25658,N_25676);
or U25832 (N_25832,N_25657,N_25789);
nor U25833 (N_25833,N_25542,N_25706);
nor U25834 (N_25834,N_25556,N_25712);
and U25835 (N_25835,N_25597,N_25750);
nand U25836 (N_25836,N_25777,N_25796);
and U25837 (N_25837,N_25736,N_25572);
nor U25838 (N_25838,N_25539,N_25632);
or U25839 (N_25839,N_25647,N_25511);
or U25840 (N_25840,N_25718,N_25699);
and U25841 (N_25841,N_25668,N_25502);
nor U25842 (N_25842,N_25641,N_25792);
nand U25843 (N_25843,N_25791,N_25749);
nand U25844 (N_25844,N_25770,N_25503);
nand U25845 (N_25845,N_25644,N_25665);
nand U25846 (N_25846,N_25555,N_25695);
nand U25847 (N_25847,N_25619,N_25506);
or U25848 (N_25848,N_25733,N_25599);
nand U25849 (N_25849,N_25663,N_25751);
nand U25850 (N_25850,N_25522,N_25735);
nand U25851 (N_25851,N_25711,N_25678);
xnor U25852 (N_25852,N_25624,N_25581);
nor U25853 (N_25853,N_25747,N_25568);
nor U25854 (N_25854,N_25652,N_25732);
xor U25855 (N_25855,N_25703,N_25524);
and U25856 (N_25856,N_25680,N_25787);
nand U25857 (N_25857,N_25633,N_25544);
and U25858 (N_25858,N_25534,N_25666);
nand U25859 (N_25859,N_25753,N_25620);
nand U25860 (N_25860,N_25518,N_25661);
nand U25861 (N_25861,N_25635,N_25710);
and U25862 (N_25862,N_25726,N_25507);
nand U25863 (N_25863,N_25769,N_25781);
or U25864 (N_25864,N_25637,N_25639);
nand U25865 (N_25865,N_25707,N_25677);
nor U25866 (N_25866,N_25782,N_25629);
nand U25867 (N_25867,N_25516,N_25551);
and U25868 (N_25868,N_25567,N_25767);
and U25869 (N_25869,N_25768,N_25640);
and U25870 (N_25870,N_25566,N_25739);
xor U25871 (N_25871,N_25618,N_25569);
and U25872 (N_25872,N_25625,N_25617);
xor U25873 (N_25873,N_25760,N_25613);
nor U25874 (N_25874,N_25508,N_25689);
nand U25875 (N_25875,N_25616,N_25744);
and U25876 (N_25876,N_25590,N_25693);
nor U25877 (N_25877,N_25681,N_25729);
xor U25878 (N_25878,N_25721,N_25596);
nor U25879 (N_25879,N_25799,N_25505);
nand U25880 (N_25880,N_25582,N_25630);
nand U25881 (N_25881,N_25691,N_25559);
and U25882 (N_25882,N_25650,N_25622);
or U25883 (N_25883,N_25558,N_25532);
nand U25884 (N_25884,N_25653,N_25771);
xor U25885 (N_25885,N_25722,N_25561);
nand U25886 (N_25886,N_25793,N_25571);
and U25887 (N_25887,N_25713,N_25724);
nand U25888 (N_25888,N_25783,N_25758);
xor U25889 (N_25889,N_25501,N_25594);
xnor U25890 (N_25890,N_25584,N_25642);
or U25891 (N_25891,N_25765,N_25794);
or U25892 (N_25892,N_25683,N_25772);
nand U25893 (N_25893,N_25595,N_25580);
xor U25894 (N_25894,N_25564,N_25755);
nor U25895 (N_25895,N_25798,N_25745);
nand U25896 (N_25896,N_25545,N_25577);
or U25897 (N_25897,N_25649,N_25519);
and U25898 (N_25898,N_25589,N_25688);
or U25899 (N_25899,N_25741,N_25779);
nor U25900 (N_25900,N_25679,N_25621);
nor U25901 (N_25901,N_25573,N_25780);
and U25902 (N_25902,N_25778,N_25686);
nand U25903 (N_25903,N_25756,N_25537);
and U25904 (N_25904,N_25788,N_25646);
nor U25905 (N_25905,N_25670,N_25738);
xor U25906 (N_25906,N_25667,N_25530);
nor U25907 (N_25907,N_25602,N_25579);
nand U25908 (N_25908,N_25790,N_25553);
nand U25909 (N_25909,N_25612,N_25605);
nor U25910 (N_25910,N_25611,N_25609);
xor U25911 (N_25911,N_25720,N_25764);
and U25912 (N_25912,N_25533,N_25696);
or U25913 (N_25913,N_25623,N_25588);
xor U25914 (N_25914,N_25655,N_25675);
nand U25915 (N_25915,N_25740,N_25531);
nand U25916 (N_25916,N_25549,N_25593);
or U25917 (N_25917,N_25550,N_25576);
or U25918 (N_25918,N_25704,N_25540);
xor U25919 (N_25919,N_25591,N_25673);
nand U25920 (N_25920,N_25552,N_25643);
or U25921 (N_25921,N_25598,N_25684);
nand U25922 (N_25922,N_25560,N_25603);
nand U25923 (N_25923,N_25562,N_25690);
and U25924 (N_25924,N_25601,N_25775);
nand U25925 (N_25925,N_25604,N_25725);
nor U25926 (N_25926,N_25674,N_25752);
nand U25927 (N_25927,N_25731,N_25583);
or U25928 (N_25928,N_25727,N_25504);
xnor U25929 (N_25929,N_25586,N_25536);
or U25930 (N_25930,N_25698,N_25526);
xor U25931 (N_25931,N_25717,N_25660);
nor U25932 (N_25932,N_25795,N_25746);
and U25933 (N_25933,N_25546,N_25672);
and U25934 (N_25934,N_25638,N_25648);
or U25935 (N_25935,N_25730,N_25669);
nor U25936 (N_25936,N_25608,N_25574);
nor U25937 (N_25937,N_25527,N_25785);
nor U25938 (N_25938,N_25645,N_25692);
xnor U25939 (N_25939,N_25659,N_25513);
and U25940 (N_25940,N_25743,N_25776);
xor U25941 (N_25941,N_25671,N_25786);
or U25942 (N_25942,N_25627,N_25797);
and U25943 (N_25943,N_25656,N_25714);
and U25944 (N_25944,N_25687,N_25742);
xnor U25945 (N_25945,N_25592,N_25515);
xor U25946 (N_25946,N_25685,N_25606);
or U25947 (N_25947,N_25654,N_25773);
and U25948 (N_25948,N_25514,N_25761);
or U25949 (N_25949,N_25543,N_25694);
and U25950 (N_25950,N_25660,N_25670);
nor U25951 (N_25951,N_25617,N_25659);
and U25952 (N_25952,N_25525,N_25533);
nor U25953 (N_25953,N_25786,N_25689);
or U25954 (N_25954,N_25609,N_25665);
and U25955 (N_25955,N_25514,N_25645);
nor U25956 (N_25956,N_25550,N_25709);
nand U25957 (N_25957,N_25513,N_25504);
nor U25958 (N_25958,N_25617,N_25709);
nand U25959 (N_25959,N_25698,N_25502);
nand U25960 (N_25960,N_25607,N_25697);
xor U25961 (N_25961,N_25600,N_25540);
nor U25962 (N_25962,N_25723,N_25528);
and U25963 (N_25963,N_25640,N_25566);
xor U25964 (N_25964,N_25799,N_25672);
nor U25965 (N_25965,N_25682,N_25575);
and U25966 (N_25966,N_25744,N_25735);
and U25967 (N_25967,N_25548,N_25625);
or U25968 (N_25968,N_25737,N_25596);
nor U25969 (N_25969,N_25752,N_25745);
and U25970 (N_25970,N_25534,N_25592);
nand U25971 (N_25971,N_25638,N_25672);
and U25972 (N_25972,N_25723,N_25770);
and U25973 (N_25973,N_25683,N_25775);
or U25974 (N_25974,N_25611,N_25687);
nor U25975 (N_25975,N_25610,N_25542);
and U25976 (N_25976,N_25792,N_25671);
nand U25977 (N_25977,N_25624,N_25728);
xor U25978 (N_25978,N_25527,N_25620);
and U25979 (N_25979,N_25614,N_25703);
and U25980 (N_25980,N_25631,N_25717);
or U25981 (N_25981,N_25718,N_25668);
nor U25982 (N_25982,N_25645,N_25596);
xnor U25983 (N_25983,N_25663,N_25727);
and U25984 (N_25984,N_25603,N_25546);
and U25985 (N_25985,N_25612,N_25600);
nand U25986 (N_25986,N_25617,N_25673);
or U25987 (N_25987,N_25755,N_25555);
nand U25988 (N_25988,N_25504,N_25798);
and U25989 (N_25989,N_25794,N_25535);
xor U25990 (N_25990,N_25701,N_25692);
and U25991 (N_25991,N_25687,N_25615);
and U25992 (N_25992,N_25707,N_25651);
nand U25993 (N_25993,N_25655,N_25527);
nand U25994 (N_25994,N_25756,N_25571);
nand U25995 (N_25995,N_25648,N_25789);
nand U25996 (N_25996,N_25646,N_25577);
nand U25997 (N_25997,N_25513,N_25760);
nand U25998 (N_25998,N_25575,N_25744);
xor U25999 (N_25999,N_25649,N_25699);
nand U26000 (N_26000,N_25636,N_25759);
xor U26001 (N_26001,N_25734,N_25510);
nand U26002 (N_26002,N_25514,N_25698);
or U26003 (N_26003,N_25580,N_25781);
and U26004 (N_26004,N_25688,N_25564);
nor U26005 (N_26005,N_25625,N_25663);
xor U26006 (N_26006,N_25583,N_25588);
nand U26007 (N_26007,N_25613,N_25745);
and U26008 (N_26008,N_25643,N_25794);
nand U26009 (N_26009,N_25566,N_25638);
nor U26010 (N_26010,N_25554,N_25657);
xnor U26011 (N_26011,N_25618,N_25518);
and U26012 (N_26012,N_25546,N_25691);
nor U26013 (N_26013,N_25638,N_25761);
and U26014 (N_26014,N_25655,N_25587);
and U26015 (N_26015,N_25511,N_25716);
nand U26016 (N_26016,N_25748,N_25669);
nand U26017 (N_26017,N_25666,N_25610);
nand U26018 (N_26018,N_25596,N_25545);
xnor U26019 (N_26019,N_25760,N_25747);
xnor U26020 (N_26020,N_25585,N_25701);
nor U26021 (N_26021,N_25624,N_25657);
and U26022 (N_26022,N_25635,N_25659);
nor U26023 (N_26023,N_25590,N_25640);
nor U26024 (N_26024,N_25619,N_25726);
nand U26025 (N_26025,N_25755,N_25672);
and U26026 (N_26026,N_25523,N_25664);
xor U26027 (N_26027,N_25752,N_25684);
xnor U26028 (N_26028,N_25750,N_25577);
xor U26029 (N_26029,N_25770,N_25662);
or U26030 (N_26030,N_25705,N_25542);
xnor U26031 (N_26031,N_25610,N_25727);
or U26032 (N_26032,N_25640,N_25737);
or U26033 (N_26033,N_25748,N_25749);
xnor U26034 (N_26034,N_25518,N_25709);
and U26035 (N_26035,N_25739,N_25621);
nor U26036 (N_26036,N_25673,N_25598);
xor U26037 (N_26037,N_25512,N_25639);
nor U26038 (N_26038,N_25707,N_25706);
or U26039 (N_26039,N_25717,N_25734);
or U26040 (N_26040,N_25691,N_25627);
xnor U26041 (N_26041,N_25741,N_25598);
or U26042 (N_26042,N_25736,N_25606);
nand U26043 (N_26043,N_25597,N_25769);
and U26044 (N_26044,N_25568,N_25642);
nand U26045 (N_26045,N_25751,N_25544);
xnor U26046 (N_26046,N_25621,N_25719);
or U26047 (N_26047,N_25503,N_25570);
and U26048 (N_26048,N_25606,N_25675);
nor U26049 (N_26049,N_25734,N_25543);
nor U26050 (N_26050,N_25553,N_25682);
nand U26051 (N_26051,N_25522,N_25787);
xor U26052 (N_26052,N_25591,N_25778);
nor U26053 (N_26053,N_25587,N_25733);
or U26054 (N_26054,N_25776,N_25714);
or U26055 (N_26055,N_25745,N_25751);
or U26056 (N_26056,N_25515,N_25552);
nand U26057 (N_26057,N_25673,N_25503);
nor U26058 (N_26058,N_25742,N_25766);
nor U26059 (N_26059,N_25630,N_25595);
nand U26060 (N_26060,N_25686,N_25547);
nand U26061 (N_26061,N_25603,N_25660);
and U26062 (N_26062,N_25584,N_25757);
and U26063 (N_26063,N_25673,N_25621);
nor U26064 (N_26064,N_25732,N_25518);
xnor U26065 (N_26065,N_25658,N_25522);
xor U26066 (N_26066,N_25716,N_25577);
and U26067 (N_26067,N_25703,N_25546);
nand U26068 (N_26068,N_25548,N_25750);
or U26069 (N_26069,N_25748,N_25790);
xor U26070 (N_26070,N_25615,N_25609);
xnor U26071 (N_26071,N_25679,N_25580);
or U26072 (N_26072,N_25519,N_25632);
nand U26073 (N_26073,N_25783,N_25503);
and U26074 (N_26074,N_25597,N_25636);
or U26075 (N_26075,N_25652,N_25665);
or U26076 (N_26076,N_25668,N_25764);
and U26077 (N_26077,N_25551,N_25517);
or U26078 (N_26078,N_25625,N_25629);
and U26079 (N_26079,N_25731,N_25569);
xor U26080 (N_26080,N_25510,N_25712);
or U26081 (N_26081,N_25679,N_25615);
nor U26082 (N_26082,N_25590,N_25708);
nand U26083 (N_26083,N_25685,N_25738);
nor U26084 (N_26084,N_25558,N_25727);
or U26085 (N_26085,N_25665,N_25798);
and U26086 (N_26086,N_25773,N_25645);
and U26087 (N_26087,N_25527,N_25730);
xnor U26088 (N_26088,N_25782,N_25741);
xor U26089 (N_26089,N_25587,N_25660);
xnor U26090 (N_26090,N_25607,N_25654);
xor U26091 (N_26091,N_25669,N_25519);
nand U26092 (N_26092,N_25565,N_25742);
xnor U26093 (N_26093,N_25650,N_25719);
and U26094 (N_26094,N_25711,N_25772);
nor U26095 (N_26095,N_25764,N_25651);
nor U26096 (N_26096,N_25678,N_25634);
nand U26097 (N_26097,N_25576,N_25540);
and U26098 (N_26098,N_25662,N_25554);
and U26099 (N_26099,N_25662,N_25732);
nand U26100 (N_26100,N_25937,N_25824);
or U26101 (N_26101,N_25988,N_25875);
xor U26102 (N_26102,N_25996,N_26083);
nand U26103 (N_26103,N_25971,N_25999);
nor U26104 (N_26104,N_25991,N_25980);
nand U26105 (N_26105,N_25908,N_26012);
nor U26106 (N_26106,N_25965,N_25821);
xnor U26107 (N_26107,N_26095,N_26059);
or U26108 (N_26108,N_25863,N_25859);
and U26109 (N_26109,N_25861,N_25833);
nand U26110 (N_26110,N_25928,N_26098);
nand U26111 (N_26111,N_25939,N_25993);
xnor U26112 (N_26112,N_26081,N_25855);
or U26113 (N_26113,N_26013,N_25942);
nand U26114 (N_26114,N_25818,N_25817);
nand U26115 (N_26115,N_25872,N_25998);
nor U26116 (N_26116,N_25843,N_26023);
or U26117 (N_26117,N_25829,N_26011);
and U26118 (N_26118,N_26033,N_25840);
nand U26119 (N_26119,N_25889,N_25888);
or U26120 (N_26120,N_25860,N_25894);
nor U26121 (N_26121,N_25816,N_25952);
xor U26122 (N_26122,N_25954,N_26064);
or U26123 (N_26123,N_26019,N_25809);
xnor U26124 (N_26124,N_26062,N_25835);
xor U26125 (N_26125,N_25885,N_26089);
nor U26126 (N_26126,N_25807,N_26021);
xnor U26127 (N_26127,N_26053,N_26007);
nor U26128 (N_26128,N_25883,N_25997);
or U26129 (N_26129,N_25819,N_25950);
nor U26130 (N_26130,N_25850,N_26017);
and U26131 (N_26131,N_25839,N_26061);
or U26132 (N_26132,N_25903,N_25895);
nor U26133 (N_26133,N_25909,N_26027);
xor U26134 (N_26134,N_25813,N_26009);
xnor U26135 (N_26135,N_25944,N_25825);
nand U26136 (N_26136,N_25880,N_25827);
nand U26137 (N_26137,N_26055,N_25987);
or U26138 (N_26138,N_25832,N_25931);
and U26139 (N_26139,N_25815,N_25856);
or U26140 (N_26140,N_26047,N_25905);
nor U26141 (N_26141,N_26058,N_26066);
or U26142 (N_26142,N_25834,N_25904);
nand U26143 (N_26143,N_26020,N_26096);
xnor U26144 (N_26144,N_25984,N_25989);
xnor U26145 (N_26145,N_25837,N_25922);
nor U26146 (N_26146,N_25853,N_25878);
xor U26147 (N_26147,N_26092,N_25990);
or U26148 (N_26148,N_26088,N_25854);
and U26149 (N_26149,N_25844,N_26090);
xor U26150 (N_26150,N_26028,N_25977);
or U26151 (N_26151,N_26016,N_26078);
and U26152 (N_26152,N_25890,N_26038);
nand U26153 (N_26153,N_25830,N_25929);
nor U26154 (N_26154,N_25899,N_26094);
nor U26155 (N_26155,N_26082,N_26071);
or U26156 (N_26156,N_25882,N_25900);
xnor U26157 (N_26157,N_26050,N_25934);
or U26158 (N_26158,N_26025,N_26070);
nor U26159 (N_26159,N_26076,N_25933);
nand U26160 (N_26160,N_26046,N_25935);
or U26161 (N_26161,N_26030,N_25969);
nor U26162 (N_26162,N_25841,N_25892);
or U26163 (N_26163,N_25992,N_25828);
nor U26164 (N_26164,N_26035,N_25955);
or U26165 (N_26165,N_25858,N_26093);
and U26166 (N_26166,N_25823,N_25930);
xor U26167 (N_26167,N_26068,N_25964);
xnor U26168 (N_26168,N_25936,N_25985);
nand U26169 (N_26169,N_26008,N_26005);
or U26170 (N_26170,N_26042,N_26080);
nand U26171 (N_26171,N_25917,N_25960);
and U26172 (N_26172,N_25868,N_26073);
nor U26173 (N_26173,N_26039,N_25877);
xnor U26174 (N_26174,N_26051,N_25864);
nand U26175 (N_26175,N_26037,N_26034);
or U26176 (N_26176,N_25804,N_25962);
xor U26177 (N_26177,N_26043,N_25921);
or U26178 (N_26178,N_25876,N_25994);
nand U26179 (N_26179,N_25978,N_25947);
xnor U26180 (N_26180,N_25867,N_25970);
and U26181 (N_26181,N_25891,N_26000);
nor U26182 (N_26182,N_26014,N_25949);
nor U26183 (N_26183,N_26079,N_25846);
and U26184 (N_26184,N_25842,N_26084);
xor U26185 (N_26185,N_25886,N_25924);
nor U26186 (N_26186,N_25948,N_25956);
or U26187 (N_26187,N_25848,N_25958);
and U26188 (N_26188,N_25851,N_26087);
nor U26189 (N_26189,N_25981,N_26048);
xor U26190 (N_26190,N_25983,N_26018);
and U26191 (N_26191,N_25866,N_26003);
nor U26192 (N_26192,N_25943,N_26065);
or U26193 (N_26193,N_26091,N_25906);
or U26194 (N_26194,N_25914,N_26004);
nand U26195 (N_26195,N_26060,N_25975);
xor U26196 (N_26196,N_25812,N_25826);
xor U26197 (N_26197,N_26067,N_25995);
nand U26198 (N_26198,N_26029,N_25814);
and U26199 (N_26199,N_25820,N_25811);
xor U26200 (N_26200,N_26069,N_25966);
xnor U26201 (N_26201,N_26045,N_25822);
or U26202 (N_26202,N_25808,N_25927);
nor U26203 (N_26203,N_25902,N_26006);
and U26204 (N_26204,N_25869,N_26022);
nor U26205 (N_26205,N_25865,N_25801);
xnor U26206 (N_26206,N_25957,N_25862);
nor U26207 (N_26207,N_25831,N_26049);
nand U26208 (N_26208,N_25896,N_25884);
and U26209 (N_26209,N_25881,N_25923);
or U26210 (N_26210,N_25845,N_26001);
or U26211 (N_26211,N_25920,N_25959);
xnor U26212 (N_26212,N_25926,N_26086);
xnor U26213 (N_26213,N_25918,N_25836);
nor U26214 (N_26214,N_26056,N_26085);
nand U26215 (N_26215,N_25951,N_25961);
nand U26216 (N_26216,N_26036,N_25873);
xor U26217 (N_26217,N_25913,N_25972);
nor U26218 (N_26218,N_25919,N_25916);
and U26219 (N_26219,N_25870,N_26032);
and U26220 (N_26220,N_25800,N_25847);
and U26221 (N_26221,N_26024,N_26041);
and U26222 (N_26222,N_25879,N_26040);
nand U26223 (N_26223,N_25940,N_25946);
xor U26224 (N_26224,N_26002,N_26099);
nor U26225 (N_26225,N_25838,N_25945);
and U26226 (N_26226,N_26015,N_25967);
nor U26227 (N_26227,N_26077,N_25986);
or U26228 (N_26228,N_25852,N_25806);
nand U26229 (N_26229,N_25874,N_26031);
nor U26230 (N_26230,N_25974,N_25805);
or U26231 (N_26231,N_25976,N_26072);
nor U26232 (N_26232,N_25907,N_25803);
or U26233 (N_26233,N_25849,N_26063);
nand U26234 (N_26234,N_26074,N_26054);
or U26235 (N_26235,N_25973,N_25898);
nor U26236 (N_26236,N_26097,N_26075);
nor U26237 (N_26237,N_25963,N_25915);
or U26238 (N_26238,N_25802,N_25932);
nor U26239 (N_26239,N_25968,N_26010);
nor U26240 (N_26240,N_26026,N_25910);
nor U26241 (N_26241,N_25953,N_25938);
or U26242 (N_26242,N_25871,N_25857);
or U26243 (N_26243,N_25810,N_25893);
nor U26244 (N_26244,N_25982,N_25901);
nor U26245 (N_26245,N_25887,N_26052);
and U26246 (N_26246,N_25925,N_26057);
xnor U26247 (N_26247,N_25897,N_26044);
and U26248 (N_26248,N_25941,N_25912);
nor U26249 (N_26249,N_25979,N_25911);
xor U26250 (N_26250,N_25960,N_26015);
nor U26251 (N_26251,N_25873,N_26016);
nor U26252 (N_26252,N_25898,N_25919);
nor U26253 (N_26253,N_25887,N_25961);
or U26254 (N_26254,N_25925,N_25984);
and U26255 (N_26255,N_25816,N_26016);
nand U26256 (N_26256,N_25862,N_25813);
nor U26257 (N_26257,N_25979,N_25813);
or U26258 (N_26258,N_26026,N_25854);
xnor U26259 (N_26259,N_25866,N_25804);
nor U26260 (N_26260,N_25879,N_26029);
xor U26261 (N_26261,N_25826,N_25806);
nand U26262 (N_26262,N_26072,N_25966);
xor U26263 (N_26263,N_26091,N_25930);
nand U26264 (N_26264,N_26022,N_25820);
xnor U26265 (N_26265,N_25829,N_25928);
nor U26266 (N_26266,N_25834,N_25913);
and U26267 (N_26267,N_25837,N_25914);
and U26268 (N_26268,N_25818,N_25859);
nand U26269 (N_26269,N_26013,N_26096);
or U26270 (N_26270,N_25865,N_25821);
nand U26271 (N_26271,N_25873,N_25900);
nor U26272 (N_26272,N_26088,N_26052);
nand U26273 (N_26273,N_25930,N_25998);
nor U26274 (N_26274,N_26052,N_26070);
nor U26275 (N_26275,N_25831,N_25877);
xor U26276 (N_26276,N_26017,N_25905);
or U26277 (N_26277,N_25992,N_26073);
nor U26278 (N_26278,N_25923,N_26096);
nor U26279 (N_26279,N_26072,N_25996);
nor U26280 (N_26280,N_25977,N_25886);
nor U26281 (N_26281,N_25868,N_26085);
and U26282 (N_26282,N_25838,N_25804);
xnor U26283 (N_26283,N_25879,N_25986);
or U26284 (N_26284,N_25906,N_25802);
nor U26285 (N_26285,N_25807,N_25861);
or U26286 (N_26286,N_26054,N_25941);
nand U26287 (N_26287,N_25973,N_26040);
and U26288 (N_26288,N_26046,N_26052);
nand U26289 (N_26289,N_25912,N_26009);
nand U26290 (N_26290,N_25870,N_25893);
nand U26291 (N_26291,N_25820,N_26025);
nor U26292 (N_26292,N_26034,N_25942);
nand U26293 (N_26293,N_25985,N_26004);
xnor U26294 (N_26294,N_26061,N_26034);
nor U26295 (N_26295,N_25983,N_26097);
and U26296 (N_26296,N_25984,N_25906);
and U26297 (N_26297,N_25936,N_25931);
or U26298 (N_26298,N_26087,N_25815);
xnor U26299 (N_26299,N_26073,N_26011);
nor U26300 (N_26300,N_25825,N_25937);
nor U26301 (N_26301,N_25926,N_26001);
nand U26302 (N_26302,N_25964,N_25930);
nand U26303 (N_26303,N_25963,N_25811);
xnor U26304 (N_26304,N_25825,N_26025);
xnor U26305 (N_26305,N_26089,N_25838);
and U26306 (N_26306,N_25879,N_25864);
nor U26307 (N_26307,N_25944,N_25933);
nand U26308 (N_26308,N_25812,N_25904);
xor U26309 (N_26309,N_25993,N_25830);
and U26310 (N_26310,N_26040,N_26028);
or U26311 (N_26311,N_26018,N_25828);
and U26312 (N_26312,N_25924,N_26085);
nand U26313 (N_26313,N_26077,N_25879);
xnor U26314 (N_26314,N_25925,N_25819);
or U26315 (N_26315,N_25827,N_25862);
xnor U26316 (N_26316,N_25951,N_25956);
nor U26317 (N_26317,N_25816,N_26024);
xnor U26318 (N_26318,N_25824,N_25805);
nand U26319 (N_26319,N_25905,N_25926);
or U26320 (N_26320,N_26058,N_26061);
xor U26321 (N_26321,N_25870,N_26060);
nor U26322 (N_26322,N_25823,N_25975);
nor U26323 (N_26323,N_26038,N_26095);
or U26324 (N_26324,N_26016,N_26044);
and U26325 (N_26325,N_25848,N_25824);
or U26326 (N_26326,N_25923,N_25892);
or U26327 (N_26327,N_25914,N_26069);
and U26328 (N_26328,N_25945,N_25910);
or U26329 (N_26329,N_25996,N_25868);
xor U26330 (N_26330,N_25949,N_25842);
or U26331 (N_26331,N_25804,N_25916);
or U26332 (N_26332,N_25855,N_25893);
xor U26333 (N_26333,N_25972,N_25925);
nor U26334 (N_26334,N_25879,N_25998);
and U26335 (N_26335,N_25913,N_25892);
nand U26336 (N_26336,N_25850,N_26006);
or U26337 (N_26337,N_25886,N_25939);
nand U26338 (N_26338,N_26058,N_25860);
xor U26339 (N_26339,N_25916,N_26098);
nor U26340 (N_26340,N_25802,N_26026);
nor U26341 (N_26341,N_25852,N_25979);
and U26342 (N_26342,N_25873,N_26097);
or U26343 (N_26343,N_25808,N_26046);
xnor U26344 (N_26344,N_25971,N_25913);
xnor U26345 (N_26345,N_25949,N_25856);
or U26346 (N_26346,N_26088,N_25848);
nand U26347 (N_26347,N_25883,N_25831);
or U26348 (N_26348,N_25972,N_26094);
nor U26349 (N_26349,N_25810,N_25979);
xnor U26350 (N_26350,N_25979,N_26033);
or U26351 (N_26351,N_26001,N_26069);
nor U26352 (N_26352,N_26005,N_25989);
xnor U26353 (N_26353,N_26081,N_25832);
xnor U26354 (N_26354,N_25871,N_25831);
xor U26355 (N_26355,N_25941,N_26084);
or U26356 (N_26356,N_25916,N_25985);
nand U26357 (N_26357,N_25986,N_25842);
xor U26358 (N_26358,N_25925,N_25968);
nand U26359 (N_26359,N_25944,N_26099);
xnor U26360 (N_26360,N_25875,N_25955);
and U26361 (N_26361,N_25992,N_25800);
xnor U26362 (N_26362,N_26037,N_25827);
nor U26363 (N_26363,N_25929,N_25910);
and U26364 (N_26364,N_25853,N_25934);
nand U26365 (N_26365,N_26084,N_26069);
or U26366 (N_26366,N_25809,N_26050);
or U26367 (N_26367,N_25835,N_26032);
and U26368 (N_26368,N_26028,N_25935);
nor U26369 (N_26369,N_25995,N_25971);
and U26370 (N_26370,N_26026,N_26021);
or U26371 (N_26371,N_25829,N_26038);
nand U26372 (N_26372,N_25995,N_26055);
nand U26373 (N_26373,N_25999,N_26085);
nand U26374 (N_26374,N_26057,N_26084);
or U26375 (N_26375,N_26070,N_25907);
or U26376 (N_26376,N_26073,N_26059);
nand U26377 (N_26377,N_25800,N_25994);
xnor U26378 (N_26378,N_26095,N_26037);
and U26379 (N_26379,N_25895,N_25910);
and U26380 (N_26380,N_25929,N_25961);
xnor U26381 (N_26381,N_25874,N_25854);
xnor U26382 (N_26382,N_26009,N_25843);
or U26383 (N_26383,N_25983,N_26079);
xnor U26384 (N_26384,N_26024,N_25811);
and U26385 (N_26385,N_25825,N_25813);
or U26386 (N_26386,N_25886,N_26035);
or U26387 (N_26387,N_25896,N_25930);
or U26388 (N_26388,N_25955,N_26010);
xnor U26389 (N_26389,N_25843,N_25958);
or U26390 (N_26390,N_25936,N_25959);
nand U26391 (N_26391,N_25864,N_25925);
or U26392 (N_26392,N_26036,N_26050);
or U26393 (N_26393,N_25986,N_26092);
nor U26394 (N_26394,N_25872,N_25921);
nor U26395 (N_26395,N_25822,N_25986);
or U26396 (N_26396,N_25992,N_25926);
or U26397 (N_26397,N_25915,N_25824);
xnor U26398 (N_26398,N_26042,N_26014);
or U26399 (N_26399,N_26096,N_25813);
nor U26400 (N_26400,N_26329,N_26283);
nand U26401 (N_26401,N_26270,N_26193);
xnor U26402 (N_26402,N_26117,N_26327);
and U26403 (N_26403,N_26299,N_26142);
or U26404 (N_26404,N_26189,N_26379);
nand U26405 (N_26405,N_26368,N_26268);
and U26406 (N_26406,N_26348,N_26230);
nand U26407 (N_26407,N_26337,N_26304);
nor U26408 (N_26408,N_26285,N_26108);
nand U26409 (N_26409,N_26264,N_26201);
nand U26410 (N_26410,N_26224,N_26282);
nand U26411 (N_26411,N_26152,N_26373);
or U26412 (N_26412,N_26111,N_26202);
and U26413 (N_26413,N_26226,N_26353);
or U26414 (N_26414,N_26294,N_26265);
or U26415 (N_26415,N_26123,N_26266);
xnor U26416 (N_26416,N_26138,N_26127);
or U26417 (N_26417,N_26100,N_26206);
nand U26418 (N_26418,N_26109,N_26252);
xnor U26419 (N_26419,N_26197,N_26317);
and U26420 (N_26420,N_26351,N_26258);
or U26421 (N_26421,N_26306,N_26195);
xor U26422 (N_26422,N_26228,N_26112);
xor U26423 (N_26423,N_26238,N_26380);
or U26424 (N_26424,N_26219,N_26101);
and U26425 (N_26425,N_26166,N_26326);
and U26426 (N_26426,N_26345,N_26204);
nor U26427 (N_26427,N_26180,N_26393);
nand U26428 (N_26428,N_26169,N_26144);
nand U26429 (N_26429,N_26274,N_26280);
xor U26430 (N_26430,N_26316,N_26208);
and U26431 (N_26431,N_26172,N_26135);
xor U26432 (N_26432,N_26207,N_26239);
or U26433 (N_26433,N_26328,N_26263);
and U26434 (N_26434,N_26255,N_26154);
xnor U26435 (N_26435,N_26205,N_26365);
xnor U26436 (N_26436,N_26250,N_26384);
nand U26437 (N_26437,N_26156,N_26107);
nand U26438 (N_26438,N_26211,N_26179);
nand U26439 (N_26439,N_26159,N_26126);
nor U26440 (N_26440,N_26158,N_26289);
and U26441 (N_26441,N_26129,N_26363);
or U26442 (N_26442,N_26340,N_26305);
nand U26443 (N_26443,N_26286,N_26291);
or U26444 (N_26444,N_26315,N_26114);
or U26445 (N_26445,N_26387,N_26355);
nor U26446 (N_26446,N_26352,N_26161);
and U26447 (N_26447,N_26377,N_26281);
xor U26448 (N_26448,N_26385,N_26396);
and U26449 (N_26449,N_26394,N_26339);
nor U26450 (N_26450,N_26350,N_26243);
xor U26451 (N_26451,N_26343,N_26139);
nor U26452 (N_26452,N_26370,N_26336);
and U26453 (N_26453,N_26269,N_26342);
and U26454 (N_26454,N_26257,N_26149);
nand U26455 (N_26455,N_26235,N_26216);
nor U26456 (N_26456,N_26386,N_26165);
nand U26457 (N_26457,N_26130,N_26227);
or U26458 (N_26458,N_26120,N_26300);
nand U26459 (N_26459,N_26332,N_26236);
xnor U26460 (N_26460,N_26381,N_26390);
nand U26461 (N_26461,N_26296,N_26247);
nand U26462 (N_26462,N_26190,N_26176);
or U26463 (N_26463,N_26178,N_26356);
or U26464 (N_26464,N_26290,N_26273);
nand U26465 (N_26465,N_26311,N_26322);
nor U26466 (N_26466,N_26103,N_26210);
nor U26467 (N_26467,N_26184,N_26200);
xnor U26468 (N_26468,N_26256,N_26106);
xnor U26469 (N_26469,N_26199,N_26369);
nor U26470 (N_26470,N_26367,N_26301);
nand U26471 (N_26471,N_26338,N_26128);
nor U26472 (N_26472,N_26341,N_26347);
nand U26473 (N_26473,N_26260,N_26163);
nor U26474 (N_26474,N_26398,N_26209);
nand U26475 (N_26475,N_26143,N_26122);
and U26476 (N_26476,N_26171,N_26335);
xnor U26477 (N_26477,N_26191,N_26357);
nand U26478 (N_26478,N_26222,N_26362);
or U26479 (N_26479,N_26364,N_26225);
nand U26480 (N_26480,N_26392,N_26221);
nand U26481 (N_26481,N_26254,N_26371);
xor U26482 (N_26482,N_26147,N_26359);
and U26483 (N_26483,N_26253,N_26249);
and U26484 (N_26484,N_26131,N_26366);
nand U26485 (N_26485,N_26185,N_26383);
nor U26486 (N_26486,N_26344,N_26167);
nand U26487 (N_26487,N_26153,N_26113);
nand U26488 (N_26488,N_26220,N_26244);
or U26489 (N_26489,N_26374,N_26376);
or U26490 (N_26490,N_26276,N_26312);
nor U26491 (N_26491,N_26331,N_26325);
xnor U26492 (N_26492,N_26375,N_26309);
and U26493 (N_26493,N_26170,N_26214);
xnor U26494 (N_26494,N_26125,N_26203);
nand U26495 (N_26495,N_26110,N_26251);
xnor U26496 (N_26496,N_26118,N_26292);
xnor U26497 (N_26497,N_26245,N_26324);
xnor U26498 (N_26498,N_26105,N_26173);
or U26499 (N_26499,N_26272,N_26288);
nand U26500 (N_26500,N_26246,N_26174);
nand U26501 (N_26501,N_26194,N_26164);
nand U26502 (N_26502,N_26104,N_26115);
nor U26503 (N_26503,N_26186,N_26229);
xor U26504 (N_26504,N_26183,N_26102);
or U26505 (N_26505,N_26287,N_26313);
or U26506 (N_26506,N_26241,N_26218);
or U26507 (N_26507,N_26389,N_26358);
nand U26508 (N_26508,N_26136,N_26133);
xnor U26509 (N_26509,N_26217,N_26297);
nand U26510 (N_26510,N_26399,N_26162);
or U26511 (N_26511,N_26334,N_26132);
nor U26512 (N_26512,N_26275,N_26215);
nor U26513 (N_26513,N_26196,N_26354);
and U26514 (N_26514,N_26278,N_26168);
xor U26515 (N_26515,N_26279,N_26372);
or U26516 (N_26516,N_26175,N_26323);
nor U26517 (N_26517,N_26124,N_26177);
or U26518 (N_26518,N_26308,N_26314);
xnor U26519 (N_26519,N_26223,N_26240);
and U26520 (N_26520,N_26333,N_26391);
xor U26521 (N_26521,N_26267,N_26187);
or U26522 (N_26522,N_26157,N_26382);
nand U26523 (N_26523,N_26192,N_26295);
and U26524 (N_26524,N_26140,N_26134);
nand U26525 (N_26525,N_26188,N_26284);
or U26526 (N_26526,N_26119,N_26198);
xor U26527 (N_26527,N_26148,N_26141);
xnor U26528 (N_26528,N_26303,N_26160);
xnor U26529 (N_26529,N_26145,N_26262);
or U26530 (N_26530,N_26307,N_26310);
and U26531 (N_26531,N_26234,N_26277);
or U26532 (N_26532,N_26121,N_26232);
and U26533 (N_26533,N_26397,N_26378);
and U26534 (N_26534,N_26182,N_26212);
and U26535 (N_26535,N_26320,N_26233);
or U26536 (N_26536,N_26231,N_26388);
xor U26537 (N_26537,N_26261,N_26321);
nand U26538 (N_26538,N_26349,N_26213);
nor U26539 (N_26539,N_26318,N_26330);
or U26540 (N_26540,N_26248,N_26181);
nand U26541 (N_26541,N_26242,N_26155);
and U26542 (N_26542,N_26319,N_26346);
and U26543 (N_26543,N_26271,N_26395);
xnor U26544 (N_26544,N_26360,N_26259);
xor U26545 (N_26545,N_26298,N_26293);
nand U26546 (N_26546,N_26302,N_26361);
xnor U26547 (N_26547,N_26150,N_26151);
or U26548 (N_26548,N_26146,N_26137);
nand U26549 (N_26549,N_26116,N_26237);
xnor U26550 (N_26550,N_26183,N_26133);
or U26551 (N_26551,N_26180,N_26381);
and U26552 (N_26552,N_26330,N_26128);
xor U26553 (N_26553,N_26165,N_26265);
and U26554 (N_26554,N_26215,N_26120);
and U26555 (N_26555,N_26218,N_26272);
nor U26556 (N_26556,N_26374,N_26178);
nor U26557 (N_26557,N_26128,N_26141);
and U26558 (N_26558,N_26272,N_26332);
nand U26559 (N_26559,N_26294,N_26379);
and U26560 (N_26560,N_26339,N_26255);
or U26561 (N_26561,N_26186,N_26146);
and U26562 (N_26562,N_26188,N_26363);
nand U26563 (N_26563,N_26143,N_26328);
nand U26564 (N_26564,N_26365,N_26337);
nor U26565 (N_26565,N_26334,N_26169);
or U26566 (N_26566,N_26320,N_26147);
nor U26567 (N_26567,N_26251,N_26307);
xor U26568 (N_26568,N_26200,N_26134);
and U26569 (N_26569,N_26328,N_26142);
and U26570 (N_26570,N_26288,N_26274);
xor U26571 (N_26571,N_26187,N_26170);
or U26572 (N_26572,N_26193,N_26361);
nand U26573 (N_26573,N_26169,N_26126);
or U26574 (N_26574,N_26314,N_26262);
xnor U26575 (N_26575,N_26149,N_26397);
nor U26576 (N_26576,N_26309,N_26124);
or U26577 (N_26577,N_26136,N_26151);
nand U26578 (N_26578,N_26355,N_26384);
nor U26579 (N_26579,N_26296,N_26387);
xnor U26580 (N_26580,N_26209,N_26237);
and U26581 (N_26581,N_26266,N_26246);
nand U26582 (N_26582,N_26212,N_26140);
and U26583 (N_26583,N_26288,N_26214);
and U26584 (N_26584,N_26153,N_26148);
and U26585 (N_26585,N_26291,N_26130);
nand U26586 (N_26586,N_26374,N_26296);
xor U26587 (N_26587,N_26156,N_26342);
and U26588 (N_26588,N_26306,N_26279);
nand U26589 (N_26589,N_26124,N_26346);
or U26590 (N_26590,N_26152,N_26267);
and U26591 (N_26591,N_26198,N_26289);
and U26592 (N_26592,N_26103,N_26361);
xor U26593 (N_26593,N_26348,N_26321);
nor U26594 (N_26594,N_26104,N_26229);
xor U26595 (N_26595,N_26126,N_26151);
and U26596 (N_26596,N_26201,N_26234);
nand U26597 (N_26597,N_26243,N_26284);
and U26598 (N_26598,N_26271,N_26368);
or U26599 (N_26599,N_26168,N_26248);
nand U26600 (N_26600,N_26273,N_26387);
and U26601 (N_26601,N_26228,N_26281);
or U26602 (N_26602,N_26321,N_26391);
or U26603 (N_26603,N_26310,N_26189);
nor U26604 (N_26604,N_26221,N_26395);
xor U26605 (N_26605,N_26299,N_26202);
and U26606 (N_26606,N_26189,N_26176);
nand U26607 (N_26607,N_26353,N_26237);
and U26608 (N_26608,N_26250,N_26256);
or U26609 (N_26609,N_26135,N_26315);
nand U26610 (N_26610,N_26365,N_26155);
xor U26611 (N_26611,N_26320,N_26350);
xor U26612 (N_26612,N_26251,N_26291);
nor U26613 (N_26613,N_26289,N_26188);
nor U26614 (N_26614,N_26146,N_26319);
nand U26615 (N_26615,N_26190,N_26281);
nand U26616 (N_26616,N_26129,N_26218);
nor U26617 (N_26617,N_26328,N_26140);
xor U26618 (N_26618,N_26312,N_26262);
or U26619 (N_26619,N_26334,N_26299);
nor U26620 (N_26620,N_26258,N_26112);
or U26621 (N_26621,N_26293,N_26399);
and U26622 (N_26622,N_26390,N_26262);
or U26623 (N_26623,N_26297,N_26225);
nor U26624 (N_26624,N_26376,N_26238);
xnor U26625 (N_26625,N_26139,N_26163);
nor U26626 (N_26626,N_26212,N_26372);
or U26627 (N_26627,N_26148,N_26135);
or U26628 (N_26628,N_26202,N_26348);
or U26629 (N_26629,N_26202,N_26320);
xnor U26630 (N_26630,N_26109,N_26329);
xnor U26631 (N_26631,N_26167,N_26153);
or U26632 (N_26632,N_26185,N_26171);
nor U26633 (N_26633,N_26129,N_26337);
xnor U26634 (N_26634,N_26303,N_26214);
and U26635 (N_26635,N_26143,N_26173);
or U26636 (N_26636,N_26225,N_26195);
nand U26637 (N_26637,N_26224,N_26356);
xnor U26638 (N_26638,N_26205,N_26132);
xnor U26639 (N_26639,N_26137,N_26145);
nand U26640 (N_26640,N_26113,N_26368);
nand U26641 (N_26641,N_26145,N_26100);
nand U26642 (N_26642,N_26288,N_26150);
or U26643 (N_26643,N_26198,N_26342);
nand U26644 (N_26644,N_26106,N_26313);
nand U26645 (N_26645,N_26392,N_26126);
or U26646 (N_26646,N_26352,N_26360);
xor U26647 (N_26647,N_26214,N_26313);
or U26648 (N_26648,N_26303,N_26276);
and U26649 (N_26649,N_26242,N_26373);
xnor U26650 (N_26650,N_26320,N_26269);
or U26651 (N_26651,N_26207,N_26295);
nand U26652 (N_26652,N_26259,N_26179);
nand U26653 (N_26653,N_26157,N_26210);
nand U26654 (N_26654,N_26285,N_26213);
xnor U26655 (N_26655,N_26186,N_26250);
or U26656 (N_26656,N_26280,N_26358);
xor U26657 (N_26657,N_26152,N_26362);
nor U26658 (N_26658,N_26129,N_26311);
nor U26659 (N_26659,N_26315,N_26230);
nand U26660 (N_26660,N_26204,N_26397);
nand U26661 (N_26661,N_26381,N_26342);
nand U26662 (N_26662,N_26252,N_26245);
and U26663 (N_26663,N_26200,N_26168);
nor U26664 (N_26664,N_26295,N_26205);
xor U26665 (N_26665,N_26310,N_26393);
nand U26666 (N_26666,N_26160,N_26192);
or U26667 (N_26667,N_26108,N_26104);
nand U26668 (N_26668,N_26237,N_26184);
and U26669 (N_26669,N_26244,N_26225);
and U26670 (N_26670,N_26381,N_26307);
xor U26671 (N_26671,N_26340,N_26293);
or U26672 (N_26672,N_26103,N_26139);
xor U26673 (N_26673,N_26338,N_26329);
and U26674 (N_26674,N_26321,N_26349);
and U26675 (N_26675,N_26280,N_26134);
or U26676 (N_26676,N_26136,N_26372);
and U26677 (N_26677,N_26289,N_26212);
nand U26678 (N_26678,N_26340,N_26105);
nand U26679 (N_26679,N_26295,N_26144);
and U26680 (N_26680,N_26183,N_26223);
and U26681 (N_26681,N_26326,N_26198);
and U26682 (N_26682,N_26271,N_26350);
nand U26683 (N_26683,N_26119,N_26208);
xnor U26684 (N_26684,N_26265,N_26157);
or U26685 (N_26685,N_26248,N_26220);
nor U26686 (N_26686,N_26167,N_26300);
nand U26687 (N_26687,N_26140,N_26126);
nand U26688 (N_26688,N_26397,N_26367);
nand U26689 (N_26689,N_26352,N_26284);
and U26690 (N_26690,N_26240,N_26179);
and U26691 (N_26691,N_26385,N_26144);
nand U26692 (N_26692,N_26238,N_26215);
nor U26693 (N_26693,N_26168,N_26194);
xnor U26694 (N_26694,N_26352,N_26311);
and U26695 (N_26695,N_26242,N_26227);
nor U26696 (N_26696,N_26315,N_26327);
xnor U26697 (N_26697,N_26243,N_26332);
nand U26698 (N_26698,N_26172,N_26288);
nor U26699 (N_26699,N_26204,N_26234);
nor U26700 (N_26700,N_26505,N_26518);
nor U26701 (N_26701,N_26613,N_26438);
nand U26702 (N_26702,N_26523,N_26415);
nor U26703 (N_26703,N_26689,N_26685);
and U26704 (N_26704,N_26629,N_26677);
xnor U26705 (N_26705,N_26420,N_26434);
xor U26706 (N_26706,N_26541,N_26458);
or U26707 (N_26707,N_26565,N_26594);
nor U26708 (N_26708,N_26563,N_26609);
xnor U26709 (N_26709,N_26534,N_26479);
and U26710 (N_26710,N_26492,N_26513);
xnor U26711 (N_26711,N_26522,N_26580);
nand U26712 (N_26712,N_26448,N_26495);
nand U26713 (N_26713,N_26583,N_26519);
or U26714 (N_26714,N_26566,N_26570);
nor U26715 (N_26715,N_26516,N_26618);
nor U26716 (N_26716,N_26668,N_26533);
xnor U26717 (N_26717,N_26605,N_26512);
xnor U26718 (N_26718,N_26648,N_26494);
or U26719 (N_26719,N_26463,N_26453);
nor U26720 (N_26720,N_26590,N_26486);
nand U26721 (N_26721,N_26466,N_26536);
or U26722 (N_26722,N_26581,N_26699);
and U26723 (N_26723,N_26655,N_26558);
xnor U26724 (N_26724,N_26527,N_26633);
and U26725 (N_26725,N_26651,N_26496);
xnor U26726 (N_26726,N_26678,N_26411);
or U26727 (N_26727,N_26625,N_26674);
or U26728 (N_26728,N_26686,N_26446);
or U26729 (N_26729,N_26690,N_26639);
xnor U26730 (N_26730,N_26669,N_26661);
nor U26731 (N_26731,N_26607,N_26652);
or U26732 (N_26732,N_26454,N_26455);
or U26733 (N_26733,N_26464,N_26471);
nor U26734 (N_26734,N_26597,N_26680);
and U26735 (N_26735,N_26428,N_26535);
nor U26736 (N_26736,N_26621,N_26435);
or U26737 (N_26737,N_26600,N_26402);
and U26738 (N_26738,N_26632,N_26620);
xnor U26739 (N_26739,N_26426,N_26596);
and U26740 (N_26740,N_26520,N_26645);
nand U26741 (N_26741,N_26490,N_26449);
nand U26742 (N_26742,N_26582,N_26658);
nor U26743 (N_26743,N_26672,N_26441);
or U26744 (N_26744,N_26663,N_26646);
xnor U26745 (N_26745,N_26657,N_26493);
nor U26746 (N_26746,N_26687,N_26511);
or U26747 (N_26747,N_26559,N_26691);
xnor U26748 (N_26748,N_26406,N_26456);
and U26749 (N_26749,N_26693,N_26514);
nand U26750 (N_26750,N_26548,N_26650);
and U26751 (N_26751,N_26575,N_26619);
xor U26752 (N_26752,N_26571,N_26465);
nand U26753 (N_26753,N_26653,N_26578);
or U26754 (N_26754,N_26612,N_26569);
nor U26755 (N_26755,N_26408,N_26637);
xnor U26756 (N_26756,N_26440,N_26521);
or U26757 (N_26757,N_26628,N_26615);
nand U26758 (N_26758,N_26662,N_26587);
nand U26759 (N_26759,N_26601,N_26537);
or U26760 (N_26760,N_26608,N_26547);
xnor U26761 (N_26761,N_26532,N_26427);
or U26762 (N_26762,N_26698,N_26515);
or U26763 (N_26763,N_26641,N_26546);
or U26764 (N_26764,N_26551,N_26526);
nand U26765 (N_26765,N_26660,N_26568);
and U26766 (N_26766,N_26598,N_26630);
xor U26767 (N_26767,N_26542,N_26412);
nand U26768 (N_26768,N_26553,N_26508);
or U26769 (N_26769,N_26517,N_26431);
and U26770 (N_26770,N_26606,N_26425);
nor U26771 (N_26771,N_26529,N_26550);
or U26772 (N_26772,N_26488,N_26401);
nand U26773 (N_26773,N_26627,N_26579);
xor U26774 (N_26774,N_26591,N_26631);
nand U26775 (N_26775,N_26642,N_26695);
or U26776 (N_26776,N_26475,N_26418);
nor U26777 (N_26777,N_26416,N_26675);
and U26778 (N_26778,N_26499,N_26483);
nor U26779 (N_26779,N_26502,N_26671);
nor U26780 (N_26780,N_26683,N_26429);
and U26781 (N_26781,N_26585,N_26626);
or U26782 (N_26782,N_26557,N_26450);
and U26783 (N_26783,N_26692,N_26422);
xor U26784 (N_26784,N_26457,N_26667);
nor U26785 (N_26785,N_26647,N_26424);
and U26786 (N_26786,N_26573,N_26610);
nand U26787 (N_26787,N_26497,N_26524);
nor U26788 (N_26788,N_26501,N_26567);
and U26789 (N_26789,N_26409,N_26577);
and U26790 (N_26790,N_26531,N_26697);
nor U26791 (N_26791,N_26696,N_26681);
and U26792 (N_26792,N_26472,N_26562);
or U26793 (N_26793,N_26623,N_26477);
and U26794 (N_26794,N_26649,N_26470);
nand U26795 (N_26795,N_26487,N_26476);
nand U26796 (N_26796,N_26407,N_26564);
nand U26797 (N_26797,N_26525,N_26554);
nor U26798 (N_26798,N_26589,N_26688);
xnor U26799 (N_26799,N_26643,N_26460);
and U26800 (N_26800,N_26481,N_26442);
xnor U26801 (N_26801,N_26538,N_26462);
or U26802 (N_26802,N_26436,N_26666);
or U26803 (N_26803,N_26510,N_26410);
and U26804 (N_26804,N_26572,N_26506);
xor U26805 (N_26805,N_26545,N_26640);
or U26806 (N_26806,N_26447,N_26588);
nand U26807 (N_26807,N_26540,N_26544);
xnor U26808 (N_26808,N_26694,N_26556);
or U26809 (N_26809,N_26430,N_26636);
and U26810 (N_26810,N_26480,N_26654);
and U26811 (N_26811,N_26445,N_26635);
xor U26812 (N_26812,N_26555,N_26676);
nor U26813 (N_26813,N_26530,N_26423);
or U26814 (N_26814,N_26638,N_26473);
nor U26815 (N_26815,N_26593,N_26414);
and U26816 (N_26816,N_26509,N_26421);
xor U26817 (N_26817,N_26659,N_26503);
xor U26818 (N_26818,N_26592,N_26439);
nor U26819 (N_26819,N_26586,N_26624);
nand U26820 (N_26820,N_26437,N_26498);
nor U26821 (N_26821,N_26507,N_26500);
and U26822 (N_26822,N_26417,N_26404);
xnor U26823 (N_26823,N_26603,N_26602);
or U26824 (N_26824,N_26413,N_26634);
xor U26825 (N_26825,N_26467,N_26644);
and U26826 (N_26826,N_26622,N_26468);
nand U26827 (N_26827,N_26539,N_26452);
or U26828 (N_26828,N_26482,N_26484);
xnor U26829 (N_26829,N_26616,N_26543);
xnor U26830 (N_26830,N_26611,N_26673);
nor U26831 (N_26831,N_26604,N_26528);
nor U26832 (N_26832,N_26682,N_26443);
or U26833 (N_26833,N_26403,N_26679);
xor U26834 (N_26834,N_26684,N_26451);
nand U26835 (N_26835,N_26400,N_26670);
nand U26836 (N_26836,N_26469,N_26489);
or U26837 (N_26837,N_26433,N_26561);
xor U26838 (N_26838,N_26664,N_26405);
nand U26839 (N_26839,N_26584,N_26432);
nor U26840 (N_26840,N_26576,N_26419);
or U26841 (N_26841,N_26656,N_26599);
or U26842 (N_26842,N_26617,N_26478);
or U26843 (N_26843,N_26461,N_26549);
nor U26844 (N_26844,N_26595,N_26459);
and U26845 (N_26845,N_26614,N_26574);
nand U26846 (N_26846,N_26485,N_26491);
or U26847 (N_26847,N_26560,N_26665);
nor U26848 (N_26848,N_26552,N_26474);
and U26849 (N_26849,N_26444,N_26504);
and U26850 (N_26850,N_26419,N_26551);
nor U26851 (N_26851,N_26641,N_26518);
nor U26852 (N_26852,N_26538,N_26456);
nand U26853 (N_26853,N_26439,N_26444);
or U26854 (N_26854,N_26503,N_26452);
nor U26855 (N_26855,N_26685,N_26618);
nor U26856 (N_26856,N_26479,N_26699);
xor U26857 (N_26857,N_26459,N_26416);
nand U26858 (N_26858,N_26660,N_26474);
nor U26859 (N_26859,N_26501,N_26672);
or U26860 (N_26860,N_26536,N_26619);
or U26861 (N_26861,N_26499,N_26635);
nand U26862 (N_26862,N_26434,N_26574);
nor U26863 (N_26863,N_26616,N_26430);
and U26864 (N_26864,N_26431,N_26562);
or U26865 (N_26865,N_26608,N_26415);
nand U26866 (N_26866,N_26639,N_26428);
nor U26867 (N_26867,N_26461,N_26587);
xnor U26868 (N_26868,N_26539,N_26492);
nand U26869 (N_26869,N_26428,N_26621);
nor U26870 (N_26870,N_26472,N_26627);
nand U26871 (N_26871,N_26476,N_26572);
or U26872 (N_26872,N_26575,N_26645);
xnor U26873 (N_26873,N_26583,N_26664);
xnor U26874 (N_26874,N_26690,N_26565);
nand U26875 (N_26875,N_26611,N_26539);
nand U26876 (N_26876,N_26521,N_26681);
and U26877 (N_26877,N_26443,N_26514);
or U26878 (N_26878,N_26495,N_26643);
xnor U26879 (N_26879,N_26679,N_26571);
or U26880 (N_26880,N_26613,N_26637);
xor U26881 (N_26881,N_26529,N_26455);
xnor U26882 (N_26882,N_26400,N_26499);
or U26883 (N_26883,N_26686,N_26605);
xor U26884 (N_26884,N_26409,N_26517);
xor U26885 (N_26885,N_26520,N_26478);
nor U26886 (N_26886,N_26621,N_26522);
nand U26887 (N_26887,N_26570,N_26643);
nor U26888 (N_26888,N_26576,N_26687);
nand U26889 (N_26889,N_26461,N_26646);
or U26890 (N_26890,N_26510,N_26579);
or U26891 (N_26891,N_26455,N_26592);
nand U26892 (N_26892,N_26637,N_26536);
nand U26893 (N_26893,N_26562,N_26646);
or U26894 (N_26894,N_26418,N_26517);
nor U26895 (N_26895,N_26688,N_26577);
nor U26896 (N_26896,N_26490,N_26624);
nor U26897 (N_26897,N_26482,N_26531);
nand U26898 (N_26898,N_26692,N_26446);
and U26899 (N_26899,N_26458,N_26607);
and U26900 (N_26900,N_26420,N_26438);
or U26901 (N_26901,N_26598,N_26509);
nor U26902 (N_26902,N_26696,N_26414);
and U26903 (N_26903,N_26637,N_26436);
xnor U26904 (N_26904,N_26612,N_26658);
or U26905 (N_26905,N_26639,N_26530);
nor U26906 (N_26906,N_26438,N_26433);
nor U26907 (N_26907,N_26478,N_26691);
and U26908 (N_26908,N_26442,N_26444);
and U26909 (N_26909,N_26513,N_26437);
nand U26910 (N_26910,N_26403,N_26454);
nand U26911 (N_26911,N_26592,N_26643);
and U26912 (N_26912,N_26405,N_26573);
or U26913 (N_26913,N_26503,N_26467);
nor U26914 (N_26914,N_26628,N_26524);
and U26915 (N_26915,N_26491,N_26422);
xor U26916 (N_26916,N_26483,N_26666);
xnor U26917 (N_26917,N_26410,N_26465);
xor U26918 (N_26918,N_26449,N_26578);
xor U26919 (N_26919,N_26490,N_26509);
or U26920 (N_26920,N_26462,N_26550);
nor U26921 (N_26921,N_26638,N_26439);
or U26922 (N_26922,N_26540,N_26631);
nand U26923 (N_26923,N_26599,N_26449);
and U26924 (N_26924,N_26530,N_26550);
and U26925 (N_26925,N_26531,N_26634);
or U26926 (N_26926,N_26613,N_26449);
and U26927 (N_26927,N_26455,N_26473);
nand U26928 (N_26928,N_26589,N_26423);
xnor U26929 (N_26929,N_26496,N_26677);
nor U26930 (N_26930,N_26578,N_26431);
xnor U26931 (N_26931,N_26483,N_26591);
or U26932 (N_26932,N_26597,N_26449);
or U26933 (N_26933,N_26626,N_26593);
and U26934 (N_26934,N_26669,N_26528);
and U26935 (N_26935,N_26456,N_26431);
or U26936 (N_26936,N_26544,N_26578);
and U26937 (N_26937,N_26580,N_26648);
or U26938 (N_26938,N_26618,N_26514);
xor U26939 (N_26939,N_26507,N_26402);
and U26940 (N_26940,N_26599,N_26576);
and U26941 (N_26941,N_26424,N_26518);
or U26942 (N_26942,N_26644,N_26620);
or U26943 (N_26943,N_26549,N_26667);
and U26944 (N_26944,N_26518,N_26451);
or U26945 (N_26945,N_26524,N_26618);
or U26946 (N_26946,N_26403,N_26584);
nand U26947 (N_26947,N_26410,N_26618);
and U26948 (N_26948,N_26687,N_26416);
and U26949 (N_26949,N_26699,N_26527);
nand U26950 (N_26950,N_26592,N_26585);
or U26951 (N_26951,N_26619,N_26405);
nor U26952 (N_26952,N_26578,N_26691);
xor U26953 (N_26953,N_26447,N_26651);
nand U26954 (N_26954,N_26516,N_26698);
and U26955 (N_26955,N_26405,N_26551);
nor U26956 (N_26956,N_26564,N_26452);
and U26957 (N_26957,N_26691,N_26491);
or U26958 (N_26958,N_26417,N_26541);
xnor U26959 (N_26959,N_26698,N_26567);
xnor U26960 (N_26960,N_26671,N_26565);
nor U26961 (N_26961,N_26612,N_26613);
nand U26962 (N_26962,N_26454,N_26443);
and U26963 (N_26963,N_26593,N_26493);
nor U26964 (N_26964,N_26505,N_26448);
xnor U26965 (N_26965,N_26549,N_26510);
or U26966 (N_26966,N_26532,N_26531);
or U26967 (N_26967,N_26424,N_26525);
nand U26968 (N_26968,N_26553,N_26482);
or U26969 (N_26969,N_26404,N_26604);
or U26970 (N_26970,N_26496,N_26658);
or U26971 (N_26971,N_26644,N_26473);
and U26972 (N_26972,N_26409,N_26435);
nand U26973 (N_26973,N_26448,N_26636);
xnor U26974 (N_26974,N_26408,N_26567);
nor U26975 (N_26975,N_26482,N_26570);
or U26976 (N_26976,N_26652,N_26634);
nor U26977 (N_26977,N_26459,N_26635);
and U26978 (N_26978,N_26637,N_26559);
nand U26979 (N_26979,N_26682,N_26526);
xnor U26980 (N_26980,N_26504,N_26616);
xor U26981 (N_26981,N_26628,N_26630);
nor U26982 (N_26982,N_26541,N_26539);
and U26983 (N_26983,N_26672,N_26442);
nand U26984 (N_26984,N_26400,N_26534);
xnor U26985 (N_26985,N_26643,N_26580);
or U26986 (N_26986,N_26505,N_26566);
or U26987 (N_26987,N_26426,N_26446);
or U26988 (N_26988,N_26559,N_26446);
nor U26989 (N_26989,N_26621,N_26659);
xnor U26990 (N_26990,N_26453,N_26630);
and U26991 (N_26991,N_26697,N_26601);
nand U26992 (N_26992,N_26578,N_26566);
xor U26993 (N_26993,N_26611,N_26663);
nor U26994 (N_26994,N_26425,N_26456);
xnor U26995 (N_26995,N_26639,N_26499);
or U26996 (N_26996,N_26611,N_26498);
or U26997 (N_26997,N_26610,N_26615);
xor U26998 (N_26998,N_26494,N_26514);
nor U26999 (N_26999,N_26652,N_26498);
nor U27000 (N_27000,N_26733,N_26934);
or U27001 (N_27001,N_26880,N_26728);
xnor U27002 (N_27002,N_26922,N_26736);
nor U27003 (N_27003,N_26890,N_26831);
xor U27004 (N_27004,N_26943,N_26755);
and U27005 (N_27005,N_26803,N_26832);
nand U27006 (N_27006,N_26778,N_26726);
and U27007 (N_27007,N_26779,N_26954);
and U27008 (N_27008,N_26788,N_26713);
nor U27009 (N_27009,N_26887,N_26798);
nor U27010 (N_27010,N_26907,N_26746);
and U27011 (N_27011,N_26870,N_26955);
and U27012 (N_27012,N_26795,N_26966);
and U27013 (N_27013,N_26792,N_26960);
nand U27014 (N_27014,N_26780,N_26867);
xor U27015 (N_27015,N_26701,N_26761);
and U27016 (N_27016,N_26857,N_26911);
xnor U27017 (N_27017,N_26808,N_26930);
or U27018 (N_27018,N_26744,N_26731);
or U27019 (N_27019,N_26716,N_26974);
or U27020 (N_27020,N_26709,N_26937);
or U27021 (N_27021,N_26727,N_26998);
and U27022 (N_27022,N_26711,N_26845);
and U27023 (N_27023,N_26723,N_26800);
nand U27024 (N_27024,N_26927,N_26988);
and U27025 (N_27025,N_26999,N_26908);
and U27026 (N_27026,N_26854,N_26707);
nor U27027 (N_27027,N_26962,N_26978);
nor U27028 (N_27028,N_26757,N_26799);
nand U27029 (N_27029,N_26714,N_26838);
nand U27030 (N_27030,N_26814,N_26985);
xnor U27031 (N_27031,N_26720,N_26920);
xor U27032 (N_27032,N_26722,N_26741);
xor U27033 (N_27033,N_26864,N_26817);
nand U27034 (N_27034,N_26902,N_26900);
nor U27035 (N_27035,N_26751,N_26967);
and U27036 (N_27036,N_26819,N_26730);
xor U27037 (N_27037,N_26840,N_26996);
nor U27038 (N_27038,N_26892,N_26929);
xnor U27039 (N_27039,N_26710,N_26956);
and U27040 (N_27040,N_26936,N_26823);
nand U27041 (N_27041,N_26993,N_26888);
and U27042 (N_27042,N_26771,N_26981);
or U27043 (N_27043,N_26853,N_26945);
nand U27044 (N_27044,N_26904,N_26891);
or U27045 (N_27045,N_26973,N_26878);
nand U27046 (N_27046,N_26813,N_26836);
nand U27047 (N_27047,N_26872,N_26980);
and U27048 (N_27048,N_26901,N_26903);
and U27049 (N_27049,N_26958,N_26706);
nor U27050 (N_27050,N_26790,N_26863);
and U27051 (N_27051,N_26932,N_26756);
nor U27052 (N_27052,N_26718,N_26747);
nor U27053 (N_27053,N_26841,N_26861);
nand U27054 (N_27054,N_26879,N_26961);
nand U27055 (N_27055,N_26989,N_26822);
nand U27056 (N_27056,N_26957,N_26804);
xnor U27057 (N_27057,N_26824,N_26812);
and U27058 (N_27058,N_26931,N_26772);
and U27059 (N_27059,N_26899,N_26940);
nand U27060 (N_27060,N_26862,N_26767);
or U27061 (N_27061,N_26721,N_26848);
xnor U27062 (N_27062,N_26882,N_26820);
or U27063 (N_27063,N_26933,N_26969);
or U27064 (N_27064,N_26830,N_26986);
and U27065 (N_27065,N_26770,N_26844);
xnor U27066 (N_27066,N_26918,N_26917);
xor U27067 (N_27067,N_26774,N_26732);
nor U27068 (N_27068,N_26811,N_26972);
and U27069 (N_27069,N_26827,N_26893);
nand U27070 (N_27070,N_26995,N_26758);
xor U27071 (N_27071,N_26729,N_26885);
nor U27072 (N_27072,N_26847,N_26786);
nor U27073 (N_27073,N_26971,N_26924);
xnor U27074 (N_27074,N_26717,N_26835);
or U27075 (N_27075,N_26963,N_26895);
nand U27076 (N_27076,N_26768,N_26821);
nor U27077 (N_27077,N_26737,N_26782);
or U27078 (N_27078,N_26865,N_26909);
or U27079 (N_27079,N_26944,N_26916);
or U27080 (N_27080,N_26816,N_26968);
or U27081 (N_27081,N_26898,N_26912);
nor U27082 (N_27082,N_26979,N_26760);
nor U27083 (N_27083,N_26914,N_26828);
and U27084 (N_27084,N_26785,N_26776);
nand U27085 (N_27085,N_26789,N_26941);
or U27086 (N_27086,N_26984,N_26705);
xor U27087 (N_27087,N_26869,N_26787);
nand U27088 (N_27088,N_26851,N_26873);
or U27089 (N_27089,N_26815,N_26951);
and U27090 (N_27090,N_26802,N_26915);
or U27091 (N_27091,N_26724,N_26715);
and U27092 (N_27092,N_26719,N_26976);
and U27093 (N_27093,N_26842,N_26807);
nand U27094 (N_27094,N_26777,N_26877);
nor U27095 (N_27095,N_26794,N_26990);
nand U27096 (N_27096,N_26743,N_26725);
and U27097 (N_27097,N_26742,N_26858);
nand U27098 (N_27098,N_26810,N_26910);
and U27099 (N_27099,N_26987,N_26806);
or U27100 (N_27100,N_26970,N_26837);
and U27101 (N_27101,N_26735,N_26991);
nand U27102 (N_27102,N_26745,N_26926);
nand U27103 (N_27103,N_26975,N_26773);
xor U27104 (N_27104,N_26818,N_26850);
or U27105 (N_27105,N_26781,N_26866);
nand U27106 (N_27106,N_26752,N_26843);
nor U27107 (N_27107,N_26754,N_26977);
or U27108 (N_27108,N_26894,N_26868);
or U27109 (N_27109,N_26938,N_26769);
nand U27110 (N_27110,N_26740,N_26905);
nand U27111 (N_27111,N_26708,N_26793);
and U27112 (N_27112,N_26791,N_26805);
or U27113 (N_27113,N_26849,N_26834);
nand U27114 (N_27114,N_26859,N_26919);
or U27115 (N_27115,N_26886,N_26856);
xor U27116 (N_27116,N_26750,N_26703);
xor U27117 (N_27117,N_26992,N_26826);
nor U27118 (N_27118,N_26734,N_26946);
or U27119 (N_27119,N_26738,N_26913);
nand U27120 (N_27120,N_26881,N_26748);
nor U27121 (N_27121,N_26852,N_26775);
xor U27122 (N_27122,N_26982,N_26925);
nand U27123 (N_27123,N_26889,N_26764);
and U27124 (N_27124,N_26876,N_26753);
or U27125 (N_27125,N_26923,N_26959);
and U27126 (N_27126,N_26801,N_26965);
or U27127 (N_27127,N_26875,N_26762);
and U27128 (N_27128,N_26947,N_26700);
or U27129 (N_27129,N_26846,N_26949);
nand U27130 (N_27130,N_26953,N_26874);
xor U27131 (N_27131,N_26759,N_26942);
and U27132 (N_27132,N_26994,N_26839);
nor U27133 (N_27133,N_26702,N_26829);
and U27134 (N_27134,N_26797,N_26809);
nand U27135 (N_27135,N_26935,N_26948);
xor U27136 (N_27136,N_26983,N_26766);
or U27137 (N_27137,N_26704,N_26883);
xnor U27138 (N_27138,N_26928,N_26884);
and U27139 (N_27139,N_26763,N_26939);
nand U27140 (N_27140,N_26739,N_26833);
nor U27141 (N_27141,N_26896,N_26897);
xnor U27142 (N_27142,N_26860,N_26783);
nand U27143 (N_27143,N_26964,N_26952);
nor U27144 (N_27144,N_26921,N_26855);
nand U27145 (N_27145,N_26749,N_26825);
nand U27146 (N_27146,N_26784,N_26906);
xor U27147 (N_27147,N_26950,N_26712);
nor U27148 (N_27148,N_26765,N_26796);
nand U27149 (N_27149,N_26871,N_26997);
nor U27150 (N_27150,N_26822,N_26934);
and U27151 (N_27151,N_26734,N_26752);
and U27152 (N_27152,N_26930,N_26924);
nor U27153 (N_27153,N_26836,N_26729);
nor U27154 (N_27154,N_26776,N_26855);
nand U27155 (N_27155,N_26756,N_26841);
or U27156 (N_27156,N_26848,N_26930);
xnor U27157 (N_27157,N_26881,N_26742);
and U27158 (N_27158,N_26939,N_26914);
nor U27159 (N_27159,N_26896,N_26808);
nand U27160 (N_27160,N_26879,N_26949);
nor U27161 (N_27161,N_26712,N_26902);
or U27162 (N_27162,N_26900,N_26978);
and U27163 (N_27163,N_26753,N_26910);
nor U27164 (N_27164,N_26999,N_26933);
xnor U27165 (N_27165,N_26779,N_26735);
or U27166 (N_27166,N_26758,N_26787);
nor U27167 (N_27167,N_26910,N_26969);
nor U27168 (N_27168,N_26977,N_26973);
xnor U27169 (N_27169,N_26824,N_26705);
and U27170 (N_27170,N_26786,N_26913);
nor U27171 (N_27171,N_26893,N_26808);
or U27172 (N_27172,N_26705,N_26729);
nand U27173 (N_27173,N_26935,N_26921);
xnor U27174 (N_27174,N_26981,N_26838);
xor U27175 (N_27175,N_26977,N_26873);
xor U27176 (N_27176,N_26981,N_26715);
nand U27177 (N_27177,N_26881,N_26735);
nor U27178 (N_27178,N_26974,N_26825);
nor U27179 (N_27179,N_26785,N_26927);
and U27180 (N_27180,N_26866,N_26930);
nor U27181 (N_27181,N_26899,N_26953);
nand U27182 (N_27182,N_26862,N_26713);
nand U27183 (N_27183,N_26906,N_26791);
and U27184 (N_27184,N_26875,N_26995);
xor U27185 (N_27185,N_26739,N_26707);
and U27186 (N_27186,N_26922,N_26802);
nand U27187 (N_27187,N_26824,N_26755);
nor U27188 (N_27188,N_26854,N_26814);
nor U27189 (N_27189,N_26886,N_26852);
and U27190 (N_27190,N_26731,N_26924);
nand U27191 (N_27191,N_26958,N_26996);
xnor U27192 (N_27192,N_26721,N_26770);
nand U27193 (N_27193,N_26976,N_26954);
nand U27194 (N_27194,N_26844,N_26767);
nand U27195 (N_27195,N_26747,N_26896);
and U27196 (N_27196,N_26767,N_26951);
xnor U27197 (N_27197,N_26976,N_26966);
xnor U27198 (N_27198,N_26761,N_26751);
or U27199 (N_27199,N_26963,N_26955);
and U27200 (N_27200,N_26764,N_26837);
xnor U27201 (N_27201,N_26794,N_26890);
or U27202 (N_27202,N_26949,N_26775);
and U27203 (N_27203,N_26954,N_26962);
and U27204 (N_27204,N_26887,N_26859);
and U27205 (N_27205,N_26887,N_26890);
and U27206 (N_27206,N_26712,N_26794);
or U27207 (N_27207,N_26931,N_26868);
or U27208 (N_27208,N_26842,N_26706);
nor U27209 (N_27209,N_26768,N_26809);
xor U27210 (N_27210,N_26741,N_26982);
xnor U27211 (N_27211,N_26725,N_26911);
or U27212 (N_27212,N_26906,N_26913);
or U27213 (N_27213,N_26915,N_26826);
nand U27214 (N_27214,N_26992,N_26764);
nor U27215 (N_27215,N_26925,N_26985);
and U27216 (N_27216,N_26720,N_26943);
nor U27217 (N_27217,N_26760,N_26832);
nand U27218 (N_27218,N_26708,N_26870);
nand U27219 (N_27219,N_26905,N_26926);
nand U27220 (N_27220,N_26759,N_26810);
xnor U27221 (N_27221,N_26867,N_26908);
and U27222 (N_27222,N_26877,N_26990);
xor U27223 (N_27223,N_26944,N_26930);
nand U27224 (N_27224,N_26878,N_26925);
or U27225 (N_27225,N_26878,N_26762);
and U27226 (N_27226,N_26823,N_26746);
and U27227 (N_27227,N_26866,N_26715);
nor U27228 (N_27228,N_26842,N_26780);
xor U27229 (N_27229,N_26781,N_26925);
nand U27230 (N_27230,N_26804,N_26726);
and U27231 (N_27231,N_26905,N_26935);
nor U27232 (N_27232,N_26971,N_26995);
xnor U27233 (N_27233,N_26756,N_26715);
nor U27234 (N_27234,N_26854,N_26703);
nand U27235 (N_27235,N_26940,N_26761);
nor U27236 (N_27236,N_26823,N_26743);
xor U27237 (N_27237,N_26971,N_26822);
or U27238 (N_27238,N_26789,N_26900);
nand U27239 (N_27239,N_26784,N_26798);
xor U27240 (N_27240,N_26901,N_26912);
nor U27241 (N_27241,N_26829,N_26772);
or U27242 (N_27242,N_26775,N_26938);
xor U27243 (N_27243,N_26932,N_26793);
nand U27244 (N_27244,N_26738,N_26819);
nand U27245 (N_27245,N_26973,N_26930);
nand U27246 (N_27246,N_26883,N_26927);
xor U27247 (N_27247,N_26944,N_26860);
or U27248 (N_27248,N_26702,N_26857);
xor U27249 (N_27249,N_26796,N_26934);
xnor U27250 (N_27250,N_26957,N_26801);
and U27251 (N_27251,N_26899,N_26725);
nand U27252 (N_27252,N_26820,N_26864);
or U27253 (N_27253,N_26878,N_26769);
xor U27254 (N_27254,N_26800,N_26832);
xnor U27255 (N_27255,N_26732,N_26918);
or U27256 (N_27256,N_26728,N_26805);
xor U27257 (N_27257,N_26953,N_26793);
and U27258 (N_27258,N_26966,N_26982);
or U27259 (N_27259,N_26933,N_26928);
or U27260 (N_27260,N_26808,N_26745);
or U27261 (N_27261,N_26756,N_26741);
or U27262 (N_27262,N_26915,N_26846);
xor U27263 (N_27263,N_26711,N_26900);
xnor U27264 (N_27264,N_26708,N_26889);
or U27265 (N_27265,N_26795,N_26968);
xnor U27266 (N_27266,N_26700,N_26869);
or U27267 (N_27267,N_26733,N_26827);
nand U27268 (N_27268,N_26834,N_26997);
xnor U27269 (N_27269,N_26752,N_26827);
or U27270 (N_27270,N_26843,N_26723);
and U27271 (N_27271,N_26978,N_26950);
or U27272 (N_27272,N_26875,N_26880);
and U27273 (N_27273,N_26957,N_26999);
xnor U27274 (N_27274,N_26914,N_26753);
nand U27275 (N_27275,N_26856,N_26978);
and U27276 (N_27276,N_26918,N_26806);
nor U27277 (N_27277,N_26954,N_26700);
nor U27278 (N_27278,N_26791,N_26918);
nor U27279 (N_27279,N_26836,N_26712);
nand U27280 (N_27280,N_26701,N_26892);
nand U27281 (N_27281,N_26978,N_26921);
or U27282 (N_27282,N_26818,N_26916);
nor U27283 (N_27283,N_26790,N_26759);
nand U27284 (N_27284,N_26707,N_26918);
or U27285 (N_27285,N_26852,N_26805);
nand U27286 (N_27286,N_26732,N_26906);
and U27287 (N_27287,N_26874,N_26857);
nor U27288 (N_27288,N_26846,N_26974);
nand U27289 (N_27289,N_26839,N_26778);
or U27290 (N_27290,N_26893,N_26755);
nand U27291 (N_27291,N_26900,N_26879);
or U27292 (N_27292,N_26890,N_26987);
or U27293 (N_27293,N_26774,N_26883);
nand U27294 (N_27294,N_26853,N_26746);
or U27295 (N_27295,N_26900,N_26729);
and U27296 (N_27296,N_26789,N_26997);
nor U27297 (N_27297,N_26726,N_26960);
or U27298 (N_27298,N_26810,N_26792);
nor U27299 (N_27299,N_26794,N_26750);
nor U27300 (N_27300,N_27105,N_27070);
or U27301 (N_27301,N_27150,N_27011);
and U27302 (N_27302,N_27025,N_27230);
nand U27303 (N_27303,N_27186,N_27182);
nand U27304 (N_27304,N_27127,N_27149);
xnor U27305 (N_27305,N_27162,N_27106);
and U27306 (N_27306,N_27014,N_27212);
and U27307 (N_27307,N_27043,N_27234);
or U27308 (N_27308,N_27282,N_27253);
xnor U27309 (N_27309,N_27130,N_27271);
xor U27310 (N_27310,N_27238,N_27024);
nor U27311 (N_27311,N_27229,N_27091);
and U27312 (N_27312,N_27272,N_27206);
nor U27313 (N_27313,N_27018,N_27075);
or U27314 (N_27314,N_27170,N_27260);
or U27315 (N_27315,N_27056,N_27210);
xor U27316 (N_27316,N_27288,N_27202);
or U27317 (N_27317,N_27211,N_27097);
nor U27318 (N_27318,N_27213,N_27079);
nand U27319 (N_27319,N_27021,N_27101);
and U27320 (N_27320,N_27051,N_27197);
nor U27321 (N_27321,N_27245,N_27246);
xor U27322 (N_27322,N_27259,N_27113);
nor U27323 (N_27323,N_27178,N_27016);
xnor U27324 (N_27324,N_27239,N_27085);
and U27325 (N_27325,N_27010,N_27279);
xor U27326 (N_27326,N_27093,N_27083);
nor U27327 (N_27327,N_27073,N_27254);
nand U27328 (N_27328,N_27166,N_27214);
or U27329 (N_27329,N_27045,N_27157);
or U27330 (N_27330,N_27129,N_27023);
xor U27331 (N_27331,N_27179,N_27019);
nor U27332 (N_27332,N_27298,N_27035);
or U27333 (N_27333,N_27071,N_27080);
xnor U27334 (N_27334,N_27276,N_27156);
nand U27335 (N_27335,N_27054,N_27123);
xor U27336 (N_27336,N_27012,N_27203);
nand U27337 (N_27337,N_27102,N_27030);
nand U27338 (N_27338,N_27022,N_27104);
and U27339 (N_27339,N_27169,N_27181);
and U27340 (N_27340,N_27152,N_27278);
nand U27341 (N_27341,N_27299,N_27161);
xor U27342 (N_27342,N_27265,N_27027);
xnor U27343 (N_27343,N_27228,N_27160);
and U27344 (N_27344,N_27001,N_27143);
xor U27345 (N_27345,N_27195,N_27068);
nor U27346 (N_27346,N_27266,N_27267);
nand U27347 (N_27347,N_27041,N_27221);
nor U27348 (N_27348,N_27120,N_27140);
xor U27349 (N_27349,N_27275,N_27227);
or U27350 (N_27350,N_27076,N_27223);
nor U27351 (N_27351,N_27167,N_27007);
or U27352 (N_27352,N_27031,N_27100);
nand U27353 (N_27353,N_27139,N_27292);
xor U27354 (N_27354,N_27126,N_27154);
and U27355 (N_27355,N_27183,N_27044);
nor U27356 (N_27356,N_27137,N_27244);
and U27357 (N_27357,N_27219,N_27231);
xor U27358 (N_27358,N_27216,N_27146);
xnor U27359 (N_27359,N_27142,N_27222);
and U27360 (N_27360,N_27060,N_27058);
nand U27361 (N_27361,N_27192,N_27037);
and U27362 (N_27362,N_27009,N_27194);
or U27363 (N_27363,N_27052,N_27115);
xor U27364 (N_27364,N_27177,N_27132);
xnor U27365 (N_27365,N_27048,N_27147);
or U27366 (N_27366,N_27198,N_27251);
and U27367 (N_27367,N_27078,N_27201);
and U27368 (N_27368,N_27050,N_27096);
nor U27369 (N_27369,N_27081,N_27233);
or U27370 (N_27370,N_27286,N_27098);
nand U27371 (N_27371,N_27066,N_27263);
nor U27372 (N_27372,N_27082,N_27042);
xnor U27373 (N_27373,N_27003,N_27165);
xor U27374 (N_27374,N_27297,N_27261);
nor U27375 (N_27375,N_27256,N_27258);
nand U27376 (N_27376,N_27188,N_27280);
xnor U27377 (N_27377,N_27122,N_27205);
or U27378 (N_27378,N_27119,N_27108);
or U27379 (N_27379,N_27099,N_27236);
and U27380 (N_27380,N_27284,N_27002);
xor U27381 (N_27381,N_27281,N_27175);
nor U27382 (N_27382,N_27061,N_27190);
or U27383 (N_27383,N_27065,N_27145);
nand U27384 (N_27384,N_27289,N_27257);
xnor U27385 (N_27385,N_27074,N_27116);
xor U27386 (N_27386,N_27028,N_27118);
nand U27387 (N_27387,N_27128,N_27013);
xor U27388 (N_27388,N_27036,N_27069);
xnor U27389 (N_27389,N_27086,N_27249);
nand U27390 (N_27390,N_27020,N_27136);
and U27391 (N_27391,N_27039,N_27172);
nor U27392 (N_27392,N_27247,N_27064);
and U27393 (N_27393,N_27243,N_27088);
and U27394 (N_27394,N_27109,N_27015);
xor U27395 (N_27395,N_27153,N_27226);
and U27396 (N_27396,N_27273,N_27200);
and U27397 (N_27397,N_27295,N_27163);
and U27398 (N_27398,N_27262,N_27224);
nor U27399 (N_27399,N_27057,N_27189);
nor U27400 (N_27400,N_27193,N_27173);
nand U27401 (N_27401,N_27270,N_27204);
nand U27402 (N_27402,N_27274,N_27092);
or U27403 (N_27403,N_27049,N_27047);
nor U27404 (N_27404,N_27138,N_27103);
and U27405 (N_27405,N_27090,N_27107);
nand U27406 (N_27406,N_27215,N_27121);
or U27407 (N_27407,N_27232,N_27144);
nand U27408 (N_27408,N_27133,N_27187);
or U27409 (N_27409,N_27084,N_27148);
nand U27410 (N_27410,N_27196,N_27117);
nor U27411 (N_27411,N_27242,N_27185);
nand U27412 (N_27412,N_27174,N_27277);
nor U27413 (N_27413,N_27134,N_27285);
nor U27414 (N_27414,N_27072,N_27255);
xnor U27415 (N_27415,N_27151,N_27269);
and U27416 (N_27416,N_27217,N_27055);
nor U27417 (N_27417,N_27112,N_27191);
and U27418 (N_27418,N_27199,N_27291);
or U27419 (N_27419,N_27124,N_27029);
nor U27420 (N_27420,N_27095,N_27158);
nor U27421 (N_27421,N_27059,N_27250);
nand U27422 (N_27422,N_27176,N_27155);
nor U27423 (N_27423,N_27026,N_27008);
and U27424 (N_27424,N_27077,N_27034);
xor U27425 (N_27425,N_27209,N_27125);
nor U27426 (N_27426,N_27287,N_27046);
xor U27427 (N_27427,N_27283,N_27111);
xor U27428 (N_27428,N_27290,N_27241);
nand U27429 (N_27429,N_27032,N_27268);
nor U27430 (N_27430,N_27218,N_27094);
nor U27431 (N_27431,N_27184,N_27252);
xor U27432 (N_27432,N_27164,N_27225);
xnor U27433 (N_27433,N_27000,N_27004);
and U27434 (N_27434,N_27264,N_27207);
and U27435 (N_27435,N_27237,N_27089);
and U27436 (N_27436,N_27294,N_27067);
or U27437 (N_27437,N_27296,N_27063);
xnor U27438 (N_27438,N_27017,N_27240);
xnor U27439 (N_27439,N_27062,N_27033);
xnor U27440 (N_27440,N_27005,N_27038);
xnor U27441 (N_27441,N_27110,N_27235);
nand U27442 (N_27442,N_27135,N_27293);
and U27443 (N_27443,N_27171,N_27053);
nor U27444 (N_27444,N_27006,N_27087);
or U27445 (N_27445,N_27159,N_27040);
nand U27446 (N_27446,N_27114,N_27168);
xor U27447 (N_27447,N_27208,N_27220);
nor U27448 (N_27448,N_27141,N_27131);
nor U27449 (N_27449,N_27248,N_27180);
or U27450 (N_27450,N_27110,N_27132);
xor U27451 (N_27451,N_27131,N_27183);
xor U27452 (N_27452,N_27186,N_27243);
and U27453 (N_27453,N_27121,N_27048);
nor U27454 (N_27454,N_27016,N_27168);
and U27455 (N_27455,N_27130,N_27075);
nand U27456 (N_27456,N_27171,N_27055);
xor U27457 (N_27457,N_27074,N_27167);
and U27458 (N_27458,N_27298,N_27026);
nand U27459 (N_27459,N_27094,N_27027);
nand U27460 (N_27460,N_27261,N_27247);
or U27461 (N_27461,N_27229,N_27152);
or U27462 (N_27462,N_27141,N_27202);
xor U27463 (N_27463,N_27253,N_27047);
xor U27464 (N_27464,N_27101,N_27025);
nand U27465 (N_27465,N_27260,N_27083);
xnor U27466 (N_27466,N_27138,N_27144);
and U27467 (N_27467,N_27146,N_27060);
xnor U27468 (N_27468,N_27264,N_27070);
or U27469 (N_27469,N_27189,N_27128);
nor U27470 (N_27470,N_27255,N_27132);
xnor U27471 (N_27471,N_27018,N_27039);
nand U27472 (N_27472,N_27187,N_27267);
xnor U27473 (N_27473,N_27207,N_27195);
or U27474 (N_27474,N_27249,N_27229);
nor U27475 (N_27475,N_27259,N_27091);
nor U27476 (N_27476,N_27290,N_27235);
xnor U27477 (N_27477,N_27286,N_27215);
and U27478 (N_27478,N_27069,N_27169);
xnor U27479 (N_27479,N_27127,N_27205);
nor U27480 (N_27480,N_27070,N_27249);
xor U27481 (N_27481,N_27295,N_27128);
nand U27482 (N_27482,N_27128,N_27187);
and U27483 (N_27483,N_27105,N_27228);
or U27484 (N_27484,N_27091,N_27003);
nand U27485 (N_27485,N_27179,N_27280);
or U27486 (N_27486,N_27293,N_27289);
nor U27487 (N_27487,N_27275,N_27283);
nor U27488 (N_27488,N_27071,N_27231);
nor U27489 (N_27489,N_27268,N_27250);
xnor U27490 (N_27490,N_27009,N_27049);
and U27491 (N_27491,N_27294,N_27100);
xnor U27492 (N_27492,N_27235,N_27154);
xor U27493 (N_27493,N_27117,N_27270);
and U27494 (N_27494,N_27253,N_27167);
xnor U27495 (N_27495,N_27214,N_27164);
or U27496 (N_27496,N_27224,N_27231);
or U27497 (N_27497,N_27037,N_27205);
or U27498 (N_27498,N_27016,N_27085);
and U27499 (N_27499,N_27164,N_27215);
xnor U27500 (N_27500,N_27149,N_27254);
or U27501 (N_27501,N_27056,N_27108);
or U27502 (N_27502,N_27019,N_27285);
and U27503 (N_27503,N_27036,N_27042);
xnor U27504 (N_27504,N_27127,N_27217);
nand U27505 (N_27505,N_27298,N_27159);
and U27506 (N_27506,N_27064,N_27218);
and U27507 (N_27507,N_27029,N_27044);
xor U27508 (N_27508,N_27160,N_27127);
nor U27509 (N_27509,N_27299,N_27009);
xor U27510 (N_27510,N_27153,N_27054);
nor U27511 (N_27511,N_27019,N_27139);
and U27512 (N_27512,N_27295,N_27249);
and U27513 (N_27513,N_27008,N_27021);
nand U27514 (N_27514,N_27099,N_27084);
xor U27515 (N_27515,N_27296,N_27222);
nand U27516 (N_27516,N_27001,N_27121);
nand U27517 (N_27517,N_27022,N_27042);
or U27518 (N_27518,N_27266,N_27023);
and U27519 (N_27519,N_27083,N_27075);
nand U27520 (N_27520,N_27225,N_27189);
and U27521 (N_27521,N_27298,N_27063);
and U27522 (N_27522,N_27048,N_27096);
xnor U27523 (N_27523,N_27099,N_27194);
xor U27524 (N_27524,N_27247,N_27051);
or U27525 (N_27525,N_27123,N_27037);
or U27526 (N_27526,N_27289,N_27010);
nand U27527 (N_27527,N_27041,N_27147);
nand U27528 (N_27528,N_27135,N_27296);
nand U27529 (N_27529,N_27094,N_27283);
xnor U27530 (N_27530,N_27030,N_27252);
nor U27531 (N_27531,N_27010,N_27152);
nor U27532 (N_27532,N_27282,N_27021);
nand U27533 (N_27533,N_27037,N_27035);
xnor U27534 (N_27534,N_27030,N_27121);
and U27535 (N_27535,N_27238,N_27165);
or U27536 (N_27536,N_27046,N_27179);
or U27537 (N_27537,N_27028,N_27068);
nor U27538 (N_27538,N_27294,N_27139);
xnor U27539 (N_27539,N_27132,N_27218);
and U27540 (N_27540,N_27001,N_27259);
and U27541 (N_27541,N_27184,N_27298);
nand U27542 (N_27542,N_27004,N_27275);
and U27543 (N_27543,N_27176,N_27006);
or U27544 (N_27544,N_27114,N_27248);
or U27545 (N_27545,N_27184,N_27234);
nand U27546 (N_27546,N_27026,N_27295);
xor U27547 (N_27547,N_27064,N_27216);
or U27548 (N_27548,N_27278,N_27293);
or U27549 (N_27549,N_27187,N_27011);
or U27550 (N_27550,N_27239,N_27121);
xnor U27551 (N_27551,N_27189,N_27181);
or U27552 (N_27552,N_27278,N_27227);
xor U27553 (N_27553,N_27027,N_27287);
nand U27554 (N_27554,N_27090,N_27095);
and U27555 (N_27555,N_27231,N_27234);
nor U27556 (N_27556,N_27015,N_27005);
xor U27557 (N_27557,N_27024,N_27079);
and U27558 (N_27558,N_27155,N_27285);
nor U27559 (N_27559,N_27088,N_27014);
nand U27560 (N_27560,N_27141,N_27171);
and U27561 (N_27561,N_27101,N_27261);
xnor U27562 (N_27562,N_27240,N_27110);
nand U27563 (N_27563,N_27094,N_27162);
and U27564 (N_27564,N_27025,N_27294);
nand U27565 (N_27565,N_27151,N_27133);
and U27566 (N_27566,N_27278,N_27284);
or U27567 (N_27567,N_27246,N_27030);
or U27568 (N_27568,N_27239,N_27050);
and U27569 (N_27569,N_27162,N_27238);
nor U27570 (N_27570,N_27252,N_27007);
nand U27571 (N_27571,N_27206,N_27190);
and U27572 (N_27572,N_27222,N_27081);
or U27573 (N_27573,N_27248,N_27030);
nand U27574 (N_27574,N_27168,N_27087);
nand U27575 (N_27575,N_27109,N_27208);
nand U27576 (N_27576,N_27179,N_27221);
nor U27577 (N_27577,N_27157,N_27116);
xor U27578 (N_27578,N_27269,N_27073);
or U27579 (N_27579,N_27269,N_27027);
nand U27580 (N_27580,N_27096,N_27127);
nor U27581 (N_27581,N_27048,N_27059);
or U27582 (N_27582,N_27211,N_27057);
and U27583 (N_27583,N_27045,N_27284);
and U27584 (N_27584,N_27106,N_27272);
xor U27585 (N_27585,N_27008,N_27123);
and U27586 (N_27586,N_27007,N_27030);
or U27587 (N_27587,N_27162,N_27239);
nand U27588 (N_27588,N_27048,N_27067);
xor U27589 (N_27589,N_27113,N_27278);
nand U27590 (N_27590,N_27159,N_27039);
nor U27591 (N_27591,N_27138,N_27218);
xor U27592 (N_27592,N_27076,N_27219);
and U27593 (N_27593,N_27051,N_27032);
and U27594 (N_27594,N_27139,N_27224);
and U27595 (N_27595,N_27229,N_27042);
xnor U27596 (N_27596,N_27299,N_27138);
nand U27597 (N_27597,N_27216,N_27033);
or U27598 (N_27598,N_27199,N_27259);
or U27599 (N_27599,N_27197,N_27137);
nor U27600 (N_27600,N_27383,N_27432);
xnor U27601 (N_27601,N_27389,N_27507);
or U27602 (N_27602,N_27365,N_27549);
xor U27603 (N_27603,N_27445,N_27550);
xnor U27604 (N_27604,N_27505,N_27311);
xor U27605 (N_27605,N_27338,N_27599);
nand U27606 (N_27606,N_27544,N_27527);
and U27607 (N_27607,N_27453,N_27334);
nor U27608 (N_27608,N_27428,N_27345);
nand U27609 (N_27609,N_27503,N_27373);
or U27610 (N_27610,N_27452,N_27476);
or U27611 (N_27611,N_27393,N_27502);
nor U27612 (N_27612,N_27440,N_27374);
or U27613 (N_27613,N_27372,N_27470);
nor U27614 (N_27614,N_27382,N_27411);
and U27615 (N_27615,N_27400,N_27519);
nor U27616 (N_27616,N_27341,N_27402);
nand U27617 (N_27617,N_27555,N_27556);
nor U27618 (N_27618,N_27590,N_27582);
and U27619 (N_27619,N_27533,N_27513);
and U27620 (N_27620,N_27315,N_27491);
or U27621 (N_27621,N_27394,N_27494);
nor U27622 (N_27622,N_27342,N_27312);
and U27623 (N_27623,N_27433,N_27427);
nor U27624 (N_27624,N_27495,N_27397);
and U27625 (N_27625,N_27306,N_27344);
or U27626 (N_27626,N_27425,N_27307);
or U27627 (N_27627,N_27329,N_27579);
and U27628 (N_27628,N_27384,N_27401);
nor U27629 (N_27629,N_27523,N_27477);
or U27630 (N_27630,N_27508,N_27352);
xnor U27631 (N_27631,N_27408,N_27593);
nand U27632 (N_27632,N_27577,N_27521);
nor U27633 (N_27633,N_27490,N_27305);
nor U27634 (N_27634,N_27461,N_27378);
nand U27635 (N_27635,N_27357,N_27359);
xor U27636 (N_27636,N_27355,N_27498);
nor U27637 (N_27637,N_27339,N_27324);
nand U27638 (N_27638,N_27443,N_27501);
nand U27639 (N_27639,N_27518,N_27569);
or U27640 (N_27640,N_27471,N_27396);
xor U27641 (N_27641,N_27540,N_27512);
nand U27642 (N_27642,N_27539,N_27541);
xnor U27643 (N_27643,N_27438,N_27412);
nor U27644 (N_27644,N_27409,N_27585);
or U27645 (N_27645,N_27573,N_27464);
nor U27646 (N_27646,N_27414,N_27459);
xnor U27647 (N_27647,N_27525,N_27514);
and U27648 (N_27648,N_27504,N_27407);
and U27649 (N_27649,N_27361,N_27472);
or U27650 (N_27650,N_27468,N_27576);
or U27651 (N_27651,N_27388,N_27422);
nand U27652 (N_27652,N_27553,N_27526);
nand U27653 (N_27653,N_27321,N_27368);
xnor U27654 (N_27654,N_27456,N_27535);
nor U27655 (N_27655,N_27435,N_27462);
and U27656 (N_27656,N_27337,N_27565);
nand U27657 (N_27657,N_27360,N_27350);
nand U27658 (N_27658,N_27302,N_27377);
nand U27659 (N_27659,N_27530,N_27482);
nand U27660 (N_27660,N_27580,N_27466);
and U27661 (N_27661,N_27387,N_27566);
xnor U27662 (N_27662,N_27586,N_27376);
and U27663 (N_27663,N_27367,N_27583);
and U27664 (N_27664,N_27568,N_27588);
and U27665 (N_27665,N_27316,N_27543);
and U27666 (N_27666,N_27354,N_27366);
nor U27667 (N_27667,N_27455,N_27493);
nand U27668 (N_27668,N_27506,N_27325);
nor U27669 (N_27669,N_27436,N_27563);
nor U27670 (N_27670,N_27591,N_27317);
xnor U27671 (N_27671,N_27310,N_27301);
xor U27672 (N_27672,N_27348,N_27390);
nor U27673 (N_27673,N_27496,N_27489);
and U27674 (N_27674,N_27536,N_27385);
xor U27675 (N_27675,N_27441,N_27564);
nand U27676 (N_27676,N_27415,N_27460);
and U27677 (N_27677,N_27347,N_27308);
nor U27678 (N_27678,N_27562,N_27446);
or U27679 (N_27679,N_27375,N_27304);
nand U27680 (N_27680,N_27353,N_27399);
nand U27681 (N_27681,N_27458,N_27370);
or U27682 (N_27682,N_27546,N_27487);
or U27683 (N_27683,N_27548,N_27333);
xor U27684 (N_27684,N_27596,N_27369);
and U27685 (N_27685,N_27392,N_27488);
and U27686 (N_27686,N_27531,N_27574);
nor U27687 (N_27687,N_27300,N_27499);
or U27688 (N_27688,N_27371,N_27450);
and U27689 (N_27689,N_27320,N_27363);
and U27690 (N_27690,N_27449,N_27303);
nand U27691 (N_27691,N_27380,N_27434);
or U27692 (N_27692,N_27484,N_27578);
or U27693 (N_27693,N_27457,N_27575);
xnor U27694 (N_27694,N_27481,N_27560);
or U27695 (N_27695,N_27485,N_27480);
xor U27696 (N_27696,N_27528,N_27358);
nand U27697 (N_27697,N_27410,N_27403);
nand U27698 (N_27698,N_27424,N_27511);
and U27699 (N_27699,N_27405,N_27572);
or U27700 (N_27700,N_27486,N_27559);
nor U27701 (N_27701,N_27581,N_27444);
nor U27702 (N_27702,N_27534,N_27537);
and U27703 (N_27703,N_27395,N_27439);
or U27704 (N_27704,N_27542,N_27515);
nand U27705 (N_27705,N_27419,N_27545);
xnor U27706 (N_27706,N_27421,N_27413);
nor U27707 (N_27707,N_27351,N_27430);
xnor U27708 (N_27708,N_27592,N_27336);
and U27709 (N_27709,N_27483,N_27510);
or U27710 (N_27710,N_27589,N_27597);
nand U27711 (N_27711,N_27538,N_27416);
nand U27712 (N_27712,N_27420,N_27492);
nand U27713 (N_27713,N_27448,N_27327);
nor U27714 (N_27714,N_27532,N_27442);
nor U27715 (N_27715,N_27429,N_27326);
and U27716 (N_27716,N_27404,N_27356);
or U27717 (N_27717,N_27349,N_27386);
and U27718 (N_27718,N_27547,N_27346);
or U27719 (N_27719,N_27509,N_27335);
and U27720 (N_27720,N_27474,N_27340);
or U27721 (N_27721,N_27465,N_27451);
xor U27722 (N_27722,N_27322,N_27331);
or U27723 (N_27723,N_27406,N_27595);
or U27724 (N_27724,N_27379,N_27516);
nor U27725 (N_27725,N_27417,N_27469);
or U27726 (N_27726,N_27423,N_27497);
nand U27727 (N_27727,N_27454,N_27551);
nand U27728 (N_27728,N_27362,N_27558);
or U27729 (N_27729,N_27522,N_27391);
nand U27730 (N_27730,N_27479,N_27557);
or U27731 (N_27731,N_27309,N_27529);
and U27732 (N_27732,N_27561,N_27447);
nand U27733 (N_27733,N_27475,N_27313);
and U27734 (N_27734,N_27520,N_27500);
or U27735 (N_27735,N_27598,N_27594);
and U27736 (N_27736,N_27463,N_27426);
or U27737 (N_27737,N_27467,N_27554);
and U27738 (N_27738,N_27524,N_27571);
nor U27739 (N_27739,N_27473,N_27364);
nor U27740 (N_27740,N_27437,N_27418);
nand U27741 (N_27741,N_27431,N_27478);
nor U27742 (N_27742,N_27319,N_27343);
and U27743 (N_27743,N_27567,N_27584);
and U27744 (N_27744,N_27517,N_27318);
or U27745 (N_27745,N_27381,N_27323);
nor U27746 (N_27746,N_27314,N_27398);
or U27747 (N_27747,N_27570,N_27328);
and U27748 (N_27748,N_27587,N_27330);
and U27749 (N_27749,N_27552,N_27332);
nand U27750 (N_27750,N_27427,N_27414);
nand U27751 (N_27751,N_27538,N_27348);
xor U27752 (N_27752,N_27478,N_27397);
nand U27753 (N_27753,N_27465,N_27553);
or U27754 (N_27754,N_27530,N_27428);
or U27755 (N_27755,N_27399,N_27429);
and U27756 (N_27756,N_27583,N_27571);
xor U27757 (N_27757,N_27310,N_27384);
and U27758 (N_27758,N_27560,N_27454);
xnor U27759 (N_27759,N_27421,N_27389);
or U27760 (N_27760,N_27400,N_27345);
nor U27761 (N_27761,N_27344,N_27594);
nor U27762 (N_27762,N_27404,N_27451);
xnor U27763 (N_27763,N_27338,N_27527);
xnor U27764 (N_27764,N_27396,N_27338);
and U27765 (N_27765,N_27430,N_27330);
xor U27766 (N_27766,N_27409,N_27389);
xor U27767 (N_27767,N_27572,N_27436);
nor U27768 (N_27768,N_27562,N_27328);
nor U27769 (N_27769,N_27379,N_27325);
or U27770 (N_27770,N_27494,N_27366);
nand U27771 (N_27771,N_27458,N_27392);
nand U27772 (N_27772,N_27544,N_27362);
xnor U27773 (N_27773,N_27339,N_27581);
xnor U27774 (N_27774,N_27504,N_27338);
nor U27775 (N_27775,N_27352,N_27301);
and U27776 (N_27776,N_27443,N_27397);
nor U27777 (N_27777,N_27301,N_27319);
xor U27778 (N_27778,N_27586,N_27383);
xnor U27779 (N_27779,N_27491,N_27489);
and U27780 (N_27780,N_27374,N_27318);
nor U27781 (N_27781,N_27334,N_27357);
nand U27782 (N_27782,N_27367,N_27313);
xor U27783 (N_27783,N_27574,N_27511);
xnor U27784 (N_27784,N_27445,N_27379);
or U27785 (N_27785,N_27363,N_27392);
xor U27786 (N_27786,N_27457,N_27321);
xnor U27787 (N_27787,N_27393,N_27302);
xnor U27788 (N_27788,N_27546,N_27386);
nand U27789 (N_27789,N_27385,N_27436);
xor U27790 (N_27790,N_27581,N_27500);
xor U27791 (N_27791,N_27356,N_27302);
or U27792 (N_27792,N_27533,N_27548);
and U27793 (N_27793,N_27554,N_27484);
and U27794 (N_27794,N_27440,N_27309);
xnor U27795 (N_27795,N_27359,N_27301);
xor U27796 (N_27796,N_27576,N_27422);
or U27797 (N_27797,N_27515,N_27514);
nor U27798 (N_27798,N_27451,N_27436);
xor U27799 (N_27799,N_27389,N_27530);
and U27800 (N_27800,N_27427,N_27570);
nand U27801 (N_27801,N_27466,N_27317);
xnor U27802 (N_27802,N_27593,N_27392);
nor U27803 (N_27803,N_27317,N_27376);
and U27804 (N_27804,N_27347,N_27481);
xnor U27805 (N_27805,N_27344,N_27579);
xor U27806 (N_27806,N_27465,N_27370);
xor U27807 (N_27807,N_27579,N_27399);
or U27808 (N_27808,N_27576,N_27538);
nand U27809 (N_27809,N_27486,N_27431);
nor U27810 (N_27810,N_27342,N_27356);
nand U27811 (N_27811,N_27453,N_27583);
or U27812 (N_27812,N_27480,N_27508);
or U27813 (N_27813,N_27549,N_27300);
nor U27814 (N_27814,N_27334,N_27308);
xnor U27815 (N_27815,N_27369,N_27456);
nand U27816 (N_27816,N_27515,N_27531);
nand U27817 (N_27817,N_27572,N_27374);
or U27818 (N_27818,N_27447,N_27563);
nand U27819 (N_27819,N_27517,N_27366);
xnor U27820 (N_27820,N_27392,N_27505);
or U27821 (N_27821,N_27346,N_27553);
nor U27822 (N_27822,N_27512,N_27376);
nand U27823 (N_27823,N_27568,N_27496);
or U27824 (N_27824,N_27428,N_27499);
and U27825 (N_27825,N_27324,N_27405);
nand U27826 (N_27826,N_27401,N_27571);
nor U27827 (N_27827,N_27559,N_27456);
nor U27828 (N_27828,N_27547,N_27520);
xnor U27829 (N_27829,N_27444,N_27578);
nor U27830 (N_27830,N_27489,N_27384);
nor U27831 (N_27831,N_27424,N_27390);
or U27832 (N_27832,N_27404,N_27322);
and U27833 (N_27833,N_27421,N_27310);
nand U27834 (N_27834,N_27515,N_27404);
or U27835 (N_27835,N_27597,N_27452);
or U27836 (N_27836,N_27570,N_27423);
or U27837 (N_27837,N_27350,N_27393);
nor U27838 (N_27838,N_27574,N_27534);
nand U27839 (N_27839,N_27591,N_27375);
and U27840 (N_27840,N_27534,N_27598);
nand U27841 (N_27841,N_27576,N_27424);
nand U27842 (N_27842,N_27425,N_27395);
nand U27843 (N_27843,N_27379,N_27506);
nor U27844 (N_27844,N_27566,N_27589);
and U27845 (N_27845,N_27378,N_27396);
nor U27846 (N_27846,N_27519,N_27482);
and U27847 (N_27847,N_27340,N_27511);
or U27848 (N_27848,N_27360,N_27488);
nor U27849 (N_27849,N_27349,N_27447);
nor U27850 (N_27850,N_27408,N_27333);
nand U27851 (N_27851,N_27550,N_27508);
and U27852 (N_27852,N_27547,N_27474);
and U27853 (N_27853,N_27445,N_27363);
or U27854 (N_27854,N_27441,N_27567);
nor U27855 (N_27855,N_27427,N_27311);
nand U27856 (N_27856,N_27537,N_27309);
xnor U27857 (N_27857,N_27463,N_27433);
or U27858 (N_27858,N_27476,N_27360);
xor U27859 (N_27859,N_27508,N_27425);
nor U27860 (N_27860,N_27365,N_27437);
or U27861 (N_27861,N_27433,N_27484);
nand U27862 (N_27862,N_27382,N_27448);
or U27863 (N_27863,N_27557,N_27394);
xnor U27864 (N_27864,N_27430,N_27325);
or U27865 (N_27865,N_27406,N_27318);
nor U27866 (N_27866,N_27364,N_27476);
nand U27867 (N_27867,N_27563,N_27585);
nand U27868 (N_27868,N_27501,N_27367);
xor U27869 (N_27869,N_27553,N_27348);
nor U27870 (N_27870,N_27550,N_27490);
nor U27871 (N_27871,N_27381,N_27452);
or U27872 (N_27872,N_27340,N_27432);
nor U27873 (N_27873,N_27401,N_27432);
xor U27874 (N_27874,N_27377,N_27489);
xnor U27875 (N_27875,N_27370,N_27481);
nor U27876 (N_27876,N_27470,N_27491);
xnor U27877 (N_27877,N_27537,N_27462);
nor U27878 (N_27878,N_27451,N_27491);
xor U27879 (N_27879,N_27341,N_27486);
nor U27880 (N_27880,N_27479,N_27528);
or U27881 (N_27881,N_27529,N_27406);
or U27882 (N_27882,N_27503,N_27345);
or U27883 (N_27883,N_27444,N_27336);
nand U27884 (N_27884,N_27378,N_27531);
and U27885 (N_27885,N_27574,N_27424);
xor U27886 (N_27886,N_27483,N_27470);
or U27887 (N_27887,N_27549,N_27458);
and U27888 (N_27888,N_27362,N_27311);
xnor U27889 (N_27889,N_27396,N_27525);
and U27890 (N_27890,N_27440,N_27453);
and U27891 (N_27891,N_27432,N_27543);
or U27892 (N_27892,N_27584,N_27301);
nand U27893 (N_27893,N_27376,N_27528);
nor U27894 (N_27894,N_27516,N_27425);
nand U27895 (N_27895,N_27558,N_27361);
or U27896 (N_27896,N_27573,N_27578);
and U27897 (N_27897,N_27311,N_27501);
xnor U27898 (N_27898,N_27547,N_27453);
and U27899 (N_27899,N_27576,N_27353);
nor U27900 (N_27900,N_27895,N_27796);
and U27901 (N_27901,N_27851,N_27630);
xor U27902 (N_27902,N_27650,N_27855);
xnor U27903 (N_27903,N_27633,N_27703);
xnor U27904 (N_27904,N_27636,N_27810);
and U27905 (N_27905,N_27876,N_27659);
nand U27906 (N_27906,N_27782,N_27727);
or U27907 (N_27907,N_27849,N_27888);
or U27908 (N_27908,N_27692,N_27770);
and U27909 (N_27909,N_27623,N_27698);
nor U27910 (N_27910,N_27629,N_27886);
nand U27911 (N_27911,N_27771,N_27774);
or U27912 (N_27912,N_27695,N_27662);
xnor U27913 (N_27913,N_27673,N_27644);
xor U27914 (N_27914,N_27688,N_27850);
nand U27915 (N_27915,N_27613,N_27658);
and U27916 (N_27916,N_27822,N_27816);
and U27917 (N_27917,N_27869,N_27844);
xor U27918 (N_27918,N_27818,N_27645);
xnor U27919 (N_27919,N_27655,N_27733);
nor U27920 (N_27920,N_27708,N_27714);
and U27921 (N_27921,N_27620,N_27606);
or U27922 (N_27922,N_27651,N_27792);
or U27923 (N_27923,N_27835,N_27853);
and U27924 (N_27924,N_27700,N_27820);
nand U27925 (N_27925,N_27762,N_27618);
xor U27926 (N_27926,N_27674,N_27772);
nor U27927 (N_27927,N_27656,N_27899);
nor U27928 (N_27928,N_27731,N_27697);
nand U27929 (N_27929,N_27631,N_27872);
xnor U27930 (N_27930,N_27778,N_27661);
and U27931 (N_27931,N_27707,N_27824);
and U27932 (N_27932,N_27775,N_27848);
xor U27933 (N_27933,N_27639,N_27632);
xor U27934 (N_27934,N_27693,N_27611);
xnor U27935 (N_27935,N_27859,N_27821);
xnor U27936 (N_27936,N_27619,N_27600);
nand U27937 (N_27937,N_27798,N_27761);
nor U27938 (N_27938,N_27654,N_27719);
xnor U27939 (N_27939,N_27829,N_27734);
or U27940 (N_27940,N_27720,N_27741);
or U27941 (N_27941,N_27825,N_27742);
or U27942 (N_27942,N_27841,N_27812);
xor U27943 (N_27943,N_27676,N_27670);
or U27944 (N_27944,N_27747,N_27802);
nand U27945 (N_27945,N_27870,N_27861);
nor U27946 (N_27946,N_27814,N_27668);
nand U27947 (N_27947,N_27682,N_27722);
or U27948 (N_27948,N_27652,N_27750);
nor U27949 (N_27949,N_27758,N_27875);
nand U27950 (N_27950,N_27787,N_27809);
nand U27951 (N_27951,N_27874,N_27681);
or U27952 (N_27952,N_27696,N_27637);
xor U27953 (N_27953,N_27799,N_27838);
nand U27954 (N_27954,N_27625,N_27601);
xnor U27955 (N_27955,N_27718,N_27826);
xor U27956 (N_27956,N_27836,N_27667);
and U27957 (N_27957,N_27789,N_27635);
nor U27958 (N_27958,N_27788,N_27884);
xor U27959 (N_27959,N_27880,N_27605);
nor U27960 (N_27960,N_27807,N_27857);
nand U27961 (N_27961,N_27828,N_27689);
or U27962 (N_27962,N_27737,N_27781);
nor U27963 (N_27963,N_27867,N_27891);
nand U27964 (N_27964,N_27843,N_27804);
and U27965 (N_27965,N_27756,N_27704);
and U27966 (N_27966,N_27705,N_27648);
xnor U27967 (N_27967,N_27759,N_27607);
and U27968 (N_27968,N_27800,N_27755);
nand U27969 (N_27969,N_27839,N_27752);
or U27970 (N_27970,N_27729,N_27678);
and U27971 (N_27971,N_27649,N_27643);
or U27972 (N_27972,N_27642,N_27602);
xor U27973 (N_27973,N_27675,N_27691);
xnor U27974 (N_27974,N_27721,N_27793);
and U27975 (N_27975,N_27783,N_27746);
nor U27976 (N_27976,N_27677,N_27864);
nand U27977 (N_27977,N_27712,N_27898);
nand U27978 (N_27978,N_27615,N_27616);
or U27979 (N_27979,N_27687,N_27711);
nor U27980 (N_27980,N_27865,N_27690);
nor U27981 (N_27981,N_27858,N_27634);
and U27982 (N_27982,N_27724,N_27827);
or U27983 (N_27983,N_27685,N_27640);
or U27984 (N_27984,N_27622,N_27866);
or U27985 (N_27985,N_27854,N_27878);
or U27986 (N_27986,N_27608,N_27686);
nor U27987 (N_27987,N_27766,N_27845);
and U27988 (N_27988,N_27887,N_27725);
or U27989 (N_27989,N_27694,N_27754);
nand U27990 (N_27990,N_27817,N_27837);
nor U27991 (N_27991,N_27834,N_27871);
and U27992 (N_27992,N_27896,N_27765);
and U27993 (N_27993,N_27868,N_27751);
and U27994 (N_27994,N_27873,N_27740);
or U27995 (N_27995,N_27815,N_27610);
or U27996 (N_27996,N_27609,N_27672);
xnor U27997 (N_27997,N_27624,N_27791);
or U27998 (N_27998,N_27883,N_27769);
xor U27999 (N_27999,N_27726,N_27663);
nand U28000 (N_28000,N_27735,N_27847);
or U28001 (N_28001,N_27790,N_27660);
or U28002 (N_28002,N_27717,N_27612);
xnor U28003 (N_28003,N_27617,N_27863);
nor U28004 (N_28004,N_27819,N_27823);
xor U28005 (N_28005,N_27780,N_27743);
nand U28006 (N_28006,N_27646,N_27763);
nand U28007 (N_28007,N_27889,N_27664);
or U28008 (N_28008,N_27683,N_27894);
xnor U28009 (N_28009,N_27715,N_27699);
and U28010 (N_28010,N_27882,N_27808);
and U28011 (N_28011,N_27877,N_27665);
nand U28012 (N_28012,N_27760,N_27753);
and U28013 (N_28013,N_27785,N_27797);
xnor U28014 (N_28014,N_27831,N_27628);
and U28015 (N_28015,N_27846,N_27768);
xnor U28016 (N_28016,N_27627,N_27786);
nor U28017 (N_28017,N_27736,N_27806);
or U28018 (N_28018,N_27749,N_27803);
xnor U28019 (N_28019,N_27892,N_27885);
nor U28020 (N_28020,N_27833,N_27745);
nor U28021 (N_28021,N_27723,N_27701);
and U28022 (N_28022,N_27710,N_27702);
and U28023 (N_28023,N_27767,N_27684);
nor U28024 (N_28024,N_27897,N_27679);
nor U28025 (N_28025,N_27795,N_27852);
nor U28026 (N_28026,N_27890,N_27779);
nor U28027 (N_28027,N_27893,N_27638);
nor U28028 (N_28028,N_27614,N_27738);
nand U28029 (N_28029,N_27709,N_27811);
or U28030 (N_28030,N_27669,N_27757);
nand U28031 (N_28031,N_27621,N_27748);
or U28032 (N_28032,N_27805,N_27641);
nor U28033 (N_28033,N_27776,N_27730);
and U28034 (N_28034,N_27647,N_27716);
nor U28035 (N_28035,N_27666,N_27626);
nand U28036 (N_28036,N_27840,N_27773);
nor U28037 (N_28037,N_27744,N_27728);
xnor U28038 (N_28038,N_27813,N_27653);
and U28039 (N_28039,N_27732,N_27739);
xor U28040 (N_28040,N_27713,N_27881);
nor U28041 (N_28041,N_27706,N_27603);
nor U28042 (N_28042,N_27794,N_27860);
nand U28043 (N_28043,N_27830,N_27604);
nor U28044 (N_28044,N_27657,N_27671);
nand U28045 (N_28045,N_27856,N_27842);
nor U28046 (N_28046,N_27777,N_27832);
nand U28047 (N_28047,N_27764,N_27801);
and U28048 (N_28048,N_27862,N_27879);
and U28049 (N_28049,N_27680,N_27784);
nand U28050 (N_28050,N_27804,N_27603);
nor U28051 (N_28051,N_27845,N_27690);
nor U28052 (N_28052,N_27805,N_27834);
nor U28053 (N_28053,N_27741,N_27736);
nand U28054 (N_28054,N_27651,N_27662);
nand U28055 (N_28055,N_27750,N_27618);
xor U28056 (N_28056,N_27839,N_27716);
and U28057 (N_28057,N_27716,N_27700);
nor U28058 (N_28058,N_27838,N_27607);
xor U28059 (N_28059,N_27736,N_27648);
or U28060 (N_28060,N_27867,N_27670);
or U28061 (N_28061,N_27683,N_27849);
nor U28062 (N_28062,N_27859,N_27759);
or U28063 (N_28063,N_27830,N_27689);
or U28064 (N_28064,N_27610,N_27724);
nand U28065 (N_28065,N_27710,N_27751);
or U28066 (N_28066,N_27794,N_27793);
nor U28067 (N_28067,N_27767,N_27807);
or U28068 (N_28068,N_27637,N_27691);
xor U28069 (N_28069,N_27677,N_27659);
xnor U28070 (N_28070,N_27654,N_27637);
or U28071 (N_28071,N_27603,N_27702);
nand U28072 (N_28072,N_27848,N_27686);
nand U28073 (N_28073,N_27691,N_27852);
or U28074 (N_28074,N_27858,N_27847);
xnor U28075 (N_28075,N_27844,N_27837);
and U28076 (N_28076,N_27778,N_27648);
and U28077 (N_28077,N_27792,N_27888);
xor U28078 (N_28078,N_27842,N_27898);
nor U28079 (N_28079,N_27791,N_27710);
xnor U28080 (N_28080,N_27691,N_27894);
or U28081 (N_28081,N_27734,N_27705);
xnor U28082 (N_28082,N_27840,N_27865);
nor U28083 (N_28083,N_27669,N_27627);
nor U28084 (N_28084,N_27659,N_27762);
nand U28085 (N_28085,N_27877,N_27745);
xnor U28086 (N_28086,N_27722,N_27794);
nand U28087 (N_28087,N_27737,N_27892);
nand U28088 (N_28088,N_27779,N_27695);
nor U28089 (N_28089,N_27785,N_27663);
and U28090 (N_28090,N_27820,N_27680);
nand U28091 (N_28091,N_27769,N_27819);
nor U28092 (N_28092,N_27816,N_27861);
nor U28093 (N_28093,N_27738,N_27617);
and U28094 (N_28094,N_27800,N_27657);
nor U28095 (N_28095,N_27878,N_27676);
xor U28096 (N_28096,N_27740,N_27671);
nor U28097 (N_28097,N_27864,N_27687);
nor U28098 (N_28098,N_27673,N_27633);
nor U28099 (N_28099,N_27817,N_27725);
nand U28100 (N_28100,N_27823,N_27757);
or U28101 (N_28101,N_27694,N_27798);
nand U28102 (N_28102,N_27684,N_27605);
or U28103 (N_28103,N_27745,N_27825);
nor U28104 (N_28104,N_27853,N_27852);
nor U28105 (N_28105,N_27631,N_27769);
xor U28106 (N_28106,N_27897,N_27622);
nand U28107 (N_28107,N_27687,N_27897);
xnor U28108 (N_28108,N_27734,N_27649);
or U28109 (N_28109,N_27697,N_27717);
nand U28110 (N_28110,N_27896,N_27629);
and U28111 (N_28111,N_27785,N_27772);
nand U28112 (N_28112,N_27688,N_27625);
xor U28113 (N_28113,N_27676,N_27808);
xor U28114 (N_28114,N_27750,N_27711);
or U28115 (N_28115,N_27851,N_27865);
or U28116 (N_28116,N_27628,N_27778);
xor U28117 (N_28117,N_27721,N_27744);
and U28118 (N_28118,N_27703,N_27714);
nand U28119 (N_28119,N_27619,N_27764);
nand U28120 (N_28120,N_27706,N_27760);
nor U28121 (N_28121,N_27635,N_27790);
xnor U28122 (N_28122,N_27861,N_27891);
xnor U28123 (N_28123,N_27836,N_27700);
nand U28124 (N_28124,N_27761,N_27659);
nor U28125 (N_28125,N_27783,N_27688);
xor U28126 (N_28126,N_27717,N_27770);
or U28127 (N_28127,N_27841,N_27891);
nand U28128 (N_28128,N_27780,N_27728);
or U28129 (N_28129,N_27686,N_27870);
nand U28130 (N_28130,N_27712,N_27851);
xnor U28131 (N_28131,N_27679,N_27678);
or U28132 (N_28132,N_27611,N_27847);
nand U28133 (N_28133,N_27669,N_27613);
xnor U28134 (N_28134,N_27600,N_27737);
and U28135 (N_28135,N_27638,N_27755);
and U28136 (N_28136,N_27724,N_27661);
and U28137 (N_28137,N_27716,N_27707);
nand U28138 (N_28138,N_27888,N_27691);
or U28139 (N_28139,N_27666,N_27879);
nand U28140 (N_28140,N_27627,N_27774);
xnor U28141 (N_28141,N_27757,N_27639);
nor U28142 (N_28142,N_27603,N_27670);
nand U28143 (N_28143,N_27807,N_27724);
nor U28144 (N_28144,N_27842,N_27603);
nand U28145 (N_28145,N_27772,N_27838);
and U28146 (N_28146,N_27805,N_27662);
nand U28147 (N_28147,N_27786,N_27842);
and U28148 (N_28148,N_27819,N_27687);
or U28149 (N_28149,N_27835,N_27830);
and U28150 (N_28150,N_27672,N_27636);
nor U28151 (N_28151,N_27800,N_27774);
xor U28152 (N_28152,N_27710,N_27804);
nor U28153 (N_28153,N_27785,N_27897);
nand U28154 (N_28154,N_27647,N_27835);
nor U28155 (N_28155,N_27777,N_27636);
nand U28156 (N_28156,N_27816,N_27670);
or U28157 (N_28157,N_27723,N_27671);
nand U28158 (N_28158,N_27677,N_27795);
and U28159 (N_28159,N_27836,N_27638);
and U28160 (N_28160,N_27601,N_27773);
nand U28161 (N_28161,N_27898,N_27853);
nand U28162 (N_28162,N_27621,N_27857);
or U28163 (N_28163,N_27703,N_27656);
nand U28164 (N_28164,N_27745,N_27771);
xnor U28165 (N_28165,N_27604,N_27857);
nand U28166 (N_28166,N_27825,N_27882);
and U28167 (N_28167,N_27810,N_27785);
nand U28168 (N_28168,N_27885,N_27817);
nand U28169 (N_28169,N_27731,N_27891);
or U28170 (N_28170,N_27752,N_27616);
nor U28171 (N_28171,N_27706,N_27842);
nor U28172 (N_28172,N_27658,N_27612);
and U28173 (N_28173,N_27739,N_27741);
nand U28174 (N_28174,N_27813,N_27717);
xor U28175 (N_28175,N_27644,N_27837);
nor U28176 (N_28176,N_27892,N_27860);
xnor U28177 (N_28177,N_27706,N_27871);
and U28178 (N_28178,N_27660,N_27601);
xnor U28179 (N_28179,N_27614,N_27608);
nand U28180 (N_28180,N_27699,N_27872);
or U28181 (N_28181,N_27807,N_27628);
or U28182 (N_28182,N_27634,N_27891);
or U28183 (N_28183,N_27639,N_27715);
and U28184 (N_28184,N_27897,N_27654);
nand U28185 (N_28185,N_27672,N_27753);
xnor U28186 (N_28186,N_27649,N_27711);
xnor U28187 (N_28187,N_27755,N_27756);
nand U28188 (N_28188,N_27648,N_27718);
nand U28189 (N_28189,N_27767,N_27812);
nor U28190 (N_28190,N_27643,N_27713);
xor U28191 (N_28191,N_27672,N_27737);
xor U28192 (N_28192,N_27777,N_27898);
xor U28193 (N_28193,N_27719,N_27640);
xor U28194 (N_28194,N_27642,N_27611);
xnor U28195 (N_28195,N_27793,N_27748);
and U28196 (N_28196,N_27801,N_27843);
nand U28197 (N_28197,N_27814,N_27635);
and U28198 (N_28198,N_27747,N_27679);
and U28199 (N_28199,N_27697,N_27695);
and U28200 (N_28200,N_28140,N_28072);
and U28201 (N_28201,N_28176,N_28148);
nand U28202 (N_28202,N_28016,N_28178);
xor U28203 (N_28203,N_28147,N_28137);
or U28204 (N_28204,N_28052,N_27989);
or U28205 (N_28205,N_28057,N_28193);
and U28206 (N_28206,N_27938,N_27908);
nand U28207 (N_28207,N_27920,N_27982);
xor U28208 (N_28208,N_27915,N_28011);
nand U28209 (N_28209,N_28063,N_28007);
xor U28210 (N_28210,N_28083,N_28146);
xnor U28211 (N_28211,N_27934,N_28032);
xor U28212 (N_28212,N_28149,N_28163);
xnor U28213 (N_28213,N_28095,N_28005);
nor U28214 (N_28214,N_28089,N_28161);
and U28215 (N_28215,N_27973,N_28003);
nand U28216 (N_28216,N_27930,N_28190);
or U28217 (N_28217,N_28069,N_28028);
nor U28218 (N_28218,N_28116,N_28145);
nand U28219 (N_28219,N_28080,N_28192);
nor U28220 (N_28220,N_27951,N_28039);
and U28221 (N_28221,N_28162,N_27994);
or U28222 (N_28222,N_28012,N_27958);
nor U28223 (N_28223,N_28025,N_28125);
xor U28224 (N_28224,N_27985,N_27931);
nor U28225 (N_28225,N_27975,N_28111);
nand U28226 (N_28226,N_28010,N_27987);
xnor U28227 (N_28227,N_28197,N_28092);
nor U28228 (N_28228,N_28041,N_28000);
nor U28229 (N_28229,N_28196,N_28076);
and U28230 (N_28230,N_28105,N_28183);
and U28231 (N_28231,N_27936,N_28094);
and U28232 (N_28232,N_27954,N_27913);
and U28233 (N_28233,N_27921,N_28188);
or U28234 (N_28234,N_27968,N_28187);
nor U28235 (N_28235,N_28048,N_28139);
and U28236 (N_28236,N_28158,N_28013);
and U28237 (N_28237,N_28086,N_28185);
and U28238 (N_28238,N_27988,N_28040);
or U28239 (N_28239,N_28033,N_27962);
and U28240 (N_28240,N_27984,N_28091);
nand U28241 (N_28241,N_28121,N_28085);
xnor U28242 (N_28242,N_28051,N_28015);
nor U28243 (N_28243,N_28023,N_27992);
nand U28244 (N_28244,N_28124,N_27910);
and U28245 (N_28245,N_27946,N_27997);
xnor U28246 (N_28246,N_28009,N_28043);
nand U28247 (N_28247,N_28002,N_28103);
nor U28248 (N_28248,N_28024,N_28014);
xor U28249 (N_28249,N_28008,N_28055);
xnor U28250 (N_28250,N_28001,N_28065);
or U28251 (N_28251,N_27903,N_28184);
nand U28252 (N_28252,N_28066,N_27952);
nand U28253 (N_28253,N_28119,N_28045);
or U28254 (N_28254,N_27965,N_28006);
nor U28255 (N_28255,N_28075,N_28042);
xor U28256 (N_28256,N_27925,N_27933);
and U28257 (N_28257,N_28198,N_28087);
nor U28258 (N_28258,N_27971,N_27947);
and U28259 (N_28259,N_28132,N_28154);
or U28260 (N_28260,N_27940,N_27977);
xnor U28261 (N_28261,N_28027,N_28068);
nor U28262 (N_28262,N_27979,N_28030);
xor U28263 (N_28263,N_27950,N_28036);
or U28264 (N_28264,N_28019,N_28159);
or U28265 (N_28265,N_28056,N_27960);
nor U28266 (N_28266,N_28177,N_28109);
nor U28267 (N_28267,N_28112,N_27990);
nor U28268 (N_28268,N_28169,N_28174);
and U28269 (N_28269,N_28070,N_28160);
xnor U28270 (N_28270,N_27981,N_27966);
or U28271 (N_28271,N_27964,N_27914);
xnor U28272 (N_28272,N_28017,N_28084);
nand U28273 (N_28273,N_27939,N_28004);
nor U28274 (N_28274,N_28079,N_27957);
nand U28275 (N_28275,N_27942,N_28191);
xnor U28276 (N_28276,N_27935,N_28021);
nand U28277 (N_28277,N_28123,N_27953);
or U28278 (N_28278,N_28133,N_27978);
xnor U28279 (N_28279,N_28060,N_27963);
nor U28280 (N_28280,N_27922,N_27926);
xor U28281 (N_28281,N_28130,N_28022);
nand U28282 (N_28282,N_27983,N_27941);
xor U28283 (N_28283,N_28117,N_28093);
and U28284 (N_28284,N_27949,N_28155);
xnor U28285 (N_28285,N_28073,N_27927);
nor U28286 (N_28286,N_28046,N_27980);
or U28287 (N_28287,N_27995,N_28071);
nand U28288 (N_28288,N_28164,N_27901);
nor U28289 (N_28289,N_28099,N_28114);
or U28290 (N_28290,N_27902,N_28143);
xor U28291 (N_28291,N_27959,N_27972);
or U28292 (N_28292,N_27928,N_27917);
and U28293 (N_28293,N_28186,N_28098);
and U28294 (N_28294,N_28077,N_28038);
and U28295 (N_28295,N_27905,N_28156);
or U28296 (N_28296,N_27906,N_28081);
or U28297 (N_28297,N_28170,N_28108);
or U28298 (N_28298,N_28053,N_28118);
nand U28299 (N_28299,N_28054,N_27974);
or U28300 (N_28300,N_27955,N_27961);
xnor U28301 (N_28301,N_27956,N_28031);
nor U28302 (N_28302,N_28067,N_27991);
and U28303 (N_28303,N_28037,N_27919);
xor U28304 (N_28304,N_28115,N_27998);
nor U28305 (N_28305,N_28113,N_27929);
nand U28306 (N_28306,N_27967,N_28062);
nand U28307 (N_28307,N_28150,N_28044);
and U28308 (N_28308,N_28047,N_27948);
and U28309 (N_28309,N_28088,N_28152);
and U28310 (N_28310,N_27937,N_28182);
nand U28311 (N_28311,N_28172,N_27909);
nor U28312 (N_28312,N_27923,N_28107);
nand U28313 (N_28313,N_28058,N_27932);
or U28314 (N_28314,N_27969,N_28144);
nand U28315 (N_28315,N_28171,N_28151);
xor U28316 (N_28316,N_28096,N_27993);
nand U28317 (N_28317,N_27918,N_27911);
and U28318 (N_28318,N_27916,N_28097);
nand U28319 (N_28319,N_28126,N_27900);
nor U28320 (N_28320,N_28167,N_28120);
nor U28321 (N_28321,N_27904,N_28074);
nand U28322 (N_28322,N_28100,N_28173);
xor U28323 (N_28323,N_28165,N_28035);
nand U28324 (N_28324,N_28127,N_28090);
nand U28325 (N_28325,N_28101,N_28034);
nor U28326 (N_28326,N_27944,N_28128);
or U28327 (N_28327,N_28102,N_28026);
xnor U28328 (N_28328,N_28064,N_28029);
or U28329 (N_28329,N_28050,N_28020);
nand U28330 (N_28330,N_28135,N_28110);
and U28331 (N_28331,N_28061,N_27924);
nor U28332 (N_28332,N_28199,N_27943);
xor U28333 (N_28333,N_28189,N_28142);
nand U28334 (N_28334,N_28179,N_28157);
xor U28335 (N_28335,N_28018,N_27970);
or U28336 (N_28336,N_28166,N_28138);
nand U28337 (N_28337,N_28134,N_27912);
or U28338 (N_28338,N_28106,N_28131);
or U28339 (N_28339,N_28104,N_28082);
or U28340 (N_28340,N_28141,N_27999);
and U28341 (N_28341,N_28059,N_28195);
nor U28342 (N_28342,N_28181,N_27996);
nand U28343 (N_28343,N_28194,N_28078);
nand U28344 (N_28344,N_28136,N_28122);
xor U28345 (N_28345,N_28175,N_27986);
or U28346 (N_28346,N_28153,N_27976);
and U28347 (N_28347,N_28180,N_27907);
xnor U28348 (N_28348,N_28168,N_27945);
or U28349 (N_28349,N_28129,N_28049);
xnor U28350 (N_28350,N_27985,N_28172);
xnor U28351 (N_28351,N_27933,N_27939);
nor U28352 (N_28352,N_27909,N_28156);
and U28353 (N_28353,N_28153,N_27902);
xor U28354 (N_28354,N_28119,N_28134);
xnor U28355 (N_28355,N_28152,N_28028);
and U28356 (N_28356,N_28046,N_28028);
xor U28357 (N_28357,N_28081,N_28164);
nor U28358 (N_28358,N_28143,N_27941);
and U28359 (N_28359,N_27909,N_27967);
nand U28360 (N_28360,N_27980,N_27978);
and U28361 (N_28361,N_28193,N_28092);
xor U28362 (N_28362,N_28031,N_28051);
and U28363 (N_28363,N_27930,N_27963);
or U28364 (N_28364,N_28151,N_28093);
xnor U28365 (N_28365,N_28140,N_27923);
xor U28366 (N_28366,N_28000,N_28161);
and U28367 (N_28367,N_28006,N_28094);
and U28368 (N_28368,N_28152,N_28012);
xor U28369 (N_28369,N_28095,N_28104);
and U28370 (N_28370,N_27986,N_28121);
xor U28371 (N_28371,N_27927,N_28018);
nand U28372 (N_28372,N_28128,N_28031);
and U28373 (N_28373,N_28030,N_27913);
and U28374 (N_28374,N_27912,N_28120);
xor U28375 (N_28375,N_28054,N_28049);
xnor U28376 (N_28376,N_27973,N_28068);
and U28377 (N_28377,N_27919,N_27945);
xor U28378 (N_28378,N_28176,N_27953);
xor U28379 (N_28379,N_27972,N_28121);
xor U28380 (N_28380,N_28046,N_28111);
and U28381 (N_28381,N_28109,N_28134);
nand U28382 (N_28382,N_28084,N_28106);
nand U28383 (N_28383,N_28030,N_27903);
or U28384 (N_28384,N_28171,N_27915);
nand U28385 (N_28385,N_27931,N_28050);
nor U28386 (N_28386,N_28173,N_27970);
nor U28387 (N_28387,N_27904,N_28052);
or U28388 (N_28388,N_27973,N_28096);
nor U28389 (N_28389,N_28025,N_28174);
nor U28390 (N_28390,N_27917,N_28031);
nor U28391 (N_28391,N_27959,N_28048);
and U28392 (N_28392,N_28198,N_28161);
nand U28393 (N_28393,N_28171,N_28113);
xor U28394 (N_28394,N_28149,N_27925);
or U28395 (N_28395,N_27978,N_28058);
nor U28396 (N_28396,N_28020,N_28086);
nor U28397 (N_28397,N_27910,N_28163);
and U28398 (N_28398,N_27903,N_27966);
and U28399 (N_28399,N_27956,N_28054);
xor U28400 (N_28400,N_28019,N_27982);
or U28401 (N_28401,N_28144,N_27919);
nand U28402 (N_28402,N_28035,N_27915);
nand U28403 (N_28403,N_27949,N_28150);
or U28404 (N_28404,N_28146,N_27988);
or U28405 (N_28405,N_28081,N_28196);
nor U28406 (N_28406,N_28189,N_27913);
nand U28407 (N_28407,N_28120,N_28148);
or U28408 (N_28408,N_28164,N_28078);
nand U28409 (N_28409,N_27905,N_27956);
or U28410 (N_28410,N_28048,N_28138);
or U28411 (N_28411,N_27972,N_28090);
nor U28412 (N_28412,N_27961,N_28051);
nor U28413 (N_28413,N_28047,N_27943);
nand U28414 (N_28414,N_28079,N_27958);
nand U28415 (N_28415,N_28072,N_27980);
nor U28416 (N_28416,N_27997,N_28060);
nand U28417 (N_28417,N_27950,N_28072);
xor U28418 (N_28418,N_27976,N_28118);
xnor U28419 (N_28419,N_28127,N_28021);
xnor U28420 (N_28420,N_28144,N_27996);
xnor U28421 (N_28421,N_28013,N_28151);
or U28422 (N_28422,N_28086,N_28141);
nand U28423 (N_28423,N_28033,N_28072);
or U28424 (N_28424,N_28168,N_28124);
nand U28425 (N_28425,N_27957,N_28166);
xor U28426 (N_28426,N_28188,N_27944);
nor U28427 (N_28427,N_28174,N_27974);
or U28428 (N_28428,N_28179,N_28169);
xor U28429 (N_28429,N_28178,N_27983);
and U28430 (N_28430,N_28138,N_28019);
xnor U28431 (N_28431,N_27900,N_28116);
or U28432 (N_28432,N_28185,N_28019);
or U28433 (N_28433,N_28157,N_27914);
nand U28434 (N_28434,N_28093,N_27983);
and U28435 (N_28435,N_28044,N_28062);
nor U28436 (N_28436,N_28094,N_28022);
nor U28437 (N_28437,N_28023,N_28132);
nand U28438 (N_28438,N_28158,N_28009);
nor U28439 (N_28439,N_28102,N_27951);
and U28440 (N_28440,N_28161,N_27992);
and U28441 (N_28441,N_27956,N_28169);
nor U28442 (N_28442,N_28081,N_28130);
xnor U28443 (N_28443,N_27952,N_28160);
xnor U28444 (N_28444,N_27939,N_28176);
and U28445 (N_28445,N_27954,N_28130);
and U28446 (N_28446,N_28143,N_28114);
or U28447 (N_28447,N_27904,N_28054);
and U28448 (N_28448,N_28010,N_28115);
and U28449 (N_28449,N_28179,N_28048);
nand U28450 (N_28450,N_28122,N_28174);
or U28451 (N_28451,N_27910,N_27918);
nand U28452 (N_28452,N_28191,N_28149);
or U28453 (N_28453,N_28094,N_27944);
nor U28454 (N_28454,N_28155,N_28011);
xnor U28455 (N_28455,N_28154,N_28016);
and U28456 (N_28456,N_28161,N_27975);
and U28457 (N_28457,N_28160,N_28177);
xnor U28458 (N_28458,N_27939,N_28177);
xnor U28459 (N_28459,N_28025,N_28077);
nor U28460 (N_28460,N_27905,N_28092);
xnor U28461 (N_28461,N_28057,N_27994);
xnor U28462 (N_28462,N_27939,N_27970);
nand U28463 (N_28463,N_27935,N_28007);
or U28464 (N_28464,N_27935,N_28127);
xor U28465 (N_28465,N_28048,N_27955);
nor U28466 (N_28466,N_28134,N_27928);
nor U28467 (N_28467,N_28016,N_28117);
and U28468 (N_28468,N_28014,N_28055);
nor U28469 (N_28469,N_28167,N_28125);
xor U28470 (N_28470,N_27952,N_28031);
and U28471 (N_28471,N_28183,N_28166);
and U28472 (N_28472,N_27935,N_28172);
and U28473 (N_28473,N_28040,N_27958);
nand U28474 (N_28474,N_28030,N_28032);
xnor U28475 (N_28475,N_28139,N_28055);
nand U28476 (N_28476,N_28109,N_28100);
nor U28477 (N_28477,N_28059,N_28129);
nor U28478 (N_28478,N_28079,N_28106);
and U28479 (N_28479,N_28108,N_28174);
or U28480 (N_28480,N_27918,N_27929);
or U28481 (N_28481,N_27912,N_27952);
xor U28482 (N_28482,N_28191,N_27946);
and U28483 (N_28483,N_27997,N_28164);
or U28484 (N_28484,N_28123,N_28026);
and U28485 (N_28485,N_27993,N_27994);
nand U28486 (N_28486,N_28136,N_27954);
nor U28487 (N_28487,N_27950,N_28101);
and U28488 (N_28488,N_27953,N_28032);
or U28489 (N_28489,N_28183,N_27975);
nor U28490 (N_28490,N_27949,N_28037);
or U28491 (N_28491,N_27905,N_27958);
nand U28492 (N_28492,N_28078,N_27967);
nor U28493 (N_28493,N_28076,N_27940);
xnor U28494 (N_28494,N_28180,N_28146);
or U28495 (N_28495,N_27953,N_28096);
and U28496 (N_28496,N_28126,N_28028);
and U28497 (N_28497,N_27992,N_27949);
xor U28498 (N_28498,N_28150,N_27914);
nand U28499 (N_28499,N_28075,N_28019);
nand U28500 (N_28500,N_28357,N_28263);
xor U28501 (N_28501,N_28283,N_28373);
and U28502 (N_28502,N_28251,N_28424);
and U28503 (N_28503,N_28402,N_28480);
or U28504 (N_28504,N_28366,N_28205);
nor U28505 (N_28505,N_28475,N_28498);
nand U28506 (N_28506,N_28355,N_28278);
nor U28507 (N_28507,N_28306,N_28238);
nor U28508 (N_28508,N_28378,N_28374);
nand U28509 (N_28509,N_28453,N_28420);
nand U28510 (N_28510,N_28339,N_28376);
xnor U28511 (N_28511,N_28409,N_28232);
and U28512 (N_28512,N_28380,N_28484);
nand U28513 (N_28513,N_28298,N_28328);
or U28514 (N_28514,N_28259,N_28395);
xor U28515 (N_28515,N_28343,N_28211);
or U28516 (N_28516,N_28220,N_28391);
nor U28517 (N_28517,N_28419,N_28264);
or U28518 (N_28518,N_28323,N_28370);
nand U28519 (N_28519,N_28294,N_28491);
xnor U28520 (N_28520,N_28312,N_28443);
xor U28521 (N_28521,N_28272,N_28321);
or U28522 (N_28522,N_28489,N_28449);
and U28523 (N_28523,N_28248,N_28299);
and U28524 (N_28524,N_28256,N_28478);
xor U28525 (N_28525,N_28315,N_28334);
nor U28526 (N_28526,N_28296,N_28254);
xnor U28527 (N_28527,N_28470,N_28445);
xor U28528 (N_28528,N_28274,N_28206);
xnor U28529 (N_28529,N_28403,N_28326);
and U28530 (N_28530,N_28266,N_28361);
nand U28531 (N_28531,N_28441,N_28246);
xor U28532 (N_28532,N_28280,N_28362);
and U28533 (N_28533,N_28432,N_28422);
xnor U28534 (N_28534,N_28468,N_28225);
nor U28535 (N_28535,N_28429,N_28457);
nand U28536 (N_28536,N_28310,N_28295);
nor U28537 (N_28537,N_28490,N_28301);
or U28538 (N_28538,N_28270,N_28426);
and U28539 (N_28539,N_28224,N_28269);
or U28540 (N_28540,N_28229,N_28358);
xor U28541 (N_28541,N_28327,N_28462);
and U28542 (N_28542,N_28239,N_28244);
and U28543 (N_28543,N_28253,N_28414);
nand U28544 (N_28544,N_28472,N_28316);
or U28545 (N_28545,N_28303,N_28284);
or U28546 (N_28546,N_28309,N_28320);
nand U28547 (N_28547,N_28203,N_28300);
nand U28548 (N_28548,N_28369,N_28435);
and U28549 (N_28549,N_28404,N_28433);
nand U28550 (N_28550,N_28285,N_28438);
or U28551 (N_28551,N_28337,N_28288);
nand U28552 (N_28552,N_28466,N_28455);
nor U28553 (N_28553,N_28410,N_28260);
nand U28554 (N_28554,N_28471,N_28473);
nand U28555 (N_28555,N_28247,N_28252);
or U28556 (N_28556,N_28495,N_28406);
and U28557 (N_28557,N_28249,N_28292);
xor U28558 (N_28558,N_28411,N_28407);
and U28559 (N_28559,N_28336,N_28387);
nor U28560 (N_28560,N_28493,N_28405);
xor U28561 (N_28561,N_28324,N_28463);
and U28562 (N_28562,N_28467,N_28322);
xor U28563 (N_28563,N_28261,N_28352);
nor U28564 (N_28564,N_28483,N_28282);
or U28565 (N_28565,N_28332,N_28434);
nor U28566 (N_28566,N_28331,N_28267);
xor U28567 (N_28567,N_28442,N_28318);
or U28568 (N_28568,N_28215,N_28250);
nor U28569 (N_28569,N_28354,N_28234);
or U28570 (N_28570,N_28221,N_28446);
xor U28571 (N_28571,N_28338,N_28486);
nand U28572 (N_28572,N_28329,N_28268);
nor U28573 (N_28573,N_28459,N_28330);
nor U28574 (N_28574,N_28262,N_28233);
or U28575 (N_28575,N_28368,N_28437);
nor U28576 (N_28576,N_28202,N_28451);
or U28577 (N_28577,N_28436,N_28237);
xor U28578 (N_28578,N_28412,N_28485);
nand U28579 (N_28579,N_28364,N_28384);
and U28580 (N_28580,N_28440,N_28290);
nand U28581 (N_28581,N_28381,N_28235);
and U28582 (N_28582,N_28350,N_28319);
or U28583 (N_28583,N_28346,N_28207);
xnor U28584 (N_28584,N_28494,N_28265);
or U28585 (N_28585,N_28421,N_28297);
xnor U28586 (N_28586,N_28231,N_28481);
and U28587 (N_28587,N_28450,N_28372);
or U28588 (N_28588,N_28499,N_28476);
nor U28589 (N_28589,N_28230,N_28277);
xnor U28590 (N_28590,N_28214,N_28305);
nor U28591 (N_28591,N_28360,N_28200);
and U28592 (N_28592,N_28430,N_28496);
nor U28593 (N_28593,N_28488,N_28210);
and U28594 (N_28594,N_28317,N_28417);
nor U28595 (N_28595,N_28273,N_28344);
xnor U28596 (N_28596,N_28477,N_28257);
and U28597 (N_28597,N_28311,N_28439);
nor U28598 (N_28598,N_28345,N_28394);
and U28599 (N_28599,N_28347,N_28335);
nand U28600 (N_28600,N_28213,N_28474);
and U28601 (N_28601,N_28465,N_28286);
and U28602 (N_28602,N_28314,N_28218);
and U28603 (N_28603,N_28386,N_28341);
nand U28604 (N_28604,N_28241,N_28464);
xnor U28605 (N_28605,N_28275,N_28397);
or U28606 (N_28606,N_28392,N_28313);
and U28607 (N_28607,N_28271,N_28209);
or U28608 (N_28608,N_28389,N_28293);
nand U28609 (N_28609,N_28398,N_28227);
xnor U28610 (N_28610,N_28418,N_28431);
xor U28611 (N_28611,N_28460,N_28348);
or U28612 (N_28612,N_28359,N_28236);
and U28613 (N_28613,N_28255,N_28365);
and U28614 (N_28614,N_28408,N_28212);
nand U28615 (N_28615,N_28388,N_28276);
xor U28616 (N_28616,N_28349,N_28492);
nand U28617 (N_28617,N_28302,N_28219);
nor U28618 (N_28618,N_28427,N_28371);
or U28619 (N_28619,N_28356,N_28379);
and U28620 (N_28620,N_28245,N_28390);
nand U28621 (N_28621,N_28385,N_28479);
xor U28622 (N_28622,N_28363,N_28208);
and U28623 (N_28623,N_28325,N_28201);
nand U28624 (N_28624,N_28482,N_28423);
nor U28625 (N_28625,N_28458,N_28353);
and U28626 (N_28626,N_28307,N_28223);
nor U28627 (N_28627,N_28279,N_28204);
nor U28628 (N_28628,N_28377,N_28242);
or U28629 (N_28629,N_28226,N_28456);
and U28630 (N_28630,N_28287,N_28469);
xnor U28631 (N_28631,N_28497,N_28382);
nand U28632 (N_28632,N_28217,N_28222);
nor U28633 (N_28633,N_28400,N_28228);
or U28634 (N_28634,N_28240,N_28304);
nor U28635 (N_28635,N_28461,N_28448);
xnor U28636 (N_28636,N_28308,N_28281);
nor U28637 (N_28637,N_28367,N_28243);
and U28638 (N_28638,N_28416,N_28258);
or U28639 (N_28639,N_28425,N_28393);
xnor U28640 (N_28640,N_28342,N_28289);
xnor U28641 (N_28641,N_28401,N_28428);
xor U28642 (N_28642,N_28396,N_28452);
nand U28643 (N_28643,N_28415,N_28399);
nor U28644 (N_28644,N_28444,N_28375);
nor U28645 (N_28645,N_28383,N_28216);
and U28646 (N_28646,N_28333,N_28487);
and U28647 (N_28647,N_28351,N_28340);
and U28648 (N_28648,N_28291,N_28447);
xor U28649 (N_28649,N_28413,N_28454);
nor U28650 (N_28650,N_28261,N_28493);
and U28651 (N_28651,N_28458,N_28422);
and U28652 (N_28652,N_28289,N_28385);
and U28653 (N_28653,N_28321,N_28364);
and U28654 (N_28654,N_28222,N_28463);
nor U28655 (N_28655,N_28289,N_28445);
nor U28656 (N_28656,N_28379,N_28237);
nand U28657 (N_28657,N_28274,N_28359);
and U28658 (N_28658,N_28327,N_28415);
and U28659 (N_28659,N_28206,N_28395);
nand U28660 (N_28660,N_28482,N_28224);
nor U28661 (N_28661,N_28410,N_28443);
or U28662 (N_28662,N_28316,N_28245);
or U28663 (N_28663,N_28462,N_28416);
or U28664 (N_28664,N_28221,N_28303);
nor U28665 (N_28665,N_28269,N_28348);
nand U28666 (N_28666,N_28486,N_28480);
nor U28667 (N_28667,N_28472,N_28274);
nand U28668 (N_28668,N_28470,N_28375);
nor U28669 (N_28669,N_28443,N_28277);
and U28670 (N_28670,N_28200,N_28314);
xnor U28671 (N_28671,N_28286,N_28489);
or U28672 (N_28672,N_28399,N_28478);
nor U28673 (N_28673,N_28347,N_28465);
or U28674 (N_28674,N_28237,N_28367);
or U28675 (N_28675,N_28415,N_28393);
and U28676 (N_28676,N_28423,N_28471);
xnor U28677 (N_28677,N_28455,N_28381);
nor U28678 (N_28678,N_28465,N_28236);
nand U28679 (N_28679,N_28475,N_28289);
or U28680 (N_28680,N_28345,N_28434);
or U28681 (N_28681,N_28458,N_28461);
or U28682 (N_28682,N_28414,N_28257);
or U28683 (N_28683,N_28497,N_28360);
nor U28684 (N_28684,N_28485,N_28276);
and U28685 (N_28685,N_28294,N_28470);
or U28686 (N_28686,N_28332,N_28201);
nor U28687 (N_28687,N_28339,N_28468);
nor U28688 (N_28688,N_28277,N_28458);
and U28689 (N_28689,N_28280,N_28247);
nor U28690 (N_28690,N_28240,N_28395);
xnor U28691 (N_28691,N_28254,N_28498);
nor U28692 (N_28692,N_28449,N_28484);
nand U28693 (N_28693,N_28279,N_28317);
nor U28694 (N_28694,N_28207,N_28301);
and U28695 (N_28695,N_28294,N_28431);
nand U28696 (N_28696,N_28235,N_28471);
nand U28697 (N_28697,N_28392,N_28248);
xor U28698 (N_28698,N_28384,N_28475);
nor U28699 (N_28699,N_28381,N_28280);
or U28700 (N_28700,N_28244,N_28328);
and U28701 (N_28701,N_28477,N_28318);
and U28702 (N_28702,N_28411,N_28286);
nor U28703 (N_28703,N_28260,N_28258);
and U28704 (N_28704,N_28214,N_28482);
xnor U28705 (N_28705,N_28350,N_28394);
nand U28706 (N_28706,N_28499,N_28249);
nand U28707 (N_28707,N_28480,N_28463);
nand U28708 (N_28708,N_28208,N_28346);
and U28709 (N_28709,N_28477,N_28242);
nor U28710 (N_28710,N_28268,N_28221);
nor U28711 (N_28711,N_28300,N_28485);
nor U28712 (N_28712,N_28398,N_28200);
and U28713 (N_28713,N_28393,N_28299);
nand U28714 (N_28714,N_28488,N_28495);
or U28715 (N_28715,N_28242,N_28343);
nor U28716 (N_28716,N_28419,N_28435);
nor U28717 (N_28717,N_28373,N_28341);
nor U28718 (N_28718,N_28403,N_28402);
or U28719 (N_28719,N_28223,N_28362);
or U28720 (N_28720,N_28482,N_28202);
nand U28721 (N_28721,N_28445,N_28400);
and U28722 (N_28722,N_28213,N_28270);
and U28723 (N_28723,N_28444,N_28473);
or U28724 (N_28724,N_28394,N_28267);
nor U28725 (N_28725,N_28360,N_28405);
xnor U28726 (N_28726,N_28213,N_28432);
xor U28727 (N_28727,N_28242,N_28307);
nor U28728 (N_28728,N_28486,N_28411);
or U28729 (N_28729,N_28278,N_28494);
or U28730 (N_28730,N_28418,N_28359);
nor U28731 (N_28731,N_28294,N_28414);
xnor U28732 (N_28732,N_28289,N_28420);
nand U28733 (N_28733,N_28424,N_28311);
xnor U28734 (N_28734,N_28438,N_28471);
nor U28735 (N_28735,N_28345,N_28231);
nand U28736 (N_28736,N_28401,N_28346);
xor U28737 (N_28737,N_28295,N_28234);
and U28738 (N_28738,N_28205,N_28387);
nor U28739 (N_28739,N_28285,N_28429);
and U28740 (N_28740,N_28447,N_28445);
and U28741 (N_28741,N_28204,N_28297);
and U28742 (N_28742,N_28285,N_28302);
or U28743 (N_28743,N_28478,N_28458);
nor U28744 (N_28744,N_28237,N_28322);
and U28745 (N_28745,N_28490,N_28455);
nand U28746 (N_28746,N_28464,N_28385);
or U28747 (N_28747,N_28453,N_28299);
or U28748 (N_28748,N_28447,N_28283);
nor U28749 (N_28749,N_28426,N_28421);
nor U28750 (N_28750,N_28446,N_28301);
nor U28751 (N_28751,N_28268,N_28465);
xor U28752 (N_28752,N_28473,N_28408);
nor U28753 (N_28753,N_28332,N_28341);
and U28754 (N_28754,N_28436,N_28246);
xnor U28755 (N_28755,N_28279,N_28346);
xnor U28756 (N_28756,N_28421,N_28362);
nand U28757 (N_28757,N_28458,N_28201);
nor U28758 (N_28758,N_28219,N_28323);
xnor U28759 (N_28759,N_28476,N_28467);
or U28760 (N_28760,N_28408,N_28494);
and U28761 (N_28761,N_28369,N_28304);
or U28762 (N_28762,N_28369,N_28321);
xnor U28763 (N_28763,N_28419,N_28210);
nor U28764 (N_28764,N_28487,N_28287);
and U28765 (N_28765,N_28425,N_28398);
xnor U28766 (N_28766,N_28313,N_28289);
nand U28767 (N_28767,N_28276,N_28492);
xnor U28768 (N_28768,N_28238,N_28337);
nor U28769 (N_28769,N_28313,N_28219);
nor U28770 (N_28770,N_28375,N_28384);
nand U28771 (N_28771,N_28375,N_28202);
xor U28772 (N_28772,N_28290,N_28232);
xnor U28773 (N_28773,N_28222,N_28394);
nand U28774 (N_28774,N_28465,N_28298);
and U28775 (N_28775,N_28237,N_28417);
and U28776 (N_28776,N_28471,N_28487);
and U28777 (N_28777,N_28368,N_28228);
nand U28778 (N_28778,N_28242,N_28400);
xor U28779 (N_28779,N_28321,N_28405);
or U28780 (N_28780,N_28376,N_28245);
and U28781 (N_28781,N_28348,N_28216);
nor U28782 (N_28782,N_28443,N_28458);
and U28783 (N_28783,N_28349,N_28287);
nor U28784 (N_28784,N_28381,N_28322);
or U28785 (N_28785,N_28406,N_28309);
or U28786 (N_28786,N_28426,N_28466);
nor U28787 (N_28787,N_28224,N_28442);
or U28788 (N_28788,N_28330,N_28219);
nor U28789 (N_28789,N_28286,N_28234);
or U28790 (N_28790,N_28340,N_28421);
or U28791 (N_28791,N_28467,N_28328);
nand U28792 (N_28792,N_28422,N_28273);
xnor U28793 (N_28793,N_28383,N_28430);
nor U28794 (N_28794,N_28239,N_28314);
nor U28795 (N_28795,N_28271,N_28259);
xor U28796 (N_28796,N_28219,N_28417);
nor U28797 (N_28797,N_28426,N_28360);
and U28798 (N_28798,N_28346,N_28212);
nor U28799 (N_28799,N_28284,N_28361);
xnor U28800 (N_28800,N_28516,N_28561);
nand U28801 (N_28801,N_28753,N_28669);
nand U28802 (N_28802,N_28577,N_28554);
and U28803 (N_28803,N_28694,N_28757);
nor U28804 (N_28804,N_28506,N_28736);
xnor U28805 (N_28805,N_28545,N_28735);
and U28806 (N_28806,N_28541,N_28713);
xnor U28807 (N_28807,N_28575,N_28630);
nor U28808 (N_28808,N_28754,N_28774);
xor U28809 (N_28809,N_28725,N_28567);
and U28810 (N_28810,N_28631,N_28717);
or U28811 (N_28811,N_28660,N_28624);
nand U28812 (N_28812,N_28626,N_28731);
nor U28813 (N_28813,N_28509,N_28776);
xor U28814 (N_28814,N_28772,N_28536);
nor U28815 (N_28815,N_28513,N_28512);
or U28816 (N_28816,N_28708,N_28720);
nand U28817 (N_28817,N_28639,N_28691);
nand U28818 (N_28818,N_28778,N_28766);
or U28819 (N_28819,N_28632,N_28685);
and U28820 (N_28820,N_28703,N_28668);
nand U28821 (N_28821,N_28553,N_28585);
xor U28822 (N_28822,N_28662,N_28781);
nor U28823 (N_28823,N_28565,N_28570);
nand U28824 (N_28824,N_28534,N_28681);
and U28825 (N_28825,N_28756,N_28775);
or U28826 (N_28826,N_28700,N_28738);
and U28827 (N_28827,N_28664,N_28785);
and U28828 (N_28828,N_28790,N_28605);
nand U28829 (N_28829,N_28634,N_28622);
or U28830 (N_28830,N_28610,N_28796);
xor U28831 (N_28831,N_28792,N_28500);
nand U28832 (N_28832,N_28549,N_28633);
and U28833 (N_28833,N_28560,N_28556);
nand U28834 (N_28834,N_28688,N_28544);
nor U28835 (N_28835,N_28730,N_28629);
and U28836 (N_28836,N_28797,N_28592);
nor U28837 (N_28837,N_28583,N_28572);
xnor U28838 (N_28838,N_28701,N_28793);
or U28839 (N_28839,N_28711,N_28682);
or U28840 (N_28840,N_28520,N_28759);
and U28841 (N_28841,N_28523,N_28696);
nand U28842 (N_28842,N_28623,N_28543);
nor U28843 (N_28843,N_28697,N_28604);
or U28844 (N_28844,N_28657,N_28744);
or U28845 (N_28845,N_28666,N_28663);
and U28846 (N_28846,N_28539,N_28524);
or U28847 (N_28847,N_28745,N_28773);
nand U28848 (N_28848,N_28680,N_28538);
and U28849 (N_28849,N_28677,N_28522);
and U28850 (N_28850,N_28727,N_28530);
xor U28851 (N_28851,N_28593,N_28659);
xnor U28852 (N_28852,N_28587,N_28640);
nor U28853 (N_28853,N_28525,N_28508);
and U28854 (N_28854,N_28645,N_28621);
or U28855 (N_28855,N_28581,N_28737);
nor U28856 (N_28856,N_28607,N_28603);
xor U28857 (N_28857,N_28765,N_28521);
xor U28858 (N_28858,N_28704,N_28692);
nand U28859 (N_28859,N_28588,N_28602);
nand U28860 (N_28860,N_28620,N_28547);
xor U28861 (N_28861,N_28637,N_28722);
nand U28862 (N_28862,N_28515,N_28580);
or U28863 (N_28863,N_28594,N_28689);
nor U28864 (N_28864,N_28528,N_28779);
and U28865 (N_28865,N_28728,N_28606);
nor U28866 (N_28866,N_28746,N_28769);
or U28867 (N_28867,N_28732,N_28527);
and U28868 (N_28868,N_28579,N_28743);
xnor U28869 (N_28869,N_28546,N_28559);
nand U28870 (N_28870,N_28652,N_28503);
xor U28871 (N_28871,N_28517,N_28676);
nand U28872 (N_28872,N_28670,N_28558);
nor U28873 (N_28873,N_28724,N_28684);
xnor U28874 (N_28874,N_28742,N_28519);
xnor U28875 (N_28875,N_28693,N_28569);
and U28876 (N_28876,N_28618,N_28564);
xor U28877 (N_28877,N_28761,N_28672);
or U28878 (N_28878,N_28683,N_28532);
and U28879 (N_28879,N_28649,N_28609);
or U28880 (N_28880,N_28574,N_28787);
and U28881 (N_28881,N_28502,N_28535);
nor U28882 (N_28882,N_28750,N_28795);
or U28883 (N_28883,N_28542,N_28642);
nor U28884 (N_28884,N_28673,N_28599);
nor U28885 (N_28885,N_28763,N_28709);
nand U28886 (N_28886,N_28764,N_28627);
nor U28887 (N_28887,N_28638,N_28576);
xor U28888 (N_28888,N_28595,N_28699);
nor U28889 (N_28889,N_28518,N_28655);
xnor U28890 (N_28890,N_28733,N_28507);
xor U28891 (N_28891,N_28562,N_28628);
nor U28892 (N_28892,N_28767,N_28589);
xor U28893 (N_28893,N_28695,N_28719);
nand U28894 (N_28894,N_28770,N_28705);
or U28895 (N_28895,N_28718,N_28531);
nand U28896 (N_28896,N_28721,N_28715);
and U28897 (N_28897,N_28714,N_28636);
and U28898 (N_28898,N_28557,N_28784);
xnor U28899 (N_28899,N_28511,N_28504);
xor U28900 (N_28900,N_28798,N_28702);
xnor U28901 (N_28901,N_28537,N_28749);
xor U28902 (N_28902,N_28578,N_28726);
or U28903 (N_28903,N_28739,N_28729);
or U28904 (N_28904,N_28679,N_28706);
and U28905 (N_28905,N_28658,N_28586);
nand U28906 (N_28906,N_28617,N_28780);
or U28907 (N_28907,N_28619,N_28650);
xor U28908 (N_28908,N_28648,N_28789);
and U28909 (N_28909,N_28551,N_28686);
or U28910 (N_28910,N_28678,N_28591);
nor U28911 (N_28911,N_28665,N_28646);
or U28912 (N_28912,N_28651,N_28616);
nand U28913 (N_28913,N_28687,N_28615);
nand U28914 (N_28914,N_28698,N_28751);
nand U28915 (N_28915,N_28654,N_28526);
xnor U28916 (N_28916,N_28771,N_28661);
nand U28917 (N_28917,N_28741,N_28710);
nand U28918 (N_28918,N_28613,N_28748);
nand U28919 (N_28919,N_28671,N_28791);
nand U28920 (N_28920,N_28734,N_28644);
xor U28921 (N_28921,N_28777,N_28600);
or U28922 (N_28922,N_28501,N_28788);
and U28923 (N_28923,N_28582,N_28740);
nand U28924 (N_28924,N_28601,N_28573);
xnor U28925 (N_28925,N_28794,N_28635);
xor U28926 (N_28926,N_28643,N_28675);
xnor U28927 (N_28927,N_28690,N_28656);
nor U28928 (N_28928,N_28598,N_28552);
and U28929 (N_28929,N_28674,N_28653);
and U28930 (N_28930,N_28548,N_28760);
or U28931 (N_28931,N_28762,N_28590);
xnor U28932 (N_28932,N_28571,N_28563);
or U28933 (N_28933,N_28614,N_28782);
nand U28934 (N_28934,N_28783,N_28799);
xor U28935 (N_28935,N_28716,N_28596);
or U28936 (N_28936,N_28568,N_28608);
and U28937 (N_28937,N_28641,N_28747);
nor U28938 (N_28938,N_28768,N_28625);
or U28939 (N_28939,N_28647,N_28597);
nor U28940 (N_28940,N_28505,N_28510);
and U28941 (N_28941,N_28612,N_28584);
nor U28942 (N_28942,N_28707,N_28555);
and U28943 (N_28943,N_28533,N_28758);
xnor U28944 (N_28944,N_28667,N_28752);
and U28945 (N_28945,N_28611,N_28723);
nand U28946 (N_28946,N_28514,N_28755);
and U28947 (N_28947,N_28786,N_28529);
xor U28948 (N_28948,N_28550,N_28540);
xnor U28949 (N_28949,N_28712,N_28566);
or U28950 (N_28950,N_28572,N_28799);
or U28951 (N_28951,N_28791,N_28763);
or U28952 (N_28952,N_28598,N_28775);
nand U28953 (N_28953,N_28526,N_28541);
and U28954 (N_28954,N_28771,N_28533);
xnor U28955 (N_28955,N_28738,N_28705);
and U28956 (N_28956,N_28735,N_28609);
and U28957 (N_28957,N_28540,N_28513);
nor U28958 (N_28958,N_28717,N_28514);
nor U28959 (N_28959,N_28792,N_28788);
or U28960 (N_28960,N_28635,N_28660);
nand U28961 (N_28961,N_28678,N_28719);
or U28962 (N_28962,N_28648,N_28680);
nor U28963 (N_28963,N_28796,N_28747);
nand U28964 (N_28964,N_28552,N_28506);
xnor U28965 (N_28965,N_28661,N_28645);
nor U28966 (N_28966,N_28634,N_28762);
xnor U28967 (N_28967,N_28701,N_28555);
nor U28968 (N_28968,N_28679,N_28778);
nor U28969 (N_28969,N_28524,N_28525);
nand U28970 (N_28970,N_28577,N_28675);
nand U28971 (N_28971,N_28716,N_28749);
xnor U28972 (N_28972,N_28547,N_28519);
nand U28973 (N_28973,N_28693,N_28783);
nor U28974 (N_28974,N_28627,N_28637);
or U28975 (N_28975,N_28612,N_28741);
or U28976 (N_28976,N_28507,N_28561);
nor U28977 (N_28977,N_28507,N_28697);
or U28978 (N_28978,N_28723,N_28748);
and U28979 (N_28979,N_28693,N_28584);
and U28980 (N_28980,N_28693,N_28560);
nand U28981 (N_28981,N_28698,N_28716);
nor U28982 (N_28982,N_28626,N_28535);
and U28983 (N_28983,N_28726,N_28793);
nor U28984 (N_28984,N_28728,N_28782);
xnor U28985 (N_28985,N_28571,N_28598);
nor U28986 (N_28986,N_28672,N_28791);
nand U28987 (N_28987,N_28758,N_28575);
and U28988 (N_28988,N_28678,N_28798);
nor U28989 (N_28989,N_28685,N_28784);
or U28990 (N_28990,N_28746,N_28657);
and U28991 (N_28991,N_28570,N_28588);
or U28992 (N_28992,N_28752,N_28780);
and U28993 (N_28993,N_28694,N_28728);
nand U28994 (N_28994,N_28761,N_28742);
or U28995 (N_28995,N_28620,N_28651);
nand U28996 (N_28996,N_28710,N_28563);
xor U28997 (N_28997,N_28587,N_28745);
xnor U28998 (N_28998,N_28659,N_28741);
xnor U28999 (N_28999,N_28559,N_28626);
xor U29000 (N_29000,N_28660,N_28640);
and U29001 (N_29001,N_28656,N_28691);
xor U29002 (N_29002,N_28513,N_28729);
xor U29003 (N_29003,N_28648,N_28654);
xnor U29004 (N_29004,N_28535,N_28569);
nand U29005 (N_29005,N_28679,N_28780);
nor U29006 (N_29006,N_28646,N_28670);
nor U29007 (N_29007,N_28512,N_28606);
or U29008 (N_29008,N_28751,N_28773);
nand U29009 (N_29009,N_28705,N_28547);
nor U29010 (N_29010,N_28623,N_28737);
and U29011 (N_29011,N_28690,N_28606);
nor U29012 (N_29012,N_28694,N_28507);
nand U29013 (N_29013,N_28746,N_28648);
nand U29014 (N_29014,N_28689,N_28603);
and U29015 (N_29015,N_28680,N_28523);
nor U29016 (N_29016,N_28640,N_28745);
nand U29017 (N_29017,N_28662,N_28554);
nor U29018 (N_29018,N_28751,N_28723);
or U29019 (N_29019,N_28697,N_28625);
xnor U29020 (N_29020,N_28543,N_28793);
nor U29021 (N_29021,N_28508,N_28716);
nor U29022 (N_29022,N_28708,N_28694);
nand U29023 (N_29023,N_28786,N_28764);
nor U29024 (N_29024,N_28536,N_28727);
xor U29025 (N_29025,N_28724,N_28581);
or U29026 (N_29026,N_28515,N_28748);
nor U29027 (N_29027,N_28786,N_28747);
nor U29028 (N_29028,N_28597,N_28649);
nor U29029 (N_29029,N_28784,N_28508);
or U29030 (N_29030,N_28506,N_28588);
nor U29031 (N_29031,N_28688,N_28794);
nand U29032 (N_29032,N_28694,N_28675);
xor U29033 (N_29033,N_28636,N_28765);
and U29034 (N_29034,N_28737,N_28671);
xnor U29035 (N_29035,N_28712,N_28615);
nor U29036 (N_29036,N_28662,N_28543);
and U29037 (N_29037,N_28732,N_28566);
xnor U29038 (N_29038,N_28700,N_28740);
xnor U29039 (N_29039,N_28627,N_28791);
or U29040 (N_29040,N_28668,N_28596);
or U29041 (N_29041,N_28791,N_28755);
xor U29042 (N_29042,N_28557,N_28599);
and U29043 (N_29043,N_28676,N_28547);
nor U29044 (N_29044,N_28610,N_28571);
nor U29045 (N_29045,N_28553,N_28711);
nand U29046 (N_29046,N_28661,N_28714);
nand U29047 (N_29047,N_28745,N_28581);
nand U29048 (N_29048,N_28564,N_28670);
xor U29049 (N_29049,N_28587,N_28730);
xnor U29050 (N_29050,N_28629,N_28762);
nor U29051 (N_29051,N_28695,N_28773);
or U29052 (N_29052,N_28789,N_28606);
nand U29053 (N_29053,N_28641,N_28586);
xnor U29054 (N_29054,N_28768,N_28627);
xnor U29055 (N_29055,N_28775,N_28539);
and U29056 (N_29056,N_28595,N_28751);
nor U29057 (N_29057,N_28528,N_28755);
nand U29058 (N_29058,N_28510,N_28659);
nand U29059 (N_29059,N_28677,N_28501);
xor U29060 (N_29060,N_28544,N_28590);
xnor U29061 (N_29061,N_28566,N_28796);
and U29062 (N_29062,N_28583,N_28714);
nor U29063 (N_29063,N_28608,N_28682);
nand U29064 (N_29064,N_28573,N_28583);
nand U29065 (N_29065,N_28751,N_28614);
and U29066 (N_29066,N_28677,N_28520);
xor U29067 (N_29067,N_28713,N_28661);
xnor U29068 (N_29068,N_28578,N_28563);
xor U29069 (N_29069,N_28747,N_28749);
or U29070 (N_29070,N_28730,N_28707);
nand U29071 (N_29071,N_28674,N_28694);
nand U29072 (N_29072,N_28585,N_28548);
xor U29073 (N_29073,N_28520,N_28588);
and U29074 (N_29074,N_28542,N_28502);
nand U29075 (N_29075,N_28574,N_28629);
xnor U29076 (N_29076,N_28541,N_28575);
nor U29077 (N_29077,N_28543,N_28631);
nand U29078 (N_29078,N_28639,N_28698);
or U29079 (N_29079,N_28557,N_28695);
nand U29080 (N_29080,N_28559,N_28734);
nand U29081 (N_29081,N_28500,N_28504);
nand U29082 (N_29082,N_28708,N_28617);
nand U29083 (N_29083,N_28678,N_28669);
or U29084 (N_29084,N_28639,N_28731);
or U29085 (N_29085,N_28686,N_28794);
or U29086 (N_29086,N_28519,N_28671);
nand U29087 (N_29087,N_28556,N_28634);
xor U29088 (N_29088,N_28590,N_28575);
nor U29089 (N_29089,N_28765,N_28729);
nand U29090 (N_29090,N_28622,N_28540);
xnor U29091 (N_29091,N_28692,N_28648);
or U29092 (N_29092,N_28686,N_28660);
and U29093 (N_29093,N_28677,N_28602);
nand U29094 (N_29094,N_28621,N_28593);
nor U29095 (N_29095,N_28651,N_28759);
and U29096 (N_29096,N_28521,N_28557);
and U29097 (N_29097,N_28785,N_28503);
xnor U29098 (N_29098,N_28675,N_28688);
or U29099 (N_29099,N_28515,N_28661);
nand U29100 (N_29100,N_29066,N_28804);
nor U29101 (N_29101,N_28869,N_29039);
xor U29102 (N_29102,N_28932,N_28902);
nand U29103 (N_29103,N_29038,N_28921);
nand U29104 (N_29104,N_28901,N_28916);
and U29105 (N_29105,N_28977,N_28981);
nand U29106 (N_29106,N_29097,N_29021);
xor U29107 (N_29107,N_29013,N_28803);
and U29108 (N_29108,N_28988,N_29011);
or U29109 (N_29109,N_28801,N_28835);
or U29110 (N_29110,N_28883,N_28989);
nor U29111 (N_29111,N_29071,N_28959);
and U29112 (N_29112,N_28837,N_28852);
nor U29113 (N_29113,N_28866,N_29088);
and U29114 (N_29114,N_28922,N_28915);
nor U29115 (N_29115,N_29030,N_29020);
nand U29116 (N_29116,N_29026,N_28944);
nand U29117 (N_29117,N_29053,N_28984);
or U29118 (N_29118,N_28888,N_28983);
nand U29119 (N_29119,N_28817,N_29082);
nor U29120 (N_29120,N_29050,N_28996);
and U29121 (N_29121,N_28894,N_29068);
and U29122 (N_29122,N_28953,N_28820);
xor U29123 (N_29123,N_29008,N_28876);
xor U29124 (N_29124,N_28830,N_28882);
nand U29125 (N_29125,N_28923,N_28897);
nand U29126 (N_29126,N_28914,N_29081);
and U29127 (N_29127,N_29083,N_28842);
xor U29128 (N_29128,N_28937,N_28873);
nor U29129 (N_29129,N_29016,N_28995);
nand U29130 (N_29130,N_28990,N_29090);
and U29131 (N_29131,N_28956,N_29095);
nand U29132 (N_29132,N_28925,N_29073);
nor U29133 (N_29133,N_28999,N_28891);
or U29134 (N_29134,N_29061,N_28834);
or U29135 (N_29135,N_28844,N_29074);
nor U29136 (N_29136,N_29063,N_29098);
nor U29137 (N_29137,N_28965,N_28920);
and U29138 (N_29138,N_29024,N_28805);
xnor U29139 (N_29139,N_29002,N_29092);
or U29140 (N_29140,N_28853,N_28872);
and U29141 (N_29141,N_28843,N_28851);
nand U29142 (N_29142,N_29091,N_29093);
nor U29143 (N_29143,N_29052,N_28946);
xnor U29144 (N_29144,N_28960,N_28951);
xor U29145 (N_29145,N_28991,N_28870);
nand U29146 (N_29146,N_28809,N_29099);
and U29147 (N_29147,N_28945,N_28881);
and U29148 (N_29148,N_29076,N_29031);
xor U29149 (N_29149,N_28847,N_29087);
xnor U29150 (N_29150,N_28807,N_29058);
and U29151 (N_29151,N_29019,N_28821);
xor U29152 (N_29152,N_28828,N_29035);
xor U29153 (N_29153,N_28884,N_28963);
xor U29154 (N_29154,N_28855,N_28848);
or U29155 (N_29155,N_28950,N_28885);
xnor U29156 (N_29156,N_28839,N_28880);
nand U29157 (N_29157,N_28856,N_28824);
and U29158 (N_29158,N_28949,N_28926);
or U29159 (N_29159,N_29014,N_28917);
nor U29160 (N_29160,N_29051,N_28841);
xor U29161 (N_29161,N_28889,N_29006);
nor U29162 (N_29162,N_29005,N_29009);
and U29163 (N_29163,N_29094,N_28955);
and U29164 (N_29164,N_28976,N_28997);
nand U29165 (N_29165,N_28970,N_28933);
nor U29166 (N_29166,N_28961,N_28971);
nor U29167 (N_29167,N_29034,N_28936);
or U29168 (N_29168,N_29084,N_28913);
nand U29169 (N_29169,N_29079,N_28934);
xor U29170 (N_29170,N_29045,N_28877);
nand U29171 (N_29171,N_29015,N_28939);
xnor U29172 (N_29172,N_28802,N_29046);
and U29173 (N_29173,N_28979,N_28980);
nand U29174 (N_29174,N_28840,N_29043);
or U29175 (N_29175,N_28886,N_29049);
nor U29176 (N_29176,N_28985,N_28947);
xor U29177 (N_29177,N_29010,N_28867);
xnor U29178 (N_29178,N_29080,N_28857);
xnor U29179 (N_29179,N_28898,N_28968);
or U29180 (N_29180,N_28940,N_29023);
and U29181 (N_29181,N_28826,N_28819);
and U29182 (N_29182,N_29070,N_28816);
and U29183 (N_29183,N_29065,N_28928);
xor U29184 (N_29184,N_28806,N_28845);
or U29185 (N_29185,N_29040,N_29089);
xor U29186 (N_29186,N_29037,N_28957);
and U29187 (N_29187,N_28864,N_28929);
nor U29188 (N_29188,N_28994,N_29000);
and U29189 (N_29189,N_28911,N_28910);
or U29190 (N_29190,N_29075,N_28827);
and U29191 (N_29191,N_28912,N_29086);
nor U29192 (N_29192,N_28909,N_29007);
nand U29193 (N_29193,N_28874,N_29057);
xor U29194 (N_29194,N_28836,N_28800);
nor U29195 (N_29195,N_29044,N_29067);
or U29196 (N_29196,N_29042,N_28906);
nor U29197 (N_29197,N_28943,N_29059);
nand U29198 (N_29198,N_28962,N_28975);
nand U29199 (N_29199,N_29085,N_28967);
nor U29200 (N_29200,N_28859,N_28927);
nand U29201 (N_29201,N_29078,N_28854);
and U29202 (N_29202,N_29032,N_28924);
and U29203 (N_29203,N_28966,N_29064);
or U29204 (N_29204,N_28905,N_29029);
xnor U29205 (N_29205,N_28993,N_28931);
or U29206 (N_29206,N_28813,N_28948);
nor U29207 (N_29207,N_29003,N_29004);
nand U29208 (N_29208,N_28938,N_29047);
nor U29209 (N_29209,N_28814,N_28903);
or U29210 (N_29210,N_28941,N_28900);
and U29211 (N_29211,N_28904,N_28863);
xnor U29212 (N_29212,N_29055,N_28942);
xor U29213 (N_29213,N_28815,N_28810);
or U29214 (N_29214,N_28879,N_28907);
and U29215 (N_29215,N_28982,N_29001);
nand U29216 (N_29216,N_28823,N_28825);
nand U29217 (N_29217,N_28838,N_29041);
and U29218 (N_29218,N_28832,N_29012);
nand U29219 (N_29219,N_28992,N_28987);
nand U29220 (N_29220,N_28812,N_29027);
xnor U29221 (N_29221,N_29018,N_28895);
nand U29222 (N_29222,N_29096,N_28998);
nand U29223 (N_29223,N_28818,N_29036);
or U29224 (N_29224,N_28887,N_28893);
and U29225 (N_29225,N_29077,N_28964);
and U29226 (N_29226,N_28822,N_28969);
nand U29227 (N_29227,N_28846,N_29069);
nand U29228 (N_29228,N_29062,N_28935);
nor U29229 (N_29229,N_28868,N_29072);
xor U29230 (N_29230,N_28958,N_28829);
or U29231 (N_29231,N_28865,N_28986);
nand U29232 (N_29232,N_29033,N_28919);
nand U29233 (N_29233,N_28831,N_28908);
nand U29234 (N_29234,N_28972,N_28878);
and U29235 (N_29235,N_28858,N_28871);
xnor U29236 (N_29236,N_28930,N_28892);
nor U29237 (N_29237,N_29056,N_28952);
or U29238 (N_29238,N_29060,N_29017);
or U29239 (N_29239,N_29054,N_28850);
and U29240 (N_29240,N_28896,N_28899);
nor U29241 (N_29241,N_29048,N_28811);
and U29242 (N_29242,N_28978,N_28861);
or U29243 (N_29243,N_28918,N_28973);
or U29244 (N_29244,N_28954,N_28862);
nor U29245 (N_29245,N_28890,N_29028);
nand U29246 (N_29246,N_28808,N_28974);
xnor U29247 (N_29247,N_29025,N_29022);
or U29248 (N_29248,N_28860,N_28833);
nand U29249 (N_29249,N_28875,N_28849);
nand U29250 (N_29250,N_28922,N_28976);
and U29251 (N_29251,N_29015,N_29035);
or U29252 (N_29252,N_29044,N_28813);
nand U29253 (N_29253,N_28858,N_28941);
nor U29254 (N_29254,N_28835,N_28888);
nand U29255 (N_29255,N_29001,N_29095);
and U29256 (N_29256,N_28914,N_28967);
nor U29257 (N_29257,N_29065,N_29068);
or U29258 (N_29258,N_29031,N_28941);
and U29259 (N_29259,N_29075,N_28962);
nor U29260 (N_29260,N_28803,N_28839);
and U29261 (N_29261,N_29073,N_28987);
nor U29262 (N_29262,N_28908,N_28888);
nand U29263 (N_29263,N_29079,N_29091);
xnor U29264 (N_29264,N_29077,N_29040);
and U29265 (N_29265,N_29052,N_28990);
xor U29266 (N_29266,N_28957,N_29029);
or U29267 (N_29267,N_28969,N_28885);
nor U29268 (N_29268,N_28884,N_28871);
or U29269 (N_29269,N_28878,N_29042);
xnor U29270 (N_29270,N_28815,N_29078);
or U29271 (N_29271,N_28848,N_28917);
or U29272 (N_29272,N_28924,N_28908);
and U29273 (N_29273,N_29045,N_29097);
nor U29274 (N_29274,N_28990,N_28894);
nor U29275 (N_29275,N_28914,N_28884);
and U29276 (N_29276,N_29053,N_28830);
or U29277 (N_29277,N_28805,N_28909);
nand U29278 (N_29278,N_28918,N_29073);
nor U29279 (N_29279,N_29022,N_29074);
xnor U29280 (N_29280,N_28940,N_28810);
xnor U29281 (N_29281,N_28804,N_29060);
xor U29282 (N_29282,N_29088,N_28977);
nand U29283 (N_29283,N_29075,N_28820);
and U29284 (N_29284,N_28984,N_28878);
or U29285 (N_29285,N_28967,N_29091);
or U29286 (N_29286,N_28862,N_28944);
nand U29287 (N_29287,N_29043,N_28862);
and U29288 (N_29288,N_29003,N_28813);
nor U29289 (N_29289,N_29009,N_28841);
and U29290 (N_29290,N_28894,N_28884);
nor U29291 (N_29291,N_28886,N_28946);
nand U29292 (N_29292,N_28996,N_28903);
and U29293 (N_29293,N_28980,N_28932);
and U29294 (N_29294,N_28881,N_28876);
nand U29295 (N_29295,N_28948,N_28941);
nand U29296 (N_29296,N_28986,N_29083);
nor U29297 (N_29297,N_29065,N_28930);
xnor U29298 (N_29298,N_29012,N_29019);
nand U29299 (N_29299,N_28815,N_28839);
xor U29300 (N_29300,N_28968,N_28879);
nand U29301 (N_29301,N_28980,N_28879);
xor U29302 (N_29302,N_28942,N_28902);
or U29303 (N_29303,N_29053,N_29074);
nor U29304 (N_29304,N_28866,N_29078);
and U29305 (N_29305,N_29020,N_29006);
and U29306 (N_29306,N_28861,N_28833);
xor U29307 (N_29307,N_28916,N_28873);
nor U29308 (N_29308,N_29087,N_28972);
xor U29309 (N_29309,N_28835,N_28936);
nor U29310 (N_29310,N_28957,N_28857);
nor U29311 (N_29311,N_28959,N_28994);
xnor U29312 (N_29312,N_28922,N_28800);
nor U29313 (N_29313,N_28856,N_29059);
and U29314 (N_29314,N_28898,N_28815);
or U29315 (N_29315,N_28963,N_28849);
xor U29316 (N_29316,N_28840,N_28838);
xnor U29317 (N_29317,N_28985,N_28999);
or U29318 (N_29318,N_29017,N_28887);
xor U29319 (N_29319,N_28957,N_28923);
xor U29320 (N_29320,N_28956,N_28843);
nand U29321 (N_29321,N_29023,N_28813);
nand U29322 (N_29322,N_28811,N_29091);
nor U29323 (N_29323,N_28985,N_29091);
xor U29324 (N_29324,N_28885,N_29002);
and U29325 (N_29325,N_29053,N_28969);
nor U29326 (N_29326,N_28956,N_28921);
nand U29327 (N_29327,N_28943,N_28929);
nand U29328 (N_29328,N_29030,N_28967);
or U29329 (N_29329,N_28917,N_29044);
nor U29330 (N_29330,N_28896,N_28908);
and U29331 (N_29331,N_28950,N_28877);
or U29332 (N_29332,N_28838,N_28812);
and U29333 (N_29333,N_28990,N_29030);
or U29334 (N_29334,N_29085,N_29014);
and U29335 (N_29335,N_29014,N_28827);
nor U29336 (N_29336,N_29013,N_28989);
and U29337 (N_29337,N_28855,N_28867);
and U29338 (N_29338,N_28831,N_28868);
and U29339 (N_29339,N_29072,N_29017);
nand U29340 (N_29340,N_28969,N_28867);
and U29341 (N_29341,N_28959,N_28832);
nor U29342 (N_29342,N_29076,N_29050);
xor U29343 (N_29343,N_28998,N_28876);
xor U29344 (N_29344,N_28892,N_29057);
nand U29345 (N_29345,N_28945,N_28878);
xor U29346 (N_29346,N_29006,N_29001);
and U29347 (N_29347,N_28967,N_28988);
nor U29348 (N_29348,N_28887,N_28969);
or U29349 (N_29349,N_29046,N_29021);
or U29350 (N_29350,N_29001,N_28956);
nand U29351 (N_29351,N_29043,N_29081);
or U29352 (N_29352,N_28913,N_28843);
and U29353 (N_29353,N_28891,N_28996);
xnor U29354 (N_29354,N_28881,N_28995);
nor U29355 (N_29355,N_28983,N_28815);
nor U29356 (N_29356,N_28886,N_28877);
or U29357 (N_29357,N_28969,N_28957);
and U29358 (N_29358,N_28824,N_28997);
xnor U29359 (N_29359,N_28813,N_28809);
nor U29360 (N_29360,N_28826,N_28974);
or U29361 (N_29361,N_29080,N_29079);
xor U29362 (N_29362,N_28983,N_29028);
or U29363 (N_29363,N_28823,N_28959);
xor U29364 (N_29364,N_29028,N_28912);
and U29365 (N_29365,N_28883,N_29036);
xor U29366 (N_29366,N_28908,N_28976);
or U29367 (N_29367,N_28994,N_29028);
or U29368 (N_29368,N_28881,N_29038);
xor U29369 (N_29369,N_28826,N_29057);
nand U29370 (N_29370,N_28817,N_28957);
or U29371 (N_29371,N_28916,N_28997);
nand U29372 (N_29372,N_29082,N_28971);
and U29373 (N_29373,N_28922,N_29078);
xnor U29374 (N_29374,N_29021,N_28941);
nor U29375 (N_29375,N_28921,N_29028);
xnor U29376 (N_29376,N_28994,N_29035);
and U29377 (N_29377,N_28894,N_29059);
or U29378 (N_29378,N_28822,N_28850);
xnor U29379 (N_29379,N_28849,N_29036);
and U29380 (N_29380,N_29085,N_28804);
nand U29381 (N_29381,N_28945,N_29090);
and U29382 (N_29382,N_28877,N_29030);
or U29383 (N_29383,N_28820,N_28959);
and U29384 (N_29384,N_29089,N_28988);
or U29385 (N_29385,N_28924,N_28861);
xnor U29386 (N_29386,N_29099,N_28994);
nor U29387 (N_29387,N_29087,N_28970);
xor U29388 (N_29388,N_28803,N_29053);
nand U29389 (N_29389,N_28899,N_28952);
xnor U29390 (N_29390,N_28954,N_28817);
nor U29391 (N_29391,N_29026,N_28955);
and U29392 (N_29392,N_29057,N_29008);
nor U29393 (N_29393,N_28823,N_28836);
nor U29394 (N_29394,N_28845,N_28808);
nand U29395 (N_29395,N_28953,N_29077);
nand U29396 (N_29396,N_28853,N_29045);
xnor U29397 (N_29397,N_29010,N_28947);
nand U29398 (N_29398,N_29047,N_28880);
xor U29399 (N_29399,N_29020,N_28940);
nand U29400 (N_29400,N_29203,N_29181);
nor U29401 (N_29401,N_29309,N_29123);
xnor U29402 (N_29402,N_29215,N_29178);
xor U29403 (N_29403,N_29352,N_29354);
nor U29404 (N_29404,N_29332,N_29127);
xor U29405 (N_29405,N_29363,N_29120);
and U29406 (N_29406,N_29209,N_29101);
nor U29407 (N_29407,N_29185,N_29349);
nand U29408 (N_29408,N_29207,N_29264);
xnor U29409 (N_29409,N_29133,N_29257);
and U29410 (N_29410,N_29293,N_29183);
nor U29411 (N_29411,N_29395,N_29102);
nor U29412 (N_29412,N_29153,N_29104);
and U29413 (N_29413,N_29139,N_29201);
nand U29414 (N_29414,N_29382,N_29384);
nand U29415 (N_29415,N_29391,N_29392);
xnor U29416 (N_29416,N_29228,N_29190);
nand U29417 (N_29417,N_29351,N_29358);
or U29418 (N_29418,N_29128,N_29344);
and U29419 (N_29419,N_29371,N_29146);
or U29420 (N_29420,N_29164,N_29166);
xor U29421 (N_29421,N_29191,N_29292);
nand U29422 (N_29422,N_29184,N_29247);
xnor U29423 (N_29423,N_29234,N_29150);
or U29424 (N_29424,N_29277,N_29223);
or U29425 (N_29425,N_29225,N_29126);
xor U29426 (N_29426,N_29140,N_29398);
or U29427 (N_29427,N_29106,N_29307);
or U29428 (N_29428,N_29243,N_29147);
or U29429 (N_29429,N_29206,N_29295);
or U29430 (N_29430,N_29130,N_29350);
nor U29431 (N_29431,N_29238,N_29271);
or U29432 (N_29432,N_29107,N_29124);
nand U29433 (N_29433,N_29219,N_29160);
xor U29434 (N_29434,N_29313,N_29226);
or U29435 (N_29435,N_29370,N_29214);
nor U29436 (N_29436,N_29348,N_29267);
nand U29437 (N_29437,N_29157,N_29205);
and U29438 (N_29438,N_29135,N_29210);
xnor U29439 (N_29439,N_29227,N_29193);
nand U29440 (N_29440,N_29156,N_29389);
and U29441 (N_29441,N_29217,N_29294);
nor U29442 (N_29442,N_29182,N_29303);
nor U29443 (N_29443,N_29194,N_29355);
nor U29444 (N_29444,N_29179,N_29317);
or U29445 (N_29445,N_29119,N_29232);
xnor U29446 (N_29446,N_29244,N_29366);
nand U29447 (N_29447,N_29270,N_29327);
and U29448 (N_29448,N_29187,N_29353);
nor U29449 (N_29449,N_29188,N_29280);
nor U29450 (N_29450,N_29200,N_29168);
xnor U29451 (N_29451,N_29186,N_29380);
or U29452 (N_29452,N_29253,N_29367);
xnor U29453 (N_29453,N_29143,N_29394);
xor U29454 (N_29454,N_29316,N_29386);
xor U29455 (N_29455,N_29290,N_29275);
and U29456 (N_29456,N_29256,N_29278);
xnor U29457 (N_29457,N_29342,N_29302);
and U29458 (N_29458,N_29326,N_29274);
nand U29459 (N_29459,N_29362,N_29279);
nand U29460 (N_29460,N_29357,N_29372);
nor U29461 (N_29461,N_29212,N_29132);
and U29462 (N_29462,N_29324,N_29121);
nand U29463 (N_29463,N_29154,N_29258);
and U29464 (N_29464,N_29231,N_29269);
nor U29465 (N_29465,N_29379,N_29388);
or U29466 (N_29466,N_29165,N_29108);
or U29467 (N_29467,N_29151,N_29211);
nor U29468 (N_29468,N_29268,N_29373);
xor U29469 (N_29469,N_29224,N_29335);
nor U29470 (N_29470,N_29115,N_29393);
xnor U29471 (N_29471,N_29310,N_29235);
nand U29472 (N_29472,N_29272,N_29174);
nor U29473 (N_29473,N_29347,N_29196);
nand U29474 (N_29474,N_29286,N_29298);
nor U29475 (N_29475,N_29237,N_29291);
nand U29476 (N_29476,N_29117,N_29301);
and U29477 (N_29477,N_29105,N_29259);
and U29478 (N_29478,N_29305,N_29399);
or U29479 (N_29479,N_29236,N_29218);
nor U29480 (N_29480,N_29314,N_29176);
nand U29481 (N_29481,N_29137,N_29281);
nor U29482 (N_29482,N_29360,N_29192);
or U29483 (N_29483,N_29375,N_29321);
xnor U29484 (N_29484,N_29131,N_29177);
nor U29485 (N_29485,N_29288,N_29377);
nand U29486 (N_29486,N_29222,N_29100);
nand U29487 (N_29487,N_29262,N_29339);
xor U29488 (N_29488,N_29296,N_29158);
xor U29489 (N_29489,N_29337,N_29122);
xnor U29490 (N_29490,N_29287,N_29263);
xor U29491 (N_29491,N_29376,N_29284);
and U29492 (N_29492,N_29361,N_29343);
and U29493 (N_29493,N_29251,N_29233);
or U29494 (N_29494,N_29246,N_29308);
nor U29495 (N_29495,N_29356,N_29159);
nor U29496 (N_29496,N_29162,N_29276);
nand U29497 (N_29497,N_29285,N_29365);
nand U29498 (N_29498,N_29282,N_29328);
nor U29499 (N_29499,N_29312,N_29374);
or U29500 (N_29500,N_29144,N_29172);
nor U29501 (N_29501,N_29112,N_29230);
or U29502 (N_29502,N_29338,N_29336);
xor U29503 (N_29503,N_29297,N_29173);
nor U29504 (N_29504,N_29323,N_29329);
nor U29505 (N_29505,N_29208,N_29289);
and U29506 (N_29506,N_29180,N_29383);
and U29507 (N_29507,N_29299,N_29204);
nor U29508 (N_29508,N_29249,N_29242);
or U29509 (N_29509,N_29129,N_29368);
nor U29510 (N_29510,N_29141,N_29239);
nand U29511 (N_29511,N_29319,N_29202);
nand U29512 (N_29512,N_29163,N_29250);
and U29513 (N_29513,N_29255,N_29378);
or U29514 (N_29514,N_29306,N_29169);
or U29515 (N_29515,N_29245,N_29300);
nand U29516 (N_29516,N_29346,N_29109);
nor U29517 (N_29517,N_29240,N_29397);
and U29518 (N_29518,N_29142,N_29229);
or U29519 (N_29519,N_29136,N_29145);
nor U29520 (N_29520,N_29216,N_29149);
and U29521 (N_29521,N_29345,N_29283);
or U29522 (N_29522,N_29364,N_29161);
nand U29523 (N_29523,N_29199,N_29125);
and U29524 (N_29524,N_29118,N_29138);
and U29525 (N_29525,N_29390,N_29273);
or U29526 (N_29526,N_29385,N_29134);
or U29527 (N_29527,N_29241,N_29265);
xnor U29528 (N_29528,N_29213,N_29334);
nand U29529 (N_29529,N_29304,N_29266);
nor U29530 (N_29530,N_29260,N_29175);
nand U29531 (N_29531,N_29148,N_29325);
nor U29532 (N_29532,N_29252,N_29359);
or U29533 (N_29533,N_29189,N_29195);
nor U29534 (N_29534,N_29248,N_29340);
nor U29535 (N_29535,N_29198,N_29170);
xnor U29536 (N_29536,N_29220,N_29315);
xnor U29537 (N_29537,N_29221,N_29381);
xor U29538 (N_29538,N_29116,N_29311);
and U29539 (N_29539,N_29387,N_29333);
and U29540 (N_29540,N_29396,N_29254);
xor U29541 (N_29541,N_29197,N_29341);
or U29542 (N_29542,N_29111,N_29155);
and U29543 (N_29543,N_29152,N_29331);
or U29544 (N_29544,N_29261,N_29103);
nor U29545 (N_29545,N_29167,N_29318);
or U29546 (N_29546,N_29110,N_29330);
xor U29547 (N_29547,N_29320,N_29113);
or U29548 (N_29548,N_29369,N_29322);
xnor U29549 (N_29549,N_29114,N_29171);
nor U29550 (N_29550,N_29252,N_29302);
or U29551 (N_29551,N_29139,N_29273);
xor U29552 (N_29552,N_29146,N_29121);
xnor U29553 (N_29553,N_29332,N_29365);
and U29554 (N_29554,N_29157,N_29166);
nand U29555 (N_29555,N_29253,N_29277);
and U29556 (N_29556,N_29354,N_29327);
and U29557 (N_29557,N_29305,N_29392);
nor U29558 (N_29558,N_29377,N_29201);
or U29559 (N_29559,N_29141,N_29380);
nor U29560 (N_29560,N_29209,N_29116);
or U29561 (N_29561,N_29399,N_29134);
nand U29562 (N_29562,N_29276,N_29358);
nand U29563 (N_29563,N_29302,N_29262);
nor U29564 (N_29564,N_29282,N_29224);
xnor U29565 (N_29565,N_29362,N_29323);
nand U29566 (N_29566,N_29100,N_29293);
and U29567 (N_29567,N_29303,N_29212);
or U29568 (N_29568,N_29298,N_29207);
nand U29569 (N_29569,N_29349,N_29298);
or U29570 (N_29570,N_29372,N_29375);
nor U29571 (N_29571,N_29370,N_29393);
nand U29572 (N_29572,N_29380,N_29172);
xor U29573 (N_29573,N_29261,N_29316);
xnor U29574 (N_29574,N_29259,N_29253);
nor U29575 (N_29575,N_29299,N_29365);
and U29576 (N_29576,N_29275,N_29177);
or U29577 (N_29577,N_29140,N_29355);
xor U29578 (N_29578,N_29360,N_29346);
nand U29579 (N_29579,N_29346,N_29238);
nor U29580 (N_29580,N_29181,N_29163);
nand U29581 (N_29581,N_29129,N_29332);
xor U29582 (N_29582,N_29313,N_29376);
and U29583 (N_29583,N_29272,N_29379);
or U29584 (N_29584,N_29314,N_29250);
nand U29585 (N_29585,N_29321,N_29283);
xor U29586 (N_29586,N_29305,N_29180);
xor U29587 (N_29587,N_29210,N_29293);
nand U29588 (N_29588,N_29205,N_29142);
nand U29589 (N_29589,N_29341,N_29379);
nor U29590 (N_29590,N_29274,N_29260);
or U29591 (N_29591,N_29125,N_29138);
and U29592 (N_29592,N_29288,N_29250);
nor U29593 (N_29593,N_29215,N_29164);
xor U29594 (N_29594,N_29351,N_29221);
xnor U29595 (N_29595,N_29302,N_29297);
nand U29596 (N_29596,N_29356,N_29177);
and U29597 (N_29597,N_29343,N_29295);
nand U29598 (N_29598,N_29374,N_29163);
and U29599 (N_29599,N_29387,N_29173);
nand U29600 (N_29600,N_29192,N_29199);
nor U29601 (N_29601,N_29328,N_29240);
xor U29602 (N_29602,N_29353,N_29157);
nand U29603 (N_29603,N_29366,N_29340);
and U29604 (N_29604,N_29177,N_29351);
and U29605 (N_29605,N_29279,N_29370);
or U29606 (N_29606,N_29272,N_29113);
or U29607 (N_29607,N_29212,N_29306);
or U29608 (N_29608,N_29118,N_29286);
xor U29609 (N_29609,N_29155,N_29104);
nand U29610 (N_29610,N_29357,N_29272);
nor U29611 (N_29611,N_29200,N_29234);
and U29612 (N_29612,N_29143,N_29379);
nand U29613 (N_29613,N_29300,N_29142);
or U29614 (N_29614,N_29299,N_29194);
or U29615 (N_29615,N_29260,N_29232);
or U29616 (N_29616,N_29384,N_29391);
and U29617 (N_29617,N_29387,N_29358);
nor U29618 (N_29618,N_29125,N_29362);
or U29619 (N_29619,N_29185,N_29143);
xnor U29620 (N_29620,N_29287,N_29341);
or U29621 (N_29621,N_29131,N_29346);
nand U29622 (N_29622,N_29212,N_29281);
xnor U29623 (N_29623,N_29212,N_29216);
or U29624 (N_29624,N_29157,N_29226);
nand U29625 (N_29625,N_29167,N_29335);
nor U29626 (N_29626,N_29285,N_29369);
xor U29627 (N_29627,N_29138,N_29206);
or U29628 (N_29628,N_29218,N_29233);
xor U29629 (N_29629,N_29350,N_29100);
nand U29630 (N_29630,N_29144,N_29376);
xnor U29631 (N_29631,N_29378,N_29260);
nor U29632 (N_29632,N_29215,N_29162);
and U29633 (N_29633,N_29166,N_29394);
or U29634 (N_29634,N_29104,N_29233);
nor U29635 (N_29635,N_29166,N_29167);
nand U29636 (N_29636,N_29243,N_29311);
nand U29637 (N_29637,N_29205,N_29362);
and U29638 (N_29638,N_29103,N_29399);
and U29639 (N_29639,N_29235,N_29284);
or U29640 (N_29640,N_29303,N_29370);
nand U29641 (N_29641,N_29359,N_29185);
and U29642 (N_29642,N_29109,N_29121);
and U29643 (N_29643,N_29188,N_29149);
xor U29644 (N_29644,N_29269,N_29133);
and U29645 (N_29645,N_29376,N_29201);
nand U29646 (N_29646,N_29359,N_29173);
nand U29647 (N_29647,N_29338,N_29123);
nand U29648 (N_29648,N_29387,N_29296);
or U29649 (N_29649,N_29166,N_29235);
and U29650 (N_29650,N_29131,N_29154);
xnor U29651 (N_29651,N_29321,N_29356);
and U29652 (N_29652,N_29133,N_29146);
nand U29653 (N_29653,N_29382,N_29373);
nor U29654 (N_29654,N_29121,N_29289);
xnor U29655 (N_29655,N_29355,N_29100);
or U29656 (N_29656,N_29109,N_29113);
or U29657 (N_29657,N_29256,N_29358);
nor U29658 (N_29658,N_29305,N_29190);
xnor U29659 (N_29659,N_29289,N_29236);
nand U29660 (N_29660,N_29165,N_29345);
nand U29661 (N_29661,N_29190,N_29235);
or U29662 (N_29662,N_29137,N_29395);
or U29663 (N_29663,N_29183,N_29132);
nand U29664 (N_29664,N_29253,N_29298);
or U29665 (N_29665,N_29249,N_29197);
nor U29666 (N_29666,N_29360,N_29398);
and U29667 (N_29667,N_29235,N_29230);
xor U29668 (N_29668,N_29166,N_29343);
nand U29669 (N_29669,N_29184,N_29392);
nor U29670 (N_29670,N_29275,N_29131);
and U29671 (N_29671,N_29124,N_29225);
xor U29672 (N_29672,N_29248,N_29246);
xor U29673 (N_29673,N_29237,N_29379);
or U29674 (N_29674,N_29116,N_29276);
nand U29675 (N_29675,N_29142,N_29395);
nor U29676 (N_29676,N_29326,N_29350);
nor U29677 (N_29677,N_29193,N_29249);
or U29678 (N_29678,N_29163,N_29170);
and U29679 (N_29679,N_29292,N_29394);
nand U29680 (N_29680,N_29373,N_29353);
nor U29681 (N_29681,N_29147,N_29133);
or U29682 (N_29682,N_29368,N_29235);
and U29683 (N_29683,N_29243,N_29269);
or U29684 (N_29684,N_29324,N_29107);
nor U29685 (N_29685,N_29312,N_29185);
xnor U29686 (N_29686,N_29271,N_29398);
xnor U29687 (N_29687,N_29197,N_29165);
or U29688 (N_29688,N_29192,N_29149);
or U29689 (N_29689,N_29176,N_29389);
and U29690 (N_29690,N_29232,N_29294);
or U29691 (N_29691,N_29101,N_29240);
nor U29692 (N_29692,N_29134,N_29106);
or U29693 (N_29693,N_29387,N_29175);
nand U29694 (N_29694,N_29348,N_29244);
xor U29695 (N_29695,N_29116,N_29200);
or U29696 (N_29696,N_29197,N_29146);
and U29697 (N_29697,N_29284,N_29330);
nor U29698 (N_29698,N_29351,N_29220);
and U29699 (N_29699,N_29156,N_29195);
xor U29700 (N_29700,N_29626,N_29612);
and U29701 (N_29701,N_29415,N_29422);
nor U29702 (N_29702,N_29649,N_29554);
xnor U29703 (N_29703,N_29417,N_29663);
xor U29704 (N_29704,N_29562,N_29569);
and U29705 (N_29705,N_29512,N_29507);
xnor U29706 (N_29706,N_29412,N_29511);
nor U29707 (N_29707,N_29441,N_29584);
and U29708 (N_29708,N_29482,N_29537);
or U29709 (N_29709,N_29401,N_29531);
nor U29710 (N_29710,N_29540,N_29407);
and U29711 (N_29711,N_29628,N_29641);
nor U29712 (N_29712,N_29518,N_29509);
xnor U29713 (N_29713,N_29520,N_29432);
and U29714 (N_29714,N_29669,N_29632);
xor U29715 (N_29715,N_29457,N_29431);
nand U29716 (N_29716,N_29434,N_29436);
or U29717 (N_29717,N_29625,N_29425);
xnor U29718 (N_29718,N_29548,N_29483);
xnor U29719 (N_29719,N_29543,N_29485);
and U29720 (N_29720,N_29501,N_29550);
or U29721 (N_29721,N_29547,N_29451);
nor U29722 (N_29722,N_29521,N_29561);
or U29723 (N_29723,N_29674,N_29536);
xor U29724 (N_29724,N_29418,N_29673);
and U29725 (N_29725,N_29533,N_29629);
nand U29726 (N_29726,N_29532,N_29410);
nor U29727 (N_29727,N_29666,N_29679);
or U29728 (N_29728,N_29620,N_29657);
and U29729 (N_29729,N_29596,N_29583);
or U29730 (N_29730,N_29403,N_29577);
xor U29731 (N_29731,N_29440,N_29650);
xnor U29732 (N_29732,N_29448,N_29559);
xnor U29733 (N_29733,N_29622,N_29426);
nor U29734 (N_29734,N_29645,N_29627);
or U29735 (N_29735,N_29579,N_29530);
or U29736 (N_29736,N_29698,N_29492);
or U29737 (N_29737,N_29670,N_29594);
nand U29738 (N_29738,N_29544,N_29662);
and U29739 (N_29739,N_29607,N_29454);
nor U29740 (N_29740,N_29499,N_29472);
nor U29741 (N_29741,N_29469,N_29664);
nand U29742 (N_29742,N_29637,N_29604);
nor U29743 (N_29743,N_29405,N_29639);
and U29744 (N_29744,N_29439,N_29466);
nand U29745 (N_29745,N_29464,N_29493);
or U29746 (N_29746,N_29661,N_29682);
xor U29747 (N_29747,N_29602,N_29456);
xor U29748 (N_29748,N_29574,N_29567);
or U29749 (N_29749,N_29406,N_29549);
and U29750 (N_29750,N_29692,N_29461);
nand U29751 (N_29751,N_29678,N_29656);
xnor U29752 (N_29752,N_29603,N_29653);
nor U29753 (N_29753,N_29502,N_29582);
and U29754 (N_29754,N_29694,N_29591);
or U29755 (N_29755,N_29595,N_29497);
and U29756 (N_29756,N_29442,N_29508);
or U29757 (N_29757,N_29465,N_29428);
xnor U29758 (N_29758,N_29654,N_29479);
nor U29759 (N_29759,N_29684,N_29546);
xnor U29760 (N_29760,N_29696,N_29560);
nand U29761 (N_29761,N_29635,N_29651);
nand U29762 (N_29762,N_29458,N_29525);
xnor U29763 (N_29763,N_29522,N_29640);
or U29764 (N_29764,N_29646,N_29459);
nor U29765 (N_29765,N_29699,N_29642);
or U29766 (N_29766,N_29437,N_29526);
and U29767 (N_29767,N_29600,N_29402);
and U29768 (N_29768,N_29572,N_29478);
or U29769 (N_29769,N_29668,N_29409);
nor U29770 (N_29770,N_29523,N_29614);
xnor U29771 (N_29771,N_29690,N_29610);
nor U29772 (N_29772,N_29423,N_29414);
xor U29773 (N_29773,N_29506,N_29580);
nor U29774 (N_29774,N_29667,N_29476);
or U29775 (N_29775,N_29613,N_29599);
and U29776 (N_29776,N_29647,N_29494);
xnor U29777 (N_29777,N_29630,N_29480);
xor U29778 (N_29778,N_29558,N_29413);
nor U29779 (N_29779,N_29564,N_29593);
nor U29780 (N_29780,N_29608,N_29644);
or U29781 (N_29781,N_29624,N_29570);
xor U29782 (N_29782,N_29488,N_29615);
xnor U29783 (N_29783,N_29611,N_29513);
xnor U29784 (N_29784,N_29424,N_29467);
nand U29785 (N_29785,N_29433,N_29427);
or U29786 (N_29786,N_29514,N_29455);
nor U29787 (N_29787,N_29585,N_29462);
and U29788 (N_29788,N_29438,N_29566);
nor U29789 (N_29789,N_29598,N_29484);
nand U29790 (N_29790,N_29697,N_29677);
and U29791 (N_29791,N_29689,N_29495);
or U29792 (N_29792,N_29634,N_29631);
nand U29793 (N_29793,N_29589,N_29452);
or U29794 (N_29794,N_29453,N_29486);
and U29795 (N_29795,N_29489,N_29515);
nand U29796 (N_29796,N_29636,N_29571);
and U29797 (N_29797,N_29450,N_29504);
xor U29798 (N_29798,N_29652,N_29538);
and U29799 (N_29799,N_29503,N_29688);
or U29800 (N_29800,N_29576,N_29552);
xor U29801 (N_29801,N_29685,N_29443);
or U29802 (N_29802,N_29643,N_29575);
xor U29803 (N_29803,N_29563,N_29655);
and U29804 (N_29804,N_29539,N_29680);
or U29805 (N_29805,N_29568,N_29545);
and U29806 (N_29806,N_29601,N_29638);
nand U29807 (N_29807,N_29542,N_29471);
xnor U29808 (N_29808,N_29619,N_29421);
and U29809 (N_29809,N_29490,N_29573);
or U29810 (N_29810,N_29460,N_29445);
xor U29811 (N_29811,N_29519,N_29404);
xor U29812 (N_29812,N_29429,N_29605);
nand U29813 (N_29813,N_29618,N_29551);
nor U29814 (N_29814,N_29633,N_29557);
nand U29815 (N_29815,N_29676,N_29474);
xor U29816 (N_29816,N_29535,N_29468);
and U29817 (N_29817,N_29477,N_29505);
xor U29818 (N_29818,N_29616,N_29617);
xnor U29819 (N_29819,N_29516,N_29444);
nand U29820 (N_29820,N_29683,N_29648);
and U29821 (N_29821,N_29587,N_29586);
xnor U29822 (N_29822,N_29491,N_29623);
xnor U29823 (N_29823,N_29411,N_29449);
and U29824 (N_29824,N_29419,N_29681);
xnor U29825 (N_29825,N_29529,N_29496);
and U29826 (N_29826,N_29416,N_29498);
nand U29827 (N_29827,N_29659,N_29510);
nor U29828 (N_29828,N_29555,N_29565);
nor U29829 (N_29829,N_29447,N_29400);
or U29830 (N_29830,N_29556,N_29446);
nor U29831 (N_29831,N_29660,N_29408);
or U29832 (N_29832,N_29470,N_29528);
nand U29833 (N_29833,N_29500,N_29695);
or U29834 (N_29834,N_29473,N_29578);
or U29835 (N_29835,N_29463,N_29606);
nand U29836 (N_29836,N_29691,N_29527);
nor U29837 (N_29837,N_29581,N_29541);
and U29838 (N_29838,N_29430,N_29665);
nor U29839 (N_29839,N_29475,N_29609);
or U29840 (N_29840,N_29592,N_29672);
xor U29841 (N_29841,N_29517,N_29675);
nor U29842 (N_29842,N_29487,N_29693);
nand U29843 (N_29843,N_29590,N_29481);
and U29844 (N_29844,N_29435,N_29686);
nand U29845 (N_29845,N_29597,N_29420);
nor U29846 (N_29846,N_29687,N_29553);
nor U29847 (N_29847,N_29621,N_29534);
xor U29848 (N_29848,N_29658,N_29671);
nand U29849 (N_29849,N_29588,N_29524);
nand U29850 (N_29850,N_29401,N_29681);
nor U29851 (N_29851,N_29413,N_29494);
and U29852 (N_29852,N_29592,N_29477);
or U29853 (N_29853,N_29644,N_29508);
nor U29854 (N_29854,N_29638,N_29449);
nand U29855 (N_29855,N_29627,N_29499);
or U29856 (N_29856,N_29645,N_29414);
or U29857 (N_29857,N_29688,N_29435);
nand U29858 (N_29858,N_29418,N_29479);
and U29859 (N_29859,N_29623,N_29609);
xnor U29860 (N_29860,N_29658,N_29641);
xor U29861 (N_29861,N_29636,N_29624);
nand U29862 (N_29862,N_29618,N_29444);
nor U29863 (N_29863,N_29459,N_29585);
nand U29864 (N_29864,N_29446,N_29505);
nor U29865 (N_29865,N_29416,N_29499);
and U29866 (N_29866,N_29590,N_29535);
or U29867 (N_29867,N_29590,N_29688);
and U29868 (N_29868,N_29455,N_29665);
and U29869 (N_29869,N_29592,N_29435);
nor U29870 (N_29870,N_29443,N_29588);
nor U29871 (N_29871,N_29697,N_29460);
nand U29872 (N_29872,N_29473,N_29566);
xnor U29873 (N_29873,N_29594,N_29625);
and U29874 (N_29874,N_29557,N_29572);
xnor U29875 (N_29875,N_29477,N_29647);
nand U29876 (N_29876,N_29699,N_29485);
xnor U29877 (N_29877,N_29631,N_29637);
or U29878 (N_29878,N_29689,N_29651);
xnor U29879 (N_29879,N_29574,N_29639);
nor U29880 (N_29880,N_29520,N_29461);
xor U29881 (N_29881,N_29500,N_29650);
and U29882 (N_29882,N_29586,N_29477);
and U29883 (N_29883,N_29482,N_29591);
or U29884 (N_29884,N_29639,N_29667);
or U29885 (N_29885,N_29508,N_29621);
nand U29886 (N_29886,N_29652,N_29475);
nand U29887 (N_29887,N_29589,N_29528);
nor U29888 (N_29888,N_29424,N_29617);
xnor U29889 (N_29889,N_29681,N_29572);
xnor U29890 (N_29890,N_29564,N_29425);
and U29891 (N_29891,N_29582,N_29431);
xnor U29892 (N_29892,N_29547,N_29508);
or U29893 (N_29893,N_29447,N_29414);
or U29894 (N_29894,N_29485,N_29685);
and U29895 (N_29895,N_29670,N_29685);
xor U29896 (N_29896,N_29442,N_29668);
nand U29897 (N_29897,N_29592,N_29503);
xnor U29898 (N_29898,N_29466,N_29588);
and U29899 (N_29899,N_29474,N_29487);
and U29900 (N_29900,N_29474,N_29612);
xnor U29901 (N_29901,N_29650,N_29549);
nor U29902 (N_29902,N_29463,N_29563);
nand U29903 (N_29903,N_29525,N_29498);
xor U29904 (N_29904,N_29437,N_29626);
or U29905 (N_29905,N_29416,N_29481);
nand U29906 (N_29906,N_29630,N_29545);
and U29907 (N_29907,N_29669,N_29444);
and U29908 (N_29908,N_29410,N_29548);
or U29909 (N_29909,N_29495,N_29630);
or U29910 (N_29910,N_29551,N_29405);
xor U29911 (N_29911,N_29608,N_29570);
or U29912 (N_29912,N_29643,N_29493);
xor U29913 (N_29913,N_29665,N_29506);
nand U29914 (N_29914,N_29566,N_29569);
xnor U29915 (N_29915,N_29435,N_29629);
nand U29916 (N_29916,N_29571,N_29637);
nand U29917 (N_29917,N_29540,N_29577);
and U29918 (N_29918,N_29410,N_29482);
nor U29919 (N_29919,N_29463,N_29523);
xnor U29920 (N_29920,N_29516,N_29592);
nand U29921 (N_29921,N_29684,N_29570);
nor U29922 (N_29922,N_29548,N_29408);
xor U29923 (N_29923,N_29469,N_29626);
nor U29924 (N_29924,N_29517,N_29539);
or U29925 (N_29925,N_29671,N_29634);
nor U29926 (N_29926,N_29484,N_29463);
or U29927 (N_29927,N_29633,N_29423);
nor U29928 (N_29928,N_29677,N_29580);
nand U29929 (N_29929,N_29465,N_29667);
nand U29930 (N_29930,N_29401,N_29586);
nand U29931 (N_29931,N_29631,N_29675);
or U29932 (N_29932,N_29525,N_29638);
and U29933 (N_29933,N_29468,N_29669);
nor U29934 (N_29934,N_29538,N_29574);
and U29935 (N_29935,N_29626,N_29537);
nor U29936 (N_29936,N_29601,N_29458);
nor U29937 (N_29937,N_29643,N_29602);
or U29938 (N_29938,N_29640,N_29680);
nand U29939 (N_29939,N_29523,N_29618);
and U29940 (N_29940,N_29509,N_29408);
nand U29941 (N_29941,N_29404,N_29545);
nor U29942 (N_29942,N_29444,N_29421);
nor U29943 (N_29943,N_29469,N_29675);
nand U29944 (N_29944,N_29651,N_29678);
and U29945 (N_29945,N_29445,N_29513);
or U29946 (N_29946,N_29473,N_29504);
nor U29947 (N_29947,N_29563,N_29475);
nor U29948 (N_29948,N_29677,N_29624);
nand U29949 (N_29949,N_29652,N_29541);
xor U29950 (N_29950,N_29469,N_29518);
nand U29951 (N_29951,N_29577,N_29625);
or U29952 (N_29952,N_29540,N_29543);
nor U29953 (N_29953,N_29567,N_29499);
nand U29954 (N_29954,N_29442,N_29561);
xnor U29955 (N_29955,N_29685,N_29409);
xnor U29956 (N_29956,N_29593,N_29601);
nor U29957 (N_29957,N_29456,N_29638);
and U29958 (N_29958,N_29625,N_29611);
or U29959 (N_29959,N_29413,N_29411);
nor U29960 (N_29960,N_29668,N_29561);
and U29961 (N_29961,N_29538,N_29677);
and U29962 (N_29962,N_29494,N_29680);
nor U29963 (N_29963,N_29469,N_29555);
and U29964 (N_29964,N_29663,N_29499);
nor U29965 (N_29965,N_29466,N_29534);
nand U29966 (N_29966,N_29695,N_29579);
xnor U29967 (N_29967,N_29475,N_29498);
xor U29968 (N_29968,N_29609,N_29400);
and U29969 (N_29969,N_29509,N_29534);
and U29970 (N_29970,N_29542,N_29526);
nor U29971 (N_29971,N_29614,N_29470);
or U29972 (N_29972,N_29617,N_29458);
nor U29973 (N_29973,N_29507,N_29417);
or U29974 (N_29974,N_29598,N_29485);
and U29975 (N_29975,N_29636,N_29536);
xor U29976 (N_29976,N_29666,N_29627);
xor U29977 (N_29977,N_29502,N_29496);
nor U29978 (N_29978,N_29420,N_29623);
nor U29979 (N_29979,N_29586,N_29673);
nand U29980 (N_29980,N_29523,N_29497);
nor U29981 (N_29981,N_29581,N_29491);
xor U29982 (N_29982,N_29626,N_29610);
nand U29983 (N_29983,N_29623,N_29688);
and U29984 (N_29984,N_29552,N_29561);
nand U29985 (N_29985,N_29599,N_29552);
and U29986 (N_29986,N_29478,N_29625);
xnor U29987 (N_29987,N_29574,N_29648);
nand U29988 (N_29988,N_29617,N_29416);
or U29989 (N_29989,N_29549,N_29640);
nor U29990 (N_29990,N_29671,N_29468);
nand U29991 (N_29991,N_29515,N_29688);
and U29992 (N_29992,N_29542,N_29538);
and U29993 (N_29993,N_29528,N_29515);
nand U29994 (N_29994,N_29602,N_29675);
nor U29995 (N_29995,N_29547,N_29448);
nand U29996 (N_29996,N_29497,N_29645);
xnor U29997 (N_29997,N_29615,N_29657);
and U29998 (N_29998,N_29504,N_29502);
nand U29999 (N_29999,N_29437,N_29645);
xnor UO_0 (O_0,N_29841,N_29908);
nand UO_1 (O_1,N_29753,N_29966);
or UO_2 (O_2,N_29961,N_29938);
or UO_3 (O_3,N_29770,N_29878);
nand UO_4 (O_4,N_29830,N_29703);
or UO_5 (O_5,N_29720,N_29858);
nor UO_6 (O_6,N_29778,N_29754);
or UO_7 (O_7,N_29779,N_29802);
xor UO_8 (O_8,N_29731,N_29928);
and UO_9 (O_9,N_29923,N_29956);
and UO_10 (O_10,N_29847,N_29888);
and UO_11 (O_11,N_29991,N_29814);
and UO_12 (O_12,N_29996,N_29846);
nand UO_13 (O_13,N_29833,N_29740);
xnor UO_14 (O_14,N_29723,N_29829);
nor UO_15 (O_15,N_29792,N_29768);
or UO_16 (O_16,N_29935,N_29948);
nor UO_17 (O_17,N_29977,N_29795);
nor UO_18 (O_18,N_29712,N_29810);
or UO_19 (O_19,N_29735,N_29895);
nand UO_20 (O_20,N_29934,N_29783);
and UO_21 (O_21,N_29827,N_29886);
or UO_22 (O_22,N_29863,N_29749);
nor UO_23 (O_23,N_29907,N_29879);
xor UO_24 (O_24,N_29839,N_29844);
xnor UO_25 (O_25,N_29949,N_29912);
and UO_26 (O_26,N_29872,N_29950);
or UO_27 (O_27,N_29741,N_29889);
nand UO_28 (O_28,N_29999,N_29724);
and UO_29 (O_29,N_29982,N_29881);
and UO_30 (O_30,N_29769,N_29992);
and UO_31 (O_31,N_29732,N_29737);
or UO_32 (O_32,N_29812,N_29859);
and UO_33 (O_33,N_29919,N_29784);
or UO_34 (O_34,N_29856,N_29817);
nor UO_35 (O_35,N_29951,N_29751);
or UO_36 (O_36,N_29954,N_29804);
nor UO_37 (O_37,N_29910,N_29945);
nor UO_38 (O_38,N_29811,N_29920);
nor UO_39 (O_39,N_29882,N_29930);
nor UO_40 (O_40,N_29794,N_29998);
xnor UO_41 (O_41,N_29845,N_29898);
and UO_42 (O_42,N_29709,N_29805);
or UO_43 (O_43,N_29867,N_29765);
or UO_44 (O_44,N_29851,N_29744);
nor UO_45 (O_45,N_29706,N_29815);
nand UO_46 (O_46,N_29902,N_29781);
or UO_47 (O_47,N_29789,N_29931);
nor UO_48 (O_48,N_29868,N_29733);
or UO_49 (O_49,N_29955,N_29965);
or UO_50 (O_50,N_29738,N_29808);
nor UO_51 (O_51,N_29979,N_29860);
or UO_52 (O_52,N_29850,N_29708);
xor UO_53 (O_53,N_29761,N_29947);
and UO_54 (O_54,N_29916,N_29757);
nand UO_55 (O_55,N_29718,N_29836);
nor UO_56 (O_56,N_29911,N_29890);
or UO_57 (O_57,N_29875,N_29906);
and UO_58 (O_58,N_29894,N_29739);
and UO_59 (O_59,N_29989,N_29974);
nand UO_60 (O_60,N_29917,N_29893);
and UO_61 (O_61,N_29866,N_29714);
nand UO_62 (O_62,N_29968,N_29832);
nand UO_63 (O_63,N_29865,N_29818);
or UO_64 (O_64,N_29942,N_29981);
nand UO_65 (O_65,N_29837,N_29800);
xor UO_66 (O_66,N_29984,N_29796);
or UO_67 (O_67,N_29755,N_29892);
nand UO_68 (O_68,N_29760,N_29873);
and UO_69 (O_69,N_29853,N_29854);
xnor UO_70 (O_70,N_29828,N_29978);
and UO_71 (O_71,N_29952,N_29785);
and UO_72 (O_72,N_29904,N_29736);
nor UO_73 (O_73,N_29710,N_29803);
or UO_74 (O_74,N_29793,N_29772);
xor UO_75 (O_75,N_29855,N_29715);
xnor UO_76 (O_76,N_29897,N_29877);
or UO_77 (O_77,N_29964,N_29993);
and UO_78 (O_78,N_29861,N_29849);
and UO_79 (O_79,N_29903,N_29990);
nor UO_80 (O_80,N_29825,N_29870);
or UO_81 (O_81,N_29936,N_29762);
and UO_82 (O_82,N_29728,N_29994);
and UO_83 (O_83,N_29767,N_29746);
nor UO_84 (O_84,N_29913,N_29786);
or UO_85 (O_85,N_29806,N_29899);
xnor UO_86 (O_86,N_29763,N_29730);
or UO_87 (O_87,N_29834,N_29941);
xnor UO_88 (O_88,N_29707,N_29972);
or UO_89 (O_89,N_29750,N_29791);
xor UO_90 (O_90,N_29776,N_29840);
nor UO_91 (O_91,N_29843,N_29716);
nand UO_92 (O_92,N_29986,N_29759);
and UO_93 (O_93,N_29819,N_29967);
xnor UO_94 (O_94,N_29742,N_29876);
and UO_95 (O_95,N_29713,N_29807);
xnor UO_96 (O_96,N_29771,N_29788);
nor UO_97 (O_97,N_29831,N_29922);
nand UO_98 (O_98,N_29959,N_29809);
xnor UO_99 (O_99,N_29727,N_29820);
or UO_100 (O_100,N_29822,N_29957);
nand UO_101 (O_101,N_29905,N_29880);
and UO_102 (O_102,N_29862,N_29777);
and UO_103 (O_103,N_29997,N_29711);
nand UO_104 (O_104,N_29801,N_29702);
nor UO_105 (O_105,N_29824,N_29960);
and UO_106 (O_106,N_29787,N_29756);
xor UO_107 (O_107,N_29891,N_29726);
xor UO_108 (O_108,N_29975,N_29857);
xnor UO_109 (O_109,N_29973,N_29752);
nand UO_110 (O_110,N_29852,N_29764);
nand UO_111 (O_111,N_29940,N_29987);
nand UO_112 (O_112,N_29971,N_29909);
or UO_113 (O_113,N_29918,N_29842);
nor UO_114 (O_114,N_29797,N_29937);
or UO_115 (O_115,N_29932,N_29705);
nand UO_116 (O_116,N_29914,N_29985);
nand UO_117 (O_117,N_29874,N_29864);
nor UO_118 (O_118,N_29915,N_29704);
and UO_119 (O_119,N_29896,N_29953);
nor UO_120 (O_120,N_29798,N_29774);
and UO_121 (O_121,N_29813,N_29983);
xor UO_122 (O_122,N_29962,N_29758);
and UO_123 (O_123,N_29944,N_29969);
nor UO_124 (O_124,N_29943,N_29823);
or UO_125 (O_125,N_29980,N_29885);
nand UO_126 (O_126,N_29725,N_29900);
nor UO_127 (O_127,N_29929,N_29924);
nand UO_128 (O_128,N_29884,N_29729);
or UO_129 (O_129,N_29719,N_29988);
and UO_130 (O_130,N_29835,N_29883);
xor UO_131 (O_131,N_29887,N_29946);
xor UO_132 (O_132,N_29926,N_29976);
or UO_133 (O_133,N_29816,N_29995);
or UO_134 (O_134,N_29826,N_29717);
xor UO_135 (O_135,N_29921,N_29958);
or UO_136 (O_136,N_29734,N_29799);
nor UO_137 (O_137,N_29780,N_29821);
or UO_138 (O_138,N_29838,N_29927);
or UO_139 (O_139,N_29871,N_29963);
nor UO_140 (O_140,N_29848,N_29933);
and UO_141 (O_141,N_29790,N_29747);
or UO_142 (O_142,N_29766,N_29721);
or UO_143 (O_143,N_29745,N_29925);
nand UO_144 (O_144,N_29775,N_29970);
or UO_145 (O_145,N_29743,N_29722);
and UO_146 (O_146,N_29782,N_29773);
or UO_147 (O_147,N_29748,N_29700);
nand UO_148 (O_148,N_29901,N_29701);
nand UO_149 (O_149,N_29939,N_29869);
nand UO_150 (O_150,N_29851,N_29891);
nand UO_151 (O_151,N_29726,N_29873);
and UO_152 (O_152,N_29979,N_29945);
xor UO_153 (O_153,N_29703,N_29758);
nand UO_154 (O_154,N_29815,N_29923);
or UO_155 (O_155,N_29823,N_29803);
and UO_156 (O_156,N_29901,N_29944);
or UO_157 (O_157,N_29774,N_29897);
nor UO_158 (O_158,N_29995,N_29993);
nor UO_159 (O_159,N_29978,N_29795);
nand UO_160 (O_160,N_29938,N_29906);
nand UO_161 (O_161,N_29905,N_29912);
or UO_162 (O_162,N_29901,N_29786);
xor UO_163 (O_163,N_29959,N_29845);
xor UO_164 (O_164,N_29968,N_29955);
nand UO_165 (O_165,N_29997,N_29742);
or UO_166 (O_166,N_29895,N_29933);
nand UO_167 (O_167,N_29722,N_29732);
xor UO_168 (O_168,N_29906,N_29921);
nand UO_169 (O_169,N_29830,N_29988);
and UO_170 (O_170,N_29769,N_29878);
nor UO_171 (O_171,N_29718,N_29740);
and UO_172 (O_172,N_29867,N_29858);
xor UO_173 (O_173,N_29815,N_29902);
xor UO_174 (O_174,N_29964,N_29826);
xor UO_175 (O_175,N_29961,N_29701);
nand UO_176 (O_176,N_29920,N_29855);
and UO_177 (O_177,N_29897,N_29994);
nand UO_178 (O_178,N_29741,N_29818);
nand UO_179 (O_179,N_29824,N_29839);
or UO_180 (O_180,N_29945,N_29767);
xnor UO_181 (O_181,N_29800,N_29702);
or UO_182 (O_182,N_29774,N_29966);
or UO_183 (O_183,N_29840,N_29767);
and UO_184 (O_184,N_29976,N_29817);
nor UO_185 (O_185,N_29846,N_29980);
xor UO_186 (O_186,N_29933,N_29909);
nor UO_187 (O_187,N_29922,N_29842);
or UO_188 (O_188,N_29839,N_29966);
nor UO_189 (O_189,N_29858,N_29875);
nor UO_190 (O_190,N_29767,N_29937);
nor UO_191 (O_191,N_29972,N_29700);
nor UO_192 (O_192,N_29723,N_29909);
xor UO_193 (O_193,N_29787,N_29739);
xnor UO_194 (O_194,N_29760,N_29882);
or UO_195 (O_195,N_29959,N_29795);
nand UO_196 (O_196,N_29822,N_29794);
or UO_197 (O_197,N_29709,N_29907);
xnor UO_198 (O_198,N_29964,N_29724);
and UO_199 (O_199,N_29925,N_29835);
nor UO_200 (O_200,N_29893,N_29873);
nand UO_201 (O_201,N_29941,N_29870);
nand UO_202 (O_202,N_29726,N_29984);
xor UO_203 (O_203,N_29893,N_29702);
and UO_204 (O_204,N_29781,N_29870);
or UO_205 (O_205,N_29877,N_29717);
and UO_206 (O_206,N_29899,N_29874);
and UO_207 (O_207,N_29941,N_29758);
or UO_208 (O_208,N_29783,N_29864);
and UO_209 (O_209,N_29909,N_29883);
and UO_210 (O_210,N_29998,N_29891);
xnor UO_211 (O_211,N_29943,N_29912);
nor UO_212 (O_212,N_29801,N_29846);
nand UO_213 (O_213,N_29716,N_29926);
xnor UO_214 (O_214,N_29933,N_29986);
and UO_215 (O_215,N_29914,N_29982);
and UO_216 (O_216,N_29784,N_29790);
or UO_217 (O_217,N_29729,N_29775);
nand UO_218 (O_218,N_29971,N_29826);
xor UO_219 (O_219,N_29720,N_29721);
xnor UO_220 (O_220,N_29760,N_29719);
or UO_221 (O_221,N_29700,N_29869);
and UO_222 (O_222,N_29871,N_29879);
nor UO_223 (O_223,N_29895,N_29806);
nor UO_224 (O_224,N_29744,N_29919);
nand UO_225 (O_225,N_29714,N_29846);
nor UO_226 (O_226,N_29907,N_29755);
and UO_227 (O_227,N_29734,N_29821);
nand UO_228 (O_228,N_29980,N_29721);
or UO_229 (O_229,N_29754,N_29868);
xnor UO_230 (O_230,N_29994,N_29773);
nor UO_231 (O_231,N_29957,N_29730);
xor UO_232 (O_232,N_29834,N_29991);
and UO_233 (O_233,N_29784,N_29730);
or UO_234 (O_234,N_29991,N_29867);
nand UO_235 (O_235,N_29805,N_29755);
xor UO_236 (O_236,N_29722,N_29817);
or UO_237 (O_237,N_29936,N_29925);
xnor UO_238 (O_238,N_29983,N_29985);
or UO_239 (O_239,N_29910,N_29803);
or UO_240 (O_240,N_29709,N_29833);
xnor UO_241 (O_241,N_29912,N_29751);
nand UO_242 (O_242,N_29718,N_29896);
and UO_243 (O_243,N_29991,N_29947);
nand UO_244 (O_244,N_29957,N_29991);
xor UO_245 (O_245,N_29975,N_29745);
nor UO_246 (O_246,N_29884,N_29798);
and UO_247 (O_247,N_29853,N_29771);
or UO_248 (O_248,N_29953,N_29844);
or UO_249 (O_249,N_29750,N_29974);
or UO_250 (O_250,N_29891,N_29811);
xnor UO_251 (O_251,N_29970,N_29749);
nand UO_252 (O_252,N_29920,N_29712);
or UO_253 (O_253,N_29757,N_29793);
nor UO_254 (O_254,N_29753,N_29981);
nor UO_255 (O_255,N_29704,N_29797);
or UO_256 (O_256,N_29814,N_29977);
nor UO_257 (O_257,N_29874,N_29835);
nand UO_258 (O_258,N_29971,N_29783);
or UO_259 (O_259,N_29755,N_29717);
or UO_260 (O_260,N_29722,N_29868);
xnor UO_261 (O_261,N_29998,N_29952);
nand UO_262 (O_262,N_29722,N_29816);
nor UO_263 (O_263,N_29881,N_29816);
nor UO_264 (O_264,N_29831,N_29797);
nor UO_265 (O_265,N_29855,N_29736);
nor UO_266 (O_266,N_29857,N_29756);
or UO_267 (O_267,N_29727,N_29845);
nand UO_268 (O_268,N_29905,N_29853);
nand UO_269 (O_269,N_29827,N_29872);
and UO_270 (O_270,N_29927,N_29721);
or UO_271 (O_271,N_29805,N_29990);
nand UO_272 (O_272,N_29875,N_29862);
xnor UO_273 (O_273,N_29954,N_29889);
and UO_274 (O_274,N_29851,N_29887);
or UO_275 (O_275,N_29889,N_29760);
xnor UO_276 (O_276,N_29893,N_29863);
nand UO_277 (O_277,N_29969,N_29897);
nor UO_278 (O_278,N_29877,N_29752);
and UO_279 (O_279,N_29959,N_29987);
nand UO_280 (O_280,N_29853,N_29909);
nor UO_281 (O_281,N_29995,N_29818);
and UO_282 (O_282,N_29980,N_29922);
nand UO_283 (O_283,N_29794,N_29956);
nor UO_284 (O_284,N_29817,N_29797);
nand UO_285 (O_285,N_29951,N_29964);
xor UO_286 (O_286,N_29812,N_29772);
and UO_287 (O_287,N_29701,N_29917);
xnor UO_288 (O_288,N_29743,N_29766);
or UO_289 (O_289,N_29775,N_29733);
nor UO_290 (O_290,N_29984,N_29771);
nand UO_291 (O_291,N_29780,N_29810);
nand UO_292 (O_292,N_29754,N_29802);
or UO_293 (O_293,N_29969,N_29721);
nor UO_294 (O_294,N_29941,N_29958);
nand UO_295 (O_295,N_29974,N_29715);
xor UO_296 (O_296,N_29942,N_29777);
xor UO_297 (O_297,N_29981,N_29941);
and UO_298 (O_298,N_29875,N_29733);
xnor UO_299 (O_299,N_29836,N_29828);
nand UO_300 (O_300,N_29979,N_29717);
nor UO_301 (O_301,N_29712,N_29776);
and UO_302 (O_302,N_29899,N_29830);
nand UO_303 (O_303,N_29865,N_29963);
nand UO_304 (O_304,N_29800,N_29731);
nor UO_305 (O_305,N_29766,N_29891);
or UO_306 (O_306,N_29716,N_29914);
nor UO_307 (O_307,N_29829,N_29901);
or UO_308 (O_308,N_29712,N_29848);
nand UO_309 (O_309,N_29934,N_29911);
or UO_310 (O_310,N_29703,N_29899);
nor UO_311 (O_311,N_29709,N_29950);
and UO_312 (O_312,N_29880,N_29902);
and UO_313 (O_313,N_29736,N_29846);
and UO_314 (O_314,N_29705,N_29966);
nor UO_315 (O_315,N_29948,N_29713);
xor UO_316 (O_316,N_29955,N_29739);
or UO_317 (O_317,N_29758,N_29920);
and UO_318 (O_318,N_29882,N_29778);
and UO_319 (O_319,N_29992,N_29740);
xor UO_320 (O_320,N_29925,N_29779);
or UO_321 (O_321,N_29889,N_29822);
nand UO_322 (O_322,N_29779,N_29719);
nand UO_323 (O_323,N_29828,N_29763);
xor UO_324 (O_324,N_29878,N_29887);
nand UO_325 (O_325,N_29719,N_29932);
or UO_326 (O_326,N_29973,N_29816);
nand UO_327 (O_327,N_29891,N_29777);
or UO_328 (O_328,N_29870,N_29908);
and UO_329 (O_329,N_29929,N_29979);
and UO_330 (O_330,N_29751,N_29879);
nand UO_331 (O_331,N_29825,N_29897);
nor UO_332 (O_332,N_29974,N_29992);
and UO_333 (O_333,N_29941,N_29980);
nor UO_334 (O_334,N_29778,N_29909);
xor UO_335 (O_335,N_29719,N_29814);
and UO_336 (O_336,N_29875,N_29857);
nand UO_337 (O_337,N_29890,N_29800);
xnor UO_338 (O_338,N_29763,N_29903);
and UO_339 (O_339,N_29701,N_29739);
nor UO_340 (O_340,N_29742,N_29814);
and UO_341 (O_341,N_29976,N_29776);
and UO_342 (O_342,N_29970,N_29913);
nor UO_343 (O_343,N_29778,N_29735);
xnor UO_344 (O_344,N_29878,N_29833);
nor UO_345 (O_345,N_29783,N_29963);
nor UO_346 (O_346,N_29952,N_29822);
or UO_347 (O_347,N_29764,N_29973);
and UO_348 (O_348,N_29728,N_29714);
and UO_349 (O_349,N_29764,N_29811);
xor UO_350 (O_350,N_29748,N_29792);
nand UO_351 (O_351,N_29899,N_29817);
or UO_352 (O_352,N_29721,N_29763);
and UO_353 (O_353,N_29832,N_29702);
nand UO_354 (O_354,N_29975,N_29898);
and UO_355 (O_355,N_29803,N_29807);
nand UO_356 (O_356,N_29709,N_29937);
nor UO_357 (O_357,N_29944,N_29961);
nor UO_358 (O_358,N_29756,N_29777);
and UO_359 (O_359,N_29874,N_29951);
xnor UO_360 (O_360,N_29859,N_29912);
xor UO_361 (O_361,N_29832,N_29899);
and UO_362 (O_362,N_29992,N_29994);
or UO_363 (O_363,N_29961,N_29893);
nand UO_364 (O_364,N_29835,N_29934);
xor UO_365 (O_365,N_29741,N_29863);
or UO_366 (O_366,N_29717,N_29914);
or UO_367 (O_367,N_29901,N_29703);
nand UO_368 (O_368,N_29781,N_29959);
nand UO_369 (O_369,N_29794,N_29994);
xor UO_370 (O_370,N_29968,N_29842);
nor UO_371 (O_371,N_29853,N_29813);
nor UO_372 (O_372,N_29897,N_29918);
and UO_373 (O_373,N_29887,N_29719);
or UO_374 (O_374,N_29771,N_29837);
nor UO_375 (O_375,N_29850,N_29743);
xnor UO_376 (O_376,N_29872,N_29796);
xor UO_377 (O_377,N_29760,N_29738);
nor UO_378 (O_378,N_29793,N_29752);
xor UO_379 (O_379,N_29814,N_29755);
nand UO_380 (O_380,N_29708,N_29909);
and UO_381 (O_381,N_29721,N_29897);
nor UO_382 (O_382,N_29715,N_29749);
xor UO_383 (O_383,N_29882,N_29707);
nor UO_384 (O_384,N_29832,N_29864);
nor UO_385 (O_385,N_29714,N_29903);
nand UO_386 (O_386,N_29759,N_29954);
or UO_387 (O_387,N_29827,N_29857);
or UO_388 (O_388,N_29714,N_29865);
xor UO_389 (O_389,N_29918,N_29883);
or UO_390 (O_390,N_29748,N_29921);
nor UO_391 (O_391,N_29708,N_29931);
nand UO_392 (O_392,N_29878,N_29860);
and UO_393 (O_393,N_29757,N_29926);
nor UO_394 (O_394,N_29916,N_29947);
and UO_395 (O_395,N_29782,N_29957);
nor UO_396 (O_396,N_29922,N_29890);
nand UO_397 (O_397,N_29931,N_29979);
nand UO_398 (O_398,N_29980,N_29905);
nor UO_399 (O_399,N_29887,N_29853);
and UO_400 (O_400,N_29925,N_29723);
nand UO_401 (O_401,N_29729,N_29969);
and UO_402 (O_402,N_29728,N_29809);
and UO_403 (O_403,N_29777,N_29878);
xnor UO_404 (O_404,N_29954,N_29776);
nand UO_405 (O_405,N_29935,N_29799);
and UO_406 (O_406,N_29846,N_29706);
or UO_407 (O_407,N_29796,N_29910);
nand UO_408 (O_408,N_29971,N_29803);
or UO_409 (O_409,N_29827,N_29890);
xor UO_410 (O_410,N_29733,N_29985);
nor UO_411 (O_411,N_29938,N_29713);
and UO_412 (O_412,N_29984,N_29980);
nand UO_413 (O_413,N_29783,N_29838);
nor UO_414 (O_414,N_29755,N_29995);
xor UO_415 (O_415,N_29903,N_29974);
and UO_416 (O_416,N_29944,N_29993);
xor UO_417 (O_417,N_29866,N_29912);
xor UO_418 (O_418,N_29810,N_29716);
or UO_419 (O_419,N_29704,N_29897);
nor UO_420 (O_420,N_29880,N_29862);
xor UO_421 (O_421,N_29956,N_29889);
and UO_422 (O_422,N_29843,N_29760);
nor UO_423 (O_423,N_29795,N_29971);
and UO_424 (O_424,N_29719,N_29905);
or UO_425 (O_425,N_29878,N_29830);
and UO_426 (O_426,N_29772,N_29895);
and UO_427 (O_427,N_29869,N_29767);
xor UO_428 (O_428,N_29857,N_29984);
or UO_429 (O_429,N_29777,N_29723);
and UO_430 (O_430,N_29739,N_29989);
nand UO_431 (O_431,N_29846,N_29830);
and UO_432 (O_432,N_29778,N_29947);
and UO_433 (O_433,N_29745,N_29826);
nor UO_434 (O_434,N_29726,N_29772);
or UO_435 (O_435,N_29825,N_29815);
nand UO_436 (O_436,N_29790,N_29738);
xnor UO_437 (O_437,N_29805,N_29792);
nand UO_438 (O_438,N_29763,N_29731);
or UO_439 (O_439,N_29864,N_29819);
nand UO_440 (O_440,N_29761,N_29940);
xor UO_441 (O_441,N_29760,N_29769);
nand UO_442 (O_442,N_29757,N_29937);
or UO_443 (O_443,N_29857,N_29949);
and UO_444 (O_444,N_29716,N_29940);
nor UO_445 (O_445,N_29865,N_29706);
nor UO_446 (O_446,N_29928,N_29983);
xnor UO_447 (O_447,N_29802,N_29993);
or UO_448 (O_448,N_29958,N_29777);
nand UO_449 (O_449,N_29907,N_29925);
or UO_450 (O_450,N_29958,N_29710);
xor UO_451 (O_451,N_29833,N_29970);
or UO_452 (O_452,N_29905,N_29865);
nand UO_453 (O_453,N_29742,N_29816);
nor UO_454 (O_454,N_29742,N_29965);
or UO_455 (O_455,N_29981,N_29845);
and UO_456 (O_456,N_29812,N_29952);
nor UO_457 (O_457,N_29767,N_29791);
or UO_458 (O_458,N_29788,N_29838);
nand UO_459 (O_459,N_29891,N_29978);
nor UO_460 (O_460,N_29798,N_29720);
or UO_461 (O_461,N_29788,N_29893);
and UO_462 (O_462,N_29980,N_29767);
and UO_463 (O_463,N_29878,N_29976);
and UO_464 (O_464,N_29880,N_29712);
nand UO_465 (O_465,N_29785,N_29745);
or UO_466 (O_466,N_29849,N_29727);
nand UO_467 (O_467,N_29774,N_29859);
or UO_468 (O_468,N_29946,N_29733);
nand UO_469 (O_469,N_29876,N_29936);
nand UO_470 (O_470,N_29808,N_29807);
and UO_471 (O_471,N_29849,N_29722);
and UO_472 (O_472,N_29992,N_29901);
or UO_473 (O_473,N_29977,N_29730);
nand UO_474 (O_474,N_29964,N_29753);
and UO_475 (O_475,N_29751,N_29913);
or UO_476 (O_476,N_29810,N_29853);
xnor UO_477 (O_477,N_29825,N_29826);
nor UO_478 (O_478,N_29875,N_29736);
xor UO_479 (O_479,N_29963,N_29756);
xnor UO_480 (O_480,N_29930,N_29807);
or UO_481 (O_481,N_29799,N_29854);
nor UO_482 (O_482,N_29729,N_29754);
and UO_483 (O_483,N_29718,N_29834);
and UO_484 (O_484,N_29855,N_29894);
or UO_485 (O_485,N_29864,N_29872);
and UO_486 (O_486,N_29706,N_29918);
or UO_487 (O_487,N_29716,N_29702);
or UO_488 (O_488,N_29966,N_29819);
nor UO_489 (O_489,N_29944,N_29952);
xor UO_490 (O_490,N_29725,N_29850);
xnor UO_491 (O_491,N_29758,N_29828);
nand UO_492 (O_492,N_29810,N_29992);
nor UO_493 (O_493,N_29911,N_29927);
and UO_494 (O_494,N_29933,N_29748);
nor UO_495 (O_495,N_29872,N_29924);
or UO_496 (O_496,N_29866,N_29792);
xor UO_497 (O_497,N_29754,N_29926);
and UO_498 (O_498,N_29800,N_29861);
nand UO_499 (O_499,N_29856,N_29950);
and UO_500 (O_500,N_29820,N_29743);
nand UO_501 (O_501,N_29915,N_29943);
or UO_502 (O_502,N_29779,N_29750);
nor UO_503 (O_503,N_29780,N_29777);
nand UO_504 (O_504,N_29776,N_29933);
nand UO_505 (O_505,N_29758,N_29810);
nand UO_506 (O_506,N_29882,N_29774);
nand UO_507 (O_507,N_29800,N_29822);
nand UO_508 (O_508,N_29774,N_29772);
and UO_509 (O_509,N_29919,N_29880);
and UO_510 (O_510,N_29711,N_29937);
and UO_511 (O_511,N_29934,N_29817);
and UO_512 (O_512,N_29793,N_29843);
or UO_513 (O_513,N_29827,N_29922);
xor UO_514 (O_514,N_29914,N_29979);
or UO_515 (O_515,N_29838,N_29971);
or UO_516 (O_516,N_29987,N_29881);
xnor UO_517 (O_517,N_29756,N_29931);
and UO_518 (O_518,N_29870,N_29714);
nand UO_519 (O_519,N_29733,N_29898);
xor UO_520 (O_520,N_29749,N_29957);
and UO_521 (O_521,N_29929,N_29746);
xor UO_522 (O_522,N_29847,N_29983);
or UO_523 (O_523,N_29999,N_29741);
xnor UO_524 (O_524,N_29881,N_29849);
xor UO_525 (O_525,N_29910,N_29791);
and UO_526 (O_526,N_29916,N_29945);
or UO_527 (O_527,N_29748,N_29898);
and UO_528 (O_528,N_29917,N_29874);
nand UO_529 (O_529,N_29896,N_29708);
xnor UO_530 (O_530,N_29705,N_29840);
or UO_531 (O_531,N_29931,N_29753);
xor UO_532 (O_532,N_29828,N_29782);
xor UO_533 (O_533,N_29744,N_29925);
and UO_534 (O_534,N_29747,N_29849);
or UO_535 (O_535,N_29907,N_29913);
or UO_536 (O_536,N_29816,N_29906);
or UO_537 (O_537,N_29969,N_29825);
xor UO_538 (O_538,N_29826,N_29830);
xor UO_539 (O_539,N_29975,N_29936);
xnor UO_540 (O_540,N_29716,N_29723);
and UO_541 (O_541,N_29854,N_29840);
nand UO_542 (O_542,N_29805,N_29726);
nand UO_543 (O_543,N_29919,N_29955);
nand UO_544 (O_544,N_29736,N_29983);
and UO_545 (O_545,N_29873,N_29812);
xnor UO_546 (O_546,N_29845,N_29833);
nor UO_547 (O_547,N_29804,N_29816);
nor UO_548 (O_548,N_29974,N_29853);
and UO_549 (O_549,N_29870,N_29752);
nand UO_550 (O_550,N_29950,N_29711);
and UO_551 (O_551,N_29775,N_29744);
and UO_552 (O_552,N_29750,N_29894);
or UO_553 (O_553,N_29787,N_29855);
xor UO_554 (O_554,N_29735,N_29898);
nor UO_555 (O_555,N_29914,N_29813);
nor UO_556 (O_556,N_29970,N_29843);
nand UO_557 (O_557,N_29925,N_29834);
and UO_558 (O_558,N_29909,N_29988);
or UO_559 (O_559,N_29822,N_29977);
nand UO_560 (O_560,N_29848,N_29990);
xnor UO_561 (O_561,N_29778,N_29868);
or UO_562 (O_562,N_29852,N_29791);
or UO_563 (O_563,N_29998,N_29923);
nor UO_564 (O_564,N_29908,N_29876);
nand UO_565 (O_565,N_29991,N_29922);
xnor UO_566 (O_566,N_29864,N_29716);
or UO_567 (O_567,N_29957,N_29884);
nor UO_568 (O_568,N_29750,N_29846);
and UO_569 (O_569,N_29834,N_29968);
and UO_570 (O_570,N_29907,N_29769);
nor UO_571 (O_571,N_29886,N_29822);
nor UO_572 (O_572,N_29789,N_29987);
nand UO_573 (O_573,N_29845,N_29892);
nor UO_574 (O_574,N_29963,N_29910);
nor UO_575 (O_575,N_29934,N_29703);
nand UO_576 (O_576,N_29713,N_29736);
nor UO_577 (O_577,N_29977,N_29933);
or UO_578 (O_578,N_29915,N_29826);
xor UO_579 (O_579,N_29866,N_29939);
and UO_580 (O_580,N_29920,N_29818);
nand UO_581 (O_581,N_29977,N_29739);
or UO_582 (O_582,N_29981,N_29905);
and UO_583 (O_583,N_29923,N_29708);
and UO_584 (O_584,N_29809,N_29960);
nand UO_585 (O_585,N_29948,N_29879);
nand UO_586 (O_586,N_29958,N_29902);
and UO_587 (O_587,N_29894,N_29926);
xor UO_588 (O_588,N_29835,N_29869);
or UO_589 (O_589,N_29939,N_29980);
or UO_590 (O_590,N_29760,N_29962);
xor UO_591 (O_591,N_29756,N_29876);
nor UO_592 (O_592,N_29762,N_29779);
xor UO_593 (O_593,N_29826,N_29945);
xor UO_594 (O_594,N_29950,N_29788);
xnor UO_595 (O_595,N_29701,N_29948);
or UO_596 (O_596,N_29945,N_29822);
or UO_597 (O_597,N_29897,N_29812);
nand UO_598 (O_598,N_29838,N_29816);
and UO_599 (O_599,N_29806,N_29873);
nor UO_600 (O_600,N_29937,N_29803);
nor UO_601 (O_601,N_29718,N_29843);
or UO_602 (O_602,N_29827,N_29797);
xor UO_603 (O_603,N_29777,N_29872);
nor UO_604 (O_604,N_29722,N_29794);
and UO_605 (O_605,N_29956,N_29780);
or UO_606 (O_606,N_29964,N_29747);
xor UO_607 (O_607,N_29847,N_29927);
xor UO_608 (O_608,N_29880,N_29770);
and UO_609 (O_609,N_29859,N_29836);
nand UO_610 (O_610,N_29747,N_29910);
and UO_611 (O_611,N_29803,N_29911);
nand UO_612 (O_612,N_29958,N_29810);
and UO_613 (O_613,N_29871,N_29796);
nor UO_614 (O_614,N_29952,N_29882);
or UO_615 (O_615,N_29782,N_29701);
nand UO_616 (O_616,N_29741,N_29859);
xor UO_617 (O_617,N_29718,N_29859);
and UO_618 (O_618,N_29815,N_29992);
nand UO_619 (O_619,N_29897,N_29839);
xor UO_620 (O_620,N_29942,N_29976);
nor UO_621 (O_621,N_29793,N_29981);
and UO_622 (O_622,N_29801,N_29749);
nand UO_623 (O_623,N_29833,N_29803);
nand UO_624 (O_624,N_29860,N_29754);
and UO_625 (O_625,N_29833,N_29828);
nor UO_626 (O_626,N_29761,N_29822);
xnor UO_627 (O_627,N_29927,N_29906);
and UO_628 (O_628,N_29894,N_29781);
and UO_629 (O_629,N_29968,N_29782);
or UO_630 (O_630,N_29889,N_29748);
xor UO_631 (O_631,N_29823,N_29804);
nor UO_632 (O_632,N_29774,N_29858);
and UO_633 (O_633,N_29719,N_29912);
nand UO_634 (O_634,N_29869,N_29866);
and UO_635 (O_635,N_29711,N_29808);
or UO_636 (O_636,N_29846,N_29785);
and UO_637 (O_637,N_29811,N_29744);
nor UO_638 (O_638,N_29913,N_29995);
nor UO_639 (O_639,N_29714,N_29898);
and UO_640 (O_640,N_29708,N_29953);
and UO_641 (O_641,N_29839,N_29710);
and UO_642 (O_642,N_29791,N_29872);
and UO_643 (O_643,N_29952,N_29927);
nand UO_644 (O_644,N_29743,N_29969);
and UO_645 (O_645,N_29791,N_29930);
nor UO_646 (O_646,N_29733,N_29740);
and UO_647 (O_647,N_29794,N_29865);
nor UO_648 (O_648,N_29848,N_29961);
and UO_649 (O_649,N_29903,N_29950);
and UO_650 (O_650,N_29767,N_29881);
and UO_651 (O_651,N_29786,N_29941);
xor UO_652 (O_652,N_29864,N_29859);
and UO_653 (O_653,N_29867,N_29711);
xor UO_654 (O_654,N_29766,N_29926);
or UO_655 (O_655,N_29736,N_29850);
and UO_656 (O_656,N_29704,N_29907);
nor UO_657 (O_657,N_29818,N_29721);
nand UO_658 (O_658,N_29996,N_29930);
and UO_659 (O_659,N_29965,N_29985);
or UO_660 (O_660,N_29951,N_29807);
xor UO_661 (O_661,N_29868,N_29893);
xnor UO_662 (O_662,N_29937,N_29726);
nor UO_663 (O_663,N_29732,N_29969);
xor UO_664 (O_664,N_29849,N_29930);
xor UO_665 (O_665,N_29761,N_29756);
nand UO_666 (O_666,N_29870,N_29902);
xnor UO_667 (O_667,N_29971,N_29988);
and UO_668 (O_668,N_29824,N_29882);
or UO_669 (O_669,N_29715,N_29987);
or UO_670 (O_670,N_29944,N_29741);
nor UO_671 (O_671,N_29726,N_29980);
and UO_672 (O_672,N_29804,N_29980);
nand UO_673 (O_673,N_29742,N_29760);
nand UO_674 (O_674,N_29816,N_29771);
nor UO_675 (O_675,N_29814,N_29999);
nand UO_676 (O_676,N_29747,N_29760);
nor UO_677 (O_677,N_29813,N_29863);
xnor UO_678 (O_678,N_29791,N_29900);
nand UO_679 (O_679,N_29950,N_29920);
xnor UO_680 (O_680,N_29763,N_29726);
nor UO_681 (O_681,N_29843,N_29860);
or UO_682 (O_682,N_29835,N_29781);
or UO_683 (O_683,N_29835,N_29794);
nand UO_684 (O_684,N_29930,N_29971);
xor UO_685 (O_685,N_29874,N_29763);
or UO_686 (O_686,N_29932,N_29842);
or UO_687 (O_687,N_29790,N_29843);
or UO_688 (O_688,N_29781,N_29860);
xnor UO_689 (O_689,N_29808,N_29974);
and UO_690 (O_690,N_29823,N_29882);
nand UO_691 (O_691,N_29736,N_29782);
or UO_692 (O_692,N_29932,N_29788);
xnor UO_693 (O_693,N_29894,N_29963);
nor UO_694 (O_694,N_29880,N_29960);
nand UO_695 (O_695,N_29925,N_29716);
xnor UO_696 (O_696,N_29847,N_29887);
and UO_697 (O_697,N_29765,N_29842);
nor UO_698 (O_698,N_29823,N_29840);
nor UO_699 (O_699,N_29806,N_29760);
nand UO_700 (O_700,N_29716,N_29889);
or UO_701 (O_701,N_29866,N_29950);
xnor UO_702 (O_702,N_29738,N_29963);
nor UO_703 (O_703,N_29772,N_29722);
and UO_704 (O_704,N_29751,N_29761);
nand UO_705 (O_705,N_29714,N_29880);
and UO_706 (O_706,N_29808,N_29716);
nor UO_707 (O_707,N_29891,N_29840);
xor UO_708 (O_708,N_29790,N_29959);
xor UO_709 (O_709,N_29956,N_29932);
or UO_710 (O_710,N_29797,N_29796);
xor UO_711 (O_711,N_29728,N_29774);
nor UO_712 (O_712,N_29815,N_29986);
nand UO_713 (O_713,N_29705,N_29743);
nand UO_714 (O_714,N_29854,N_29972);
and UO_715 (O_715,N_29794,N_29748);
or UO_716 (O_716,N_29955,N_29905);
and UO_717 (O_717,N_29817,N_29801);
nand UO_718 (O_718,N_29902,N_29968);
nand UO_719 (O_719,N_29908,N_29820);
nand UO_720 (O_720,N_29854,N_29887);
nor UO_721 (O_721,N_29895,N_29718);
or UO_722 (O_722,N_29861,N_29785);
xnor UO_723 (O_723,N_29847,N_29753);
nand UO_724 (O_724,N_29839,N_29904);
and UO_725 (O_725,N_29709,N_29863);
nor UO_726 (O_726,N_29960,N_29747);
nor UO_727 (O_727,N_29991,N_29835);
or UO_728 (O_728,N_29702,N_29973);
nor UO_729 (O_729,N_29938,N_29923);
nor UO_730 (O_730,N_29844,N_29837);
and UO_731 (O_731,N_29992,N_29703);
xnor UO_732 (O_732,N_29861,N_29822);
nand UO_733 (O_733,N_29848,N_29971);
or UO_734 (O_734,N_29989,N_29704);
and UO_735 (O_735,N_29995,N_29732);
and UO_736 (O_736,N_29740,N_29995);
or UO_737 (O_737,N_29951,N_29995);
and UO_738 (O_738,N_29982,N_29780);
and UO_739 (O_739,N_29883,N_29855);
xnor UO_740 (O_740,N_29834,N_29721);
nand UO_741 (O_741,N_29791,N_29831);
xnor UO_742 (O_742,N_29729,N_29862);
nor UO_743 (O_743,N_29873,N_29795);
xor UO_744 (O_744,N_29999,N_29922);
and UO_745 (O_745,N_29889,N_29773);
nand UO_746 (O_746,N_29845,N_29876);
xnor UO_747 (O_747,N_29735,N_29844);
xnor UO_748 (O_748,N_29723,N_29845);
nor UO_749 (O_749,N_29714,N_29774);
nor UO_750 (O_750,N_29988,N_29737);
or UO_751 (O_751,N_29704,N_29967);
nand UO_752 (O_752,N_29950,N_29978);
nor UO_753 (O_753,N_29972,N_29904);
nand UO_754 (O_754,N_29802,N_29922);
and UO_755 (O_755,N_29800,N_29886);
nor UO_756 (O_756,N_29863,N_29800);
xor UO_757 (O_757,N_29780,N_29830);
xnor UO_758 (O_758,N_29841,N_29810);
nand UO_759 (O_759,N_29796,N_29869);
xor UO_760 (O_760,N_29988,N_29755);
and UO_761 (O_761,N_29834,N_29711);
nor UO_762 (O_762,N_29803,N_29718);
or UO_763 (O_763,N_29743,N_29802);
and UO_764 (O_764,N_29841,N_29876);
nor UO_765 (O_765,N_29959,N_29832);
nand UO_766 (O_766,N_29802,N_29958);
nand UO_767 (O_767,N_29801,N_29962);
and UO_768 (O_768,N_29896,N_29863);
xnor UO_769 (O_769,N_29847,N_29879);
and UO_770 (O_770,N_29846,N_29712);
nand UO_771 (O_771,N_29735,N_29814);
or UO_772 (O_772,N_29828,N_29872);
xnor UO_773 (O_773,N_29820,N_29868);
nand UO_774 (O_774,N_29806,N_29809);
xor UO_775 (O_775,N_29704,N_29796);
xor UO_776 (O_776,N_29808,N_29844);
and UO_777 (O_777,N_29902,N_29959);
nor UO_778 (O_778,N_29958,N_29957);
nor UO_779 (O_779,N_29949,N_29813);
xor UO_780 (O_780,N_29756,N_29863);
nor UO_781 (O_781,N_29987,N_29742);
nand UO_782 (O_782,N_29970,N_29825);
or UO_783 (O_783,N_29964,N_29782);
or UO_784 (O_784,N_29827,N_29998);
and UO_785 (O_785,N_29909,N_29942);
nand UO_786 (O_786,N_29754,N_29703);
or UO_787 (O_787,N_29910,N_29877);
and UO_788 (O_788,N_29881,N_29862);
nor UO_789 (O_789,N_29854,N_29893);
nor UO_790 (O_790,N_29744,N_29876);
nor UO_791 (O_791,N_29756,N_29708);
and UO_792 (O_792,N_29957,N_29952);
and UO_793 (O_793,N_29761,N_29842);
nor UO_794 (O_794,N_29986,N_29923);
or UO_795 (O_795,N_29776,N_29838);
nor UO_796 (O_796,N_29858,N_29852);
xnor UO_797 (O_797,N_29879,N_29829);
or UO_798 (O_798,N_29970,N_29751);
nor UO_799 (O_799,N_29844,N_29820);
and UO_800 (O_800,N_29984,N_29869);
or UO_801 (O_801,N_29774,N_29969);
nand UO_802 (O_802,N_29774,N_29990);
and UO_803 (O_803,N_29765,N_29939);
nand UO_804 (O_804,N_29762,N_29826);
nor UO_805 (O_805,N_29863,N_29978);
nor UO_806 (O_806,N_29850,N_29702);
nand UO_807 (O_807,N_29892,N_29883);
xor UO_808 (O_808,N_29973,N_29868);
nand UO_809 (O_809,N_29804,N_29734);
nand UO_810 (O_810,N_29717,N_29863);
xor UO_811 (O_811,N_29779,N_29946);
xor UO_812 (O_812,N_29969,N_29987);
nor UO_813 (O_813,N_29977,N_29708);
nor UO_814 (O_814,N_29795,N_29906);
and UO_815 (O_815,N_29881,N_29774);
or UO_816 (O_816,N_29778,N_29918);
xor UO_817 (O_817,N_29722,N_29809);
nor UO_818 (O_818,N_29995,N_29811);
and UO_819 (O_819,N_29990,N_29851);
and UO_820 (O_820,N_29915,N_29797);
or UO_821 (O_821,N_29888,N_29940);
nand UO_822 (O_822,N_29892,N_29903);
or UO_823 (O_823,N_29700,N_29717);
or UO_824 (O_824,N_29873,N_29904);
xnor UO_825 (O_825,N_29867,N_29732);
and UO_826 (O_826,N_29889,N_29909);
nand UO_827 (O_827,N_29817,N_29994);
nand UO_828 (O_828,N_29707,N_29907);
nor UO_829 (O_829,N_29954,N_29743);
and UO_830 (O_830,N_29799,N_29700);
or UO_831 (O_831,N_29995,N_29793);
nand UO_832 (O_832,N_29714,N_29700);
nand UO_833 (O_833,N_29916,N_29937);
or UO_834 (O_834,N_29985,N_29966);
or UO_835 (O_835,N_29752,N_29900);
nand UO_836 (O_836,N_29929,N_29898);
nand UO_837 (O_837,N_29825,N_29849);
and UO_838 (O_838,N_29726,N_29876);
xnor UO_839 (O_839,N_29860,N_29726);
xor UO_840 (O_840,N_29895,N_29782);
nor UO_841 (O_841,N_29856,N_29975);
nand UO_842 (O_842,N_29708,N_29700);
xnor UO_843 (O_843,N_29761,N_29959);
nor UO_844 (O_844,N_29848,N_29745);
nor UO_845 (O_845,N_29761,N_29891);
nor UO_846 (O_846,N_29755,N_29775);
nand UO_847 (O_847,N_29865,N_29877);
nand UO_848 (O_848,N_29857,N_29780);
nor UO_849 (O_849,N_29828,N_29912);
and UO_850 (O_850,N_29783,N_29853);
nor UO_851 (O_851,N_29774,N_29997);
nor UO_852 (O_852,N_29964,N_29769);
nor UO_853 (O_853,N_29936,N_29894);
and UO_854 (O_854,N_29857,N_29701);
nor UO_855 (O_855,N_29822,N_29762);
or UO_856 (O_856,N_29799,N_29970);
nor UO_857 (O_857,N_29716,N_29985);
or UO_858 (O_858,N_29895,N_29785);
xnor UO_859 (O_859,N_29930,N_29726);
or UO_860 (O_860,N_29823,N_29716);
nor UO_861 (O_861,N_29906,N_29736);
nand UO_862 (O_862,N_29860,N_29819);
nand UO_863 (O_863,N_29746,N_29957);
nor UO_864 (O_864,N_29974,N_29987);
or UO_865 (O_865,N_29875,N_29824);
nor UO_866 (O_866,N_29732,N_29794);
nand UO_867 (O_867,N_29997,N_29948);
or UO_868 (O_868,N_29750,N_29834);
or UO_869 (O_869,N_29885,N_29936);
or UO_870 (O_870,N_29845,N_29900);
xnor UO_871 (O_871,N_29997,N_29951);
nor UO_872 (O_872,N_29821,N_29779);
and UO_873 (O_873,N_29721,N_29967);
nor UO_874 (O_874,N_29755,N_29769);
xnor UO_875 (O_875,N_29921,N_29788);
nor UO_876 (O_876,N_29753,N_29787);
nor UO_877 (O_877,N_29885,N_29749);
nand UO_878 (O_878,N_29970,N_29941);
nor UO_879 (O_879,N_29848,N_29760);
nor UO_880 (O_880,N_29703,N_29791);
nor UO_881 (O_881,N_29732,N_29977);
nand UO_882 (O_882,N_29873,N_29723);
nand UO_883 (O_883,N_29907,N_29874);
and UO_884 (O_884,N_29791,N_29746);
nor UO_885 (O_885,N_29945,N_29914);
nor UO_886 (O_886,N_29883,N_29977);
nor UO_887 (O_887,N_29965,N_29878);
or UO_888 (O_888,N_29939,N_29948);
nor UO_889 (O_889,N_29741,N_29796);
nand UO_890 (O_890,N_29845,N_29852);
xnor UO_891 (O_891,N_29923,N_29787);
nor UO_892 (O_892,N_29779,N_29927);
xor UO_893 (O_893,N_29987,N_29862);
nand UO_894 (O_894,N_29937,N_29894);
nor UO_895 (O_895,N_29966,N_29934);
nand UO_896 (O_896,N_29742,N_29933);
or UO_897 (O_897,N_29894,N_29764);
nor UO_898 (O_898,N_29707,N_29927);
xor UO_899 (O_899,N_29933,N_29887);
and UO_900 (O_900,N_29994,N_29813);
nand UO_901 (O_901,N_29864,N_29898);
nor UO_902 (O_902,N_29712,N_29789);
nor UO_903 (O_903,N_29704,N_29763);
nor UO_904 (O_904,N_29944,N_29866);
or UO_905 (O_905,N_29743,N_29893);
nand UO_906 (O_906,N_29945,N_29941);
xor UO_907 (O_907,N_29868,N_29721);
nor UO_908 (O_908,N_29771,N_29735);
and UO_909 (O_909,N_29949,N_29791);
or UO_910 (O_910,N_29758,N_29829);
and UO_911 (O_911,N_29745,N_29916);
or UO_912 (O_912,N_29832,N_29922);
nor UO_913 (O_913,N_29973,N_29782);
nand UO_914 (O_914,N_29741,N_29960);
nor UO_915 (O_915,N_29754,N_29893);
and UO_916 (O_916,N_29971,N_29953);
or UO_917 (O_917,N_29995,N_29795);
or UO_918 (O_918,N_29892,N_29738);
nor UO_919 (O_919,N_29767,N_29972);
nor UO_920 (O_920,N_29841,N_29923);
nor UO_921 (O_921,N_29835,N_29734);
xor UO_922 (O_922,N_29758,N_29739);
nor UO_923 (O_923,N_29794,N_29805);
and UO_924 (O_924,N_29876,N_29725);
or UO_925 (O_925,N_29753,N_29938);
and UO_926 (O_926,N_29708,N_29863);
nand UO_927 (O_927,N_29833,N_29863);
and UO_928 (O_928,N_29883,N_29820);
xnor UO_929 (O_929,N_29740,N_29779);
nor UO_930 (O_930,N_29879,N_29910);
nor UO_931 (O_931,N_29825,N_29876);
and UO_932 (O_932,N_29761,N_29845);
xnor UO_933 (O_933,N_29859,N_29944);
xor UO_934 (O_934,N_29768,N_29733);
nor UO_935 (O_935,N_29828,N_29901);
nor UO_936 (O_936,N_29993,N_29911);
xor UO_937 (O_937,N_29902,N_29775);
xnor UO_938 (O_938,N_29733,N_29848);
and UO_939 (O_939,N_29760,N_29995);
xnor UO_940 (O_940,N_29804,N_29948);
and UO_941 (O_941,N_29722,N_29956);
and UO_942 (O_942,N_29979,N_29773);
nor UO_943 (O_943,N_29892,N_29747);
nand UO_944 (O_944,N_29971,N_29976);
or UO_945 (O_945,N_29723,N_29878);
or UO_946 (O_946,N_29782,N_29868);
and UO_947 (O_947,N_29705,N_29829);
or UO_948 (O_948,N_29832,N_29861);
and UO_949 (O_949,N_29913,N_29958);
nor UO_950 (O_950,N_29741,N_29931);
and UO_951 (O_951,N_29728,N_29761);
nor UO_952 (O_952,N_29772,N_29948);
or UO_953 (O_953,N_29736,N_29809);
nor UO_954 (O_954,N_29758,N_29892);
nor UO_955 (O_955,N_29920,N_29913);
or UO_956 (O_956,N_29832,N_29888);
or UO_957 (O_957,N_29983,N_29712);
xnor UO_958 (O_958,N_29822,N_29789);
xor UO_959 (O_959,N_29948,N_29899);
and UO_960 (O_960,N_29935,N_29976);
or UO_961 (O_961,N_29720,N_29818);
xnor UO_962 (O_962,N_29936,N_29884);
nor UO_963 (O_963,N_29837,N_29952);
xor UO_964 (O_964,N_29976,N_29718);
or UO_965 (O_965,N_29974,N_29884);
and UO_966 (O_966,N_29918,N_29960);
or UO_967 (O_967,N_29872,N_29829);
xnor UO_968 (O_968,N_29868,N_29740);
and UO_969 (O_969,N_29735,N_29943);
nand UO_970 (O_970,N_29785,N_29722);
xnor UO_971 (O_971,N_29853,N_29939);
xnor UO_972 (O_972,N_29904,N_29815);
xnor UO_973 (O_973,N_29900,N_29905);
or UO_974 (O_974,N_29841,N_29772);
xnor UO_975 (O_975,N_29899,N_29828);
xnor UO_976 (O_976,N_29738,N_29964);
xnor UO_977 (O_977,N_29923,N_29718);
nand UO_978 (O_978,N_29804,N_29744);
or UO_979 (O_979,N_29705,N_29965);
nor UO_980 (O_980,N_29835,N_29995);
or UO_981 (O_981,N_29843,N_29822);
or UO_982 (O_982,N_29856,N_29864);
and UO_983 (O_983,N_29831,N_29873);
nand UO_984 (O_984,N_29899,N_29743);
xnor UO_985 (O_985,N_29844,N_29772);
xor UO_986 (O_986,N_29789,N_29811);
nor UO_987 (O_987,N_29726,N_29817);
nand UO_988 (O_988,N_29786,N_29973);
nand UO_989 (O_989,N_29896,N_29957);
nand UO_990 (O_990,N_29835,N_29913);
nor UO_991 (O_991,N_29756,N_29856);
nand UO_992 (O_992,N_29752,N_29736);
nor UO_993 (O_993,N_29752,N_29943);
xnor UO_994 (O_994,N_29978,N_29700);
nor UO_995 (O_995,N_29772,N_29947);
and UO_996 (O_996,N_29810,N_29733);
nand UO_997 (O_997,N_29717,N_29767);
xor UO_998 (O_998,N_29708,N_29984);
and UO_999 (O_999,N_29845,N_29922);
nand UO_1000 (O_1000,N_29958,N_29837);
nor UO_1001 (O_1001,N_29850,N_29885);
nand UO_1002 (O_1002,N_29993,N_29752);
nor UO_1003 (O_1003,N_29961,N_29746);
nand UO_1004 (O_1004,N_29718,N_29951);
nor UO_1005 (O_1005,N_29912,N_29973);
nand UO_1006 (O_1006,N_29903,N_29912);
xnor UO_1007 (O_1007,N_29905,N_29898);
or UO_1008 (O_1008,N_29880,N_29997);
nand UO_1009 (O_1009,N_29788,N_29915);
nand UO_1010 (O_1010,N_29789,N_29904);
or UO_1011 (O_1011,N_29736,N_29723);
xor UO_1012 (O_1012,N_29899,N_29873);
nor UO_1013 (O_1013,N_29932,N_29938);
nand UO_1014 (O_1014,N_29773,N_29839);
or UO_1015 (O_1015,N_29791,N_29970);
and UO_1016 (O_1016,N_29915,N_29755);
or UO_1017 (O_1017,N_29995,N_29805);
xnor UO_1018 (O_1018,N_29777,N_29832);
and UO_1019 (O_1019,N_29954,N_29837);
and UO_1020 (O_1020,N_29914,N_29852);
nand UO_1021 (O_1021,N_29938,N_29774);
xor UO_1022 (O_1022,N_29976,N_29822);
xnor UO_1023 (O_1023,N_29912,N_29716);
and UO_1024 (O_1024,N_29760,N_29922);
xnor UO_1025 (O_1025,N_29923,N_29884);
or UO_1026 (O_1026,N_29914,N_29935);
nor UO_1027 (O_1027,N_29790,N_29992);
nor UO_1028 (O_1028,N_29996,N_29723);
and UO_1029 (O_1029,N_29786,N_29967);
and UO_1030 (O_1030,N_29721,N_29800);
xnor UO_1031 (O_1031,N_29874,N_29993);
and UO_1032 (O_1032,N_29965,N_29903);
nand UO_1033 (O_1033,N_29814,N_29852);
xor UO_1034 (O_1034,N_29975,N_29893);
nor UO_1035 (O_1035,N_29777,N_29805);
nor UO_1036 (O_1036,N_29757,N_29724);
or UO_1037 (O_1037,N_29800,N_29959);
xor UO_1038 (O_1038,N_29860,N_29926);
and UO_1039 (O_1039,N_29950,N_29955);
or UO_1040 (O_1040,N_29871,N_29894);
nand UO_1041 (O_1041,N_29723,N_29769);
or UO_1042 (O_1042,N_29897,N_29962);
xor UO_1043 (O_1043,N_29791,N_29773);
and UO_1044 (O_1044,N_29932,N_29704);
or UO_1045 (O_1045,N_29726,N_29958);
nand UO_1046 (O_1046,N_29756,N_29972);
xnor UO_1047 (O_1047,N_29961,N_29707);
and UO_1048 (O_1048,N_29937,N_29881);
xnor UO_1049 (O_1049,N_29728,N_29837);
nand UO_1050 (O_1050,N_29725,N_29940);
nor UO_1051 (O_1051,N_29751,N_29853);
xnor UO_1052 (O_1052,N_29984,N_29908);
or UO_1053 (O_1053,N_29926,N_29993);
nand UO_1054 (O_1054,N_29980,N_29966);
nand UO_1055 (O_1055,N_29783,N_29960);
nand UO_1056 (O_1056,N_29912,N_29784);
and UO_1057 (O_1057,N_29965,N_29733);
nor UO_1058 (O_1058,N_29779,N_29911);
nand UO_1059 (O_1059,N_29966,N_29943);
or UO_1060 (O_1060,N_29951,N_29864);
nand UO_1061 (O_1061,N_29814,N_29976);
nand UO_1062 (O_1062,N_29862,N_29980);
nor UO_1063 (O_1063,N_29898,N_29944);
nor UO_1064 (O_1064,N_29709,N_29728);
nand UO_1065 (O_1065,N_29825,N_29796);
xnor UO_1066 (O_1066,N_29863,N_29938);
and UO_1067 (O_1067,N_29846,N_29967);
nand UO_1068 (O_1068,N_29727,N_29885);
or UO_1069 (O_1069,N_29788,N_29734);
xor UO_1070 (O_1070,N_29927,N_29830);
nor UO_1071 (O_1071,N_29969,N_29807);
nand UO_1072 (O_1072,N_29855,N_29785);
and UO_1073 (O_1073,N_29729,N_29903);
nor UO_1074 (O_1074,N_29785,N_29807);
or UO_1075 (O_1075,N_29771,N_29854);
xnor UO_1076 (O_1076,N_29716,N_29719);
or UO_1077 (O_1077,N_29705,N_29993);
xnor UO_1078 (O_1078,N_29886,N_29854);
nor UO_1079 (O_1079,N_29974,N_29905);
or UO_1080 (O_1080,N_29748,N_29934);
nor UO_1081 (O_1081,N_29772,N_29751);
nor UO_1082 (O_1082,N_29984,N_29919);
xnor UO_1083 (O_1083,N_29862,N_29811);
xor UO_1084 (O_1084,N_29783,N_29904);
or UO_1085 (O_1085,N_29894,N_29730);
nor UO_1086 (O_1086,N_29716,N_29870);
and UO_1087 (O_1087,N_29709,N_29806);
and UO_1088 (O_1088,N_29883,N_29839);
xor UO_1089 (O_1089,N_29944,N_29869);
xor UO_1090 (O_1090,N_29994,N_29875);
or UO_1091 (O_1091,N_29806,N_29891);
and UO_1092 (O_1092,N_29901,N_29888);
and UO_1093 (O_1093,N_29795,N_29877);
xor UO_1094 (O_1094,N_29789,N_29738);
xor UO_1095 (O_1095,N_29718,N_29986);
and UO_1096 (O_1096,N_29949,N_29864);
nor UO_1097 (O_1097,N_29711,N_29804);
xnor UO_1098 (O_1098,N_29882,N_29736);
and UO_1099 (O_1099,N_29935,N_29845);
nor UO_1100 (O_1100,N_29747,N_29721);
and UO_1101 (O_1101,N_29894,N_29841);
or UO_1102 (O_1102,N_29918,N_29914);
nor UO_1103 (O_1103,N_29754,N_29743);
nand UO_1104 (O_1104,N_29868,N_29862);
xnor UO_1105 (O_1105,N_29967,N_29831);
nand UO_1106 (O_1106,N_29967,N_29785);
nand UO_1107 (O_1107,N_29800,N_29793);
nor UO_1108 (O_1108,N_29705,N_29976);
xor UO_1109 (O_1109,N_29828,N_29997);
or UO_1110 (O_1110,N_29999,N_29849);
nand UO_1111 (O_1111,N_29834,N_29935);
or UO_1112 (O_1112,N_29967,N_29944);
nor UO_1113 (O_1113,N_29754,N_29747);
nand UO_1114 (O_1114,N_29864,N_29910);
nand UO_1115 (O_1115,N_29798,N_29748);
and UO_1116 (O_1116,N_29706,N_29920);
nand UO_1117 (O_1117,N_29704,N_29961);
nand UO_1118 (O_1118,N_29766,N_29816);
nand UO_1119 (O_1119,N_29913,N_29766);
nand UO_1120 (O_1120,N_29814,N_29776);
xnor UO_1121 (O_1121,N_29949,N_29919);
nor UO_1122 (O_1122,N_29914,N_29943);
xor UO_1123 (O_1123,N_29855,N_29822);
or UO_1124 (O_1124,N_29966,N_29910);
and UO_1125 (O_1125,N_29858,N_29816);
and UO_1126 (O_1126,N_29838,N_29749);
and UO_1127 (O_1127,N_29968,N_29733);
and UO_1128 (O_1128,N_29946,N_29755);
nor UO_1129 (O_1129,N_29760,N_29856);
or UO_1130 (O_1130,N_29887,N_29899);
nor UO_1131 (O_1131,N_29861,N_29856);
and UO_1132 (O_1132,N_29872,N_29903);
or UO_1133 (O_1133,N_29850,N_29813);
nand UO_1134 (O_1134,N_29763,N_29896);
nand UO_1135 (O_1135,N_29947,N_29862);
or UO_1136 (O_1136,N_29927,N_29741);
and UO_1137 (O_1137,N_29902,N_29744);
xor UO_1138 (O_1138,N_29755,N_29780);
and UO_1139 (O_1139,N_29892,N_29846);
and UO_1140 (O_1140,N_29742,N_29963);
or UO_1141 (O_1141,N_29773,N_29894);
or UO_1142 (O_1142,N_29773,N_29840);
or UO_1143 (O_1143,N_29782,N_29799);
and UO_1144 (O_1144,N_29776,N_29918);
or UO_1145 (O_1145,N_29970,N_29741);
or UO_1146 (O_1146,N_29819,N_29916);
and UO_1147 (O_1147,N_29804,N_29894);
or UO_1148 (O_1148,N_29793,N_29810);
or UO_1149 (O_1149,N_29852,N_29752);
nor UO_1150 (O_1150,N_29833,N_29926);
or UO_1151 (O_1151,N_29996,N_29909);
xor UO_1152 (O_1152,N_29880,N_29800);
or UO_1153 (O_1153,N_29712,N_29832);
or UO_1154 (O_1154,N_29766,N_29894);
nand UO_1155 (O_1155,N_29879,N_29839);
or UO_1156 (O_1156,N_29833,N_29887);
or UO_1157 (O_1157,N_29728,N_29888);
or UO_1158 (O_1158,N_29917,N_29835);
xnor UO_1159 (O_1159,N_29740,N_29987);
nor UO_1160 (O_1160,N_29982,N_29734);
and UO_1161 (O_1161,N_29976,N_29830);
nand UO_1162 (O_1162,N_29849,N_29779);
or UO_1163 (O_1163,N_29791,N_29856);
or UO_1164 (O_1164,N_29942,N_29905);
nand UO_1165 (O_1165,N_29967,N_29927);
xor UO_1166 (O_1166,N_29897,N_29944);
or UO_1167 (O_1167,N_29788,N_29807);
nand UO_1168 (O_1168,N_29891,N_29966);
xor UO_1169 (O_1169,N_29911,N_29881);
xor UO_1170 (O_1170,N_29742,N_29991);
or UO_1171 (O_1171,N_29992,N_29878);
or UO_1172 (O_1172,N_29917,N_29952);
nand UO_1173 (O_1173,N_29948,N_29783);
nor UO_1174 (O_1174,N_29883,N_29997);
nor UO_1175 (O_1175,N_29831,N_29766);
nand UO_1176 (O_1176,N_29746,N_29958);
nor UO_1177 (O_1177,N_29893,N_29978);
nor UO_1178 (O_1178,N_29840,N_29730);
nand UO_1179 (O_1179,N_29713,N_29937);
nor UO_1180 (O_1180,N_29783,N_29987);
or UO_1181 (O_1181,N_29871,N_29946);
nor UO_1182 (O_1182,N_29749,N_29830);
nand UO_1183 (O_1183,N_29782,N_29844);
and UO_1184 (O_1184,N_29736,N_29956);
and UO_1185 (O_1185,N_29821,N_29924);
or UO_1186 (O_1186,N_29734,N_29747);
and UO_1187 (O_1187,N_29800,N_29954);
nand UO_1188 (O_1188,N_29975,N_29853);
or UO_1189 (O_1189,N_29916,N_29717);
and UO_1190 (O_1190,N_29719,N_29888);
nor UO_1191 (O_1191,N_29900,N_29772);
or UO_1192 (O_1192,N_29861,N_29776);
nor UO_1193 (O_1193,N_29937,N_29931);
nor UO_1194 (O_1194,N_29862,N_29840);
nand UO_1195 (O_1195,N_29957,N_29837);
xnor UO_1196 (O_1196,N_29774,N_29760);
nand UO_1197 (O_1197,N_29857,N_29957);
xnor UO_1198 (O_1198,N_29946,N_29943);
nand UO_1199 (O_1199,N_29870,N_29985);
nor UO_1200 (O_1200,N_29906,N_29738);
nand UO_1201 (O_1201,N_29886,N_29944);
xor UO_1202 (O_1202,N_29929,N_29770);
or UO_1203 (O_1203,N_29984,N_29752);
and UO_1204 (O_1204,N_29889,N_29807);
xor UO_1205 (O_1205,N_29807,N_29753);
and UO_1206 (O_1206,N_29941,N_29954);
or UO_1207 (O_1207,N_29925,N_29732);
nand UO_1208 (O_1208,N_29786,N_29887);
xnor UO_1209 (O_1209,N_29944,N_29724);
nand UO_1210 (O_1210,N_29958,N_29806);
or UO_1211 (O_1211,N_29924,N_29811);
and UO_1212 (O_1212,N_29897,N_29756);
nand UO_1213 (O_1213,N_29864,N_29913);
nor UO_1214 (O_1214,N_29895,N_29960);
nor UO_1215 (O_1215,N_29921,N_29772);
or UO_1216 (O_1216,N_29901,N_29999);
or UO_1217 (O_1217,N_29944,N_29973);
and UO_1218 (O_1218,N_29912,N_29837);
xnor UO_1219 (O_1219,N_29992,N_29889);
and UO_1220 (O_1220,N_29936,N_29758);
or UO_1221 (O_1221,N_29843,N_29879);
nand UO_1222 (O_1222,N_29926,N_29964);
or UO_1223 (O_1223,N_29934,N_29985);
and UO_1224 (O_1224,N_29942,N_29756);
xor UO_1225 (O_1225,N_29811,N_29893);
nand UO_1226 (O_1226,N_29765,N_29717);
and UO_1227 (O_1227,N_29957,N_29783);
xnor UO_1228 (O_1228,N_29937,N_29766);
nand UO_1229 (O_1229,N_29777,N_29846);
nand UO_1230 (O_1230,N_29933,N_29914);
nand UO_1231 (O_1231,N_29977,N_29748);
nand UO_1232 (O_1232,N_29721,N_29869);
and UO_1233 (O_1233,N_29928,N_29926);
xnor UO_1234 (O_1234,N_29924,N_29940);
xnor UO_1235 (O_1235,N_29730,N_29923);
nor UO_1236 (O_1236,N_29991,N_29897);
or UO_1237 (O_1237,N_29788,N_29985);
or UO_1238 (O_1238,N_29755,N_29831);
or UO_1239 (O_1239,N_29806,N_29706);
nor UO_1240 (O_1240,N_29856,N_29829);
xnor UO_1241 (O_1241,N_29749,N_29790);
nand UO_1242 (O_1242,N_29928,N_29751);
nor UO_1243 (O_1243,N_29941,N_29778);
or UO_1244 (O_1244,N_29798,N_29846);
or UO_1245 (O_1245,N_29930,N_29754);
nand UO_1246 (O_1246,N_29965,N_29729);
nor UO_1247 (O_1247,N_29974,N_29796);
nor UO_1248 (O_1248,N_29764,N_29837);
and UO_1249 (O_1249,N_29824,N_29747);
or UO_1250 (O_1250,N_29777,N_29860);
nand UO_1251 (O_1251,N_29715,N_29780);
xnor UO_1252 (O_1252,N_29867,N_29918);
or UO_1253 (O_1253,N_29967,N_29941);
or UO_1254 (O_1254,N_29814,N_29788);
nor UO_1255 (O_1255,N_29738,N_29894);
or UO_1256 (O_1256,N_29738,N_29811);
nor UO_1257 (O_1257,N_29869,N_29948);
nand UO_1258 (O_1258,N_29906,N_29799);
nor UO_1259 (O_1259,N_29772,N_29857);
or UO_1260 (O_1260,N_29966,N_29965);
nand UO_1261 (O_1261,N_29996,N_29709);
nand UO_1262 (O_1262,N_29840,N_29886);
nand UO_1263 (O_1263,N_29791,N_29923);
nor UO_1264 (O_1264,N_29787,N_29911);
nand UO_1265 (O_1265,N_29892,N_29704);
and UO_1266 (O_1266,N_29800,N_29770);
nand UO_1267 (O_1267,N_29773,N_29712);
nor UO_1268 (O_1268,N_29714,N_29778);
xnor UO_1269 (O_1269,N_29898,N_29749);
nor UO_1270 (O_1270,N_29744,N_29749);
xnor UO_1271 (O_1271,N_29916,N_29843);
xnor UO_1272 (O_1272,N_29884,N_29955);
nor UO_1273 (O_1273,N_29917,N_29842);
or UO_1274 (O_1274,N_29722,N_29759);
or UO_1275 (O_1275,N_29775,N_29741);
and UO_1276 (O_1276,N_29737,N_29731);
and UO_1277 (O_1277,N_29799,N_29844);
nor UO_1278 (O_1278,N_29984,N_29700);
nand UO_1279 (O_1279,N_29933,N_29924);
nor UO_1280 (O_1280,N_29858,N_29920);
or UO_1281 (O_1281,N_29966,N_29745);
and UO_1282 (O_1282,N_29825,N_29728);
nor UO_1283 (O_1283,N_29778,N_29803);
nor UO_1284 (O_1284,N_29823,N_29895);
and UO_1285 (O_1285,N_29759,N_29823);
or UO_1286 (O_1286,N_29702,N_29927);
and UO_1287 (O_1287,N_29987,N_29772);
and UO_1288 (O_1288,N_29848,N_29947);
nand UO_1289 (O_1289,N_29751,N_29856);
nor UO_1290 (O_1290,N_29718,N_29906);
nor UO_1291 (O_1291,N_29944,N_29707);
xor UO_1292 (O_1292,N_29891,N_29983);
and UO_1293 (O_1293,N_29874,N_29756);
nand UO_1294 (O_1294,N_29755,N_29936);
xor UO_1295 (O_1295,N_29920,N_29719);
or UO_1296 (O_1296,N_29803,N_29935);
nor UO_1297 (O_1297,N_29828,N_29711);
nor UO_1298 (O_1298,N_29960,N_29707);
or UO_1299 (O_1299,N_29810,N_29864);
nand UO_1300 (O_1300,N_29796,N_29967);
xnor UO_1301 (O_1301,N_29861,N_29712);
or UO_1302 (O_1302,N_29843,N_29730);
and UO_1303 (O_1303,N_29792,N_29951);
xnor UO_1304 (O_1304,N_29994,N_29715);
or UO_1305 (O_1305,N_29909,N_29767);
and UO_1306 (O_1306,N_29725,N_29703);
or UO_1307 (O_1307,N_29927,N_29816);
or UO_1308 (O_1308,N_29928,N_29816);
or UO_1309 (O_1309,N_29874,N_29748);
and UO_1310 (O_1310,N_29866,N_29943);
and UO_1311 (O_1311,N_29796,N_29978);
nand UO_1312 (O_1312,N_29831,N_29896);
nand UO_1313 (O_1313,N_29930,N_29766);
xor UO_1314 (O_1314,N_29895,N_29889);
nor UO_1315 (O_1315,N_29762,N_29792);
and UO_1316 (O_1316,N_29824,N_29725);
and UO_1317 (O_1317,N_29820,N_29976);
or UO_1318 (O_1318,N_29860,N_29906);
nor UO_1319 (O_1319,N_29892,N_29991);
or UO_1320 (O_1320,N_29799,N_29867);
or UO_1321 (O_1321,N_29890,N_29718);
nand UO_1322 (O_1322,N_29928,N_29872);
nand UO_1323 (O_1323,N_29765,N_29959);
nor UO_1324 (O_1324,N_29961,N_29831);
nand UO_1325 (O_1325,N_29795,N_29917);
xor UO_1326 (O_1326,N_29881,N_29773);
xor UO_1327 (O_1327,N_29792,N_29874);
and UO_1328 (O_1328,N_29770,N_29885);
xnor UO_1329 (O_1329,N_29985,N_29993);
or UO_1330 (O_1330,N_29782,N_29745);
nor UO_1331 (O_1331,N_29813,N_29962);
nand UO_1332 (O_1332,N_29894,N_29971);
nand UO_1333 (O_1333,N_29727,N_29776);
or UO_1334 (O_1334,N_29945,N_29709);
xor UO_1335 (O_1335,N_29748,N_29908);
nor UO_1336 (O_1336,N_29767,N_29971);
xor UO_1337 (O_1337,N_29904,N_29963);
nor UO_1338 (O_1338,N_29936,N_29931);
or UO_1339 (O_1339,N_29757,N_29990);
nor UO_1340 (O_1340,N_29763,N_29920);
or UO_1341 (O_1341,N_29748,N_29931);
or UO_1342 (O_1342,N_29754,N_29855);
xor UO_1343 (O_1343,N_29869,N_29832);
xor UO_1344 (O_1344,N_29948,N_29700);
nor UO_1345 (O_1345,N_29910,N_29777);
or UO_1346 (O_1346,N_29729,N_29741);
xnor UO_1347 (O_1347,N_29965,N_29773);
and UO_1348 (O_1348,N_29820,N_29969);
and UO_1349 (O_1349,N_29998,N_29764);
or UO_1350 (O_1350,N_29849,N_29811);
nor UO_1351 (O_1351,N_29718,N_29914);
and UO_1352 (O_1352,N_29855,N_29728);
or UO_1353 (O_1353,N_29859,N_29708);
nor UO_1354 (O_1354,N_29704,N_29820);
nor UO_1355 (O_1355,N_29846,N_29804);
nor UO_1356 (O_1356,N_29703,N_29979);
xnor UO_1357 (O_1357,N_29771,N_29965);
nor UO_1358 (O_1358,N_29849,N_29833);
and UO_1359 (O_1359,N_29817,N_29808);
or UO_1360 (O_1360,N_29982,N_29741);
nor UO_1361 (O_1361,N_29924,N_29901);
nor UO_1362 (O_1362,N_29761,N_29970);
and UO_1363 (O_1363,N_29874,N_29980);
nor UO_1364 (O_1364,N_29853,N_29968);
nand UO_1365 (O_1365,N_29982,N_29727);
xnor UO_1366 (O_1366,N_29889,N_29780);
xor UO_1367 (O_1367,N_29783,N_29859);
or UO_1368 (O_1368,N_29862,N_29705);
nor UO_1369 (O_1369,N_29975,N_29983);
xnor UO_1370 (O_1370,N_29859,N_29871);
and UO_1371 (O_1371,N_29982,N_29871);
nand UO_1372 (O_1372,N_29997,N_29841);
or UO_1373 (O_1373,N_29907,N_29882);
nand UO_1374 (O_1374,N_29817,N_29759);
xor UO_1375 (O_1375,N_29993,N_29969);
nor UO_1376 (O_1376,N_29774,N_29782);
nand UO_1377 (O_1377,N_29847,N_29885);
nand UO_1378 (O_1378,N_29887,N_29826);
or UO_1379 (O_1379,N_29871,N_29721);
or UO_1380 (O_1380,N_29745,N_29865);
xor UO_1381 (O_1381,N_29811,N_29854);
or UO_1382 (O_1382,N_29911,N_29969);
xnor UO_1383 (O_1383,N_29787,N_29750);
and UO_1384 (O_1384,N_29804,N_29805);
nand UO_1385 (O_1385,N_29994,N_29768);
or UO_1386 (O_1386,N_29920,N_29984);
nand UO_1387 (O_1387,N_29983,N_29830);
or UO_1388 (O_1388,N_29927,N_29777);
xor UO_1389 (O_1389,N_29885,N_29945);
and UO_1390 (O_1390,N_29822,N_29834);
nand UO_1391 (O_1391,N_29767,N_29721);
nor UO_1392 (O_1392,N_29746,N_29798);
and UO_1393 (O_1393,N_29729,N_29702);
nand UO_1394 (O_1394,N_29875,N_29874);
or UO_1395 (O_1395,N_29948,N_29888);
nand UO_1396 (O_1396,N_29870,N_29766);
nand UO_1397 (O_1397,N_29931,N_29779);
nor UO_1398 (O_1398,N_29973,N_29847);
nor UO_1399 (O_1399,N_29910,N_29881);
xor UO_1400 (O_1400,N_29901,N_29931);
nor UO_1401 (O_1401,N_29799,N_29982);
nand UO_1402 (O_1402,N_29894,N_29805);
or UO_1403 (O_1403,N_29718,N_29751);
or UO_1404 (O_1404,N_29994,N_29882);
and UO_1405 (O_1405,N_29838,N_29929);
nand UO_1406 (O_1406,N_29926,N_29790);
nor UO_1407 (O_1407,N_29975,N_29796);
nor UO_1408 (O_1408,N_29795,N_29842);
or UO_1409 (O_1409,N_29718,N_29948);
and UO_1410 (O_1410,N_29731,N_29853);
xnor UO_1411 (O_1411,N_29789,N_29968);
and UO_1412 (O_1412,N_29922,N_29750);
or UO_1413 (O_1413,N_29758,N_29754);
nand UO_1414 (O_1414,N_29880,N_29721);
and UO_1415 (O_1415,N_29747,N_29969);
and UO_1416 (O_1416,N_29830,N_29785);
or UO_1417 (O_1417,N_29970,N_29940);
xnor UO_1418 (O_1418,N_29916,N_29897);
or UO_1419 (O_1419,N_29856,N_29989);
and UO_1420 (O_1420,N_29897,N_29822);
or UO_1421 (O_1421,N_29987,N_29950);
nand UO_1422 (O_1422,N_29831,N_29852);
or UO_1423 (O_1423,N_29954,N_29767);
or UO_1424 (O_1424,N_29722,N_29940);
xor UO_1425 (O_1425,N_29713,N_29742);
nor UO_1426 (O_1426,N_29845,N_29932);
xor UO_1427 (O_1427,N_29884,N_29956);
nor UO_1428 (O_1428,N_29909,N_29799);
and UO_1429 (O_1429,N_29815,N_29834);
nor UO_1430 (O_1430,N_29782,N_29783);
and UO_1431 (O_1431,N_29857,N_29932);
xnor UO_1432 (O_1432,N_29825,N_29925);
nor UO_1433 (O_1433,N_29730,N_29807);
nand UO_1434 (O_1434,N_29728,N_29823);
nor UO_1435 (O_1435,N_29912,N_29902);
and UO_1436 (O_1436,N_29900,N_29763);
nor UO_1437 (O_1437,N_29795,N_29975);
nand UO_1438 (O_1438,N_29998,N_29973);
nand UO_1439 (O_1439,N_29786,N_29963);
and UO_1440 (O_1440,N_29831,N_29977);
or UO_1441 (O_1441,N_29798,N_29713);
or UO_1442 (O_1442,N_29921,N_29741);
or UO_1443 (O_1443,N_29916,N_29734);
nand UO_1444 (O_1444,N_29884,N_29908);
xor UO_1445 (O_1445,N_29770,N_29784);
nand UO_1446 (O_1446,N_29786,N_29914);
and UO_1447 (O_1447,N_29926,N_29987);
nand UO_1448 (O_1448,N_29799,N_29923);
or UO_1449 (O_1449,N_29729,N_29723);
nand UO_1450 (O_1450,N_29944,N_29712);
nand UO_1451 (O_1451,N_29905,N_29747);
or UO_1452 (O_1452,N_29874,N_29737);
or UO_1453 (O_1453,N_29959,N_29732);
nor UO_1454 (O_1454,N_29854,N_29821);
and UO_1455 (O_1455,N_29821,N_29942);
and UO_1456 (O_1456,N_29909,N_29725);
nand UO_1457 (O_1457,N_29945,N_29733);
or UO_1458 (O_1458,N_29716,N_29842);
and UO_1459 (O_1459,N_29834,N_29915);
nand UO_1460 (O_1460,N_29833,N_29961);
and UO_1461 (O_1461,N_29713,N_29782);
nand UO_1462 (O_1462,N_29942,N_29797);
nand UO_1463 (O_1463,N_29838,N_29797);
nor UO_1464 (O_1464,N_29792,N_29994);
or UO_1465 (O_1465,N_29826,N_29808);
or UO_1466 (O_1466,N_29891,N_29866);
and UO_1467 (O_1467,N_29886,N_29710);
nor UO_1468 (O_1468,N_29774,N_29930);
nor UO_1469 (O_1469,N_29888,N_29909);
nand UO_1470 (O_1470,N_29972,N_29882);
and UO_1471 (O_1471,N_29830,N_29915);
xnor UO_1472 (O_1472,N_29877,N_29883);
nor UO_1473 (O_1473,N_29740,N_29746);
xor UO_1474 (O_1474,N_29806,N_29833);
and UO_1475 (O_1475,N_29839,N_29910);
or UO_1476 (O_1476,N_29757,N_29996);
xor UO_1477 (O_1477,N_29700,N_29970);
nor UO_1478 (O_1478,N_29977,N_29852);
or UO_1479 (O_1479,N_29950,N_29841);
and UO_1480 (O_1480,N_29774,N_29850);
and UO_1481 (O_1481,N_29965,N_29983);
or UO_1482 (O_1482,N_29772,N_29905);
xnor UO_1483 (O_1483,N_29713,N_29844);
nor UO_1484 (O_1484,N_29812,N_29929);
and UO_1485 (O_1485,N_29978,N_29722);
nor UO_1486 (O_1486,N_29943,N_29716);
nand UO_1487 (O_1487,N_29735,N_29815);
nor UO_1488 (O_1488,N_29801,N_29857);
nor UO_1489 (O_1489,N_29988,N_29876);
nand UO_1490 (O_1490,N_29972,N_29731);
nand UO_1491 (O_1491,N_29857,N_29956);
nor UO_1492 (O_1492,N_29750,N_29982);
or UO_1493 (O_1493,N_29768,N_29916);
nor UO_1494 (O_1494,N_29828,N_29876);
or UO_1495 (O_1495,N_29816,N_29905);
xnor UO_1496 (O_1496,N_29954,N_29700);
xnor UO_1497 (O_1497,N_29949,N_29775);
xor UO_1498 (O_1498,N_29747,N_29793);
nor UO_1499 (O_1499,N_29891,N_29793);
xnor UO_1500 (O_1500,N_29719,N_29778);
nand UO_1501 (O_1501,N_29740,N_29760);
nor UO_1502 (O_1502,N_29977,N_29866);
xnor UO_1503 (O_1503,N_29830,N_29871);
xor UO_1504 (O_1504,N_29721,N_29792);
or UO_1505 (O_1505,N_29957,N_29848);
or UO_1506 (O_1506,N_29875,N_29741);
xnor UO_1507 (O_1507,N_29714,N_29760);
xnor UO_1508 (O_1508,N_29999,N_29890);
xor UO_1509 (O_1509,N_29953,N_29770);
or UO_1510 (O_1510,N_29923,N_29820);
nand UO_1511 (O_1511,N_29886,N_29962);
and UO_1512 (O_1512,N_29815,N_29770);
xor UO_1513 (O_1513,N_29922,N_29720);
and UO_1514 (O_1514,N_29880,N_29813);
nand UO_1515 (O_1515,N_29713,N_29786);
nand UO_1516 (O_1516,N_29976,N_29863);
nand UO_1517 (O_1517,N_29883,N_29920);
nand UO_1518 (O_1518,N_29946,N_29786);
xor UO_1519 (O_1519,N_29984,N_29949);
and UO_1520 (O_1520,N_29804,N_29927);
nand UO_1521 (O_1521,N_29973,N_29777);
xnor UO_1522 (O_1522,N_29768,N_29931);
nand UO_1523 (O_1523,N_29957,N_29831);
or UO_1524 (O_1524,N_29747,N_29840);
nor UO_1525 (O_1525,N_29736,N_29908);
or UO_1526 (O_1526,N_29902,N_29964);
xor UO_1527 (O_1527,N_29845,N_29799);
nor UO_1528 (O_1528,N_29907,N_29721);
nor UO_1529 (O_1529,N_29977,N_29832);
and UO_1530 (O_1530,N_29990,N_29931);
nand UO_1531 (O_1531,N_29740,N_29935);
or UO_1532 (O_1532,N_29999,N_29863);
or UO_1533 (O_1533,N_29838,N_29731);
or UO_1534 (O_1534,N_29861,N_29818);
nand UO_1535 (O_1535,N_29897,N_29956);
and UO_1536 (O_1536,N_29809,N_29774);
nand UO_1537 (O_1537,N_29879,N_29850);
or UO_1538 (O_1538,N_29976,N_29721);
xnor UO_1539 (O_1539,N_29728,N_29755);
nand UO_1540 (O_1540,N_29895,N_29873);
and UO_1541 (O_1541,N_29815,N_29772);
nor UO_1542 (O_1542,N_29853,N_29886);
nand UO_1543 (O_1543,N_29780,N_29869);
xor UO_1544 (O_1544,N_29896,N_29712);
and UO_1545 (O_1545,N_29984,N_29724);
and UO_1546 (O_1546,N_29922,N_29923);
xor UO_1547 (O_1547,N_29992,N_29764);
nor UO_1548 (O_1548,N_29975,N_29994);
or UO_1549 (O_1549,N_29796,N_29777);
nor UO_1550 (O_1550,N_29831,N_29816);
nor UO_1551 (O_1551,N_29874,N_29807);
and UO_1552 (O_1552,N_29700,N_29919);
nand UO_1553 (O_1553,N_29998,N_29824);
and UO_1554 (O_1554,N_29717,N_29947);
or UO_1555 (O_1555,N_29828,N_29983);
nand UO_1556 (O_1556,N_29948,N_29719);
xnor UO_1557 (O_1557,N_29837,N_29739);
and UO_1558 (O_1558,N_29955,N_29766);
nor UO_1559 (O_1559,N_29808,N_29951);
or UO_1560 (O_1560,N_29761,N_29747);
and UO_1561 (O_1561,N_29984,N_29805);
nand UO_1562 (O_1562,N_29935,N_29904);
and UO_1563 (O_1563,N_29994,N_29988);
and UO_1564 (O_1564,N_29827,N_29907);
nand UO_1565 (O_1565,N_29818,N_29757);
nor UO_1566 (O_1566,N_29970,N_29725);
and UO_1567 (O_1567,N_29729,N_29995);
and UO_1568 (O_1568,N_29772,N_29981);
and UO_1569 (O_1569,N_29962,N_29808);
xnor UO_1570 (O_1570,N_29791,N_29809);
or UO_1571 (O_1571,N_29710,N_29919);
nor UO_1572 (O_1572,N_29768,N_29914);
nor UO_1573 (O_1573,N_29759,N_29850);
and UO_1574 (O_1574,N_29739,N_29848);
nand UO_1575 (O_1575,N_29927,N_29936);
nor UO_1576 (O_1576,N_29757,N_29961);
nor UO_1577 (O_1577,N_29896,N_29752);
nand UO_1578 (O_1578,N_29723,N_29992);
nor UO_1579 (O_1579,N_29917,N_29942);
and UO_1580 (O_1580,N_29921,N_29743);
xor UO_1581 (O_1581,N_29917,N_29820);
nor UO_1582 (O_1582,N_29949,N_29872);
xor UO_1583 (O_1583,N_29908,N_29818);
nand UO_1584 (O_1584,N_29963,N_29701);
xnor UO_1585 (O_1585,N_29840,N_29713);
or UO_1586 (O_1586,N_29971,N_29847);
xor UO_1587 (O_1587,N_29974,N_29776);
nor UO_1588 (O_1588,N_29812,N_29760);
and UO_1589 (O_1589,N_29987,N_29946);
nand UO_1590 (O_1590,N_29955,N_29975);
nor UO_1591 (O_1591,N_29810,N_29744);
or UO_1592 (O_1592,N_29803,N_29862);
and UO_1593 (O_1593,N_29982,N_29941);
or UO_1594 (O_1594,N_29777,N_29835);
nor UO_1595 (O_1595,N_29970,N_29965);
or UO_1596 (O_1596,N_29796,N_29850);
and UO_1597 (O_1597,N_29787,N_29852);
and UO_1598 (O_1598,N_29895,N_29941);
nand UO_1599 (O_1599,N_29926,N_29940);
nor UO_1600 (O_1600,N_29764,N_29896);
and UO_1601 (O_1601,N_29970,N_29990);
or UO_1602 (O_1602,N_29860,N_29953);
and UO_1603 (O_1603,N_29937,N_29990);
nand UO_1604 (O_1604,N_29937,N_29763);
nand UO_1605 (O_1605,N_29861,N_29789);
and UO_1606 (O_1606,N_29768,N_29980);
nor UO_1607 (O_1607,N_29998,N_29959);
or UO_1608 (O_1608,N_29810,N_29811);
nor UO_1609 (O_1609,N_29934,N_29822);
nand UO_1610 (O_1610,N_29894,N_29905);
nand UO_1611 (O_1611,N_29959,N_29960);
nand UO_1612 (O_1612,N_29986,N_29912);
and UO_1613 (O_1613,N_29744,N_29918);
xnor UO_1614 (O_1614,N_29754,N_29755);
and UO_1615 (O_1615,N_29915,N_29769);
nand UO_1616 (O_1616,N_29955,N_29752);
nor UO_1617 (O_1617,N_29881,N_29953);
xnor UO_1618 (O_1618,N_29845,N_29741);
or UO_1619 (O_1619,N_29987,N_29960);
or UO_1620 (O_1620,N_29702,N_29943);
or UO_1621 (O_1621,N_29861,N_29700);
or UO_1622 (O_1622,N_29846,N_29741);
xor UO_1623 (O_1623,N_29761,N_29991);
and UO_1624 (O_1624,N_29860,N_29708);
nand UO_1625 (O_1625,N_29878,N_29990);
nand UO_1626 (O_1626,N_29738,N_29822);
nand UO_1627 (O_1627,N_29844,N_29754);
xnor UO_1628 (O_1628,N_29792,N_29821);
or UO_1629 (O_1629,N_29991,N_29731);
or UO_1630 (O_1630,N_29728,N_29864);
nand UO_1631 (O_1631,N_29901,N_29708);
nor UO_1632 (O_1632,N_29923,N_29768);
and UO_1633 (O_1633,N_29836,N_29817);
nor UO_1634 (O_1634,N_29884,N_29990);
nand UO_1635 (O_1635,N_29898,N_29947);
and UO_1636 (O_1636,N_29724,N_29951);
or UO_1637 (O_1637,N_29823,N_29995);
nor UO_1638 (O_1638,N_29749,N_29927);
xor UO_1639 (O_1639,N_29957,N_29943);
xor UO_1640 (O_1640,N_29767,N_29799);
or UO_1641 (O_1641,N_29837,N_29818);
nand UO_1642 (O_1642,N_29906,N_29994);
or UO_1643 (O_1643,N_29808,N_29955);
nand UO_1644 (O_1644,N_29981,N_29825);
nor UO_1645 (O_1645,N_29849,N_29728);
and UO_1646 (O_1646,N_29864,N_29816);
nand UO_1647 (O_1647,N_29719,N_29848);
nor UO_1648 (O_1648,N_29960,N_29909);
nor UO_1649 (O_1649,N_29910,N_29856);
nor UO_1650 (O_1650,N_29949,N_29928);
nand UO_1651 (O_1651,N_29985,N_29997);
and UO_1652 (O_1652,N_29878,N_29727);
and UO_1653 (O_1653,N_29704,N_29985);
nand UO_1654 (O_1654,N_29980,N_29998);
and UO_1655 (O_1655,N_29717,N_29933);
nand UO_1656 (O_1656,N_29927,N_29886);
or UO_1657 (O_1657,N_29865,N_29934);
nor UO_1658 (O_1658,N_29979,N_29868);
nor UO_1659 (O_1659,N_29720,N_29797);
or UO_1660 (O_1660,N_29919,N_29716);
and UO_1661 (O_1661,N_29702,N_29916);
nor UO_1662 (O_1662,N_29712,N_29981);
or UO_1663 (O_1663,N_29926,N_29920);
and UO_1664 (O_1664,N_29869,N_29808);
nand UO_1665 (O_1665,N_29849,N_29819);
or UO_1666 (O_1666,N_29939,N_29860);
nand UO_1667 (O_1667,N_29750,N_29900);
nand UO_1668 (O_1668,N_29871,N_29733);
nor UO_1669 (O_1669,N_29963,N_29784);
or UO_1670 (O_1670,N_29858,N_29893);
xnor UO_1671 (O_1671,N_29748,N_29736);
nand UO_1672 (O_1672,N_29740,N_29739);
xnor UO_1673 (O_1673,N_29976,N_29960);
or UO_1674 (O_1674,N_29872,N_29755);
or UO_1675 (O_1675,N_29762,N_29772);
xnor UO_1676 (O_1676,N_29917,N_29771);
nor UO_1677 (O_1677,N_29731,N_29825);
or UO_1678 (O_1678,N_29717,N_29874);
and UO_1679 (O_1679,N_29895,N_29836);
or UO_1680 (O_1680,N_29958,N_29758);
or UO_1681 (O_1681,N_29966,N_29912);
or UO_1682 (O_1682,N_29706,N_29709);
nor UO_1683 (O_1683,N_29906,N_29709);
nor UO_1684 (O_1684,N_29762,N_29769);
and UO_1685 (O_1685,N_29724,N_29804);
or UO_1686 (O_1686,N_29942,N_29868);
and UO_1687 (O_1687,N_29995,N_29876);
and UO_1688 (O_1688,N_29841,N_29700);
and UO_1689 (O_1689,N_29815,N_29715);
or UO_1690 (O_1690,N_29718,N_29714);
nand UO_1691 (O_1691,N_29795,N_29813);
nor UO_1692 (O_1692,N_29875,N_29990);
or UO_1693 (O_1693,N_29750,N_29979);
or UO_1694 (O_1694,N_29953,N_29806);
or UO_1695 (O_1695,N_29968,N_29867);
and UO_1696 (O_1696,N_29824,N_29749);
or UO_1697 (O_1697,N_29821,N_29997);
or UO_1698 (O_1698,N_29736,N_29957);
and UO_1699 (O_1699,N_29748,N_29879);
xor UO_1700 (O_1700,N_29879,N_29818);
nand UO_1701 (O_1701,N_29933,N_29978);
nand UO_1702 (O_1702,N_29965,N_29935);
nor UO_1703 (O_1703,N_29874,N_29708);
and UO_1704 (O_1704,N_29802,N_29847);
or UO_1705 (O_1705,N_29852,N_29850);
nor UO_1706 (O_1706,N_29715,N_29830);
nor UO_1707 (O_1707,N_29946,N_29716);
xor UO_1708 (O_1708,N_29894,N_29811);
and UO_1709 (O_1709,N_29745,N_29722);
nor UO_1710 (O_1710,N_29889,N_29818);
nand UO_1711 (O_1711,N_29949,N_29871);
nand UO_1712 (O_1712,N_29996,N_29827);
nand UO_1713 (O_1713,N_29731,N_29823);
nand UO_1714 (O_1714,N_29810,N_29968);
or UO_1715 (O_1715,N_29911,N_29841);
nor UO_1716 (O_1716,N_29960,N_29767);
or UO_1717 (O_1717,N_29964,N_29859);
or UO_1718 (O_1718,N_29703,N_29824);
nand UO_1719 (O_1719,N_29706,N_29974);
nand UO_1720 (O_1720,N_29707,N_29829);
and UO_1721 (O_1721,N_29979,N_29720);
and UO_1722 (O_1722,N_29976,N_29794);
xor UO_1723 (O_1723,N_29748,N_29749);
or UO_1724 (O_1724,N_29815,N_29888);
xor UO_1725 (O_1725,N_29703,N_29771);
nor UO_1726 (O_1726,N_29962,N_29769);
xor UO_1727 (O_1727,N_29766,N_29712);
nand UO_1728 (O_1728,N_29802,N_29805);
and UO_1729 (O_1729,N_29889,N_29854);
nor UO_1730 (O_1730,N_29712,N_29929);
and UO_1731 (O_1731,N_29814,N_29870);
nand UO_1732 (O_1732,N_29779,N_29732);
and UO_1733 (O_1733,N_29948,N_29702);
and UO_1734 (O_1734,N_29875,N_29843);
nor UO_1735 (O_1735,N_29972,N_29807);
nor UO_1736 (O_1736,N_29828,N_29823);
nor UO_1737 (O_1737,N_29981,N_29999);
nand UO_1738 (O_1738,N_29992,N_29885);
nand UO_1739 (O_1739,N_29934,N_29710);
nand UO_1740 (O_1740,N_29712,N_29949);
nand UO_1741 (O_1741,N_29943,N_29884);
nand UO_1742 (O_1742,N_29782,N_29984);
nand UO_1743 (O_1743,N_29861,N_29869);
or UO_1744 (O_1744,N_29780,N_29878);
nor UO_1745 (O_1745,N_29911,N_29749);
or UO_1746 (O_1746,N_29895,N_29881);
nand UO_1747 (O_1747,N_29809,N_29802);
or UO_1748 (O_1748,N_29713,N_29957);
nand UO_1749 (O_1749,N_29824,N_29879);
nand UO_1750 (O_1750,N_29944,N_29880);
and UO_1751 (O_1751,N_29938,N_29810);
or UO_1752 (O_1752,N_29890,N_29900);
xor UO_1753 (O_1753,N_29984,N_29836);
and UO_1754 (O_1754,N_29852,N_29913);
xor UO_1755 (O_1755,N_29972,N_29955);
xnor UO_1756 (O_1756,N_29778,N_29715);
nor UO_1757 (O_1757,N_29986,N_29731);
or UO_1758 (O_1758,N_29889,N_29739);
xnor UO_1759 (O_1759,N_29900,N_29950);
and UO_1760 (O_1760,N_29789,N_29710);
xnor UO_1761 (O_1761,N_29806,N_29725);
xor UO_1762 (O_1762,N_29890,N_29925);
nor UO_1763 (O_1763,N_29729,N_29839);
and UO_1764 (O_1764,N_29818,N_29867);
and UO_1765 (O_1765,N_29808,N_29785);
nor UO_1766 (O_1766,N_29969,N_29719);
nor UO_1767 (O_1767,N_29818,N_29983);
xnor UO_1768 (O_1768,N_29923,N_29739);
xnor UO_1769 (O_1769,N_29831,N_29878);
nor UO_1770 (O_1770,N_29958,N_29744);
and UO_1771 (O_1771,N_29903,N_29818);
or UO_1772 (O_1772,N_29756,N_29740);
nand UO_1773 (O_1773,N_29704,N_29881);
or UO_1774 (O_1774,N_29722,N_29962);
and UO_1775 (O_1775,N_29752,N_29991);
and UO_1776 (O_1776,N_29947,N_29880);
nor UO_1777 (O_1777,N_29976,N_29765);
and UO_1778 (O_1778,N_29929,N_29832);
nand UO_1779 (O_1779,N_29867,N_29751);
xor UO_1780 (O_1780,N_29773,N_29729);
nor UO_1781 (O_1781,N_29756,N_29719);
nor UO_1782 (O_1782,N_29798,N_29776);
xor UO_1783 (O_1783,N_29954,N_29945);
xnor UO_1784 (O_1784,N_29769,N_29927);
nand UO_1785 (O_1785,N_29759,N_29865);
nand UO_1786 (O_1786,N_29914,N_29988);
nand UO_1787 (O_1787,N_29791,N_29766);
and UO_1788 (O_1788,N_29924,N_29873);
nand UO_1789 (O_1789,N_29875,N_29914);
or UO_1790 (O_1790,N_29827,N_29809);
xnor UO_1791 (O_1791,N_29824,N_29853);
nor UO_1792 (O_1792,N_29806,N_29816);
nor UO_1793 (O_1793,N_29864,N_29814);
xor UO_1794 (O_1794,N_29787,N_29920);
or UO_1795 (O_1795,N_29708,N_29818);
and UO_1796 (O_1796,N_29743,N_29780);
and UO_1797 (O_1797,N_29790,N_29997);
and UO_1798 (O_1798,N_29957,N_29733);
and UO_1799 (O_1799,N_29789,N_29746);
or UO_1800 (O_1800,N_29985,N_29722);
or UO_1801 (O_1801,N_29738,N_29703);
xor UO_1802 (O_1802,N_29806,N_29949);
nor UO_1803 (O_1803,N_29991,N_29755);
or UO_1804 (O_1804,N_29933,N_29716);
nor UO_1805 (O_1805,N_29958,N_29770);
and UO_1806 (O_1806,N_29793,N_29853);
and UO_1807 (O_1807,N_29996,N_29748);
xnor UO_1808 (O_1808,N_29800,N_29727);
or UO_1809 (O_1809,N_29741,N_29953);
nand UO_1810 (O_1810,N_29984,N_29714);
and UO_1811 (O_1811,N_29773,N_29940);
nor UO_1812 (O_1812,N_29910,N_29734);
nor UO_1813 (O_1813,N_29797,N_29769);
nand UO_1814 (O_1814,N_29807,N_29777);
nand UO_1815 (O_1815,N_29863,N_29771);
or UO_1816 (O_1816,N_29850,N_29857);
and UO_1817 (O_1817,N_29718,N_29963);
or UO_1818 (O_1818,N_29995,N_29994);
nor UO_1819 (O_1819,N_29818,N_29958);
and UO_1820 (O_1820,N_29760,N_29789);
xnor UO_1821 (O_1821,N_29742,N_29817);
nor UO_1822 (O_1822,N_29747,N_29741);
nor UO_1823 (O_1823,N_29993,N_29728);
nor UO_1824 (O_1824,N_29893,N_29945);
or UO_1825 (O_1825,N_29905,N_29778);
xor UO_1826 (O_1826,N_29818,N_29834);
xor UO_1827 (O_1827,N_29999,N_29968);
xor UO_1828 (O_1828,N_29939,N_29856);
or UO_1829 (O_1829,N_29939,N_29930);
and UO_1830 (O_1830,N_29703,N_29961);
and UO_1831 (O_1831,N_29875,N_29761);
and UO_1832 (O_1832,N_29953,N_29763);
nand UO_1833 (O_1833,N_29762,N_29842);
xnor UO_1834 (O_1834,N_29949,N_29837);
and UO_1835 (O_1835,N_29767,N_29800);
nand UO_1836 (O_1836,N_29719,N_29949);
xor UO_1837 (O_1837,N_29959,N_29910);
xnor UO_1838 (O_1838,N_29862,N_29910);
and UO_1839 (O_1839,N_29856,N_29837);
or UO_1840 (O_1840,N_29860,N_29752);
and UO_1841 (O_1841,N_29906,N_29723);
and UO_1842 (O_1842,N_29743,N_29836);
nand UO_1843 (O_1843,N_29934,N_29973);
nand UO_1844 (O_1844,N_29943,N_29986);
and UO_1845 (O_1845,N_29931,N_29956);
xnor UO_1846 (O_1846,N_29797,N_29867);
nor UO_1847 (O_1847,N_29866,N_29999);
nor UO_1848 (O_1848,N_29976,N_29884);
nor UO_1849 (O_1849,N_29897,N_29752);
or UO_1850 (O_1850,N_29933,N_29985);
nor UO_1851 (O_1851,N_29776,N_29843);
and UO_1852 (O_1852,N_29875,N_29864);
nand UO_1853 (O_1853,N_29927,N_29724);
xnor UO_1854 (O_1854,N_29890,N_29868);
nor UO_1855 (O_1855,N_29816,N_29849);
xnor UO_1856 (O_1856,N_29865,N_29758);
and UO_1857 (O_1857,N_29716,N_29987);
xnor UO_1858 (O_1858,N_29884,N_29853);
or UO_1859 (O_1859,N_29862,N_29781);
and UO_1860 (O_1860,N_29801,N_29983);
xor UO_1861 (O_1861,N_29973,N_29705);
nand UO_1862 (O_1862,N_29994,N_29788);
or UO_1863 (O_1863,N_29759,N_29747);
nand UO_1864 (O_1864,N_29955,N_29780);
nand UO_1865 (O_1865,N_29999,N_29832);
xnor UO_1866 (O_1866,N_29849,N_29967);
nor UO_1867 (O_1867,N_29756,N_29883);
or UO_1868 (O_1868,N_29778,N_29750);
nand UO_1869 (O_1869,N_29708,N_29754);
nor UO_1870 (O_1870,N_29706,N_29741);
and UO_1871 (O_1871,N_29869,N_29703);
or UO_1872 (O_1872,N_29918,N_29887);
nor UO_1873 (O_1873,N_29726,N_29762);
nor UO_1874 (O_1874,N_29926,N_29742);
nand UO_1875 (O_1875,N_29785,N_29753);
or UO_1876 (O_1876,N_29902,N_29974);
nand UO_1877 (O_1877,N_29992,N_29997);
xnor UO_1878 (O_1878,N_29848,N_29770);
and UO_1879 (O_1879,N_29783,N_29842);
xor UO_1880 (O_1880,N_29955,N_29998);
or UO_1881 (O_1881,N_29869,N_29888);
nand UO_1882 (O_1882,N_29772,N_29920);
or UO_1883 (O_1883,N_29879,N_29981);
xor UO_1884 (O_1884,N_29859,N_29925);
or UO_1885 (O_1885,N_29771,N_29916);
xnor UO_1886 (O_1886,N_29811,N_29755);
nand UO_1887 (O_1887,N_29774,N_29727);
nor UO_1888 (O_1888,N_29764,N_29962);
nor UO_1889 (O_1889,N_29771,N_29924);
or UO_1890 (O_1890,N_29789,N_29825);
or UO_1891 (O_1891,N_29911,N_29805);
or UO_1892 (O_1892,N_29852,N_29768);
or UO_1893 (O_1893,N_29893,N_29720);
and UO_1894 (O_1894,N_29933,N_29738);
nand UO_1895 (O_1895,N_29719,N_29725);
xor UO_1896 (O_1896,N_29733,N_29944);
xnor UO_1897 (O_1897,N_29983,N_29995);
xor UO_1898 (O_1898,N_29976,N_29846);
nor UO_1899 (O_1899,N_29804,N_29813);
or UO_1900 (O_1900,N_29991,N_29852);
nor UO_1901 (O_1901,N_29937,N_29899);
nand UO_1902 (O_1902,N_29742,N_29784);
nor UO_1903 (O_1903,N_29871,N_29911);
xnor UO_1904 (O_1904,N_29728,N_29997);
nand UO_1905 (O_1905,N_29955,N_29941);
nand UO_1906 (O_1906,N_29988,N_29771);
nand UO_1907 (O_1907,N_29942,N_29885);
nand UO_1908 (O_1908,N_29829,N_29862);
nand UO_1909 (O_1909,N_29772,N_29911);
nor UO_1910 (O_1910,N_29856,N_29996);
nor UO_1911 (O_1911,N_29701,N_29931);
nand UO_1912 (O_1912,N_29849,N_29888);
or UO_1913 (O_1913,N_29726,N_29901);
nor UO_1914 (O_1914,N_29933,N_29945);
or UO_1915 (O_1915,N_29924,N_29928);
or UO_1916 (O_1916,N_29849,N_29994);
or UO_1917 (O_1917,N_29939,N_29855);
and UO_1918 (O_1918,N_29764,N_29984);
nor UO_1919 (O_1919,N_29976,N_29886);
or UO_1920 (O_1920,N_29932,N_29753);
nand UO_1921 (O_1921,N_29833,N_29951);
or UO_1922 (O_1922,N_29889,N_29781);
or UO_1923 (O_1923,N_29952,N_29932);
nand UO_1924 (O_1924,N_29897,N_29801);
and UO_1925 (O_1925,N_29710,N_29856);
or UO_1926 (O_1926,N_29999,N_29727);
xor UO_1927 (O_1927,N_29858,N_29877);
and UO_1928 (O_1928,N_29791,N_29715);
nand UO_1929 (O_1929,N_29839,N_29701);
nand UO_1930 (O_1930,N_29946,N_29995);
xnor UO_1931 (O_1931,N_29701,N_29745);
xnor UO_1932 (O_1932,N_29906,N_29957);
nor UO_1933 (O_1933,N_29841,N_29733);
and UO_1934 (O_1934,N_29873,N_29823);
or UO_1935 (O_1935,N_29903,N_29951);
nand UO_1936 (O_1936,N_29984,N_29848);
nand UO_1937 (O_1937,N_29975,N_29995);
and UO_1938 (O_1938,N_29875,N_29764);
or UO_1939 (O_1939,N_29781,N_29896);
nor UO_1940 (O_1940,N_29886,N_29829);
nor UO_1941 (O_1941,N_29837,N_29738);
nor UO_1942 (O_1942,N_29737,N_29818);
and UO_1943 (O_1943,N_29760,N_29949);
and UO_1944 (O_1944,N_29709,N_29832);
nor UO_1945 (O_1945,N_29935,N_29779);
or UO_1946 (O_1946,N_29879,N_29935);
or UO_1947 (O_1947,N_29802,N_29954);
nor UO_1948 (O_1948,N_29982,N_29732);
xnor UO_1949 (O_1949,N_29875,N_29750);
xnor UO_1950 (O_1950,N_29879,N_29949);
nand UO_1951 (O_1951,N_29869,N_29821);
nor UO_1952 (O_1952,N_29950,N_29771);
nand UO_1953 (O_1953,N_29825,N_29882);
or UO_1954 (O_1954,N_29795,N_29853);
or UO_1955 (O_1955,N_29862,N_29855);
nor UO_1956 (O_1956,N_29893,N_29735);
nand UO_1957 (O_1957,N_29716,N_29759);
and UO_1958 (O_1958,N_29900,N_29707);
nor UO_1959 (O_1959,N_29835,N_29811);
nand UO_1960 (O_1960,N_29727,N_29991);
xnor UO_1961 (O_1961,N_29918,N_29958);
and UO_1962 (O_1962,N_29707,N_29895);
and UO_1963 (O_1963,N_29894,N_29997);
and UO_1964 (O_1964,N_29816,N_29723);
and UO_1965 (O_1965,N_29739,N_29700);
xnor UO_1966 (O_1966,N_29802,N_29982);
nand UO_1967 (O_1967,N_29765,N_29807);
nand UO_1968 (O_1968,N_29770,N_29980);
nand UO_1969 (O_1969,N_29715,N_29745);
xnor UO_1970 (O_1970,N_29816,N_29896);
xor UO_1971 (O_1971,N_29914,N_29867);
or UO_1972 (O_1972,N_29867,N_29764);
nand UO_1973 (O_1973,N_29966,N_29802);
nand UO_1974 (O_1974,N_29918,N_29954);
xor UO_1975 (O_1975,N_29929,N_29796);
nor UO_1976 (O_1976,N_29736,N_29768);
nor UO_1977 (O_1977,N_29808,N_29756);
nand UO_1978 (O_1978,N_29892,N_29938);
or UO_1979 (O_1979,N_29775,N_29894);
xnor UO_1980 (O_1980,N_29778,N_29805);
or UO_1981 (O_1981,N_29784,N_29797);
or UO_1982 (O_1982,N_29999,N_29754);
nor UO_1983 (O_1983,N_29999,N_29780);
nor UO_1984 (O_1984,N_29731,N_29978);
or UO_1985 (O_1985,N_29794,N_29802);
or UO_1986 (O_1986,N_29878,N_29957);
and UO_1987 (O_1987,N_29909,N_29937);
nand UO_1988 (O_1988,N_29831,N_29847);
nor UO_1989 (O_1989,N_29891,N_29971);
xor UO_1990 (O_1990,N_29985,N_29829);
and UO_1991 (O_1991,N_29719,N_29974);
nor UO_1992 (O_1992,N_29858,N_29950);
and UO_1993 (O_1993,N_29744,N_29910);
nand UO_1994 (O_1994,N_29789,N_29725);
xnor UO_1995 (O_1995,N_29905,N_29804);
xnor UO_1996 (O_1996,N_29894,N_29886);
or UO_1997 (O_1997,N_29765,N_29987);
and UO_1998 (O_1998,N_29702,N_29828);
or UO_1999 (O_1999,N_29915,N_29843);
xnor UO_2000 (O_2000,N_29880,N_29926);
and UO_2001 (O_2001,N_29808,N_29872);
nand UO_2002 (O_2002,N_29836,N_29825);
nand UO_2003 (O_2003,N_29891,N_29730);
xor UO_2004 (O_2004,N_29920,N_29742);
or UO_2005 (O_2005,N_29798,N_29819);
xor UO_2006 (O_2006,N_29774,N_29750);
xnor UO_2007 (O_2007,N_29916,N_29942);
nand UO_2008 (O_2008,N_29829,N_29826);
nand UO_2009 (O_2009,N_29821,N_29896);
nand UO_2010 (O_2010,N_29711,N_29772);
nand UO_2011 (O_2011,N_29940,N_29972);
xnor UO_2012 (O_2012,N_29982,N_29874);
nor UO_2013 (O_2013,N_29871,N_29944);
nand UO_2014 (O_2014,N_29897,N_29900);
or UO_2015 (O_2015,N_29939,N_29851);
nor UO_2016 (O_2016,N_29864,N_29840);
xnor UO_2017 (O_2017,N_29729,N_29791);
or UO_2018 (O_2018,N_29940,N_29831);
and UO_2019 (O_2019,N_29905,N_29850);
nand UO_2020 (O_2020,N_29891,N_29940);
or UO_2021 (O_2021,N_29775,N_29849);
and UO_2022 (O_2022,N_29751,N_29803);
xnor UO_2023 (O_2023,N_29962,N_29752);
xnor UO_2024 (O_2024,N_29795,N_29761);
nand UO_2025 (O_2025,N_29993,N_29998);
nor UO_2026 (O_2026,N_29974,N_29847);
and UO_2027 (O_2027,N_29960,N_29753);
xnor UO_2028 (O_2028,N_29806,N_29713);
nor UO_2029 (O_2029,N_29798,N_29722);
or UO_2030 (O_2030,N_29807,N_29827);
xor UO_2031 (O_2031,N_29706,N_29848);
or UO_2032 (O_2032,N_29732,N_29708);
nand UO_2033 (O_2033,N_29799,N_29865);
xor UO_2034 (O_2034,N_29929,N_29780);
nand UO_2035 (O_2035,N_29916,N_29920);
and UO_2036 (O_2036,N_29780,N_29742);
nand UO_2037 (O_2037,N_29892,N_29799);
nor UO_2038 (O_2038,N_29745,N_29748);
and UO_2039 (O_2039,N_29991,N_29704);
xor UO_2040 (O_2040,N_29717,N_29721);
or UO_2041 (O_2041,N_29853,N_29925);
and UO_2042 (O_2042,N_29723,N_29849);
nor UO_2043 (O_2043,N_29838,N_29710);
nor UO_2044 (O_2044,N_29883,N_29864);
and UO_2045 (O_2045,N_29721,N_29715);
xnor UO_2046 (O_2046,N_29993,N_29988);
and UO_2047 (O_2047,N_29744,N_29733);
nor UO_2048 (O_2048,N_29902,N_29905);
nor UO_2049 (O_2049,N_29987,N_29972);
nor UO_2050 (O_2050,N_29805,N_29901);
xnor UO_2051 (O_2051,N_29782,N_29906);
or UO_2052 (O_2052,N_29750,N_29861);
or UO_2053 (O_2053,N_29851,N_29916);
and UO_2054 (O_2054,N_29958,N_29831);
nor UO_2055 (O_2055,N_29787,N_29793);
and UO_2056 (O_2056,N_29727,N_29757);
nor UO_2057 (O_2057,N_29926,N_29858);
nand UO_2058 (O_2058,N_29994,N_29938);
or UO_2059 (O_2059,N_29842,N_29845);
xor UO_2060 (O_2060,N_29974,N_29834);
nor UO_2061 (O_2061,N_29836,N_29919);
nand UO_2062 (O_2062,N_29969,N_29762);
nand UO_2063 (O_2063,N_29847,N_29977);
xor UO_2064 (O_2064,N_29976,N_29791);
nor UO_2065 (O_2065,N_29934,N_29986);
xor UO_2066 (O_2066,N_29804,N_29829);
nor UO_2067 (O_2067,N_29881,N_29794);
xor UO_2068 (O_2068,N_29986,N_29749);
nor UO_2069 (O_2069,N_29784,N_29788);
and UO_2070 (O_2070,N_29744,N_29716);
nor UO_2071 (O_2071,N_29719,N_29997);
or UO_2072 (O_2072,N_29827,N_29719);
or UO_2073 (O_2073,N_29929,N_29960);
xnor UO_2074 (O_2074,N_29821,N_29886);
nand UO_2075 (O_2075,N_29870,N_29756);
nand UO_2076 (O_2076,N_29719,N_29860);
xnor UO_2077 (O_2077,N_29867,N_29946);
and UO_2078 (O_2078,N_29903,N_29970);
nand UO_2079 (O_2079,N_29936,N_29820);
nand UO_2080 (O_2080,N_29887,N_29756);
xnor UO_2081 (O_2081,N_29946,N_29956);
nor UO_2082 (O_2082,N_29937,N_29722);
or UO_2083 (O_2083,N_29946,N_29892);
nor UO_2084 (O_2084,N_29939,N_29777);
and UO_2085 (O_2085,N_29940,N_29932);
nor UO_2086 (O_2086,N_29918,N_29806);
xnor UO_2087 (O_2087,N_29957,N_29988);
and UO_2088 (O_2088,N_29795,N_29803);
xor UO_2089 (O_2089,N_29860,N_29808);
or UO_2090 (O_2090,N_29803,N_29868);
xor UO_2091 (O_2091,N_29706,N_29954);
and UO_2092 (O_2092,N_29846,N_29911);
xnor UO_2093 (O_2093,N_29935,N_29814);
nand UO_2094 (O_2094,N_29870,N_29866);
nand UO_2095 (O_2095,N_29765,N_29931);
and UO_2096 (O_2096,N_29726,N_29976);
xnor UO_2097 (O_2097,N_29796,N_29701);
xnor UO_2098 (O_2098,N_29865,N_29907);
or UO_2099 (O_2099,N_29997,N_29745);
or UO_2100 (O_2100,N_29824,N_29918);
nor UO_2101 (O_2101,N_29946,N_29804);
and UO_2102 (O_2102,N_29745,N_29949);
nand UO_2103 (O_2103,N_29953,N_29842);
and UO_2104 (O_2104,N_29811,N_29768);
nand UO_2105 (O_2105,N_29976,N_29864);
and UO_2106 (O_2106,N_29822,N_29870);
and UO_2107 (O_2107,N_29995,N_29950);
nor UO_2108 (O_2108,N_29955,N_29750);
xnor UO_2109 (O_2109,N_29954,N_29842);
nand UO_2110 (O_2110,N_29812,N_29961);
nand UO_2111 (O_2111,N_29987,N_29702);
nor UO_2112 (O_2112,N_29809,N_29983);
xor UO_2113 (O_2113,N_29816,N_29821);
nor UO_2114 (O_2114,N_29762,N_29859);
and UO_2115 (O_2115,N_29935,N_29944);
nand UO_2116 (O_2116,N_29777,N_29737);
or UO_2117 (O_2117,N_29933,N_29715);
or UO_2118 (O_2118,N_29759,N_29999);
or UO_2119 (O_2119,N_29919,N_29711);
and UO_2120 (O_2120,N_29989,N_29783);
and UO_2121 (O_2121,N_29710,N_29759);
nor UO_2122 (O_2122,N_29920,N_29752);
or UO_2123 (O_2123,N_29728,N_29868);
nand UO_2124 (O_2124,N_29704,N_29997);
and UO_2125 (O_2125,N_29811,N_29936);
nor UO_2126 (O_2126,N_29892,N_29926);
and UO_2127 (O_2127,N_29896,N_29892);
nor UO_2128 (O_2128,N_29758,N_29974);
or UO_2129 (O_2129,N_29747,N_29885);
and UO_2130 (O_2130,N_29778,N_29771);
xnor UO_2131 (O_2131,N_29722,N_29865);
nor UO_2132 (O_2132,N_29999,N_29745);
xor UO_2133 (O_2133,N_29834,N_29864);
xnor UO_2134 (O_2134,N_29919,N_29781);
nor UO_2135 (O_2135,N_29805,N_29758);
nand UO_2136 (O_2136,N_29766,N_29974);
and UO_2137 (O_2137,N_29960,N_29817);
and UO_2138 (O_2138,N_29782,N_29796);
nor UO_2139 (O_2139,N_29907,N_29878);
xnor UO_2140 (O_2140,N_29846,N_29895);
xor UO_2141 (O_2141,N_29709,N_29925);
nand UO_2142 (O_2142,N_29865,N_29743);
and UO_2143 (O_2143,N_29845,N_29882);
nand UO_2144 (O_2144,N_29997,N_29998);
or UO_2145 (O_2145,N_29971,N_29771);
xnor UO_2146 (O_2146,N_29925,N_29861);
nand UO_2147 (O_2147,N_29767,N_29865);
nor UO_2148 (O_2148,N_29966,N_29908);
and UO_2149 (O_2149,N_29917,N_29729);
or UO_2150 (O_2150,N_29780,N_29884);
and UO_2151 (O_2151,N_29820,N_29736);
nor UO_2152 (O_2152,N_29904,N_29798);
nor UO_2153 (O_2153,N_29759,N_29893);
or UO_2154 (O_2154,N_29811,N_29809);
xnor UO_2155 (O_2155,N_29812,N_29988);
nand UO_2156 (O_2156,N_29987,N_29966);
xnor UO_2157 (O_2157,N_29958,N_29791);
or UO_2158 (O_2158,N_29867,N_29713);
nand UO_2159 (O_2159,N_29706,N_29965);
xor UO_2160 (O_2160,N_29915,N_29975);
xor UO_2161 (O_2161,N_29838,N_29949);
and UO_2162 (O_2162,N_29976,N_29821);
or UO_2163 (O_2163,N_29838,N_29923);
and UO_2164 (O_2164,N_29876,N_29905);
nand UO_2165 (O_2165,N_29887,N_29978);
nor UO_2166 (O_2166,N_29926,N_29922);
or UO_2167 (O_2167,N_29974,N_29904);
nor UO_2168 (O_2168,N_29822,N_29808);
xnor UO_2169 (O_2169,N_29942,N_29980);
xor UO_2170 (O_2170,N_29896,N_29935);
or UO_2171 (O_2171,N_29745,N_29808);
nand UO_2172 (O_2172,N_29918,N_29785);
nor UO_2173 (O_2173,N_29907,N_29832);
and UO_2174 (O_2174,N_29886,N_29873);
nand UO_2175 (O_2175,N_29799,N_29945);
and UO_2176 (O_2176,N_29955,N_29872);
xor UO_2177 (O_2177,N_29972,N_29808);
xnor UO_2178 (O_2178,N_29881,N_29804);
xnor UO_2179 (O_2179,N_29706,N_29792);
nor UO_2180 (O_2180,N_29716,N_29901);
or UO_2181 (O_2181,N_29848,N_29950);
nand UO_2182 (O_2182,N_29810,N_29794);
xnor UO_2183 (O_2183,N_29968,N_29800);
or UO_2184 (O_2184,N_29897,N_29712);
nor UO_2185 (O_2185,N_29731,N_29939);
xnor UO_2186 (O_2186,N_29974,N_29923);
xnor UO_2187 (O_2187,N_29945,N_29750);
and UO_2188 (O_2188,N_29866,N_29764);
nor UO_2189 (O_2189,N_29745,N_29829);
nand UO_2190 (O_2190,N_29953,N_29775);
nor UO_2191 (O_2191,N_29798,N_29778);
xor UO_2192 (O_2192,N_29953,N_29883);
and UO_2193 (O_2193,N_29833,N_29892);
xor UO_2194 (O_2194,N_29821,N_29860);
nor UO_2195 (O_2195,N_29826,N_29889);
nor UO_2196 (O_2196,N_29874,N_29930);
and UO_2197 (O_2197,N_29727,N_29832);
xor UO_2198 (O_2198,N_29716,N_29706);
nor UO_2199 (O_2199,N_29875,N_29891);
or UO_2200 (O_2200,N_29856,N_29924);
nor UO_2201 (O_2201,N_29935,N_29855);
xnor UO_2202 (O_2202,N_29785,N_29809);
xor UO_2203 (O_2203,N_29977,N_29865);
and UO_2204 (O_2204,N_29955,N_29912);
and UO_2205 (O_2205,N_29884,N_29968);
and UO_2206 (O_2206,N_29851,N_29877);
nor UO_2207 (O_2207,N_29769,N_29791);
or UO_2208 (O_2208,N_29711,N_29802);
xnor UO_2209 (O_2209,N_29857,N_29837);
or UO_2210 (O_2210,N_29964,N_29893);
or UO_2211 (O_2211,N_29874,N_29958);
nor UO_2212 (O_2212,N_29989,N_29951);
nand UO_2213 (O_2213,N_29704,N_29748);
or UO_2214 (O_2214,N_29922,N_29772);
or UO_2215 (O_2215,N_29968,N_29852);
xor UO_2216 (O_2216,N_29978,N_29980);
and UO_2217 (O_2217,N_29766,N_29986);
or UO_2218 (O_2218,N_29930,N_29804);
or UO_2219 (O_2219,N_29927,N_29915);
or UO_2220 (O_2220,N_29705,N_29895);
or UO_2221 (O_2221,N_29908,N_29927);
nand UO_2222 (O_2222,N_29974,N_29879);
or UO_2223 (O_2223,N_29895,N_29896);
and UO_2224 (O_2224,N_29887,N_29994);
xnor UO_2225 (O_2225,N_29811,N_29952);
or UO_2226 (O_2226,N_29946,N_29756);
and UO_2227 (O_2227,N_29818,N_29947);
xnor UO_2228 (O_2228,N_29738,N_29740);
nor UO_2229 (O_2229,N_29805,N_29815);
nor UO_2230 (O_2230,N_29995,N_29771);
nand UO_2231 (O_2231,N_29969,N_29792);
nand UO_2232 (O_2232,N_29747,N_29902);
or UO_2233 (O_2233,N_29875,N_29927);
xnor UO_2234 (O_2234,N_29975,N_29718);
and UO_2235 (O_2235,N_29755,N_29957);
nand UO_2236 (O_2236,N_29789,N_29876);
xnor UO_2237 (O_2237,N_29941,N_29748);
nor UO_2238 (O_2238,N_29753,N_29730);
and UO_2239 (O_2239,N_29866,N_29759);
and UO_2240 (O_2240,N_29936,N_29919);
nor UO_2241 (O_2241,N_29978,N_29849);
nor UO_2242 (O_2242,N_29974,N_29705);
and UO_2243 (O_2243,N_29977,N_29719);
and UO_2244 (O_2244,N_29827,N_29937);
nor UO_2245 (O_2245,N_29998,N_29854);
and UO_2246 (O_2246,N_29960,N_29866);
nor UO_2247 (O_2247,N_29895,N_29831);
xnor UO_2248 (O_2248,N_29814,N_29703);
nand UO_2249 (O_2249,N_29778,N_29960);
xor UO_2250 (O_2250,N_29905,N_29899);
and UO_2251 (O_2251,N_29972,N_29780);
or UO_2252 (O_2252,N_29848,N_29967);
xor UO_2253 (O_2253,N_29731,N_29762);
nor UO_2254 (O_2254,N_29765,N_29927);
and UO_2255 (O_2255,N_29793,N_29932);
nor UO_2256 (O_2256,N_29973,N_29994);
nand UO_2257 (O_2257,N_29800,N_29934);
nor UO_2258 (O_2258,N_29828,N_29948);
nor UO_2259 (O_2259,N_29932,N_29988);
nand UO_2260 (O_2260,N_29971,N_29886);
nand UO_2261 (O_2261,N_29700,N_29857);
nand UO_2262 (O_2262,N_29731,N_29739);
xnor UO_2263 (O_2263,N_29929,N_29915);
xor UO_2264 (O_2264,N_29721,N_29819);
xor UO_2265 (O_2265,N_29763,N_29827);
nor UO_2266 (O_2266,N_29930,N_29720);
nor UO_2267 (O_2267,N_29888,N_29991);
nand UO_2268 (O_2268,N_29749,N_29968);
nor UO_2269 (O_2269,N_29999,N_29708);
and UO_2270 (O_2270,N_29715,N_29929);
and UO_2271 (O_2271,N_29960,N_29763);
nor UO_2272 (O_2272,N_29899,N_29898);
nor UO_2273 (O_2273,N_29824,N_29921);
or UO_2274 (O_2274,N_29922,N_29956);
or UO_2275 (O_2275,N_29985,N_29918);
or UO_2276 (O_2276,N_29809,N_29709);
or UO_2277 (O_2277,N_29851,N_29710);
or UO_2278 (O_2278,N_29763,N_29816);
and UO_2279 (O_2279,N_29905,N_29884);
nand UO_2280 (O_2280,N_29843,N_29910);
nand UO_2281 (O_2281,N_29871,N_29910);
and UO_2282 (O_2282,N_29721,N_29993);
xnor UO_2283 (O_2283,N_29891,N_29753);
or UO_2284 (O_2284,N_29939,N_29829);
xor UO_2285 (O_2285,N_29858,N_29861);
nor UO_2286 (O_2286,N_29854,N_29908);
or UO_2287 (O_2287,N_29914,N_29795);
nor UO_2288 (O_2288,N_29852,N_29865);
and UO_2289 (O_2289,N_29763,N_29805);
nor UO_2290 (O_2290,N_29995,N_29998);
xor UO_2291 (O_2291,N_29964,N_29710);
nand UO_2292 (O_2292,N_29811,N_29927);
nand UO_2293 (O_2293,N_29755,N_29711);
xor UO_2294 (O_2294,N_29811,N_29938);
xnor UO_2295 (O_2295,N_29906,N_29726);
and UO_2296 (O_2296,N_29744,N_29836);
and UO_2297 (O_2297,N_29979,N_29866);
or UO_2298 (O_2298,N_29738,N_29932);
nor UO_2299 (O_2299,N_29962,N_29916);
nand UO_2300 (O_2300,N_29820,N_29919);
xor UO_2301 (O_2301,N_29774,N_29856);
and UO_2302 (O_2302,N_29917,N_29972);
nor UO_2303 (O_2303,N_29742,N_29726);
nand UO_2304 (O_2304,N_29998,N_29867);
xor UO_2305 (O_2305,N_29948,N_29751);
nor UO_2306 (O_2306,N_29978,N_29847);
xnor UO_2307 (O_2307,N_29724,N_29791);
and UO_2308 (O_2308,N_29976,N_29747);
and UO_2309 (O_2309,N_29995,N_29770);
and UO_2310 (O_2310,N_29929,N_29931);
nand UO_2311 (O_2311,N_29799,N_29711);
nor UO_2312 (O_2312,N_29968,N_29783);
nand UO_2313 (O_2313,N_29933,N_29973);
xnor UO_2314 (O_2314,N_29940,N_29805);
and UO_2315 (O_2315,N_29925,N_29896);
xnor UO_2316 (O_2316,N_29933,N_29915);
nand UO_2317 (O_2317,N_29857,N_29974);
and UO_2318 (O_2318,N_29883,N_29844);
and UO_2319 (O_2319,N_29953,N_29835);
and UO_2320 (O_2320,N_29826,N_29746);
xnor UO_2321 (O_2321,N_29719,N_29816);
nand UO_2322 (O_2322,N_29707,N_29791);
nand UO_2323 (O_2323,N_29831,N_29965);
or UO_2324 (O_2324,N_29792,N_29751);
nor UO_2325 (O_2325,N_29733,N_29851);
xnor UO_2326 (O_2326,N_29891,N_29700);
or UO_2327 (O_2327,N_29745,N_29760);
nand UO_2328 (O_2328,N_29797,N_29917);
and UO_2329 (O_2329,N_29900,N_29817);
or UO_2330 (O_2330,N_29990,N_29885);
nor UO_2331 (O_2331,N_29799,N_29961);
nor UO_2332 (O_2332,N_29771,N_29742);
xor UO_2333 (O_2333,N_29939,N_29967);
or UO_2334 (O_2334,N_29972,N_29927);
nand UO_2335 (O_2335,N_29902,N_29835);
and UO_2336 (O_2336,N_29936,N_29845);
nor UO_2337 (O_2337,N_29740,N_29777);
xor UO_2338 (O_2338,N_29893,N_29922);
nand UO_2339 (O_2339,N_29820,N_29815);
nand UO_2340 (O_2340,N_29983,N_29894);
or UO_2341 (O_2341,N_29966,N_29883);
nand UO_2342 (O_2342,N_29892,N_29826);
nor UO_2343 (O_2343,N_29987,N_29992);
nor UO_2344 (O_2344,N_29935,N_29943);
nor UO_2345 (O_2345,N_29711,N_29865);
xor UO_2346 (O_2346,N_29874,N_29754);
and UO_2347 (O_2347,N_29955,N_29976);
or UO_2348 (O_2348,N_29804,N_29981);
nor UO_2349 (O_2349,N_29821,N_29914);
nand UO_2350 (O_2350,N_29958,N_29872);
and UO_2351 (O_2351,N_29762,N_29839);
nand UO_2352 (O_2352,N_29772,N_29819);
nor UO_2353 (O_2353,N_29949,N_29844);
xor UO_2354 (O_2354,N_29802,N_29923);
and UO_2355 (O_2355,N_29996,N_29784);
nand UO_2356 (O_2356,N_29702,N_29708);
or UO_2357 (O_2357,N_29847,N_29936);
or UO_2358 (O_2358,N_29777,N_29930);
nand UO_2359 (O_2359,N_29723,N_29766);
xnor UO_2360 (O_2360,N_29736,N_29939);
nor UO_2361 (O_2361,N_29880,N_29762);
xor UO_2362 (O_2362,N_29896,N_29704);
and UO_2363 (O_2363,N_29929,N_29885);
or UO_2364 (O_2364,N_29826,N_29722);
or UO_2365 (O_2365,N_29766,N_29823);
and UO_2366 (O_2366,N_29888,N_29737);
or UO_2367 (O_2367,N_29884,N_29802);
or UO_2368 (O_2368,N_29876,N_29896);
xnor UO_2369 (O_2369,N_29799,N_29907);
nor UO_2370 (O_2370,N_29953,N_29781);
or UO_2371 (O_2371,N_29769,N_29775);
or UO_2372 (O_2372,N_29870,N_29871);
xnor UO_2373 (O_2373,N_29990,N_29873);
xnor UO_2374 (O_2374,N_29745,N_29875);
xnor UO_2375 (O_2375,N_29770,N_29860);
xor UO_2376 (O_2376,N_29731,N_29944);
or UO_2377 (O_2377,N_29729,N_29968);
nor UO_2378 (O_2378,N_29982,N_29994);
nor UO_2379 (O_2379,N_29734,N_29847);
nor UO_2380 (O_2380,N_29850,N_29959);
xor UO_2381 (O_2381,N_29865,N_29803);
and UO_2382 (O_2382,N_29981,N_29898);
xor UO_2383 (O_2383,N_29888,N_29905);
nand UO_2384 (O_2384,N_29841,N_29713);
and UO_2385 (O_2385,N_29909,N_29970);
xor UO_2386 (O_2386,N_29931,N_29921);
nand UO_2387 (O_2387,N_29747,N_29766);
nor UO_2388 (O_2388,N_29827,N_29976);
or UO_2389 (O_2389,N_29829,N_29885);
and UO_2390 (O_2390,N_29802,N_29849);
and UO_2391 (O_2391,N_29927,N_29708);
xor UO_2392 (O_2392,N_29834,N_29936);
xnor UO_2393 (O_2393,N_29895,N_29740);
or UO_2394 (O_2394,N_29951,N_29836);
and UO_2395 (O_2395,N_29903,N_29853);
xor UO_2396 (O_2396,N_29877,N_29852);
and UO_2397 (O_2397,N_29897,N_29850);
nand UO_2398 (O_2398,N_29911,N_29861);
and UO_2399 (O_2399,N_29912,N_29867);
xnor UO_2400 (O_2400,N_29703,N_29871);
or UO_2401 (O_2401,N_29985,N_29789);
xnor UO_2402 (O_2402,N_29891,N_29734);
or UO_2403 (O_2403,N_29928,N_29782);
or UO_2404 (O_2404,N_29755,N_29737);
nor UO_2405 (O_2405,N_29842,N_29967);
and UO_2406 (O_2406,N_29717,N_29857);
or UO_2407 (O_2407,N_29803,N_29883);
and UO_2408 (O_2408,N_29775,N_29954);
nand UO_2409 (O_2409,N_29865,N_29781);
or UO_2410 (O_2410,N_29720,N_29761);
xnor UO_2411 (O_2411,N_29713,N_29983);
or UO_2412 (O_2412,N_29728,N_29740);
xnor UO_2413 (O_2413,N_29966,N_29964);
and UO_2414 (O_2414,N_29736,N_29903);
nand UO_2415 (O_2415,N_29971,N_29707);
and UO_2416 (O_2416,N_29909,N_29953);
or UO_2417 (O_2417,N_29979,N_29766);
and UO_2418 (O_2418,N_29949,N_29892);
nor UO_2419 (O_2419,N_29703,N_29737);
or UO_2420 (O_2420,N_29974,N_29956);
and UO_2421 (O_2421,N_29779,N_29822);
nand UO_2422 (O_2422,N_29743,N_29714);
nand UO_2423 (O_2423,N_29800,N_29915);
or UO_2424 (O_2424,N_29780,N_29848);
or UO_2425 (O_2425,N_29890,N_29833);
nand UO_2426 (O_2426,N_29775,N_29929);
and UO_2427 (O_2427,N_29956,N_29727);
nand UO_2428 (O_2428,N_29785,N_29988);
xor UO_2429 (O_2429,N_29753,N_29704);
and UO_2430 (O_2430,N_29814,N_29911);
xor UO_2431 (O_2431,N_29988,N_29790);
nor UO_2432 (O_2432,N_29937,N_29908);
nand UO_2433 (O_2433,N_29878,N_29987);
nor UO_2434 (O_2434,N_29750,N_29901);
nor UO_2435 (O_2435,N_29751,N_29915);
or UO_2436 (O_2436,N_29804,N_29889);
nor UO_2437 (O_2437,N_29935,N_29748);
and UO_2438 (O_2438,N_29944,N_29777);
nor UO_2439 (O_2439,N_29835,N_29992);
nor UO_2440 (O_2440,N_29732,N_29863);
nor UO_2441 (O_2441,N_29793,N_29707);
nor UO_2442 (O_2442,N_29853,N_29812);
or UO_2443 (O_2443,N_29853,N_29954);
and UO_2444 (O_2444,N_29838,N_29709);
and UO_2445 (O_2445,N_29765,N_29982);
or UO_2446 (O_2446,N_29885,N_29961);
nor UO_2447 (O_2447,N_29927,N_29836);
and UO_2448 (O_2448,N_29837,N_29829);
or UO_2449 (O_2449,N_29912,N_29785);
xor UO_2450 (O_2450,N_29975,N_29803);
or UO_2451 (O_2451,N_29890,N_29873);
xnor UO_2452 (O_2452,N_29920,N_29908);
nand UO_2453 (O_2453,N_29777,N_29957);
nor UO_2454 (O_2454,N_29777,N_29961);
or UO_2455 (O_2455,N_29843,N_29858);
nand UO_2456 (O_2456,N_29951,N_29941);
or UO_2457 (O_2457,N_29923,N_29879);
nand UO_2458 (O_2458,N_29856,N_29824);
nand UO_2459 (O_2459,N_29709,N_29910);
or UO_2460 (O_2460,N_29869,N_29727);
or UO_2461 (O_2461,N_29826,N_29884);
nand UO_2462 (O_2462,N_29862,N_29888);
xor UO_2463 (O_2463,N_29733,N_29820);
nand UO_2464 (O_2464,N_29808,N_29818);
and UO_2465 (O_2465,N_29856,N_29934);
or UO_2466 (O_2466,N_29943,N_29861);
nor UO_2467 (O_2467,N_29791,N_29898);
nor UO_2468 (O_2468,N_29877,N_29831);
nor UO_2469 (O_2469,N_29753,N_29896);
or UO_2470 (O_2470,N_29729,N_29869);
and UO_2471 (O_2471,N_29801,N_29771);
or UO_2472 (O_2472,N_29702,N_29819);
and UO_2473 (O_2473,N_29718,N_29964);
xor UO_2474 (O_2474,N_29840,N_29778);
nand UO_2475 (O_2475,N_29780,N_29901);
nor UO_2476 (O_2476,N_29983,N_29829);
nand UO_2477 (O_2477,N_29706,N_29878);
nand UO_2478 (O_2478,N_29860,N_29743);
xnor UO_2479 (O_2479,N_29978,N_29792);
nor UO_2480 (O_2480,N_29863,N_29859);
nand UO_2481 (O_2481,N_29834,N_29897);
nor UO_2482 (O_2482,N_29894,N_29785);
nand UO_2483 (O_2483,N_29812,N_29749);
xor UO_2484 (O_2484,N_29947,N_29739);
and UO_2485 (O_2485,N_29939,N_29733);
and UO_2486 (O_2486,N_29741,N_29961);
or UO_2487 (O_2487,N_29752,N_29706);
xnor UO_2488 (O_2488,N_29814,N_29988);
nand UO_2489 (O_2489,N_29744,N_29950);
or UO_2490 (O_2490,N_29814,N_29851);
xnor UO_2491 (O_2491,N_29828,N_29952);
or UO_2492 (O_2492,N_29724,N_29744);
and UO_2493 (O_2493,N_29732,N_29936);
xnor UO_2494 (O_2494,N_29782,N_29715);
or UO_2495 (O_2495,N_29877,N_29975);
or UO_2496 (O_2496,N_29819,N_29991);
nand UO_2497 (O_2497,N_29950,N_29765);
nand UO_2498 (O_2498,N_29847,N_29994);
or UO_2499 (O_2499,N_29968,N_29883);
nor UO_2500 (O_2500,N_29805,N_29892);
nor UO_2501 (O_2501,N_29992,N_29977);
xor UO_2502 (O_2502,N_29954,N_29772);
nor UO_2503 (O_2503,N_29841,N_29973);
xor UO_2504 (O_2504,N_29883,N_29716);
and UO_2505 (O_2505,N_29909,N_29792);
xnor UO_2506 (O_2506,N_29873,N_29917);
nor UO_2507 (O_2507,N_29721,N_29966);
nand UO_2508 (O_2508,N_29783,N_29719);
nand UO_2509 (O_2509,N_29963,N_29714);
xor UO_2510 (O_2510,N_29800,N_29937);
nor UO_2511 (O_2511,N_29942,N_29895);
nor UO_2512 (O_2512,N_29984,N_29894);
nor UO_2513 (O_2513,N_29985,N_29976);
nor UO_2514 (O_2514,N_29888,N_29897);
xnor UO_2515 (O_2515,N_29911,N_29973);
and UO_2516 (O_2516,N_29827,N_29803);
or UO_2517 (O_2517,N_29930,N_29846);
nand UO_2518 (O_2518,N_29979,N_29863);
nand UO_2519 (O_2519,N_29796,N_29941);
nor UO_2520 (O_2520,N_29895,N_29794);
and UO_2521 (O_2521,N_29796,N_29760);
nor UO_2522 (O_2522,N_29751,N_29731);
nand UO_2523 (O_2523,N_29886,N_29704);
nand UO_2524 (O_2524,N_29744,N_29882);
or UO_2525 (O_2525,N_29754,N_29953);
nand UO_2526 (O_2526,N_29710,N_29914);
xnor UO_2527 (O_2527,N_29872,N_29790);
or UO_2528 (O_2528,N_29988,N_29953);
nand UO_2529 (O_2529,N_29967,N_29806);
nand UO_2530 (O_2530,N_29729,N_29961);
nand UO_2531 (O_2531,N_29996,N_29939);
nand UO_2532 (O_2532,N_29996,N_29728);
and UO_2533 (O_2533,N_29780,N_29897);
nor UO_2534 (O_2534,N_29985,N_29700);
and UO_2535 (O_2535,N_29761,N_29922);
and UO_2536 (O_2536,N_29739,N_29747);
nor UO_2537 (O_2537,N_29946,N_29904);
and UO_2538 (O_2538,N_29777,N_29971);
or UO_2539 (O_2539,N_29905,N_29704);
or UO_2540 (O_2540,N_29708,N_29726);
or UO_2541 (O_2541,N_29841,N_29988);
nand UO_2542 (O_2542,N_29821,N_29946);
xor UO_2543 (O_2543,N_29748,N_29896);
nor UO_2544 (O_2544,N_29991,N_29798);
nand UO_2545 (O_2545,N_29991,N_29989);
nand UO_2546 (O_2546,N_29867,N_29717);
and UO_2547 (O_2547,N_29718,N_29793);
or UO_2548 (O_2548,N_29870,N_29817);
xnor UO_2549 (O_2549,N_29907,N_29745);
and UO_2550 (O_2550,N_29721,N_29764);
and UO_2551 (O_2551,N_29732,N_29956);
or UO_2552 (O_2552,N_29861,N_29722);
and UO_2553 (O_2553,N_29783,N_29932);
nand UO_2554 (O_2554,N_29893,N_29848);
nor UO_2555 (O_2555,N_29710,N_29702);
xor UO_2556 (O_2556,N_29946,N_29790);
nand UO_2557 (O_2557,N_29713,N_29829);
or UO_2558 (O_2558,N_29779,N_29721);
nor UO_2559 (O_2559,N_29940,N_29944);
nand UO_2560 (O_2560,N_29963,N_29954);
xnor UO_2561 (O_2561,N_29799,N_29847);
nor UO_2562 (O_2562,N_29991,N_29730);
xnor UO_2563 (O_2563,N_29945,N_29782);
nor UO_2564 (O_2564,N_29849,N_29784);
or UO_2565 (O_2565,N_29863,N_29929);
nor UO_2566 (O_2566,N_29779,N_29795);
or UO_2567 (O_2567,N_29947,N_29954);
or UO_2568 (O_2568,N_29961,N_29734);
xnor UO_2569 (O_2569,N_29712,N_29940);
nor UO_2570 (O_2570,N_29989,N_29768);
nor UO_2571 (O_2571,N_29723,N_29863);
nand UO_2572 (O_2572,N_29814,N_29736);
nor UO_2573 (O_2573,N_29726,N_29956);
nand UO_2574 (O_2574,N_29774,N_29757);
xnor UO_2575 (O_2575,N_29909,N_29850);
nand UO_2576 (O_2576,N_29847,N_29884);
nor UO_2577 (O_2577,N_29981,N_29872);
nor UO_2578 (O_2578,N_29890,N_29773);
nand UO_2579 (O_2579,N_29807,N_29935);
xnor UO_2580 (O_2580,N_29931,N_29743);
xor UO_2581 (O_2581,N_29843,N_29920);
nor UO_2582 (O_2582,N_29991,N_29751);
xnor UO_2583 (O_2583,N_29977,N_29928);
or UO_2584 (O_2584,N_29976,N_29962);
nand UO_2585 (O_2585,N_29777,N_29972);
nand UO_2586 (O_2586,N_29762,N_29979);
nor UO_2587 (O_2587,N_29828,N_29722);
or UO_2588 (O_2588,N_29909,N_29809);
and UO_2589 (O_2589,N_29984,N_29925);
nor UO_2590 (O_2590,N_29950,N_29747);
nand UO_2591 (O_2591,N_29815,N_29889);
and UO_2592 (O_2592,N_29727,N_29798);
nor UO_2593 (O_2593,N_29881,N_29770);
nand UO_2594 (O_2594,N_29926,N_29954);
nand UO_2595 (O_2595,N_29746,N_29702);
nor UO_2596 (O_2596,N_29953,N_29700);
nand UO_2597 (O_2597,N_29708,N_29763);
nor UO_2598 (O_2598,N_29805,N_29721);
nor UO_2599 (O_2599,N_29847,N_29870);
or UO_2600 (O_2600,N_29983,N_29990);
and UO_2601 (O_2601,N_29772,N_29918);
nor UO_2602 (O_2602,N_29751,N_29848);
and UO_2603 (O_2603,N_29966,N_29748);
nor UO_2604 (O_2604,N_29992,N_29786);
nand UO_2605 (O_2605,N_29769,N_29923);
nor UO_2606 (O_2606,N_29961,N_29782);
nand UO_2607 (O_2607,N_29943,N_29712);
nor UO_2608 (O_2608,N_29881,N_29950);
or UO_2609 (O_2609,N_29858,N_29790);
nand UO_2610 (O_2610,N_29942,N_29706);
and UO_2611 (O_2611,N_29841,N_29807);
or UO_2612 (O_2612,N_29791,N_29869);
xnor UO_2613 (O_2613,N_29964,N_29903);
xnor UO_2614 (O_2614,N_29814,N_29924);
nor UO_2615 (O_2615,N_29700,N_29819);
or UO_2616 (O_2616,N_29790,N_29741);
or UO_2617 (O_2617,N_29956,N_29766);
xnor UO_2618 (O_2618,N_29737,N_29879);
or UO_2619 (O_2619,N_29994,N_29934);
xnor UO_2620 (O_2620,N_29825,N_29952);
xnor UO_2621 (O_2621,N_29849,N_29936);
nand UO_2622 (O_2622,N_29745,N_29930);
or UO_2623 (O_2623,N_29897,N_29976);
nor UO_2624 (O_2624,N_29954,N_29928);
nand UO_2625 (O_2625,N_29940,N_29728);
xnor UO_2626 (O_2626,N_29821,N_29814);
nand UO_2627 (O_2627,N_29810,N_29966);
nor UO_2628 (O_2628,N_29785,N_29810);
xor UO_2629 (O_2629,N_29867,N_29749);
or UO_2630 (O_2630,N_29980,N_29774);
nand UO_2631 (O_2631,N_29732,N_29907);
nor UO_2632 (O_2632,N_29788,N_29853);
xnor UO_2633 (O_2633,N_29895,N_29746);
or UO_2634 (O_2634,N_29833,N_29894);
nand UO_2635 (O_2635,N_29713,N_29825);
and UO_2636 (O_2636,N_29835,N_29978);
and UO_2637 (O_2637,N_29777,N_29843);
nand UO_2638 (O_2638,N_29901,N_29990);
nand UO_2639 (O_2639,N_29886,N_29922);
nor UO_2640 (O_2640,N_29790,N_29844);
nor UO_2641 (O_2641,N_29838,N_29811);
nor UO_2642 (O_2642,N_29758,N_29982);
or UO_2643 (O_2643,N_29715,N_29951);
nor UO_2644 (O_2644,N_29940,N_29904);
nor UO_2645 (O_2645,N_29814,N_29987);
or UO_2646 (O_2646,N_29917,N_29946);
and UO_2647 (O_2647,N_29966,N_29831);
or UO_2648 (O_2648,N_29928,N_29843);
and UO_2649 (O_2649,N_29915,N_29786);
xor UO_2650 (O_2650,N_29758,N_29867);
and UO_2651 (O_2651,N_29713,N_29953);
xor UO_2652 (O_2652,N_29831,N_29871);
or UO_2653 (O_2653,N_29904,N_29939);
xnor UO_2654 (O_2654,N_29837,N_29979);
xor UO_2655 (O_2655,N_29853,N_29862);
xnor UO_2656 (O_2656,N_29942,N_29853);
and UO_2657 (O_2657,N_29711,N_29869);
nand UO_2658 (O_2658,N_29751,N_29723);
nor UO_2659 (O_2659,N_29858,N_29928);
nor UO_2660 (O_2660,N_29975,N_29887);
nand UO_2661 (O_2661,N_29907,N_29859);
nand UO_2662 (O_2662,N_29872,N_29910);
and UO_2663 (O_2663,N_29817,N_29735);
and UO_2664 (O_2664,N_29742,N_29982);
nand UO_2665 (O_2665,N_29742,N_29747);
and UO_2666 (O_2666,N_29882,N_29754);
and UO_2667 (O_2667,N_29712,N_29921);
or UO_2668 (O_2668,N_29937,N_29814);
nor UO_2669 (O_2669,N_29816,N_29826);
or UO_2670 (O_2670,N_29812,N_29954);
nand UO_2671 (O_2671,N_29728,N_29787);
and UO_2672 (O_2672,N_29764,N_29714);
and UO_2673 (O_2673,N_29903,N_29938);
xor UO_2674 (O_2674,N_29965,N_29926);
nor UO_2675 (O_2675,N_29847,N_29915);
and UO_2676 (O_2676,N_29963,N_29988);
or UO_2677 (O_2677,N_29707,N_29996);
and UO_2678 (O_2678,N_29866,N_29905);
nand UO_2679 (O_2679,N_29785,N_29977);
and UO_2680 (O_2680,N_29944,N_29876);
xnor UO_2681 (O_2681,N_29943,N_29720);
nor UO_2682 (O_2682,N_29952,N_29746);
nor UO_2683 (O_2683,N_29792,N_29710);
and UO_2684 (O_2684,N_29966,N_29727);
nor UO_2685 (O_2685,N_29906,N_29764);
nand UO_2686 (O_2686,N_29910,N_29719);
nand UO_2687 (O_2687,N_29828,N_29942);
nor UO_2688 (O_2688,N_29772,N_29957);
nand UO_2689 (O_2689,N_29953,N_29983);
nand UO_2690 (O_2690,N_29894,N_29827);
xnor UO_2691 (O_2691,N_29932,N_29813);
nand UO_2692 (O_2692,N_29943,N_29747);
nand UO_2693 (O_2693,N_29926,N_29813);
nand UO_2694 (O_2694,N_29818,N_29859);
and UO_2695 (O_2695,N_29973,N_29825);
nand UO_2696 (O_2696,N_29794,N_29969);
xnor UO_2697 (O_2697,N_29795,N_29875);
xor UO_2698 (O_2698,N_29893,N_29929);
nor UO_2699 (O_2699,N_29915,N_29997);
nand UO_2700 (O_2700,N_29999,N_29994);
nor UO_2701 (O_2701,N_29732,N_29917);
or UO_2702 (O_2702,N_29984,N_29932);
xor UO_2703 (O_2703,N_29764,N_29902);
nor UO_2704 (O_2704,N_29892,N_29831);
and UO_2705 (O_2705,N_29745,N_29755);
or UO_2706 (O_2706,N_29766,N_29837);
or UO_2707 (O_2707,N_29966,N_29904);
and UO_2708 (O_2708,N_29782,N_29856);
xnor UO_2709 (O_2709,N_29890,N_29866);
nor UO_2710 (O_2710,N_29757,N_29754);
xnor UO_2711 (O_2711,N_29727,N_29822);
xor UO_2712 (O_2712,N_29901,N_29781);
and UO_2713 (O_2713,N_29823,N_29814);
or UO_2714 (O_2714,N_29969,N_29881);
xnor UO_2715 (O_2715,N_29852,N_29964);
nand UO_2716 (O_2716,N_29993,N_29981);
nor UO_2717 (O_2717,N_29870,N_29953);
xor UO_2718 (O_2718,N_29958,N_29859);
and UO_2719 (O_2719,N_29704,N_29866);
or UO_2720 (O_2720,N_29732,N_29802);
or UO_2721 (O_2721,N_29947,N_29844);
nor UO_2722 (O_2722,N_29789,N_29809);
nor UO_2723 (O_2723,N_29882,N_29897);
nand UO_2724 (O_2724,N_29783,N_29770);
nor UO_2725 (O_2725,N_29881,N_29785);
or UO_2726 (O_2726,N_29805,N_29993);
nand UO_2727 (O_2727,N_29855,N_29974);
nand UO_2728 (O_2728,N_29856,N_29954);
or UO_2729 (O_2729,N_29878,N_29766);
xnor UO_2730 (O_2730,N_29841,N_29965);
nor UO_2731 (O_2731,N_29966,N_29924);
xor UO_2732 (O_2732,N_29983,N_29976);
nor UO_2733 (O_2733,N_29823,N_29998);
or UO_2734 (O_2734,N_29704,N_29809);
and UO_2735 (O_2735,N_29881,N_29909);
nor UO_2736 (O_2736,N_29713,N_29748);
nand UO_2737 (O_2737,N_29777,N_29806);
xnor UO_2738 (O_2738,N_29835,N_29819);
or UO_2739 (O_2739,N_29866,N_29795);
nand UO_2740 (O_2740,N_29783,N_29870);
nand UO_2741 (O_2741,N_29758,N_29831);
nand UO_2742 (O_2742,N_29739,N_29761);
and UO_2743 (O_2743,N_29801,N_29891);
or UO_2744 (O_2744,N_29958,N_29712);
or UO_2745 (O_2745,N_29854,N_29760);
and UO_2746 (O_2746,N_29819,N_29920);
or UO_2747 (O_2747,N_29998,N_29705);
nand UO_2748 (O_2748,N_29700,N_29787);
or UO_2749 (O_2749,N_29874,N_29910);
or UO_2750 (O_2750,N_29952,N_29708);
nand UO_2751 (O_2751,N_29964,N_29918);
or UO_2752 (O_2752,N_29774,N_29929);
nor UO_2753 (O_2753,N_29876,N_29861);
nor UO_2754 (O_2754,N_29839,N_29714);
xnor UO_2755 (O_2755,N_29764,N_29900);
nand UO_2756 (O_2756,N_29758,N_29926);
nand UO_2757 (O_2757,N_29884,N_29863);
xnor UO_2758 (O_2758,N_29953,N_29732);
and UO_2759 (O_2759,N_29761,N_29773);
nand UO_2760 (O_2760,N_29953,N_29877);
xor UO_2761 (O_2761,N_29792,N_29965);
and UO_2762 (O_2762,N_29993,N_29815);
or UO_2763 (O_2763,N_29755,N_29958);
xor UO_2764 (O_2764,N_29932,N_29892);
nand UO_2765 (O_2765,N_29871,N_29723);
or UO_2766 (O_2766,N_29767,N_29837);
nor UO_2767 (O_2767,N_29713,N_29928);
nor UO_2768 (O_2768,N_29884,N_29785);
or UO_2769 (O_2769,N_29987,N_29918);
xnor UO_2770 (O_2770,N_29783,N_29736);
xnor UO_2771 (O_2771,N_29777,N_29886);
nor UO_2772 (O_2772,N_29834,N_29909);
or UO_2773 (O_2773,N_29743,N_29790);
xor UO_2774 (O_2774,N_29804,N_29856);
nand UO_2775 (O_2775,N_29793,N_29900);
or UO_2776 (O_2776,N_29816,N_29943);
nand UO_2777 (O_2777,N_29739,N_29903);
nor UO_2778 (O_2778,N_29781,N_29756);
or UO_2779 (O_2779,N_29729,N_29739);
nand UO_2780 (O_2780,N_29767,N_29714);
or UO_2781 (O_2781,N_29842,N_29899);
xor UO_2782 (O_2782,N_29900,N_29989);
and UO_2783 (O_2783,N_29952,N_29762);
and UO_2784 (O_2784,N_29856,N_29994);
or UO_2785 (O_2785,N_29956,N_29844);
or UO_2786 (O_2786,N_29943,N_29805);
or UO_2787 (O_2787,N_29780,N_29796);
or UO_2788 (O_2788,N_29938,N_29884);
nand UO_2789 (O_2789,N_29764,N_29778);
xor UO_2790 (O_2790,N_29776,N_29719);
nor UO_2791 (O_2791,N_29874,N_29742);
or UO_2792 (O_2792,N_29794,N_29747);
and UO_2793 (O_2793,N_29884,N_29999);
or UO_2794 (O_2794,N_29798,N_29896);
and UO_2795 (O_2795,N_29812,N_29723);
and UO_2796 (O_2796,N_29938,N_29711);
or UO_2797 (O_2797,N_29765,N_29745);
and UO_2798 (O_2798,N_29780,N_29758);
nand UO_2799 (O_2799,N_29872,N_29941);
nand UO_2800 (O_2800,N_29762,N_29930);
or UO_2801 (O_2801,N_29900,N_29726);
or UO_2802 (O_2802,N_29867,N_29956);
and UO_2803 (O_2803,N_29939,N_29762);
nor UO_2804 (O_2804,N_29938,N_29763);
nand UO_2805 (O_2805,N_29981,N_29951);
nand UO_2806 (O_2806,N_29929,N_29967);
xor UO_2807 (O_2807,N_29975,N_29969);
or UO_2808 (O_2808,N_29783,N_29821);
or UO_2809 (O_2809,N_29851,N_29997);
xnor UO_2810 (O_2810,N_29995,N_29800);
xor UO_2811 (O_2811,N_29940,N_29768);
or UO_2812 (O_2812,N_29868,N_29824);
or UO_2813 (O_2813,N_29794,N_29752);
and UO_2814 (O_2814,N_29712,N_29764);
or UO_2815 (O_2815,N_29726,N_29713);
and UO_2816 (O_2816,N_29966,N_29874);
nand UO_2817 (O_2817,N_29925,N_29757);
nor UO_2818 (O_2818,N_29871,N_29897);
or UO_2819 (O_2819,N_29945,N_29868);
and UO_2820 (O_2820,N_29708,N_29910);
nor UO_2821 (O_2821,N_29750,N_29840);
xnor UO_2822 (O_2822,N_29934,N_29999);
nand UO_2823 (O_2823,N_29790,N_29982);
nand UO_2824 (O_2824,N_29887,N_29787);
nand UO_2825 (O_2825,N_29739,N_29935);
nand UO_2826 (O_2826,N_29765,N_29736);
or UO_2827 (O_2827,N_29795,N_29823);
and UO_2828 (O_2828,N_29993,N_29923);
and UO_2829 (O_2829,N_29748,N_29812);
or UO_2830 (O_2830,N_29900,N_29716);
nand UO_2831 (O_2831,N_29717,N_29835);
and UO_2832 (O_2832,N_29803,N_29780);
or UO_2833 (O_2833,N_29755,N_29817);
xor UO_2834 (O_2834,N_29992,N_29827);
xor UO_2835 (O_2835,N_29762,N_29920);
and UO_2836 (O_2836,N_29704,N_29890);
nand UO_2837 (O_2837,N_29937,N_29734);
and UO_2838 (O_2838,N_29747,N_29805);
nor UO_2839 (O_2839,N_29834,N_29844);
nand UO_2840 (O_2840,N_29828,N_29979);
nand UO_2841 (O_2841,N_29931,N_29893);
nand UO_2842 (O_2842,N_29816,N_29913);
or UO_2843 (O_2843,N_29894,N_29843);
and UO_2844 (O_2844,N_29946,N_29893);
xor UO_2845 (O_2845,N_29764,N_29727);
xnor UO_2846 (O_2846,N_29992,N_29989);
or UO_2847 (O_2847,N_29796,N_29904);
and UO_2848 (O_2848,N_29802,N_29763);
and UO_2849 (O_2849,N_29768,N_29873);
and UO_2850 (O_2850,N_29920,N_29717);
nor UO_2851 (O_2851,N_29951,N_29736);
and UO_2852 (O_2852,N_29823,N_29950);
or UO_2853 (O_2853,N_29949,N_29965);
xor UO_2854 (O_2854,N_29978,N_29753);
nor UO_2855 (O_2855,N_29959,N_29709);
nand UO_2856 (O_2856,N_29813,N_29991);
and UO_2857 (O_2857,N_29974,N_29916);
or UO_2858 (O_2858,N_29737,N_29957);
nor UO_2859 (O_2859,N_29834,N_29849);
and UO_2860 (O_2860,N_29940,N_29816);
xnor UO_2861 (O_2861,N_29937,N_29735);
nor UO_2862 (O_2862,N_29910,N_29783);
and UO_2863 (O_2863,N_29956,N_29805);
nand UO_2864 (O_2864,N_29864,N_29821);
xnor UO_2865 (O_2865,N_29976,N_29704);
nor UO_2866 (O_2866,N_29777,N_29938);
or UO_2867 (O_2867,N_29803,N_29939);
and UO_2868 (O_2868,N_29792,N_29896);
nor UO_2869 (O_2869,N_29889,N_29964);
or UO_2870 (O_2870,N_29794,N_29842);
nand UO_2871 (O_2871,N_29976,N_29771);
or UO_2872 (O_2872,N_29919,N_29803);
xor UO_2873 (O_2873,N_29899,N_29979);
and UO_2874 (O_2874,N_29831,N_29963);
and UO_2875 (O_2875,N_29885,N_29744);
and UO_2876 (O_2876,N_29713,N_29908);
xnor UO_2877 (O_2877,N_29943,N_29839);
nand UO_2878 (O_2878,N_29795,N_29952);
nor UO_2879 (O_2879,N_29938,N_29719);
and UO_2880 (O_2880,N_29811,N_29987);
nor UO_2881 (O_2881,N_29914,N_29883);
nand UO_2882 (O_2882,N_29767,N_29761);
and UO_2883 (O_2883,N_29847,N_29954);
nand UO_2884 (O_2884,N_29724,N_29865);
xor UO_2885 (O_2885,N_29852,N_29733);
xnor UO_2886 (O_2886,N_29933,N_29796);
and UO_2887 (O_2887,N_29733,N_29707);
nand UO_2888 (O_2888,N_29820,N_29942);
and UO_2889 (O_2889,N_29871,N_29761);
nand UO_2890 (O_2890,N_29874,N_29844);
or UO_2891 (O_2891,N_29966,N_29728);
and UO_2892 (O_2892,N_29932,N_29745);
or UO_2893 (O_2893,N_29908,N_29835);
nor UO_2894 (O_2894,N_29903,N_29769);
and UO_2895 (O_2895,N_29915,N_29899);
xnor UO_2896 (O_2896,N_29997,N_29700);
nand UO_2897 (O_2897,N_29775,N_29838);
xnor UO_2898 (O_2898,N_29979,N_29728);
or UO_2899 (O_2899,N_29726,N_29883);
xor UO_2900 (O_2900,N_29915,N_29872);
and UO_2901 (O_2901,N_29933,N_29791);
or UO_2902 (O_2902,N_29807,N_29994);
nor UO_2903 (O_2903,N_29757,N_29837);
or UO_2904 (O_2904,N_29894,N_29834);
nand UO_2905 (O_2905,N_29795,N_29851);
xor UO_2906 (O_2906,N_29909,N_29831);
and UO_2907 (O_2907,N_29808,N_29839);
nor UO_2908 (O_2908,N_29871,N_29779);
nor UO_2909 (O_2909,N_29735,N_29986);
nor UO_2910 (O_2910,N_29942,N_29835);
nand UO_2911 (O_2911,N_29729,N_29837);
or UO_2912 (O_2912,N_29786,N_29765);
nor UO_2913 (O_2913,N_29801,N_29837);
and UO_2914 (O_2914,N_29737,N_29974);
or UO_2915 (O_2915,N_29996,N_29858);
xnor UO_2916 (O_2916,N_29709,N_29865);
xnor UO_2917 (O_2917,N_29900,N_29804);
xor UO_2918 (O_2918,N_29806,N_29820);
xor UO_2919 (O_2919,N_29929,N_29750);
or UO_2920 (O_2920,N_29753,N_29903);
nor UO_2921 (O_2921,N_29979,N_29851);
and UO_2922 (O_2922,N_29949,N_29842);
nor UO_2923 (O_2923,N_29822,N_29874);
xor UO_2924 (O_2924,N_29877,N_29929);
and UO_2925 (O_2925,N_29716,N_29849);
and UO_2926 (O_2926,N_29955,N_29921);
and UO_2927 (O_2927,N_29792,N_29766);
nor UO_2928 (O_2928,N_29877,N_29993);
xnor UO_2929 (O_2929,N_29968,N_29838);
or UO_2930 (O_2930,N_29723,N_29719);
nor UO_2931 (O_2931,N_29774,N_29982);
or UO_2932 (O_2932,N_29854,N_29932);
xnor UO_2933 (O_2933,N_29798,N_29772);
xnor UO_2934 (O_2934,N_29868,N_29947);
xor UO_2935 (O_2935,N_29843,N_29952);
nor UO_2936 (O_2936,N_29831,N_29833);
nor UO_2937 (O_2937,N_29882,N_29843);
or UO_2938 (O_2938,N_29930,N_29739);
and UO_2939 (O_2939,N_29993,N_29918);
and UO_2940 (O_2940,N_29880,N_29824);
and UO_2941 (O_2941,N_29932,N_29829);
xnor UO_2942 (O_2942,N_29998,N_29719);
nor UO_2943 (O_2943,N_29713,N_29758);
or UO_2944 (O_2944,N_29902,N_29869);
nor UO_2945 (O_2945,N_29773,N_29897);
xnor UO_2946 (O_2946,N_29716,N_29984);
xor UO_2947 (O_2947,N_29823,N_29715);
nand UO_2948 (O_2948,N_29953,N_29906);
nand UO_2949 (O_2949,N_29830,N_29994);
nor UO_2950 (O_2950,N_29767,N_29874);
nor UO_2951 (O_2951,N_29769,N_29827);
nor UO_2952 (O_2952,N_29945,N_29985);
xor UO_2953 (O_2953,N_29769,N_29906);
nand UO_2954 (O_2954,N_29877,N_29782);
and UO_2955 (O_2955,N_29908,N_29976);
or UO_2956 (O_2956,N_29885,N_29710);
nand UO_2957 (O_2957,N_29713,N_29830);
nor UO_2958 (O_2958,N_29703,N_29851);
and UO_2959 (O_2959,N_29743,N_29724);
and UO_2960 (O_2960,N_29868,N_29751);
and UO_2961 (O_2961,N_29805,N_29862);
and UO_2962 (O_2962,N_29732,N_29974);
xnor UO_2963 (O_2963,N_29710,N_29734);
nor UO_2964 (O_2964,N_29984,N_29820);
nand UO_2965 (O_2965,N_29852,N_29849);
nand UO_2966 (O_2966,N_29772,N_29848);
or UO_2967 (O_2967,N_29831,N_29769);
nor UO_2968 (O_2968,N_29797,N_29999);
or UO_2969 (O_2969,N_29856,N_29816);
nor UO_2970 (O_2970,N_29803,N_29741);
nand UO_2971 (O_2971,N_29998,N_29913);
nor UO_2972 (O_2972,N_29797,N_29871);
and UO_2973 (O_2973,N_29906,N_29793);
xor UO_2974 (O_2974,N_29701,N_29868);
xnor UO_2975 (O_2975,N_29883,N_29930);
nand UO_2976 (O_2976,N_29780,N_29804);
xnor UO_2977 (O_2977,N_29892,N_29700);
nand UO_2978 (O_2978,N_29987,N_29710);
xnor UO_2979 (O_2979,N_29997,N_29835);
nor UO_2980 (O_2980,N_29988,N_29918);
nor UO_2981 (O_2981,N_29767,N_29821);
nor UO_2982 (O_2982,N_29815,N_29763);
and UO_2983 (O_2983,N_29948,N_29910);
nand UO_2984 (O_2984,N_29773,N_29947);
nor UO_2985 (O_2985,N_29808,N_29901);
or UO_2986 (O_2986,N_29980,N_29900);
xnor UO_2987 (O_2987,N_29729,N_29959);
nand UO_2988 (O_2988,N_29704,N_29839);
nand UO_2989 (O_2989,N_29968,N_29855);
and UO_2990 (O_2990,N_29995,N_29705);
xor UO_2991 (O_2991,N_29983,N_29949);
or UO_2992 (O_2992,N_29827,N_29801);
nor UO_2993 (O_2993,N_29965,N_29875);
xnor UO_2994 (O_2994,N_29711,N_29826);
nor UO_2995 (O_2995,N_29911,N_29916);
xor UO_2996 (O_2996,N_29892,N_29873);
and UO_2997 (O_2997,N_29774,N_29903);
or UO_2998 (O_2998,N_29739,N_29866);
or UO_2999 (O_2999,N_29823,N_29864);
nor UO_3000 (O_3000,N_29727,N_29955);
xor UO_3001 (O_3001,N_29766,N_29751);
xor UO_3002 (O_3002,N_29859,N_29950);
nor UO_3003 (O_3003,N_29771,N_29943);
nand UO_3004 (O_3004,N_29907,N_29724);
nor UO_3005 (O_3005,N_29934,N_29869);
and UO_3006 (O_3006,N_29896,N_29984);
nand UO_3007 (O_3007,N_29744,N_29801);
or UO_3008 (O_3008,N_29831,N_29899);
nand UO_3009 (O_3009,N_29700,N_29973);
nor UO_3010 (O_3010,N_29784,N_29974);
xnor UO_3011 (O_3011,N_29939,N_29911);
and UO_3012 (O_3012,N_29813,N_29820);
and UO_3013 (O_3013,N_29743,N_29859);
or UO_3014 (O_3014,N_29979,N_29909);
nor UO_3015 (O_3015,N_29893,N_29933);
nand UO_3016 (O_3016,N_29987,N_29807);
nor UO_3017 (O_3017,N_29970,N_29897);
xor UO_3018 (O_3018,N_29916,N_29830);
xnor UO_3019 (O_3019,N_29965,N_29963);
nor UO_3020 (O_3020,N_29912,N_29896);
xor UO_3021 (O_3021,N_29723,N_29945);
nor UO_3022 (O_3022,N_29940,N_29976);
nor UO_3023 (O_3023,N_29879,N_29715);
or UO_3024 (O_3024,N_29763,N_29773);
or UO_3025 (O_3025,N_29998,N_29895);
or UO_3026 (O_3026,N_29755,N_29855);
nand UO_3027 (O_3027,N_29834,N_29881);
xnor UO_3028 (O_3028,N_29816,N_29720);
xor UO_3029 (O_3029,N_29705,N_29985);
nor UO_3030 (O_3030,N_29946,N_29881);
nor UO_3031 (O_3031,N_29711,N_29811);
xor UO_3032 (O_3032,N_29780,N_29960);
nor UO_3033 (O_3033,N_29984,N_29927);
xor UO_3034 (O_3034,N_29814,N_29890);
or UO_3035 (O_3035,N_29727,N_29758);
nor UO_3036 (O_3036,N_29767,N_29878);
nand UO_3037 (O_3037,N_29940,N_29975);
nand UO_3038 (O_3038,N_29880,N_29737);
xnor UO_3039 (O_3039,N_29714,N_29703);
xnor UO_3040 (O_3040,N_29969,N_29781);
nand UO_3041 (O_3041,N_29780,N_29752);
nor UO_3042 (O_3042,N_29824,N_29724);
xnor UO_3043 (O_3043,N_29808,N_29909);
or UO_3044 (O_3044,N_29875,N_29729);
nand UO_3045 (O_3045,N_29712,N_29803);
nor UO_3046 (O_3046,N_29891,N_29873);
xor UO_3047 (O_3047,N_29955,N_29856);
or UO_3048 (O_3048,N_29748,N_29786);
nand UO_3049 (O_3049,N_29715,N_29907);
nand UO_3050 (O_3050,N_29812,N_29822);
or UO_3051 (O_3051,N_29769,N_29985);
nand UO_3052 (O_3052,N_29929,N_29705);
xnor UO_3053 (O_3053,N_29922,N_29975);
or UO_3054 (O_3054,N_29957,N_29843);
nand UO_3055 (O_3055,N_29839,N_29935);
nand UO_3056 (O_3056,N_29793,N_29909);
nor UO_3057 (O_3057,N_29843,N_29937);
nor UO_3058 (O_3058,N_29965,N_29832);
nand UO_3059 (O_3059,N_29800,N_29983);
xor UO_3060 (O_3060,N_29776,N_29721);
nor UO_3061 (O_3061,N_29757,N_29866);
xor UO_3062 (O_3062,N_29939,N_29929);
and UO_3063 (O_3063,N_29751,N_29722);
nand UO_3064 (O_3064,N_29853,N_29927);
nor UO_3065 (O_3065,N_29722,N_29708);
and UO_3066 (O_3066,N_29966,N_29803);
xnor UO_3067 (O_3067,N_29876,N_29826);
nand UO_3068 (O_3068,N_29814,N_29922);
nor UO_3069 (O_3069,N_29983,N_29951);
xor UO_3070 (O_3070,N_29987,N_29978);
and UO_3071 (O_3071,N_29954,N_29857);
and UO_3072 (O_3072,N_29768,N_29767);
nand UO_3073 (O_3073,N_29757,N_29775);
or UO_3074 (O_3074,N_29809,N_29879);
nand UO_3075 (O_3075,N_29755,N_29964);
nor UO_3076 (O_3076,N_29958,N_29786);
nor UO_3077 (O_3077,N_29772,N_29838);
xnor UO_3078 (O_3078,N_29874,N_29862);
or UO_3079 (O_3079,N_29795,N_29855);
and UO_3080 (O_3080,N_29751,N_29744);
and UO_3081 (O_3081,N_29970,N_29729);
and UO_3082 (O_3082,N_29826,N_29709);
and UO_3083 (O_3083,N_29759,N_29796);
and UO_3084 (O_3084,N_29751,N_29919);
and UO_3085 (O_3085,N_29993,N_29780);
xnor UO_3086 (O_3086,N_29866,N_29978);
or UO_3087 (O_3087,N_29812,N_29900);
xor UO_3088 (O_3088,N_29896,N_29709);
or UO_3089 (O_3089,N_29855,N_29959);
or UO_3090 (O_3090,N_29809,N_29963);
and UO_3091 (O_3091,N_29893,N_29958);
nor UO_3092 (O_3092,N_29729,N_29733);
nor UO_3093 (O_3093,N_29876,N_29996);
nand UO_3094 (O_3094,N_29987,N_29979);
xnor UO_3095 (O_3095,N_29712,N_29705);
nand UO_3096 (O_3096,N_29852,N_29920);
nand UO_3097 (O_3097,N_29822,N_29944);
xnor UO_3098 (O_3098,N_29856,N_29758);
and UO_3099 (O_3099,N_29844,N_29842);
or UO_3100 (O_3100,N_29748,N_29789);
nand UO_3101 (O_3101,N_29831,N_29884);
nand UO_3102 (O_3102,N_29922,N_29853);
and UO_3103 (O_3103,N_29900,N_29855);
or UO_3104 (O_3104,N_29753,N_29926);
or UO_3105 (O_3105,N_29921,N_29814);
nor UO_3106 (O_3106,N_29754,N_29857);
or UO_3107 (O_3107,N_29962,N_29790);
nor UO_3108 (O_3108,N_29934,N_29727);
nor UO_3109 (O_3109,N_29728,N_29903);
nor UO_3110 (O_3110,N_29790,N_29805);
nor UO_3111 (O_3111,N_29968,N_29745);
or UO_3112 (O_3112,N_29775,N_29853);
nor UO_3113 (O_3113,N_29904,N_29997);
or UO_3114 (O_3114,N_29861,N_29878);
nand UO_3115 (O_3115,N_29884,N_29914);
nand UO_3116 (O_3116,N_29807,N_29781);
nand UO_3117 (O_3117,N_29870,N_29989);
nand UO_3118 (O_3118,N_29913,N_29948);
and UO_3119 (O_3119,N_29700,N_29738);
xor UO_3120 (O_3120,N_29916,N_29809);
xnor UO_3121 (O_3121,N_29917,N_29742);
and UO_3122 (O_3122,N_29829,N_29778);
or UO_3123 (O_3123,N_29906,N_29837);
and UO_3124 (O_3124,N_29815,N_29979);
and UO_3125 (O_3125,N_29864,N_29793);
xor UO_3126 (O_3126,N_29815,N_29896);
nor UO_3127 (O_3127,N_29723,N_29709);
xor UO_3128 (O_3128,N_29952,N_29984);
xor UO_3129 (O_3129,N_29783,N_29826);
nor UO_3130 (O_3130,N_29963,N_29724);
nand UO_3131 (O_3131,N_29795,N_29938);
or UO_3132 (O_3132,N_29825,N_29745);
or UO_3133 (O_3133,N_29857,N_29877);
nor UO_3134 (O_3134,N_29710,N_29925);
nand UO_3135 (O_3135,N_29777,N_29716);
and UO_3136 (O_3136,N_29858,N_29891);
nor UO_3137 (O_3137,N_29755,N_29762);
nand UO_3138 (O_3138,N_29711,N_29952);
xnor UO_3139 (O_3139,N_29960,N_29919);
nand UO_3140 (O_3140,N_29764,N_29754);
nor UO_3141 (O_3141,N_29756,N_29802);
xor UO_3142 (O_3142,N_29785,N_29940);
or UO_3143 (O_3143,N_29900,N_29865);
xnor UO_3144 (O_3144,N_29811,N_29704);
or UO_3145 (O_3145,N_29731,N_29876);
and UO_3146 (O_3146,N_29793,N_29986);
xnor UO_3147 (O_3147,N_29796,N_29765);
and UO_3148 (O_3148,N_29969,N_29848);
xor UO_3149 (O_3149,N_29975,N_29941);
or UO_3150 (O_3150,N_29800,N_29909);
xor UO_3151 (O_3151,N_29788,N_29731);
and UO_3152 (O_3152,N_29721,N_29959);
nor UO_3153 (O_3153,N_29773,N_29856);
or UO_3154 (O_3154,N_29955,N_29935);
xnor UO_3155 (O_3155,N_29873,N_29758);
nand UO_3156 (O_3156,N_29856,N_29925);
or UO_3157 (O_3157,N_29873,N_29921);
and UO_3158 (O_3158,N_29957,N_29869);
nor UO_3159 (O_3159,N_29702,N_29869);
nand UO_3160 (O_3160,N_29923,N_29891);
or UO_3161 (O_3161,N_29943,N_29731);
or UO_3162 (O_3162,N_29954,N_29788);
xor UO_3163 (O_3163,N_29757,N_29747);
nor UO_3164 (O_3164,N_29885,N_29965);
xnor UO_3165 (O_3165,N_29785,N_29893);
xor UO_3166 (O_3166,N_29820,N_29732);
or UO_3167 (O_3167,N_29907,N_29871);
or UO_3168 (O_3168,N_29724,N_29796);
nand UO_3169 (O_3169,N_29881,N_29957);
or UO_3170 (O_3170,N_29721,N_29854);
and UO_3171 (O_3171,N_29718,N_29959);
and UO_3172 (O_3172,N_29953,N_29912);
and UO_3173 (O_3173,N_29723,N_29803);
and UO_3174 (O_3174,N_29890,N_29894);
xnor UO_3175 (O_3175,N_29931,N_29961);
xnor UO_3176 (O_3176,N_29988,N_29793);
and UO_3177 (O_3177,N_29864,N_29933);
nor UO_3178 (O_3178,N_29912,N_29868);
xor UO_3179 (O_3179,N_29990,N_29818);
xor UO_3180 (O_3180,N_29726,N_29943);
and UO_3181 (O_3181,N_29857,N_29891);
and UO_3182 (O_3182,N_29886,N_29957);
nor UO_3183 (O_3183,N_29702,N_29849);
or UO_3184 (O_3184,N_29927,N_29770);
and UO_3185 (O_3185,N_29777,N_29905);
and UO_3186 (O_3186,N_29982,N_29963);
nor UO_3187 (O_3187,N_29755,N_29851);
or UO_3188 (O_3188,N_29807,N_29910);
nor UO_3189 (O_3189,N_29877,N_29873);
xnor UO_3190 (O_3190,N_29882,N_29797);
and UO_3191 (O_3191,N_29766,N_29869);
nor UO_3192 (O_3192,N_29842,N_29923);
or UO_3193 (O_3193,N_29740,N_29813);
or UO_3194 (O_3194,N_29977,N_29915);
nand UO_3195 (O_3195,N_29977,N_29854);
or UO_3196 (O_3196,N_29722,N_29998);
xor UO_3197 (O_3197,N_29770,N_29829);
and UO_3198 (O_3198,N_29749,N_29979);
or UO_3199 (O_3199,N_29728,N_29808);
nand UO_3200 (O_3200,N_29798,N_29910);
nand UO_3201 (O_3201,N_29767,N_29947);
nor UO_3202 (O_3202,N_29905,N_29879);
and UO_3203 (O_3203,N_29723,N_29907);
nand UO_3204 (O_3204,N_29924,N_29781);
or UO_3205 (O_3205,N_29904,N_29995);
or UO_3206 (O_3206,N_29971,N_29743);
xor UO_3207 (O_3207,N_29934,N_29853);
nand UO_3208 (O_3208,N_29711,N_29893);
xnor UO_3209 (O_3209,N_29797,N_29759);
nor UO_3210 (O_3210,N_29750,N_29876);
nand UO_3211 (O_3211,N_29812,N_29752);
nand UO_3212 (O_3212,N_29759,N_29981);
and UO_3213 (O_3213,N_29741,N_29752);
nand UO_3214 (O_3214,N_29806,N_29959);
or UO_3215 (O_3215,N_29981,N_29790);
nor UO_3216 (O_3216,N_29718,N_29744);
xnor UO_3217 (O_3217,N_29860,N_29731);
and UO_3218 (O_3218,N_29937,N_29768);
or UO_3219 (O_3219,N_29886,N_29828);
or UO_3220 (O_3220,N_29828,N_29708);
nor UO_3221 (O_3221,N_29894,N_29725);
nand UO_3222 (O_3222,N_29976,N_29982);
xnor UO_3223 (O_3223,N_29774,N_29993);
nor UO_3224 (O_3224,N_29725,N_29728);
nand UO_3225 (O_3225,N_29820,N_29725);
or UO_3226 (O_3226,N_29911,N_29859);
nand UO_3227 (O_3227,N_29726,N_29878);
or UO_3228 (O_3228,N_29806,N_29910);
nand UO_3229 (O_3229,N_29826,N_29763);
nand UO_3230 (O_3230,N_29865,N_29933);
or UO_3231 (O_3231,N_29842,N_29775);
nand UO_3232 (O_3232,N_29706,N_29876);
or UO_3233 (O_3233,N_29739,N_29768);
nor UO_3234 (O_3234,N_29959,N_29945);
xor UO_3235 (O_3235,N_29711,N_29993);
or UO_3236 (O_3236,N_29931,N_29964);
or UO_3237 (O_3237,N_29779,N_29785);
xnor UO_3238 (O_3238,N_29994,N_29708);
or UO_3239 (O_3239,N_29726,N_29719);
or UO_3240 (O_3240,N_29802,N_29995);
nand UO_3241 (O_3241,N_29864,N_29944);
nand UO_3242 (O_3242,N_29983,N_29835);
or UO_3243 (O_3243,N_29777,N_29912);
or UO_3244 (O_3244,N_29983,N_29788);
or UO_3245 (O_3245,N_29821,N_29911);
nand UO_3246 (O_3246,N_29897,N_29961);
and UO_3247 (O_3247,N_29945,N_29726);
or UO_3248 (O_3248,N_29850,N_29745);
nor UO_3249 (O_3249,N_29984,N_29723);
nand UO_3250 (O_3250,N_29874,N_29904);
or UO_3251 (O_3251,N_29972,N_29905);
or UO_3252 (O_3252,N_29841,N_29956);
xnor UO_3253 (O_3253,N_29707,N_29738);
or UO_3254 (O_3254,N_29839,N_29739);
or UO_3255 (O_3255,N_29708,N_29890);
or UO_3256 (O_3256,N_29757,N_29977);
or UO_3257 (O_3257,N_29860,N_29920);
and UO_3258 (O_3258,N_29940,N_29845);
nor UO_3259 (O_3259,N_29746,N_29744);
and UO_3260 (O_3260,N_29834,N_29785);
nand UO_3261 (O_3261,N_29988,N_29987);
nor UO_3262 (O_3262,N_29929,N_29945);
nor UO_3263 (O_3263,N_29700,N_29895);
nand UO_3264 (O_3264,N_29760,N_29810);
nand UO_3265 (O_3265,N_29908,N_29861);
nor UO_3266 (O_3266,N_29867,N_29921);
nand UO_3267 (O_3267,N_29770,N_29974);
nor UO_3268 (O_3268,N_29714,N_29821);
and UO_3269 (O_3269,N_29793,N_29901);
xor UO_3270 (O_3270,N_29740,N_29970);
xnor UO_3271 (O_3271,N_29981,N_29715);
nor UO_3272 (O_3272,N_29978,N_29732);
nand UO_3273 (O_3273,N_29892,N_29719);
nor UO_3274 (O_3274,N_29829,N_29907);
and UO_3275 (O_3275,N_29711,N_29805);
xnor UO_3276 (O_3276,N_29826,N_29802);
nor UO_3277 (O_3277,N_29828,N_29995);
xnor UO_3278 (O_3278,N_29891,N_29727);
and UO_3279 (O_3279,N_29778,N_29998);
nor UO_3280 (O_3280,N_29853,N_29805);
and UO_3281 (O_3281,N_29975,N_29712);
xnor UO_3282 (O_3282,N_29789,N_29793);
or UO_3283 (O_3283,N_29749,N_29720);
and UO_3284 (O_3284,N_29978,N_29897);
and UO_3285 (O_3285,N_29812,N_29858);
nor UO_3286 (O_3286,N_29788,N_29702);
and UO_3287 (O_3287,N_29990,N_29996);
xnor UO_3288 (O_3288,N_29718,N_29705);
or UO_3289 (O_3289,N_29998,N_29963);
nor UO_3290 (O_3290,N_29794,N_29729);
nor UO_3291 (O_3291,N_29703,N_29957);
nand UO_3292 (O_3292,N_29864,N_29745);
nand UO_3293 (O_3293,N_29856,N_29960);
or UO_3294 (O_3294,N_29763,N_29749);
and UO_3295 (O_3295,N_29972,N_29946);
nand UO_3296 (O_3296,N_29708,N_29867);
nor UO_3297 (O_3297,N_29909,N_29907);
or UO_3298 (O_3298,N_29809,N_29814);
or UO_3299 (O_3299,N_29955,N_29928);
nand UO_3300 (O_3300,N_29809,N_29782);
nand UO_3301 (O_3301,N_29852,N_29758);
xnor UO_3302 (O_3302,N_29841,N_29761);
or UO_3303 (O_3303,N_29901,N_29835);
and UO_3304 (O_3304,N_29809,N_29980);
or UO_3305 (O_3305,N_29883,N_29979);
nand UO_3306 (O_3306,N_29749,N_29910);
xnor UO_3307 (O_3307,N_29834,N_29817);
and UO_3308 (O_3308,N_29940,N_29738);
xor UO_3309 (O_3309,N_29888,N_29750);
xor UO_3310 (O_3310,N_29717,N_29901);
and UO_3311 (O_3311,N_29765,N_29818);
xnor UO_3312 (O_3312,N_29862,N_29774);
xnor UO_3313 (O_3313,N_29942,N_29873);
nor UO_3314 (O_3314,N_29905,N_29708);
nand UO_3315 (O_3315,N_29869,N_29967);
nor UO_3316 (O_3316,N_29935,N_29735);
xnor UO_3317 (O_3317,N_29826,N_29962);
xnor UO_3318 (O_3318,N_29716,N_29866);
and UO_3319 (O_3319,N_29974,N_29760);
xnor UO_3320 (O_3320,N_29862,N_29975);
or UO_3321 (O_3321,N_29768,N_29754);
nor UO_3322 (O_3322,N_29983,N_29885);
nor UO_3323 (O_3323,N_29825,N_29985);
nand UO_3324 (O_3324,N_29945,N_29843);
and UO_3325 (O_3325,N_29883,N_29845);
nor UO_3326 (O_3326,N_29799,N_29977);
nor UO_3327 (O_3327,N_29838,N_29995);
nand UO_3328 (O_3328,N_29835,N_29791);
nor UO_3329 (O_3329,N_29989,N_29718);
and UO_3330 (O_3330,N_29952,N_29928);
xnor UO_3331 (O_3331,N_29918,N_29909);
nand UO_3332 (O_3332,N_29990,N_29744);
xor UO_3333 (O_3333,N_29729,N_29960);
nand UO_3334 (O_3334,N_29744,N_29991);
nor UO_3335 (O_3335,N_29717,N_29831);
xor UO_3336 (O_3336,N_29857,N_29790);
xnor UO_3337 (O_3337,N_29943,N_29780);
nand UO_3338 (O_3338,N_29777,N_29816);
or UO_3339 (O_3339,N_29847,N_29726);
or UO_3340 (O_3340,N_29792,N_29835);
and UO_3341 (O_3341,N_29778,N_29710);
nor UO_3342 (O_3342,N_29868,N_29734);
nand UO_3343 (O_3343,N_29776,N_29791);
xnor UO_3344 (O_3344,N_29963,N_29835);
or UO_3345 (O_3345,N_29816,N_29947);
and UO_3346 (O_3346,N_29971,N_29903);
xor UO_3347 (O_3347,N_29883,N_29927);
nor UO_3348 (O_3348,N_29778,N_29777);
xor UO_3349 (O_3349,N_29720,N_29775);
and UO_3350 (O_3350,N_29975,N_29996);
nand UO_3351 (O_3351,N_29781,N_29772);
nor UO_3352 (O_3352,N_29726,N_29709);
nand UO_3353 (O_3353,N_29747,N_29821);
xnor UO_3354 (O_3354,N_29749,N_29783);
and UO_3355 (O_3355,N_29787,N_29904);
nand UO_3356 (O_3356,N_29843,N_29908);
and UO_3357 (O_3357,N_29847,N_29930);
xor UO_3358 (O_3358,N_29828,N_29987);
nand UO_3359 (O_3359,N_29985,N_29779);
xnor UO_3360 (O_3360,N_29828,N_29937);
and UO_3361 (O_3361,N_29713,N_29714);
nor UO_3362 (O_3362,N_29778,N_29762);
nor UO_3363 (O_3363,N_29990,N_29888);
or UO_3364 (O_3364,N_29989,N_29995);
xnor UO_3365 (O_3365,N_29711,N_29737);
nand UO_3366 (O_3366,N_29702,N_29744);
and UO_3367 (O_3367,N_29778,N_29801);
xnor UO_3368 (O_3368,N_29936,N_29770);
xnor UO_3369 (O_3369,N_29937,N_29761);
and UO_3370 (O_3370,N_29739,N_29780);
nor UO_3371 (O_3371,N_29841,N_29745);
and UO_3372 (O_3372,N_29902,N_29855);
nor UO_3373 (O_3373,N_29813,N_29960);
nor UO_3374 (O_3374,N_29988,N_29835);
nor UO_3375 (O_3375,N_29969,N_29824);
or UO_3376 (O_3376,N_29707,N_29976);
xnor UO_3377 (O_3377,N_29907,N_29749);
nand UO_3378 (O_3378,N_29898,N_29857);
nor UO_3379 (O_3379,N_29812,N_29722);
or UO_3380 (O_3380,N_29747,N_29701);
nor UO_3381 (O_3381,N_29740,N_29796);
xor UO_3382 (O_3382,N_29858,N_29967);
and UO_3383 (O_3383,N_29985,N_29923);
xnor UO_3384 (O_3384,N_29738,N_29824);
nand UO_3385 (O_3385,N_29803,N_29947);
nor UO_3386 (O_3386,N_29795,N_29802);
nand UO_3387 (O_3387,N_29921,N_29945);
and UO_3388 (O_3388,N_29865,N_29849);
nor UO_3389 (O_3389,N_29981,N_29735);
or UO_3390 (O_3390,N_29934,N_29790);
and UO_3391 (O_3391,N_29905,N_29810);
or UO_3392 (O_3392,N_29807,N_29871);
or UO_3393 (O_3393,N_29841,N_29820);
and UO_3394 (O_3394,N_29959,N_29746);
nor UO_3395 (O_3395,N_29988,N_29774);
nand UO_3396 (O_3396,N_29765,N_29824);
xnor UO_3397 (O_3397,N_29992,N_29940);
and UO_3398 (O_3398,N_29789,N_29715);
and UO_3399 (O_3399,N_29904,N_29723);
or UO_3400 (O_3400,N_29798,N_29959);
nor UO_3401 (O_3401,N_29993,N_29989);
and UO_3402 (O_3402,N_29983,N_29900);
nand UO_3403 (O_3403,N_29915,N_29928);
xnor UO_3404 (O_3404,N_29864,N_29888);
or UO_3405 (O_3405,N_29912,N_29876);
and UO_3406 (O_3406,N_29756,N_29826);
or UO_3407 (O_3407,N_29784,N_29946);
xor UO_3408 (O_3408,N_29724,N_29916);
and UO_3409 (O_3409,N_29781,N_29944);
nor UO_3410 (O_3410,N_29949,N_29991);
or UO_3411 (O_3411,N_29989,N_29841);
xnor UO_3412 (O_3412,N_29861,N_29946);
and UO_3413 (O_3413,N_29917,N_29828);
and UO_3414 (O_3414,N_29892,N_29874);
nand UO_3415 (O_3415,N_29831,N_29753);
nor UO_3416 (O_3416,N_29910,N_29849);
nor UO_3417 (O_3417,N_29989,N_29907);
and UO_3418 (O_3418,N_29866,N_29808);
and UO_3419 (O_3419,N_29707,N_29896);
and UO_3420 (O_3420,N_29814,N_29984);
and UO_3421 (O_3421,N_29905,N_29759);
nand UO_3422 (O_3422,N_29857,N_29913);
nand UO_3423 (O_3423,N_29948,N_29952);
xor UO_3424 (O_3424,N_29886,N_29764);
xor UO_3425 (O_3425,N_29831,N_29997);
xor UO_3426 (O_3426,N_29926,N_29809);
and UO_3427 (O_3427,N_29955,N_29788);
or UO_3428 (O_3428,N_29912,N_29976);
nand UO_3429 (O_3429,N_29956,N_29757);
nor UO_3430 (O_3430,N_29894,N_29969);
nor UO_3431 (O_3431,N_29849,N_29968);
nor UO_3432 (O_3432,N_29871,N_29770);
and UO_3433 (O_3433,N_29745,N_29735);
nand UO_3434 (O_3434,N_29794,N_29928);
nor UO_3435 (O_3435,N_29853,N_29882);
or UO_3436 (O_3436,N_29840,N_29827);
nand UO_3437 (O_3437,N_29756,N_29833);
nor UO_3438 (O_3438,N_29923,N_29777);
xor UO_3439 (O_3439,N_29993,N_29930);
nor UO_3440 (O_3440,N_29709,N_29821);
xnor UO_3441 (O_3441,N_29741,N_29894);
nor UO_3442 (O_3442,N_29959,N_29750);
or UO_3443 (O_3443,N_29854,N_29868);
or UO_3444 (O_3444,N_29791,N_29995);
nor UO_3445 (O_3445,N_29715,N_29718);
nand UO_3446 (O_3446,N_29889,N_29709);
and UO_3447 (O_3447,N_29787,N_29979);
xnor UO_3448 (O_3448,N_29970,N_29873);
and UO_3449 (O_3449,N_29885,N_29934);
xor UO_3450 (O_3450,N_29946,N_29963);
xor UO_3451 (O_3451,N_29843,N_29896);
or UO_3452 (O_3452,N_29779,N_29851);
and UO_3453 (O_3453,N_29745,N_29820);
xnor UO_3454 (O_3454,N_29908,N_29953);
nand UO_3455 (O_3455,N_29990,N_29803);
and UO_3456 (O_3456,N_29994,N_29713);
xor UO_3457 (O_3457,N_29786,N_29822);
nand UO_3458 (O_3458,N_29795,N_29894);
and UO_3459 (O_3459,N_29761,N_29755);
nand UO_3460 (O_3460,N_29965,N_29788);
and UO_3461 (O_3461,N_29873,N_29911);
nand UO_3462 (O_3462,N_29800,N_29717);
or UO_3463 (O_3463,N_29887,N_29779);
nand UO_3464 (O_3464,N_29848,N_29709);
or UO_3465 (O_3465,N_29701,N_29718);
nor UO_3466 (O_3466,N_29804,N_29891);
or UO_3467 (O_3467,N_29846,N_29844);
and UO_3468 (O_3468,N_29724,N_29766);
nand UO_3469 (O_3469,N_29873,N_29901);
and UO_3470 (O_3470,N_29990,N_29961);
xnor UO_3471 (O_3471,N_29851,N_29918);
xor UO_3472 (O_3472,N_29950,N_29891);
nor UO_3473 (O_3473,N_29881,N_29702);
nand UO_3474 (O_3474,N_29800,N_29792);
xor UO_3475 (O_3475,N_29981,N_29869);
nor UO_3476 (O_3476,N_29904,N_29718);
and UO_3477 (O_3477,N_29758,N_29860);
and UO_3478 (O_3478,N_29723,N_29804);
nor UO_3479 (O_3479,N_29739,N_29764);
nand UO_3480 (O_3480,N_29717,N_29887);
nor UO_3481 (O_3481,N_29833,N_29820);
or UO_3482 (O_3482,N_29710,N_29722);
xnor UO_3483 (O_3483,N_29978,N_29782);
nor UO_3484 (O_3484,N_29983,N_29775);
xor UO_3485 (O_3485,N_29913,N_29715);
or UO_3486 (O_3486,N_29877,N_29778);
and UO_3487 (O_3487,N_29933,N_29906);
and UO_3488 (O_3488,N_29887,N_29821);
xor UO_3489 (O_3489,N_29787,N_29896);
xor UO_3490 (O_3490,N_29924,N_29853);
xnor UO_3491 (O_3491,N_29950,N_29984);
and UO_3492 (O_3492,N_29850,N_29881);
xnor UO_3493 (O_3493,N_29744,N_29786);
nand UO_3494 (O_3494,N_29962,N_29848);
and UO_3495 (O_3495,N_29826,N_29809);
nor UO_3496 (O_3496,N_29844,N_29902);
or UO_3497 (O_3497,N_29752,N_29744);
xnor UO_3498 (O_3498,N_29880,N_29975);
nor UO_3499 (O_3499,N_29766,N_29807);
endmodule