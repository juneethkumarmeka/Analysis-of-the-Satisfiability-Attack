module basic_2500_25000_3000_40_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_1904,In_555);
nand U1 (N_1,In_2297,In_1453);
xor U2 (N_2,In_1825,In_2305);
nand U3 (N_3,In_2346,In_2436);
and U4 (N_4,In_1788,In_2034);
nand U5 (N_5,In_359,In_2475);
or U6 (N_6,In_2342,In_146);
or U7 (N_7,In_2158,In_2263);
xor U8 (N_8,In_1546,In_416);
xor U9 (N_9,In_1879,In_1727);
or U10 (N_10,In_180,In_1387);
and U11 (N_11,In_376,In_1228);
nor U12 (N_12,In_726,In_363);
or U13 (N_13,In_1814,In_2347);
nand U14 (N_14,In_1654,In_640);
xor U15 (N_15,In_1821,In_988);
nand U16 (N_16,In_621,In_1745);
xnor U17 (N_17,In_1327,In_2292);
and U18 (N_18,In_1051,In_868);
nand U19 (N_19,In_2366,In_1310);
and U20 (N_20,In_1160,In_195);
or U21 (N_21,In_1886,In_410);
nand U22 (N_22,In_2382,In_1021);
xnor U23 (N_23,In_685,In_1774);
xnor U24 (N_24,In_684,In_183);
and U25 (N_25,In_1043,In_508);
or U26 (N_26,In_2384,In_2179);
xor U27 (N_27,In_152,In_1783);
nor U28 (N_28,In_1065,In_1437);
or U29 (N_29,In_1036,In_631);
nor U30 (N_30,In_1349,In_2211);
xor U31 (N_31,In_1206,In_979);
nor U32 (N_32,In_2268,In_905);
and U33 (N_33,In_861,In_2145);
nand U34 (N_34,In_1584,In_58);
nor U35 (N_35,In_1278,In_112);
nor U36 (N_36,In_891,In_468);
nand U37 (N_37,In_1171,In_1232);
nand U38 (N_38,In_2444,In_1011);
and U39 (N_39,In_297,In_397);
or U40 (N_40,In_2479,In_423);
or U41 (N_41,In_1279,In_435);
or U42 (N_42,In_617,In_2368);
nor U43 (N_43,In_1460,In_1353);
nor U44 (N_44,In_51,In_762);
xnor U45 (N_45,In_1236,In_386);
xor U46 (N_46,In_249,In_810);
nor U47 (N_47,In_1418,In_1342);
or U48 (N_48,In_501,In_179);
or U49 (N_49,In_2044,In_1448);
xor U50 (N_50,In_831,In_437);
xor U51 (N_51,In_1817,In_924);
or U52 (N_52,In_1970,In_1713);
nand U53 (N_53,In_2089,In_299);
nand U54 (N_54,In_2328,In_2473);
nand U55 (N_55,In_2418,In_191);
and U56 (N_56,In_709,In_1081);
nand U57 (N_57,In_239,In_969);
nor U58 (N_58,In_2279,In_147);
or U59 (N_59,In_2023,In_2293);
and U60 (N_60,In_61,In_68);
and U61 (N_61,In_2282,In_371);
and U62 (N_62,In_2280,In_502);
or U63 (N_63,In_405,In_571);
and U64 (N_64,In_2326,In_288);
xnor U65 (N_65,In_2140,In_1810);
xnor U66 (N_66,In_1633,In_926);
or U67 (N_67,In_1072,In_1020);
and U68 (N_68,In_497,In_851);
nand U69 (N_69,In_674,In_2001);
and U70 (N_70,In_449,In_1956);
and U71 (N_71,In_1594,In_1145);
and U72 (N_72,In_2141,In_521);
xnor U73 (N_73,In_624,In_770);
or U74 (N_74,In_2430,In_1608);
or U75 (N_75,In_190,In_2197);
and U76 (N_76,In_1264,In_226);
and U77 (N_77,In_2483,In_753);
and U78 (N_78,In_1335,In_1990);
or U79 (N_79,In_1307,In_433);
nor U80 (N_80,In_2274,In_379);
and U81 (N_81,In_671,In_138);
nor U82 (N_82,In_1960,In_2083);
or U83 (N_83,In_546,In_1069);
or U84 (N_84,In_1842,In_593);
and U85 (N_85,In_258,In_157);
xor U86 (N_86,In_2148,In_1419);
xor U87 (N_87,In_1019,In_948);
nand U88 (N_88,In_1473,In_400);
and U89 (N_89,In_2101,In_750);
and U90 (N_90,In_2397,In_149);
and U91 (N_91,In_2312,In_1256);
xnor U92 (N_92,In_1626,In_1263);
and U93 (N_93,In_1988,In_2228);
xnor U94 (N_94,In_615,In_1589);
nand U95 (N_95,In_2039,In_2269);
xnor U96 (N_96,In_2106,In_535);
nand U97 (N_97,In_908,In_520);
nand U98 (N_98,In_2370,In_1405);
nand U99 (N_99,In_479,In_2434);
xor U100 (N_100,In_2116,In_610);
nand U101 (N_101,In_185,In_1499);
xnor U102 (N_102,In_121,In_724);
xor U103 (N_103,In_1911,In_2307);
nand U104 (N_104,In_1028,In_395);
or U105 (N_105,In_1314,In_2469);
nand U106 (N_106,In_2287,In_389);
nor U107 (N_107,In_1404,In_616);
and U108 (N_108,In_1916,In_1134);
nor U109 (N_109,In_852,In_1406);
xnor U110 (N_110,In_1846,In_2017);
nor U111 (N_111,In_1106,In_879);
xnor U112 (N_112,In_1482,In_1903);
and U113 (N_113,In_1112,In_2332);
xnor U114 (N_114,In_1966,In_602);
nor U115 (N_115,In_1940,In_1005);
nor U116 (N_116,In_1557,In_528);
nor U117 (N_117,In_773,In_1796);
or U118 (N_118,In_2435,In_1196);
nor U119 (N_119,In_344,In_2353);
nand U120 (N_120,In_1052,In_1304);
xor U121 (N_121,In_1484,In_2308);
nor U122 (N_122,In_1386,In_1086);
xnor U123 (N_123,In_590,In_2363);
and U124 (N_124,In_768,In_1959);
and U125 (N_125,In_767,In_377);
or U126 (N_126,In_2372,In_282);
or U127 (N_127,In_106,In_693);
xnor U128 (N_128,In_369,In_1010);
or U129 (N_129,In_345,In_1420);
and U130 (N_130,In_983,In_1619);
xor U131 (N_131,In_116,In_655);
or U132 (N_132,In_336,In_2086);
and U133 (N_133,In_2240,In_1138);
xor U134 (N_134,In_1739,In_1229);
nand U135 (N_135,In_242,In_2136);
xor U136 (N_136,In_1362,In_2427);
or U137 (N_137,In_622,In_572);
nand U138 (N_138,In_1175,In_2431);
xor U139 (N_139,In_1298,In_2053);
and U140 (N_140,In_2388,In_1276);
xnor U141 (N_141,In_692,In_62);
nor U142 (N_142,In_1850,In_862);
xor U143 (N_143,In_2360,In_273);
nor U144 (N_144,In_1471,In_1492);
and U145 (N_145,In_1260,In_17);
and U146 (N_146,In_1318,In_504);
xor U147 (N_147,In_2210,In_2040);
and U148 (N_148,In_718,In_135);
and U149 (N_149,In_557,In_7);
or U150 (N_150,In_1359,In_1122);
nor U151 (N_151,In_156,In_2213);
nand U152 (N_152,In_579,In_1835);
or U153 (N_153,In_2168,In_1189);
and U154 (N_154,In_764,In_2152);
and U155 (N_155,In_343,In_1408);
and U156 (N_156,In_1672,In_970);
nand U157 (N_157,In_399,In_1500);
or U158 (N_158,In_488,In_1925);
nand U159 (N_159,In_148,In_974);
nor U160 (N_160,In_1429,In_1383);
or U161 (N_161,In_1695,In_13);
xor U162 (N_162,In_2077,In_1870);
xor U163 (N_163,In_2171,In_366);
nor U164 (N_164,In_1114,In_719);
xor U165 (N_165,In_1928,In_517);
and U166 (N_166,In_1169,In_206);
nand U167 (N_167,In_1939,In_2357);
or U168 (N_168,In_442,In_1737);
and U169 (N_169,In_1248,In_1816);
or U170 (N_170,In_2462,In_2003);
nor U171 (N_171,In_943,In_2095);
nand U172 (N_172,In_1528,In_1348);
and U173 (N_173,In_1535,In_1168);
or U174 (N_174,In_954,In_492);
and U175 (N_175,In_1198,In_796);
nor U176 (N_176,In_1214,In_663);
or U177 (N_177,In_1035,In_317);
nand U178 (N_178,In_474,In_1901);
nor U179 (N_179,In_1451,In_1024);
and U180 (N_180,In_1489,In_1213);
xnor U181 (N_181,In_1670,In_1380);
nand U182 (N_182,In_1631,In_141);
and U183 (N_183,In_986,In_686);
and U184 (N_184,In_1937,In_2072);
nor U185 (N_185,In_2195,In_989);
xnor U186 (N_186,In_2409,In_1747);
xor U187 (N_187,In_2183,In_303);
nor U188 (N_188,In_2385,In_2407);
or U189 (N_189,In_1666,In_2371);
nand U190 (N_190,In_165,In_2311);
xnor U191 (N_191,In_478,In_814);
xor U192 (N_192,In_122,In_2439);
nor U193 (N_193,In_1819,In_1332);
and U194 (N_194,In_415,In_743);
nand U195 (N_195,In_1391,In_9);
nor U196 (N_196,In_37,In_1501);
nor U197 (N_197,In_1438,In_248);
and U198 (N_198,In_722,In_1431);
xor U199 (N_199,In_976,In_637);
nor U200 (N_200,In_702,In_2313);
and U201 (N_201,In_1597,In_115);
or U202 (N_202,In_1470,In_688);
and U203 (N_203,In_503,In_930);
nand U204 (N_204,In_1186,In_1055);
and U205 (N_205,In_1881,In_475);
or U206 (N_206,In_964,In_1365);
xor U207 (N_207,In_1250,In_1140);
nand U208 (N_208,In_1709,In_644);
and U209 (N_209,In_319,In_470);
or U210 (N_210,In_199,In_2399);
xor U211 (N_211,In_623,In_421);
nor U212 (N_212,In_1211,In_154);
or U213 (N_213,In_71,In_2383);
xor U214 (N_214,In_1132,In_496);
and U215 (N_215,In_1262,In_1892);
nor U216 (N_216,In_364,In_394);
nand U217 (N_217,In_599,In_654);
nor U218 (N_218,In_2154,In_2122);
nand U219 (N_219,In_2099,In_782);
and U220 (N_220,In_2190,In_279);
and U221 (N_221,In_125,In_963);
or U222 (N_222,In_2309,In_1258);
nor U223 (N_223,In_2425,In_747);
xor U224 (N_224,In_1675,In_2163);
xnor U225 (N_225,In_698,In_283);
and U226 (N_226,In_830,In_204);
and U227 (N_227,In_1797,In_1170);
or U228 (N_228,In_1325,In_537);
and U229 (N_229,In_2013,In_1883);
or U230 (N_230,In_917,In_177);
and U231 (N_231,In_2481,In_1301);
nand U232 (N_232,In_162,In_2005);
and U233 (N_233,In_1822,In_245);
or U234 (N_234,In_1933,In_102);
and U235 (N_235,In_251,In_2193);
xnor U236 (N_236,In_1893,In_1195);
or U237 (N_237,In_716,In_1854);
or U238 (N_238,In_824,In_1203);
and U239 (N_239,In_775,In_2369);
xnor U240 (N_240,In_2432,In_2164);
and U241 (N_241,In_853,In_920);
nor U242 (N_242,In_1372,In_1120);
nor U243 (N_243,In_2079,In_1147);
xnor U244 (N_244,In_613,In_788);
xor U245 (N_245,In_213,In_1234);
nand U246 (N_246,In_63,In_1126);
nor U247 (N_247,In_1309,In_1895);
and U248 (N_248,In_1366,In_357);
and U249 (N_249,In_2488,In_131);
and U250 (N_250,In_1139,In_2087);
nand U251 (N_251,In_1746,In_316);
nor U252 (N_252,In_524,In_2225);
nor U253 (N_253,In_1617,In_666);
nor U254 (N_254,In_1510,In_1936);
xnor U255 (N_255,In_270,In_1433);
xor U256 (N_256,In_1804,In_1566);
or U257 (N_257,In_2146,In_839);
or U258 (N_258,In_1179,In_22);
nand U259 (N_259,In_1423,In_1048);
nand U260 (N_260,In_1071,In_1215);
xnor U261 (N_261,In_1524,In_1678);
nand U262 (N_262,In_257,In_143);
nor U263 (N_263,In_1285,In_605);
xnor U264 (N_264,In_2173,In_2375);
or U265 (N_265,In_2258,In_1770);
and U266 (N_266,In_2172,In_1539);
and U267 (N_267,In_967,In_1743);
and U268 (N_268,In_261,In_913);
nand U269 (N_269,In_8,In_1656);
nor U270 (N_270,In_1523,In_1286);
and U271 (N_271,In_2286,In_2285);
nor U272 (N_272,In_2215,In_1917);
nand U273 (N_273,In_292,In_816);
or U274 (N_274,In_232,In_2075);
nor U275 (N_275,In_2204,In_1981);
xor U276 (N_276,In_2111,In_2440);
and U277 (N_277,In_1582,In_578);
nor U278 (N_278,In_2461,In_1121);
or U279 (N_279,In_123,In_153);
nor U280 (N_280,In_2496,In_25);
and U281 (N_281,In_1089,In_1130);
xor U282 (N_282,In_79,In_929);
and U283 (N_283,In_1664,In_651);
nor U284 (N_284,In_401,In_406);
nand U285 (N_285,In_396,In_2466);
xor U286 (N_286,In_779,In_1467);
nand U287 (N_287,In_255,In_2214);
and U288 (N_288,In_227,In_456);
xnor U289 (N_289,In_2203,In_1426);
and U290 (N_290,In_1908,In_889);
or U291 (N_291,In_438,In_1650);
or U292 (N_292,In_2236,In_1156);
xor U293 (N_293,In_337,In_809);
nor U294 (N_294,In_1809,In_2042);
nor U295 (N_295,In_2008,In_792);
or U296 (N_296,In_2242,In_88);
and U297 (N_297,In_445,In_778);
or U298 (N_298,In_1943,In_2069);
xor U299 (N_299,In_374,In_2247);
nor U300 (N_300,In_1001,In_2120);
nor U301 (N_301,In_43,In_1934);
and U302 (N_302,In_661,In_2177);
nor U303 (N_303,In_2149,In_916);
xor U304 (N_304,In_2390,In_734);
xor U305 (N_305,In_407,In_937);
nor U306 (N_306,In_1843,In_2043);
xor U307 (N_307,In_1100,In_3);
nand U308 (N_308,In_660,In_2422);
xor U309 (N_309,In_2392,In_178);
xor U310 (N_310,In_2337,In_1708);
nand U311 (N_311,In_1000,In_1830);
or U312 (N_312,In_745,In_133);
xnor U313 (N_313,In_720,In_1866);
or U314 (N_314,In_1980,In_1536);
nand U315 (N_315,In_1253,In_1292);
nor U316 (N_316,In_525,In_432);
nor U317 (N_317,In_1085,In_1974);
xor U318 (N_318,In_1720,In_950);
nor U319 (N_319,In_701,In_1345);
xnor U320 (N_320,In_1136,In_1355);
or U321 (N_321,In_538,In_1172);
xor U322 (N_322,In_334,In_1642);
or U323 (N_323,In_1410,In_2374);
nor U324 (N_324,In_931,In_67);
or U325 (N_325,In_2314,In_1519);
and U326 (N_326,In_936,In_2088);
nor U327 (N_327,In_2386,In_2445);
nor U328 (N_328,In_927,In_310);
xnor U329 (N_329,In_1046,In_1158);
nand U330 (N_330,In_2202,In_1671);
nor U331 (N_331,In_1369,In_2150);
xor U332 (N_332,In_2248,In_1515);
nor U333 (N_333,In_1224,In_342);
xnor U334 (N_334,In_834,In_365);
nor U335 (N_335,In_1620,In_844);
nor U336 (N_336,In_2170,In_1151);
nor U337 (N_337,In_275,In_2319);
nor U338 (N_338,In_2381,In_540);
nor U339 (N_339,In_1063,In_928);
nand U340 (N_340,In_1090,In_1984);
xnor U341 (N_341,In_2019,In_733);
nand U342 (N_342,In_139,In_558);
xor U343 (N_343,In_1469,In_1636);
or U344 (N_344,In_55,In_2151);
xor U345 (N_345,In_550,In_163);
xnor U346 (N_346,In_2414,In_188);
and U347 (N_347,In_164,In_269);
nor U348 (N_348,In_2271,In_2379);
and U349 (N_349,In_1047,In_296);
or U350 (N_350,In_2446,In_895);
and U351 (N_351,In_1946,In_1311);
xor U352 (N_352,In_1299,In_1876);
or U353 (N_353,In_2284,In_1768);
or U354 (N_354,In_117,In_975);
nor U355 (N_355,In_1367,In_424);
and U356 (N_356,In_2118,In_1861);
or U357 (N_357,In_495,In_2333);
xor U358 (N_358,In_265,In_1390);
and U359 (N_359,In_1702,In_1697);
xor U360 (N_360,In_980,In_1689);
and U361 (N_361,In_1381,In_527);
nor U362 (N_362,In_471,In_1498);
and U363 (N_363,In_1780,In_1658);
nand U364 (N_364,In_1385,In_874);
and U365 (N_365,In_1765,In_1014);
and U366 (N_366,In_324,In_1906);
nor U367 (N_367,In_2201,In_1623);
xor U368 (N_368,In_901,In_2054);
nor U369 (N_369,In_1176,In_2220);
nor U370 (N_370,In_113,In_1871);
or U371 (N_371,In_114,In_1167);
or U372 (N_372,In_2108,In_1572);
or U373 (N_373,In_990,In_65);
nand U374 (N_374,In_2250,In_1481);
xnor U375 (N_375,In_267,In_783);
xnor U376 (N_376,In_1534,In_1401);
nor U377 (N_377,In_1660,In_1017);
or U378 (N_378,In_2103,In_570);
nand U379 (N_379,In_444,In_1856);
and U380 (N_380,In_910,In_477);
and U381 (N_381,In_327,In_2102);
nor U382 (N_382,In_715,In_2124);
and U383 (N_383,In_1267,In_448);
and U384 (N_384,In_634,In_2223);
nor U385 (N_385,In_2480,In_2254);
nand U386 (N_386,In_29,In_500);
xor U387 (N_387,In_1973,In_2185);
or U388 (N_388,In_2402,In_877);
xnor U389 (N_389,In_1583,In_211);
nor U390 (N_390,In_320,In_1143);
xnor U391 (N_391,In_1696,In_1518);
or U392 (N_392,In_210,In_1596);
and U393 (N_393,In_266,In_315);
or U394 (N_394,In_1360,In_2272);
nand U395 (N_395,In_34,In_2066);
xnor U396 (N_396,In_2014,In_1096);
nand U397 (N_397,In_789,In_2335);
nor U398 (N_398,In_1605,In_1905);
nand U399 (N_399,In_1769,In_2352);
nor U400 (N_400,In_829,In_295);
xor U401 (N_401,In_1744,In_1165);
nand U402 (N_402,In_2090,In_1480);
nand U403 (N_403,In_1986,In_1358);
nor U404 (N_404,In_938,In_104);
and U405 (N_405,In_1789,In_464);
nor U406 (N_406,In_821,In_1734);
and U407 (N_407,In_1845,In_757);
nor U408 (N_408,In_899,In_1514);
nand U409 (N_409,In_291,In_218);
nor U410 (N_410,In_1957,In_1907);
and U411 (N_411,In_1479,In_2464);
nor U412 (N_412,In_1700,In_1926);
nor U413 (N_413,In_2156,In_515);
and U414 (N_414,In_1873,In_2161);
and U415 (N_415,In_679,In_473);
or U416 (N_416,In_1125,In_403);
and U417 (N_417,In_1268,In_1097);
or U418 (N_418,In_285,In_977);
or U419 (N_419,In_2252,In_1627);
nor U420 (N_420,In_739,In_1409);
nand U421 (N_421,In_561,In_289);
and U422 (N_422,In_2249,In_1613);
nor U423 (N_423,In_574,In_428);
nor U424 (N_424,In_194,In_1338);
nand U425 (N_425,In_635,In_33);
nor U426 (N_426,In_1199,In_441);
xnor U427 (N_427,In_2051,In_959);
xor U428 (N_428,In_1287,In_1091);
xnor U429 (N_429,In_375,In_83);
xnor U430 (N_430,In_1251,In_1254);
nor U431 (N_431,In_1651,In_1899);
or U432 (N_432,In_680,In_1512);
nor U433 (N_433,In_2021,In_1975);
nand U434 (N_434,In_801,In_1961);
nor U435 (N_435,In_518,In_2266);
nor U436 (N_436,In_1392,In_669);
nand U437 (N_437,In_689,In_1150);
xor U438 (N_438,In_1162,In_765);
and U439 (N_439,In_708,In_919);
and U440 (N_440,In_695,In_1771);
or U441 (N_441,In_1612,In_922);
or U442 (N_442,In_494,In_1828);
or U443 (N_443,In_595,In_1823);
nor U444 (N_444,In_347,In_47);
nand U445 (N_445,In_1412,In_1979);
or U446 (N_446,In_2007,In_1399);
xnor U447 (N_447,In_507,In_2270);
or U448 (N_448,In_559,In_124);
or U449 (N_449,In_1885,In_1108);
nand U450 (N_450,In_1204,In_166);
and U451 (N_451,In_1424,In_754);
and U452 (N_452,In_1067,In_81);
nor U453 (N_453,In_549,In_1773);
and U454 (N_454,In_781,In_2472);
xnor U455 (N_455,In_1305,In_1131);
xnor U456 (N_456,In_1354,In_890);
nand U457 (N_457,In_1949,In_1398);
nor U458 (N_458,In_2234,In_1416);
and U459 (N_459,In_32,In_1245);
and U460 (N_460,In_2405,In_547);
and U461 (N_461,In_1261,In_2377);
xnor U462 (N_462,In_1351,In_385);
nor U463 (N_463,In_1294,In_2091);
nand U464 (N_464,In_828,In_1303);
or U465 (N_465,In_2343,In_1124);
nand U466 (N_466,In_690,In_128);
nor U467 (N_467,In_706,In_2294);
nor U468 (N_468,In_1364,In_2437);
and U469 (N_469,In_85,In_2094);
xnor U470 (N_470,In_431,In_961);
xnor U471 (N_471,In_216,In_545);
nor U472 (N_472,In_27,In_996);
xor U473 (N_473,In_1686,In_66);
nand U474 (N_474,In_2394,In_56);
nor U475 (N_475,In_482,In_2334);
nor U476 (N_476,In_126,In_1860);
xnor U477 (N_477,In_1606,In_2174);
nand U478 (N_478,In_513,In_221);
or U479 (N_479,In_78,In_2303);
nor U480 (N_480,In_656,In_462);
or U481 (N_481,In_417,In_888);
or U482 (N_482,In_75,In_2486);
nand U483 (N_483,In_531,In_2081);
nor U484 (N_484,In_212,In_1368);
nor U485 (N_485,In_923,In_667);
and U486 (N_486,In_949,In_944);
nand U487 (N_487,In_169,In_1266);
xnor U488 (N_488,In_703,In_848);
nor U489 (N_489,In_1802,In_1087);
and U490 (N_490,In_268,In_1187);
nand U491 (N_491,In_2046,In_873);
or U492 (N_492,In_1182,In_1867);
and U493 (N_493,In_921,In_2497);
or U494 (N_494,In_1503,In_457);
or U495 (N_495,In_962,In_170);
or U496 (N_496,In_639,In_958);
or U497 (N_497,In_1761,In_2045);
xnor U498 (N_498,In_2126,In_800);
xor U499 (N_499,In_568,In_677);
xor U500 (N_500,In_1756,In_2096);
or U501 (N_501,In_1025,In_618);
xor U502 (N_502,In_1238,In_804);
and U503 (N_503,In_742,In_150);
nor U504 (N_504,In_1989,In_451);
and U505 (N_505,In_90,In_175);
nor U506 (N_506,In_1750,In_1992);
or U507 (N_507,In_1598,In_567);
and U508 (N_508,In_340,In_1505);
and U509 (N_509,In_682,In_484);
nor U510 (N_510,In_2485,In_201);
or U511 (N_511,In_1283,In_1791);
xor U512 (N_512,In_493,In_1754);
nand U513 (N_513,In_1552,In_2018);
xor U514 (N_514,In_2457,In_1897);
and U515 (N_515,In_1948,In_2356);
xnor U516 (N_516,In_1983,In_607);
and U517 (N_517,In_93,In_611);
or U518 (N_518,In_2376,In_1545);
or U519 (N_519,In_2028,In_1184);
nand U520 (N_520,In_1356,In_2246);
xnor U521 (N_521,In_362,In_2135);
nand U522 (N_522,In_1591,In_353);
nand U523 (N_523,In_2325,In_1246);
nor U524 (N_524,In_1725,In_903);
nor U525 (N_525,In_82,In_57);
nor U526 (N_526,In_1760,In_746);
nor U527 (N_527,In_1513,In_628);
or U528 (N_528,In_1425,In_2238);
and U529 (N_529,In_1079,In_1938);
or U530 (N_530,In_1882,In_2256);
nand U531 (N_531,In_1622,In_2459);
or U532 (N_532,In_1083,In_1994);
xnor U533 (N_533,In_803,In_1319);
or U534 (N_534,In_575,In_1472);
nand U535 (N_535,In_2059,In_653);
and U536 (N_536,In_1075,In_192);
xnor U537 (N_537,In_314,In_1726);
and U538 (N_538,In_642,In_1630);
and U539 (N_539,In_1890,In_243);
and U540 (N_540,In_1235,In_1565);
and U541 (N_541,In_1221,In_1443);
and U542 (N_542,In_312,In_1447);
nor U543 (N_543,In_1703,In_1243);
and U544 (N_544,In_346,In_1653);
or U545 (N_545,In_1914,In_993);
or U546 (N_546,In_1554,In_2109);
nor U547 (N_547,In_1296,In_1084);
and U548 (N_548,In_2365,In_939);
nor U549 (N_549,In_1508,In_1680);
or U550 (N_550,In_1297,In_459);
nor U551 (N_551,In_1638,In_1913);
nor U552 (N_552,In_2037,In_1643);
nor U553 (N_553,In_1998,In_1615);
or U554 (N_554,In_832,In_902);
or U555 (N_555,In_912,In_1909);
nand U556 (N_556,In_736,In_1935);
and U557 (N_557,In_1450,In_1915);
nand U558 (N_558,In_2216,In_349);
or U559 (N_559,In_2160,In_2463);
xnor U560 (N_560,In_358,In_325);
nand U561 (N_561,In_355,In_2056);
nand U562 (N_562,In_1334,In_1436);
xnor U563 (N_563,In_2092,In_42);
nor U564 (N_564,In_730,In_11);
nor U565 (N_565,In_2306,In_1592);
or U566 (N_566,In_2080,In_1040);
nor U567 (N_567,In_887,In_91);
nand U568 (N_568,In_1293,In_38);
and U569 (N_569,In_1076,In_509);
and U570 (N_570,In_1985,In_2350);
xor U571 (N_571,In_40,In_39);
and U572 (N_572,In_231,In_46);
xnor U573 (N_573,In_633,In_18);
and U574 (N_574,In_54,In_196);
xor U575 (N_575,In_1833,In_1377);
nand U576 (N_576,In_1661,In_1153);
and U577 (N_577,In_1969,In_73);
and U578 (N_578,In_1838,In_1060);
or U579 (N_579,In_2295,In_1764);
or U580 (N_580,In_869,In_994);
or U581 (N_581,In_305,In_499);
nand U582 (N_582,In_110,In_2192);
or U583 (N_583,In_1857,In_544);
and U584 (N_584,In_1417,In_1029);
nor U585 (N_585,In_907,In_1078);
nor U586 (N_586,In_1865,In_1647);
xor U587 (N_587,In_2487,In_2396);
and U588 (N_588,In_2331,In_2029);
or U589 (N_589,In_418,In_696);
nor U590 (N_590,In_512,In_592);
nor U591 (N_591,In_1240,In_1101);
nor U592 (N_592,In_352,In_1152);
or U593 (N_593,In_897,In_2257);
and U594 (N_594,In_2082,In_2499);
or U595 (N_595,In_1724,In_2355);
and U596 (N_596,In_1009,In_807);
and U597 (N_597,In_2318,In_404);
xor U598 (N_598,In_1588,In_608);
nand U599 (N_599,In_2323,In_193);
and U600 (N_600,In_254,In_2212);
xnor U601 (N_601,In_1149,In_823);
xor U602 (N_602,In_1226,In_250);
xnor U603 (N_603,In_2208,In_652);
nor U604 (N_604,In_1687,In_1103);
xnor U605 (N_605,In_1963,In_1123);
nor U606 (N_606,In_1662,In_1230);
or U607 (N_607,In_1434,In_2221);
xnor U608 (N_608,In_1851,In_1070);
nor U609 (N_609,In_1640,In_712);
nor U610 (N_610,In_1648,In_612);
xor U611 (N_611,In_960,In_1690);
nand U612 (N_612,In_1506,In_2226);
xnor U613 (N_613,In_1782,In_260);
xnor U614 (N_614,In_1058,In_1601);
xnor U615 (N_615,In_1414,In_217);
nand U616 (N_616,In_1407,In_1316);
nor U617 (N_617,In_259,In_553);
nand U618 (N_618,In_1558,In_2478);
or U619 (N_619,In_1275,In_1655);
or U620 (N_620,In_168,In_2327);
nand U621 (N_621,In_414,In_2442);
xnor U622 (N_622,In_333,In_92);
xor U623 (N_623,In_749,In_80);
xor U624 (N_624,In_202,In_2489);
or U625 (N_625,In_543,In_665);
xnor U626 (N_626,N_575,N_492);
and U627 (N_627,In_1629,In_1529);
xor U628 (N_628,In_2358,N_164);
and U629 (N_629,In_2239,In_45);
nor U630 (N_630,In_1559,In_108);
and U631 (N_631,N_567,In_2498);
or U632 (N_632,N_499,In_1787);
or U633 (N_633,In_1273,N_163);
nand U634 (N_634,N_420,In_1556);
xor U635 (N_635,In_1766,In_2467);
nand U636 (N_636,In_815,N_204);
nand U637 (N_637,In_384,In_393);
xor U638 (N_638,In_409,In_1632);
xor U639 (N_639,In_1201,In_956);
nor U640 (N_640,In_2367,N_353);
nand U641 (N_641,N_476,N_45);
or U642 (N_642,N_230,In_893);
xnor U643 (N_643,N_558,In_1497);
or U644 (N_644,In_2074,N_310);
xnor U645 (N_645,In_2,In_1952);
xnor U646 (N_646,N_159,In_1485);
or U647 (N_647,In_1891,In_228);
and U648 (N_648,In_1637,In_134);
nand U649 (N_649,In_284,N_79);
nor U650 (N_650,In_1008,In_446);
nand U651 (N_651,N_516,In_1698);
nor U652 (N_652,N_463,N_308);
nor U653 (N_653,In_1894,N_324);
and U654 (N_654,In_530,In_576);
and U655 (N_655,N_211,N_252);
nand U656 (N_656,In_1784,N_238);
nand U657 (N_657,N_202,In_2495);
and U658 (N_658,N_98,N_113);
or U659 (N_659,N_43,N_320);
or U660 (N_660,In_1731,N_377);
xor U661 (N_661,N_446,In_1762);
nand U662 (N_662,N_604,In_1714);
nor U663 (N_663,N_70,N_160);
xor U664 (N_664,In_307,In_886);
xor U665 (N_665,N_534,In_1553);
nor U666 (N_666,In_563,N_341);
xor U667 (N_667,N_148,In_588);
nor U668 (N_668,In_1549,In_426);
nand U669 (N_669,N_169,In_1717);
and U670 (N_670,N_17,In_1066);
xor U671 (N_671,In_48,N_187);
or U672 (N_672,In_2474,In_2449);
xor U673 (N_673,In_1781,N_245);
nand U674 (N_674,In_1954,N_24);
xor U675 (N_675,In_1255,In_1525);
and U676 (N_676,N_454,In_2020);
nor U677 (N_677,In_797,In_1921);
nor U678 (N_678,In_609,N_360);
and U679 (N_679,In_1544,N_125);
nor U680 (N_680,In_2421,In_856);
xor U681 (N_681,In_1600,In_577);
xor U682 (N_682,In_529,In_1271);
or U683 (N_683,In_1971,N_514);
and U684 (N_684,N_331,In_2006);
and U685 (N_685,In_802,In_1965);
nand U686 (N_686,N_158,In_72);
nand U687 (N_687,N_88,In_1329);
or U688 (N_688,N_3,In_472);
and U689 (N_689,N_440,In_668);
and U690 (N_690,In_1045,In_1449);
nand U691 (N_691,N_594,N_268);
xnor U692 (N_692,In_704,In_12);
xnor U693 (N_693,N_546,In_2301);
nor U694 (N_694,In_2322,In_833);
or U695 (N_695,In_1037,N_123);
or U696 (N_696,N_497,N_274);
nor U697 (N_697,In_274,In_522);
nand U698 (N_698,In_1688,In_19);
xor U699 (N_699,In_1628,In_1639);
xnor U700 (N_700,N_387,In_1900);
or U701 (N_701,In_995,In_35);
and U702 (N_702,N_355,In_200);
nand U703 (N_703,In_1738,In_2477);
nand U704 (N_704,In_822,In_2235);
xnor U705 (N_705,In_2471,In_738);
and U706 (N_706,In_1073,In_1621);
or U707 (N_707,In_1379,In_717);
nand U708 (N_708,N_299,In_2143);
or U709 (N_709,N_343,In_795);
nand U710 (N_710,In_1459,In_313);
and U711 (N_711,In_843,In_915);
and U712 (N_712,In_137,In_1042);
xor U713 (N_713,N_115,In_1324);
nor U714 (N_714,N_478,In_1452);
nor U715 (N_715,In_2338,In_918);
nand U716 (N_716,In_2416,In_1942);
and U717 (N_717,In_294,In_1241);
nand U718 (N_718,N_347,In_650);
nor U719 (N_719,N_176,In_370);
nand U720 (N_720,In_2070,N_263);
nand U721 (N_721,In_691,N_40);
or U722 (N_722,N_325,In_984);
nand U723 (N_723,In_229,In_1454);
nor U724 (N_724,N_501,In_1002);
and U725 (N_725,In_1652,In_287);
or U726 (N_726,In_1044,In_2100);
or U727 (N_727,In_900,In_1464);
nand U728 (N_728,In_301,N_445);
nor U729 (N_729,In_1635,In_1701);
xor U730 (N_730,In_1968,In_641);
xor U731 (N_731,In_882,In_2482);
nor U732 (N_732,In_699,In_2196);
xnor U733 (N_733,In_2310,In_997);
and U734 (N_734,In_1223,In_672);
and U735 (N_735,N_511,N_46);
or U736 (N_736,In_1030,In_1210);
and U737 (N_737,N_303,In_554);
nor U738 (N_738,N_216,In_1333);
nand U739 (N_739,In_790,N_412);
xnor U740 (N_740,N_578,N_498);
and U741 (N_741,In_2026,N_536);
nand U742 (N_742,In_587,In_1411);
nand U743 (N_743,In_1728,In_2373);
or U744 (N_744,In_1749,In_2232);
and U745 (N_745,N_162,In_2451);
or U746 (N_746,In_772,N_590);
and U747 (N_747,N_337,In_187);
nand U748 (N_748,In_318,In_2494);
nor U749 (N_749,N_471,In_581);
xor U750 (N_750,In_220,In_322);
nand U751 (N_751,In_1679,In_1093);
xor U752 (N_752,N_488,N_402);
nor U753 (N_753,In_1190,In_5);
nand U754 (N_754,In_1208,In_721);
nor U755 (N_755,In_619,In_1603);
nand U756 (N_756,N_539,In_1562);
or U757 (N_757,N_515,In_1922);
and U758 (N_758,N_103,In_565);
or U759 (N_759,N_519,In_1964);
or U760 (N_760,In_429,In_367);
and U761 (N_761,N_393,In_247);
or U762 (N_762,In_311,In_1183);
nand U763 (N_763,In_413,In_103);
and U764 (N_764,In_1099,In_2107);
and U765 (N_765,In_1840,In_2491);
nand U766 (N_766,N_205,N_396);
or U767 (N_767,N_80,N_434);
nand U768 (N_768,N_455,In_2167);
nor U769 (N_769,N_431,In_1586);
nor U770 (N_770,In_1803,In_1997);
xor U771 (N_771,In_26,In_1291);
or U772 (N_772,In_514,N_260);
and U773 (N_773,In_1494,In_2490);
or U774 (N_774,In_2267,In_2476);
nand U775 (N_775,In_158,In_2316);
nor U776 (N_776,In_1347,N_87);
or U777 (N_777,In_1712,N_117);
nand U778 (N_778,In_1777,In_1027);
nand U779 (N_779,In_562,In_1242);
xnor U780 (N_780,In_2128,N_623);
xnor U781 (N_781,N_99,In_1222);
or U782 (N_782,In_573,In_647);
xnor U783 (N_783,In_766,In_2063);
nor U784 (N_784,N_266,In_2378);
nand U785 (N_785,In_1474,In_52);
or U786 (N_786,In_569,In_1733);
nor U787 (N_787,N_452,In_884);
and U788 (N_788,In_491,In_1736);
xnor U789 (N_789,In_1445,In_326);
nand U790 (N_790,N_109,In_1476);
xnor U791 (N_791,In_1312,In_203);
and U792 (N_792,N_541,N_551);
nor U793 (N_793,In_145,In_1995);
nand U794 (N_794,N_180,In_453);
xnor U795 (N_795,N_562,In_664);
nand U796 (N_796,In_2058,N_36);
nor U797 (N_797,In_167,In_1799);
and U798 (N_798,In_460,In_28);
nand U799 (N_799,N_240,N_329);
nand U800 (N_800,In_1018,In_1269);
or U801 (N_801,In_2057,In_1013);
xnor U802 (N_802,N_411,In_1945);
nor U803 (N_803,In_24,In_1699);
nand U804 (N_804,In_1382,In_2255);
nor U805 (N_805,In_1509,In_1321);
or U806 (N_806,In_2067,In_1958);
and U807 (N_807,In_1326,In_985);
xor U808 (N_808,In_234,In_252);
xor U809 (N_809,In_1538,In_1763);
nand U810 (N_810,N_466,In_1927);
xnor U811 (N_811,N_383,In_1676);
nor U812 (N_812,In_859,In_2153);
nor U813 (N_813,In_1146,In_818);
nor U814 (N_814,In_171,In_2180);
and U815 (N_815,N_177,In_981);
nor U816 (N_816,In_186,In_1463);
xor U817 (N_817,N_91,In_878);
or U818 (N_818,N_249,In_1322);
or U819 (N_819,In_812,N_119);
xnor U820 (N_820,In_871,In_785);
or U821 (N_821,N_624,In_373);
or U822 (N_822,In_398,In_434);
xnor U823 (N_823,In_854,In_2078);
nor U824 (N_824,N_469,N_610);
and U825 (N_825,In_1721,In_2391);
and U826 (N_826,In_744,N_365);
xnor U827 (N_827,N_582,N_602);
nand U828 (N_828,In_2304,In_381);
nor U829 (N_829,N_357,In_2032);
nor U830 (N_830,In_1691,N_267);
nor U831 (N_831,In_205,In_1795);
or U832 (N_832,N_132,N_116);
xnor U833 (N_833,In_1793,In_1173);
or U834 (N_834,In_2320,In_1350);
xnor U835 (N_835,In_2068,In_1953);
or U836 (N_836,In_2400,In_1006);
and U837 (N_837,In_1502,In_941);
xor U838 (N_838,N_285,N_384);
or U839 (N_839,In_487,N_592);
nor U840 (N_840,In_2395,In_636);
xnor U841 (N_841,In_1004,In_2419);
xnor U842 (N_842,In_2061,In_1868);
and U843 (N_843,N_559,In_1920);
xor U844 (N_844,In_1581,In_97);
and U845 (N_845,N_231,In_1288);
nand U846 (N_846,N_447,In_1880);
nor U847 (N_847,In_2138,N_203);
nor U848 (N_848,N_53,In_629);
and U849 (N_849,In_2341,In_1339);
xor U850 (N_850,In_978,In_176);
nand U851 (N_851,In_486,In_1315);
nand U852 (N_852,In_539,N_618);
nor U853 (N_853,In_2336,In_41);
xnor U854 (N_854,In_1864,In_2380);
nor U855 (N_855,In_2025,In_159);
nor U856 (N_856,In_1910,In_2302);
xnor U857 (N_857,In_2155,N_246);
nor U858 (N_858,N_529,N_376);
xor U859 (N_859,In_1641,N_588);
xnor U860 (N_860,In_2404,In_2441);
xor U861 (N_861,In_1681,In_430);
and U862 (N_862,In_1488,In_2176);
and U863 (N_863,N_547,In_1003);
xor U864 (N_864,N_151,In_700);
and U865 (N_865,In_1962,N_195);
nand U866 (N_866,N_2,In_1328);
or U867 (N_867,In_402,In_2052);
xor U868 (N_868,In_489,In_1604);
nor U869 (N_869,In_1659,N_253);
or U870 (N_870,In_1128,N_467);
or U871 (N_871,In_1039,In_2413);
and U872 (N_872,In_1374,N_112);
and U873 (N_873,In_1602,N_143);
nand U874 (N_874,N_100,N_483);
xor U875 (N_875,In_1778,In_447);
nor U876 (N_876,In_1142,In_1343);
nor U877 (N_877,N_366,N_198);
and U878 (N_878,In_2401,In_1668);
xor U879 (N_879,N_401,N_316);
nand U880 (N_880,N_1,N_102);
nor U881 (N_881,N_419,In_1154);
nand U882 (N_882,In_1402,In_799);
nand U883 (N_883,In_293,N_385);
or U884 (N_884,In_1225,N_97);
or U885 (N_885,In_1759,In_1872);
and U886 (N_886,In_1023,In_876);
nor U887 (N_887,N_149,In_214);
nand U888 (N_888,N_287,In_2038);
and U889 (N_889,In_1863,In_1813);
xor U890 (N_890,In_1444,In_390);
and U891 (N_891,N_146,In_2041);
xnor U892 (N_892,In_127,In_1155);
or U893 (N_893,In_626,N_386);
nand U894 (N_894,N_429,In_589);
nor U895 (N_895,N_206,In_1996);
xnor U896 (N_896,N_405,In_583);
xnor U897 (N_897,In_1576,In_161);
or U898 (N_898,N_229,N_281);
or U899 (N_899,N_83,In_2010);
xnor U900 (N_900,In_1239,In_526);
and U901 (N_901,In_662,In_933);
and U902 (N_902,N_225,In_1839);
or U903 (N_903,N_38,In_209);
nor U904 (N_904,In_15,In_2283);
nand U905 (N_905,N_493,In_233);
xnor U906 (N_906,In_2219,In_2073);
or U907 (N_907,In_1707,In_263);
nand U908 (N_908,N_407,In_1207);
or U909 (N_909,N_453,In_1133);
nand U910 (N_910,In_1693,In_173);
or U911 (N_911,N_389,N_334);
nand U912 (N_912,In_1259,In_1849);
xor U913 (N_913,N_133,In_1477);
nor U914 (N_914,In_1188,In_1977);
xor U915 (N_915,In_2460,N_394);
xor U916 (N_916,N_489,N_537);
and U917 (N_917,N_156,In_761);
nor U918 (N_918,In_53,In_69);
or U919 (N_919,In_348,N_52);
nor U920 (N_920,In_857,In_1775);
and U921 (N_921,In_1041,In_368);
xnor U922 (N_922,In_1233,N_577);
and U923 (N_923,N_239,N_185);
nor U924 (N_924,N_472,N_166);
xnor U925 (N_925,In_1456,In_272);
xor U926 (N_926,N_586,In_1533);
nor U927 (N_927,In_351,In_673);
and U928 (N_928,In_511,In_2281);
nor U929 (N_929,In_329,N_542);
and U930 (N_930,In_1102,In_281);
and U931 (N_931,In_2470,In_2002);
nand U932 (N_932,N_378,In_1137);
and U933 (N_933,In_1094,N_256);
nor U934 (N_934,N_73,In_1373);
xnor U935 (N_935,In_1331,N_410);
or U936 (N_936,In_264,In_675);
or U937 (N_937,N_349,In_1607);
xnor U938 (N_938,In_276,N_291);
and U939 (N_939,In_836,N_556);
or U940 (N_940,N_600,In_1991);
and U941 (N_941,In_262,N_172);
or U942 (N_942,N_0,In_476);
or U943 (N_943,In_1077,In_1806);
nor U944 (N_944,In_1896,N_505);
nor U945 (N_945,N_186,N_278);
or U946 (N_946,N_335,In_1578);
xnor U947 (N_947,In_1166,In_711);
and U948 (N_948,In_2340,In_942);
nor U949 (N_949,N_363,In_1413);
or U950 (N_950,N_94,N_219);
and U951 (N_951,N_5,In_332);
nand U952 (N_952,N_155,N_527);
and U953 (N_953,In_973,In_1466);
nor U954 (N_954,In_1435,In_1375);
and U955 (N_955,N_352,In_208);
xor U956 (N_956,In_1573,In_1859);
or U957 (N_957,In_534,In_1742);
and U958 (N_958,In_99,N_120);
and U959 (N_959,In_1370,In_1371);
and U960 (N_960,In_44,In_1683);
or U961 (N_961,In_1716,In_1520);
or U962 (N_962,In_2387,In_59);
or U963 (N_963,In_298,In_36);
nor U964 (N_964,In_951,In_2132);
nor U965 (N_965,In_911,N_364);
xor U966 (N_966,N_438,In_450);
or U967 (N_967,In_1824,N_190);
xnor U968 (N_968,In_731,In_2110);
xor U969 (N_969,N_222,In_542);
nand U970 (N_970,In_174,In_649);
xor U971 (N_971,In_817,N_171);
nor U972 (N_972,N_328,N_545);
and U973 (N_973,In_1415,In_331);
and U974 (N_974,In_2429,In_21);
nor U975 (N_975,N_241,In_1107);
nand U976 (N_976,In_2093,In_286);
nor U977 (N_977,N_284,In_2104);
or U978 (N_978,In_872,In_748);
nor U979 (N_979,In_1669,N_197);
and U980 (N_980,N_68,N_479);
xnor U981 (N_981,In_2458,In_241);
nand U982 (N_982,In_1530,In_1022);
nor U983 (N_983,In_935,In_278);
xnor U984 (N_984,In_787,In_0);
nand U985 (N_985,In_1918,In_1098);
or U986 (N_986,N_212,In_551);
or U987 (N_987,In_1531,In_306);
and U988 (N_988,N_425,In_1858);
xor U989 (N_989,N_242,N_276);
and U990 (N_990,N_596,In_2229);
or U991 (N_991,In_105,In_945);
nand U992 (N_992,N_354,In_2137);
and U993 (N_993,N_39,In_759);
nand U994 (N_994,In_244,N_482);
nand U995 (N_995,N_259,In_940);
xnor U996 (N_996,In_2121,In_1599);
nor U997 (N_997,In_966,In_1685);
nand U998 (N_998,In_1068,In_1191);
xnor U999 (N_999,In_2181,N_75);
xnor U1000 (N_1000,In_223,In_2484);
or U1001 (N_1001,In_566,In_1847);
nor U1002 (N_1002,In_465,N_236);
or U1003 (N_1003,In_794,N_50);
nand U1004 (N_1004,In_222,In_600);
xnor U1005 (N_1005,In_2349,N_369);
nor U1006 (N_1006,In_2237,In_335);
nor U1007 (N_1007,In_2450,N_29);
nand U1008 (N_1008,In_2127,In_1317);
or U1009 (N_1009,In_934,In_1252);
or U1010 (N_1010,In_1088,In_2217);
nand U1011 (N_1011,In_1618,N_404);
nand U1012 (N_1012,In_1430,In_971);
xnor U1013 (N_1013,In_2423,In_598);
and U1014 (N_1014,In_2024,N_174);
xor U1015 (N_1015,N_290,N_548);
nor U1016 (N_1016,In_2415,N_196);
nor U1017 (N_1017,In_614,N_318);
xor U1018 (N_1018,In_2035,N_114);
or U1019 (N_1019,In_627,N_294);
and U1020 (N_1020,In_1832,N_168);
and U1021 (N_1021,N_33,In_728);
or U1022 (N_1022,N_430,In_533);
or U1023 (N_1023,N_327,In_1490);
or U1024 (N_1024,In_1290,In_290);
and U1025 (N_1025,In_1852,In_1007);
xnor U1026 (N_1026,In_1164,In_1446);
or U1027 (N_1027,In_64,In_892);
and U1028 (N_1028,In_670,N_314);
or U1029 (N_1029,N_561,N_579);
or U1030 (N_1030,In_308,In_760);
or U1031 (N_1031,N_8,N_258);
xor U1032 (N_1032,N_544,N_111);
nand U1033 (N_1033,In_2277,In_2159);
xor U1034 (N_1034,N_477,In_60);
nand U1035 (N_1035,In_838,In_1080);
nand U1036 (N_1036,In_2452,In_302);
xnor U1037 (N_1037,In_2065,In_2206);
or U1038 (N_1038,In_1521,N_587);
nand U1039 (N_1039,In_1212,In_280);
nand U1040 (N_1040,In_1673,In_865);
nand U1041 (N_1041,In_1987,In_532);
nand U1042 (N_1042,N_603,N_459);
or U1043 (N_1043,In_1478,In_658);
and U1044 (N_1044,N_591,In_1468);
nor U1045 (N_1045,N_126,In_860);
and U1046 (N_1046,In_2191,In_1898);
nand U1047 (N_1047,N_210,In_339);
nand U1048 (N_1048,In_2433,In_235);
nand U1049 (N_1049,N_153,N_484);
nor U1050 (N_1050,N_20,In_1624);
nand U1051 (N_1051,In_2016,In_372);
and U1052 (N_1052,N_509,In_1730);
xor U1053 (N_1053,In_1400,In_1116);
or U1054 (N_1054,In_763,In_1735);
xor U1055 (N_1055,N_63,N_475);
nor U1056 (N_1056,In_1220,In_1855);
nand U1057 (N_1057,N_423,N_295);
or U1058 (N_1058,In_1439,In_1507);
nand U1059 (N_1059,N_315,In_480);
or U1060 (N_1060,In_436,N_279);
or U1061 (N_1061,In_1197,In_84);
nor U1062 (N_1062,In_2493,In_1848);
xor U1063 (N_1063,In_1200,N_442);
and U1064 (N_1064,N_494,N_14);
nand U1065 (N_1065,In_2131,In_1772);
xor U1066 (N_1066,In_808,N_332);
nor U1067 (N_1067,In_1313,In_1826);
xor U1068 (N_1068,In_2389,In_1104);
nor U1069 (N_1069,N_76,In_1740);
xnor U1070 (N_1070,In_2315,N_262);
nor U1071 (N_1071,In_1571,In_2299);
xor U1072 (N_1072,N_15,In_1192);
nand U1073 (N_1073,N_304,N_234);
or U1074 (N_1074,N_311,N_191);
or U1075 (N_1075,In_707,In_2406);
nand U1076 (N_1076,In_1185,In_2076);
nor U1077 (N_1077,In_1853,In_443);
xor U1078 (N_1078,N_69,In_1395);
and U1079 (N_1079,In_1976,In_1547);
and U1080 (N_1080,N_508,In_2443);
xor U1081 (N_1081,N_408,In_1034);
xor U1082 (N_1082,In_2009,In_74);
and U1083 (N_1083,In_2408,In_1219);
nor U1084 (N_1084,N_565,N_271);
and U1085 (N_1085,In_2114,N_48);
xor U1086 (N_1086,In_237,In_1888);
or U1087 (N_1087,In_354,In_740);
nand U1088 (N_1088,In_972,In_189);
nand U1089 (N_1089,N_533,N_131);
nor U1090 (N_1090,In_1491,In_1644);
xnor U1091 (N_1091,In_1144,N_382);
or U1092 (N_1092,In_1805,In_253);
nand U1093 (N_1093,N_221,In_4);
xnor U1094 (N_1094,In_1827,In_678);
nand U1095 (N_1095,N_495,N_368);
xor U1096 (N_1096,In_20,In_2162);
and U1097 (N_1097,In_2182,In_914);
or U1098 (N_1098,N_62,In_2027);
nor U1099 (N_1099,In_1931,N_549);
xor U1100 (N_1100,N_283,N_173);
nor U1101 (N_1101,In_1032,In_898);
nor U1102 (N_1102,In_1493,N_86);
nand U1103 (N_1103,In_240,In_2224);
or U1104 (N_1104,N_179,N_250);
or U1105 (N_1105,In_2264,In_1569);
nand U1106 (N_1106,In_1595,N_480);
nand U1107 (N_1107,In_1320,In_1148);
and U1108 (N_1108,In_2428,N_107);
or U1109 (N_1109,In_1336,In_2133);
nand U1110 (N_1110,N_273,N_362);
xnor U1111 (N_1111,In_49,N_457);
nor U1112 (N_1112,In_338,In_1403);
and U1113 (N_1113,N_520,In_1831);
xnor U1114 (N_1114,In_1902,In_548);
nor U1115 (N_1115,N_130,In_2227);
nor U1116 (N_1116,In_1455,In_1247);
nand U1117 (N_1117,In_132,In_1527);
or U1118 (N_1118,In_732,N_21);
xor U1119 (N_1119,N_35,In_2084);
xor U1120 (N_1120,N_142,N_323);
nand U1121 (N_1121,In_1344,In_867);
or U1122 (N_1122,N_400,In_516);
or U1123 (N_1123,In_1462,In_946);
xor U1124 (N_1124,In_2112,In_1786);
and U1125 (N_1125,N_12,N_108);
and U1126 (N_1126,In_94,In_23);
nand U1127 (N_1127,In_2230,In_2398);
and U1128 (N_1128,In_1776,In_2420);
nand U1129 (N_1129,N_140,In_1428);
and U1130 (N_1130,In_1932,In_2207);
and U1131 (N_1131,N_289,N_348);
or U1132 (N_1132,In_111,In_2411);
and U1133 (N_1133,In_741,N_433);
nor U1134 (N_1134,In_1947,In_1205);
nor U1135 (N_1135,In_300,In_2119);
nor U1136 (N_1136,In_2244,N_518);
and U1137 (N_1137,In_350,N_583);
nor U1138 (N_1138,In_1161,N_614);
xnor U1139 (N_1139,In_1792,N_25);
or U1140 (N_1140,In_2447,In_771);
or U1141 (N_1141,In_826,In_422);
xnor U1142 (N_1142,In_1389,N_601);
or U1143 (N_1143,N_233,In_50);
and U1144 (N_1144,N_522,In_2033);
or U1145 (N_1145,In_1216,In_552);
or U1146 (N_1146,In_2273,In_1575);
and U1147 (N_1147,In_604,In_391);
and U1148 (N_1148,In_2157,In_2260);
nand U1149 (N_1149,In_786,In_1563);
or U1150 (N_1150,N_557,In_1929);
or U1151 (N_1151,In_309,In_1495);
nor U1152 (N_1152,In_76,In_2115);
nor U1153 (N_1153,N_312,In_1614);
and U1154 (N_1154,N_57,In_2134);
or U1155 (N_1155,In_723,In_687);
nand U1156 (N_1156,In_277,In_2187);
nor U1157 (N_1157,N_64,In_1231);
nand U1158 (N_1158,In_1684,In_835);
nor U1159 (N_1159,N_322,In_380);
nand U1160 (N_1160,In_755,In_107);
xnor U1161 (N_1161,N_566,In_1141);
xnor U1162 (N_1162,In_2465,In_356);
nor U1163 (N_1163,In_992,In_142);
and U1164 (N_1164,In_523,N_622);
xnor U1165 (N_1165,In_452,In_1016);
and U1166 (N_1166,In_1517,In_1993);
and U1167 (N_1167,In_2454,N_612);
or U1168 (N_1168,N_374,N_451);
and U1169 (N_1169,N_563,In_378);
or U1170 (N_1170,N_532,In_1800);
nand U1171 (N_1171,In_1257,N_31);
nand U1172 (N_1172,In_1378,In_466);
or U1173 (N_1173,N_456,In_2178);
nand U1174 (N_1174,In_955,N_61);
nor U1175 (N_1175,In_1543,In_820);
xor U1176 (N_1176,In_2117,In_1585);
xnor U1177 (N_1177,In_1059,In_1376);
or U1178 (N_1178,In_1590,In_1062);
nor U1179 (N_1179,N_6,In_1394);
xor U1180 (N_1180,In_705,N_4);
nor U1181 (N_1181,N_358,In_1300);
or U1182 (N_1182,In_224,N_503);
nor U1183 (N_1183,In_1741,N_154);
xor U1184 (N_1184,In_1798,In_880);
and U1185 (N_1185,N_178,N_269);
or U1186 (N_1186,N_96,N_106);
nand U1187 (N_1187,In_2049,N_395);
nor U1188 (N_1188,In_1634,In_140);
xor U1189 (N_1189,N_189,In_1346);
nand U1190 (N_1190,N_350,In_1461);
or U1191 (N_1191,In_1753,In_1237);
nand U1192 (N_1192,N_255,In_1729);
nor U1193 (N_1193,N_530,In_1723);
or U1194 (N_1194,N_71,N_550);
nor U1195 (N_1195,In_304,In_681);
and U1196 (N_1196,In_2062,In_2455);
nor U1197 (N_1197,N_428,In_1950);
or U1198 (N_1198,In_1807,N_237);
or U1199 (N_1199,In_1174,In_1878);
xnor U1200 (N_1200,In_2345,N_417);
nand U1201 (N_1201,In_2064,N_621);
and U1202 (N_1202,In_594,In_454);
xor U1203 (N_1203,N_306,In_1050);
xor U1204 (N_1204,In_1982,N_85);
and U1205 (N_1205,N_504,In_519);
nor U1206 (N_1206,In_2105,In_2351);
nor U1207 (N_1207,In_1561,In_1388);
nand U1208 (N_1208,In_1092,N_616);
xor U1209 (N_1209,N_406,N_37);
or U1210 (N_1210,In_1580,In_2278);
and U1211 (N_1211,In_172,In_89);
xnor U1212 (N_1212,In_847,N_421);
nand U1213 (N_1213,N_339,N_344);
nor U1214 (N_1214,In_2189,In_2194);
and U1215 (N_1215,In_1483,N_481);
nand U1216 (N_1216,In_2438,N_517);
nor U1217 (N_1217,N_568,N_286);
or U1218 (N_1218,N_399,In_1625);
xnor U1219 (N_1219,N_345,N_16);
xor U1220 (N_1220,N_375,In_1157);
or U1221 (N_1221,In_591,N_124);
and U1222 (N_1222,N_89,N_597);
or U1223 (N_1223,In_467,N_7);
and U1224 (N_1224,N_464,In_2426);
xor U1225 (N_1225,In_2139,N_93);
and U1226 (N_1226,N_104,In_1486);
or U1227 (N_1227,N_129,N_620);
nor U1228 (N_1228,In_2289,In_2199);
nor U1229 (N_1229,In_1281,N_317);
nand U1230 (N_1230,In_2321,In_505);
and U1231 (N_1231,In_2403,In_1751);
or U1232 (N_1232,In_2060,In_2209);
nor U1233 (N_1233,In_1442,N_531);
and U1234 (N_1234,In_1397,In_1421);
nand U1235 (N_1235,In_87,N_121);
and U1236 (N_1236,In_1722,N_147);
or U1237 (N_1237,N_184,N_572);
nor U1238 (N_1238,In_841,N_569);
and U1239 (N_1239,In_2344,N_486);
xnor U1240 (N_1240,N_58,In_1038);
nor U1241 (N_1241,In_1551,N_462);
nand U1242 (N_1242,N_28,In_952);
nand U1243 (N_1243,In_2198,In_714);
nor U1244 (N_1244,In_1053,In_1732);
nor U1245 (N_1245,N_56,N_608);
nand U1246 (N_1246,In_1280,N_65);
nor U1247 (N_1247,N_261,N_571);
nand U1248 (N_1248,In_560,In_420);
and U1249 (N_1249,N_496,In_1427);
nand U1250 (N_1250,In_1363,N_254);
xnor U1251 (N_1251,N_1028,In_1441);
or U1252 (N_1252,In_2410,N_18);
and U1253 (N_1253,In_1341,N_137);
xnor U1254 (N_1254,In_1113,In_256);
or U1255 (N_1255,In_1282,In_1323);
and U1256 (N_1256,N_643,N_1073);
nor U1257 (N_1257,N_1096,In_735);
nand U1258 (N_1258,N_218,N_1170);
nor U1259 (N_1259,N_441,N_424);
or U1260 (N_1260,In_1875,N_1112);
xnor U1261 (N_1261,N_1060,N_251);
and U1262 (N_1262,N_649,N_10);
xor U1263 (N_1263,In_1705,In_2298);
nor U1264 (N_1264,In_419,N_1199);
nand U1265 (N_1265,N_752,In_230);
or U1266 (N_1266,N_409,N_982);
and U1267 (N_1267,N_666,N_753);
xnor U1268 (N_1268,N_792,N_667);
nand U1269 (N_1269,N_1119,In_1340);
xnor U1270 (N_1270,N_977,N_609);
nand U1271 (N_1271,N_1074,N_1143);
nor U1272 (N_1272,N_653,N_656);
nand U1273 (N_1273,In_2031,In_2288);
and U1274 (N_1274,N_683,N_1233);
xor U1275 (N_1275,In_1834,N_1144);
nor U1276 (N_1276,N_1120,N_766);
or U1277 (N_1277,N_502,N_300);
nand U1278 (N_1278,In_1537,N_1080);
xnor U1279 (N_1279,N_804,N_746);
nand U1280 (N_1280,In_411,N_809);
and U1281 (N_1281,N_1042,N_826);
or U1282 (N_1282,N_1240,N_817);
nand U1283 (N_1283,N_892,N_832);
or U1284 (N_1284,N_413,N_974);
nand U1285 (N_1285,N_1129,N_903);
nor U1286 (N_1286,N_1141,In_1054);
xor U1287 (N_1287,N_432,N_1017);
or U1288 (N_1288,N_1039,N_1215);
or U1289 (N_1289,N_1205,In_1119);
or U1290 (N_1290,N_759,N_896);
or U1291 (N_1291,N_1196,N_1207);
xor U1292 (N_1292,N_914,N_1086);
nand U1293 (N_1293,N_936,N_1146);
and U1294 (N_1294,N_491,N_474);
and U1295 (N_1295,N_678,N_722);
and U1296 (N_1296,N_118,N_34);
nand U1297 (N_1297,In_2359,In_1270);
xnor U1298 (N_1298,N_760,N_909);
nand U1299 (N_1299,In_1227,N_427);
xor U1300 (N_1300,In_2348,N_786);
nor U1301 (N_1301,N_1116,N_593);
nand U1302 (N_1302,In_1277,N_1235);
nand U1303 (N_1303,N_980,N_1037);
or U1304 (N_1304,N_30,N_448);
nand U1305 (N_1305,N_975,In_182);
nand U1306 (N_1306,In_1715,N_776);
or U1307 (N_1307,N_26,In_864);
nor U1308 (N_1308,In_119,N_770);
and U1309 (N_1309,N_967,In_541);
and U1310 (N_1310,N_625,In_906);
nor U1311 (N_1311,N_538,In_1667);
xor U1312 (N_1312,In_725,In_1244);
xor U1313 (N_1313,N_443,N_500);
nor U1314 (N_1314,N_1072,N_661);
or U1315 (N_1315,N_1181,N_805);
or U1316 (N_1316,In_2218,In_683);
nand U1317 (N_1317,In_751,In_2233);
or U1318 (N_1318,N_956,N_67);
xnor U1319 (N_1319,N_1043,In_1193);
and U1320 (N_1320,N_1157,In_1475);
nor U1321 (N_1321,N_771,In_883);
nand U1322 (N_1322,N_1230,In_904);
nand U1323 (N_1323,In_1649,N_881);
xnor U1324 (N_1324,N_782,N_877);
or U1325 (N_1325,N_1133,In_1361);
nor U1326 (N_1326,N_1122,In_596);
and U1327 (N_1327,N_19,In_2362);
nor U1328 (N_1328,N_906,N_1049);
nand U1329 (N_1329,N_1204,N_659);
and U1330 (N_1330,In_855,N_972);
xor U1331 (N_1331,In_2166,N_183);
nand U1332 (N_1332,N_460,In_1815);
xnor U1333 (N_1333,N_800,N_640);
nor U1334 (N_1334,N_866,N_599);
and U1335 (N_1335,In_932,N_338);
xnor U1336 (N_1336,N_13,N_861);
or U1337 (N_1337,N_330,N_1203);
nand U1338 (N_1338,N_390,In_2259);
nor U1339 (N_1339,N_869,In_1031);
or U1340 (N_1340,N_657,N_1176);
or U1341 (N_1341,N_1171,In_1181);
nand U1342 (N_1342,N_938,N_638);
nor U1343 (N_1343,N_747,N_574);
xnor U1344 (N_1344,N_929,In_1884);
and U1345 (N_1345,N_1218,N_822);
nor U1346 (N_1346,In_1560,N_54);
or U1347 (N_1347,N_1100,N_783);
and U1348 (N_1348,In_2125,N_1022);
nor U1349 (N_1349,N_372,N_847);
xnor U1350 (N_1350,N_1241,In_1568);
nand U1351 (N_1351,N_885,N_860);
and U1352 (N_1352,In_1272,N_1082);
nand U1353 (N_1353,In_1694,In_6);
and U1354 (N_1354,N_55,In_849);
and U1355 (N_1355,In_1677,N_1193);
and U1356 (N_1356,In_894,N_644);
xnor U1357 (N_1357,N_333,In_2317);
xor U1358 (N_1358,N_207,N_1111);
and U1359 (N_1359,N_926,N_1046);
xnor U1360 (N_1360,N_1154,N_450);
nand U1361 (N_1361,N_1016,In_2364);
and U1362 (N_1362,N_1234,N_757);
nor U1363 (N_1363,N_435,In_2261);
and U1364 (N_1364,N_490,N_228);
nand U1365 (N_1365,N_662,In_2165);
nand U1366 (N_1366,In_30,N_652);
and U1367 (N_1367,N_762,In_1555);
nand U1368 (N_1368,N_1109,N_1209);
xnor U1369 (N_1369,In_840,In_756);
nand U1370 (N_1370,In_2262,N_1062);
xor U1371 (N_1371,In_10,N_1058);
nand U1372 (N_1372,N_848,N_1076);
nor U1373 (N_1373,In_1748,N_1167);
xor U1374 (N_1374,N_672,N_619);
nor U1375 (N_1375,N_192,N_951);
and U1376 (N_1376,N_90,In_1177);
nand U1377 (N_1377,In_86,In_98);
xor U1378 (N_1378,In_14,In_825);
and U1379 (N_1379,In_737,N_750);
nand U1380 (N_1380,In_2291,In_1540);
or U1381 (N_1381,In_1330,N_1186);
nor U1382 (N_1382,N_917,In_1541);
nand U1383 (N_1383,N_704,N_895);
and U1384 (N_1384,N_581,N_1145);
nor U1385 (N_1385,N_175,N_684);
nor U1386 (N_1386,N_1114,N_803);
nand U1387 (N_1387,In_2265,N_962);
nor U1388 (N_1388,In_630,N_952);
and U1389 (N_1389,N_9,N_1012);
nor U1390 (N_1390,In_842,In_2047);
xor U1391 (N_1391,N_699,N_1142);
and U1392 (N_1392,N_1106,In_1611);
nor U1393 (N_1393,N_418,In_806);
and U1394 (N_1394,N_883,N_912);
xnor U1395 (N_1395,N_1174,In_1550);
xor U1396 (N_1396,In_1396,N_841);
and U1397 (N_1397,In_1284,In_1274);
and U1398 (N_1398,N_277,N_188);
nor U1399 (N_1399,N_874,N_953);
and U1400 (N_1400,N_305,In_2468);
or U1401 (N_1401,In_1159,N_751);
nor U1402 (N_1402,N_971,In_2205);
xnor U1403 (N_1403,In_798,In_2251);
nand U1404 (N_1404,In_100,N_969);
nor U1405 (N_1405,N_973,N_1032);
nand U1406 (N_1406,N_380,N_820);
and U1407 (N_1407,N_930,In_1837);
nor U1408 (N_1408,In_1110,In_151);
nor U1409 (N_1409,N_51,N_837);
nand U1410 (N_1410,N_1011,In_1930);
nor U1411 (N_1411,N_1208,N_1224);
and U1412 (N_1412,N_979,N_1041);
nor U1413 (N_1413,N_1030,In_238);
or U1414 (N_1414,N_74,N_1151);
nand U1415 (N_1415,N_302,N_617);
and U1416 (N_1416,N_1138,N_996);
nor U1417 (N_1417,In_2243,N_887);
xnor U1418 (N_1418,N_677,N_937);
and U1419 (N_1419,N_416,N_1038);
or U1420 (N_1420,In_1012,N_993);
nor U1421 (N_1421,N_1020,In_597);
nor U1422 (N_1422,In_1440,N_921);
nand U1423 (N_1423,N_651,In_1757);
or U1424 (N_1424,N_1110,In_1249);
xor U1425 (N_1425,In_982,N_816);
nand U1426 (N_1426,In_197,In_2448);
nand U1427 (N_1427,N_414,N_243);
nor U1428 (N_1428,N_674,N_829);
nor U1429 (N_1429,In_1357,N_1088);
or U1430 (N_1430,In_1209,In_2098);
xor U1431 (N_1431,N_1162,N_729);
xnor U1432 (N_1432,N_415,In_1711);
and U1433 (N_1433,N_642,N_724);
and U1434 (N_1434,N_890,In_120);
or U1435 (N_1435,In_1095,N_984);
or U1436 (N_1436,In_1117,N_1191);
or U1437 (N_1437,N_1136,N_695);
and U1438 (N_1438,In_2241,In_2129);
nand U1439 (N_1439,N_598,In_1593);
or U1440 (N_1440,N_626,N_629);
nor U1441 (N_1441,N_646,N_1212);
nand U1442 (N_1442,N_827,N_908);
and U1443 (N_1443,In_1393,N_473);
xnor U1444 (N_1444,N_585,N_227);
or U1445 (N_1445,In_1511,N_1081);
nor U1446 (N_1446,N_1090,N_444);
or U1447 (N_1447,N_1068,N_781);
xor U1448 (N_1448,In_777,N_1093);
or U1449 (N_1449,In_2036,N_806);
nand U1450 (N_1450,N_1201,N_66);
or U1451 (N_1451,In_1869,N_436);
xnor U1452 (N_1452,N_1244,N_403);
nor U1453 (N_1453,N_808,N_1226);
nand U1454 (N_1454,N_1147,N_145);
nand U1455 (N_1455,N_999,N_247);
nand U1456 (N_1456,In_1,N_796);
and U1457 (N_1457,In_1178,N_1025);
nor U1458 (N_1458,N_1014,N_945);
or U1459 (N_1459,N_1211,N_878);
or U1460 (N_1460,N_388,N_867);
nand U1461 (N_1461,N_1220,N_201);
or U1462 (N_1462,In_96,N_948);
xnor U1463 (N_1463,N_955,N_1001);
and U1464 (N_1464,N_765,N_690);
or U1465 (N_1465,N_1057,N_1095);
nor U1466 (N_1466,N_510,N_723);
and U1467 (N_1467,N_1187,In_632);
nand U1468 (N_1468,N_864,N_1034);
nor U1469 (N_1469,N_373,N_1121);
and U1470 (N_1470,In_827,In_144);
nor U1471 (N_1471,N_193,N_580);
and U1472 (N_1472,N_232,N_136);
xor U1473 (N_1473,N_833,N_995);
or U1474 (N_1474,N_351,N_576);
xor U1475 (N_1475,N_697,In_330);
or U1476 (N_1476,N_22,N_1031);
or U1477 (N_1477,N_946,In_2393);
xnor U1478 (N_1478,N_1108,In_925);
nand U1479 (N_1479,In_1337,In_2015);
xnor U1480 (N_1480,N_981,In_1217);
or U1481 (N_1481,In_710,In_77);
nor U1482 (N_1482,N_288,N_1155);
or U1483 (N_1483,N_144,N_42);
or U1484 (N_1484,N_850,N_1113);
xnor U1485 (N_1485,N_554,N_978);
or U1486 (N_1486,N_714,In_1794);
nand U1487 (N_1487,N_1243,N_1015);
or U1488 (N_1488,In_1811,N_1149);
nor U1489 (N_1489,N_1177,N_127);
and U1490 (N_1490,N_741,N_465);
nand U1491 (N_1491,N_507,N_902);
nand U1492 (N_1492,N_910,N_899);
nand U1493 (N_1493,In_2330,In_1522);
and U1494 (N_1494,In_207,N_1078);
xor U1495 (N_1495,N_813,N_888);
and U1496 (N_1496,In_1015,N_788);
and U1497 (N_1497,In_657,N_342);
or U1498 (N_1498,N_811,In_1718);
nand U1499 (N_1499,In_1352,In_1862);
xnor U1500 (N_1500,N_1127,N_968);
or U1501 (N_1501,N_990,In_1516);
xnor U1502 (N_1502,N_679,N_834);
and U1503 (N_1503,In_1923,In_1663);
nor U1504 (N_1504,In_2456,N_718);
and U1505 (N_1505,N_1105,N_1019);
xor U1506 (N_1506,N_60,N_105);
nand U1507 (N_1507,In_1432,N_1045);
nand U1508 (N_1508,N_745,N_641);
xnor U1509 (N_1509,In_2412,N_1228);
xor U1510 (N_1510,In_2130,In_536);
and U1511 (N_1511,N_138,N_669);
xor U1512 (N_1512,N_680,N_992);
xor U1513 (N_1513,N_1024,In_383);
xor U1514 (N_1514,In_236,In_246);
nor U1515 (N_1515,N_849,N_226);
or U1516 (N_1516,N_1169,N_670);
xnor U1517 (N_1517,In_774,In_1967);
and U1518 (N_1518,N_710,N_1159);
or U1519 (N_1519,N_727,In_387);
nand U1520 (N_1520,N_1064,N_754);
nand U1521 (N_1521,N_135,N_842);
nand U1522 (N_1522,N_919,In_1674);
and U1523 (N_1523,N_470,In_1567);
nor U1524 (N_1524,N_725,In_837);
nor U1525 (N_1525,In_1074,N_959);
and U1526 (N_1526,In_1941,In_2085);
nand U1527 (N_1527,In_1458,N_859);
or U1528 (N_1528,N_655,In_1841);
or U1529 (N_1529,In_2200,N_506);
and U1530 (N_1530,In_412,In_461);
and U1531 (N_1531,In_1785,N_731);
nor U1532 (N_1532,In_620,N_1160);
or U1533 (N_1533,N_1231,N_898);
xor U1534 (N_1534,In_811,N_214);
nand U1535 (N_1535,In_580,In_1587);
and U1536 (N_1536,N_924,N_844);
nor U1537 (N_1537,N_1188,In_1061);
xnor U1538 (N_1538,In_805,In_483);
xor U1539 (N_1539,N_647,N_701);
or U1540 (N_1540,In_2245,In_863);
and U1541 (N_1541,N_595,N_940);
or U1542 (N_1542,N_139,In_225);
nand U1543 (N_1543,N_884,In_215);
and U1544 (N_1544,N_391,N_1249);
nand U1545 (N_1545,In_957,N_1164);
nand U1546 (N_1546,N_1216,N_468);
xnor U1547 (N_1547,N_853,In_388);
xnor U1548 (N_1548,N_540,N_1128);
nand U1549 (N_1549,In_1570,N_686);
nand U1550 (N_1550,N_720,N_685);
or U1551 (N_1551,N_735,In_485);
xor U1552 (N_1552,In_1105,N_292);
or U1553 (N_1553,In_1616,In_819);
nor U1554 (N_1554,In_793,N_282);
nand U1555 (N_1555,N_645,In_1924);
xor U1556 (N_1556,N_1238,N_27);
nand U1557 (N_1557,N_769,N_728);
xnor U1558 (N_1558,N_1236,N_1229);
and U1559 (N_1559,N_82,N_880);
and U1560 (N_1560,N_733,N_862);
xor U1561 (N_1561,In_991,N_857);
nor U1562 (N_1562,In_1710,N_692);
or U1563 (N_1563,N_1013,N_293);
xnor U1564 (N_1564,N_900,N_526);
and U1565 (N_1565,N_458,N_1056);
xnor U1566 (N_1566,In_1610,N_681);
nor U1567 (N_1567,In_1465,In_1064);
and U1568 (N_1568,N_707,N_1101);
and U1569 (N_1569,N_821,In_713);
nor U1570 (N_1570,N_1223,In_784);
nor U1571 (N_1571,N_789,N_868);
or U1572 (N_1572,In_845,In_1755);
nor U1573 (N_1573,N_1202,N_326);
nand U1574 (N_1574,N_181,N_957);
nand U1575 (N_1575,In_1609,N_1172);
and U1576 (N_1576,N_814,N_758);
xor U1577 (N_1577,In_184,N_931);
xnor U1578 (N_1578,N_854,N_1148);
and U1579 (N_1579,N_1123,In_1129);
nand U1580 (N_1580,In_2113,N_426);
nand U1581 (N_1581,N_611,N_1194);
or U1582 (N_1582,In_1767,N_705);
xor U1583 (N_1583,N_1183,In_2361);
xor U1584 (N_1584,In_694,In_155);
xor U1585 (N_1585,N_1227,In_1127);
nor U1586 (N_1586,N_818,In_31);
nand U1587 (N_1587,In_645,N_1050);
xnor U1588 (N_1588,In_1135,N_110);
or U1589 (N_1589,N_694,N_1185);
nor U1590 (N_1590,N_872,N_1214);
nor U1591 (N_1591,In_2188,In_1526);
nand U1592 (N_1592,In_1919,N_976);
and U1593 (N_1593,N_1097,In_498);
xnor U1594 (N_1594,N_756,N_852);
xnor U1595 (N_1595,N_23,N_59);
and U1596 (N_1596,In_469,In_160);
and U1597 (N_1597,N_703,In_603);
and U1598 (N_1598,N_298,N_1166);
xor U1599 (N_1599,N_904,In_2071);
and U1600 (N_1600,N_671,In_2275);
nand U1601 (N_1601,N_791,N_772);
nor U1602 (N_1602,In_1801,N_698);
nor U1603 (N_1603,N_665,N_856);
nand U1604 (N_1604,In_1944,N_1006);
xor U1605 (N_1605,N_487,N_960);
nand U1606 (N_1606,In_1829,N_950);
nor U1607 (N_1607,N_1210,N_627);
nor U1608 (N_1608,N_1225,In_752);
nor U1609 (N_1609,N_966,In_1665);
nand U1610 (N_1610,N_863,N_301);
nor U1611 (N_1611,In_458,N_1152);
or U1612 (N_1612,N_223,N_944);
or U1613 (N_1613,N_49,In_676);
or U1614 (N_1614,N_812,N_319);
and U1615 (N_1615,N_346,N_1091);
and U1616 (N_1616,N_573,N_660);
nor U1617 (N_1617,In_1289,N_706);
and U1618 (N_1618,In_585,N_632);
or U1619 (N_1619,In_2147,N_911);
xor U1620 (N_1620,N_128,N_737);
nor U1621 (N_1621,N_631,N_700);
nand U1622 (N_1622,In_1808,N_918);
or U1623 (N_1623,In_909,N_987);
nor U1624 (N_1624,In_1790,N_779);
nand U1625 (N_1625,N_768,N_839);
nor U1626 (N_1626,N_650,N_1222);
or U1627 (N_1627,N_248,N_709);
or U1628 (N_1628,N_835,N_553);
and U1629 (N_1629,N_77,N_1124);
nor U1630 (N_1630,N_1132,In_965);
nand U1631 (N_1631,N_648,N_570);
or U1632 (N_1632,N_297,In_2142);
and U1633 (N_1633,N_964,N_1010);
xnor U1634 (N_1634,N_635,In_2186);
nor U1635 (N_1635,N_528,In_646);
nand U1636 (N_1636,N_1232,N_876);
and U1637 (N_1637,N_734,In_1532);
nor U1638 (N_1638,N_235,N_1069);
nand U1639 (N_1639,N_846,In_1504);
nor U1640 (N_1640,In_846,N_1156);
nand U1641 (N_1641,In_858,In_1218);
nor U1642 (N_1642,N_1065,In_490);
and U1643 (N_1643,N_711,N_889);
nor U1644 (N_1644,N_934,N_913);
and U1645 (N_1645,In_659,N_1173);
or U1646 (N_1646,N_965,In_2011);
and U1647 (N_1647,N_668,In_2276);
xor U1648 (N_1648,In_729,N_1000);
and U1649 (N_1649,N_865,N_1066);
and U1650 (N_1650,N_615,N_161);
xor U1651 (N_1651,N_1180,N_658);
nand U1652 (N_1652,N_157,N_954);
xnor U1653 (N_1653,In_70,N_244);
nand U1654 (N_1654,N_200,N_1048);
nand U1655 (N_1655,In_271,In_1692);
xor U1656 (N_1656,In_947,In_2050);
and U1657 (N_1657,N_81,In_1758);
nand U1658 (N_1658,N_449,In_2097);
nand U1659 (N_1659,N_702,N_1070);
nor U1660 (N_1660,N_970,In_1752);
or U1661 (N_1661,N_1248,N_721);
nand U1662 (N_1662,N_1071,In_361);
and U1663 (N_1663,N_209,N_825);
nand U1664 (N_1664,In_1577,N_1165);
or U1665 (N_1665,N_122,In_1111);
xor U1666 (N_1666,N_691,N_359);
and U1667 (N_1667,In_463,In_582);
xnor U1668 (N_1668,In_2453,N_199);
xnor U1669 (N_1669,In_896,N_1040);
or U1670 (N_1670,N_716,N_828);
xor U1671 (N_1671,N_521,In_850);
or U1672 (N_1672,In_181,N_336);
nor U1673 (N_1673,N_606,N_1059);
xor U1674 (N_1674,N_675,In_556);
or U1675 (N_1675,In_1579,N_893);
or U1676 (N_1676,In_1818,N_764);
or U1677 (N_1677,N_1200,In_1457);
and U1678 (N_1678,N_1206,N_555);
xnor U1679 (N_1679,N_84,N_744);
nand U1680 (N_1680,N_1131,In_2354);
nand U1681 (N_1681,In_1877,N_361);
or U1682 (N_1682,N_916,N_1197);
and U1683 (N_1683,N_605,In_776);
nor U1684 (N_1684,N_264,In_1951);
xor U1685 (N_1685,N_664,N_1246);
nor U1686 (N_1686,In_1978,In_2424);
and U1687 (N_1687,In_118,N_1099);
nor U1688 (N_1688,In_2222,N_810);
nand U1689 (N_1689,In_625,In_584);
nor U1690 (N_1690,In_1082,N_1021);
and U1691 (N_1691,N_152,In_1889);
or U1692 (N_1692,In_2123,N_749);
nand U1693 (N_1693,In_1719,N_1125);
nand U1694 (N_1694,N_220,In_2492);
and U1695 (N_1695,N_636,N_307);
xor U1696 (N_1696,N_607,N_313);
nor U1697 (N_1697,In_1704,N_693);
nand U1698 (N_1698,In_1657,N_961);
nand U1699 (N_1699,N_739,N_1083);
nor U1700 (N_1700,N_998,N_958);
and U1701 (N_1701,N_732,N_715);
nor U1702 (N_1702,N_1079,N_32);
nand U1703 (N_1703,N_1061,In_758);
xor U1704 (N_1704,N_799,N_1098);
xnor U1705 (N_1705,N_708,N_807);
and U1706 (N_1706,N_935,N_523);
and U1707 (N_1707,In_321,N_1052);
and U1708 (N_1708,In_1844,N_763);
xnor U1709 (N_1709,N_1077,N_823);
or U1710 (N_1710,N_47,N_840);
xnor U1711 (N_1711,N_933,N_907);
xnor U1712 (N_1712,In_1115,N_824);
or U1713 (N_1713,N_730,N_1023);
or U1714 (N_1714,N_485,N_1115);
nand U1715 (N_1715,N_985,N_1150);
nor U1716 (N_1716,N_726,N_272);
nand U1717 (N_1717,N_95,In_2048);
xor U1718 (N_1718,N_1029,In_791);
or U1719 (N_1719,N_1003,N_639);
or U1720 (N_1720,N_1026,In_130);
or U1721 (N_1721,N_513,In_564);
nor U1722 (N_1722,N_543,In_440);
and U1723 (N_1723,N_949,In_1422);
nor U1724 (N_1724,N_774,N_1245);
nand U1725 (N_1725,In_95,N_736);
or U1726 (N_1726,In_648,In_392);
nor U1727 (N_1727,N_381,N_309);
and U1728 (N_1728,N_215,N_392);
xor U1729 (N_1729,N_1158,In_2022);
nor U1730 (N_1730,N_182,In_1646);
nand U1731 (N_1731,N_787,In_1295);
or U1732 (N_1732,N_795,N_1103);
and U1733 (N_1733,In_1202,N_1135);
xor U1734 (N_1734,In_2329,N_794);
nand U1735 (N_1735,In_2300,N_855);
xor U1736 (N_1736,In_866,In_1487);
or U1737 (N_1737,N_905,N_742);
nand U1738 (N_1738,N_994,N_845);
nor U1739 (N_1739,In_998,N_873);
nor U1740 (N_1740,N_92,N_1008);
nand U1741 (N_1741,In_341,In_2184);
nand U1742 (N_1742,N_897,N_843);
nor U1743 (N_1743,N_1242,In_1308);
xnor U1744 (N_1744,In_427,In_382);
nor U1745 (N_1745,In_1118,In_2144);
or U1746 (N_1746,N_712,N_696);
and U1747 (N_1747,N_1051,N_340);
nor U1748 (N_1748,N_630,N_524);
or U1749 (N_1749,N_830,In_2339);
xor U1750 (N_1750,N_886,N_943);
nor U1751 (N_1751,In_109,In_2000);
xnor U1752 (N_1752,N_1002,In_408);
nor U1753 (N_1753,N_988,N_1184);
nor U1754 (N_1754,N_923,N_628);
xnor U1755 (N_1755,N_552,In_2030);
and U1756 (N_1756,N_1044,In_1887);
nand U1757 (N_1757,N_748,N_321);
or U1758 (N_1758,N_780,N_208);
xnor U1759 (N_1759,N_894,In_1912);
and U1760 (N_1760,In_2231,N_1134);
and U1761 (N_1761,N_1033,N_775);
xnor U1762 (N_1762,In_1836,N_170);
nor U1763 (N_1763,In_2004,N_134);
nand U1764 (N_1764,In_1874,N_1007);
xor U1765 (N_1765,In_1564,In_439);
or U1766 (N_1766,In_987,N_1163);
nand U1767 (N_1767,In_2012,N_963);
or U1768 (N_1768,N_1140,In_1049);
nand U1769 (N_1769,N_265,N_713);
xnor U1770 (N_1770,N_891,N_1067);
xor U1771 (N_1771,N_1084,N_922);
xnor U1772 (N_1772,N_1035,In_2055);
and U1773 (N_1773,N_41,In_2175);
nand U1774 (N_1774,In_1056,N_997);
and U1775 (N_1775,N_1175,N_1189);
nor U1776 (N_1776,N_831,N_901);
nor U1777 (N_1777,N_1237,N_939);
and U1778 (N_1778,N_213,N_1027);
or U1779 (N_1779,In_219,In_813);
and U1780 (N_1780,N_1054,N_439);
and U1781 (N_1781,N_871,N_761);
xnor U1782 (N_1782,N_564,N_986);
xnor U1783 (N_1783,N_1130,In_2169);
nand U1784 (N_1784,N_270,In_643);
nor U1785 (N_1785,N_1221,N_1092);
or U1786 (N_1786,N_1047,N_257);
nand U1787 (N_1787,In_1194,N_535);
xnor U1788 (N_1788,In_198,In_2290);
xor U1789 (N_1789,In_510,N_1179);
nand U1790 (N_1790,N_1087,N_1178);
or U1791 (N_1791,In_1306,In_360);
nand U1792 (N_1792,N_767,N_1126);
xor U1793 (N_1793,N_633,In_999);
nor U1794 (N_1794,N_676,N_379);
nor U1795 (N_1795,In_1999,In_129);
nand U1796 (N_1796,N_654,N_717);
nand U1797 (N_1797,In_136,In_1033);
or U1798 (N_1798,N_370,In_481);
xnor U1799 (N_1799,N_167,N_1161);
nor U1800 (N_1800,N_1195,In_780);
nand U1801 (N_1801,In_1163,N_275);
nand U1802 (N_1802,N_1102,N_1018);
and U1803 (N_1803,N_777,N_1192);
nand U1804 (N_1804,N_296,N_11);
nand U1805 (N_1805,N_525,N_44);
nor U1806 (N_1806,N_838,N_1009);
xor U1807 (N_1807,In_1109,In_323);
nand U1808 (N_1808,In_1026,N_512);
or U1809 (N_1809,N_875,N_773);
nor U1810 (N_1810,N_560,In_870);
nor U1811 (N_1811,N_1118,N_688);
and U1812 (N_1812,N_687,N_858);
xor U1813 (N_1813,N_1168,In_1955);
nor U1814 (N_1814,In_1812,N_740);
xor U1815 (N_1815,N_367,In_1706);
and U1816 (N_1816,In_601,N_1089);
nor U1817 (N_1817,N_1085,N_793);
nor U1818 (N_1818,N_925,N_1104);
xor U1819 (N_1819,N_1139,N_790);
or U1820 (N_1820,N_778,N_719);
or U1821 (N_1821,N_801,In_727);
nand U1822 (N_1822,N_371,N_1107);
nand U1823 (N_1823,N_785,In_328);
xor U1824 (N_1824,In_1302,In_455);
nor U1825 (N_1825,N_1198,N_634);
xnor U1826 (N_1826,N_738,In_881);
or U1827 (N_1827,N_1063,In_1384);
and U1828 (N_1828,N_217,N_78);
and U1829 (N_1829,N_682,N_991);
and U1830 (N_1830,N_851,N_927);
nor U1831 (N_1831,In_1574,In_506);
xor U1832 (N_1832,N_920,In_1265);
nor U1833 (N_1833,N_1075,In_1779);
nand U1834 (N_1834,N_397,N_1137);
xnor U1835 (N_1835,N_1217,N_1094);
nand U1836 (N_1836,In_2253,N_915);
or U1837 (N_1837,In_1542,N_165);
and U1838 (N_1838,N_673,N_1247);
xnor U1839 (N_1839,In_875,N_836);
nor U1840 (N_1840,N_1036,In_769);
nor U1841 (N_1841,N_1219,N_932);
nor U1842 (N_1842,N_663,In_1548);
or U1843 (N_1843,In_1682,In_586);
nand U1844 (N_1844,N_194,N_797);
xor U1845 (N_1845,N_613,In_425);
xor U1846 (N_1846,N_1182,N_1117);
or U1847 (N_1847,In_1057,N_1005);
nand U1848 (N_1848,N_947,N_72);
or U1849 (N_1849,N_437,In_1645);
nor U1850 (N_1850,N_802,In_1180);
nand U1851 (N_1851,N_356,N_941);
nand U1852 (N_1852,N_461,N_101);
or U1853 (N_1853,In_16,N_1053);
or U1854 (N_1854,In_638,N_983);
xor U1855 (N_1855,N_870,N_398);
nand U1856 (N_1856,N_743,In_606);
nor U1857 (N_1857,N_882,In_101);
or U1858 (N_1858,N_1239,In_1496);
xor U1859 (N_1859,N_989,N_224);
xor U1860 (N_1860,In_953,N_1190);
nand U1861 (N_1861,In_1820,N_1153);
xnor U1862 (N_1862,N_798,N_819);
nor U1863 (N_1863,N_755,N_422);
and U1864 (N_1864,N_928,N_689);
and U1865 (N_1865,In_2296,N_1055);
nand U1866 (N_1866,N_879,N_637);
nand U1867 (N_1867,In_1972,In_885);
and U1868 (N_1868,In_697,N_1004);
xnor U1869 (N_1869,N_1213,N_784);
nor U1870 (N_1870,N_815,N_584);
nand U1871 (N_1871,In_2417,In_2324);
and U1872 (N_1872,N_280,N_589);
nor U1873 (N_1873,N_942,N_150);
xor U1874 (N_1874,In_968,N_141);
or U1875 (N_1875,N_1311,N_1442);
nor U1876 (N_1876,N_1649,N_1280);
or U1877 (N_1877,N_1752,N_1449);
nor U1878 (N_1878,N_1750,N_1406);
nor U1879 (N_1879,N_1781,N_1317);
and U1880 (N_1880,N_1509,N_1265);
or U1881 (N_1881,N_1809,N_1467);
or U1882 (N_1882,N_1388,N_1636);
nand U1883 (N_1883,N_1275,N_1641);
nand U1884 (N_1884,N_1721,N_1692);
and U1885 (N_1885,N_1375,N_1776);
nor U1886 (N_1886,N_1592,N_1686);
xor U1887 (N_1887,N_1754,N_1260);
nand U1888 (N_1888,N_1550,N_1552);
and U1889 (N_1889,N_1476,N_1354);
and U1890 (N_1890,N_1570,N_1766);
nor U1891 (N_1891,N_1489,N_1832);
and U1892 (N_1892,N_1808,N_1846);
nand U1893 (N_1893,N_1409,N_1800);
nor U1894 (N_1894,N_1868,N_1432);
nor U1895 (N_1895,N_1748,N_1296);
xor U1896 (N_1896,N_1820,N_1517);
and U1897 (N_1897,N_1500,N_1605);
and U1898 (N_1898,N_1431,N_1870);
nand U1899 (N_1899,N_1333,N_1510);
and U1900 (N_1900,N_1858,N_1305);
and U1901 (N_1901,N_1697,N_1606);
and U1902 (N_1902,N_1586,N_1661);
xor U1903 (N_1903,N_1698,N_1745);
or U1904 (N_1904,N_1775,N_1612);
and U1905 (N_1905,N_1370,N_1648);
and U1906 (N_1906,N_1443,N_1621);
nand U1907 (N_1907,N_1380,N_1768);
nand U1908 (N_1908,N_1471,N_1310);
and U1909 (N_1909,N_1864,N_1600);
and U1910 (N_1910,N_1741,N_1717);
and U1911 (N_1911,N_1321,N_1787);
nand U1912 (N_1912,N_1282,N_1426);
or U1913 (N_1913,N_1546,N_1695);
and U1914 (N_1914,N_1620,N_1734);
xnor U1915 (N_1915,N_1325,N_1551);
nor U1916 (N_1916,N_1849,N_1299);
nor U1917 (N_1917,N_1503,N_1462);
and U1918 (N_1918,N_1323,N_1516);
nand U1919 (N_1919,N_1716,N_1292);
nor U1920 (N_1920,N_1785,N_1491);
and U1921 (N_1921,N_1535,N_1690);
and U1922 (N_1922,N_1660,N_1414);
and U1923 (N_1923,N_1663,N_1278);
xor U1924 (N_1924,N_1297,N_1378);
nor U1925 (N_1925,N_1304,N_1587);
nand U1926 (N_1926,N_1344,N_1543);
nand U1927 (N_1927,N_1658,N_1622);
and U1928 (N_1928,N_1420,N_1682);
nor U1929 (N_1929,N_1330,N_1392);
nand U1930 (N_1930,N_1839,N_1677);
xor U1931 (N_1931,N_1367,N_1261);
nand U1932 (N_1932,N_1457,N_1525);
nor U1933 (N_1933,N_1404,N_1687);
xor U1934 (N_1934,N_1450,N_1867);
nor U1935 (N_1935,N_1508,N_1316);
xnor U1936 (N_1936,N_1685,N_1684);
and U1937 (N_1937,N_1396,N_1482);
xnor U1938 (N_1938,N_1593,N_1262);
or U1939 (N_1939,N_1738,N_1564);
and U1940 (N_1940,N_1637,N_1788);
nor U1941 (N_1941,N_1329,N_1258);
or U1942 (N_1942,N_1452,N_1324);
or U1943 (N_1943,N_1514,N_1633);
nand U1944 (N_1944,N_1873,N_1712);
nor U1945 (N_1945,N_1328,N_1521);
and U1946 (N_1946,N_1838,N_1263);
or U1947 (N_1947,N_1363,N_1368);
nand U1948 (N_1948,N_1577,N_1290);
xor U1949 (N_1949,N_1713,N_1287);
xnor U1950 (N_1950,N_1607,N_1831);
xnor U1951 (N_1951,N_1585,N_1553);
or U1952 (N_1952,N_1408,N_1594);
xnor U1953 (N_1953,N_1519,N_1722);
or U1954 (N_1954,N_1447,N_1761);
or U1955 (N_1955,N_1411,N_1778);
and U1956 (N_1956,N_1495,N_1731);
or U1957 (N_1957,N_1665,N_1478);
nor U1958 (N_1958,N_1874,N_1861);
nand U1959 (N_1959,N_1298,N_1494);
xor U1960 (N_1960,N_1827,N_1609);
xnor U1961 (N_1961,N_1430,N_1259);
xor U1962 (N_1962,N_1817,N_1705);
or U1963 (N_1963,N_1554,N_1751);
xor U1964 (N_1964,N_1309,N_1456);
and U1965 (N_1965,N_1853,N_1353);
xor U1966 (N_1966,N_1582,N_1739);
or U1967 (N_1967,N_1847,N_1529);
or U1968 (N_1968,N_1611,N_1446);
and U1969 (N_1969,N_1528,N_1373);
xnor U1970 (N_1970,N_1374,N_1691);
or U1971 (N_1971,N_1294,N_1301);
xor U1972 (N_1972,N_1393,N_1279);
xnor U1973 (N_1973,N_1589,N_1340);
and U1974 (N_1974,N_1556,N_1657);
or U1975 (N_1975,N_1773,N_1436);
nor U1976 (N_1976,N_1782,N_1771);
xor U1977 (N_1977,N_1357,N_1567);
nor U1978 (N_1978,N_1578,N_1531);
xor U1979 (N_1979,N_1410,N_1557);
xor U1980 (N_1980,N_1696,N_1810);
nand U1981 (N_1981,N_1295,N_1327);
and U1982 (N_1982,N_1616,N_1670);
nand U1983 (N_1983,N_1271,N_1512);
xnor U1984 (N_1984,N_1473,N_1459);
and U1985 (N_1985,N_1399,N_1255);
xor U1986 (N_1986,N_1797,N_1477);
nand U1987 (N_1987,N_1326,N_1439);
xor U1988 (N_1988,N_1719,N_1451);
nand U1989 (N_1989,N_1866,N_1850);
nand U1990 (N_1990,N_1701,N_1822);
or U1991 (N_1991,N_1569,N_1795);
or U1992 (N_1992,N_1842,N_1837);
xor U1993 (N_1993,N_1575,N_1400);
or U1994 (N_1994,N_1726,N_1794);
nor U1995 (N_1995,N_1490,N_1863);
or U1996 (N_1996,N_1843,N_1848);
and U1997 (N_1997,N_1468,N_1799);
nand U1998 (N_1998,N_1427,N_1798);
xnor U1999 (N_1999,N_1707,N_1454);
or U2000 (N_2000,N_1656,N_1763);
xnor U2001 (N_2001,N_1421,N_1676);
and U2002 (N_2002,N_1497,N_1816);
xor U2003 (N_2003,N_1654,N_1683);
nand U2004 (N_2004,N_1267,N_1276);
nand U2005 (N_2005,N_1617,N_1461);
nand U2006 (N_2006,N_1384,N_1610);
nor U2007 (N_2007,N_1505,N_1804);
nand U2008 (N_2008,N_1708,N_1520);
nor U2009 (N_2009,N_1308,N_1693);
nor U2010 (N_2010,N_1407,N_1671);
or U2011 (N_2011,N_1869,N_1472);
and U2012 (N_2012,N_1549,N_1428);
or U2013 (N_2013,N_1780,N_1285);
and U2014 (N_2014,N_1742,N_1253);
xnor U2015 (N_2015,N_1591,N_1563);
nand U2016 (N_2016,N_1540,N_1349);
or U2017 (N_2017,N_1257,N_1424);
nand U2018 (N_2018,N_1796,N_1283);
nor U2019 (N_2019,N_1437,N_1281);
and U2020 (N_2020,N_1678,N_1581);
nand U2021 (N_2021,N_1448,N_1523);
and U2022 (N_2022,N_1642,N_1562);
or U2023 (N_2023,N_1635,N_1499);
and U2024 (N_2024,N_1871,N_1312);
nor U2025 (N_2025,N_1830,N_1250);
xor U2026 (N_2026,N_1845,N_1627);
xor U2027 (N_2027,N_1366,N_1792);
xor U2028 (N_2028,N_1560,N_1835);
nand U2029 (N_2029,N_1545,N_1624);
xor U2030 (N_2030,N_1706,N_1568);
or U2031 (N_2031,N_1433,N_1851);
nand U2032 (N_2032,N_1369,N_1727);
and U2033 (N_2033,N_1429,N_1416);
and U2034 (N_2034,N_1479,N_1615);
nand U2035 (N_2035,N_1856,N_1595);
nand U2036 (N_2036,N_1361,N_1371);
and U2037 (N_2037,N_1266,N_1632);
or U2038 (N_2038,N_1815,N_1653);
or U2039 (N_2039,N_1802,N_1288);
and U2040 (N_2040,N_1664,N_1526);
nor U2041 (N_2041,N_1537,N_1302);
xnor U2042 (N_2042,N_1710,N_1498);
and U2043 (N_2043,N_1320,N_1511);
xor U2044 (N_2044,N_1558,N_1694);
xor U2045 (N_2045,N_1355,N_1854);
or U2046 (N_2046,N_1791,N_1756);
nand U2047 (N_2047,N_1565,N_1474);
nand U2048 (N_2048,N_1566,N_1645);
nand U2049 (N_2049,N_1662,N_1358);
nor U2050 (N_2050,N_1572,N_1732);
nor U2051 (N_2051,N_1669,N_1372);
xnor U2052 (N_2052,N_1397,N_1524);
nand U2053 (N_2053,N_1395,N_1415);
or U2054 (N_2054,N_1533,N_1646);
or U2055 (N_2055,N_1840,N_1322);
nand U2056 (N_2056,N_1501,N_1862);
or U2057 (N_2057,N_1453,N_1650);
xor U2058 (N_2058,N_1762,N_1680);
xor U2059 (N_2059,N_1289,N_1619);
or U2060 (N_2060,N_1484,N_1507);
and U2061 (N_2061,N_1826,N_1640);
xnor U2062 (N_2062,N_1841,N_1655);
nor U2063 (N_2063,N_1573,N_1291);
or U2064 (N_2064,N_1651,N_1613);
or U2065 (N_2065,N_1814,N_1597);
and U2066 (N_2066,N_1718,N_1382);
nand U2067 (N_2067,N_1749,N_1688);
xor U2068 (N_2068,N_1379,N_1737);
nor U2069 (N_2069,N_1269,N_1438);
xnor U2070 (N_2070,N_1376,N_1347);
or U2071 (N_2071,N_1398,N_1747);
or U2072 (N_2072,N_1541,N_1532);
or U2073 (N_2073,N_1647,N_1760);
nand U2074 (N_2074,N_1307,N_1784);
nand U2075 (N_2075,N_1674,N_1689);
nand U2076 (N_2076,N_1381,N_1643);
nand U2077 (N_2077,N_1336,N_1590);
nand U2078 (N_2078,N_1348,N_1576);
xor U2079 (N_2079,N_1769,N_1383);
nor U2080 (N_2080,N_1534,N_1755);
nand U2081 (N_2081,N_1821,N_1805);
xor U2082 (N_2082,N_1793,N_1639);
or U2083 (N_2083,N_1389,N_1390);
and U2084 (N_2084,N_1332,N_1487);
and U2085 (N_2085,N_1483,N_1659);
nand U2086 (N_2086,N_1496,N_1789);
nor U2087 (N_2087,N_1359,N_1772);
nor U2088 (N_2088,N_1634,N_1352);
xor U2089 (N_2089,N_1828,N_1724);
nand U2090 (N_2090,N_1865,N_1542);
or U2091 (N_2091,N_1273,N_1583);
nand U2092 (N_2092,N_1264,N_1356);
nor U2093 (N_2093,N_1801,N_1405);
xnor U2094 (N_2094,N_1720,N_1602);
and U2095 (N_2095,N_1740,N_1391);
or U2096 (N_2096,N_1422,N_1387);
nand U2097 (N_2097,N_1811,N_1628);
and U2098 (N_2098,N_1711,N_1458);
and U2099 (N_2099,N_1714,N_1274);
or U2100 (N_2100,N_1819,N_1777);
and U2101 (N_2101,N_1444,N_1588);
nand U2102 (N_2102,N_1603,N_1758);
xnor U2103 (N_2103,N_1855,N_1625);
xnor U2104 (N_2104,N_1402,N_1859);
xor U2105 (N_2105,N_1277,N_1790);
xnor U2106 (N_2106,N_1723,N_1702);
and U2107 (N_2107,N_1544,N_1813);
or U2108 (N_2108,N_1481,N_1715);
or U2109 (N_2109,N_1825,N_1728);
xnor U2110 (N_2110,N_1403,N_1704);
or U2111 (N_2111,N_1440,N_1360);
xnor U2112 (N_2112,N_1284,N_1770);
nor U2113 (N_2113,N_1759,N_1744);
nand U2114 (N_2114,N_1824,N_1337);
nor U2115 (N_2115,N_1493,N_1315);
nor U2116 (N_2116,N_1425,N_1608);
and U2117 (N_2117,N_1823,N_1580);
xor U2118 (N_2118,N_1596,N_1303);
or U2119 (N_2119,N_1774,N_1571);
or U2120 (N_2120,N_1584,N_1419);
or U2121 (N_2121,N_1538,N_1806);
nand U2122 (N_2122,N_1365,N_1527);
xor U2123 (N_2123,N_1377,N_1699);
nand U2124 (N_2124,N_1644,N_1548);
nor U2125 (N_2125,N_1362,N_1435);
xnor U2126 (N_2126,N_1547,N_1679);
xnor U2127 (N_2127,N_1631,N_1786);
or U2128 (N_2128,N_1466,N_1256);
xor U2129 (N_2129,N_1506,N_1486);
xnor U2130 (N_2130,N_1675,N_1735);
and U2131 (N_2131,N_1530,N_1539);
or U2132 (N_2132,N_1492,N_1629);
or U2133 (N_2133,N_1252,N_1757);
or U2134 (N_2134,N_1339,N_1672);
xnor U2135 (N_2135,N_1767,N_1350);
xnor U2136 (N_2136,N_1729,N_1618);
nor U2137 (N_2137,N_1441,N_1574);
or U2138 (N_2138,N_1765,N_1346);
nand U2139 (N_2139,N_1681,N_1251);
xor U2140 (N_2140,N_1518,N_1555);
xnor U2141 (N_2141,N_1319,N_1836);
nand U2142 (N_2142,N_1413,N_1599);
xor U2143 (N_2143,N_1872,N_1725);
xor U2144 (N_2144,N_1286,N_1614);
nand U2145 (N_2145,N_1668,N_1626);
nor U2146 (N_2146,N_1746,N_1561);
xor U2147 (N_2147,N_1385,N_1475);
nor U2148 (N_2148,N_1464,N_1364);
xor U2149 (N_2149,N_1667,N_1351);
and U2150 (N_2150,N_1254,N_1604);
or U2151 (N_2151,N_1343,N_1469);
nor U2152 (N_2152,N_1536,N_1652);
or U2153 (N_2153,N_1513,N_1673);
and U2154 (N_2154,N_1504,N_1833);
nand U2155 (N_2155,N_1700,N_1293);
nand U2156 (N_2156,N_1730,N_1386);
nand U2157 (N_2157,N_1522,N_1463);
xor U2158 (N_2158,N_1342,N_1434);
or U2159 (N_2159,N_1807,N_1703);
nor U2160 (N_2160,N_1579,N_1709);
xnor U2161 (N_2161,N_1341,N_1331);
and U2162 (N_2162,N_1779,N_1313);
xor U2163 (N_2163,N_1394,N_1857);
xnor U2164 (N_2164,N_1803,N_1338);
nor U2165 (N_2165,N_1559,N_1834);
nand U2166 (N_2166,N_1268,N_1753);
nand U2167 (N_2167,N_1306,N_1334);
nand U2168 (N_2168,N_1445,N_1829);
nor U2169 (N_2169,N_1318,N_1812);
nor U2170 (N_2170,N_1300,N_1412);
nand U2171 (N_2171,N_1601,N_1783);
xnor U2172 (N_2172,N_1418,N_1630);
or U2173 (N_2173,N_1480,N_1417);
nand U2174 (N_2174,N_1485,N_1470);
nand U2175 (N_2175,N_1818,N_1423);
or U2176 (N_2176,N_1460,N_1860);
nor U2177 (N_2177,N_1852,N_1272);
nor U2178 (N_2178,N_1335,N_1314);
nor U2179 (N_2179,N_1743,N_1736);
and U2180 (N_2180,N_1465,N_1502);
and U2181 (N_2181,N_1623,N_1764);
and U2182 (N_2182,N_1345,N_1270);
xor U2183 (N_2183,N_1666,N_1598);
or U2184 (N_2184,N_1638,N_1455);
or U2185 (N_2185,N_1844,N_1488);
or U2186 (N_2186,N_1733,N_1401);
nor U2187 (N_2187,N_1515,N_1514);
and U2188 (N_2188,N_1581,N_1644);
and U2189 (N_2189,N_1307,N_1434);
or U2190 (N_2190,N_1351,N_1383);
xnor U2191 (N_2191,N_1781,N_1556);
nand U2192 (N_2192,N_1547,N_1575);
nand U2193 (N_2193,N_1296,N_1483);
xor U2194 (N_2194,N_1380,N_1467);
nor U2195 (N_2195,N_1283,N_1672);
nor U2196 (N_2196,N_1279,N_1420);
and U2197 (N_2197,N_1867,N_1506);
nor U2198 (N_2198,N_1283,N_1433);
xnor U2199 (N_2199,N_1820,N_1310);
nand U2200 (N_2200,N_1759,N_1826);
nor U2201 (N_2201,N_1557,N_1386);
nand U2202 (N_2202,N_1275,N_1607);
nor U2203 (N_2203,N_1537,N_1298);
or U2204 (N_2204,N_1502,N_1698);
nand U2205 (N_2205,N_1325,N_1312);
xnor U2206 (N_2206,N_1425,N_1550);
or U2207 (N_2207,N_1283,N_1273);
or U2208 (N_2208,N_1690,N_1808);
and U2209 (N_2209,N_1253,N_1736);
xor U2210 (N_2210,N_1663,N_1681);
or U2211 (N_2211,N_1301,N_1735);
nand U2212 (N_2212,N_1508,N_1449);
and U2213 (N_2213,N_1267,N_1869);
nand U2214 (N_2214,N_1809,N_1340);
and U2215 (N_2215,N_1347,N_1850);
or U2216 (N_2216,N_1410,N_1632);
xor U2217 (N_2217,N_1824,N_1631);
xnor U2218 (N_2218,N_1317,N_1676);
or U2219 (N_2219,N_1592,N_1711);
xnor U2220 (N_2220,N_1645,N_1827);
nor U2221 (N_2221,N_1546,N_1629);
or U2222 (N_2222,N_1767,N_1497);
xnor U2223 (N_2223,N_1475,N_1411);
xnor U2224 (N_2224,N_1581,N_1870);
or U2225 (N_2225,N_1675,N_1416);
and U2226 (N_2226,N_1748,N_1831);
nor U2227 (N_2227,N_1734,N_1396);
nor U2228 (N_2228,N_1410,N_1431);
nor U2229 (N_2229,N_1602,N_1694);
nor U2230 (N_2230,N_1308,N_1256);
or U2231 (N_2231,N_1461,N_1524);
or U2232 (N_2232,N_1686,N_1685);
nand U2233 (N_2233,N_1475,N_1593);
nor U2234 (N_2234,N_1745,N_1706);
nor U2235 (N_2235,N_1808,N_1559);
xor U2236 (N_2236,N_1504,N_1643);
xor U2237 (N_2237,N_1560,N_1378);
nor U2238 (N_2238,N_1816,N_1854);
nand U2239 (N_2239,N_1334,N_1689);
and U2240 (N_2240,N_1520,N_1375);
xnor U2241 (N_2241,N_1479,N_1522);
xor U2242 (N_2242,N_1715,N_1774);
nand U2243 (N_2243,N_1302,N_1770);
nor U2244 (N_2244,N_1678,N_1504);
nand U2245 (N_2245,N_1835,N_1689);
xnor U2246 (N_2246,N_1559,N_1869);
nand U2247 (N_2247,N_1616,N_1284);
xor U2248 (N_2248,N_1423,N_1793);
nor U2249 (N_2249,N_1277,N_1278);
or U2250 (N_2250,N_1848,N_1713);
xor U2251 (N_2251,N_1547,N_1614);
and U2252 (N_2252,N_1408,N_1821);
or U2253 (N_2253,N_1614,N_1528);
xor U2254 (N_2254,N_1437,N_1363);
nor U2255 (N_2255,N_1785,N_1643);
xor U2256 (N_2256,N_1253,N_1601);
nor U2257 (N_2257,N_1389,N_1829);
and U2258 (N_2258,N_1701,N_1837);
or U2259 (N_2259,N_1462,N_1608);
nor U2260 (N_2260,N_1408,N_1478);
or U2261 (N_2261,N_1501,N_1864);
nor U2262 (N_2262,N_1275,N_1730);
and U2263 (N_2263,N_1743,N_1365);
xnor U2264 (N_2264,N_1402,N_1663);
xnor U2265 (N_2265,N_1636,N_1284);
or U2266 (N_2266,N_1550,N_1668);
nand U2267 (N_2267,N_1387,N_1643);
xnor U2268 (N_2268,N_1587,N_1719);
and U2269 (N_2269,N_1369,N_1253);
and U2270 (N_2270,N_1726,N_1781);
xor U2271 (N_2271,N_1646,N_1335);
nor U2272 (N_2272,N_1856,N_1475);
nand U2273 (N_2273,N_1668,N_1836);
nand U2274 (N_2274,N_1850,N_1771);
nor U2275 (N_2275,N_1813,N_1588);
xor U2276 (N_2276,N_1250,N_1608);
nor U2277 (N_2277,N_1814,N_1520);
nand U2278 (N_2278,N_1345,N_1657);
nor U2279 (N_2279,N_1842,N_1736);
xnor U2280 (N_2280,N_1470,N_1625);
xnor U2281 (N_2281,N_1813,N_1549);
and U2282 (N_2282,N_1838,N_1529);
nor U2283 (N_2283,N_1438,N_1858);
and U2284 (N_2284,N_1631,N_1699);
and U2285 (N_2285,N_1766,N_1561);
nor U2286 (N_2286,N_1254,N_1735);
or U2287 (N_2287,N_1663,N_1839);
and U2288 (N_2288,N_1671,N_1721);
nand U2289 (N_2289,N_1643,N_1558);
xor U2290 (N_2290,N_1714,N_1597);
and U2291 (N_2291,N_1318,N_1343);
nand U2292 (N_2292,N_1751,N_1331);
or U2293 (N_2293,N_1560,N_1699);
nor U2294 (N_2294,N_1397,N_1278);
and U2295 (N_2295,N_1516,N_1512);
nand U2296 (N_2296,N_1509,N_1620);
xor U2297 (N_2297,N_1824,N_1813);
xnor U2298 (N_2298,N_1821,N_1831);
nor U2299 (N_2299,N_1863,N_1448);
or U2300 (N_2300,N_1542,N_1336);
or U2301 (N_2301,N_1311,N_1771);
and U2302 (N_2302,N_1511,N_1493);
xnor U2303 (N_2303,N_1700,N_1722);
or U2304 (N_2304,N_1474,N_1271);
nor U2305 (N_2305,N_1421,N_1831);
and U2306 (N_2306,N_1777,N_1563);
and U2307 (N_2307,N_1767,N_1368);
xnor U2308 (N_2308,N_1656,N_1764);
or U2309 (N_2309,N_1327,N_1868);
and U2310 (N_2310,N_1846,N_1448);
or U2311 (N_2311,N_1676,N_1727);
xnor U2312 (N_2312,N_1586,N_1258);
xor U2313 (N_2313,N_1774,N_1491);
nor U2314 (N_2314,N_1699,N_1255);
nand U2315 (N_2315,N_1443,N_1838);
nand U2316 (N_2316,N_1695,N_1627);
xor U2317 (N_2317,N_1636,N_1667);
xnor U2318 (N_2318,N_1623,N_1300);
nor U2319 (N_2319,N_1862,N_1411);
nor U2320 (N_2320,N_1272,N_1764);
or U2321 (N_2321,N_1796,N_1601);
or U2322 (N_2322,N_1656,N_1532);
xor U2323 (N_2323,N_1588,N_1811);
nand U2324 (N_2324,N_1359,N_1542);
nor U2325 (N_2325,N_1688,N_1456);
and U2326 (N_2326,N_1754,N_1866);
nor U2327 (N_2327,N_1387,N_1310);
or U2328 (N_2328,N_1275,N_1556);
and U2329 (N_2329,N_1558,N_1428);
nor U2330 (N_2330,N_1641,N_1466);
and U2331 (N_2331,N_1669,N_1862);
xor U2332 (N_2332,N_1332,N_1442);
nor U2333 (N_2333,N_1663,N_1396);
or U2334 (N_2334,N_1436,N_1799);
and U2335 (N_2335,N_1374,N_1571);
and U2336 (N_2336,N_1427,N_1395);
nor U2337 (N_2337,N_1415,N_1514);
and U2338 (N_2338,N_1554,N_1366);
or U2339 (N_2339,N_1453,N_1551);
nand U2340 (N_2340,N_1417,N_1782);
xnor U2341 (N_2341,N_1661,N_1549);
nand U2342 (N_2342,N_1872,N_1669);
nor U2343 (N_2343,N_1424,N_1540);
xnor U2344 (N_2344,N_1719,N_1605);
or U2345 (N_2345,N_1789,N_1515);
or U2346 (N_2346,N_1567,N_1287);
nor U2347 (N_2347,N_1747,N_1745);
nor U2348 (N_2348,N_1554,N_1531);
and U2349 (N_2349,N_1605,N_1599);
or U2350 (N_2350,N_1354,N_1720);
xnor U2351 (N_2351,N_1639,N_1513);
xor U2352 (N_2352,N_1550,N_1543);
xor U2353 (N_2353,N_1869,N_1397);
or U2354 (N_2354,N_1660,N_1563);
or U2355 (N_2355,N_1614,N_1595);
xor U2356 (N_2356,N_1412,N_1801);
or U2357 (N_2357,N_1736,N_1614);
nor U2358 (N_2358,N_1665,N_1832);
xor U2359 (N_2359,N_1816,N_1815);
and U2360 (N_2360,N_1403,N_1736);
nand U2361 (N_2361,N_1572,N_1448);
xor U2362 (N_2362,N_1562,N_1515);
nand U2363 (N_2363,N_1496,N_1464);
xnor U2364 (N_2364,N_1801,N_1657);
nand U2365 (N_2365,N_1487,N_1706);
nand U2366 (N_2366,N_1537,N_1492);
and U2367 (N_2367,N_1502,N_1357);
and U2368 (N_2368,N_1263,N_1660);
xor U2369 (N_2369,N_1514,N_1826);
or U2370 (N_2370,N_1420,N_1726);
xor U2371 (N_2371,N_1399,N_1432);
or U2372 (N_2372,N_1732,N_1874);
nand U2373 (N_2373,N_1651,N_1694);
xnor U2374 (N_2374,N_1329,N_1370);
and U2375 (N_2375,N_1771,N_1737);
and U2376 (N_2376,N_1480,N_1353);
nand U2377 (N_2377,N_1625,N_1824);
nor U2378 (N_2378,N_1485,N_1530);
or U2379 (N_2379,N_1486,N_1528);
or U2380 (N_2380,N_1696,N_1565);
xnor U2381 (N_2381,N_1791,N_1699);
and U2382 (N_2382,N_1717,N_1738);
nand U2383 (N_2383,N_1421,N_1738);
nand U2384 (N_2384,N_1772,N_1707);
xor U2385 (N_2385,N_1380,N_1290);
or U2386 (N_2386,N_1302,N_1270);
nand U2387 (N_2387,N_1851,N_1786);
nor U2388 (N_2388,N_1406,N_1680);
xnor U2389 (N_2389,N_1647,N_1480);
xor U2390 (N_2390,N_1286,N_1320);
nor U2391 (N_2391,N_1638,N_1815);
xnor U2392 (N_2392,N_1407,N_1744);
and U2393 (N_2393,N_1676,N_1594);
xnor U2394 (N_2394,N_1337,N_1301);
and U2395 (N_2395,N_1362,N_1720);
or U2396 (N_2396,N_1703,N_1599);
and U2397 (N_2397,N_1579,N_1799);
xor U2398 (N_2398,N_1817,N_1334);
xor U2399 (N_2399,N_1554,N_1385);
xor U2400 (N_2400,N_1872,N_1469);
nand U2401 (N_2401,N_1594,N_1711);
nor U2402 (N_2402,N_1359,N_1591);
or U2403 (N_2403,N_1811,N_1352);
xnor U2404 (N_2404,N_1704,N_1317);
xnor U2405 (N_2405,N_1505,N_1288);
or U2406 (N_2406,N_1873,N_1430);
nand U2407 (N_2407,N_1373,N_1722);
or U2408 (N_2408,N_1400,N_1453);
nand U2409 (N_2409,N_1552,N_1854);
xnor U2410 (N_2410,N_1849,N_1490);
xnor U2411 (N_2411,N_1332,N_1580);
and U2412 (N_2412,N_1514,N_1479);
xor U2413 (N_2413,N_1494,N_1301);
nor U2414 (N_2414,N_1873,N_1331);
nand U2415 (N_2415,N_1797,N_1487);
nor U2416 (N_2416,N_1680,N_1350);
xnor U2417 (N_2417,N_1597,N_1859);
nor U2418 (N_2418,N_1801,N_1793);
nor U2419 (N_2419,N_1793,N_1757);
nand U2420 (N_2420,N_1467,N_1611);
nand U2421 (N_2421,N_1424,N_1331);
or U2422 (N_2422,N_1637,N_1733);
and U2423 (N_2423,N_1494,N_1284);
and U2424 (N_2424,N_1345,N_1393);
and U2425 (N_2425,N_1467,N_1617);
and U2426 (N_2426,N_1415,N_1681);
or U2427 (N_2427,N_1626,N_1251);
nor U2428 (N_2428,N_1734,N_1376);
and U2429 (N_2429,N_1477,N_1394);
nand U2430 (N_2430,N_1446,N_1856);
or U2431 (N_2431,N_1462,N_1645);
xnor U2432 (N_2432,N_1483,N_1821);
nand U2433 (N_2433,N_1798,N_1430);
nand U2434 (N_2434,N_1683,N_1668);
and U2435 (N_2435,N_1421,N_1627);
xnor U2436 (N_2436,N_1826,N_1822);
xnor U2437 (N_2437,N_1524,N_1680);
nand U2438 (N_2438,N_1700,N_1866);
xor U2439 (N_2439,N_1368,N_1354);
nor U2440 (N_2440,N_1570,N_1548);
or U2441 (N_2441,N_1298,N_1528);
or U2442 (N_2442,N_1410,N_1323);
and U2443 (N_2443,N_1276,N_1539);
and U2444 (N_2444,N_1645,N_1293);
nor U2445 (N_2445,N_1698,N_1542);
xor U2446 (N_2446,N_1311,N_1637);
xnor U2447 (N_2447,N_1797,N_1692);
and U2448 (N_2448,N_1395,N_1455);
nor U2449 (N_2449,N_1431,N_1396);
or U2450 (N_2450,N_1836,N_1371);
xor U2451 (N_2451,N_1343,N_1345);
nor U2452 (N_2452,N_1587,N_1503);
or U2453 (N_2453,N_1406,N_1425);
or U2454 (N_2454,N_1298,N_1495);
and U2455 (N_2455,N_1641,N_1824);
xor U2456 (N_2456,N_1575,N_1496);
and U2457 (N_2457,N_1362,N_1367);
nor U2458 (N_2458,N_1841,N_1581);
nor U2459 (N_2459,N_1847,N_1355);
or U2460 (N_2460,N_1708,N_1609);
nor U2461 (N_2461,N_1529,N_1656);
xnor U2462 (N_2462,N_1844,N_1337);
and U2463 (N_2463,N_1691,N_1351);
and U2464 (N_2464,N_1386,N_1412);
xnor U2465 (N_2465,N_1556,N_1571);
nor U2466 (N_2466,N_1429,N_1750);
xor U2467 (N_2467,N_1519,N_1798);
and U2468 (N_2468,N_1539,N_1413);
or U2469 (N_2469,N_1732,N_1258);
or U2470 (N_2470,N_1720,N_1532);
xor U2471 (N_2471,N_1657,N_1692);
and U2472 (N_2472,N_1642,N_1621);
and U2473 (N_2473,N_1521,N_1252);
or U2474 (N_2474,N_1452,N_1527);
or U2475 (N_2475,N_1609,N_1327);
xor U2476 (N_2476,N_1353,N_1348);
nor U2477 (N_2477,N_1361,N_1390);
and U2478 (N_2478,N_1321,N_1421);
nor U2479 (N_2479,N_1331,N_1660);
or U2480 (N_2480,N_1295,N_1577);
or U2481 (N_2481,N_1829,N_1335);
or U2482 (N_2482,N_1654,N_1828);
xor U2483 (N_2483,N_1784,N_1738);
xor U2484 (N_2484,N_1422,N_1655);
xnor U2485 (N_2485,N_1779,N_1516);
and U2486 (N_2486,N_1302,N_1283);
nand U2487 (N_2487,N_1595,N_1767);
nand U2488 (N_2488,N_1379,N_1796);
nor U2489 (N_2489,N_1287,N_1751);
nor U2490 (N_2490,N_1461,N_1479);
or U2491 (N_2491,N_1587,N_1675);
or U2492 (N_2492,N_1641,N_1843);
nor U2493 (N_2493,N_1450,N_1684);
nor U2494 (N_2494,N_1334,N_1393);
and U2495 (N_2495,N_1341,N_1457);
nand U2496 (N_2496,N_1752,N_1821);
nor U2497 (N_2497,N_1697,N_1624);
nor U2498 (N_2498,N_1868,N_1634);
nand U2499 (N_2499,N_1409,N_1435);
nand U2500 (N_2500,N_1928,N_2151);
nand U2501 (N_2501,N_2141,N_1979);
nor U2502 (N_2502,N_2128,N_2467);
and U2503 (N_2503,N_2180,N_1876);
xnor U2504 (N_2504,N_2013,N_2118);
nand U2505 (N_2505,N_1887,N_2428);
nor U2506 (N_2506,N_2033,N_2014);
nand U2507 (N_2507,N_1878,N_1888);
or U2508 (N_2508,N_2086,N_2288);
nand U2509 (N_2509,N_1918,N_2370);
and U2510 (N_2510,N_2201,N_2134);
xor U2511 (N_2511,N_2457,N_1974);
and U2512 (N_2512,N_1972,N_2373);
or U2513 (N_2513,N_1892,N_2414);
nor U2514 (N_2514,N_2055,N_2101);
xor U2515 (N_2515,N_2442,N_2439);
and U2516 (N_2516,N_2179,N_2406);
and U2517 (N_2517,N_1963,N_2483);
nor U2518 (N_2518,N_1895,N_1916);
or U2519 (N_2519,N_2224,N_1880);
xnor U2520 (N_2520,N_2066,N_2408);
nand U2521 (N_2521,N_2424,N_2072);
and U2522 (N_2522,N_1894,N_2423);
nand U2523 (N_2523,N_2181,N_1884);
or U2524 (N_2524,N_2355,N_2000);
or U2525 (N_2525,N_2311,N_1975);
and U2526 (N_2526,N_1898,N_1993);
or U2527 (N_2527,N_2427,N_2052);
and U2528 (N_2528,N_2475,N_2229);
or U2529 (N_2529,N_1981,N_2167);
or U2530 (N_2530,N_2160,N_2271);
xnor U2531 (N_2531,N_2473,N_2460);
or U2532 (N_2532,N_2076,N_1966);
nand U2533 (N_2533,N_1907,N_2144);
nand U2534 (N_2534,N_2148,N_2218);
xnor U2535 (N_2535,N_2105,N_2253);
nor U2536 (N_2536,N_2312,N_1978);
or U2537 (N_2537,N_2278,N_2178);
nor U2538 (N_2538,N_2411,N_2327);
and U2539 (N_2539,N_2074,N_2447);
nor U2540 (N_2540,N_1909,N_2410);
or U2541 (N_2541,N_2137,N_2195);
and U2542 (N_2542,N_2097,N_2333);
or U2543 (N_2543,N_1930,N_2315);
nand U2544 (N_2544,N_2497,N_2035);
xor U2545 (N_2545,N_2202,N_2413);
nand U2546 (N_2546,N_2003,N_2368);
nor U2547 (N_2547,N_2028,N_2234);
xor U2548 (N_2548,N_2479,N_2356);
and U2549 (N_2549,N_2015,N_2210);
nand U2550 (N_2550,N_2170,N_2245);
or U2551 (N_2551,N_2319,N_2383);
nand U2552 (N_2552,N_2317,N_2109);
nand U2553 (N_2553,N_2166,N_2081);
nor U2554 (N_2554,N_2030,N_1990);
or U2555 (N_2555,N_2261,N_2477);
xor U2556 (N_2556,N_2269,N_2274);
and U2557 (N_2557,N_2207,N_2173);
or U2558 (N_2558,N_2126,N_2443);
or U2559 (N_2559,N_2495,N_2259);
and U2560 (N_2560,N_2197,N_2045);
or U2561 (N_2561,N_2132,N_2082);
xor U2562 (N_2562,N_2029,N_2021);
and U2563 (N_2563,N_2283,N_1905);
nand U2564 (N_2564,N_2272,N_2092);
and U2565 (N_2565,N_2068,N_2380);
nand U2566 (N_2566,N_2049,N_2051);
and U2567 (N_2567,N_2250,N_2042);
or U2568 (N_2568,N_2230,N_2268);
xor U2569 (N_2569,N_2194,N_2484);
and U2570 (N_2570,N_2114,N_2240);
nor U2571 (N_2571,N_2330,N_2139);
and U2572 (N_2572,N_1908,N_2112);
nand U2573 (N_2573,N_2256,N_2418);
nor U2574 (N_2574,N_2110,N_2407);
and U2575 (N_2575,N_2270,N_2405);
and U2576 (N_2576,N_1915,N_2184);
nand U2577 (N_2577,N_2307,N_2306);
nand U2578 (N_2578,N_2249,N_1951);
or U2579 (N_2579,N_1931,N_2205);
and U2580 (N_2580,N_2353,N_1935);
or U2581 (N_2581,N_2108,N_2191);
nor U2582 (N_2582,N_2438,N_2059);
nor U2583 (N_2583,N_2212,N_2192);
or U2584 (N_2584,N_1970,N_2449);
nand U2585 (N_2585,N_2220,N_2378);
nor U2586 (N_2586,N_2396,N_1983);
and U2587 (N_2587,N_1943,N_2446);
or U2588 (N_2588,N_1954,N_1911);
and U2589 (N_2589,N_2369,N_2285);
nand U2590 (N_2590,N_2247,N_2417);
nor U2591 (N_2591,N_2064,N_2496);
nand U2592 (N_2592,N_2119,N_2236);
or U2593 (N_2593,N_2102,N_2208);
and U2594 (N_2594,N_2083,N_2206);
and U2595 (N_2595,N_2241,N_2388);
or U2596 (N_2596,N_2481,N_2214);
xor U2597 (N_2597,N_2279,N_2031);
nor U2598 (N_2598,N_2493,N_2142);
nand U2599 (N_2599,N_1960,N_1988);
nand U2600 (N_2600,N_2222,N_2290);
xnor U2601 (N_2601,N_2155,N_2273);
nor U2602 (N_2602,N_2093,N_2337);
nor U2603 (N_2603,N_2041,N_2252);
nand U2604 (N_2604,N_2070,N_1901);
or U2605 (N_2605,N_1929,N_2091);
xnor U2606 (N_2606,N_1937,N_2100);
or U2607 (N_2607,N_1881,N_1940);
or U2608 (N_2608,N_2024,N_2131);
xnor U2609 (N_2609,N_2164,N_1999);
xor U2610 (N_2610,N_1923,N_2060);
and U2611 (N_2611,N_2302,N_2352);
and U2612 (N_2612,N_2482,N_2303);
and U2613 (N_2613,N_2043,N_2019);
nand U2614 (N_2614,N_1984,N_2080);
and U2615 (N_2615,N_2163,N_2329);
nand U2616 (N_2616,N_1998,N_2006);
nor U2617 (N_2617,N_2403,N_2275);
and U2618 (N_2618,N_2498,N_2153);
or U2619 (N_2619,N_2314,N_2172);
xor U2620 (N_2620,N_2300,N_2350);
or U2621 (N_2621,N_2186,N_2204);
or U2622 (N_2622,N_2088,N_2198);
nand U2623 (N_2623,N_1921,N_1939);
or U2624 (N_2624,N_1936,N_1977);
nand U2625 (N_2625,N_1971,N_2298);
nand U2626 (N_2626,N_1958,N_2200);
or U2627 (N_2627,N_1945,N_2171);
or U2628 (N_2628,N_1961,N_2152);
or U2629 (N_2629,N_2010,N_2293);
and U2630 (N_2630,N_2099,N_2254);
xnor U2631 (N_2631,N_2367,N_2140);
nor U2632 (N_2632,N_2382,N_2359);
and U2633 (N_2633,N_2436,N_2239);
xnor U2634 (N_2634,N_2340,N_1980);
nand U2635 (N_2635,N_2426,N_2287);
or U2636 (N_2636,N_2044,N_1885);
xnor U2637 (N_2637,N_1956,N_2089);
xnor U2638 (N_2638,N_2429,N_1946);
nor U2639 (N_2639,N_2313,N_1897);
and U2640 (N_2640,N_2103,N_2494);
nor U2641 (N_2641,N_2113,N_2299);
nor U2642 (N_2642,N_2096,N_1917);
xnor U2643 (N_2643,N_2161,N_2464);
xor U2644 (N_2644,N_1889,N_2393);
and U2645 (N_2645,N_2231,N_2162);
xnor U2646 (N_2646,N_2296,N_2223);
nor U2647 (N_2647,N_2156,N_2491);
and U2648 (N_2648,N_2468,N_2372);
and U2649 (N_2649,N_2478,N_1882);
nor U2650 (N_2650,N_1982,N_2343);
xnor U2651 (N_2651,N_2430,N_1969);
nand U2652 (N_2652,N_2216,N_2437);
and U2653 (N_2653,N_2005,N_1950);
xor U2654 (N_2654,N_2242,N_2445);
nand U2655 (N_2655,N_2190,N_2384);
nor U2656 (N_2656,N_2122,N_2415);
and U2657 (N_2657,N_2090,N_2264);
and U2658 (N_2658,N_1959,N_2219);
nor U2659 (N_2659,N_2281,N_2387);
or U2660 (N_2660,N_2169,N_1987);
xnor U2661 (N_2661,N_1891,N_2098);
nand U2662 (N_2662,N_1913,N_2360);
nor U2663 (N_2663,N_2046,N_1991);
or U2664 (N_2664,N_2276,N_1944);
nor U2665 (N_2665,N_2036,N_2196);
and U2666 (N_2666,N_2133,N_2316);
nor U2667 (N_2667,N_2463,N_2107);
nor U2668 (N_2668,N_2130,N_2432);
xor U2669 (N_2669,N_2398,N_1957);
and U2670 (N_2670,N_2165,N_2363);
nor U2671 (N_2671,N_2129,N_2348);
nand U2672 (N_2672,N_2004,N_1900);
nor U2673 (N_2673,N_2402,N_2435);
xor U2674 (N_2674,N_2053,N_2379);
nand U2675 (N_2675,N_2087,N_2255);
nand U2676 (N_2676,N_2357,N_1906);
xnor U2677 (N_2677,N_2025,N_2111);
nand U2678 (N_2678,N_2094,N_2489);
xor U2679 (N_2679,N_2002,N_2048);
xor U2680 (N_2680,N_1886,N_2323);
xnor U2681 (N_2681,N_2263,N_2347);
nand U2682 (N_2682,N_2412,N_2084);
or U2683 (N_2683,N_2326,N_2400);
nand U2684 (N_2684,N_2331,N_1997);
and U2685 (N_2685,N_1992,N_2085);
and U2686 (N_2686,N_2027,N_1903);
nor U2687 (N_2687,N_2469,N_2039);
nand U2688 (N_2688,N_2017,N_1942);
xor U2689 (N_2689,N_2282,N_2462);
or U2690 (N_2690,N_2433,N_1962);
nand U2691 (N_2691,N_2374,N_2095);
nor U2692 (N_2692,N_2174,N_2375);
and U2693 (N_2693,N_1904,N_2257);
xor U2694 (N_2694,N_2221,N_1965);
xnor U2695 (N_2695,N_2371,N_1976);
xnor U2696 (N_2696,N_1947,N_2354);
nor U2697 (N_2697,N_2452,N_1922);
or U2698 (N_2698,N_2203,N_2136);
and U2699 (N_2699,N_1964,N_2310);
xor U2700 (N_2700,N_2168,N_2286);
nor U2701 (N_2701,N_2381,N_2104);
or U2702 (N_2702,N_2365,N_2425);
xnor U2703 (N_2703,N_2305,N_2488);
nor U2704 (N_2704,N_2386,N_2016);
xnor U2705 (N_2705,N_2007,N_1985);
xnor U2706 (N_2706,N_2078,N_2459);
xor U2707 (N_2707,N_2244,N_2358);
xor U2708 (N_2708,N_2487,N_2232);
and U2709 (N_2709,N_1899,N_2260);
and U2710 (N_2710,N_2038,N_2040);
nor U2711 (N_2711,N_2309,N_2001);
nand U2712 (N_2712,N_2338,N_2154);
or U2713 (N_2713,N_2177,N_1994);
xor U2714 (N_2714,N_1890,N_2434);
or U2715 (N_2715,N_2009,N_2146);
xor U2716 (N_2716,N_2420,N_1967);
xnor U2717 (N_2717,N_1925,N_2486);
or U2718 (N_2718,N_2235,N_1932);
nor U2719 (N_2719,N_2292,N_2441);
and U2720 (N_2720,N_2377,N_2193);
xor U2721 (N_2721,N_2077,N_2409);
xnor U2722 (N_2722,N_1989,N_2349);
and U2723 (N_2723,N_2472,N_1941);
nor U2724 (N_2724,N_2280,N_1927);
xor U2725 (N_2725,N_2320,N_2318);
or U2726 (N_2726,N_2061,N_2490);
xor U2727 (N_2727,N_2054,N_2440);
nand U2728 (N_2728,N_2183,N_2277);
or U2729 (N_2729,N_1896,N_2233);
nand U2730 (N_2730,N_2116,N_2150);
and U2731 (N_2731,N_2421,N_2149);
nor U2732 (N_2732,N_1919,N_2453);
or U2733 (N_2733,N_1996,N_1914);
xnor U2734 (N_2734,N_1973,N_2262);
or U2735 (N_2735,N_2401,N_2125);
nand U2736 (N_2736,N_2390,N_1893);
and U2737 (N_2737,N_2158,N_2325);
or U2738 (N_2738,N_2215,N_2011);
or U2739 (N_2739,N_1910,N_2332);
xor U2740 (N_2740,N_2243,N_2079);
and U2741 (N_2741,N_2361,N_2335);
xor U2742 (N_2742,N_2385,N_2022);
nand U2743 (N_2743,N_2344,N_1953);
nor U2744 (N_2744,N_2291,N_2456);
xnor U2745 (N_2745,N_2265,N_2336);
xnor U2746 (N_2746,N_2366,N_2056);
nor U2747 (N_2747,N_2461,N_1926);
and U2748 (N_2748,N_2322,N_2444);
or U2749 (N_2749,N_1948,N_2227);
or U2750 (N_2750,N_2284,N_2023);
nand U2751 (N_2751,N_1938,N_2238);
and U2752 (N_2752,N_2115,N_2419);
nor U2753 (N_2753,N_2159,N_2334);
nor U2754 (N_2754,N_2058,N_2188);
or U2755 (N_2755,N_2189,N_2034);
or U2756 (N_2756,N_2211,N_2182);
xor U2757 (N_2757,N_2145,N_1995);
xnor U2758 (N_2758,N_2339,N_2289);
and U2759 (N_2759,N_2012,N_2185);
nor U2760 (N_2760,N_2450,N_2364);
or U2761 (N_2761,N_2328,N_2321);
nor U2762 (N_2762,N_1955,N_2431);
nor U2763 (N_2763,N_2213,N_1986);
nand U2764 (N_2764,N_2251,N_2106);
xnor U2765 (N_2765,N_2397,N_2127);
or U2766 (N_2766,N_2448,N_2217);
and U2767 (N_2767,N_2399,N_2458);
or U2768 (N_2768,N_2020,N_2075);
nand U2769 (N_2769,N_2047,N_1933);
nand U2770 (N_2770,N_2304,N_2237);
nand U2771 (N_2771,N_2451,N_2258);
and U2772 (N_2772,N_2228,N_2492);
and U2773 (N_2773,N_1883,N_1924);
nor U2774 (N_2774,N_2404,N_2480);
and U2775 (N_2775,N_2341,N_2135);
and U2776 (N_2776,N_2138,N_2123);
nand U2777 (N_2777,N_2121,N_2465);
or U2778 (N_2778,N_2324,N_2226);
nor U2779 (N_2779,N_2471,N_2362);
or U2780 (N_2780,N_2037,N_2209);
and U2781 (N_2781,N_2225,N_1902);
nor U2782 (N_2782,N_2267,N_2476);
nand U2783 (N_2783,N_2147,N_2474);
nand U2784 (N_2784,N_2065,N_2067);
and U2785 (N_2785,N_2301,N_2143);
or U2786 (N_2786,N_2470,N_2485);
or U2787 (N_2787,N_2050,N_2308);
and U2788 (N_2788,N_2394,N_2294);
nand U2789 (N_2789,N_2032,N_2455);
nor U2790 (N_2790,N_2351,N_1920);
nand U2791 (N_2791,N_2454,N_2416);
or U2792 (N_2792,N_2062,N_2346);
or U2793 (N_2793,N_2422,N_2392);
nand U2794 (N_2794,N_2187,N_2295);
nor U2795 (N_2795,N_2073,N_2026);
nor U2796 (N_2796,N_1875,N_1952);
and U2797 (N_2797,N_2008,N_2246);
or U2798 (N_2798,N_2124,N_2499);
and U2799 (N_2799,N_2345,N_1912);
or U2800 (N_2800,N_2063,N_2176);
xnor U2801 (N_2801,N_2266,N_2395);
xnor U2802 (N_2802,N_2248,N_2376);
or U2803 (N_2803,N_1949,N_2120);
xnor U2804 (N_2804,N_1934,N_2069);
nand U2805 (N_2805,N_2297,N_1879);
nand U2806 (N_2806,N_2117,N_1968);
or U2807 (N_2807,N_2018,N_2391);
and U2808 (N_2808,N_1877,N_2071);
and U2809 (N_2809,N_2466,N_2175);
xor U2810 (N_2810,N_2057,N_2342);
xnor U2811 (N_2811,N_2157,N_2199);
nor U2812 (N_2812,N_2389,N_2388);
and U2813 (N_2813,N_2413,N_2463);
xnor U2814 (N_2814,N_2235,N_2170);
and U2815 (N_2815,N_2105,N_2404);
or U2816 (N_2816,N_2476,N_2132);
nor U2817 (N_2817,N_2241,N_2037);
nand U2818 (N_2818,N_2469,N_1892);
nor U2819 (N_2819,N_2039,N_2225);
or U2820 (N_2820,N_2247,N_2036);
nand U2821 (N_2821,N_2420,N_2157);
nor U2822 (N_2822,N_2214,N_2117);
and U2823 (N_2823,N_2240,N_2479);
xnor U2824 (N_2824,N_2471,N_2026);
or U2825 (N_2825,N_2193,N_2125);
xnor U2826 (N_2826,N_2435,N_2376);
nand U2827 (N_2827,N_1970,N_2459);
nand U2828 (N_2828,N_2106,N_2434);
xor U2829 (N_2829,N_2406,N_1899);
or U2830 (N_2830,N_1971,N_1932);
or U2831 (N_2831,N_2211,N_2069);
or U2832 (N_2832,N_2247,N_2254);
and U2833 (N_2833,N_1889,N_2327);
or U2834 (N_2834,N_2240,N_2000);
nand U2835 (N_2835,N_2024,N_2034);
nand U2836 (N_2836,N_2003,N_1979);
nand U2837 (N_2837,N_2089,N_2025);
nand U2838 (N_2838,N_2051,N_2176);
or U2839 (N_2839,N_2290,N_2140);
or U2840 (N_2840,N_2183,N_2064);
nor U2841 (N_2841,N_2443,N_2375);
or U2842 (N_2842,N_2161,N_2398);
or U2843 (N_2843,N_2465,N_1996);
nor U2844 (N_2844,N_2294,N_2367);
nand U2845 (N_2845,N_2246,N_2236);
nand U2846 (N_2846,N_2302,N_2279);
nor U2847 (N_2847,N_2055,N_2398);
xor U2848 (N_2848,N_2460,N_1885);
nand U2849 (N_2849,N_2139,N_2087);
nand U2850 (N_2850,N_2114,N_1936);
xor U2851 (N_2851,N_1878,N_2376);
nand U2852 (N_2852,N_1896,N_2073);
and U2853 (N_2853,N_2084,N_1990);
nor U2854 (N_2854,N_2272,N_2070);
nand U2855 (N_2855,N_2221,N_2271);
or U2856 (N_2856,N_2333,N_2297);
or U2857 (N_2857,N_2075,N_2205);
nand U2858 (N_2858,N_1936,N_2079);
or U2859 (N_2859,N_2473,N_2285);
xnor U2860 (N_2860,N_2064,N_2424);
nand U2861 (N_2861,N_1891,N_2024);
nand U2862 (N_2862,N_2048,N_1992);
and U2863 (N_2863,N_2331,N_2319);
nor U2864 (N_2864,N_2168,N_2022);
nand U2865 (N_2865,N_2063,N_2334);
and U2866 (N_2866,N_1960,N_2141);
xor U2867 (N_2867,N_2049,N_2304);
xor U2868 (N_2868,N_1919,N_1921);
nand U2869 (N_2869,N_2188,N_2199);
nand U2870 (N_2870,N_2193,N_2038);
xor U2871 (N_2871,N_2110,N_1937);
nor U2872 (N_2872,N_2061,N_1955);
and U2873 (N_2873,N_2334,N_1972);
or U2874 (N_2874,N_2354,N_2307);
or U2875 (N_2875,N_2469,N_2157);
or U2876 (N_2876,N_2379,N_2475);
nand U2877 (N_2877,N_2304,N_2088);
nand U2878 (N_2878,N_2240,N_2191);
nor U2879 (N_2879,N_1956,N_2387);
xor U2880 (N_2880,N_2328,N_2355);
or U2881 (N_2881,N_2069,N_2454);
xor U2882 (N_2882,N_2000,N_2209);
xnor U2883 (N_2883,N_2173,N_2323);
nor U2884 (N_2884,N_2064,N_2258);
nor U2885 (N_2885,N_2332,N_2197);
and U2886 (N_2886,N_2105,N_2373);
nor U2887 (N_2887,N_2189,N_2146);
xnor U2888 (N_2888,N_2025,N_2236);
xor U2889 (N_2889,N_2472,N_2416);
nor U2890 (N_2890,N_1988,N_2429);
and U2891 (N_2891,N_2128,N_2064);
and U2892 (N_2892,N_2224,N_1952);
and U2893 (N_2893,N_2081,N_2438);
and U2894 (N_2894,N_2341,N_2142);
xnor U2895 (N_2895,N_2235,N_2126);
xnor U2896 (N_2896,N_2279,N_2112);
nor U2897 (N_2897,N_2279,N_2320);
and U2898 (N_2898,N_2356,N_2439);
nand U2899 (N_2899,N_2442,N_2138);
and U2900 (N_2900,N_2197,N_2314);
and U2901 (N_2901,N_2054,N_2334);
or U2902 (N_2902,N_2344,N_2160);
nor U2903 (N_2903,N_1906,N_2400);
and U2904 (N_2904,N_1939,N_2271);
nand U2905 (N_2905,N_1967,N_2484);
and U2906 (N_2906,N_2246,N_2497);
and U2907 (N_2907,N_2481,N_2142);
and U2908 (N_2908,N_1915,N_1966);
and U2909 (N_2909,N_2484,N_1880);
or U2910 (N_2910,N_2401,N_2033);
and U2911 (N_2911,N_1905,N_1985);
xor U2912 (N_2912,N_2115,N_2024);
xor U2913 (N_2913,N_2045,N_1984);
or U2914 (N_2914,N_2392,N_2144);
xnor U2915 (N_2915,N_2353,N_2168);
nor U2916 (N_2916,N_2257,N_2305);
and U2917 (N_2917,N_1960,N_2171);
nor U2918 (N_2918,N_1986,N_2263);
xor U2919 (N_2919,N_2326,N_2497);
xnor U2920 (N_2920,N_2342,N_2279);
xnor U2921 (N_2921,N_2053,N_2099);
xor U2922 (N_2922,N_2354,N_1945);
xor U2923 (N_2923,N_2192,N_2283);
and U2924 (N_2924,N_2233,N_2184);
xor U2925 (N_2925,N_2354,N_2076);
xor U2926 (N_2926,N_2360,N_2240);
and U2927 (N_2927,N_2095,N_2385);
or U2928 (N_2928,N_2167,N_2118);
or U2929 (N_2929,N_2191,N_2181);
nor U2930 (N_2930,N_2285,N_2186);
or U2931 (N_2931,N_2109,N_2219);
nand U2932 (N_2932,N_2225,N_2263);
nor U2933 (N_2933,N_2432,N_2348);
nand U2934 (N_2934,N_2419,N_2441);
and U2935 (N_2935,N_1894,N_2234);
or U2936 (N_2936,N_1991,N_2440);
and U2937 (N_2937,N_2441,N_2065);
nor U2938 (N_2938,N_1954,N_2461);
xor U2939 (N_2939,N_2347,N_2341);
nor U2940 (N_2940,N_2211,N_1961);
or U2941 (N_2941,N_2322,N_2294);
nor U2942 (N_2942,N_2149,N_1937);
nor U2943 (N_2943,N_1997,N_2337);
and U2944 (N_2944,N_2341,N_2365);
xnor U2945 (N_2945,N_2152,N_2167);
nand U2946 (N_2946,N_2464,N_2397);
nand U2947 (N_2947,N_1883,N_2488);
nor U2948 (N_2948,N_2349,N_2229);
nand U2949 (N_2949,N_1977,N_2083);
and U2950 (N_2950,N_2056,N_2310);
xnor U2951 (N_2951,N_2494,N_2101);
and U2952 (N_2952,N_2365,N_1883);
xnor U2953 (N_2953,N_2033,N_2118);
or U2954 (N_2954,N_1882,N_2152);
nor U2955 (N_2955,N_2360,N_2083);
xnor U2956 (N_2956,N_2487,N_2475);
nand U2957 (N_2957,N_2353,N_2416);
nand U2958 (N_2958,N_2229,N_2205);
and U2959 (N_2959,N_2195,N_2025);
xnor U2960 (N_2960,N_2047,N_1975);
nand U2961 (N_2961,N_2131,N_2044);
xnor U2962 (N_2962,N_1982,N_2122);
and U2963 (N_2963,N_2201,N_2486);
nand U2964 (N_2964,N_2084,N_2176);
and U2965 (N_2965,N_2403,N_2493);
xor U2966 (N_2966,N_2382,N_2291);
nor U2967 (N_2967,N_1920,N_2166);
xor U2968 (N_2968,N_2009,N_2243);
nor U2969 (N_2969,N_2171,N_2412);
nand U2970 (N_2970,N_2012,N_2167);
and U2971 (N_2971,N_2007,N_2408);
or U2972 (N_2972,N_2402,N_2351);
nand U2973 (N_2973,N_2125,N_2089);
and U2974 (N_2974,N_2327,N_2220);
xnor U2975 (N_2975,N_2122,N_2160);
xnor U2976 (N_2976,N_1948,N_2456);
xnor U2977 (N_2977,N_1974,N_2040);
xor U2978 (N_2978,N_2269,N_2434);
nand U2979 (N_2979,N_2302,N_2009);
or U2980 (N_2980,N_2257,N_2093);
nand U2981 (N_2981,N_2320,N_2305);
nor U2982 (N_2982,N_2386,N_2256);
or U2983 (N_2983,N_1895,N_2487);
or U2984 (N_2984,N_2316,N_2361);
nand U2985 (N_2985,N_1927,N_2400);
xnor U2986 (N_2986,N_1962,N_2487);
nand U2987 (N_2987,N_2328,N_1976);
nor U2988 (N_2988,N_2020,N_2333);
nand U2989 (N_2989,N_2152,N_2411);
or U2990 (N_2990,N_2127,N_2469);
or U2991 (N_2991,N_1987,N_1886);
nor U2992 (N_2992,N_2069,N_2331);
xor U2993 (N_2993,N_2271,N_2399);
xnor U2994 (N_2994,N_2461,N_2034);
and U2995 (N_2995,N_2408,N_2277);
xor U2996 (N_2996,N_2020,N_2367);
xor U2997 (N_2997,N_2311,N_1937);
xnor U2998 (N_2998,N_2373,N_2379);
nor U2999 (N_2999,N_2311,N_2181);
and U3000 (N_3000,N_2032,N_2102);
nand U3001 (N_3001,N_2282,N_1928);
or U3002 (N_3002,N_1907,N_2322);
and U3003 (N_3003,N_2067,N_2319);
or U3004 (N_3004,N_1915,N_2127);
and U3005 (N_3005,N_2081,N_2304);
or U3006 (N_3006,N_2025,N_2140);
or U3007 (N_3007,N_1935,N_2130);
and U3008 (N_3008,N_2113,N_2105);
xnor U3009 (N_3009,N_2059,N_2100);
and U3010 (N_3010,N_2211,N_2105);
and U3011 (N_3011,N_2320,N_2182);
nor U3012 (N_3012,N_2060,N_1924);
and U3013 (N_3013,N_2397,N_2047);
nand U3014 (N_3014,N_2338,N_2374);
or U3015 (N_3015,N_2146,N_2406);
nand U3016 (N_3016,N_2310,N_2309);
xnor U3017 (N_3017,N_1961,N_2464);
nand U3018 (N_3018,N_2006,N_2420);
xnor U3019 (N_3019,N_2042,N_1900);
or U3020 (N_3020,N_2426,N_1949);
or U3021 (N_3021,N_1879,N_2091);
nand U3022 (N_3022,N_2237,N_2387);
nand U3023 (N_3023,N_2182,N_2374);
and U3024 (N_3024,N_1950,N_2165);
or U3025 (N_3025,N_1940,N_2290);
nor U3026 (N_3026,N_2009,N_2246);
or U3027 (N_3027,N_1893,N_1919);
and U3028 (N_3028,N_2408,N_2335);
and U3029 (N_3029,N_2119,N_2289);
nand U3030 (N_3030,N_2247,N_2083);
and U3031 (N_3031,N_1915,N_2365);
nor U3032 (N_3032,N_2411,N_2242);
or U3033 (N_3033,N_2495,N_2034);
xnor U3034 (N_3034,N_2112,N_2223);
nand U3035 (N_3035,N_2357,N_2179);
nand U3036 (N_3036,N_2366,N_2104);
and U3037 (N_3037,N_2497,N_2457);
nand U3038 (N_3038,N_1988,N_2415);
or U3039 (N_3039,N_2310,N_1926);
and U3040 (N_3040,N_2325,N_2477);
or U3041 (N_3041,N_1932,N_2307);
nand U3042 (N_3042,N_2381,N_1995);
nor U3043 (N_3043,N_1902,N_2345);
nand U3044 (N_3044,N_2258,N_2117);
or U3045 (N_3045,N_2158,N_2207);
xor U3046 (N_3046,N_2010,N_1975);
or U3047 (N_3047,N_2048,N_2242);
xor U3048 (N_3048,N_2023,N_2337);
or U3049 (N_3049,N_2220,N_2045);
nor U3050 (N_3050,N_2413,N_2380);
and U3051 (N_3051,N_2383,N_2214);
or U3052 (N_3052,N_2249,N_2086);
nand U3053 (N_3053,N_2282,N_1921);
and U3054 (N_3054,N_2477,N_2017);
xnor U3055 (N_3055,N_2302,N_2007);
xor U3056 (N_3056,N_2083,N_2152);
nand U3057 (N_3057,N_1987,N_2356);
and U3058 (N_3058,N_2481,N_2199);
and U3059 (N_3059,N_2356,N_2115);
and U3060 (N_3060,N_1957,N_2384);
and U3061 (N_3061,N_2062,N_1953);
nand U3062 (N_3062,N_2071,N_1909);
nand U3063 (N_3063,N_2109,N_2343);
xor U3064 (N_3064,N_1909,N_2340);
xnor U3065 (N_3065,N_2011,N_1878);
xnor U3066 (N_3066,N_2054,N_2487);
and U3067 (N_3067,N_2145,N_2106);
nand U3068 (N_3068,N_2482,N_1922);
nand U3069 (N_3069,N_1966,N_2253);
or U3070 (N_3070,N_1953,N_2334);
and U3071 (N_3071,N_1920,N_2440);
or U3072 (N_3072,N_2301,N_1913);
nand U3073 (N_3073,N_1879,N_1966);
nand U3074 (N_3074,N_2499,N_1912);
and U3075 (N_3075,N_2014,N_2496);
nor U3076 (N_3076,N_2407,N_2116);
or U3077 (N_3077,N_2290,N_2196);
nand U3078 (N_3078,N_2425,N_2315);
xor U3079 (N_3079,N_1905,N_2273);
nand U3080 (N_3080,N_2157,N_2378);
or U3081 (N_3081,N_2315,N_2077);
xnor U3082 (N_3082,N_1892,N_2315);
nor U3083 (N_3083,N_2264,N_2140);
or U3084 (N_3084,N_2484,N_2140);
nand U3085 (N_3085,N_2115,N_2048);
xor U3086 (N_3086,N_1971,N_2222);
and U3087 (N_3087,N_2318,N_1990);
and U3088 (N_3088,N_2384,N_2034);
or U3089 (N_3089,N_1879,N_1951);
nor U3090 (N_3090,N_2092,N_2224);
nand U3091 (N_3091,N_1987,N_1999);
or U3092 (N_3092,N_1898,N_2000);
nor U3093 (N_3093,N_2229,N_2079);
xor U3094 (N_3094,N_2326,N_2178);
nand U3095 (N_3095,N_2171,N_2298);
xnor U3096 (N_3096,N_2463,N_2424);
and U3097 (N_3097,N_2293,N_1996);
xor U3098 (N_3098,N_2439,N_2339);
and U3099 (N_3099,N_2168,N_2050);
or U3100 (N_3100,N_2204,N_1984);
and U3101 (N_3101,N_2425,N_2456);
nand U3102 (N_3102,N_2452,N_2483);
xor U3103 (N_3103,N_1876,N_2197);
or U3104 (N_3104,N_2499,N_2161);
or U3105 (N_3105,N_2129,N_1941);
xor U3106 (N_3106,N_2439,N_2256);
nand U3107 (N_3107,N_2040,N_1949);
nor U3108 (N_3108,N_2151,N_2322);
or U3109 (N_3109,N_2262,N_2164);
nand U3110 (N_3110,N_2103,N_2015);
and U3111 (N_3111,N_2112,N_2161);
or U3112 (N_3112,N_1927,N_2076);
nor U3113 (N_3113,N_2065,N_2376);
xnor U3114 (N_3114,N_2334,N_2006);
nand U3115 (N_3115,N_2181,N_2076);
nand U3116 (N_3116,N_2166,N_2406);
xor U3117 (N_3117,N_2012,N_1942);
nor U3118 (N_3118,N_2053,N_1965);
nor U3119 (N_3119,N_1989,N_2339);
xor U3120 (N_3120,N_2288,N_2405);
nand U3121 (N_3121,N_2485,N_2017);
and U3122 (N_3122,N_2104,N_2054);
nand U3123 (N_3123,N_2374,N_2198);
xor U3124 (N_3124,N_2050,N_2326);
and U3125 (N_3125,N_2799,N_2670);
nor U3126 (N_3126,N_2815,N_2854);
or U3127 (N_3127,N_2642,N_3064);
or U3128 (N_3128,N_2794,N_2676);
nand U3129 (N_3129,N_2833,N_2659);
nor U3130 (N_3130,N_2719,N_2737);
or U3131 (N_3131,N_2714,N_3085);
or U3132 (N_3132,N_2554,N_2955);
nand U3133 (N_3133,N_2764,N_2996);
xnor U3134 (N_3134,N_2739,N_2848);
or U3135 (N_3135,N_2920,N_2548);
nor U3136 (N_3136,N_3047,N_2699);
nor U3137 (N_3137,N_3031,N_2513);
nor U3138 (N_3138,N_2929,N_2767);
nor U3139 (N_3139,N_2805,N_2504);
or U3140 (N_3140,N_2564,N_2705);
or U3141 (N_3141,N_2656,N_3083);
xnor U3142 (N_3142,N_3104,N_2568);
nand U3143 (N_3143,N_2536,N_2661);
or U3144 (N_3144,N_2570,N_2840);
xnor U3145 (N_3145,N_3110,N_3001);
and U3146 (N_3146,N_2509,N_3079);
or U3147 (N_3147,N_2587,N_2851);
and U3148 (N_3148,N_3045,N_2911);
xnor U3149 (N_3149,N_2766,N_2763);
or U3150 (N_3150,N_2663,N_3086);
or U3151 (N_3151,N_2567,N_2586);
xor U3152 (N_3152,N_2639,N_3005);
xnor U3153 (N_3153,N_2557,N_2876);
nand U3154 (N_3154,N_2745,N_3032);
nor U3155 (N_3155,N_2643,N_2753);
xnor U3156 (N_3156,N_2776,N_3072);
nand U3157 (N_3157,N_2600,N_2706);
xor U3158 (N_3158,N_3101,N_2665);
nand U3159 (N_3159,N_2521,N_3108);
nand U3160 (N_3160,N_2510,N_2878);
or U3161 (N_3161,N_2960,N_3010);
and U3162 (N_3162,N_2980,N_2680);
and U3163 (N_3163,N_3002,N_2507);
xor U3164 (N_3164,N_2725,N_2779);
xor U3165 (N_3165,N_2566,N_2875);
nor U3166 (N_3166,N_2762,N_2723);
nand U3167 (N_3167,N_2900,N_2826);
xor U3168 (N_3168,N_3092,N_2597);
or U3169 (N_3169,N_2824,N_2910);
and U3170 (N_3170,N_2844,N_3078);
nor U3171 (N_3171,N_3118,N_2654);
nand U3172 (N_3172,N_2651,N_3048);
and U3173 (N_3173,N_3068,N_2538);
or U3174 (N_3174,N_2653,N_2615);
or U3175 (N_3175,N_2619,N_2914);
nor U3176 (N_3176,N_2608,N_2730);
nor U3177 (N_3177,N_2899,N_2593);
nand U3178 (N_3178,N_2853,N_2944);
and U3179 (N_3179,N_2527,N_3076);
nand U3180 (N_3180,N_2704,N_2674);
or U3181 (N_3181,N_2817,N_2750);
and U3182 (N_3182,N_3013,N_2894);
and U3183 (N_3183,N_3063,N_2873);
or U3184 (N_3184,N_2720,N_2971);
or U3185 (N_3185,N_2585,N_2519);
nor U3186 (N_3186,N_2939,N_2821);
nor U3187 (N_3187,N_2591,N_2685);
and U3188 (N_3188,N_2865,N_3023);
and U3189 (N_3189,N_2917,N_2697);
and U3190 (N_3190,N_2775,N_2648);
and U3191 (N_3191,N_2916,N_2930);
and U3192 (N_3192,N_2967,N_2992);
nor U3193 (N_3193,N_2603,N_2921);
or U3194 (N_3194,N_2769,N_2842);
nand U3195 (N_3195,N_2777,N_2636);
nand U3196 (N_3196,N_2502,N_2781);
or U3197 (N_3197,N_2890,N_2517);
and U3198 (N_3198,N_2846,N_2617);
xor U3199 (N_3199,N_2933,N_2578);
nor U3200 (N_3200,N_2695,N_2728);
or U3201 (N_3201,N_2556,N_2631);
and U3202 (N_3202,N_3030,N_2647);
or U3203 (N_3203,N_2547,N_2668);
or U3204 (N_3204,N_2713,N_2868);
nand U3205 (N_3205,N_2925,N_2645);
nor U3206 (N_3206,N_2732,N_3006);
xor U3207 (N_3207,N_3046,N_3016);
and U3208 (N_3208,N_2823,N_2908);
or U3209 (N_3209,N_2870,N_2516);
nor U3210 (N_3210,N_2828,N_2523);
and U3211 (N_3211,N_2688,N_2816);
nand U3212 (N_3212,N_2679,N_2748);
nor U3213 (N_3213,N_3107,N_3082);
nand U3214 (N_3214,N_2666,N_2683);
nand U3215 (N_3215,N_2582,N_3040);
and U3216 (N_3216,N_2512,N_2864);
or U3217 (N_3217,N_2847,N_2742);
nor U3218 (N_3218,N_3009,N_2596);
nor U3219 (N_3219,N_2788,N_2956);
and U3220 (N_3220,N_3119,N_2958);
and U3221 (N_3221,N_2595,N_2809);
and U3222 (N_3222,N_2797,N_2711);
nor U3223 (N_3223,N_2698,N_2687);
or U3224 (N_3224,N_3115,N_3065);
xnor U3225 (N_3225,N_2918,N_3094);
or U3226 (N_3226,N_2827,N_2551);
xnor U3227 (N_3227,N_2752,N_2852);
nor U3228 (N_3228,N_3051,N_2975);
nand U3229 (N_3229,N_3035,N_2795);
and U3230 (N_3230,N_3088,N_3116);
xnor U3231 (N_3231,N_2624,N_2961);
or U3232 (N_3232,N_2858,N_2838);
nor U3233 (N_3233,N_2985,N_2681);
nor U3234 (N_3234,N_2877,N_3060);
xor U3235 (N_3235,N_2501,N_2924);
xnor U3236 (N_3236,N_2998,N_2667);
nor U3237 (N_3237,N_3084,N_2834);
nand U3238 (N_3238,N_2758,N_2690);
nand U3239 (N_3239,N_2829,N_2987);
xor U3240 (N_3240,N_3049,N_2581);
nor U3241 (N_3241,N_2907,N_2796);
nand U3242 (N_3242,N_3120,N_2935);
and U3243 (N_3243,N_3012,N_2822);
nand U3244 (N_3244,N_2791,N_3112);
xor U3245 (N_3245,N_2717,N_3096);
nor U3246 (N_3246,N_2880,N_2773);
and U3247 (N_3247,N_2601,N_2802);
and U3248 (N_3248,N_2729,N_2740);
or U3249 (N_3249,N_3003,N_2830);
nand U3250 (N_3250,N_2923,N_2895);
xnor U3251 (N_3251,N_2574,N_3089);
and U3252 (N_3252,N_2818,N_2633);
or U3253 (N_3253,N_2966,N_2912);
and U3254 (N_3254,N_2937,N_2979);
and U3255 (N_3255,N_2563,N_2500);
and U3256 (N_3256,N_3097,N_2530);
or U3257 (N_3257,N_2938,N_2810);
or U3258 (N_3258,N_2941,N_2771);
and U3259 (N_3259,N_2575,N_2902);
xnor U3260 (N_3260,N_2843,N_2526);
or U3261 (N_3261,N_2889,N_2760);
nor U3262 (N_3262,N_2522,N_2727);
xnor U3263 (N_3263,N_2897,N_2977);
nand U3264 (N_3264,N_2855,N_2784);
nor U3265 (N_3265,N_2707,N_2820);
xor U3266 (N_3266,N_2637,N_2814);
nor U3267 (N_3267,N_2936,N_2808);
nor U3268 (N_3268,N_3123,N_2803);
nand U3269 (N_3269,N_2630,N_3095);
nand U3270 (N_3270,N_2589,N_2678);
nand U3271 (N_3271,N_2850,N_2959);
or U3272 (N_3272,N_2550,N_2628);
nor U3273 (N_3273,N_3022,N_2761);
nand U3274 (N_3274,N_2528,N_2609);
xor U3275 (N_3275,N_2515,N_2555);
nand U3276 (N_3276,N_2614,N_3020);
xnor U3277 (N_3277,N_3058,N_2755);
nand U3278 (N_3278,N_2590,N_2968);
xnor U3279 (N_3279,N_2765,N_3093);
and U3280 (N_3280,N_2849,N_2896);
or U3281 (N_3281,N_2943,N_2525);
nor U3282 (N_3282,N_2859,N_2743);
nand U3283 (N_3283,N_2533,N_2726);
and U3284 (N_3284,N_2613,N_3024);
xor U3285 (N_3285,N_2986,N_2673);
xor U3286 (N_3286,N_2542,N_2905);
nand U3287 (N_3287,N_2552,N_3066);
or U3288 (N_3288,N_3117,N_2749);
xnor U3289 (N_3289,N_2592,N_3056);
xnor U3290 (N_3290,N_2942,N_2731);
nand U3291 (N_3291,N_2928,N_2598);
or U3292 (N_3292,N_2560,N_2543);
or U3293 (N_3293,N_2825,N_3122);
or U3294 (N_3294,N_2511,N_2759);
nor U3295 (N_3295,N_2997,N_3021);
and U3296 (N_3296,N_2839,N_2789);
nor U3297 (N_3297,N_2952,N_2620);
nor U3298 (N_3298,N_2804,N_3121);
nand U3299 (N_3299,N_2583,N_2774);
nand U3300 (N_3300,N_3050,N_3103);
and U3301 (N_3301,N_2904,N_2709);
nand U3302 (N_3302,N_2863,N_3113);
nand U3303 (N_3303,N_2915,N_2622);
and U3304 (N_3304,N_3008,N_2607);
nand U3305 (N_3305,N_2879,N_2945);
nor U3306 (N_3306,N_3037,N_3102);
and U3307 (N_3307,N_2638,N_2577);
xnor U3308 (N_3308,N_2991,N_2783);
or U3309 (N_3309,N_3015,N_2972);
or U3310 (N_3310,N_2708,N_2541);
xnor U3311 (N_3311,N_3027,N_2953);
xor U3312 (N_3312,N_3038,N_2520);
or U3313 (N_3313,N_2976,N_2934);
or U3314 (N_3314,N_2835,N_2800);
nand U3315 (N_3315,N_2983,N_2508);
nor U3316 (N_3316,N_2872,N_2993);
nand U3317 (N_3317,N_2768,N_2995);
nand U3318 (N_3318,N_3124,N_2963);
xor U3319 (N_3319,N_2922,N_3109);
xor U3320 (N_3320,N_3033,N_3061);
xor U3321 (N_3321,N_2701,N_3025);
xor U3322 (N_3322,N_2957,N_2950);
nand U3323 (N_3323,N_2886,N_3081);
nand U3324 (N_3324,N_2506,N_2696);
and U3325 (N_3325,N_2571,N_2580);
or U3326 (N_3326,N_2724,N_2505);
xnor U3327 (N_3327,N_2691,N_2909);
nand U3328 (N_3328,N_3074,N_3090);
xnor U3329 (N_3329,N_2990,N_2883);
xnor U3330 (N_3330,N_2532,N_2962);
nand U3331 (N_3331,N_2514,N_2632);
nor U3332 (N_3332,N_2994,N_2801);
and U3333 (N_3333,N_2634,N_2970);
or U3334 (N_3334,N_2931,N_2832);
xor U3335 (N_3335,N_2888,N_2901);
or U3336 (N_3336,N_2792,N_2569);
and U3337 (N_3337,N_2841,N_2721);
xnor U3338 (N_3338,N_2741,N_3106);
nor U3339 (N_3339,N_3087,N_2862);
or U3340 (N_3340,N_2669,N_2984);
nand U3341 (N_3341,N_2973,N_2671);
xnor U3342 (N_3342,N_2616,N_2565);
or U3343 (N_3343,N_3070,N_2735);
and U3344 (N_3344,N_2602,N_2887);
and U3345 (N_3345,N_3034,N_2964);
nand U3346 (N_3346,N_2756,N_2926);
nor U3347 (N_3347,N_3100,N_2641);
and U3348 (N_3348,N_2734,N_3091);
xor U3349 (N_3349,N_3080,N_2747);
nand U3350 (N_3350,N_2710,N_2682);
nor U3351 (N_3351,N_2594,N_2540);
nand U3352 (N_3352,N_2785,N_2549);
nor U3353 (N_3353,N_3053,N_2629);
and U3354 (N_3354,N_2780,N_2529);
xnor U3355 (N_3355,N_2626,N_2693);
nor U3356 (N_3356,N_3039,N_2866);
or U3357 (N_3357,N_3062,N_3105);
xor U3358 (N_3358,N_2715,N_2584);
nor U3359 (N_3359,N_2874,N_2546);
xnor U3360 (N_3360,N_2787,N_2657);
and U3361 (N_3361,N_2524,N_2702);
xor U3362 (N_3362,N_2625,N_2978);
or U3363 (N_3363,N_2989,N_3007);
or U3364 (N_3364,N_2965,N_3043);
and U3365 (N_3365,N_2778,N_2845);
xnor U3366 (N_3366,N_2819,N_2757);
nor U3367 (N_3367,N_2738,N_2553);
xor U3368 (N_3368,N_2885,N_3067);
or U3369 (N_3369,N_2919,N_2660);
nor U3370 (N_3370,N_2712,N_2718);
nor U3371 (N_3371,N_2621,N_2932);
xor U3372 (N_3372,N_2605,N_3052);
xor U3373 (N_3373,N_2545,N_2982);
or U3374 (N_3374,N_2535,N_2686);
nand U3375 (N_3375,N_2947,N_2969);
xnor U3376 (N_3376,N_2646,N_2867);
xnor U3377 (N_3377,N_2627,N_2981);
and U3378 (N_3378,N_3019,N_3073);
or U3379 (N_3379,N_2798,N_3041);
nor U3380 (N_3380,N_2949,N_2531);
xor U3381 (N_3381,N_2974,N_2793);
xnor U3382 (N_3382,N_3069,N_2812);
or U3383 (N_3383,N_2611,N_2898);
nand U3384 (N_3384,N_2837,N_2503);
or U3385 (N_3385,N_2836,N_2612);
nand U3386 (N_3386,N_2813,N_2951);
xnor U3387 (N_3387,N_2988,N_2882);
xnor U3388 (N_3388,N_3042,N_2618);
nand U3389 (N_3389,N_2662,N_2623);
and U3390 (N_3390,N_2658,N_3011);
and U3391 (N_3391,N_3044,N_2999);
or U3392 (N_3392,N_2856,N_3036);
nand U3393 (N_3393,N_2650,N_2562);
nand U3394 (N_3394,N_2572,N_2893);
and U3395 (N_3395,N_2954,N_2689);
nand U3396 (N_3396,N_2640,N_2579);
or U3397 (N_3397,N_2744,N_2694);
nand U3398 (N_3398,N_2561,N_2881);
or U3399 (N_3399,N_2606,N_2716);
nor U3400 (N_3400,N_2675,N_2644);
xor U3401 (N_3401,N_3057,N_2940);
and U3402 (N_3402,N_2677,N_2736);
xor U3403 (N_3403,N_2576,N_2703);
nor U3404 (N_3404,N_2807,N_3000);
and U3405 (N_3405,N_3098,N_2537);
or U3406 (N_3406,N_3018,N_2733);
and U3407 (N_3407,N_2746,N_3059);
and U3408 (N_3408,N_2588,N_2751);
nand U3409 (N_3409,N_2892,N_2754);
nor U3410 (N_3410,N_2558,N_2573);
nor U3411 (N_3411,N_3054,N_2946);
and U3412 (N_3412,N_2672,N_2722);
xnor U3413 (N_3413,N_3017,N_2684);
xnor U3414 (N_3414,N_2649,N_2806);
nor U3415 (N_3415,N_2869,N_3026);
nor U3416 (N_3416,N_2770,N_2906);
or U3417 (N_3417,N_2655,N_3014);
and U3418 (N_3418,N_2635,N_2927);
nor U3419 (N_3419,N_3055,N_3004);
nand U3420 (N_3420,N_2884,N_2871);
nor U3421 (N_3421,N_2948,N_2652);
nand U3422 (N_3422,N_2559,N_3075);
nand U3423 (N_3423,N_2664,N_2700);
nand U3424 (N_3424,N_2544,N_2772);
xor U3425 (N_3425,N_2610,N_3111);
xor U3426 (N_3426,N_2534,N_2604);
and U3427 (N_3427,N_2913,N_3114);
nor U3428 (N_3428,N_2782,N_2891);
or U3429 (N_3429,N_3071,N_2831);
and U3430 (N_3430,N_2599,N_2790);
nor U3431 (N_3431,N_3077,N_2539);
nand U3432 (N_3432,N_2857,N_2861);
nand U3433 (N_3433,N_2692,N_3099);
nand U3434 (N_3434,N_3028,N_2903);
nor U3435 (N_3435,N_2786,N_2518);
nor U3436 (N_3436,N_3029,N_2811);
nor U3437 (N_3437,N_2860,N_2747);
nor U3438 (N_3438,N_2601,N_2841);
nor U3439 (N_3439,N_2533,N_2801);
and U3440 (N_3440,N_2852,N_2518);
and U3441 (N_3441,N_2976,N_2673);
nor U3442 (N_3442,N_2522,N_3068);
and U3443 (N_3443,N_3022,N_3049);
xnor U3444 (N_3444,N_2693,N_2712);
or U3445 (N_3445,N_2658,N_3052);
nor U3446 (N_3446,N_2738,N_2849);
or U3447 (N_3447,N_2953,N_3084);
and U3448 (N_3448,N_2949,N_2855);
or U3449 (N_3449,N_2798,N_3115);
nand U3450 (N_3450,N_2631,N_3082);
and U3451 (N_3451,N_2661,N_2738);
nand U3452 (N_3452,N_2500,N_2644);
nand U3453 (N_3453,N_2729,N_2916);
and U3454 (N_3454,N_2599,N_3051);
nor U3455 (N_3455,N_2727,N_2791);
nor U3456 (N_3456,N_2927,N_2898);
nand U3457 (N_3457,N_2974,N_3031);
nor U3458 (N_3458,N_2890,N_2779);
and U3459 (N_3459,N_2799,N_2633);
nand U3460 (N_3460,N_2535,N_2768);
or U3461 (N_3461,N_2833,N_3121);
xnor U3462 (N_3462,N_2987,N_2977);
nor U3463 (N_3463,N_2981,N_2667);
and U3464 (N_3464,N_3062,N_2997);
xor U3465 (N_3465,N_2624,N_2967);
and U3466 (N_3466,N_2979,N_2719);
nor U3467 (N_3467,N_2856,N_3059);
and U3468 (N_3468,N_3041,N_2773);
nor U3469 (N_3469,N_2839,N_2826);
and U3470 (N_3470,N_2510,N_2799);
and U3471 (N_3471,N_2978,N_2968);
nor U3472 (N_3472,N_3095,N_2945);
nand U3473 (N_3473,N_2589,N_2731);
nand U3474 (N_3474,N_3122,N_2604);
nor U3475 (N_3475,N_3041,N_3047);
and U3476 (N_3476,N_2730,N_2548);
or U3477 (N_3477,N_2564,N_2855);
or U3478 (N_3478,N_3124,N_2755);
nor U3479 (N_3479,N_2912,N_2843);
and U3480 (N_3480,N_2963,N_2912);
nand U3481 (N_3481,N_2579,N_2801);
nor U3482 (N_3482,N_2929,N_2551);
and U3483 (N_3483,N_2672,N_3109);
and U3484 (N_3484,N_2626,N_2848);
nor U3485 (N_3485,N_2887,N_2651);
and U3486 (N_3486,N_2636,N_3114);
xor U3487 (N_3487,N_2880,N_2831);
nor U3488 (N_3488,N_2688,N_2875);
and U3489 (N_3489,N_2779,N_2506);
and U3490 (N_3490,N_2964,N_2565);
xor U3491 (N_3491,N_2966,N_2909);
or U3492 (N_3492,N_3123,N_2777);
nor U3493 (N_3493,N_3092,N_2867);
and U3494 (N_3494,N_2518,N_3066);
and U3495 (N_3495,N_2667,N_2826);
nand U3496 (N_3496,N_2807,N_2944);
nor U3497 (N_3497,N_2933,N_2616);
or U3498 (N_3498,N_2670,N_3101);
and U3499 (N_3499,N_2775,N_2691);
and U3500 (N_3500,N_2976,N_2971);
xor U3501 (N_3501,N_2641,N_2534);
nor U3502 (N_3502,N_3045,N_2963);
nand U3503 (N_3503,N_2821,N_3004);
and U3504 (N_3504,N_2771,N_2604);
or U3505 (N_3505,N_2762,N_2995);
xor U3506 (N_3506,N_3082,N_2652);
and U3507 (N_3507,N_3014,N_2647);
nor U3508 (N_3508,N_2604,N_2580);
and U3509 (N_3509,N_2910,N_2661);
nand U3510 (N_3510,N_2558,N_2552);
nand U3511 (N_3511,N_2584,N_2735);
nor U3512 (N_3512,N_2877,N_2745);
nor U3513 (N_3513,N_2870,N_2907);
nand U3514 (N_3514,N_2799,N_2926);
xor U3515 (N_3515,N_3105,N_2922);
xor U3516 (N_3516,N_2682,N_2598);
xor U3517 (N_3517,N_2607,N_3118);
xnor U3518 (N_3518,N_2900,N_2583);
nand U3519 (N_3519,N_2605,N_2944);
nand U3520 (N_3520,N_2501,N_2519);
nand U3521 (N_3521,N_2601,N_2870);
nand U3522 (N_3522,N_2780,N_3000);
and U3523 (N_3523,N_2715,N_2774);
or U3524 (N_3524,N_2644,N_2937);
and U3525 (N_3525,N_2548,N_3028);
or U3526 (N_3526,N_2533,N_2654);
xor U3527 (N_3527,N_2879,N_3121);
xor U3528 (N_3528,N_2761,N_2795);
and U3529 (N_3529,N_2717,N_2630);
and U3530 (N_3530,N_2683,N_2847);
and U3531 (N_3531,N_2976,N_2580);
or U3532 (N_3532,N_3079,N_2578);
nor U3533 (N_3533,N_3057,N_2925);
nor U3534 (N_3534,N_3024,N_2995);
nand U3535 (N_3535,N_2517,N_2577);
nor U3536 (N_3536,N_2693,N_2612);
and U3537 (N_3537,N_2795,N_2745);
and U3538 (N_3538,N_2971,N_2730);
or U3539 (N_3539,N_2971,N_2644);
nor U3540 (N_3540,N_3081,N_2792);
nand U3541 (N_3541,N_2834,N_3057);
nand U3542 (N_3542,N_2718,N_2668);
xor U3543 (N_3543,N_3005,N_3027);
nand U3544 (N_3544,N_2551,N_2789);
and U3545 (N_3545,N_2744,N_2584);
and U3546 (N_3546,N_2742,N_2935);
xnor U3547 (N_3547,N_2770,N_3005);
or U3548 (N_3548,N_2638,N_2508);
and U3549 (N_3549,N_2955,N_2753);
nor U3550 (N_3550,N_2522,N_2516);
and U3551 (N_3551,N_2983,N_2560);
and U3552 (N_3552,N_3026,N_2533);
xnor U3553 (N_3553,N_3106,N_2854);
nor U3554 (N_3554,N_2656,N_2642);
nor U3555 (N_3555,N_2901,N_2722);
and U3556 (N_3556,N_3014,N_2874);
nand U3557 (N_3557,N_2973,N_2605);
or U3558 (N_3558,N_2591,N_2629);
and U3559 (N_3559,N_2874,N_2715);
nand U3560 (N_3560,N_2689,N_2536);
nand U3561 (N_3561,N_2610,N_2536);
nand U3562 (N_3562,N_2838,N_3106);
or U3563 (N_3563,N_3084,N_2940);
and U3564 (N_3564,N_2770,N_2569);
nor U3565 (N_3565,N_2720,N_3075);
nor U3566 (N_3566,N_2507,N_2622);
xor U3567 (N_3567,N_3020,N_2661);
nand U3568 (N_3568,N_2715,N_3071);
xor U3569 (N_3569,N_3043,N_2775);
and U3570 (N_3570,N_2823,N_2730);
nor U3571 (N_3571,N_2632,N_2832);
and U3572 (N_3572,N_2630,N_3082);
and U3573 (N_3573,N_3009,N_2624);
or U3574 (N_3574,N_2538,N_2720);
xor U3575 (N_3575,N_2791,N_2718);
xor U3576 (N_3576,N_2858,N_3001);
xnor U3577 (N_3577,N_2856,N_2607);
xor U3578 (N_3578,N_2986,N_2871);
nor U3579 (N_3579,N_2775,N_2534);
nor U3580 (N_3580,N_3027,N_3068);
xnor U3581 (N_3581,N_2536,N_2618);
nor U3582 (N_3582,N_2752,N_3029);
or U3583 (N_3583,N_2549,N_2889);
xor U3584 (N_3584,N_2805,N_3045);
nand U3585 (N_3585,N_2910,N_2923);
nor U3586 (N_3586,N_2523,N_3002);
or U3587 (N_3587,N_2775,N_2810);
or U3588 (N_3588,N_2621,N_2735);
and U3589 (N_3589,N_2970,N_3011);
or U3590 (N_3590,N_2629,N_2988);
nand U3591 (N_3591,N_2721,N_2701);
xor U3592 (N_3592,N_2646,N_2555);
xnor U3593 (N_3593,N_3111,N_2526);
xor U3594 (N_3594,N_3023,N_2578);
nor U3595 (N_3595,N_2695,N_2992);
or U3596 (N_3596,N_2588,N_2846);
nand U3597 (N_3597,N_2884,N_2629);
and U3598 (N_3598,N_2533,N_3090);
or U3599 (N_3599,N_2884,N_3015);
nor U3600 (N_3600,N_2999,N_2539);
nand U3601 (N_3601,N_2639,N_2893);
nor U3602 (N_3602,N_2856,N_2874);
nand U3603 (N_3603,N_2600,N_2888);
xnor U3604 (N_3604,N_2648,N_2754);
xor U3605 (N_3605,N_3112,N_2842);
or U3606 (N_3606,N_2529,N_3063);
and U3607 (N_3607,N_2766,N_3101);
nor U3608 (N_3608,N_2718,N_2914);
and U3609 (N_3609,N_2733,N_2886);
nor U3610 (N_3610,N_3071,N_2586);
nor U3611 (N_3611,N_2654,N_2638);
and U3612 (N_3612,N_2648,N_2985);
nand U3613 (N_3613,N_2627,N_2956);
or U3614 (N_3614,N_2979,N_2701);
nor U3615 (N_3615,N_3107,N_3050);
nand U3616 (N_3616,N_2548,N_2793);
xor U3617 (N_3617,N_2645,N_2874);
or U3618 (N_3618,N_2893,N_3001);
nor U3619 (N_3619,N_2698,N_2776);
and U3620 (N_3620,N_2753,N_2729);
nor U3621 (N_3621,N_2612,N_2910);
xnor U3622 (N_3622,N_2804,N_2665);
nand U3623 (N_3623,N_3066,N_2768);
or U3624 (N_3624,N_2804,N_2589);
xnor U3625 (N_3625,N_2508,N_2665);
nand U3626 (N_3626,N_2585,N_2742);
and U3627 (N_3627,N_3014,N_2710);
xor U3628 (N_3628,N_3084,N_2605);
nand U3629 (N_3629,N_2674,N_2709);
and U3630 (N_3630,N_2546,N_2838);
or U3631 (N_3631,N_2605,N_2684);
or U3632 (N_3632,N_3045,N_2718);
nor U3633 (N_3633,N_2814,N_2590);
or U3634 (N_3634,N_3030,N_2610);
nor U3635 (N_3635,N_2622,N_2619);
nor U3636 (N_3636,N_2660,N_3112);
and U3637 (N_3637,N_2771,N_3089);
or U3638 (N_3638,N_2856,N_3094);
nor U3639 (N_3639,N_2623,N_2608);
or U3640 (N_3640,N_3001,N_2825);
and U3641 (N_3641,N_2660,N_2646);
nand U3642 (N_3642,N_2947,N_2888);
or U3643 (N_3643,N_2895,N_3053);
xor U3644 (N_3644,N_2514,N_2533);
and U3645 (N_3645,N_3022,N_2843);
nor U3646 (N_3646,N_3071,N_2900);
and U3647 (N_3647,N_2598,N_2963);
nand U3648 (N_3648,N_2881,N_2779);
and U3649 (N_3649,N_2544,N_2782);
nor U3650 (N_3650,N_3117,N_2855);
nor U3651 (N_3651,N_3006,N_2862);
and U3652 (N_3652,N_2949,N_2807);
and U3653 (N_3653,N_2771,N_2874);
nand U3654 (N_3654,N_2959,N_2875);
or U3655 (N_3655,N_3092,N_2551);
or U3656 (N_3656,N_2995,N_2833);
and U3657 (N_3657,N_2717,N_2658);
nor U3658 (N_3658,N_2670,N_2903);
or U3659 (N_3659,N_2761,N_2644);
nor U3660 (N_3660,N_2783,N_3011);
nand U3661 (N_3661,N_2537,N_3048);
xnor U3662 (N_3662,N_3047,N_2921);
nand U3663 (N_3663,N_3098,N_3076);
or U3664 (N_3664,N_2672,N_2961);
nor U3665 (N_3665,N_3016,N_3092);
nor U3666 (N_3666,N_2698,N_2683);
and U3667 (N_3667,N_2957,N_2556);
nand U3668 (N_3668,N_2588,N_2643);
and U3669 (N_3669,N_2572,N_2616);
nand U3670 (N_3670,N_2839,N_2933);
and U3671 (N_3671,N_2502,N_2907);
or U3672 (N_3672,N_2643,N_2536);
xor U3673 (N_3673,N_2993,N_2603);
xnor U3674 (N_3674,N_3032,N_2533);
nor U3675 (N_3675,N_2984,N_2755);
nor U3676 (N_3676,N_2698,N_3068);
nor U3677 (N_3677,N_3078,N_2941);
nand U3678 (N_3678,N_3097,N_2767);
or U3679 (N_3679,N_2843,N_2835);
nor U3680 (N_3680,N_2615,N_2819);
and U3681 (N_3681,N_2601,N_3009);
xor U3682 (N_3682,N_2735,N_2818);
xnor U3683 (N_3683,N_2528,N_2932);
xnor U3684 (N_3684,N_3096,N_2678);
xnor U3685 (N_3685,N_3094,N_2553);
nor U3686 (N_3686,N_2950,N_2746);
nand U3687 (N_3687,N_2937,N_2860);
and U3688 (N_3688,N_3039,N_2876);
or U3689 (N_3689,N_2708,N_3094);
nand U3690 (N_3690,N_2565,N_2555);
and U3691 (N_3691,N_2902,N_2555);
nor U3692 (N_3692,N_2767,N_2692);
and U3693 (N_3693,N_2602,N_2629);
and U3694 (N_3694,N_2604,N_2779);
nor U3695 (N_3695,N_2920,N_2838);
nor U3696 (N_3696,N_3024,N_2631);
xnor U3697 (N_3697,N_2657,N_2872);
or U3698 (N_3698,N_2885,N_2665);
and U3699 (N_3699,N_2915,N_2584);
or U3700 (N_3700,N_3045,N_2550);
nand U3701 (N_3701,N_2603,N_3066);
xnor U3702 (N_3702,N_3027,N_2896);
or U3703 (N_3703,N_2719,N_2598);
nand U3704 (N_3704,N_2895,N_2947);
or U3705 (N_3705,N_3045,N_3117);
xor U3706 (N_3706,N_2770,N_2774);
xnor U3707 (N_3707,N_2517,N_2881);
xor U3708 (N_3708,N_2715,N_2753);
or U3709 (N_3709,N_2985,N_2954);
nor U3710 (N_3710,N_2723,N_2954);
or U3711 (N_3711,N_2964,N_2535);
nor U3712 (N_3712,N_2624,N_2852);
and U3713 (N_3713,N_2959,N_3003);
or U3714 (N_3714,N_2926,N_2961);
nor U3715 (N_3715,N_2736,N_3064);
xor U3716 (N_3716,N_3051,N_2537);
or U3717 (N_3717,N_2873,N_2867);
nand U3718 (N_3718,N_2875,N_2656);
or U3719 (N_3719,N_3038,N_2819);
or U3720 (N_3720,N_2576,N_3102);
xnor U3721 (N_3721,N_2509,N_2897);
and U3722 (N_3722,N_2521,N_2820);
nand U3723 (N_3723,N_2994,N_2828);
nor U3724 (N_3724,N_2567,N_3098);
xor U3725 (N_3725,N_2563,N_2632);
or U3726 (N_3726,N_2767,N_3064);
or U3727 (N_3727,N_2619,N_3037);
nand U3728 (N_3728,N_2984,N_2909);
xor U3729 (N_3729,N_3108,N_3014);
nor U3730 (N_3730,N_2651,N_2868);
and U3731 (N_3731,N_2756,N_2980);
and U3732 (N_3732,N_2500,N_2813);
xnor U3733 (N_3733,N_3068,N_2551);
nor U3734 (N_3734,N_2927,N_2659);
or U3735 (N_3735,N_3067,N_2761);
or U3736 (N_3736,N_2654,N_2628);
or U3737 (N_3737,N_2957,N_3010);
xor U3738 (N_3738,N_2673,N_2547);
nor U3739 (N_3739,N_2693,N_2611);
nand U3740 (N_3740,N_3033,N_3048);
or U3741 (N_3741,N_2645,N_2669);
xor U3742 (N_3742,N_2633,N_3086);
nand U3743 (N_3743,N_2652,N_2613);
and U3744 (N_3744,N_3091,N_2579);
xnor U3745 (N_3745,N_3105,N_2676);
nand U3746 (N_3746,N_2800,N_3050);
xor U3747 (N_3747,N_2705,N_2778);
nor U3748 (N_3748,N_3074,N_2623);
nand U3749 (N_3749,N_2646,N_3076);
xnor U3750 (N_3750,N_3293,N_3134);
xor U3751 (N_3751,N_3494,N_3423);
or U3752 (N_3752,N_3712,N_3150);
or U3753 (N_3753,N_3718,N_3282);
nand U3754 (N_3754,N_3379,N_3402);
and U3755 (N_3755,N_3335,N_3462);
nor U3756 (N_3756,N_3298,N_3260);
nor U3757 (N_3757,N_3355,N_3395);
and U3758 (N_3758,N_3160,N_3146);
nor U3759 (N_3759,N_3653,N_3204);
nor U3760 (N_3760,N_3680,N_3378);
or U3761 (N_3761,N_3655,N_3634);
nor U3762 (N_3762,N_3201,N_3565);
xor U3763 (N_3763,N_3276,N_3745);
xnor U3764 (N_3764,N_3420,N_3301);
nand U3765 (N_3765,N_3314,N_3598);
nor U3766 (N_3766,N_3589,N_3631);
and U3767 (N_3767,N_3461,N_3400);
or U3768 (N_3768,N_3261,N_3579);
and U3769 (N_3769,N_3645,N_3135);
or U3770 (N_3770,N_3733,N_3270);
nor U3771 (N_3771,N_3453,N_3251);
and U3772 (N_3772,N_3452,N_3376);
nor U3773 (N_3773,N_3370,N_3695);
xor U3774 (N_3774,N_3515,N_3361);
nor U3775 (N_3775,N_3303,N_3235);
or U3776 (N_3776,N_3384,N_3677);
nor U3777 (N_3777,N_3585,N_3366);
nand U3778 (N_3778,N_3648,N_3299);
xnor U3779 (N_3779,N_3536,N_3243);
and U3780 (N_3780,N_3467,N_3180);
nand U3781 (N_3781,N_3621,N_3309);
nor U3782 (N_3782,N_3573,N_3560);
nand U3783 (N_3783,N_3422,N_3222);
and U3784 (N_3784,N_3432,N_3702);
and U3785 (N_3785,N_3709,N_3548);
nand U3786 (N_3786,N_3182,N_3721);
nor U3787 (N_3787,N_3140,N_3212);
xor U3788 (N_3788,N_3698,N_3673);
or U3789 (N_3789,N_3392,N_3224);
xor U3790 (N_3790,N_3491,N_3255);
or U3791 (N_3791,N_3343,N_3318);
nand U3792 (N_3792,N_3678,N_3509);
nand U3793 (N_3793,N_3143,N_3390);
or U3794 (N_3794,N_3728,N_3337);
and U3795 (N_3795,N_3660,N_3741);
and U3796 (N_3796,N_3531,N_3170);
xnor U3797 (N_3797,N_3271,N_3538);
nand U3798 (N_3798,N_3528,N_3177);
and U3799 (N_3799,N_3288,N_3389);
nand U3800 (N_3800,N_3502,N_3574);
nand U3801 (N_3801,N_3372,N_3597);
nor U3802 (N_3802,N_3722,N_3264);
nand U3803 (N_3803,N_3186,N_3247);
nand U3804 (N_3804,N_3425,N_3200);
xnor U3805 (N_3805,N_3273,N_3697);
nand U3806 (N_3806,N_3525,N_3628);
or U3807 (N_3807,N_3441,N_3162);
and U3808 (N_3808,N_3209,N_3612);
and U3809 (N_3809,N_3351,N_3691);
and U3810 (N_3810,N_3693,N_3521);
and U3811 (N_3811,N_3369,N_3316);
nand U3812 (N_3812,N_3662,N_3620);
or U3813 (N_3813,N_3320,N_3486);
or U3814 (N_3814,N_3717,N_3307);
and U3815 (N_3815,N_3469,N_3562);
xnor U3816 (N_3816,N_3375,N_3158);
xor U3817 (N_3817,N_3207,N_3541);
nor U3818 (N_3818,N_3147,N_3606);
nor U3819 (N_3819,N_3687,N_3321);
xnor U3820 (N_3820,N_3367,N_3252);
or U3821 (N_3821,N_3383,N_3128);
and U3822 (N_3822,N_3381,N_3688);
nand U3823 (N_3823,N_3426,N_3743);
nand U3824 (N_3824,N_3216,N_3468);
nor U3825 (N_3825,N_3694,N_3557);
or U3826 (N_3826,N_3411,N_3704);
xnor U3827 (N_3827,N_3446,N_3568);
nor U3828 (N_3828,N_3668,N_3340);
and U3829 (N_3829,N_3380,N_3516);
or U3830 (N_3830,N_3644,N_3311);
nand U3831 (N_3831,N_3403,N_3600);
and U3832 (N_3832,N_3415,N_3591);
and U3833 (N_3833,N_3664,N_3749);
xor U3834 (N_3834,N_3213,N_3386);
and U3835 (N_3835,N_3746,N_3592);
and U3836 (N_3836,N_3163,N_3310);
nand U3837 (N_3837,N_3191,N_3176);
xnor U3838 (N_3838,N_3338,N_3399);
and U3839 (N_3839,N_3342,N_3626);
xnor U3840 (N_3840,N_3168,N_3167);
and U3841 (N_3841,N_3195,N_3734);
or U3842 (N_3842,N_3608,N_3666);
and U3843 (N_3843,N_3667,N_3483);
xor U3844 (N_3844,N_3129,N_3454);
xnor U3845 (N_3845,N_3493,N_3393);
nand U3846 (N_3846,N_3187,N_3363);
and U3847 (N_3847,N_3481,N_3735);
xnor U3848 (N_3848,N_3545,N_3409);
or U3849 (N_3849,N_3582,N_3642);
nand U3850 (N_3850,N_3546,N_3569);
nand U3851 (N_3851,N_3277,N_3157);
or U3852 (N_3852,N_3701,N_3561);
or U3853 (N_3853,N_3617,N_3269);
nand U3854 (N_3854,N_3249,N_3661);
and U3855 (N_3855,N_3513,N_3387);
and U3856 (N_3856,N_3239,N_3529);
xnor U3857 (N_3857,N_3442,N_3604);
xor U3858 (N_3858,N_3679,N_3322);
nand U3859 (N_3859,N_3711,N_3499);
nand U3860 (N_3860,N_3506,N_3496);
xnor U3861 (N_3861,N_3268,N_3744);
nand U3862 (N_3862,N_3543,N_3527);
nand U3863 (N_3863,N_3570,N_3488);
or U3864 (N_3864,N_3226,N_3285);
xor U3865 (N_3865,N_3306,N_3256);
and U3866 (N_3866,N_3517,N_3127);
and U3867 (N_3867,N_3246,N_3726);
xor U3868 (N_3868,N_3723,N_3328);
nor U3869 (N_3869,N_3391,N_3401);
nor U3870 (N_3870,N_3535,N_3736);
nor U3871 (N_3871,N_3473,N_3374);
nand U3872 (N_3872,N_3339,N_3184);
and U3873 (N_3873,N_3312,N_3331);
xnor U3874 (N_3874,N_3413,N_3737);
nand U3875 (N_3875,N_3408,N_3194);
or U3876 (N_3876,N_3192,N_3166);
nor U3877 (N_3877,N_3287,N_3482);
xor U3878 (N_3878,N_3333,N_3319);
xor U3879 (N_3879,N_3497,N_3629);
nand U3880 (N_3880,N_3263,N_3555);
and U3881 (N_3881,N_3705,N_3669);
or U3882 (N_3882,N_3296,N_3344);
nor U3883 (N_3883,N_3281,N_3739);
nand U3884 (N_3884,N_3325,N_3706);
or U3885 (N_3885,N_3149,N_3689);
nor U3886 (N_3886,N_3699,N_3272);
nand U3887 (N_3887,N_3447,N_3500);
and U3888 (N_3888,N_3421,N_3586);
nand U3889 (N_3889,N_3394,N_3225);
xnor U3890 (N_3890,N_3730,N_3443);
or U3891 (N_3891,N_3148,N_3266);
nor U3892 (N_3892,N_3231,N_3715);
xor U3893 (N_3893,N_3475,N_3650);
or U3894 (N_3894,N_3466,N_3259);
or U3895 (N_3895,N_3512,N_3397);
nand U3896 (N_3896,N_3365,N_3278);
and U3897 (N_3897,N_3171,N_3313);
and U3898 (N_3898,N_3405,N_3508);
nor U3899 (N_3899,N_3242,N_3199);
nand U3900 (N_3900,N_3532,N_3720);
xnor U3901 (N_3901,N_3554,N_3690);
and U3902 (N_3902,N_3202,N_3430);
nand U3903 (N_3903,N_3738,N_3605);
and U3904 (N_3904,N_3435,N_3639);
or U3905 (N_3905,N_3424,N_3233);
or U3906 (N_3906,N_3610,N_3220);
nand U3907 (N_3907,N_3707,N_3710);
and U3908 (N_3908,N_3302,N_3125);
xnor U3909 (N_3909,N_3388,N_3358);
or U3910 (N_3910,N_3323,N_3507);
or U3911 (N_3911,N_3248,N_3294);
nor U3912 (N_3912,N_3197,N_3474);
and U3913 (N_3913,N_3254,N_3601);
or U3914 (N_3914,N_3613,N_3641);
xnor U3915 (N_3915,N_3151,N_3286);
or U3916 (N_3916,N_3492,N_3412);
nand U3917 (N_3917,N_3464,N_3317);
and U3918 (N_3918,N_3593,N_3185);
and U3919 (N_3919,N_3686,N_3649);
xnor U3920 (N_3920,N_3161,N_3336);
xnor U3921 (N_3921,N_3652,N_3228);
and U3922 (N_3922,N_3627,N_3131);
and U3923 (N_3923,N_3700,N_3329);
nor U3924 (N_3924,N_3484,N_3537);
nor U3925 (N_3925,N_3681,N_3159);
nand U3926 (N_3926,N_3139,N_3732);
nor U3927 (N_3927,N_3208,N_3245);
xor U3928 (N_3928,N_3189,N_3183);
xnor U3929 (N_3929,N_3250,N_3164);
or U3930 (N_3930,N_3410,N_3217);
or U3931 (N_3931,N_3657,N_3144);
nor U3932 (N_3932,N_3382,N_3126);
and U3933 (N_3933,N_3427,N_3172);
or U3934 (N_3934,N_3615,N_3571);
and U3935 (N_3935,N_3190,N_3364);
nand U3936 (N_3936,N_3352,N_3227);
and U3937 (N_3937,N_3471,N_3637);
nor U3938 (N_3938,N_3614,N_3575);
xnor U3939 (N_3939,N_3547,N_3457);
nor U3940 (N_3940,N_3132,N_3658);
nor U3941 (N_3941,N_3324,N_3616);
nor U3942 (N_3942,N_3280,N_3439);
or U3943 (N_3943,N_3154,N_3326);
nand U3944 (N_3944,N_3623,N_3459);
nor U3945 (N_3945,N_3193,N_3747);
nor U3946 (N_3946,N_3206,N_3713);
nor U3947 (N_3947,N_3740,N_3211);
nor U3948 (N_3948,N_3692,N_3451);
and U3949 (N_3949,N_3479,N_3156);
and U3950 (N_3950,N_3433,N_3350);
or U3951 (N_3951,N_3330,N_3542);
nor U3952 (N_3952,N_3708,N_3472);
or U3953 (N_3953,N_3334,N_3179);
nand U3954 (N_3954,N_3456,N_3152);
nor U3955 (N_3955,N_3232,N_3354);
or U3956 (N_3956,N_3345,N_3463);
or U3957 (N_3957,N_3214,N_3520);
nor U3958 (N_3958,N_3262,N_3414);
and U3959 (N_3959,N_3581,N_3240);
nand U3960 (N_3960,N_3373,N_3449);
nor U3961 (N_3961,N_3341,N_3534);
xor U3962 (N_3962,N_3181,N_3670);
xor U3963 (N_3963,N_3275,N_3210);
and U3964 (N_3964,N_3611,N_3609);
xnor U3965 (N_3965,N_3539,N_3327);
or U3966 (N_3966,N_3619,N_3141);
nor U3967 (N_3967,N_3267,N_3284);
and U3968 (N_3968,N_3455,N_3362);
and U3969 (N_3969,N_3289,N_3596);
nor U3970 (N_3970,N_3643,N_3503);
and U3971 (N_3971,N_3523,N_3460);
nor U3972 (N_3972,N_3522,N_3419);
xnor U3973 (N_3973,N_3279,N_3607);
nand U3974 (N_3974,N_3404,N_3510);
nor U3975 (N_3975,N_3188,N_3137);
nand U3976 (N_3976,N_3636,N_3297);
and U3977 (N_3977,N_3238,N_3489);
nand U3978 (N_3978,N_3450,N_3651);
nand U3979 (N_3979,N_3377,N_3725);
xnor U3980 (N_3980,N_3654,N_3130);
or U3981 (N_3981,N_3742,N_3685);
and U3982 (N_3982,N_3549,N_3274);
or U3983 (N_3983,N_3429,N_3458);
and U3984 (N_3984,N_3175,N_3576);
or U3985 (N_3985,N_3136,N_3635);
nand U3986 (N_3986,N_3360,N_3748);
or U3987 (N_3987,N_3544,N_3353);
and U3988 (N_3988,N_3359,N_3504);
xor U3989 (N_3989,N_3622,N_3526);
or U3990 (N_3990,N_3169,N_3646);
or U3991 (N_3991,N_3672,N_3518);
nor U3992 (N_3992,N_3418,N_3292);
nor U3993 (N_3993,N_3203,N_3656);
nand U3994 (N_3994,N_3599,N_3253);
or U3995 (N_3995,N_3524,N_3445);
nand U3996 (N_3996,N_3564,N_3476);
and U3997 (N_3997,N_3501,N_3553);
and U3998 (N_3998,N_3398,N_3556);
nor U3999 (N_3999,N_3142,N_3145);
and U4000 (N_4000,N_3205,N_3237);
xnor U4001 (N_4001,N_3514,N_3416);
nand U4002 (N_4002,N_3349,N_3487);
and U4003 (N_4003,N_3716,N_3674);
xnor U4004 (N_4004,N_3230,N_3198);
nor U4005 (N_4005,N_3584,N_3552);
or U4006 (N_4006,N_3229,N_3724);
and U4007 (N_4007,N_3567,N_3434);
nand U4008 (N_4008,N_3583,N_3407);
xor U4009 (N_4009,N_3540,N_3165);
nand U4010 (N_4010,N_3223,N_3236);
and U4011 (N_4011,N_3566,N_3703);
or U4012 (N_4012,N_3625,N_3219);
nand U4013 (N_4013,N_3602,N_3417);
or U4014 (N_4014,N_3244,N_3218);
xnor U4015 (N_4015,N_3663,N_3647);
nand U4016 (N_4016,N_3638,N_3511);
nand U4017 (N_4017,N_3133,N_3580);
nand U4018 (N_4018,N_3385,N_3174);
xor U4019 (N_4019,N_3665,N_3221);
xor U4020 (N_4020,N_3550,N_3283);
xor U4021 (N_4021,N_3258,N_3348);
or U4022 (N_4022,N_3173,N_3485);
nor U4023 (N_4023,N_3257,N_3587);
nor U4024 (N_4024,N_3315,N_3498);
nor U4025 (N_4025,N_3618,N_3624);
or U4026 (N_4026,N_3308,N_3490);
xor U4027 (N_4027,N_3572,N_3632);
xnor U4028 (N_4028,N_3590,N_3234);
and U4029 (N_4029,N_3640,N_3671);
or U4030 (N_4030,N_3530,N_3371);
xor U4031 (N_4031,N_3347,N_3346);
and U4032 (N_4032,N_3676,N_3551);
nand U4033 (N_4033,N_3241,N_3630);
nor U4034 (N_4034,N_3696,N_3505);
or U4035 (N_4035,N_3588,N_3431);
xnor U4036 (N_4036,N_3495,N_3436);
xnor U4037 (N_4037,N_3729,N_3477);
and U4038 (N_4038,N_3558,N_3633);
and U4039 (N_4039,N_3215,N_3480);
nor U4040 (N_4040,N_3438,N_3682);
or U4041 (N_4041,N_3603,N_3406);
nand U4042 (N_4042,N_3304,N_3300);
and U4043 (N_4043,N_3196,N_3155);
nor U4044 (N_4044,N_3731,N_3357);
xor U4045 (N_4045,N_3683,N_3332);
or U4046 (N_4046,N_3559,N_3519);
xnor U4047 (N_4047,N_3594,N_3675);
or U4048 (N_4048,N_3153,N_3714);
nand U4049 (N_4049,N_3305,N_3368);
nand U4050 (N_4050,N_3444,N_3396);
or U4051 (N_4051,N_3465,N_3684);
nor U4052 (N_4052,N_3291,N_3437);
nand U4053 (N_4053,N_3595,N_3178);
xnor U4054 (N_4054,N_3727,N_3533);
nor U4055 (N_4055,N_3428,N_3578);
xnor U4056 (N_4056,N_3659,N_3577);
nand U4057 (N_4057,N_3440,N_3265);
xor U4058 (N_4058,N_3290,N_3356);
and U4059 (N_4059,N_3478,N_3448);
nand U4060 (N_4060,N_3563,N_3138);
and U4061 (N_4061,N_3719,N_3295);
or U4062 (N_4062,N_3470,N_3643);
or U4063 (N_4063,N_3537,N_3647);
and U4064 (N_4064,N_3438,N_3648);
and U4065 (N_4065,N_3135,N_3557);
and U4066 (N_4066,N_3134,N_3563);
or U4067 (N_4067,N_3399,N_3678);
xnor U4068 (N_4068,N_3217,N_3584);
or U4069 (N_4069,N_3332,N_3175);
xnor U4070 (N_4070,N_3655,N_3211);
and U4071 (N_4071,N_3453,N_3168);
nand U4072 (N_4072,N_3489,N_3552);
and U4073 (N_4073,N_3748,N_3405);
and U4074 (N_4074,N_3216,N_3125);
xor U4075 (N_4075,N_3670,N_3539);
and U4076 (N_4076,N_3511,N_3460);
or U4077 (N_4077,N_3741,N_3339);
and U4078 (N_4078,N_3500,N_3536);
nand U4079 (N_4079,N_3393,N_3563);
nand U4080 (N_4080,N_3202,N_3523);
nor U4081 (N_4081,N_3152,N_3175);
nor U4082 (N_4082,N_3381,N_3592);
or U4083 (N_4083,N_3685,N_3322);
and U4084 (N_4084,N_3498,N_3690);
nor U4085 (N_4085,N_3704,N_3290);
xnor U4086 (N_4086,N_3301,N_3663);
or U4087 (N_4087,N_3561,N_3596);
nor U4088 (N_4088,N_3329,N_3737);
and U4089 (N_4089,N_3601,N_3649);
nor U4090 (N_4090,N_3619,N_3578);
nand U4091 (N_4091,N_3525,N_3394);
or U4092 (N_4092,N_3554,N_3204);
xnor U4093 (N_4093,N_3160,N_3412);
nand U4094 (N_4094,N_3677,N_3136);
and U4095 (N_4095,N_3310,N_3684);
nor U4096 (N_4096,N_3201,N_3637);
or U4097 (N_4097,N_3293,N_3439);
xnor U4098 (N_4098,N_3565,N_3645);
and U4099 (N_4099,N_3271,N_3596);
nand U4100 (N_4100,N_3674,N_3406);
nor U4101 (N_4101,N_3358,N_3396);
xnor U4102 (N_4102,N_3556,N_3705);
xnor U4103 (N_4103,N_3690,N_3234);
xnor U4104 (N_4104,N_3212,N_3679);
or U4105 (N_4105,N_3682,N_3498);
nor U4106 (N_4106,N_3421,N_3222);
nor U4107 (N_4107,N_3229,N_3230);
and U4108 (N_4108,N_3670,N_3185);
nor U4109 (N_4109,N_3516,N_3407);
and U4110 (N_4110,N_3622,N_3153);
and U4111 (N_4111,N_3194,N_3400);
xor U4112 (N_4112,N_3662,N_3453);
or U4113 (N_4113,N_3172,N_3478);
xnor U4114 (N_4114,N_3395,N_3235);
nand U4115 (N_4115,N_3349,N_3178);
or U4116 (N_4116,N_3442,N_3265);
and U4117 (N_4117,N_3131,N_3555);
or U4118 (N_4118,N_3557,N_3249);
nor U4119 (N_4119,N_3438,N_3188);
nand U4120 (N_4120,N_3160,N_3201);
nand U4121 (N_4121,N_3342,N_3356);
or U4122 (N_4122,N_3536,N_3330);
and U4123 (N_4123,N_3365,N_3322);
nor U4124 (N_4124,N_3514,N_3405);
nand U4125 (N_4125,N_3440,N_3218);
and U4126 (N_4126,N_3229,N_3726);
xor U4127 (N_4127,N_3285,N_3735);
nor U4128 (N_4128,N_3428,N_3608);
nor U4129 (N_4129,N_3387,N_3718);
or U4130 (N_4130,N_3632,N_3507);
nand U4131 (N_4131,N_3739,N_3650);
xnor U4132 (N_4132,N_3595,N_3591);
xor U4133 (N_4133,N_3404,N_3391);
or U4134 (N_4134,N_3625,N_3269);
nand U4135 (N_4135,N_3406,N_3292);
nand U4136 (N_4136,N_3397,N_3264);
and U4137 (N_4137,N_3220,N_3739);
or U4138 (N_4138,N_3161,N_3335);
xor U4139 (N_4139,N_3641,N_3734);
nor U4140 (N_4140,N_3240,N_3697);
or U4141 (N_4141,N_3171,N_3565);
and U4142 (N_4142,N_3214,N_3657);
nand U4143 (N_4143,N_3632,N_3440);
xor U4144 (N_4144,N_3670,N_3544);
nand U4145 (N_4145,N_3183,N_3364);
xnor U4146 (N_4146,N_3251,N_3482);
or U4147 (N_4147,N_3570,N_3292);
or U4148 (N_4148,N_3670,N_3519);
nor U4149 (N_4149,N_3616,N_3156);
or U4150 (N_4150,N_3396,N_3470);
nor U4151 (N_4151,N_3327,N_3511);
nand U4152 (N_4152,N_3629,N_3203);
or U4153 (N_4153,N_3686,N_3530);
or U4154 (N_4154,N_3471,N_3166);
nor U4155 (N_4155,N_3435,N_3155);
xor U4156 (N_4156,N_3749,N_3172);
nor U4157 (N_4157,N_3363,N_3229);
or U4158 (N_4158,N_3414,N_3697);
and U4159 (N_4159,N_3134,N_3413);
or U4160 (N_4160,N_3126,N_3312);
nand U4161 (N_4161,N_3468,N_3225);
nand U4162 (N_4162,N_3607,N_3559);
xor U4163 (N_4163,N_3653,N_3296);
and U4164 (N_4164,N_3392,N_3282);
and U4165 (N_4165,N_3240,N_3367);
or U4166 (N_4166,N_3727,N_3142);
or U4167 (N_4167,N_3178,N_3337);
and U4168 (N_4168,N_3321,N_3374);
xnor U4169 (N_4169,N_3373,N_3129);
and U4170 (N_4170,N_3699,N_3184);
nor U4171 (N_4171,N_3641,N_3619);
xor U4172 (N_4172,N_3246,N_3465);
or U4173 (N_4173,N_3745,N_3273);
nand U4174 (N_4174,N_3748,N_3305);
or U4175 (N_4175,N_3326,N_3185);
xnor U4176 (N_4176,N_3278,N_3665);
xor U4177 (N_4177,N_3460,N_3725);
xor U4178 (N_4178,N_3430,N_3475);
or U4179 (N_4179,N_3486,N_3749);
xor U4180 (N_4180,N_3723,N_3579);
nand U4181 (N_4181,N_3601,N_3471);
nor U4182 (N_4182,N_3452,N_3282);
or U4183 (N_4183,N_3427,N_3638);
and U4184 (N_4184,N_3643,N_3654);
xnor U4185 (N_4185,N_3424,N_3215);
and U4186 (N_4186,N_3128,N_3355);
nor U4187 (N_4187,N_3292,N_3679);
nand U4188 (N_4188,N_3440,N_3417);
or U4189 (N_4189,N_3249,N_3284);
and U4190 (N_4190,N_3740,N_3525);
nor U4191 (N_4191,N_3208,N_3610);
nor U4192 (N_4192,N_3565,N_3163);
xnor U4193 (N_4193,N_3582,N_3612);
and U4194 (N_4194,N_3356,N_3355);
xor U4195 (N_4195,N_3425,N_3695);
nand U4196 (N_4196,N_3650,N_3263);
or U4197 (N_4197,N_3600,N_3444);
and U4198 (N_4198,N_3367,N_3687);
nand U4199 (N_4199,N_3530,N_3516);
and U4200 (N_4200,N_3152,N_3447);
nor U4201 (N_4201,N_3701,N_3640);
xor U4202 (N_4202,N_3166,N_3220);
or U4203 (N_4203,N_3261,N_3139);
xnor U4204 (N_4204,N_3671,N_3277);
nor U4205 (N_4205,N_3557,N_3147);
or U4206 (N_4206,N_3476,N_3221);
or U4207 (N_4207,N_3197,N_3187);
nor U4208 (N_4208,N_3586,N_3462);
and U4209 (N_4209,N_3666,N_3657);
xor U4210 (N_4210,N_3228,N_3574);
nand U4211 (N_4211,N_3352,N_3660);
or U4212 (N_4212,N_3552,N_3716);
and U4213 (N_4213,N_3350,N_3591);
nor U4214 (N_4214,N_3446,N_3614);
xnor U4215 (N_4215,N_3156,N_3155);
xnor U4216 (N_4216,N_3578,N_3195);
nand U4217 (N_4217,N_3663,N_3656);
and U4218 (N_4218,N_3343,N_3372);
or U4219 (N_4219,N_3198,N_3669);
xor U4220 (N_4220,N_3551,N_3441);
nand U4221 (N_4221,N_3347,N_3399);
or U4222 (N_4222,N_3460,N_3249);
nor U4223 (N_4223,N_3547,N_3666);
nor U4224 (N_4224,N_3295,N_3726);
xor U4225 (N_4225,N_3130,N_3611);
xnor U4226 (N_4226,N_3198,N_3272);
nor U4227 (N_4227,N_3263,N_3673);
nand U4228 (N_4228,N_3389,N_3195);
and U4229 (N_4229,N_3341,N_3701);
and U4230 (N_4230,N_3747,N_3353);
xor U4231 (N_4231,N_3390,N_3167);
and U4232 (N_4232,N_3665,N_3173);
nand U4233 (N_4233,N_3534,N_3326);
xor U4234 (N_4234,N_3245,N_3547);
nor U4235 (N_4235,N_3606,N_3379);
xor U4236 (N_4236,N_3314,N_3691);
nand U4237 (N_4237,N_3589,N_3735);
xor U4238 (N_4238,N_3420,N_3465);
and U4239 (N_4239,N_3353,N_3490);
nor U4240 (N_4240,N_3406,N_3670);
nor U4241 (N_4241,N_3493,N_3191);
nor U4242 (N_4242,N_3231,N_3376);
nand U4243 (N_4243,N_3691,N_3365);
xnor U4244 (N_4244,N_3510,N_3461);
nor U4245 (N_4245,N_3374,N_3177);
and U4246 (N_4246,N_3486,N_3437);
nand U4247 (N_4247,N_3585,N_3535);
and U4248 (N_4248,N_3544,N_3739);
or U4249 (N_4249,N_3476,N_3367);
and U4250 (N_4250,N_3386,N_3398);
and U4251 (N_4251,N_3352,N_3454);
nand U4252 (N_4252,N_3236,N_3377);
nor U4253 (N_4253,N_3588,N_3377);
and U4254 (N_4254,N_3568,N_3170);
xor U4255 (N_4255,N_3374,N_3425);
or U4256 (N_4256,N_3541,N_3520);
nor U4257 (N_4257,N_3588,N_3332);
xor U4258 (N_4258,N_3320,N_3579);
and U4259 (N_4259,N_3656,N_3200);
nand U4260 (N_4260,N_3622,N_3158);
nor U4261 (N_4261,N_3355,N_3331);
and U4262 (N_4262,N_3547,N_3707);
xnor U4263 (N_4263,N_3684,N_3451);
nand U4264 (N_4264,N_3668,N_3575);
or U4265 (N_4265,N_3379,N_3314);
nand U4266 (N_4266,N_3695,N_3656);
nor U4267 (N_4267,N_3722,N_3626);
nor U4268 (N_4268,N_3201,N_3211);
xnor U4269 (N_4269,N_3416,N_3170);
and U4270 (N_4270,N_3473,N_3230);
nand U4271 (N_4271,N_3135,N_3439);
xnor U4272 (N_4272,N_3217,N_3261);
xor U4273 (N_4273,N_3270,N_3296);
or U4274 (N_4274,N_3246,N_3430);
nand U4275 (N_4275,N_3245,N_3183);
nor U4276 (N_4276,N_3335,N_3698);
xor U4277 (N_4277,N_3515,N_3561);
and U4278 (N_4278,N_3558,N_3722);
nand U4279 (N_4279,N_3485,N_3220);
and U4280 (N_4280,N_3304,N_3685);
nand U4281 (N_4281,N_3268,N_3683);
xor U4282 (N_4282,N_3323,N_3489);
or U4283 (N_4283,N_3387,N_3413);
xnor U4284 (N_4284,N_3735,N_3146);
xnor U4285 (N_4285,N_3296,N_3578);
nand U4286 (N_4286,N_3241,N_3432);
nor U4287 (N_4287,N_3255,N_3207);
xor U4288 (N_4288,N_3361,N_3414);
xor U4289 (N_4289,N_3155,N_3730);
or U4290 (N_4290,N_3605,N_3165);
or U4291 (N_4291,N_3250,N_3277);
nor U4292 (N_4292,N_3558,N_3201);
and U4293 (N_4293,N_3310,N_3331);
xnor U4294 (N_4294,N_3392,N_3144);
xor U4295 (N_4295,N_3152,N_3538);
or U4296 (N_4296,N_3143,N_3667);
or U4297 (N_4297,N_3565,N_3342);
xnor U4298 (N_4298,N_3260,N_3334);
or U4299 (N_4299,N_3527,N_3399);
nor U4300 (N_4300,N_3740,N_3205);
nand U4301 (N_4301,N_3705,N_3357);
nand U4302 (N_4302,N_3645,N_3187);
nor U4303 (N_4303,N_3546,N_3686);
nor U4304 (N_4304,N_3680,N_3187);
xnor U4305 (N_4305,N_3219,N_3307);
xor U4306 (N_4306,N_3667,N_3661);
and U4307 (N_4307,N_3394,N_3736);
nor U4308 (N_4308,N_3565,N_3622);
xor U4309 (N_4309,N_3375,N_3218);
nand U4310 (N_4310,N_3361,N_3403);
and U4311 (N_4311,N_3242,N_3369);
nor U4312 (N_4312,N_3387,N_3176);
xnor U4313 (N_4313,N_3627,N_3156);
and U4314 (N_4314,N_3562,N_3128);
nand U4315 (N_4315,N_3569,N_3461);
nand U4316 (N_4316,N_3681,N_3214);
nand U4317 (N_4317,N_3415,N_3546);
or U4318 (N_4318,N_3505,N_3481);
nand U4319 (N_4319,N_3139,N_3669);
and U4320 (N_4320,N_3571,N_3277);
or U4321 (N_4321,N_3560,N_3236);
and U4322 (N_4322,N_3482,N_3322);
and U4323 (N_4323,N_3487,N_3506);
nand U4324 (N_4324,N_3577,N_3275);
nand U4325 (N_4325,N_3195,N_3531);
nand U4326 (N_4326,N_3719,N_3638);
and U4327 (N_4327,N_3195,N_3261);
nor U4328 (N_4328,N_3479,N_3747);
or U4329 (N_4329,N_3468,N_3237);
and U4330 (N_4330,N_3707,N_3361);
or U4331 (N_4331,N_3436,N_3602);
nor U4332 (N_4332,N_3698,N_3749);
nor U4333 (N_4333,N_3257,N_3640);
nor U4334 (N_4334,N_3284,N_3542);
or U4335 (N_4335,N_3697,N_3268);
or U4336 (N_4336,N_3313,N_3218);
or U4337 (N_4337,N_3458,N_3658);
or U4338 (N_4338,N_3573,N_3516);
and U4339 (N_4339,N_3197,N_3324);
and U4340 (N_4340,N_3374,N_3285);
nand U4341 (N_4341,N_3749,N_3744);
nor U4342 (N_4342,N_3405,N_3430);
or U4343 (N_4343,N_3247,N_3600);
xnor U4344 (N_4344,N_3235,N_3629);
nand U4345 (N_4345,N_3703,N_3537);
or U4346 (N_4346,N_3582,N_3484);
nor U4347 (N_4347,N_3343,N_3545);
or U4348 (N_4348,N_3247,N_3206);
xnor U4349 (N_4349,N_3741,N_3490);
nand U4350 (N_4350,N_3703,N_3511);
nand U4351 (N_4351,N_3432,N_3526);
or U4352 (N_4352,N_3541,N_3709);
xnor U4353 (N_4353,N_3508,N_3265);
or U4354 (N_4354,N_3259,N_3676);
and U4355 (N_4355,N_3214,N_3544);
and U4356 (N_4356,N_3379,N_3511);
nor U4357 (N_4357,N_3744,N_3440);
nor U4358 (N_4358,N_3555,N_3528);
nor U4359 (N_4359,N_3326,N_3474);
and U4360 (N_4360,N_3356,N_3363);
or U4361 (N_4361,N_3685,N_3610);
nand U4362 (N_4362,N_3125,N_3321);
and U4363 (N_4363,N_3190,N_3582);
or U4364 (N_4364,N_3673,N_3514);
xnor U4365 (N_4365,N_3419,N_3173);
nor U4366 (N_4366,N_3374,N_3369);
xnor U4367 (N_4367,N_3537,N_3683);
and U4368 (N_4368,N_3680,N_3388);
xor U4369 (N_4369,N_3584,N_3165);
xnor U4370 (N_4370,N_3330,N_3127);
nor U4371 (N_4371,N_3234,N_3517);
or U4372 (N_4372,N_3336,N_3339);
and U4373 (N_4373,N_3644,N_3126);
or U4374 (N_4374,N_3197,N_3413);
nor U4375 (N_4375,N_4059,N_4024);
nand U4376 (N_4376,N_4084,N_3951);
nor U4377 (N_4377,N_4270,N_3945);
or U4378 (N_4378,N_3788,N_3810);
nand U4379 (N_4379,N_3978,N_3787);
and U4380 (N_4380,N_3928,N_4208);
and U4381 (N_4381,N_3864,N_4302);
and U4382 (N_4382,N_4345,N_4049);
or U4383 (N_4383,N_4115,N_3897);
and U4384 (N_4384,N_3910,N_3896);
xor U4385 (N_4385,N_4308,N_3819);
nand U4386 (N_4386,N_3801,N_3992);
and U4387 (N_4387,N_4187,N_4040);
xor U4388 (N_4388,N_4082,N_4317);
nor U4389 (N_4389,N_3957,N_3922);
or U4390 (N_4390,N_3885,N_3880);
nand U4391 (N_4391,N_4031,N_4069);
or U4392 (N_4392,N_4287,N_3994);
nand U4393 (N_4393,N_3866,N_3777);
xor U4394 (N_4394,N_4130,N_4075);
xnor U4395 (N_4395,N_4001,N_3848);
nor U4396 (N_4396,N_3867,N_3861);
nand U4397 (N_4397,N_4291,N_4335);
or U4398 (N_4398,N_4227,N_3751);
or U4399 (N_4399,N_4285,N_4260);
nand U4400 (N_4400,N_3981,N_4177);
or U4401 (N_4401,N_4361,N_3761);
or U4402 (N_4402,N_3937,N_4117);
xnor U4403 (N_4403,N_4062,N_4162);
or U4404 (N_4404,N_3758,N_4307);
or U4405 (N_4405,N_4102,N_4172);
xor U4406 (N_4406,N_3927,N_3948);
and U4407 (N_4407,N_4171,N_3956);
or U4408 (N_4408,N_3841,N_4006);
nand U4409 (N_4409,N_3825,N_4201);
xor U4410 (N_4410,N_4222,N_3915);
and U4411 (N_4411,N_4267,N_3916);
xor U4412 (N_4412,N_3862,N_4218);
nor U4413 (N_4413,N_4211,N_3795);
or U4414 (N_4414,N_3934,N_4044);
or U4415 (N_4415,N_4026,N_3844);
and U4416 (N_4416,N_3797,N_4093);
nand U4417 (N_4417,N_4158,N_4119);
nand U4418 (N_4418,N_4118,N_4078);
xnor U4419 (N_4419,N_4165,N_4322);
or U4420 (N_4420,N_3813,N_3771);
nand U4421 (N_4421,N_4089,N_4099);
or U4422 (N_4422,N_3925,N_4304);
nand U4423 (N_4423,N_4209,N_4163);
xor U4424 (N_4424,N_3857,N_4116);
xor U4425 (N_4425,N_3832,N_3838);
or U4426 (N_4426,N_3875,N_4139);
and U4427 (N_4427,N_4124,N_4083);
xnor U4428 (N_4428,N_4330,N_4202);
and U4429 (N_4429,N_4252,N_4255);
xnor U4430 (N_4430,N_3851,N_4053);
and U4431 (N_4431,N_3886,N_4297);
nand U4432 (N_4432,N_4253,N_4323);
and U4433 (N_4433,N_3939,N_3753);
nor U4434 (N_4434,N_4238,N_4166);
nor U4435 (N_4435,N_4348,N_4232);
and U4436 (N_4436,N_4319,N_3828);
nand U4437 (N_4437,N_4245,N_3871);
nand U4438 (N_4438,N_3873,N_4101);
or U4439 (N_4439,N_4204,N_4045);
nor U4440 (N_4440,N_4284,N_4217);
nor U4441 (N_4441,N_3970,N_4196);
xnor U4442 (N_4442,N_3966,N_3865);
and U4443 (N_4443,N_3878,N_4262);
and U4444 (N_4444,N_4157,N_4122);
nor U4445 (N_4445,N_3911,N_3772);
xor U4446 (N_4446,N_4133,N_4242);
and U4447 (N_4447,N_3755,N_3764);
xnor U4448 (N_4448,N_4339,N_3997);
xnor U4449 (N_4449,N_4243,N_4263);
nor U4450 (N_4450,N_3768,N_4344);
nor U4451 (N_4451,N_4336,N_4364);
nor U4452 (N_4452,N_4250,N_4257);
or U4453 (N_4453,N_4184,N_3954);
xnor U4454 (N_4454,N_4025,N_4131);
nand U4455 (N_4455,N_4015,N_4363);
and U4456 (N_4456,N_3996,N_4220);
and U4457 (N_4457,N_3808,N_4321);
nand U4458 (N_4458,N_4318,N_4332);
nor U4459 (N_4459,N_3998,N_4090);
xnor U4460 (N_4460,N_3993,N_4138);
xor U4461 (N_4461,N_3868,N_3863);
xnor U4462 (N_4462,N_4316,N_4000);
nor U4463 (N_4463,N_4228,N_3932);
nor U4464 (N_4464,N_3971,N_3952);
nand U4465 (N_4465,N_3960,N_4215);
nor U4466 (N_4466,N_4343,N_3869);
nor U4467 (N_4467,N_4074,N_4351);
nand U4468 (N_4468,N_3858,N_4023);
nor U4469 (N_4469,N_3909,N_3923);
xnor U4470 (N_4470,N_3983,N_4374);
or U4471 (N_4471,N_4106,N_3890);
nor U4472 (N_4472,N_3982,N_4098);
nor U4473 (N_4473,N_3941,N_4367);
and U4474 (N_4474,N_4362,N_3756);
and U4475 (N_4475,N_3826,N_4181);
and U4476 (N_4476,N_4047,N_4065);
or U4477 (N_4477,N_4096,N_4290);
xor U4478 (N_4478,N_4027,N_4155);
xnor U4479 (N_4479,N_4070,N_4142);
or U4480 (N_4480,N_3955,N_4219);
nor U4481 (N_4481,N_4055,N_4046);
and U4482 (N_4482,N_4173,N_3822);
or U4483 (N_4483,N_3882,N_3750);
nand U4484 (N_4484,N_3892,N_4340);
nand U4485 (N_4485,N_4246,N_4357);
nand U4486 (N_4486,N_3965,N_4016);
and U4487 (N_4487,N_3818,N_4329);
and U4488 (N_4488,N_4085,N_4347);
nor U4489 (N_4489,N_4301,N_4239);
or U4490 (N_4490,N_3918,N_3985);
and U4491 (N_4491,N_3847,N_4300);
nor U4492 (N_4492,N_3906,N_4033);
and U4493 (N_4493,N_3969,N_4261);
nor U4494 (N_4494,N_4198,N_3975);
xor U4495 (N_4495,N_4273,N_4146);
xor U4496 (N_4496,N_3814,N_4052);
nand U4497 (N_4497,N_3933,N_4058);
nand U4498 (N_4498,N_3762,N_4168);
xnor U4499 (N_4499,N_4354,N_3757);
xor U4500 (N_4500,N_4128,N_3840);
nor U4501 (N_4501,N_3977,N_4152);
nor U4502 (N_4502,N_4254,N_4210);
xor U4503 (N_4503,N_4141,N_3999);
or U4504 (N_4504,N_3926,N_3876);
or U4505 (N_4505,N_4022,N_3835);
or U4506 (N_4506,N_4021,N_4009);
and U4507 (N_4507,N_4034,N_4154);
nand U4508 (N_4508,N_3799,N_3782);
or U4509 (N_4509,N_3831,N_4278);
and U4510 (N_4510,N_4236,N_4226);
nor U4511 (N_4511,N_3779,N_4274);
xnor U4512 (N_4512,N_3806,N_4327);
or U4513 (N_4513,N_3938,N_4043);
and U4514 (N_4514,N_4160,N_4346);
nand U4515 (N_4515,N_4235,N_4003);
or U4516 (N_4516,N_4081,N_3776);
nand U4517 (N_4517,N_4237,N_4071);
xnor U4518 (N_4518,N_4352,N_4234);
nand U4519 (N_4519,N_3907,N_4265);
nor U4520 (N_4520,N_4275,N_3839);
xnor U4521 (N_4521,N_4251,N_3827);
nor U4522 (N_4522,N_4143,N_3765);
and U4523 (N_4523,N_3879,N_3846);
nor U4524 (N_4524,N_4064,N_3903);
and U4525 (N_4525,N_3791,N_4080);
or U4526 (N_4526,N_4097,N_4174);
xor U4527 (N_4527,N_3780,N_3843);
and U4528 (N_4528,N_3986,N_4331);
nor U4529 (N_4529,N_4060,N_3769);
or U4530 (N_4530,N_4079,N_4121);
and U4531 (N_4531,N_4303,N_3794);
nand U4532 (N_4532,N_4258,N_4193);
nor U4533 (N_4533,N_4061,N_3856);
or U4534 (N_4534,N_3754,N_3943);
or U4535 (N_4535,N_4135,N_4140);
nand U4536 (N_4536,N_4032,N_4276);
nand U4537 (N_4537,N_3770,N_4191);
nand U4538 (N_4538,N_3947,N_4249);
nor U4539 (N_4539,N_4073,N_3789);
and U4540 (N_4540,N_3908,N_4004);
nor U4541 (N_4541,N_4372,N_3920);
and U4542 (N_4542,N_4145,N_4180);
and U4543 (N_4543,N_4126,N_4298);
and U4544 (N_4544,N_3834,N_3919);
nor U4545 (N_4545,N_4183,N_4175);
xor U4546 (N_4546,N_4153,N_3887);
nor U4547 (N_4547,N_4159,N_4342);
or U4548 (N_4548,N_4008,N_4150);
or U4549 (N_4549,N_3800,N_4048);
xnor U4550 (N_4550,N_4067,N_4076);
or U4551 (N_4551,N_3859,N_4068);
or U4552 (N_4552,N_4086,N_4014);
xor U4553 (N_4553,N_4100,N_4216);
xor U4554 (N_4554,N_4286,N_3924);
xnor U4555 (N_4555,N_4259,N_4203);
nor U4556 (N_4556,N_4292,N_4056);
xor U4557 (N_4557,N_3914,N_3902);
nand U4558 (N_4558,N_4305,N_4030);
or U4559 (N_4559,N_4013,N_3823);
nand U4560 (N_4560,N_3854,N_4179);
and U4561 (N_4561,N_3901,N_4029);
and U4562 (N_4562,N_4206,N_4349);
or U4563 (N_4563,N_4360,N_3785);
xnor U4564 (N_4564,N_3895,N_4314);
xnor U4565 (N_4565,N_3898,N_4077);
or U4566 (N_4566,N_4256,N_4041);
nor U4567 (N_4567,N_3766,N_4095);
xor U4568 (N_4568,N_4266,N_4019);
and U4569 (N_4569,N_4170,N_3815);
nand U4570 (N_4570,N_4350,N_4248);
or U4571 (N_4571,N_4371,N_3833);
and U4572 (N_4572,N_4137,N_3817);
nor U4573 (N_4573,N_3883,N_3968);
and U4574 (N_4574,N_4366,N_3963);
or U4575 (N_4575,N_4365,N_4205);
nand U4576 (N_4576,N_4315,N_4294);
nand U4577 (N_4577,N_4221,N_4167);
nand U4578 (N_4578,N_3989,N_4088);
or U4579 (N_4579,N_3974,N_4229);
and U4580 (N_4580,N_3917,N_4185);
and U4581 (N_4581,N_3803,N_3767);
or U4582 (N_4582,N_4194,N_4247);
xnor U4583 (N_4583,N_4151,N_4296);
nand U4584 (N_4584,N_3942,N_3881);
nand U4585 (N_4585,N_3760,N_4334);
and U4586 (N_4586,N_3784,N_4109);
or U4587 (N_4587,N_3773,N_3891);
xnor U4588 (N_4588,N_4231,N_3913);
nor U4589 (N_4589,N_3872,N_4156);
or U4590 (N_4590,N_4223,N_4309);
and U4591 (N_4591,N_4272,N_4199);
nor U4592 (N_4592,N_3991,N_3976);
and U4593 (N_4593,N_4178,N_3964);
and U4594 (N_4594,N_3940,N_4105);
xor U4595 (N_4595,N_4012,N_4295);
and U4596 (N_4596,N_3820,N_4063);
nor U4597 (N_4597,N_3829,N_4050);
xnor U4598 (N_4598,N_3790,N_3775);
and U4599 (N_4599,N_4212,N_4104);
nor U4600 (N_4600,N_3912,N_4127);
and U4601 (N_4601,N_3812,N_4188);
nor U4602 (N_4602,N_3946,N_4103);
nand U4603 (N_4603,N_3781,N_3936);
nor U4604 (N_4604,N_4005,N_4092);
or U4605 (N_4605,N_4164,N_4369);
or U4606 (N_4606,N_4368,N_3959);
and U4607 (N_4607,N_4241,N_3763);
and U4608 (N_4608,N_4010,N_4018);
xnor U4609 (N_4609,N_3953,N_3830);
and U4610 (N_4610,N_4312,N_4149);
nor U4611 (N_4611,N_3816,N_3893);
nand U4612 (N_4612,N_3984,N_4281);
or U4613 (N_4613,N_4333,N_4356);
and U4614 (N_4614,N_4240,N_4147);
nand U4615 (N_4615,N_4039,N_3798);
nor U4616 (N_4616,N_3811,N_4176);
nor U4617 (N_4617,N_3855,N_4224);
or U4618 (N_4618,N_3850,N_4072);
nor U4619 (N_4619,N_3889,N_4011);
nand U4620 (N_4620,N_4268,N_3824);
xor U4621 (N_4621,N_3929,N_4186);
and U4622 (N_4622,N_4197,N_4017);
or U4623 (N_4623,N_4114,N_4373);
or U4624 (N_4624,N_4038,N_3884);
nor U4625 (N_4625,N_3849,N_4036);
or U4626 (N_4626,N_3836,N_3874);
or U4627 (N_4627,N_4190,N_3900);
or U4628 (N_4628,N_4337,N_4112);
xnor U4629 (N_4629,N_3950,N_4283);
nand U4630 (N_4630,N_3870,N_4214);
nor U4631 (N_4631,N_4113,N_4355);
nand U4632 (N_4632,N_4037,N_4299);
and U4633 (N_4633,N_3759,N_4324);
nor U4634 (N_4634,N_3987,N_4002);
nor U4635 (N_4635,N_3752,N_4051);
nand U4636 (N_4636,N_3904,N_4233);
nor U4637 (N_4637,N_4328,N_4148);
or U4638 (N_4638,N_4192,N_4313);
or U4639 (N_4639,N_4195,N_3888);
or U4640 (N_4640,N_4213,N_4182);
or U4641 (N_4641,N_3973,N_3853);
nor U4642 (N_4642,N_4279,N_3990);
xor U4643 (N_4643,N_3921,N_4007);
xor U4644 (N_4644,N_4341,N_4244);
nor U4645 (N_4645,N_4271,N_3821);
xor U4646 (N_4646,N_3778,N_4107);
and U4647 (N_4647,N_3796,N_3805);
or U4648 (N_4648,N_4353,N_3860);
nand U4649 (N_4649,N_4042,N_3988);
or U4650 (N_4650,N_4035,N_3979);
xnor U4651 (N_4651,N_3842,N_4289);
nor U4652 (N_4652,N_4123,N_3980);
or U4653 (N_4653,N_4125,N_3894);
nand U4654 (N_4654,N_3967,N_4320);
nor U4655 (N_4655,N_4325,N_4277);
xor U4656 (N_4656,N_4280,N_4134);
or U4657 (N_4657,N_3935,N_4310);
or U4658 (N_4658,N_4200,N_4132);
nand U4659 (N_4659,N_4054,N_4110);
nor U4660 (N_4660,N_3792,N_4358);
xnor U4661 (N_4661,N_3961,N_3972);
nor U4662 (N_4662,N_4230,N_3944);
xor U4663 (N_4663,N_3877,N_4057);
and U4664 (N_4664,N_4129,N_4264);
nand U4665 (N_4665,N_4359,N_3995);
xor U4666 (N_4666,N_4066,N_3931);
and U4667 (N_4667,N_3845,N_4087);
nor U4668 (N_4668,N_3837,N_4144);
or U4669 (N_4669,N_4370,N_3930);
and U4670 (N_4670,N_3905,N_3793);
nand U4671 (N_4671,N_3786,N_4293);
or U4672 (N_4672,N_3852,N_3802);
or U4673 (N_4673,N_4225,N_3807);
and U4674 (N_4674,N_4108,N_4161);
or U4675 (N_4675,N_4136,N_4094);
or U4676 (N_4676,N_4120,N_3962);
or U4677 (N_4677,N_4269,N_4169);
and U4678 (N_4678,N_4306,N_4020);
nor U4679 (N_4679,N_3783,N_4207);
or U4680 (N_4680,N_3949,N_3804);
xor U4681 (N_4681,N_4028,N_4338);
nand U4682 (N_4682,N_4189,N_3809);
nand U4683 (N_4683,N_4091,N_3899);
nor U4684 (N_4684,N_3958,N_4288);
and U4685 (N_4685,N_4282,N_4111);
xor U4686 (N_4686,N_4326,N_4311);
nor U4687 (N_4687,N_3774,N_4358);
xor U4688 (N_4688,N_3855,N_4110);
or U4689 (N_4689,N_4330,N_4325);
and U4690 (N_4690,N_4293,N_4183);
or U4691 (N_4691,N_4150,N_4348);
or U4692 (N_4692,N_4213,N_3804);
or U4693 (N_4693,N_4172,N_4302);
nor U4694 (N_4694,N_4062,N_3930);
xnor U4695 (N_4695,N_3895,N_4115);
and U4696 (N_4696,N_3945,N_4121);
nor U4697 (N_4697,N_4076,N_4352);
or U4698 (N_4698,N_3962,N_4179);
nand U4699 (N_4699,N_4354,N_3853);
or U4700 (N_4700,N_4372,N_4076);
and U4701 (N_4701,N_4262,N_3857);
nand U4702 (N_4702,N_4000,N_4012);
xnor U4703 (N_4703,N_4273,N_4027);
nand U4704 (N_4704,N_3756,N_4293);
and U4705 (N_4705,N_3952,N_4059);
xnor U4706 (N_4706,N_4041,N_4356);
or U4707 (N_4707,N_4202,N_3850);
xnor U4708 (N_4708,N_3782,N_4207);
nor U4709 (N_4709,N_4162,N_4364);
nand U4710 (N_4710,N_4210,N_4293);
xor U4711 (N_4711,N_4018,N_4201);
and U4712 (N_4712,N_4241,N_4141);
xor U4713 (N_4713,N_4177,N_4353);
and U4714 (N_4714,N_3829,N_3801);
and U4715 (N_4715,N_3994,N_4345);
or U4716 (N_4716,N_3899,N_4269);
xnor U4717 (N_4717,N_4191,N_4110);
and U4718 (N_4718,N_4043,N_4104);
nor U4719 (N_4719,N_4163,N_3807);
nand U4720 (N_4720,N_4136,N_3768);
or U4721 (N_4721,N_4236,N_4292);
and U4722 (N_4722,N_4025,N_3820);
or U4723 (N_4723,N_4283,N_4181);
xor U4724 (N_4724,N_4181,N_3844);
nor U4725 (N_4725,N_4271,N_4369);
nand U4726 (N_4726,N_3777,N_3896);
nand U4727 (N_4727,N_3771,N_3926);
nor U4728 (N_4728,N_4176,N_3943);
nand U4729 (N_4729,N_3799,N_4333);
nand U4730 (N_4730,N_4139,N_4051);
or U4731 (N_4731,N_3874,N_3781);
xnor U4732 (N_4732,N_4348,N_3791);
and U4733 (N_4733,N_3815,N_4301);
nor U4734 (N_4734,N_4128,N_4287);
and U4735 (N_4735,N_3851,N_4158);
or U4736 (N_4736,N_4275,N_4069);
nor U4737 (N_4737,N_4146,N_4340);
and U4738 (N_4738,N_3821,N_4333);
nor U4739 (N_4739,N_4196,N_4254);
or U4740 (N_4740,N_4212,N_4096);
xor U4741 (N_4741,N_3836,N_4333);
or U4742 (N_4742,N_3880,N_3914);
nand U4743 (N_4743,N_4299,N_4202);
nand U4744 (N_4744,N_3929,N_4334);
and U4745 (N_4745,N_4233,N_4354);
nor U4746 (N_4746,N_3926,N_3891);
and U4747 (N_4747,N_4148,N_4192);
nand U4748 (N_4748,N_4079,N_3768);
and U4749 (N_4749,N_3767,N_4186);
nor U4750 (N_4750,N_3889,N_4143);
or U4751 (N_4751,N_3895,N_4156);
nand U4752 (N_4752,N_4130,N_3918);
and U4753 (N_4753,N_4231,N_4108);
nor U4754 (N_4754,N_3860,N_3903);
xnor U4755 (N_4755,N_4053,N_4149);
nand U4756 (N_4756,N_4046,N_4111);
or U4757 (N_4757,N_4203,N_3995);
xnor U4758 (N_4758,N_3911,N_4234);
and U4759 (N_4759,N_3957,N_4190);
xor U4760 (N_4760,N_3788,N_3767);
or U4761 (N_4761,N_4031,N_4289);
nand U4762 (N_4762,N_3831,N_4002);
nand U4763 (N_4763,N_4265,N_4153);
nor U4764 (N_4764,N_4239,N_4039);
nor U4765 (N_4765,N_4100,N_4323);
xor U4766 (N_4766,N_4035,N_3977);
or U4767 (N_4767,N_4133,N_4315);
and U4768 (N_4768,N_4173,N_4154);
and U4769 (N_4769,N_4173,N_3946);
xnor U4770 (N_4770,N_3796,N_4215);
and U4771 (N_4771,N_4020,N_4266);
or U4772 (N_4772,N_3864,N_4016);
nand U4773 (N_4773,N_3755,N_3914);
xor U4774 (N_4774,N_4107,N_3971);
nor U4775 (N_4775,N_3901,N_3765);
xor U4776 (N_4776,N_4192,N_4297);
or U4777 (N_4777,N_3923,N_3905);
nor U4778 (N_4778,N_4185,N_4188);
nand U4779 (N_4779,N_3958,N_4272);
xnor U4780 (N_4780,N_4249,N_4078);
nand U4781 (N_4781,N_4201,N_4202);
nand U4782 (N_4782,N_4367,N_3835);
nand U4783 (N_4783,N_4047,N_4259);
nand U4784 (N_4784,N_4266,N_3837);
and U4785 (N_4785,N_4092,N_3798);
nand U4786 (N_4786,N_4201,N_3855);
nor U4787 (N_4787,N_3800,N_4139);
xor U4788 (N_4788,N_4151,N_4099);
xnor U4789 (N_4789,N_3973,N_3941);
nor U4790 (N_4790,N_3756,N_3856);
nand U4791 (N_4791,N_4078,N_4343);
xnor U4792 (N_4792,N_3986,N_4281);
or U4793 (N_4793,N_4255,N_3809);
and U4794 (N_4794,N_4204,N_3901);
or U4795 (N_4795,N_4353,N_4316);
xnor U4796 (N_4796,N_3974,N_4300);
or U4797 (N_4797,N_4143,N_3981);
nor U4798 (N_4798,N_4311,N_3911);
nor U4799 (N_4799,N_3980,N_4077);
or U4800 (N_4800,N_4317,N_3892);
nand U4801 (N_4801,N_4224,N_4294);
xor U4802 (N_4802,N_3797,N_4374);
nor U4803 (N_4803,N_4102,N_4243);
nand U4804 (N_4804,N_4260,N_4118);
xor U4805 (N_4805,N_4188,N_3896);
or U4806 (N_4806,N_3999,N_4167);
nor U4807 (N_4807,N_3781,N_4273);
nor U4808 (N_4808,N_4104,N_3789);
nor U4809 (N_4809,N_4143,N_3948);
and U4810 (N_4810,N_4304,N_4066);
xor U4811 (N_4811,N_4021,N_4108);
and U4812 (N_4812,N_4126,N_3826);
and U4813 (N_4813,N_4362,N_3824);
nor U4814 (N_4814,N_3953,N_4101);
or U4815 (N_4815,N_3997,N_4052);
xnor U4816 (N_4816,N_4228,N_4019);
nand U4817 (N_4817,N_4133,N_4268);
xnor U4818 (N_4818,N_3833,N_3945);
and U4819 (N_4819,N_3935,N_4165);
xnor U4820 (N_4820,N_4315,N_4208);
xor U4821 (N_4821,N_3859,N_3941);
xnor U4822 (N_4822,N_3969,N_4072);
xor U4823 (N_4823,N_3885,N_3776);
and U4824 (N_4824,N_4259,N_3916);
or U4825 (N_4825,N_4327,N_3914);
xor U4826 (N_4826,N_4257,N_4245);
nor U4827 (N_4827,N_4334,N_4147);
nand U4828 (N_4828,N_3965,N_4356);
nor U4829 (N_4829,N_4121,N_4333);
xnor U4830 (N_4830,N_3973,N_4256);
nand U4831 (N_4831,N_4006,N_4133);
xor U4832 (N_4832,N_3805,N_3972);
or U4833 (N_4833,N_3954,N_3989);
xor U4834 (N_4834,N_4084,N_4001);
and U4835 (N_4835,N_4227,N_4186);
nand U4836 (N_4836,N_4291,N_3982);
or U4837 (N_4837,N_3913,N_4084);
or U4838 (N_4838,N_4244,N_4188);
or U4839 (N_4839,N_4261,N_3915);
xor U4840 (N_4840,N_4150,N_3858);
and U4841 (N_4841,N_3905,N_4026);
nor U4842 (N_4842,N_4174,N_4306);
nand U4843 (N_4843,N_4374,N_3987);
or U4844 (N_4844,N_3790,N_4234);
nor U4845 (N_4845,N_4308,N_3908);
xnor U4846 (N_4846,N_4075,N_4259);
xnor U4847 (N_4847,N_3833,N_4233);
and U4848 (N_4848,N_4021,N_4317);
and U4849 (N_4849,N_4333,N_4359);
xnor U4850 (N_4850,N_3907,N_4206);
nand U4851 (N_4851,N_4301,N_4032);
nand U4852 (N_4852,N_4152,N_4187);
or U4853 (N_4853,N_3757,N_3810);
or U4854 (N_4854,N_4263,N_4373);
and U4855 (N_4855,N_3983,N_4194);
or U4856 (N_4856,N_3766,N_3781);
nor U4857 (N_4857,N_3787,N_4333);
or U4858 (N_4858,N_4144,N_3980);
xnor U4859 (N_4859,N_3933,N_4301);
and U4860 (N_4860,N_4313,N_3808);
and U4861 (N_4861,N_4307,N_4086);
xnor U4862 (N_4862,N_4371,N_4075);
and U4863 (N_4863,N_4032,N_4124);
nor U4864 (N_4864,N_3755,N_4156);
nand U4865 (N_4865,N_3871,N_4349);
nand U4866 (N_4866,N_4004,N_3887);
xor U4867 (N_4867,N_4101,N_3924);
and U4868 (N_4868,N_4259,N_3836);
nand U4869 (N_4869,N_4285,N_4221);
and U4870 (N_4870,N_3804,N_3951);
or U4871 (N_4871,N_3916,N_3796);
nor U4872 (N_4872,N_3921,N_4093);
xnor U4873 (N_4873,N_4244,N_3829);
nor U4874 (N_4874,N_4056,N_3968);
nor U4875 (N_4875,N_3954,N_3933);
and U4876 (N_4876,N_4183,N_4085);
xor U4877 (N_4877,N_4343,N_4001);
nand U4878 (N_4878,N_3824,N_3842);
nand U4879 (N_4879,N_3812,N_3908);
nor U4880 (N_4880,N_4036,N_4118);
xor U4881 (N_4881,N_4263,N_4225);
and U4882 (N_4882,N_4007,N_4049);
and U4883 (N_4883,N_4024,N_3959);
nand U4884 (N_4884,N_3915,N_3815);
nand U4885 (N_4885,N_4179,N_4007);
or U4886 (N_4886,N_3782,N_3920);
xor U4887 (N_4887,N_3900,N_4012);
or U4888 (N_4888,N_4350,N_4341);
or U4889 (N_4889,N_3786,N_3868);
or U4890 (N_4890,N_4083,N_4323);
nand U4891 (N_4891,N_3834,N_4334);
nand U4892 (N_4892,N_3779,N_4315);
xor U4893 (N_4893,N_3756,N_4109);
or U4894 (N_4894,N_3884,N_4101);
or U4895 (N_4895,N_4091,N_3896);
or U4896 (N_4896,N_4005,N_3989);
nand U4897 (N_4897,N_4181,N_3778);
nand U4898 (N_4898,N_3955,N_4046);
nor U4899 (N_4899,N_4288,N_4332);
xor U4900 (N_4900,N_3873,N_4269);
and U4901 (N_4901,N_4065,N_4354);
nor U4902 (N_4902,N_4351,N_3996);
nor U4903 (N_4903,N_4098,N_4056);
or U4904 (N_4904,N_4052,N_3909);
nand U4905 (N_4905,N_3896,N_3904);
xnor U4906 (N_4906,N_3779,N_4352);
nand U4907 (N_4907,N_4053,N_3930);
or U4908 (N_4908,N_4215,N_4264);
nand U4909 (N_4909,N_4310,N_4072);
xnor U4910 (N_4910,N_3969,N_4265);
or U4911 (N_4911,N_4174,N_3874);
or U4912 (N_4912,N_3917,N_4290);
nand U4913 (N_4913,N_4043,N_4029);
nand U4914 (N_4914,N_3976,N_3778);
nor U4915 (N_4915,N_4370,N_4127);
or U4916 (N_4916,N_4070,N_3914);
nor U4917 (N_4917,N_3939,N_3834);
or U4918 (N_4918,N_3906,N_4206);
xnor U4919 (N_4919,N_4290,N_3863);
nand U4920 (N_4920,N_4151,N_4304);
and U4921 (N_4921,N_3978,N_4043);
nor U4922 (N_4922,N_3776,N_3904);
xnor U4923 (N_4923,N_3763,N_4350);
nand U4924 (N_4924,N_3771,N_3893);
nor U4925 (N_4925,N_4274,N_4080);
or U4926 (N_4926,N_3939,N_4234);
or U4927 (N_4927,N_3975,N_3777);
and U4928 (N_4928,N_3978,N_3990);
nand U4929 (N_4929,N_3763,N_4349);
and U4930 (N_4930,N_4286,N_4290);
nor U4931 (N_4931,N_4186,N_3913);
or U4932 (N_4932,N_4145,N_3781);
xor U4933 (N_4933,N_4159,N_4270);
nand U4934 (N_4934,N_4113,N_3907);
nand U4935 (N_4935,N_3998,N_4360);
nor U4936 (N_4936,N_3874,N_3820);
xnor U4937 (N_4937,N_3831,N_3990);
or U4938 (N_4938,N_4181,N_4221);
or U4939 (N_4939,N_3774,N_4323);
xor U4940 (N_4940,N_4134,N_3966);
xor U4941 (N_4941,N_4027,N_4036);
nor U4942 (N_4942,N_4132,N_4119);
xor U4943 (N_4943,N_3884,N_3810);
and U4944 (N_4944,N_3774,N_4066);
nand U4945 (N_4945,N_4089,N_4283);
nor U4946 (N_4946,N_4051,N_3828);
or U4947 (N_4947,N_3868,N_4023);
nand U4948 (N_4948,N_4185,N_4373);
nor U4949 (N_4949,N_4011,N_4224);
xnor U4950 (N_4950,N_3966,N_3905);
nand U4951 (N_4951,N_3920,N_4022);
xnor U4952 (N_4952,N_4009,N_3891);
nor U4953 (N_4953,N_3971,N_3789);
nor U4954 (N_4954,N_4167,N_3918);
or U4955 (N_4955,N_3984,N_4257);
nand U4956 (N_4956,N_3944,N_4297);
xnor U4957 (N_4957,N_4047,N_4163);
xor U4958 (N_4958,N_4151,N_3791);
xor U4959 (N_4959,N_4157,N_3811);
nand U4960 (N_4960,N_4360,N_3800);
nor U4961 (N_4961,N_3893,N_4042);
and U4962 (N_4962,N_3906,N_4007);
nor U4963 (N_4963,N_4205,N_4190);
or U4964 (N_4964,N_3960,N_4161);
nand U4965 (N_4965,N_4273,N_4363);
nor U4966 (N_4966,N_4105,N_4347);
or U4967 (N_4967,N_4265,N_4239);
or U4968 (N_4968,N_4067,N_4183);
and U4969 (N_4969,N_3980,N_4356);
xor U4970 (N_4970,N_4279,N_4288);
nand U4971 (N_4971,N_4078,N_3930);
nand U4972 (N_4972,N_3935,N_3789);
nor U4973 (N_4973,N_3922,N_4335);
nand U4974 (N_4974,N_3962,N_4273);
nor U4975 (N_4975,N_4180,N_3993);
or U4976 (N_4976,N_4129,N_4150);
and U4977 (N_4977,N_4151,N_3789);
nand U4978 (N_4978,N_3958,N_4344);
or U4979 (N_4979,N_4245,N_4266);
and U4980 (N_4980,N_4155,N_4119);
nor U4981 (N_4981,N_3803,N_4221);
or U4982 (N_4982,N_4332,N_4365);
nor U4983 (N_4983,N_4297,N_4236);
nand U4984 (N_4984,N_3803,N_3974);
nand U4985 (N_4985,N_3992,N_4070);
nand U4986 (N_4986,N_4056,N_4285);
xor U4987 (N_4987,N_4019,N_3947);
nand U4988 (N_4988,N_4055,N_4373);
or U4989 (N_4989,N_4242,N_4116);
and U4990 (N_4990,N_3969,N_4299);
nand U4991 (N_4991,N_3983,N_3754);
nand U4992 (N_4992,N_4295,N_3914);
or U4993 (N_4993,N_3993,N_4349);
nand U4994 (N_4994,N_3943,N_3824);
nand U4995 (N_4995,N_4104,N_3930);
nand U4996 (N_4996,N_3975,N_4281);
nor U4997 (N_4997,N_3889,N_3773);
or U4998 (N_4998,N_3750,N_4017);
or U4999 (N_4999,N_3882,N_4355);
and U5000 (N_5000,N_4848,N_4853);
or U5001 (N_5001,N_4912,N_4390);
or U5002 (N_5002,N_4464,N_4667);
xnor U5003 (N_5003,N_4773,N_4463);
nor U5004 (N_5004,N_4566,N_4849);
or U5005 (N_5005,N_4658,N_4775);
xor U5006 (N_5006,N_4488,N_4842);
or U5007 (N_5007,N_4649,N_4602);
nor U5008 (N_5008,N_4962,N_4731);
nor U5009 (N_5009,N_4690,N_4948);
nand U5010 (N_5010,N_4445,N_4578);
and U5011 (N_5011,N_4951,N_4722);
or U5012 (N_5012,N_4659,N_4622);
and U5013 (N_5013,N_4983,N_4791);
and U5014 (N_5014,N_4507,N_4890);
or U5015 (N_5015,N_4556,N_4902);
xnor U5016 (N_5016,N_4819,N_4618);
and U5017 (N_5017,N_4917,N_4614);
or U5018 (N_5018,N_4748,N_4531);
nand U5019 (N_5019,N_4715,N_4854);
nor U5020 (N_5020,N_4899,N_4650);
xor U5021 (N_5021,N_4898,N_4877);
nand U5022 (N_5022,N_4936,N_4817);
nor U5023 (N_5023,N_4502,N_4975);
or U5024 (N_5024,N_4519,N_4694);
nand U5025 (N_5025,N_4993,N_4816);
xor U5026 (N_5026,N_4830,N_4453);
and U5027 (N_5027,N_4674,N_4527);
xnor U5028 (N_5028,N_4812,N_4794);
nand U5029 (N_5029,N_4553,N_4423);
nor U5030 (N_5030,N_4668,N_4711);
xor U5031 (N_5031,N_4868,N_4508);
nor U5032 (N_5032,N_4472,N_4823);
and U5033 (N_5033,N_4678,N_4414);
nand U5034 (N_5034,N_4561,N_4687);
nor U5035 (N_5035,N_4485,N_4834);
nand U5036 (N_5036,N_4953,N_4500);
and U5037 (N_5037,N_4511,N_4473);
or U5038 (N_5038,N_4451,N_4883);
xor U5039 (N_5039,N_4944,N_4610);
or U5040 (N_5040,N_4872,N_4763);
nor U5041 (N_5041,N_4987,N_4856);
and U5042 (N_5042,N_4406,N_4394);
nor U5043 (N_5043,N_4478,N_4870);
nand U5044 (N_5044,N_4528,N_4664);
and U5045 (N_5045,N_4728,N_4847);
or U5046 (N_5046,N_4846,N_4892);
and U5047 (N_5047,N_4805,N_4539);
and U5048 (N_5048,N_4956,N_4484);
and U5049 (N_5049,N_4720,N_4851);
and U5050 (N_5050,N_4729,N_4441);
xnor U5051 (N_5051,N_4879,N_4810);
nor U5052 (N_5052,N_4671,N_4928);
or U5053 (N_5053,N_4882,N_4557);
or U5054 (N_5054,N_4613,N_4867);
xnor U5055 (N_5055,N_4803,N_4981);
nor U5056 (N_5056,N_4384,N_4798);
nor U5057 (N_5057,N_4437,N_4654);
nand U5058 (N_5058,N_4754,N_4638);
or U5059 (N_5059,N_4918,N_4996);
and U5060 (N_5060,N_4696,N_4818);
nor U5061 (N_5061,N_4706,N_4564);
or U5062 (N_5062,N_4838,N_4376);
or U5063 (N_5063,N_4946,N_4621);
nor U5064 (N_5064,N_4583,N_4767);
and U5065 (N_5065,N_4685,N_4637);
nor U5066 (N_5066,N_4560,N_4477);
xor U5067 (N_5067,N_4426,N_4777);
or U5068 (N_5068,N_4814,N_4516);
and U5069 (N_5069,N_4859,N_4753);
nand U5070 (N_5070,N_4875,N_4701);
xnor U5071 (N_5071,N_4547,N_4465);
nand U5072 (N_5072,N_4629,N_4417);
nand U5073 (N_5073,N_4934,N_4733);
xor U5074 (N_5074,N_4703,N_4525);
or U5075 (N_5075,N_4660,N_4933);
and U5076 (N_5076,N_4985,N_4448);
xnor U5077 (N_5077,N_4433,N_4494);
or U5078 (N_5078,N_4765,N_4693);
nor U5079 (N_5079,N_4392,N_4549);
nor U5080 (N_5080,N_4474,N_4863);
nand U5081 (N_5081,N_4970,N_4761);
nor U5082 (N_5082,N_4862,N_4735);
xor U5083 (N_5083,N_4626,N_4976);
nor U5084 (N_5084,N_4977,N_4513);
nor U5085 (N_5085,N_4570,N_4554);
nor U5086 (N_5086,N_4772,N_4861);
nand U5087 (N_5087,N_4904,N_4876);
or U5088 (N_5088,N_4689,N_4866);
nand U5089 (N_5089,N_4957,N_4375);
or U5090 (N_5090,N_4852,N_4959);
and U5091 (N_5091,N_4497,N_4895);
nand U5092 (N_5092,N_4466,N_4776);
or U5093 (N_5093,N_4579,N_4921);
xor U5094 (N_5094,N_4691,N_4808);
or U5095 (N_5095,N_4881,N_4692);
nand U5096 (N_5096,N_4961,N_4672);
or U5097 (N_5097,N_4480,N_4438);
and U5098 (N_5098,N_4670,N_4782);
or U5099 (N_5099,N_4718,N_4546);
or U5100 (N_5100,N_4771,N_4572);
and U5101 (N_5101,N_4815,N_4865);
nor U5102 (N_5102,N_4841,N_4617);
or U5103 (N_5103,N_4491,N_4990);
nand U5104 (N_5104,N_4790,N_4945);
xor U5105 (N_5105,N_4585,N_4683);
nor U5106 (N_5106,N_4586,N_4590);
nand U5107 (N_5107,N_4927,N_4398);
or U5108 (N_5108,N_4829,N_4404);
nor U5109 (N_5109,N_4379,N_4475);
nor U5110 (N_5110,N_4608,N_4955);
xor U5111 (N_5111,N_4545,N_4575);
and U5112 (N_5112,N_4732,N_4965);
xnor U5113 (N_5113,N_4991,N_4529);
xnor U5114 (N_5114,N_4385,N_4897);
nand U5115 (N_5115,N_4709,N_4986);
nor U5116 (N_5116,N_4434,N_4643);
nand U5117 (N_5117,N_4843,N_4938);
nand U5118 (N_5118,N_4869,N_4537);
or U5119 (N_5119,N_4653,N_4391);
and U5120 (N_5120,N_4682,N_4960);
xor U5121 (N_5121,N_4966,N_4551);
nand U5122 (N_5122,N_4542,N_4787);
xor U5123 (N_5123,N_4874,N_4383);
and U5124 (N_5124,N_4901,N_4958);
nor U5125 (N_5125,N_4992,N_4721);
and U5126 (N_5126,N_4630,N_4697);
and U5127 (N_5127,N_4850,N_4871);
or U5128 (N_5128,N_4745,N_4532);
nand U5129 (N_5129,N_4884,N_4781);
or U5130 (N_5130,N_4467,N_4736);
xnor U5131 (N_5131,N_4571,N_4793);
and U5132 (N_5132,N_4710,N_4459);
and U5133 (N_5133,N_4967,N_4786);
xnor U5134 (N_5134,N_4624,N_4909);
xnor U5135 (N_5135,N_4700,N_4496);
and U5136 (N_5136,N_4483,N_4926);
or U5137 (N_5137,N_4616,N_4601);
xnor U5138 (N_5138,N_4964,N_4755);
nand U5139 (N_5139,N_4569,N_4397);
xor U5140 (N_5140,N_4481,N_4886);
nand U5141 (N_5141,N_4625,N_4717);
and U5142 (N_5142,N_4550,N_4646);
nand U5143 (N_5143,N_4925,N_4908);
nor U5144 (N_5144,N_4386,N_4768);
and U5145 (N_5145,N_4752,N_4963);
or U5146 (N_5146,N_4597,N_4400);
xnor U5147 (N_5147,N_4971,N_4792);
xor U5148 (N_5148,N_4778,N_4587);
and U5149 (N_5149,N_4673,N_4639);
xor U5150 (N_5150,N_4840,N_4825);
and U5151 (N_5151,N_4517,N_4640);
nor U5152 (N_5152,N_4422,N_4647);
nor U5153 (N_5153,N_4974,N_4835);
and U5154 (N_5154,N_4424,N_4446);
and U5155 (N_5155,N_4929,N_4656);
or U5156 (N_5156,N_4439,N_4450);
and U5157 (N_5157,N_4797,N_4739);
xor U5158 (N_5158,N_4760,N_4452);
nor U5159 (N_5159,N_4666,N_4455);
or U5160 (N_5160,N_4893,N_4913);
or U5161 (N_5161,N_4609,N_4563);
xnor U5162 (N_5162,N_4980,N_4381);
xor U5163 (N_5163,N_4695,N_4430);
or U5164 (N_5164,N_4801,N_4503);
and U5165 (N_5165,N_4506,N_4774);
or U5166 (N_5166,N_4836,N_4675);
nand U5167 (N_5167,N_4458,N_4395);
nand U5168 (N_5168,N_4628,N_4454);
and U5169 (N_5169,N_4416,N_4995);
nor U5170 (N_5170,N_4600,N_4538);
nor U5171 (N_5171,N_4512,N_4943);
or U5172 (N_5172,N_4495,N_4581);
nand U5173 (N_5173,N_4418,N_4584);
or U5174 (N_5174,N_4930,N_4443);
and U5175 (N_5175,N_4730,N_4950);
xnor U5176 (N_5176,N_4833,N_4839);
nor U5177 (N_5177,N_4663,N_4620);
or U5178 (N_5178,N_4482,N_4419);
nor U5179 (N_5179,N_4651,N_4704);
xnor U5180 (N_5180,N_4820,N_4489);
and U5181 (N_5181,N_4442,N_4914);
and U5182 (N_5182,N_4758,N_4521);
or U5183 (N_5183,N_4744,N_4509);
xnor U5184 (N_5184,N_4716,N_4574);
nand U5185 (N_5185,N_4724,N_4501);
and U5186 (N_5186,N_4631,N_4471);
or U5187 (N_5187,N_4410,N_4747);
nand U5188 (N_5188,N_4676,N_4727);
or U5189 (N_5189,N_4492,N_4734);
nor U5190 (N_5190,N_4799,N_4526);
nor U5191 (N_5191,N_4611,N_4447);
nand U5192 (N_5192,N_4800,N_4552);
and U5193 (N_5193,N_4903,N_4952);
nand U5194 (N_5194,N_4470,N_4669);
and U5195 (N_5195,N_4636,N_4415);
and U5196 (N_5196,N_4476,N_4811);
nand U5197 (N_5197,N_4920,N_4873);
and U5198 (N_5198,N_4807,N_4662);
and U5199 (N_5199,N_4947,N_4510);
xor U5200 (N_5200,N_4919,N_4708);
nor U5201 (N_5201,N_4606,N_4954);
or U5202 (N_5202,N_4702,N_4393);
or U5203 (N_5203,N_4746,N_4982);
or U5204 (N_5204,N_4707,N_4407);
nor U5205 (N_5205,N_4937,N_4589);
or U5206 (N_5206,N_4555,N_4887);
xnor U5207 (N_5207,N_4828,N_4940);
xnor U5208 (N_5208,N_4837,N_4741);
or U5209 (N_5209,N_4409,N_4699);
or U5210 (N_5210,N_4648,N_4738);
xor U5211 (N_5211,N_4607,N_4534);
or U5212 (N_5212,N_4661,N_4742);
and U5213 (N_5213,N_4523,N_4860);
or U5214 (N_5214,N_4988,N_4421);
xnor U5215 (N_5215,N_4380,N_4905);
and U5216 (N_5216,N_4594,N_4541);
xor U5217 (N_5217,N_4493,N_4845);
nand U5218 (N_5218,N_4764,N_4479);
nor U5219 (N_5219,N_4535,N_4922);
nand U5220 (N_5220,N_4428,N_4878);
xnor U5221 (N_5221,N_4759,N_4558);
and U5222 (N_5222,N_4827,N_4723);
or U5223 (N_5223,N_4998,N_4468);
and U5224 (N_5224,N_4499,N_4994);
and U5225 (N_5225,N_4677,N_4725);
and U5226 (N_5226,N_4377,N_4425);
nand U5227 (N_5227,N_4462,N_4619);
nand U5228 (N_5228,N_4411,N_4688);
or U5229 (N_5229,N_4968,N_4524);
and U5230 (N_5230,N_4824,N_4681);
nand U5231 (N_5231,N_4813,N_4796);
and U5232 (N_5232,N_4749,N_4916);
nor U5233 (N_5233,N_4931,N_4680);
nor U5234 (N_5234,N_4655,N_4858);
nand U5235 (N_5235,N_4632,N_4915);
and U5236 (N_5236,N_4864,N_4504);
nand U5237 (N_5237,N_4889,N_4740);
xnor U5238 (N_5238,N_4779,N_4456);
nand U5239 (N_5239,N_4888,N_4573);
nand U5240 (N_5240,N_4644,N_4568);
xnor U5241 (N_5241,N_4530,N_4487);
and U5242 (N_5242,N_4979,N_4972);
nand U5243 (N_5243,N_4429,N_4457);
and U5244 (N_5244,N_4461,N_4577);
nor U5245 (N_5245,N_4652,N_4596);
nand U5246 (N_5246,N_4378,N_4978);
nand U5247 (N_5247,N_4907,N_4855);
nor U5248 (N_5248,N_4408,N_4427);
or U5249 (N_5249,N_4548,N_4780);
nor U5250 (N_5250,N_4382,N_4770);
xnor U5251 (N_5251,N_4783,N_4420);
or U5252 (N_5252,N_4784,N_4633);
xor U5253 (N_5253,N_4844,N_4540);
nand U5254 (N_5254,N_4396,N_4891);
nor U5255 (N_5255,N_4440,N_4543);
or U5256 (N_5256,N_4603,N_4665);
nand U5257 (N_5257,N_4989,N_4822);
and U5258 (N_5258,N_4387,N_4941);
and U5259 (N_5259,N_4911,N_4460);
and U5260 (N_5260,N_4756,N_4949);
or U5261 (N_5261,N_4806,N_4591);
nand U5262 (N_5262,N_4490,N_4896);
or U5263 (N_5263,N_4785,N_4705);
xor U5264 (N_5264,N_4762,N_4412);
or U5265 (N_5265,N_4788,N_4562);
and U5266 (N_5266,N_4515,N_4469);
nand U5267 (N_5267,N_4932,N_4592);
nand U5268 (N_5268,N_4520,N_4795);
or U5269 (N_5269,N_4559,N_4580);
xnor U5270 (N_5270,N_4679,N_4743);
and U5271 (N_5271,N_4615,N_4627);
and U5272 (N_5272,N_4684,N_4885);
nand U5273 (N_5273,N_4498,N_4900);
xor U5274 (N_5274,N_4726,N_4831);
xor U5275 (N_5275,N_4536,N_4402);
xor U5276 (N_5276,N_4514,N_4604);
nand U5277 (N_5277,N_4449,N_4737);
and U5278 (N_5278,N_4894,N_4789);
or U5279 (N_5279,N_4595,N_4769);
and U5280 (N_5280,N_4802,N_4969);
nor U5281 (N_5281,N_4973,N_4388);
xor U5282 (N_5282,N_4605,N_4857);
or U5283 (N_5283,N_4750,N_4751);
and U5284 (N_5284,N_4999,N_4804);
xnor U5285 (N_5285,N_4576,N_4623);
or U5286 (N_5286,N_4598,N_4924);
xnor U5287 (N_5287,N_4880,N_4984);
nor U5288 (N_5288,N_4567,N_4939);
nor U5289 (N_5289,N_4935,N_4399);
nand U5290 (N_5290,N_4686,N_4588);
xor U5291 (N_5291,N_4657,N_4906);
nand U5292 (N_5292,N_4719,N_4444);
nor U5293 (N_5293,N_4436,N_4582);
nor U5294 (N_5294,N_4635,N_4544);
and U5295 (N_5295,N_4403,N_4809);
and U5296 (N_5296,N_4712,N_4713);
nor U5297 (N_5297,N_4593,N_4698);
and U5298 (N_5298,N_4486,N_4634);
nor U5299 (N_5299,N_4565,N_4923);
nor U5300 (N_5300,N_4641,N_4405);
or U5301 (N_5301,N_4389,N_4435);
and U5302 (N_5302,N_4642,N_4645);
nand U5303 (N_5303,N_4757,N_4505);
or U5304 (N_5304,N_4910,N_4714);
or U5305 (N_5305,N_4401,N_4832);
nor U5306 (N_5306,N_4518,N_4612);
nand U5307 (N_5307,N_4533,N_4766);
nor U5308 (N_5308,N_4942,N_4599);
nor U5309 (N_5309,N_4432,N_4431);
or U5310 (N_5310,N_4522,N_4997);
xnor U5311 (N_5311,N_4821,N_4413);
nand U5312 (N_5312,N_4826,N_4741);
xor U5313 (N_5313,N_4735,N_4920);
and U5314 (N_5314,N_4977,N_4930);
xnor U5315 (N_5315,N_4988,N_4750);
nand U5316 (N_5316,N_4756,N_4518);
xnor U5317 (N_5317,N_4786,N_4478);
nand U5318 (N_5318,N_4977,N_4485);
or U5319 (N_5319,N_4392,N_4667);
nor U5320 (N_5320,N_4680,N_4716);
or U5321 (N_5321,N_4979,N_4529);
and U5322 (N_5322,N_4478,N_4994);
or U5323 (N_5323,N_4933,N_4855);
and U5324 (N_5324,N_4680,N_4550);
xnor U5325 (N_5325,N_4452,N_4814);
nor U5326 (N_5326,N_4937,N_4704);
nor U5327 (N_5327,N_4584,N_4562);
or U5328 (N_5328,N_4834,N_4943);
xnor U5329 (N_5329,N_4768,N_4738);
or U5330 (N_5330,N_4769,N_4526);
nor U5331 (N_5331,N_4929,N_4914);
xnor U5332 (N_5332,N_4969,N_4950);
nand U5333 (N_5333,N_4693,N_4927);
nor U5334 (N_5334,N_4712,N_4680);
or U5335 (N_5335,N_4436,N_4494);
nand U5336 (N_5336,N_4486,N_4771);
xor U5337 (N_5337,N_4599,N_4490);
nand U5338 (N_5338,N_4616,N_4382);
or U5339 (N_5339,N_4552,N_4783);
and U5340 (N_5340,N_4534,N_4752);
or U5341 (N_5341,N_4482,N_4406);
and U5342 (N_5342,N_4523,N_4629);
and U5343 (N_5343,N_4577,N_4546);
and U5344 (N_5344,N_4695,N_4795);
nand U5345 (N_5345,N_4462,N_4448);
nand U5346 (N_5346,N_4458,N_4894);
xor U5347 (N_5347,N_4610,N_4793);
nand U5348 (N_5348,N_4618,N_4627);
nor U5349 (N_5349,N_4740,N_4426);
and U5350 (N_5350,N_4892,N_4611);
and U5351 (N_5351,N_4950,N_4967);
nor U5352 (N_5352,N_4759,N_4756);
nor U5353 (N_5353,N_4583,N_4620);
and U5354 (N_5354,N_4699,N_4970);
xor U5355 (N_5355,N_4946,N_4821);
xnor U5356 (N_5356,N_4705,N_4881);
nor U5357 (N_5357,N_4576,N_4377);
and U5358 (N_5358,N_4538,N_4657);
and U5359 (N_5359,N_4829,N_4738);
nor U5360 (N_5360,N_4672,N_4462);
and U5361 (N_5361,N_4843,N_4709);
nor U5362 (N_5362,N_4702,N_4783);
xnor U5363 (N_5363,N_4770,N_4527);
nand U5364 (N_5364,N_4829,N_4571);
xnor U5365 (N_5365,N_4482,N_4505);
nand U5366 (N_5366,N_4882,N_4623);
and U5367 (N_5367,N_4790,N_4986);
xnor U5368 (N_5368,N_4751,N_4534);
or U5369 (N_5369,N_4478,N_4522);
or U5370 (N_5370,N_4894,N_4390);
nor U5371 (N_5371,N_4395,N_4802);
nand U5372 (N_5372,N_4984,N_4596);
nand U5373 (N_5373,N_4457,N_4952);
and U5374 (N_5374,N_4456,N_4562);
xnor U5375 (N_5375,N_4621,N_4945);
nand U5376 (N_5376,N_4882,N_4583);
and U5377 (N_5377,N_4667,N_4918);
xnor U5378 (N_5378,N_4836,N_4889);
and U5379 (N_5379,N_4546,N_4696);
nor U5380 (N_5380,N_4480,N_4935);
xor U5381 (N_5381,N_4831,N_4586);
nand U5382 (N_5382,N_4492,N_4780);
or U5383 (N_5383,N_4872,N_4789);
nor U5384 (N_5384,N_4872,N_4449);
and U5385 (N_5385,N_4777,N_4460);
or U5386 (N_5386,N_4658,N_4533);
or U5387 (N_5387,N_4731,N_4387);
xnor U5388 (N_5388,N_4739,N_4844);
or U5389 (N_5389,N_4390,N_4864);
nand U5390 (N_5390,N_4786,N_4477);
xor U5391 (N_5391,N_4637,N_4448);
xor U5392 (N_5392,N_4859,N_4744);
or U5393 (N_5393,N_4977,N_4623);
nand U5394 (N_5394,N_4985,N_4678);
or U5395 (N_5395,N_4679,N_4878);
xnor U5396 (N_5396,N_4556,N_4901);
nor U5397 (N_5397,N_4636,N_4533);
or U5398 (N_5398,N_4920,N_4647);
and U5399 (N_5399,N_4441,N_4988);
and U5400 (N_5400,N_4612,N_4398);
nor U5401 (N_5401,N_4875,N_4924);
nor U5402 (N_5402,N_4979,N_4581);
or U5403 (N_5403,N_4927,N_4800);
xor U5404 (N_5404,N_4476,N_4787);
xnor U5405 (N_5405,N_4720,N_4968);
nor U5406 (N_5406,N_4922,N_4839);
nor U5407 (N_5407,N_4606,N_4815);
nand U5408 (N_5408,N_4835,N_4925);
xor U5409 (N_5409,N_4611,N_4379);
or U5410 (N_5410,N_4405,N_4451);
nor U5411 (N_5411,N_4376,N_4650);
and U5412 (N_5412,N_4958,N_4684);
xor U5413 (N_5413,N_4473,N_4727);
nor U5414 (N_5414,N_4534,N_4555);
nand U5415 (N_5415,N_4916,N_4759);
or U5416 (N_5416,N_4659,N_4941);
nand U5417 (N_5417,N_4401,N_4741);
nor U5418 (N_5418,N_4673,N_4378);
nand U5419 (N_5419,N_4795,N_4897);
and U5420 (N_5420,N_4511,N_4767);
or U5421 (N_5421,N_4782,N_4573);
or U5422 (N_5422,N_4421,N_4580);
xnor U5423 (N_5423,N_4522,N_4473);
and U5424 (N_5424,N_4559,N_4890);
or U5425 (N_5425,N_4859,N_4766);
or U5426 (N_5426,N_4792,N_4603);
nor U5427 (N_5427,N_4555,N_4661);
or U5428 (N_5428,N_4450,N_4841);
xnor U5429 (N_5429,N_4550,N_4918);
xnor U5430 (N_5430,N_4886,N_4874);
and U5431 (N_5431,N_4443,N_4711);
or U5432 (N_5432,N_4404,N_4492);
or U5433 (N_5433,N_4923,N_4891);
xnor U5434 (N_5434,N_4912,N_4515);
nand U5435 (N_5435,N_4812,N_4461);
nand U5436 (N_5436,N_4893,N_4480);
nor U5437 (N_5437,N_4995,N_4998);
xnor U5438 (N_5438,N_4956,N_4549);
and U5439 (N_5439,N_4467,N_4985);
nor U5440 (N_5440,N_4831,N_4815);
xnor U5441 (N_5441,N_4601,N_4639);
xor U5442 (N_5442,N_4736,N_4926);
or U5443 (N_5443,N_4540,N_4768);
xnor U5444 (N_5444,N_4650,N_4539);
or U5445 (N_5445,N_4490,N_4829);
and U5446 (N_5446,N_4810,N_4640);
nor U5447 (N_5447,N_4498,N_4399);
nand U5448 (N_5448,N_4744,N_4647);
and U5449 (N_5449,N_4788,N_4695);
nand U5450 (N_5450,N_4493,N_4608);
nand U5451 (N_5451,N_4394,N_4762);
and U5452 (N_5452,N_4768,N_4975);
and U5453 (N_5453,N_4889,N_4739);
nor U5454 (N_5454,N_4765,N_4375);
nor U5455 (N_5455,N_4693,N_4532);
nand U5456 (N_5456,N_4947,N_4699);
nor U5457 (N_5457,N_4869,N_4610);
nand U5458 (N_5458,N_4779,N_4734);
nor U5459 (N_5459,N_4862,N_4539);
xor U5460 (N_5460,N_4822,N_4562);
nor U5461 (N_5461,N_4481,N_4535);
xor U5462 (N_5462,N_4564,N_4877);
nand U5463 (N_5463,N_4521,N_4653);
xnor U5464 (N_5464,N_4407,N_4652);
and U5465 (N_5465,N_4650,N_4531);
and U5466 (N_5466,N_4657,N_4641);
nand U5467 (N_5467,N_4637,N_4584);
nand U5468 (N_5468,N_4413,N_4664);
nand U5469 (N_5469,N_4895,N_4396);
nand U5470 (N_5470,N_4386,N_4851);
and U5471 (N_5471,N_4484,N_4752);
and U5472 (N_5472,N_4412,N_4947);
nand U5473 (N_5473,N_4461,N_4875);
and U5474 (N_5474,N_4609,N_4847);
nand U5475 (N_5475,N_4826,N_4386);
nor U5476 (N_5476,N_4604,N_4529);
xnor U5477 (N_5477,N_4756,N_4534);
nand U5478 (N_5478,N_4585,N_4475);
nor U5479 (N_5479,N_4650,N_4994);
nand U5480 (N_5480,N_4877,N_4750);
or U5481 (N_5481,N_4645,N_4407);
and U5482 (N_5482,N_4574,N_4750);
nor U5483 (N_5483,N_4383,N_4408);
nor U5484 (N_5484,N_4651,N_4557);
nor U5485 (N_5485,N_4681,N_4543);
and U5486 (N_5486,N_4970,N_4473);
nor U5487 (N_5487,N_4912,N_4559);
and U5488 (N_5488,N_4812,N_4628);
or U5489 (N_5489,N_4743,N_4585);
nor U5490 (N_5490,N_4394,N_4898);
and U5491 (N_5491,N_4763,N_4874);
or U5492 (N_5492,N_4408,N_4582);
and U5493 (N_5493,N_4750,N_4583);
nor U5494 (N_5494,N_4983,N_4675);
or U5495 (N_5495,N_4981,N_4739);
xnor U5496 (N_5496,N_4853,N_4464);
and U5497 (N_5497,N_4758,N_4452);
nand U5498 (N_5498,N_4455,N_4676);
nor U5499 (N_5499,N_4418,N_4452);
xor U5500 (N_5500,N_4633,N_4663);
or U5501 (N_5501,N_4434,N_4694);
xnor U5502 (N_5502,N_4395,N_4553);
xnor U5503 (N_5503,N_4723,N_4989);
and U5504 (N_5504,N_4994,N_4381);
and U5505 (N_5505,N_4756,N_4838);
or U5506 (N_5506,N_4602,N_4509);
nand U5507 (N_5507,N_4613,N_4951);
nor U5508 (N_5508,N_4507,N_4429);
or U5509 (N_5509,N_4797,N_4920);
and U5510 (N_5510,N_4803,N_4564);
nand U5511 (N_5511,N_4535,N_4392);
nor U5512 (N_5512,N_4408,N_4738);
xnor U5513 (N_5513,N_4868,N_4695);
or U5514 (N_5514,N_4769,N_4443);
nand U5515 (N_5515,N_4673,N_4935);
nor U5516 (N_5516,N_4546,N_4766);
xor U5517 (N_5517,N_4810,N_4920);
xor U5518 (N_5518,N_4724,N_4913);
xnor U5519 (N_5519,N_4670,N_4544);
nand U5520 (N_5520,N_4805,N_4411);
nand U5521 (N_5521,N_4692,N_4960);
nand U5522 (N_5522,N_4641,N_4776);
nor U5523 (N_5523,N_4807,N_4940);
nor U5524 (N_5524,N_4633,N_4509);
nor U5525 (N_5525,N_4702,N_4951);
nand U5526 (N_5526,N_4579,N_4649);
xnor U5527 (N_5527,N_4984,N_4495);
nor U5528 (N_5528,N_4457,N_4525);
xnor U5529 (N_5529,N_4693,N_4567);
nand U5530 (N_5530,N_4838,N_4802);
nor U5531 (N_5531,N_4477,N_4922);
and U5532 (N_5532,N_4851,N_4506);
nor U5533 (N_5533,N_4579,N_4524);
and U5534 (N_5534,N_4995,N_4555);
or U5535 (N_5535,N_4742,N_4559);
or U5536 (N_5536,N_4761,N_4868);
and U5537 (N_5537,N_4996,N_4721);
xor U5538 (N_5538,N_4493,N_4522);
xor U5539 (N_5539,N_4460,N_4738);
or U5540 (N_5540,N_4791,N_4689);
nand U5541 (N_5541,N_4993,N_4991);
xnor U5542 (N_5542,N_4724,N_4547);
or U5543 (N_5543,N_4793,N_4436);
or U5544 (N_5544,N_4958,N_4670);
nand U5545 (N_5545,N_4616,N_4884);
and U5546 (N_5546,N_4949,N_4672);
and U5547 (N_5547,N_4692,N_4668);
or U5548 (N_5548,N_4411,N_4770);
and U5549 (N_5549,N_4494,N_4666);
or U5550 (N_5550,N_4881,N_4802);
nand U5551 (N_5551,N_4476,N_4939);
nand U5552 (N_5552,N_4865,N_4591);
or U5553 (N_5553,N_4615,N_4899);
nand U5554 (N_5554,N_4603,N_4462);
nand U5555 (N_5555,N_4904,N_4906);
nor U5556 (N_5556,N_4956,N_4438);
nor U5557 (N_5557,N_4577,N_4930);
nand U5558 (N_5558,N_4408,N_4795);
or U5559 (N_5559,N_4392,N_4446);
nor U5560 (N_5560,N_4644,N_4377);
or U5561 (N_5561,N_4962,N_4916);
nor U5562 (N_5562,N_4593,N_4426);
nor U5563 (N_5563,N_4997,N_4630);
nand U5564 (N_5564,N_4666,N_4817);
or U5565 (N_5565,N_4598,N_4897);
nand U5566 (N_5566,N_4759,N_4908);
xor U5567 (N_5567,N_4769,N_4792);
nor U5568 (N_5568,N_4626,N_4478);
nor U5569 (N_5569,N_4704,N_4772);
or U5570 (N_5570,N_4588,N_4719);
xor U5571 (N_5571,N_4577,N_4915);
nor U5572 (N_5572,N_4806,N_4717);
nor U5573 (N_5573,N_4673,N_4455);
nand U5574 (N_5574,N_4541,N_4416);
and U5575 (N_5575,N_4417,N_4512);
xor U5576 (N_5576,N_4654,N_4735);
and U5577 (N_5577,N_4773,N_4983);
nor U5578 (N_5578,N_4736,N_4590);
nor U5579 (N_5579,N_4648,N_4792);
nor U5580 (N_5580,N_4498,N_4514);
or U5581 (N_5581,N_4604,N_4614);
nor U5582 (N_5582,N_4659,N_4885);
nand U5583 (N_5583,N_4465,N_4868);
and U5584 (N_5584,N_4651,N_4433);
nand U5585 (N_5585,N_4519,N_4631);
or U5586 (N_5586,N_4654,N_4918);
xor U5587 (N_5587,N_4980,N_4962);
xor U5588 (N_5588,N_4721,N_4955);
or U5589 (N_5589,N_4640,N_4383);
nand U5590 (N_5590,N_4563,N_4467);
or U5591 (N_5591,N_4592,N_4893);
xnor U5592 (N_5592,N_4663,N_4691);
and U5593 (N_5593,N_4771,N_4797);
and U5594 (N_5594,N_4587,N_4646);
nor U5595 (N_5595,N_4818,N_4802);
nand U5596 (N_5596,N_4776,N_4485);
and U5597 (N_5597,N_4481,N_4949);
and U5598 (N_5598,N_4375,N_4599);
xor U5599 (N_5599,N_4694,N_4823);
nand U5600 (N_5600,N_4562,N_4851);
and U5601 (N_5601,N_4736,N_4722);
nand U5602 (N_5602,N_4566,N_4906);
or U5603 (N_5603,N_4847,N_4510);
nor U5604 (N_5604,N_4445,N_4928);
nand U5605 (N_5605,N_4871,N_4445);
nand U5606 (N_5606,N_4947,N_4473);
nor U5607 (N_5607,N_4972,N_4558);
and U5608 (N_5608,N_4528,N_4970);
xor U5609 (N_5609,N_4713,N_4701);
xor U5610 (N_5610,N_4863,N_4995);
or U5611 (N_5611,N_4458,N_4445);
nand U5612 (N_5612,N_4532,N_4718);
xor U5613 (N_5613,N_4992,N_4747);
or U5614 (N_5614,N_4968,N_4682);
nand U5615 (N_5615,N_4570,N_4951);
nor U5616 (N_5616,N_4981,N_4682);
xor U5617 (N_5617,N_4632,N_4673);
and U5618 (N_5618,N_4858,N_4409);
nor U5619 (N_5619,N_4526,N_4555);
xor U5620 (N_5620,N_4768,N_4830);
nand U5621 (N_5621,N_4761,N_4545);
nor U5622 (N_5622,N_4940,N_4673);
nor U5623 (N_5623,N_4397,N_4446);
or U5624 (N_5624,N_4703,N_4986);
xor U5625 (N_5625,N_5336,N_5398);
or U5626 (N_5626,N_5231,N_5470);
xnor U5627 (N_5627,N_5441,N_5192);
and U5628 (N_5628,N_5224,N_5418);
xor U5629 (N_5629,N_5606,N_5431);
nand U5630 (N_5630,N_5613,N_5512);
xnor U5631 (N_5631,N_5251,N_5303);
or U5632 (N_5632,N_5330,N_5164);
nand U5633 (N_5633,N_5202,N_5474);
or U5634 (N_5634,N_5346,N_5268);
nand U5635 (N_5635,N_5435,N_5142);
or U5636 (N_5636,N_5439,N_5307);
or U5637 (N_5637,N_5280,N_5538);
nand U5638 (N_5638,N_5056,N_5298);
nand U5639 (N_5639,N_5543,N_5326);
and U5640 (N_5640,N_5552,N_5456);
and U5641 (N_5641,N_5479,N_5577);
nor U5642 (N_5642,N_5249,N_5507);
nand U5643 (N_5643,N_5375,N_5215);
nor U5644 (N_5644,N_5378,N_5272);
and U5645 (N_5645,N_5173,N_5328);
or U5646 (N_5646,N_5476,N_5460);
or U5647 (N_5647,N_5137,N_5354);
or U5648 (N_5648,N_5109,N_5103);
or U5649 (N_5649,N_5132,N_5491);
and U5650 (N_5650,N_5089,N_5603);
or U5651 (N_5651,N_5204,N_5135);
and U5652 (N_5652,N_5172,N_5419);
or U5653 (N_5653,N_5558,N_5128);
nor U5654 (N_5654,N_5434,N_5495);
nor U5655 (N_5655,N_5310,N_5526);
or U5656 (N_5656,N_5285,N_5221);
xnor U5657 (N_5657,N_5390,N_5533);
nand U5658 (N_5658,N_5565,N_5403);
nor U5659 (N_5659,N_5194,N_5034);
and U5660 (N_5660,N_5212,N_5542);
nor U5661 (N_5661,N_5339,N_5246);
nand U5662 (N_5662,N_5047,N_5529);
nor U5663 (N_5663,N_5304,N_5352);
and U5664 (N_5664,N_5466,N_5196);
nand U5665 (N_5665,N_5550,N_5027);
and U5666 (N_5666,N_5618,N_5373);
and U5667 (N_5667,N_5010,N_5499);
nand U5668 (N_5668,N_5551,N_5138);
and U5669 (N_5669,N_5168,N_5450);
nand U5670 (N_5670,N_5487,N_5174);
and U5671 (N_5671,N_5165,N_5457);
xor U5672 (N_5672,N_5124,N_5623);
or U5673 (N_5673,N_5360,N_5535);
nor U5674 (N_5674,N_5478,N_5093);
nor U5675 (N_5675,N_5404,N_5199);
and U5676 (N_5676,N_5241,N_5388);
nand U5677 (N_5677,N_5144,N_5155);
xor U5678 (N_5678,N_5154,N_5362);
or U5679 (N_5679,N_5019,N_5170);
nor U5680 (N_5680,N_5073,N_5448);
nand U5681 (N_5681,N_5157,N_5006);
and U5682 (N_5682,N_5070,N_5355);
and U5683 (N_5683,N_5218,N_5277);
nor U5684 (N_5684,N_5544,N_5227);
xor U5685 (N_5685,N_5140,N_5454);
xor U5686 (N_5686,N_5267,N_5209);
nand U5687 (N_5687,N_5306,N_5119);
and U5688 (N_5688,N_5036,N_5396);
or U5689 (N_5689,N_5193,N_5051);
and U5690 (N_5690,N_5412,N_5503);
nor U5691 (N_5691,N_5402,N_5610);
and U5692 (N_5692,N_5275,N_5294);
or U5693 (N_5693,N_5612,N_5120);
nand U5694 (N_5694,N_5033,N_5320);
xnor U5695 (N_5695,N_5545,N_5270);
nor U5696 (N_5696,N_5541,N_5601);
xor U5697 (N_5697,N_5621,N_5079);
nand U5698 (N_5698,N_5096,N_5585);
nand U5699 (N_5699,N_5149,N_5175);
or U5700 (N_5700,N_5094,N_5185);
nor U5701 (N_5701,N_5325,N_5077);
nor U5702 (N_5702,N_5208,N_5205);
xnor U5703 (N_5703,N_5127,N_5288);
nor U5704 (N_5704,N_5332,N_5554);
nor U5705 (N_5705,N_5501,N_5335);
xnor U5706 (N_5706,N_5438,N_5483);
xnor U5707 (N_5707,N_5314,N_5167);
or U5708 (N_5708,N_5222,N_5578);
nand U5709 (N_5709,N_5557,N_5287);
and U5710 (N_5710,N_5570,N_5453);
or U5711 (N_5711,N_5020,N_5568);
or U5712 (N_5712,N_5273,N_5300);
and U5713 (N_5713,N_5058,N_5248);
nor U5714 (N_5714,N_5133,N_5615);
xor U5715 (N_5715,N_5038,N_5050);
and U5716 (N_5716,N_5031,N_5236);
and U5717 (N_5717,N_5350,N_5293);
nand U5718 (N_5718,N_5265,N_5309);
nor U5719 (N_5719,N_5177,N_5032);
nor U5720 (N_5720,N_5245,N_5413);
nor U5721 (N_5721,N_5493,N_5593);
nand U5722 (N_5722,N_5343,N_5214);
nor U5723 (N_5723,N_5598,N_5030);
xnor U5724 (N_5724,N_5116,N_5420);
nor U5725 (N_5725,N_5587,N_5281);
nor U5726 (N_5726,N_5594,N_5382);
nand U5727 (N_5727,N_5387,N_5411);
or U5728 (N_5728,N_5282,N_5000);
nor U5729 (N_5729,N_5301,N_5409);
nand U5730 (N_5730,N_5092,N_5376);
nand U5731 (N_5731,N_5226,N_5455);
nor U5732 (N_5732,N_5292,N_5059);
and U5733 (N_5733,N_5283,N_5473);
nand U5734 (N_5734,N_5257,N_5098);
or U5735 (N_5735,N_5276,N_5024);
nor U5736 (N_5736,N_5088,N_5083);
and U5737 (N_5737,N_5572,N_5337);
and U5738 (N_5738,N_5481,N_5009);
or U5739 (N_5739,N_5596,N_5406);
nor U5740 (N_5740,N_5198,N_5134);
nand U5741 (N_5741,N_5423,N_5016);
nand U5742 (N_5742,N_5415,N_5525);
and U5743 (N_5743,N_5148,N_5297);
or U5744 (N_5744,N_5506,N_5039);
xor U5745 (N_5745,N_5443,N_5482);
nand U5746 (N_5746,N_5232,N_5296);
or U5747 (N_5747,N_5106,N_5527);
or U5748 (N_5748,N_5317,N_5494);
xor U5749 (N_5749,N_5468,N_5052);
nand U5750 (N_5750,N_5284,N_5452);
nand U5751 (N_5751,N_5562,N_5429);
and U5752 (N_5752,N_5123,N_5595);
nand U5753 (N_5753,N_5136,N_5216);
xor U5754 (N_5754,N_5130,N_5367);
nand U5755 (N_5755,N_5159,N_5129);
nand U5756 (N_5756,N_5053,N_5278);
nor U5757 (N_5757,N_5417,N_5291);
xor U5758 (N_5758,N_5044,N_5054);
nand U5759 (N_5759,N_5080,N_5421);
or U5760 (N_5760,N_5611,N_5061);
and U5761 (N_5761,N_5266,N_5023);
or U5762 (N_5762,N_5449,N_5514);
and U5763 (N_5763,N_5437,N_5139);
nand U5764 (N_5764,N_5472,N_5290);
and U5765 (N_5765,N_5581,N_5008);
or U5766 (N_5766,N_5146,N_5046);
nand U5767 (N_5767,N_5622,N_5536);
nor U5768 (N_5768,N_5260,N_5171);
or U5769 (N_5769,N_5446,N_5496);
nand U5770 (N_5770,N_5012,N_5381);
nand U5771 (N_5771,N_5101,N_5502);
or U5772 (N_5772,N_5107,N_5063);
or U5773 (N_5773,N_5189,N_5005);
xor U5774 (N_5774,N_5097,N_5004);
xnor U5775 (N_5775,N_5584,N_5340);
xnor U5776 (N_5776,N_5111,N_5011);
and U5777 (N_5777,N_5416,N_5131);
nor U5778 (N_5778,N_5255,N_5179);
and U5779 (N_5779,N_5108,N_5197);
or U5780 (N_5780,N_5385,N_5424);
and U5781 (N_5781,N_5607,N_5374);
nor U5782 (N_5782,N_5141,N_5289);
or U5783 (N_5783,N_5516,N_5254);
xnor U5784 (N_5784,N_5567,N_5219);
xor U5785 (N_5785,N_5321,N_5384);
or U5786 (N_5786,N_5341,N_5395);
or U5787 (N_5787,N_5201,N_5488);
nor U5788 (N_5788,N_5256,N_5263);
or U5789 (N_5789,N_5361,N_5329);
xor U5790 (N_5790,N_5313,N_5143);
nand U5791 (N_5791,N_5546,N_5153);
nand U5792 (N_5792,N_5068,N_5041);
xor U5793 (N_5793,N_5553,N_5549);
xnor U5794 (N_5794,N_5532,N_5069);
nand U5795 (N_5795,N_5162,N_5002);
or U5796 (N_5796,N_5345,N_5117);
or U5797 (N_5797,N_5055,N_5427);
nand U5798 (N_5798,N_5104,N_5407);
nor U5799 (N_5799,N_5025,N_5357);
and U5800 (N_5800,N_5286,N_5334);
nor U5801 (N_5801,N_5566,N_5178);
or U5802 (N_5802,N_5436,N_5299);
nor U5803 (N_5803,N_5302,N_5014);
nand U5804 (N_5804,N_5017,N_5353);
or U5805 (N_5805,N_5368,N_5377);
or U5806 (N_5806,N_5405,N_5308);
or U5807 (N_5807,N_5616,N_5391);
xnor U5808 (N_5808,N_5358,N_5344);
and U5809 (N_5809,N_5191,N_5045);
and U5810 (N_5810,N_5370,N_5327);
xnor U5811 (N_5811,N_5105,N_5576);
xor U5812 (N_5812,N_5084,N_5430);
nand U5813 (N_5813,N_5166,N_5590);
or U5814 (N_5814,N_5180,N_5331);
nand U5815 (N_5815,N_5071,N_5062);
nand U5816 (N_5816,N_5564,N_5262);
nor U5817 (N_5817,N_5145,N_5264);
xnor U5818 (N_5818,N_5190,N_5312);
xnor U5819 (N_5819,N_5239,N_5181);
or U5820 (N_5820,N_5095,N_5086);
nor U5821 (N_5821,N_5515,N_5234);
nor U5822 (N_5822,N_5614,N_5509);
xnor U5823 (N_5823,N_5579,N_5349);
nor U5824 (N_5824,N_5161,N_5573);
and U5825 (N_5825,N_5575,N_5351);
xor U5826 (N_5826,N_5559,N_5015);
nor U5827 (N_5827,N_5067,N_5305);
or U5828 (N_5828,N_5311,N_5432);
and U5829 (N_5829,N_5447,N_5235);
nor U5830 (N_5830,N_5486,N_5492);
or U5831 (N_5831,N_5158,N_5469);
and U5832 (N_5832,N_5480,N_5467);
xnor U5833 (N_5833,N_5237,N_5091);
and U5834 (N_5834,N_5534,N_5600);
nor U5835 (N_5835,N_5003,N_5065);
xnor U5836 (N_5836,N_5490,N_5521);
nand U5837 (N_5837,N_5125,N_5078);
nor U5838 (N_5838,N_5115,N_5605);
or U5839 (N_5839,N_5364,N_5592);
or U5840 (N_5840,N_5497,N_5026);
nand U5841 (N_5841,N_5464,N_5114);
nor U5842 (N_5842,N_5022,N_5574);
xor U5843 (N_5843,N_5356,N_5323);
and U5844 (N_5844,N_5414,N_5445);
nor U5845 (N_5845,N_5150,N_5258);
or U5846 (N_5846,N_5118,N_5090);
and U5847 (N_5847,N_5505,N_5617);
and U5848 (N_5848,N_5518,N_5583);
nor U5849 (N_5849,N_5485,N_5560);
xnor U5850 (N_5850,N_5064,N_5540);
nand U5851 (N_5851,N_5066,N_5184);
and U5852 (N_5852,N_5333,N_5548);
xor U5853 (N_5853,N_5571,N_5524);
xor U5854 (N_5854,N_5624,N_5348);
or U5855 (N_5855,N_5425,N_5458);
or U5856 (N_5856,N_5028,N_5187);
or U5857 (N_5857,N_5207,N_5608);
nor U5858 (N_5858,N_5182,N_5569);
nor U5859 (N_5859,N_5253,N_5126);
nor U5860 (N_5860,N_5539,N_5556);
nand U5861 (N_5861,N_5463,N_5229);
xor U5862 (N_5862,N_5510,N_5233);
or U5863 (N_5863,N_5206,N_5408);
and U5864 (N_5864,N_5599,N_5271);
xor U5865 (N_5865,N_5604,N_5049);
and U5866 (N_5866,N_5589,N_5243);
xor U5867 (N_5867,N_5561,N_5359);
nor U5868 (N_5868,N_5394,N_5244);
xnor U5869 (N_5869,N_5471,N_5082);
or U5870 (N_5870,N_5160,N_5322);
nand U5871 (N_5871,N_5588,N_5563);
nand U5872 (N_5872,N_5440,N_5001);
xor U5873 (N_5873,N_5156,N_5318);
and U5874 (N_5874,N_5152,N_5007);
nor U5875 (N_5875,N_5230,N_5081);
nand U5876 (N_5876,N_5465,N_5511);
nand U5877 (N_5877,N_5528,N_5547);
and U5878 (N_5878,N_5057,N_5462);
or U5879 (N_5879,N_5250,N_5371);
nor U5880 (N_5880,N_5113,N_5484);
or U5881 (N_5881,N_5169,N_5225);
nor U5882 (N_5882,N_5461,N_5021);
and U5883 (N_5883,N_5163,N_5085);
nor U5884 (N_5884,N_5043,N_5295);
nor U5885 (N_5885,N_5099,N_5217);
or U5886 (N_5886,N_5151,N_5074);
nor U5887 (N_5887,N_5520,N_5517);
nand U5888 (N_5888,N_5338,N_5386);
nand U5889 (N_5889,N_5220,N_5238);
or U5890 (N_5890,N_5347,N_5279);
and U5891 (N_5891,N_5397,N_5075);
nor U5892 (N_5892,N_5498,N_5203);
xor U5893 (N_5893,N_5620,N_5087);
nand U5894 (N_5894,N_5223,N_5242);
and U5895 (N_5895,N_5580,N_5228);
nand U5896 (N_5896,N_5112,N_5324);
and U5897 (N_5897,N_5316,N_5513);
nor U5898 (N_5898,N_5319,N_5372);
or U5899 (N_5899,N_5048,N_5186);
nand U5900 (N_5900,N_5619,N_5428);
and U5901 (N_5901,N_5389,N_5500);
and U5902 (N_5902,N_5530,N_5060);
and U5903 (N_5903,N_5200,N_5100);
nor U5904 (N_5904,N_5076,N_5013);
nand U5905 (N_5905,N_5602,N_5029);
or U5906 (N_5906,N_5401,N_5121);
xnor U5907 (N_5907,N_5147,N_5379);
and U5908 (N_5908,N_5110,N_5261);
nand U5909 (N_5909,N_5591,N_5537);
or U5910 (N_5910,N_5426,N_5040);
xor U5911 (N_5911,N_5363,N_5042);
xor U5912 (N_5912,N_5422,N_5508);
or U5913 (N_5913,N_5442,N_5475);
nand U5914 (N_5914,N_5176,N_5400);
xnor U5915 (N_5915,N_5451,N_5519);
nand U5916 (N_5916,N_5582,N_5213);
and U5917 (N_5917,N_5555,N_5410);
or U5918 (N_5918,N_5210,N_5342);
nand U5919 (N_5919,N_5609,N_5240);
nor U5920 (N_5920,N_5315,N_5035);
nand U5921 (N_5921,N_5597,N_5444);
xor U5922 (N_5922,N_5183,N_5369);
nand U5923 (N_5923,N_5274,N_5489);
nor U5924 (N_5924,N_5247,N_5037);
nor U5925 (N_5925,N_5269,N_5366);
or U5926 (N_5926,N_5383,N_5252);
nor U5927 (N_5927,N_5018,N_5072);
and U5928 (N_5928,N_5433,N_5393);
nor U5929 (N_5929,N_5380,N_5459);
nand U5930 (N_5930,N_5531,N_5399);
or U5931 (N_5931,N_5259,N_5522);
xnor U5932 (N_5932,N_5195,N_5586);
or U5933 (N_5933,N_5392,N_5477);
nand U5934 (N_5934,N_5365,N_5122);
nand U5935 (N_5935,N_5211,N_5102);
nand U5936 (N_5936,N_5188,N_5504);
or U5937 (N_5937,N_5523,N_5316);
xor U5938 (N_5938,N_5453,N_5496);
xnor U5939 (N_5939,N_5622,N_5142);
nand U5940 (N_5940,N_5131,N_5555);
and U5941 (N_5941,N_5320,N_5282);
xnor U5942 (N_5942,N_5466,N_5013);
xnor U5943 (N_5943,N_5269,N_5401);
and U5944 (N_5944,N_5259,N_5426);
nand U5945 (N_5945,N_5545,N_5594);
nand U5946 (N_5946,N_5042,N_5586);
nand U5947 (N_5947,N_5155,N_5196);
nand U5948 (N_5948,N_5203,N_5483);
or U5949 (N_5949,N_5543,N_5423);
xnor U5950 (N_5950,N_5445,N_5321);
nand U5951 (N_5951,N_5114,N_5160);
xor U5952 (N_5952,N_5612,N_5385);
and U5953 (N_5953,N_5110,N_5517);
nand U5954 (N_5954,N_5007,N_5469);
and U5955 (N_5955,N_5396,N_5235);
or U5956 (N_5956,N_5244,N_5623);
nand U5957 (N_5957,N_5468,N_5032);
nor U5958 (N_5958,N_5452,N_5426);
xnor U5959 (N_5959,N_5185,N_5368);
xor U5960 (N_5960,N_5076,N_5397);
and U5961 (N_5961,N_5400,N_5612);
nand U5962 (N_5962,N_5019,N_5066);
nand U5963 (N_5963,N_5098,N_5387);
nor U5964 (N_5964,N_5546,N_5057);
and U5965 (N_5965,N_5268,N_5397);
or U5966 (N_5966,N_5447,N_5187);
nand U5967 (N_5967,N_5323,N_5251);
and U5968 (N_5968,N_5287,N_5014);
and U5969 (N_5969,N_5416,N_5207);
or U5970 (N_5970,N_5601,N_5438);
nand U5971 (N_5971,N_5421,N_5548);
nor U5972 (N_5972,N_5586,N_5240);
or U5973 (N_5973,N_5194,N_5557);
and U5974 (N_5974,N_5444,N_5279);
or U5975 (N_5975,N_5477,N_5235);
and U5976 (N_5976,N_5609,N_5547);
xnor U5977 (N_5977,N_5365,N_5107);
nand U5978 (N_5978,N_5230,N_5366);
xor U5979 (N_5979,N_5286,N_5586);
or U5980 (N_5980,N_5109,N_5300);
xor U5981 (N_5981,N_5422,N_5507);
xor U5982 (N_5982,N_5567,N_5088);
nand U5983 (N_5983,N_5369,N_5409);
and U5984 (N_5984,N_5270,N_5122);
nor U5985 (N_5985,N_5187,N_5140);
nand U5986 (N_5986,N_5389,N_5224);
nor U5987 (N_5987,N_5248,N_5152);
and U5988 (N_5988,N_5478,N_5544);
nor U5989 (N_5989,N_5153,N_5381);
nand U5990 (N_5990,N_5616,N_5481);
xnor U5991 (N_5991,N_5594,N_5044);
and U5992 (N_5992,N_5194,N_5226);
and U5993 (N_5993,N_5145,N_5371);
and U5994 (N_5994,N_5252,N_5533);
nor U5995 (N_5995,N_5393,N_5424);
or U5996 (N_5996,N_5221,N_5173);
xnor U5997 (N_5997,N_5146,N_5005);
or U5998 (N_5998,N_5305,N_5273);
xnor U5999 (N_5999,N_5529,N_5024);
or U6000 (N_6000,N_5400,N_5075);
nand U6001 (N_6001,N_5571,N_5008);
or U6002 (N_6002,N_5570,N_5331);
or U6003 (N_6003,N_5255,N_5077);
and U6004 (N_6004,N_5451,N_5583);
nor U6005 (N_6005,N_5517,N_5567);
xor U6006 (N_6006,N_5322,N_5312);
and U6007 (N_6007,N_5041,N_5187);
and U6008 (N_6008,N_5589,N_5595);
or U6009 (N_6009,N_5001,N_5488);
xnor U6010 (N_6010,N_5309,N_5554);
nand U6011 (N_6011,N_5128,N_5160);
and U6012 (N_6012,N_5343,N_5108);
or U6013 (N_6013,N_5006,N_5349);
xor U6014 (N_6014,N_5076,N_5185);
or U6015 (N_6015,N_5434,N_5543);
nor U6016 (N_6016,N_5371,N_5150);
xnor U6017 (N_6017,N_5017,N_5039);
and U6018 (N_6018,N_5616,N_5141);
and U6019 (N_6019,N_5515,N_5363);
or U6020 (N_6020,N_5187,N_5536);
xnor U6021 (N_6021,N_5485,N_5282);
and U6022 (N_6022,N_5601,N_5132);
xnor U6023 (N_6023,N_5613,N_5488);
xnor U6024 (N_6024,N_5401,N_5585);
and U6025 (N_6025,N_5033,N_5175);
or U6026 (N_6026,N_5329,N_5032);
or U6027 (N_6027,N_5475,N_5562);
xor U6028 (N_6028,N_5192,N_5497);
and U6029 (N_6029,N_5173,N_5104);
nor U6030 (N_6030,N_5274,N_5276);
xnor U6031 (N_6031,N_5523,N_5230);
nor U6032 (N_6032,N_5444,N_5064);
nor U6033 (N_6033,N_5309,N_5529);
nand U6034 (N_6034,N_5266,N_5106);
xnor U6035 (N_6035,N_5238,N_5225);
nor U6036 (N_6036,N_5135,N_5216);
and U6037 (N_6037,N_5337,N_5037);
xor U6038 (N_6038,N_5416,N_5519);
nor U6039 (N_6039,N_5579,N_5157);
xnor U6040 (N_6040,N_5460,N_5613);
or U6041 (N_6041,N_5216,N_5342);
nand U6042 (N_6042,N_5576,N_5247);
and U6043 (N_6043,N_5618,N_5138);
or U6044 (N_6044,N_5544,N_5128);
nor U6045 (N_6045,N_5337,N_5246);
nor U6046 (N_6046,N_5621,N_5514);
nor U6047 (N_6047,N_5047,N_5564);
nor U6048 (N_6048,N_5209,N_5164);
nand U6049 (N_6049,N_5035,N_5140);
or U6050 (N_6050,N_5215,N_5144);
xor U6051 (N_6051,N_5248,N_5424);
or U6052 (N_6052,N_5265,N_5220);
or U6053 (N_6053,N_5273,N_5133);
xnor U6054 (N_6054,N_5267,N_5430);
nor U6055 (N_6055,N_5207,N_5216);
nor U6056 (N_6056,N_5603,N_5186);
and U6057 (N_6057,N_5427,N_5299);
nor U6058 (N_6058,N_5261,N_5014);
and U6059 (N_6059,N_5070,N_5296);
nand U6060 (N_6060,N_5473,N_5308);
nand U6061 (N_6061,N_5350,N_5228);
and U6062 (N_6062,N_5141,N_5165);
nor U6063 (N_6063,N_5460,N_5481);
nor U6064 (N_6064,N_5555,N_5533);
or U6065 (N_6065,N_5213,N_5123);
nor U6066 (N_6066,N_5155,N_5505);
and U6067 (N_6067,N_5583,N_5192);
or U6068 (N_6068,N_5021,N_5134);
xor U6069 (N_6069,N_5119,N_5058);
and U6070 (N_6070,N_5241,N_5408);
and U6071 (N_6071,N_5530,N_5097);
nor U6072 (N_6072,N_5252,N_5489);
or U6073 (N_6073,N_5399,N_5043);
nor U6074 (N_6074,N_5400,N_5034);
and U6075 (N_6075,N_5101,N_5246);
nand U6076 (N_6076,N_5285,N_5256);
nand U6077 (N_6077,N_5388,N_5112);
xor U6078 (N_6078,N_5454,N_5195);
nand U6079 (N_6079,N_5212,N_5367);
nor U6080 (N_6080,N_5265,N_5351);
xnor U6081 (N_6081,N_5058,N_5143);
xor U6082 (N_6082,N_5105,N_5139);
and U6083 (N_6083,N_5393,N_5098);
nand U6084 (N_6084,N_5153,N_5457);
and U6085 (N_6085,N_5368,N_5227);
or U6086 (N_6086,N_5113,N_5125);
nor U6087 (N_6087,N_5591,N_5007);
nor U6088 (N_6088,N_5078,N_5521);
or U6089 (N_6089,N_5007,N_5032);
nand U6090 (N_6090,N_5573,N_5225);
and U6091 (N_6091,N_5285,N_5353);
nor U6092 (N_6092,N_5442,N_5578);
and U6093 (N_6093,N_5414,N_5204);
nor U6094 (N_6094,N_5369,N_5014);
xor U6095 (N_6095,N_5553,N_5585);
and U6096 (N_6096,N_5353,N_5119);
or U6097 (N_6097,N_5108,N_5159);
and U6098 (N_6098,N_5281,N_5623);
nor U6099 (N_6099,N_5066,N_5339);
and U6100 (N_6100,N_5204,N_5020);
nor U6101 (N_6101,N_5280,N_5142);
nor U6102 (N_6102,N_5177,N_5498);
nand U6103 (N_6103,N_5455,N_5222);
xnor U6104 (N_6104,N_5335,N_5540);
nor U6105 (N_6105,N_5119,N_5017);
nand U6106 (N_6106,N_5037,N_5539);
nor U6107 (N_6107,N_5185,N_5429);
and U6108 (N_6108,N_5403,N_5442);
xor U6109 (N_6109,N_5037,N_5192);
nor U6110 (N_6110,N_5329,N_5264);
nor U6111 (N_6111,N_5588,N_5599);
and U6112 (N_6112,N_5531,N_5043);
nand U6113 (N_6113,N_5021,N_5469);
nand U6114 (N_6114,N_5515,N_5322);
xnor U6115 (N_6115,N_5277,N_5129);
or U6116 (N_6116,N_5088,N_5493);
nand U6117 (N_6117,N_5320,N_5618);
nand U6118 (N_6118,N_5182,N_5479);
or U6119 (N_6119,N_5164,N_5490);
or U6120 (N_6120,N_5484,N_5108);
nand U6121 (N_6121,N_5146,N_5374);
and U6122 (N_6122,N_5134,N_5253);
and U6123 (N_6123,N_5150,N_5202);
nor U6124 (N_6124,N_5502,N_5057);
nand U6125 (N_6125,N_5339,N_5542);
xnor U6126 (N_6126,N_5523,N_5282);
and U6127 (N_6127,N_5171,N_5402);
or U6128 (N_6128,N_5591,N_5115);
nand U6129 (N_6129,N_5024,N_5395);
nand U6130 (N_6130,N_5264,N_5064);
nor U6131 (N_6131,N_5028,N_5378);
or U6132 (N_6132,N_5611,N_5000);
nor U6133 (N_6133,N_5561,N_5102);
nor U6134 (N_6134,N_5276,N_5212);
or U6135 (N_6135,N_5527,N_5305);
and U6136 (N_6136,N_5439,N_5462);
nor U6137 (N_6137,N_5215,N_5263);
and U6138 (N_6138,N_5598,N_5020);
and U6139 (N_6139,N_5478,N_5126);
or U6140 (N_6140,N_5318,N_5495);
xor U6141 (N_6141,N_5338,N_5348);
nor U6142 (N_6142,N_5006,N_5516);
xnor U6143 (N_6143,N_5334,N_5421);
nor U6144 (N_6144,N_5003,N_5331);
nor U6145 (N_6145,N_5030,N_5441);
nor U6146 (N_6146,N_5285,N_5196);
and U6147 (N_6147,N_5144,N_5576);
xor U6148 (N_6148,N_5579,N_5442);
nand U6149 (N_6149,N_5481,N_5278);
xnor U6150 (N_6150,N_5554,N_5261);
nand U6151 (N_6151,N_5118,N_5586);
and U6152 (N_6152,N_5183,N_5227);
or U6153 (N_6153,N_5347,N_5397);
or U6154 (N_6154,N_5218,N_5084);
or U6155 (N_6155,N_5436,N_5581);
xnor U6156 (N_6156,N_5201,N_5153);
and U6157 (N_6157,N_5317,N_5171);
or U6158 (N_6158,N_5098,N_5567);
and U6159 (N_6159,N_5059,N_5135);
or U6160 (N_6160,N_5087,N_5407);
nor U6161 (N_6161,N_5317,N_5273);
xnor U6162 (N_6162,N_5151,N_5597);
or U6163 (N_6163,N_5321,N_5376);
or U6164 (N_6164,N_5392,N_5261);
nand U6165 (N_6165,N_5005,N_5002);
xnor U6166 (N_6166,N_5366,N_5543);
nor U6167 (N_6167,N_5353,N_5189);
nor U6168 (N_6168,N_5540,N_5065);
or U6169 (N_6169,N_5161,N_5009);
xnor U6170 (N_6170,N_5356,N_5505);
xnor U6171 (N_6171,N_5189,N_5290);
and U6172 (N_6172,N_5186,N_5300);
nor U6173 (N_6173,N_5514,N_5330);
or U6174 (N_6174,N_5157,N_5232);
nand U6175 (N_6175,N_5537,N_5531);
and U6176 (N_6176,N_5088,N_5223);
xnor U6177 (N_6177,N_5061,N_5182);
or U6178 (N_6178,N_5187,N_5334);
xor U6179 (N_6179,N_5037,N_5003);
nor U6180 (N_6180,N_5141,N_5149);
nand U6181 (N_6181,N_5493,N_5263);
or U6182 (N_6182,N_5134,N_5276);
and U6183 (N_6183,N_5038,N_5572);
nand U6184 (N_6184,N_5415,N_5040);
nor U6185 (N_6185,N_5353,N_5234);
xor U6186 (N_6186,N_5305,N_5495);
xnor U6187 (N_6187,N_5439,N_5141);
xor U6188 (N_6188,N_5179,N_5047);
or U6189 (N_6189,N_5621,N_5087);
xnor U6190 (N_6190,N_5188,N_5065);
xnor U6191 (N_6191,N_5128,N_5456);
and U6192 (N_6192,N_5413,N_5192);
xnor U6193 (N_6193,N_5190,N_5397);
nor U6194 (N_6194,N_5388,N_5138);
nor U6195 (N_6195,N_5304,N_5500);
xor U6196 (N_6196,N_5359,N_5286);
nor U6197 (N_6197,N_5256,N_5502);
xnor U6198 (N_6198,N_5088,N_5106);
nand U6199 (N_6199,N_5042,N_5320);
nor U6200 (N_6200,N_5596,N_5369);
xor U6201 (N_6201,N_5470,N_5455);
xor U6202 (N_6202,N_5137,N_5223);
and U6203 (N_6203,N_5514,N_5024);
nor U6204 (N_6204,N_5243,N_5075);
or U6205 (N_6205,N_5157,N_5074);
nand U6206 (N_6206,N_5250,N_5515);
nor U6207 (N_6207,N_5145,N_5398);
xnor U6208 (N_6208,N_5134,N_5211);
nor U6209 (N_6209,N_5624,N_5503);
and U6210 (N_6210,N_5026,N_5442);
and U6211 (N_6211,N_5529,N_5123);
or U6212 (N_6212,N_5490,N_5601);
xor U6213 (N_6213,N_5157,N_5222);
and U6214 (N_6214,N_5511,N_5146);
nand U6215 (N_6215,N_5244,N_5128);
and U6216 (N_6216,N_5566,N_5293);
nand U6217 (N_6217,N_5022,N_5489);
nor U6218 (N_6218,N_5021,N_5066);
or U6219 (N_6219,N_5098,N_5535);
nor U6220 (N_6220,N_5362,N_5591);
nor U6221 (N_6221,N_5618,N_5188);
xnor U6222 (N_6222,N_5215,N_5589);
and U6223 (N_6223,N_5109,N_5018);
nand U6224 (N_6224,N_5451,N_5453);
or U6225 (N_6225,N_5576,N_5242);
nor U6226 (N_6226,N_5236,N_5214);
or U6227 (N_6227,N_5271,N_5153);
xnor U6228 (N_6228,N_5304,N_5022);
and U6229 (N_6229,N_5118,N_5391);
xor U6230 (N_6230,N_5076,N_5525);
nor U6231 (N_6231,N_5076,N_5533);
xor U6232 (N_6232,N_5477,N_5029);
xor U6233 (N_6233,N_5464,N_5486);
nor U6234 (N_6234,N_5280,N_5452);
nor U6235 (N_6235,N_5555,N_5051);
nand U6236 (N_6236,N_5312,N_5003);
nor U6237 (N_6237,N_5173,N_5429);
nand U6238 (N_6238,N_5361,N_5402);
nand U6239 (N_6239,N_5085,N_5057);
and U6240 (N_6240,N_5579,N_5471);
nand U6241 (N_6241,N_5481,N_5153);
or U6242 (N_6242,N_5348,N_5572);
xor U6243 (N_6243,N_5504,N_5361);
or U6244 (N_6244,N_5400,N_5349);
and U6245 (N_6245,N_5047,N_5231);
and U6246 (N_6246,N_5121,N_5390);
nor U6247 (N_6247,N_5052,N_5002);
and U6248 (N_6248,N_5360,N_5068);
or U6249 (N_6249,N_5346,N_5014);
xnor U6250 (N_6250,N_6082,N_5732);
nand U6251 (N_6251,N_5711,N_5660);
or U6252 (N_6252,N_5943,N_6060);
nor U6253 (N_6253,N_5892,N_5995);
and U6254 (N_6254,N_6166,N_5749);
nor U6255 (N_6255,N_6225,N_5735);
nand U6256 (N_6256,N_6046,N_6196);
and U6257 (N_6257,N_5885,N_6138);
and U6258 (N_6258,N_6001,N_5987);
and U6259 (N_6259,N_5716,N_5811);
xnor U6260 (N_6260,N_6213,N_5993);
xnor U6261 (N_6261,N_5858,N_6154);
nor U6262 (N_6262,N_5849,N_5954);
xor U6263 (N_6263,N_6158,N_5707);
xnor U6264 (N_6264,N_6179,N_5780);
xnor U6265 (N_6265,N_5742,N_5709);
nand U6266 (N_6266,N_5775,N_6110);
nor U6267 (N_6267,N_5792,N_6209);
or U6268 (N_6268,N_6047,N_6002);
or U6269 (N_6269,N_5673,N_5700);
nor U6270 (N_6270,N_5865,N_6059);
or U6271 (N_6271,N_5848,N_6030);
or U6272 (N_6272,N_5836,N_5837);
or U6273 (N_6273,N_6193,N_5766);
or U6274 (N_6274,N_6122,N_5840);
xor U6275 (N_6275,N_5860,N_6100);
and U6276 (N_6276,N_5650,N_6086);
and U6277 (N_6277,N_5701,N_5908);
or U6278 (N_6278,N_6147,N_6029);
or U6279 (N_6279,N_5887,N_6164);
nor U6280 (N_6280,N_5740,N_6071);
or U6281 (N_6281,N_6113,N_6244);
nor U6282 (N_6282,N_5714,N_6243);
xnor U6283 (N_6283,N_5658,N_5875);
nand U6284 (N_6284,N_5758,N_6211);
nand U6285 (N_6285,N_5656,N_5910);
and U6286 (N_6286,N_6024,N_6098);
xnor U6287 (N_6287,N_5893,N_5816);
or U6288 (N_6288,N_5654,N_5730);
nand U6289 (N_6289,N_5924,N_5917);
and U6290 (N_6290,N_6016,N_6067);
or U6291 (N_6291,N_6177,N_6132);
xnor U6292 (N_6292,N_5810,N_5722);
nor U6293 (N_6293,N_6136,N_6124);
xnor U6294 (N_6294,N_6176,N_5713);
nor U6295 (N_6295,N_5876,N_5867);
nand U6296 (N_6296,N_5643,N_6246);
or U6297 (N_6297,N_5747,N_6237);
nor U6298 (N_6298,N_6068,N_6129);
and U6299 (N_6299,N_6148,N_5774);
nor U6300 (N_6300,N_5677,N_5838);
or U6301 (N_6301,N_5659,N_5800);
xor U6302 (N_6302,N_6008,N_5681);
or U6303 (N_6303,N_5955,N_5771);
nor U6304 (N_6304,N_5731,N_5894);
xor U6305 (N_6305,N_5990,N_6131);
nand U6306 (N_6306,N_5630,N_5627);
nor U6307 (N_6307,N_5631,N_5895);
nor U6308 (N_6308,N_5717,N_5920);
xnor U6309 (N_6309,N_5765,N_5914);
nor U6310 (N_6310,N_6052,N_6201);
or U6311 (N_6311,N_5632,N_6037);
nor U6312 (N_6312,N_5915,N_6162);
xnor U6313 (N_6313,N_5845,N_5842);
or U6314 (N_6314,N_6096,N_5980);
xnor U6315 (N_6315,N_5853,N_5657);
and U6316 (N_6316,N_5629,N_5738);
xor U6317 (N_6317,N_5695,N_6218);
nand U6318 (N_6318,N_5906,N_6224);
xor U6319 (N_6319,N_6116,N_6019);
nand U6320 (N_6320,N_5830,N_6123);
xor U6321 (N_6321,N_5704,N_5667);
nand U6322 (N_6322,N_6161,N_6175);
or U6323 (N_6323,N_5922,N_5739);
or U6324 (N_6324,N_6007,N_6012);
or U6325 (N_6325,N_6080,N_6157);
nor U6326 (N_6326,N_5851,N_5689);
or U6327 (N_6327,N_5850,N_5970);
nor U6328 (N_6328,N_6040,N_5905);
nor U6329 (N_6329,N_5690,N_6222);
or U6330 (N_6330,N_6145,N_5813);
xor U6331 (N_6331,N_6069,N_6079);
nand U6332 (N_6332,N_6010,N_5769);
nand U6333 (N_6333,N_5823,N_6039);
or U6334 (N_6334,N_5699,N_5685);
and U6335 (N_6335,N_5821,N_6167);
nand U6336 (N_6336,N_6054,N_6089);
or U6337 (N_6337,N_5641,N_5957);
nor U6338 (N_6338,N_5818,N_6202);
nor U6339 (N_6339,N_5642,N_5975);
or U6340 (N_6340,N_5686,N_5934);
or U6341 (N_6341,N_5812,N_6018);
and U6342 (N_6342,N_5814,N_5972);
nand U6343 (N_6343,N_5904,N_5844);
and U6344 (N_6344,N_5947,N_6107);
and U6345 (N_6345,N_5843,N_5804);
or U6346 (N_6346,N_5918,N_5940);
and U6347 (N_6347,N_6231,N_6185);
xor U6348 (N_6348,N_6173,N_6205);
nand U6349 (N_6349,N_6045,N_5856);
or U6350 (N_6350,N_6005,N_5662);
nand U6351 (N_6351,N_5978,N_6027);
nor U6352 (N_6352,N_5694,N_5863);
nor U6353 (N_6353,N_5712,N_5808);
nand U6354 (N_6354,N_5870,N_5839);
or U6355 (N_6355,N_6076,N_6223);
nor U6356 (N_6356,N_6014,N_5764);
xor U6357 (N_6357,N_5637,N_6017);
nor U6358 (N_6358,N_5859,N_5974);
or U6359 (N_6359,N_6233,N_5734);
and U6360 (N_6360,N_6153,N_5939);
nand U6361 (N_6361,N_5973,N_5669);
xor U6362 (N_6362,N_6190,N_5628);
or U6363 (N_6363,N_5799,N_5687);
and U6364 (N_6364,N_5756,N_6245);
nand U6365 (N_6365,N_6065,N_6150);
nand U6366 (N_6366,N_6200,N_5919);
nor U6367 (N_6367,N_6178,N_6084);
nor U6368 (N_6368,N_5877,N_5868);
and U6369 (N_6369,N_5929,N_5959);
or U6370 (N_6370,N_6044,N_5889);
nand U6371 (N_6371,N_5753,N_6187);
or U6372 (N_6372,N_5761,N_5744);
nor U6373 (N_6373,N_6104,N_6035);
nor U6374 (N_6374,N_5805,N_5933);
xor U6375 (N_6375,N_6056,N_5796);
nor U6376 (N_6376,N_6151,N_5666);
nand U6377 (N_6377,N_6058,N_5748);
xor U6378 (N_6378,N_5896,N_5646);
nand U6379 (N_6379,N_6064,N_6133);
or U6380 (N_6380,N_5872,N_5634);
xnor U6381 (N_6381,N_6048,N_5942);
nand U6382 (N_6382,N_6234,N_6235);
or U6383 (N_6383,N_5930,N_6249);
xor U6384 (N_6384,N_5785,N_6183);
and U6385 (N_6385,N_5652,N_5854);
xnor U6386 (N_6386,N_5724,N_5790);
or U6387 (N_6387,N_5997,N_5871);
and U6388 (N_6388,N_5971,N_5831);
xor U6389 (N_6389,N_5626,N_5874);
nand U6390 (N_6390,N_5991,N_6043);
nand U6391 (N_6391,N_6051,N_6191);
and U6392 (N_6392,N_6203,N_5788);
nand U6393 (N_6393,N_6006,N_6165);
and U6394 (N_6394,N_6011,N_5952);
xnor U6395 (N_6395,N_6214,N_6057);
and U6396 (N_6396,N_6220,N_5902);
nor U6397 (N_6397,N_6152,N_5625);
and U6398 (N_6398,N_6228,N_5819);
nor U6399 (N_6399,N_5644,N_5638);
or U6400 (N_6400,N_5981,N_5710);
xor U6401 (N_6401,N_6236,N_5891);
or U6402 (N_6402,N_5721,N_6090);
xnor U6403 (N_6403,N_6119,N_6210);
nor U6404 (N_6404,N_6171,N_6066);
nor U6405 (N_6405,N_6240,N_6004);
nor U6406 (N_6406,N_5679,N_6112);
nand U6407 (N_6407,N_5963,N_5697);
nor U6408 (N_6408,N_5873,N_5647);
or U6409 (N_6409,N_5960,N_5862);
nor U6410 (N_6410,N_5635,N_6031);
nor U6411 (N_6411,N_6070,N_6074);
nor U6412 (N_6412,N_6195,N_6168);
nor U6413 (N_6413,N_6118,N_5882);
or U6414 (N_6414,N_5757,N_5852);
and U6415 (N_6415,N_5857,N_5988);
nor U6416 (N_6416,N_5855,N_6239);
or U6417 (N_6417,N_5822,N_5928);
or U6418 (N_6418,N_5648,N_5898);
or U6419 (N_6419,N_6063,N_5983);
xnor U6420 (N_6420,N_5633,N_5977);
nand U6421 (N_6421,N_5664,N_5976);
and U6422 (N_6422,N_6127,N_5961);
nor U6423 (N_6423,N_5782,N_6053);
nor U6424 (N_6424,N_6221,N_5936);
or U6425 (N_6425,N_6186,N_5797);
and U6426 (N_6426,N_6212,N_5706);
xor U6427 (N_6427,N_6182,N_6207);
nor U6428 (N_6428,N_5846,N_5927);
and U6429 (N_6429,N_5807,N_6038);
nor U6430 (N_6430,N_6003,N_5682);
nand U6431 (N_6431,N_6026,N_6238);
or U6432 (N_6432,N_6219,N_6134);
nor U6433 (N_6433,N_6033,N_5937);
and U6434 (N_6434,N_6117,N_5880);
nand U6435 (N_6435,N_5678,N_5789);
xor U6436 (N_6436,N_5639,N_5941);
nand U6437 (N_6437,N_5826,N_5878);
nand U6438 (N_6438,N_6242,N_5921);
or U6439 (N_6439,N_5802,N_6083);
nor U6440 (N_6440,N_5696,N_5938);
xnor U6441 (N_6441,N_5786,N_6232);
nand U6442 (N_6442,N_5817,N_6049);
or U6443 (N_6443,N_6075,N_6130);
nand U6444 (N_6444,N_5994,N_6072);
or U6445 (N_6445,N_5967,N_6102);
nor U6446 (N_6446,N_5835,N_5645);
nor U6447 (N_6447,N_5798,N_6229);
nor U6448 (N_6448,N_6188,N_5864);
and U6449 (N_6449,N_6120,N_5890);
and U6450 (N_6450,N_6143,N_5661);
or U6451 (N_6451,N_6140,N_5999);
and U6452 (N_6452,N_5932,N_6174);
nand U6453 (N_6453,N_5897,N_5841);
or U6454 (N_6454,N_6170,N_5760);
nor U6455 (N_6455,N_5965,N_6189);
xor U6456 (N_6456,N_6103,N_5801);
nand U6457 (N_6457,N_5825,N_6204);
nand U6458 (N_6458,N_5698,N_6169);
and U6459 (N_6459,N_5665,N_6055);
nand U6460 (N_6460,N_6241,N_5705);
or U6461 (N_6461,N_5833,N_5672);
and U6462 (N_6462,N_5779,N_5773);
and U6463 (N_6463,N_6216,N_5829);
or U6464 (N_6464,N_5777,N_6036);
xnor U6465 (N_6465,N_6105,N_5916);
or U6466 (N_6466,N_5718,N_5985);
nor U6467 (N_6467,N_5886,N_5725);
xnor U6468 (N_6468,N_5989,N_5945);
and U6469 (N_6469,N_5969,N_5900);
xor U6470 (N_6470,N_6226,N_6156);
nand U6471 (N_6471,N_6081,N_5772);
xnor U6472 (N_6472,N_5884,N_5762);
nor U6473 (N_6473,N_6013,N_5733);
xnor U6474 (N_6474,N_5888,N_5719);
and U6475 (N_6475,N_5692,N_5913);
nor U6476 (N_6476,N_6172,N_5815);
and U6477 (N_6477,N_5684,N_5794);
nor U6478 (N_6478,N_5741,N_5827);
or U6479 (N_6479,N_6227,N_5834);
nor U6480 (N_6480,N_5931,N_5676);
or U6481 (N_6481,N_5795,N_6198);
or U6482 (N_6482,N_5746,N_6128);
nand U6483 (N_6483,N_6093,N_5754);
or U6484 (N_6484,N_6199,N_5640);
xor U6485 (N_6485,N_5728,N_5926);
nor U6486 (N_6486,N_5883,N_5743);
nor U6487 (N_6487,N_5737,N_5968);
nand U6488 (N_6488,N_5778,N_6042);
nand U6489 (N_6489,N_5745,N_5680);
nand U6490 (N_6490,N_5751,N_5636);
nor U6491 (N_6491,N_6115,N_5683);
nor U6492 (N_6492,N_6073,N_5675);
or U6493 (N_6493,N_5951,N_6099);
xor U6494 (N_6494,N_6181,N_5726);
nand U6495 (N_6495,N_6184,N_5966);
xnor U6496 (N_6496,N_6230,N_6215);
xnor U6497 (N_6497,N_5979,N_5953);
or U6498 (N_6498,N_6139,N_6088);
nor U6499 (N_6499,N_5776,N_5693);
and U6500 (N_6500,N_5787,N_6208);
nand U6501 (N_6501,N_5655,N_5964);
or U6502 (N_6502,N_6000,N_6087);
nand U6503 (N_6503,N_5702,N_5824);
nand U6504 (N_6504,N_5768,N_5729);
nor U6505 (N_6505,N_6111,N_5907);
and U6506 (N_6506,N_6125,N_5668);
or U6507 (N_6507,N_5791,N_6023);
xor U6508 (N_6508,N_6097,N_5901);
nor U6509 (N_6509,N_5653,N_6009);
nor U6510 (N_6510,N_6248,N_6126);
nand U6511 (N_6511,N_6022,N_5911);
or U6512 (N_6512,N_5923,N_6109);
nand U6513 (N_6513,N_6091,N_6137);
nand U6514 (N_6514,N_6159,N_6085);
or U6515 (N_6515,N_5663,N_5651);
xor U6516 (N_6516,N_5763,N_6034);
nand U6517 (N_6517,N_5671,N_6032);
nor U6518 (N_6518,N_5767,N_6101);
and U6519 (N_6519,N_6155,N_5832);
nand U6520 (N_6520,N_6015,N_6021);
nor U6521 (N_6521,N_5708,N_5723);
or U6522 (N_6522,N_5949,N_5861);
nand U6523 (N_6523,N_5828,N_5946);
or U6524 (N_6524,N_5727,N_5986);
nor U6525 (N_6525,N_5755,N_5962);
nand U6526 (N_6526,N_6163,N_5809);
xnor U6527 (N_6527,N_5703,N_6206);
and U6528 (N_6528,N_5806,N_5869);
nor U6529 (N_6529,N_6160,N_6078);
xnor U6530 (N_6530,N_6028,N_5948);
and U6531 (N_6531,N_5649,N_5688);
or U6532 (N_6532,N_5935,N_5866);
nor U6533 (N_6533,N_5715,N_6025);
xor U6534 (N_6534,N_5950,N_5752);
or U6535 (N_6535,N_5996,N_6217);
nor U6536 (N_6536,N_6194,N_5720);
and U6537 (N_6537,N_5674,N_6050);
or U6538 (N_6538,N_5881,N_6041);
nand U6539 (N_6539,N_5759,N_6149);
nor U6540 (N_6540,N_6146,N_6114);
or U6541 (N_6541,N_5958,N_5781);
and U6542 (N_6542,N_5670,N_5793);
xnor U6543 (N_6543,N_5750,N_6061);
nand U6544 (N_6544,N_5912,N_6141);
xor U6545 (N_6545,N_6135,N_6247);
nand U6546 (N_6546,N_5770,N_5984);
nor U6547 (N_6547,N_6197,N_6095);
xor U6548 (N_6548,N_5982,N_6192);
nand U6549 (N_6549,N_6094,N_6077);
and U6550 (N_6550,N_6144,N_6092);
xor U6551 (N_6551,N_6106,N_5992);
or U6552 (N_6552,N_5803,N_6108);
and U6553 (N_6553,N_6142,N_5784);
or U6554 (N_6554,N_5820,N_6180);
or U6555 (N_6555,N_6020,N_5903);
or U6556 (N_6556,N_5691,N_5944);
or U6557 (N_6557,N_6062,N_5736);
and U6558 (N_6558,N_5879,N_5956);
xor U6559 (N_6559,N_5847,N_5783);
nor U6560 (N_6560,N_5998,N_6121);
xor U6561 (N_6561,N_5909,N_5925);
xnor U6562 (N_6562,N_5899,N_6240);
or U6563 (N_6563,N_5945,N_5835);
nor U6564 (N_6564,N_6053,N_5829);
xnor U6565 (N_6565,N_5693,N_6222);
xor U6566 (N_6566,N_5794,N_5649);
nand U6567 (N_6567,N_6154,N_6007);
or U6568 (N_6568,N_5753,N_5742);
nand U6569 (N_6569,N_5947,N_5972);
nor U6570 (N_6570,N_6111,N_5909);
nand U6571 (N_6571,N_6213,N_6214);
or U6572 (N_6572,N_5717,N_5814);
or U6573 (N_6573,N_6190,N_6231);
or U6574 (N_6574,N_6138,N_6139);
nor U6575 (N_6575,N_5956,N_5804);
xor U6576 (N_6576,N_5883,N_6032);
xor U6577 (N_6577,N_5831,N_5752);
nand U6578 (N_6578,N_5951,N_5727);
and U6579 (N_6579,N_6206,N_5757);
or U6580 (N_6580,N_5659,N_5799);
xor U6581 (N_6581,N_5786,N_6166);
nor U6582 (N_6582,N_5748,N_6102);
nand U6583 (N_6583,N_6233,N_6075);
and U6584 (N_6584,N_5975,N_6075);
nor U6585 (N_6585,N_5670,N_6242);
and U6586 (N_6586,N_5957,N_5839);
or U6587 (N_6587,N_5856,N_6000);
xnor U6588 (N_6588,N_5974,N_5626);
and U6589 (N_6589,N_6184,N_5815);
and U6590 (N_6590,N_5957,N_5772);
or U6591 (N_6591,N_6185,N_5798);
xor U6592 (N_6592,N_5629,N_6023);
and U6593 (N_6593,N_6027,N_6057);
nand U6594 (N_6594,N_6145,N_5647);
and U6595 (N_6595,N_5992,N_5840);
and U6596 (N_6596,N_5976,N_6023);
and U6597 (N_6597,N_6090,N_5872);
xor U6598 (N_6598,N_6231,N_5731);
nand U6599 (N_6599,N_5944,N_6235);
nor U6600 (N_6600,N_5727,N_6088);
nand U6601 (N_6601,N_5745,N_5888);
nor U6602 (N_6602,N_6113,N_6114);
xnor U6603 (N_6603,N_6247,N_6114);
xor U6604 (N_6604,N_5705,N_5998);
or U6605 (N_6605,N_6198,N_5813);
or U6606 (N_6606,N_6126,N_6104);
nor U6607 (N_6607,N_5861,N_6184);
xor U6608 (N_6608,N_5969,N_5650);
or U6609 (N_6609,N_5801,N_6237);
and U6610 (N_6610,N_5800,N_6126);
and U6611 (N_6611,N_6177,N_5730);
xor U6612 (N_6612,N_5933,N_6184);
nor U6613 (N_6613,N_5728,N_6210);
or U6614 (N_6614,N_5713,N_6132);
and U6615 (N_6615,N_6181,N_6171);
nor U6616 (N_6616,N_5986,N_5817);
nor U6617 (N_6617,N_5758,N_5779);
nor U6618 (N_6618,N_5816,N_6111);
nand U6619 (N_6619,N_5946,N_5907);
and U6620 (N_6620,N_6196,N_5694);
xor U6621 (N_6621,N_6072,N_5746);
nand U6622 (N_6622,N_6114,N_6079);
and U6623 (N_6623,N_5877,N_6246);
and U6624 (N_6624,N_5958,N_5996);
or U6625 (N_6625,N_6077,N_5808);
nand U6626 (N_6626,N_5852,N_6152);
nor U6627 (N_6627,N_5689,N_6113);
xor U6628 (N_6628,N_5961,N_5700);
nor U6629 (N_6629,N_6228,N_5749);
nor U6630 (N_6630,N_6220,N_6246);
and U6631 (N_6631,N_6041,N_5947);
nor U6632 (N_6632,N_5700,N_5712);
nor U6633 (N_6633,N_5963,N_6030);
xnor U6634 (N_6634,N_6042,N_5912);
nand U6635 (N_6635,N_5946,N_5668);
xnor U6636 (N_6636,N_6115,N_5953);
nand U6637 (N_6637,N_5893,N_6128);
xor U6638 (N_6638,N_5656,N_6102);
and U6639 (N_6639,N_5727,N_6163);
nand U6640 (N_6640,N_6153,N_5944);
nor U6641 (N_6641,N_5765,N_5961);
xor U6642 (N_6642,N_5786,N_5773);
xnor U6643 (N_6643,N_5980,N_5796);
xnor U6644 (N_6644,N_6105,N_6056);
or U6645 (N_6645,N_5640,N_6001);
nor U6646 (N_6646,N_5962,N_5977);
xnor U6647 (N_6647,N_5941,N_5714);
or U6648 (N_6648,N_6178,N_5996);
nor U6649 (N_6649,N_5935,N_5709);
nand U6650 (N_6650,N_6083,N_5835);
xnor U6651 (N_6651,N_5781,N_6225);
xnor U6652 (N_6652,N_5709,N_6042);
and U6653 (N_6653,N_5701,N_6170);
or U6654 (N_6654,N_6116,N_5803);
and U6655 (N_6655,N_5661,N_5748);
or U6656 (N_6656,N_5781,N_5850);
and U6657 (N_6657,N_5633,N_5809);
and U6658 (N_6658,N_5915,N_5767);
nor U6659 (N_6659,N_6052,N_5705);
and U6660 (N_6660,N_6019,N_5969);
nand U6661 (N_6661,N_6221,N_5842);
nor U6662 (N_6662,N_6148,N_6103);
nor U6663 (N_6663,N_5876,N_6069);
and U6664 (N_6664,N_6018,N_5643);
nor U6665 (N_6665,N_5971,N_6109);
and U6666 (N_6666,N_5806,N_5688);
or U6667 (N_6667,N_6178,N_6216);
or U6668 (N_6668,N_6193,N_5992);
nor U6669 (N_6669,N_6029,N_6097);
or U6670 (N_6670,N_5694,N_5781);
nor U6671 (N_6671,N_5861,N_5826);
nand U6672 (N_6672,N_6018,N_5960);
and U6673 (N_6673,N_5642,N_5941);
nand U6674 (N_6674,N_5808,N_5741);
nor U6675 (N_6675,N_6091,N_5747);
nand U6676 (N_6676,N_5713,N_5872);
xor U6677 (N_6677,N_5950,N_5969);
xnor U6678 (N_6678,N_6100,N_6176);
nand U6679 (N_6679,N_5628,N_5960);
nand U6680 (N_6680,N_5700,N_5807);
xnor U6681 (N_6681,N_6173,N_6079);
nor U6682 (N_6682,N_5685,N_6012);
nor U6683 (N_6683,N_5715,N_6038);
or U6684 (N_6684,N_6092,N_5965);
xnor U6685 (N_6685,N_5879,N_5932);
and U6686 (N_6686,N_5761,N_6089);
xnor U6687 (N_6687,N_5843,N_6229);
and U6688 (N_6688,N_6206,N_6212);
or U6689 (N_6689,N_5897,N_5980);
or U6690 (N_6690,N_5954,N_6165);
xor U6691 (N_6691,N_5831,N_5882);
and U6692 (N_6692,N_6141,N_5958);
nor U6693 (N_6693,N_5630,N_6094);
or U6694 (N_6694,N_5763,N_6029);
or U6695 (N_6695,N_5741,N_5651);
nand U6696 (N_6696,N_5696,N_5828);
nand U6697 (N_6697,N_5745,N_6084);
and U6698 (N_6698,N_6061,N_6126);
and U6699 (N_6699,N_5757,N_5676);
or U6700 (N_6700,N_6126,N_5962);
nand U6701 (N_6701,N_5654,N_5842);
xor U6702 (N_6702,N_6119,N_5859);
nand U6703 (N_6703,N_5813,N_5815);
xor U6704 (N_6704,N_5952,N_5751);
nor U6705 (N_6705,N_6178,N_5798);
nand U6706 (N_6706,N_5668,N_5884);
or U6707 (N_6707,N_6179,N_5943);
or U6708 (N_6708,N_6169,N_5627);
or U6709 (N_6709,N_5734,N_5745);
or U6710 (N_6710,N_6012,N_5729);
nand U6711 (N_6711,N_5844,N_6072);
nor U6712 (N_6712,N_6112,N_6139);
xor U6713 (N_6713,N_6194,N_5981);
nor U6714 (N_6714,N_6076,N_5809);
nand U6715 (N_6715,N_5702,N_5629);
nor U6716 (N_6716,N_6055,N_5699);
or U6717 (N_6717,N_6223,N_6226);
or U6718 (N_6718,N_6222,N_5789);
and U6719 (N_6719,N_5819,N_5814);
nor U6720 (N_6720,N_5656,N_5635);
and U6721 (N_6721,N_5967,N_5795);
and U6722 (N_6722,N_5691,N_6101);
or U6723 (N_6723,N_5987,N_5977);
and U6724 (N_6724,N_6244,N_6115);
and U6725 (N_6725,N_5703,N_5725);
nand U6726 (N_6726,N_5958,N_5811);
xnor U6727 (N_6727,N_6190,N_5899);
or U6728 (N_6728,N_5980,N_6009);
nand U6729 (N_6729,N_6078,N_6231);
nand U6730 (N_6730,N_5641,N_5661);
nand U6731 (N_6731,N_6008,N_6209);
xnor U6732 (N_6732,N_6005,N_6092);
nand U6733 (N_6733,N_5896,N_5851);
nor U6734 (N_6734,N_5838,N_6193);
or U6735 (N_6735,N_6114,N_6043);
and U6736 (N_6736,N_6186,N_5673);
nor U6737 (N_6737,N_6159,N_5700);
or U6738 (N_6738,N_5832,N_5970);
nand U6739 (N_6739,N_5783,N_5792);
nand U6740 (N_6740,N_6217,N_5697);
xnor U6741 (N_6741,N_5790,N_6129);
or U6742 (N_6742,N_6199,N_6105);
nand U6743 (N_6743,N_6124,N_6217);
xnor U6744 (N_6744,N_5746,N_5977);
or U6745 (N_6745,N_5723,N_5775);
xor U6746 (N_6746,N_5773,N_5951);
or U6747 (N_6747,N_5938,N_5660);
or U6748 (N_6748,N_5642,N_5745);
xnor U6749 (N_6749,N_5818,N_5896);
nor U6750 (N_6750,N_6005,N_5778);
nor U6751 (N_6751,N_5802,N_5805);
nor U6752 (N_6752,N_6159,N_6183);
and U6753 (N_6753,N_5756,N_6119);
and U6754 (N_6754,N_5985,N_6148);
nor U6755 (N_6755,N_6096,N_5690);
nand U6756 (N_6756,N_6172,N_6195);
nand U6757 (N_6757,N_5804,N_6208);
nor U6758 (N_6758,N_5625,N_6082);
xnor U6759 (N_6759,N_5875,N_5873);
and U6760 (N_6760,N_5819,N_6154);
nor U6761 (N_6761,N_5959,N_6219);
xnor U6762 (N_6762,N_5845,N_5945);
or U6763 (N_6763,N_5634,N_5657);
nor U6764 (N_6764,N_6128,N_5913);
nand U6765 (N_6765,N_5706,N_5971);
nor U6766 (N_6766,N_5836,N_6228);
nor U6767 (N_6767,N_5798,N_5809);
nor U6768 (N_6768,N_5877,N_5959);
and U6769 (N_6769,N_5797,N_5631);
xnor U6770 (N_6770,N_5951,N_6182);
nand U6771 (N_6771,N_6080,N_5883);
nor U6772 (N_6772,N_5727,N_6012);
or U6773 (N_6773,N_6198,N_5767);
nor U6774 (N_6774,N_5721,N_5665);
and U6775 (N_6775,N_6237,N_5650);
and U6776 (N_6776,N_5706,N_6155);
or U6777 (N_6777,N_5931,N_5705);
xnor U6778 (N_6778,N_6005,N_5636);
nand U6779 (N_6779,N_6079,N_5800);
xor U6780 (N_6780,N_6240,N_6051);
xor U6781 (N_6781,N_5717,N_6008);
nand U6782 (N_6782,N_6249,N_6024);
nand U6783 (N_6783,N_6194,N_5685);
or U6784 (N_6784,N_5767,N_5740);
and U6785 (N_6785,N_6243,N_5972);
xnor U6786 (N_6786,N_5740,N_6130);
nand U6787 (N_6787,N_5847,N_6118);
nor U6788 (N_6788,N_6247,N_5833);
xnor U6789 (N_6789,N_6232,N_5812);
or U6790 (N_6790,N_6078,N_5974);
nor U6791 (N_6791,N_5645,N_6168);
xnor U6792 (N_6792,N_5858,N_5698);
nand U6793 (N_6793,N_6070,N_5829);
and U6794 (N_6794,N_5636,N_5906);
xnor U6795 (N_6795,N_6012,N_5962);
and U6796 (N_6796,N_5823,N_6110);
or U6797 (N_6797,N_5980,N_6069);
or U6798 (N_6798,N_5630,N_5982);
xor U6799 (N_6799,N_6217,N_5656);
nand U6800 (N_6800,N_5957,N_6221);
and U6801 (N_6801,N_5952,N_6122);
nor U6802 (N_6802,N_6120,N_6248);
nand U6803 (N_6803,N_6008,N_5712);
nor U6804 (N_6804,N_5951,N_6177);
nand U6805 (N_6805,N_6176,N_5783);
or U6806 (N_6806,N_6159,N_5688);
xnor U6807 (N_6807,N_5839,N_5767);
nor U6808 (N_6808,N_6009,N_5783);
and U6809 (N_6809,N_5833,N_6173);
and U6810 (N_6810,N_6009,N_5734);
xnor U6811 (N_6811,N_5681,N_5947);
or U6812 (N_6812,N_5697,N_5779);
xnor U6813 (N_6813,N_5885,N_5741);
nor U6814 (N_6814,N_6146,N_6231);
or U6815 (N_6815,N_6106,N_5950);
nor U6816 (N_6816,N_6134,N_5727);
nor U6817 (N_6817,N_6053,N_5648);
and U6818 (N_6818,N_6150,N_5840);
and U6819 (N_6819,N_5677,N_5744);
nand U6820 (N_6820,N_6193,N_5756);
xnor U6821 (N_6821,N_6217,N_5750);
and U6822 (N_6822,N_5783,N_6061);
nand U6823 (N_6823,N_6141,N_5790);
and U6824 (N_6824,N_5941,N_5853);
xnor U6825 (N_6825,N_6160,N_6102);
xor U6826 (N_6826,N_5914,N_5679);
and U6827 (N_6827,N_5776,N_5985);
nand U6828 (N_6828,N_6212,N_6138);
nor U6829 (N_6829,N_6029,N_5784);
xor U6830 (N_6830,N_5965,N_5952);
xnor U6831 (N_6831,N_5676,N_6150);
nand U6832 (N_6832,N_5859,N_5719);
xnor U6833 (N_6833,N_5913,N_5921);
nand U6834 (N_6834,N_5643,N_6109);
nor U6835 (N_6835,N_5729,N_5693);
or U6836 (N_6836,N_6008,N_5802);
xor U6837 (N_6837,N_5907,N_5625);
and U6838 (N_6838,N_5985,N_6222);
nand U6839 (N_6839,N_5785,N_5689);
nor U6840 (N_6840,N_6230,N_6161);
nor U6841 (N_6841,N_5879,N_5819);
and U6842 (N_6842,N_5911,N_6184);
or U6843 (N_6843,N_6018,N_6072);
nor U6844 (N_6844,N_6183,N_6127);
nand U6845 (N_6845,N_5964,N_5759);
nand U6846 (N_6846,N_5928,N_5979);
nor U6847 (N_6847,N_6044,N_5829);
or U6848 (N_6848,N_5883,N_5965);
nor U6849 (N_6849,N_6172,N_5705);
nor U6850 (N_6850,N_6228,N_5894);
nor U6851 (N_6851,N_5727,N_6239);
xnor U6852 (N_6852,N_5875,N_5769);
and U6853 (N_6853,N_6141,N_5990);
and U6854 (N_6854,N_5695,N_6000);
and U6855 (N_6855,N_5875,N_6063);
or U6856 (N_6856,N_6109,N_6225);
nand U6857 (N_6857,N_6236,N_6244);
and U6858 (N_6858,N_5965,N_5798);
and U6859 (N_6859,N_5985,N_5850);
and U6860 (N_6860,N_5870,N_6042);
or U6861 (N_6861,N_5650,N_5938);
or U6862 (N_6862,N_5794,N_5643);
nor U6863 (N_6863,N_5645,N_5677);
and U6864 (N_6864,N_5658,N_5771);
nor U6865 (N_6865,N_6233,N_5930);
xor U6866 (N_6866,N_6224,N_5964);
xnor U6867 (N_6867,N_6235,N_5740);
nor U6868 (N_6868,N_5740,N_6087);
xnor U6869 (N_6869,N_6228,N_6154);
nor U6870 (N_6870,N_5981,N_6125);
nand U6871 (N_6871,N_5861,N_6170);
nor U6872 (N_6872,N_6149,N_6116);
xor U6873 (N_6873,N_5811,N_5653);
xor U6874 (N_6874,N_6155,N_6063);
nand U6875 (N_6875,N_6855,N_6543);
xor U6876 (N_6876,N_6685,N_6724);
nor U6877 (N_6877,N_6250,N_6824);
and U6878 (N_6878,N_6415,N_6421);
nand U6879 (N_6879,N_6255,N_6683);
nand U6880 (N_6880,N_6578,N_6536);
xnor U6881 (N_6881,N_6258,N_6831);
and U6882 (N_6882,N_6570,N_6350);
and U6883 (N_6883,N_6299,N_6719);
nand U6884 (N_6884,N_6443,N_6615);
xnor U6885 (N_6885,N_6655,N_6446);
nor U6886 (N_6886,N_6846,N_6254);
xor U6887 (N_6887,N_6376,N_6865);
nor U6888 (N_6888,N_6342,N_6505);
xor U6889 (N_6889,N_6745,N_6352);
xor U6890 (N_6890,N_6348,N_6811);
nor U6891 (N_6891,N_6436,N_6432);
nand U6892 (N_6892,N_6413,N_6703);
or U6893 (N_6893,N_6334,N_6288);
or U6894 (N_6894,N_6868,N_6861);
or U6895 (N_6895,N_6765,N_6409);
xor U6896 (N_6896,N_6704,N_6457);
or U6897 (N_6897,N_6266,N_6656);
nand U6898 (N_6898,N_6662,N_6616);
xor U6899 (N_6899,N_6510,N_6571);
xor U6900 (N_6900,N_6291,N_6315);
nor U6901 (N_6901,N_6509,N_6261);
and U6902 (N_6902,N_6821,N_6489);
and U6903 (N_6903,N_6274,N_6406);
or U6904 (N_6904,N_6838,N_6650);
and U6905 (N_6905,N_6462,N_6608);
nand U6906 (N_6906,N_6337,N_6309);
nand U6907 (N_6907,N_6641,N_6279);
and U6908 (N_6908,N_6374,N_6734);
nand U6909 (N_6909,N_6872,N_6874);
nor U6910 (N_6910,N_6711,N_6358);
nor U6911 (N_6911,N_6722,N_6568);
nand U6912 (N_6912,N_6466,N_6714);
nor U6913 (N_6913,N_6682,N_6325);
nor U6914 (N_6914,N_6692,N_6272);
nand U6915 (N_6915,N_6486,N_6481);
or U6916 (N_6916,N_6773,N_6527);
xor U6917 (N_6917,N_6648,N_6638);
nor U6918 (N_6918,N_6524,N_6857);
xnor U6919 (N_6919,N_6252,N_6414);
nand U6920 (N_6920,N_6517,N_6806);
nor U6921 (N_6921,N_6307,N_6465);
and U6922 (N_6922,N_6265,N_6329);
or U6923 (N_6923,N_6424,N_6444);
nand U6924 (N_6924,N_6754,N_6269);
xor U6925 (N_6925,N_6384,N_6845);
or U6926 (N_6926,N_6805,N_6675);
xnor U6927 (N_6927,N_6774,N_6270);
xor U6928 (N_6928,N_6796,N_6725);
and U6929 (N_6929,N_6530,N_6470);
and U6930 (N_6930,N_6706,N_6364);
or U6931 (N_6931,N_6775,N_6686);
xor U6932 (N_6932,N_6324,N_6472);
and U6933 (N_6933,N_6800,N_6469);
nand U6934 (N_6934,N_6825,N_6416);
nand U6935 (N_6935,N_6295,N_6437);
nand U6936 (N_6936,N_6627,N_6873);
xor U6937 (N_6937,N_6684,N_6625);
or U6938 (N_6938,N_6849,N_6493);
nor U6939 (N_6939,N_6271,N_6532);
xor U6940 (N_6940,N_6689,N_6296);
and U6941 (N_6941,N_6643,N_6582);
nor U6942 (N_6942,N_6764,N_6757);
nor U6943 (N_6943,N_6665,N_6856);
nor U6944 (N_6944,N_6626,N_6817);
and U6945 (N_6945,N_6508,N_6426);
xnor U6946 (N_6946,N_6435,N_6769);
nand U6947 (N_6947,N_6564,N_6450);
nor U6948 (N_6948,N_6736,N_6577);
or U6949 (N_6949,N_6488,N_6726);
nand U6950 (N_6950,N_6776,N_6807);
or U6951 (N_6951,N_6506,N_6397);
nor U6952 (N_6952,N_6283,N_6474);
nor U6953 (N_6953,N_6460,N_6318);
nand U6954 (N_6954,N_6576,N_6447);
and U6955 (N_6955,N_6546,N_6672);
or U6956 (N_6956,N_6553,N_6671);
xor U6957 (N_6957,N_6306,N_6669);
nor U6958 (N_6958,N_6287,N_6778);
nor U6959 (N_6959,N_6630,N_6268);
nand U6960 (N_6960,N_6727,N_6293);
xor U6961 (N_6961,N_6308,N_6585);
nand U6962 (N_6962,N_6870,N_6741);
and U6963 (N_6963,N_6407,N_6558);
and U6964 (N_6964,N_6368,N_6834);
xor U6965 (N_6965,N_6353,N_6783);
nor U6966 (N_6966,N_6850,N_6814);
and U6967 (N_6967,N_6526,N_6499);
nor U6968 (N_6968,N_6747,N_6439);
nor U6969 (N_6969,N_6702,N_6781);
nor U6970 (N_6970,N_6761,N_6289);
nor U6971 (N_6971,N_6750,N_6634);
or U6972 (N_6972,N_6476,N_6678);
and U6973 (N_6973,N_6590,N_6664);
and U6974 (N_6974,N_6323,N_6471);
and U6975 (N_6975,N_6535,N_6452);
and U6976 (N_6976,N_6304,N_6561);
and U6977 (N_6977,N_6605,N_6848);
nor U6978 (N_6978,N_6322,N_6297);
xor U6979 (N_6979,N_6592,N_6673);
or U6980 (N_6980,N_6319,N_6565);
nand U6981 (N_6981,N_6789,N_6496);
nor U6982 (N_6982,N_6441,N_6812);
and U6983 (N_6983,N_6534,N_6300);
or U6984 (N_6984,N_6263,N_6431);
nand U6985 (N_6985,N_6760,N_6584);
and U6986 (N_6986,N_6273,N_6646);
or U6987 (N_6987,N_6813,N_6835);
nor U6988 (N_6988,N_6539,N_6393);
xor U6989 (N_6989,N_6310,N_6455);
nor U6990 (N_6990,N_6713,N_6645);
and U6991 (N_6991,N_6788,N_6339);
nand U6992 (N_6992,N_6867,N_6573);
or U6993 (N_6993,N_6380,N_6687);
or U6994 (N_6994,N_6385,N_6448);
xnor U6995 (N_6995,N_6787,N_6328);
nor U6996 (N_6996,N_6779,N_6858);
nand U6997 (N_6997,N_6823,N_6483);
or U6998 (N_6998,N_6541,N_6494);
and U6999 (N_6999,N_6631,N_6808);
xor U7000 (N_7000,N_6795,N_6251);
or U7001 (N_7001,N_6351,N_6567);
and U7002 (N_7002,N_6402,N_6338);
nand U7003 (N_7003,N_6737,N_6609);
xor U7004 (N_7004,N_6302,N_6696);
xnor U7005 (N_7005,N_6679,N_6259);
nand U7006 (N_7006,N_6497,N_6349);
or U7007 (N_7007,N_6286,N_6516);
and U7008 (N_7008,N_6639,N_6528);
nor U7009 (N_7009,N_6600,N_6738);
xnor U7010 (N_7010,N_6604,N_6749);
or U7011 (N_7011,N_6670,N_6451);
xnor U7012 (N_7012,N_6477,N_6359);
and U7013 (N_7013,N_6365,N_6828);
nand U7014 (N_7014,N_6552,N_6700);
nor U7015 (N_7015,N_6491,N_6453);
xnor U7016 (N_7016,N_6635,N_6336);
or U7017 (N_7017,N_6820,N_6705);
and U7018 (N_7018,N_6390,N_6716);
and U7019 (N_7019,N_6332,N_6628);
or U7020 (N_7020,N_6559,N_6490);
and U7021 (N_7021,N_6378,N_6511);
or U7022 (N_7022,N_6373,N_6624);
xor U7023 (N_7023,N_6657,N_6369);
or U7024 (N_7024,N_6709,N_6386);
and U7025 (N_7025,N_6518,N_6396);
xnor U7026 (N_7026,N_6556,N_6440);
nor U7027 (N_7027,N_6575,N_6545);
xor U7028 (N_7028,N_6740,N_6382);
and U7029 (N_7029,N_6732,N_6801);
xor U7030 (N_7030,N_6459,N_6581);
nand U7031 (N_7031,N_6859,N_6537);
nand U7032 (N_7032,N_6548,N_6377);
nand U7033 (N_7033,N_6412,N_6791);
or U7034 (N_7034,N_6341,N_6723);
or U7035 (N_7035,N_6305,N_6357);
or U7036 (N_7036,N_6387,N_6809);
or U7037 (N_7037,N_6544,N_6837);
xor U7038 (N_7038,N_6829,N_6320);
nor U7039 (N_7039,N_6601,N_6843);
xnor U7040 (N_7040,N_6479,N_6542);
nor U7041 (N_7041,N_6599,N_6697);
nand U7042 (N_7042,N_6758,N_6613);
xor U7043 (N_7043,N_6316,N_6693);
nand U7044 (N_7044,N_6840,N_6822);
and U7045 (N_7045,N_6422,N_6411);
xor U7046 (N_7046,N_6547,N_6851);
and U7047 (N_7047,N_6473,N_6563);
and U7048 (N_7048,N_6560,N_6404);
nor U7049 (N_7049,N_6520,N_6438);
nand U7050 (N_7050,N_6854,N_6772);
nand U7051 (N_7051,N_6294,N_6449);
and U7052 (N_7052,N_6344,N_6588);
nand U7053 (N_7053,N_6549,N_6718);
nand U7054 (N_7054,N_6862,N_6731);
and U7055 (N_7055,N_6580,N_6652);
or U7056 (N_7056,N_6832,N_6729);
nand U7057 (N_7057,N_6504,N_6456);
and U7058 (N_7058,N_6793,N_6503);
nor U7059 (N_7059,N_6383,N_6852);
nor U7060 (N_7060,N_6802,N_6589);
or U7061 (N_7061,N_6388,N_6744);
nand U7062 (N_7062,N_6792,N_6445);
xnor U7063 (N_7063,N_6400,N_6429);
xor U7064 (N_7064,N_6555,N_6391);
xnor U7065 (N_7065,N_6654,N_6554);
nand U7066 (N_7066,N_6428,N_6816);
nor U7067 (N_7067,N_6830,N_6701);
nand U7068 (N_7068,N_6484,N_6661);
xnor U7069 (N_7069,N_6458,N_6253);
nor U7070 (N_7070,N_6644,N_6658);
xnor U7071 (N_7071,N_6607,N_6743);
nand U7072 (N_7072,N_6410,N_6755);
xor U7073 (N_7073,N_6538,N_6695);
nor U7074 (N_7074,N_6540,N_6420);
xnor U7075 (N_7075,N_6612,N_6777);
and U7076 (N_7076,N_6770,N_6333);
or U7077 (N_7077,N_6482,N_6620);
nand U7078 (N_7078,N_6264,N_6844);
xnor U7079 (N_7079,N_6756,N_6434);
xor U7080 (N_7080,N_6794,N_6401);
and U7081 (N_7081,N_6529,N_6298);
nand U7082 (N_7082,N_6767,N_6395);
nor U7083 (N_7083,N_6636,N_6677);
nand U7084 (N_7084,N_6523,N_6694);
or U7085 (N_7085,N_6804,N_6690);
xnor U7086 (N_7086,N_6321,N_6871);
nand U7087 (N_7087,N_6782,N_6798);
xnor U7088 (N_7088,N_6810,N_6853);
and U7089 (N_7089,N_6784,N_6464);
nand U7090 (N_7090,N_6591,N_6715);
nor U7091 (N_7091,N_6361,N_6282);
or U7092 (N_7092,N_6863,N_6717);
nor U7093 (N_7093,N_6721,N_6403);
xor U7094 (N_7094,N_6587,N_6733);
nor U7095 (N_7095,N_6619,N_6399);
nand U7096 (N_7096,N_6500,N_6864);
nor U7097 (N_7097,N_6623,N_6467);
xor U7098 (N_7098,N_6818,N_6819);
xor U7099 (N_7099,N_6618,N_6728);
or U7100 (N_7100,N_6340,N_6317);
and U7101 (N_7101,N_6640,N_6839);
xnor U7102 (N_7102,N_6280,N_6290);
nand U7103 (N_7103,N_6311,N_6372);
and U7104 (N_7104,N_6492,N_6389);
nand U7105 (N_7105,N_6674,N_6551);
and U7106 (N_7106,N_6487,N_6468);
xor U7107 (N_7107,N_6593,N_6771);
nand U7108 (N_7108,N_6423,N_6768);
or U7109 (N_7109,N_6569,N_6292);
nor U7110 (N_7110,N_6327,N_6419);
or U7111 (N_7111,N_6262,N_6507);
and U7112 (N_7112,N_6680,N_6501);
and U7113 (N_7113,N_6281,N_6394);
nor U7114 (N_7114,N_6427,N_6277);
xor U7115 (N_7115,N_6346,N_6276);
xnor U7116 (N_7116,N_6785,N_6356);
xnor U7117 (N_7117,N_6417,N_6360);
and U7118 (N_7118,N_6405,N_6475);
xor U7119 (N_7119,N_6660,N_6594);
nand U7120 (N_7120,N_6659,N_6596);
and U7121 (N_7121,N_6710,N_6312);
and U7122 (N_7122,N_6866,N_6256);
xor U7123 (N_7123,N_6614,N_6275);
and U7124 (N_7124,N_6666,N_6786);
nor U7125 (N_7125,N_6514,N_6533);
xnor U7126 (N_7126,N_6301,N_6257);
nor U7127 (N_7127,N_6478,N_6566);
xor U7128 (N_7128,N_6367,N_6842);
or U7129 (N_7129,N_6803,N_6330);
or U7130 (N_7130,N_6285,N_6629);
xnor U7131 (N_7131,N_6495,N_6681);
nor U7132 (N_7132,N_6699,N_6498);
nor U7133 (N_7133,N_6314,N_6597);
and U7134 (N_7134,N_6739,N_6512);
and U7135 (N_7135,N_6335,N_6833);
and U7136 (N_7136,N_6611,N_6519);
and U7137 (N_7137,N_6622,N_6521);
or U7138 (N_7138,N_6347,N_6430);
or U7139 (N_7139,N_6485,N_6780);
xor U7140 (N_7140,N_6762,N_6730);
or U7141 (N_7141,N_6642,N_6433);
or U7142 (N_7142,N_6392,N_6284);
nand U7143 (N_7143,N_6647,N_6610);
xor U7144 (N_7144,N_6637,N_6550);
nor U7145 (N_7145,N_6326,N_6751);
and U7146 (N_7146,N_6363,N_6742);
nand U7147 (N_7147,N_6408,N_6278);
and U7148 (N_7148,N_6797,N_6841);
nor U7149 (N_7149,N_6463,N_6746);
and U7150 (N_7150,N_6418,N_6720);
nand U7151 (N_7151,N_6708,N_6748);
nor U7152 (N_7152,N_6502,N_6525);
nand U7153 (N_7153,N_6260,N_6354);
xor U7154 (N_7154,N_6815,N_6375);
nor U7155 (N_7155,N_6370,N_6313);
or U7156 (N_7156,N_6676,N_6602);
or U7157 (N_7157,N_6454,N_6766);
or U7158 (N_7158,N_6371,N_6598);
xnor U7159 (N_7159,N_6869,N_6759);
nand U7160 (N_7160,N_6595,N_6653);
xor U7161 (N_7161,N_6586,N_6617);
xor U7162 (N_7162,N_6621,N_6799);
or U7163 (N_7163,N_6633,N_6267);
or U7164 (N_7164,N_6827,N_6847);
and U7165 (N_7165,N_6442,N_6355);
nand U7166 (N_7166,N_6632,N_6398);
xnor U7167 (N_7167,N_6515,N_6860);
and U7168 (N_7168,N_6763,N_6688);
xnor U7169 (N_7169,N_6522,N_6707);
xnor U7170 (N_7170,N_6480,N_6362);
and U7171 (N_7171,N_6667,N_6331);
or U7172 (N_7172,N_6691,N_6379);
nor U7173 (N_7173,N_6698,N_6649);
or U7174 (N_7174,N_6557,N_6712);
xnor U7175 (N_7175,N_6381,N_6836);
nor U7176 (N_7176,N_6425,N_6663);
nand U7177 (N_7177,N_6790,N_6735);
xor U7178 (N_7178,N_6572,N_6752);
nor U7179 (N_7179,N_6579,N_6562);
or U7180 (N_7180,N_6606,N_6366);
nor U7181 (N_7181,N_6753,N_6583);
nor U7182 (N_7182,N_6651,N_6668);
or U7183 (N_7183,N_6531,N_6603);
nor U7184 (N_7184,N_6345,N_6513);
and U7185 (N_7185,N_6303,N_6826);
and U7186 (N_7186,N_6574,N_6461);
or U7187 (N_7187,N_6343,N_6522);
nor U7188 (N_7188,N_6829,N_6716);
nor U7189 (N_7189,N_6306,N_6398);
nor U7190 (N_7190,N_6386,N_6392);
nand U7191 (N_7191,N_6509,N_6633);
and U7192 (N_7192,N_6315,N_6771);
nor U7193 (N_7193,N_6700,N_6771);
or U7194 (N_7194,N_6609,N_6773);
nor U7195 (N_7195,N_6719,N_6717);
and U7196 (N_7196,N_6381,N_6804);
or U7197 (N_7197,N_6870,N_6653);
xnor U7198 (N_7198,N_6375,N_6607);
xor U7199 (N_7199,N_6699,N_6345);
nor U7200 (N_7200,N_6376,N_6517);
or U7201 (N_7201,N_6467,N_6651);
and U7202 (N_7202,N_6805,N_6466);
nand U7203 (N_7203,N_6587,N_6779);
or U7204 (N_7204,N_6369,N_6277);
or U7205 (N_7205,N_6284,N_6665);
nand U7206 (N_7206,N_6675,N_6511);
nor U7207 (N_7207,N_6553,N_6741);
xnor U7208 (N_7208,N_6416,N_6271);
nand U7209 (N_7209,N_6565,N_6251);
xnor U7210 (N_7210,N_6639,N_6771);
or U7211 (N_7211,N_6362,N_6409);
and U7212 (N_7212,N_6453,N_6763);
nor U7213 (N_7213,N_6672,N_6477);
or U7214 (N_7214,N_6869,N_6781);
and U7215 (N_7215,N_6709,N_6606);
nand U7216 (N_7216,N_6820,N_6670);
and U7217 (N_7217,N_6865,N_6351);
nand U7218 (N_7218,N_6780,N_6379);
and U7219 (N_7219,N_6696,N_6844);
nor U7220 (N_7220,N_6275,N_6674);
nor U7221 (N_7221,N_6828,N_6664);
nor U7222 (N_7222,N_6795,N_6637);
nor U7223 (N_7223,N_6734,N_6674);
nor U7224 (N_7224,N_6541,N_6348);
or U7225 (N_7225,N_6258,N_6480);
or U7226 (N_7226,N_6452,N_6313);
nor U7227 (N_7227,N_6519,N_6278);
nor U7228 (N_7228,N_6326,N_6504);
and U7229 (N_7229,N_6283,N_6824);
or U7230 (N_7230,N_6373,N_6819);
nand U7231 (N_7231,N_6774,N_6718);
or U7232 (N_7232,N_6857,N_6321);
and U7233 (N_7233,N_6491,N_6342);
or U7234 (N_7234,N_6508,N_6481);
and U7235 (N_7235,N_6506,N_6574);
xnor U7236 (N_7236,N_6387,N_6547);
xor U7237 (N_7237,N_6778,N_6458);
xor U7238 (N_7238,N_6535,N_6338);
xor U7239 (N_7239,N_6738,N_6439);
nand U7240 (N_7240,N_6370,N_6365);
nand U7241 (N_7241,N_6361,N_6733);
or U7242 (N_7242,N_6535,N_6505);
and U7243 (N_7243,N_6799,N_6841);
nand U7244 (N_7244,N_6521,N_6658);
or U7245 (N_7245,N_6597,N_6251);
nand U7246 (N_7246,N_6673,N_6419);
nand U7247 (N_7247,N_6691,N_6865);
or U7248 (N_7248,N_6573,N_6270);
nor U7249 (N_7249,N_6367,N_6419);
nor U7250 (N_7250,N_6281,N_6705);
xnor U7251 (N_7251,N_6476,N_6666);
nand U7252 (N_7252,N_6686,N_6262);
and U7253 (N_7253,N_6523,N_6250);
and U7254 (N_7254,N_6423,N_6522);
xnor U7255 (N_7255,N_6759,N_6443);
and U7256 (N_7256,N_6296,N_6443);
or U7257 (N_7257,N_6401,N_6545);
xnor U7258 (N_7258,N_6593,N_6822);
xnor U7259 (N_7259,N_6837,N_6688);
xnor U7260 (N_7260,N_6290,N_6536);
xor U7261 (N_7261,N_6483,N_6493);
xnor U7262 (N_7262,N_6266,N_6346);
and U7263 (N_7263,N_6310,N_6671);
nand U7264 (N_7264,N_6317,N_6302);
nor U7265 (N_7265,N_6456,N_6251);
xnor U7266 (N_7266,N_6355,N_6656);
nor U7267 (N_7267,N_6782,N_6837);
xnor U7268 (N_7268,N_6386,N_6364);
xor U7269 (N_7269,N_6423,N_6539);
nor U7270 (N_7270,N_6648,N_6828);
nor U7271 (N_7271,N_6409,N_6604);
nand U7272 (N_7272,N_6863,N_6512);
and U7273 (N_7273,N_6753,N_6568);
and U7274 (N_7274,N_6328,N_6667);
or U7275 (N_7275,N_6465,N_6261);
nor U7276 (N_7276,N_6359,N_6583);
nand U7277 (N_7277,N_6340,N_6790);
xor U7278 (N_7278,N_6712,N_6619);
xnor U7279 (N_7279,N_6703,N_6547);
xnor U7280 (N_7280,N_6552,N_6433);
nor U7281 (N_7281,N_6567,N_6737);
xor U7282 (N_7282,N_6307,N_6844);
nor U7283 (N_7283,N_6293,N_6586);
nor U7284 (N_7284,N_6384,N_6778);
or U7285 (N_7285,N_6786,N_6808);
xor U7286 (N_7286,N_6335,N_6464);
nor U7287 (N_7287,N_6743,N_6689);
nand U7288 (N_7288,N_6832,N_6301);
or U7289 (N_7289,N_6324,N_6418);
nand U7290 (N_7290,N_6835,N_6568);
or U7291 (N_7291,N_6540,N_6816);
xnor U7292 (N_7292,N_6638,N_6314);
nand U7293 (N_7293,N_6530,N_6628);
or U7294 (N_7294,N_6482,N_6814);
or U7295 (N_7295,N_6453,N_6868);
xnor U7296 (N_7296,N_6378,N_6498);
nand U7297 (N_7297,N_6731,N_6776);
xor U7298 (N_7298,N_6363,N_6610);
nand U7299 (N_7299,N_6680,N_6487);
or U7300 (N_7300,N_6848,N_6869);
nor U7301 (N_7301,N_6666,N_6787);
nand U7302 (N_7302,N_6637,N_6441);
and U7303 (N_7303,N_6801,N_6762);
or U7304 (N_7304,N_6665,N_6684);
xor U7305 (N_7305,N_6275,N_6662);
and U7306 (N_7306,N_6263,N_6610);
xor U7307 (N_7307,N_6579,N_6395);
and U7308 (N_7308,N_6873,N_6421);
or U7309 (N_7309,N_6562,N_6539);
nor U7310 (N_7310,N_6357,N_6549);
and U7311 (N_7311,N_6385,N_6294);
xnor U7312 (N_7312,N_6299,N_6490);
or U7313 (N_7313,N_6564,N_6519);
nor U7314 (N_7314,N_6460,N_6431);
or U7315 (N_7315,N_6465,N_6762);
nor U7316 (N_7316,N_6764,N_6740);
or U7317 (N_7317,N_6407,N_6740);
and U7318 (N_7318,N_6404,N_6322);
or U7319 (N_7319,N_6293,N_6781);
or U7320 (N_7320,N_6357,N_6278);
nand U7321 (N_7321,N_6584,N_6255);
xor U7322 (N_7322,N_6524,N_6453);
xnor U7323 (N_7323,N_6678,N_6590);
and U7324 (N_7324,N_6305,N_6811);
or U7325 (N_7325,N_6688,N_6799);
and U7326 (N_7326,N_6565,N_6456);
and U7327 (N_7327,N_6724,N_6358);
nor U7328 (N_7328,N_6544,N_6633);
xor U7329 (N_7329,N_6816,N_6763);
or U7330 (N_7330,N_6498,N_6860);
nand U7331 (N_7331,N_6353,N_6437);
nand U7332 (N_7332,N_6407,N_6424);
and U7333 (N_7333,N_6303,N_6515);
nand U7334 (N_7334,N_6366,N_6623);
xnor U7335 (N_7335,N_6794,N_6552);
nand U7336 (N_7336,N_6412,N_6292);
nand U7337 (N_7337,N_6359,N_6743);
or U7338 (N_7338,N_6632,N_6851);
or U7339 (N_7339,N_6303,N_6847);
xor U7340 (N_7340,N_6657,N_6360);
or U7341 (N_7341,N_6333,N_6400);
or U7342 (N_7342,N_6860,N_6473);
nand U7343 (N_7343,N_6250,N_6577);
nand U7344 (N_7344,N_6472,N_6804);
and U7345 (N_7345,N_6326,N_6379);
nor U7346 (N_7346,N_6592,N_6682);
and U7347 (N_7347,N_6325,N_6441);
xor U7348 (N_7348,N_6467,N_6767);
nand U7349 (N_7349,N_6463,N_6811);
nand U7350 (N_7350,N_6543,N_6834);
xor U7351 (N_7351,N_6525,N_6689);
nor U7352 (N_7352,N_6493,N_6434);
xnor U7353 (N_7353,N_6390,N_6846);
or U7354 (N_7354,N_6512,N_6651);
xnor U7355 (N_7355,N_6545,N_6706);
nand U7356 (N_7356,N_6665,N_6833);
xor U7357 (N_7357,N_6799,N_6570);
nor U7358 (N_7358,N_6558,N_6677);
xor U7359 (N_7359,N_6620,N_6747);
and U7360 (N_7360,N_6809,N_6649);
and U7361 (N_7361,N_6460,N_6639);
and U7362 (N_7362,N_6852,N_6390);
nand U7363 (N_7363,N_6398,N_6278);
or U7364 (N_7364,N_6423,N_6407);
and U7365 (N_7365,N_6749,N_6569);
or U7366 (N_7366,N_6827,N_6783);
nor U7367 (N_7367,N_6610,N_6764);
nand U7368 (N_7368,N_6289,N_6608);
xor U7369 (N_7369,N_6868,N_6818);
or U7370 (N_7370,N_6650,N_6329);
nor U7371 (N_7371,N_6479,N_6356);
nand U7372 (N_7372,N_6640,N_6439);
and U7373 (N_7373,N_6684,N_6412);
and U7374 (N_7374,N_6611,N_6649);
and U7375 (N_7375,N_6467,N_6462);
or U7376 (N_7376,N_6584,N_6646);
nand U7377 (N_7377,N_6747,N_6408);
or U7378 (N_7378,N_6757,N_6375);
and U7379 (N_7379,N_6479,N_6526);
or U7380 (N_7380,N_6827,N_6807);
or U7381 (N_7381,N_6695,N_6409);
xor U7382 (N_7382,N_6751,N_6402);
nand U7383 (N_7383,N_6510,N_6720);
nor U7384 (N_7384,N_6709,N_6566);
and U7385 (N_7385,N_6434,N_6835);
or U7386 (N_7386,N_6826,N_6725);
xor U7387 (N_7387,N_6455,N_6337);
or U7388 (N_7388,N_6747,N_6460);
nand U7389 (N_7389,N_6631,N_6730);
nor U7390 (N_7390,N_6364,N_6464);
or U7391 (N_7391,N_6518,N_6788);
xnor U7392 (N_7392,N_6548,N_6826);
or U7393 (N_7393,N_6774,N_6767);
or U7394 (N_7394,N_6614,N_6460);
xor U7395 (N_7395,N_6647,N_6593);
nor U7396 (N_7396,N_6682,N_6863);
xor U7397 (N_7397,N_6706,N_6737);
xnor U7398 (N_7398,N_6440,N_6320);
nand U7399 (N_7399,N_6468,N_6422);
xor U7400 (N_7400,N_6595,N_6643);
xnor U7401 (N_7401,N_6781,N_6642);
and U7402 (N_7402,N_6668,N_6252);
or U7403 (N_7403,N_6396,N_6742);
or U7404 (N_7404,N_6478,N_6674);
nor U7405 (N_7405,N_6809,N_6733);
and U7406 (N_7406,N_6660,N_6563);
xor U7407 (N_7407,N_6643,N_6355);
nor U7408 (N_7408,N_6353,N_6283);
or U7409 (N_7409,N_6395,N_6380);
nor U7410 (N_7410,N_6440,N_6845);
or U7411 (N_7411,N_6526,N_6270);
or U7412 (N_7412,N_6462,N_6321);
and U7413 (N_7413,N_6377,N_6333);
nand U7414 (N_7414,N_6583,N_6326);
xnor U7415 (N_7415,N_6258,N_6778);
nand U7416 (N_7416,N_6371,N_6593);
nor U7417 (N_7417,N_6711,N_6766);
xor U7418 (N_7418,N_6253,N_6404);
xnor U7419 (N_7419,N_6820,N_6673);
or U7420 (N_7420,N_6385,N_6827);
or U7421 (N_7421,N_6319,N_6665);
or U7422 (N_7422,N_6294,N_6500);
nor U7423 (N_7423,N_6305,N_6796);
or U7424 (N_7424,N_6333,N_6288);
or U7425 (N_7425,N_6383,N_6758);
or U7426 (N_7426,N_6280,N_6536);
or U7427 (N_7427,N_6747,N_6815);
nor U7428 (N_7428,N_6861,N_6381);
nor U7429 (N_7429,N_6716,N_6808);
nand U7430 (N_7430,N_6321,N_6398);
and U7431 (N_7431,N_6540,N_6342);
or U7432 (N_7432,N_6558,N_6406);
and U7433 (N_7433,N_6849,N_6341);
nand U7434 (N_7434,N_6349,N_6871);
xnor U7435 (N_7435,N_6726,N_6309);
or U7436 (N_7436,N_6390,N_6671);
and U7437 (N_7437,N_6668,N_6285);
and U7438 (N_7438,N_6757,N_6707);
or U7439 (N_7439,N_6390,N_6398);
xor U7440 (N_7440,N_6524,N_6868);
nand U7441 (N_7441,N_6388,N_6791);
or U7442 (N_7442,N_6274,N_6471);
and U7443 (N_7443,N_6598,N_6715);
or U7444 (N_7444,N_6797,N_6574);
nor U7445 (N_7445,N_6395,N_6559);
nand U7446 (N_7446,N_6347,N_6564);
or U7447 (N_7447,N_6298,N_6797);
xnor U7448 (N_7448,N_6255,N_6440);
nand U7449 (N_7449,N_6335,N_6338);
nand U7450 (N_7450,N_6398,N_6769);
or U7451 (N_7451,N_6454,N_6527);
nor U7452 (N_7452,N_6461,N_6478);
and U7453 (N_7453,N_6731,N_6516);
and U7454 (N_7454,N_6870,N_6701);
and U7455 (N_7455,N_6813,N_6832);
and U7456 (N_7456,N_6769,N_6546);
nor U7457 (N_7457,N_6661,N_6345);
nand U7458 (N_7458,N_6748,N_6451);
and U7459 (N_7459,N_6364,N_6294);
and U7460 (N_7460,N_6285,N_6295);
nand U7461 (N_7461,N_6728,N_6753);
nor U7462 (N_7462,N_6571,N_6755);
nor U7463 (N_7463,N_6680,N_6662);
nor U7464 (N_7464,N_6332,N_6526);
or U7465 (N_7465,N_6869,N_6839);
and U7466 (N_7466,N_6416,N_6301);
nand U7467 (N_7467,N_6817,N_6399);
xor U7468 (N_7468,N_6342,N_6538);
and U7469 (N_7469,N_6560,N_6340);
xor U7470 (N_7470,N_6565,N_6513);
or U7471 (N_7471,N_6357,N_6726);
nand U7472 (N_7472,N_6318,N_6873);
and U7473 (N_7473,N_6275,N_6773);
nand U7474 (N_7474,N_6764,N_6382);
nand U7475 (N_7475,N_6518,N_6692);
nor U7476 (N_7476,N_6358,N_6344);
or U7477 (N_7477,N_6836,N_6822);
and U7478 (N_7478,N_6648,N_6692);
nand U7479 (N_7479,N_6385,N_6318);
and U7480 (N_7480,N_6407,N_6863);
or U7481 (N_7481,N_6457,N_6461);
nand U7482 (N_7482,N_6844,N_6404);
or U7483 (N_7483,N_6655,N_6757);
nand U7484 (N_7484,N_6318,N_6272);
nand U7485 (N_7485,N_6789,N_6477);
nand U7486 (N_7486,N_6517,N_6819);
or U7487 (N_7487,N_6315,N_6633);
and U7488 (N_7488,N_6262,N_6332);
nand U7489 (N_7489,N_6770,N_6563);
xor U7490 (N_7490,N_6279,N_6461);
and U7491 (N_7491,N_6692,N_6860);
nor U7492 (N_7492,N_6259,N_6561);
xor U7493 (N_7493,N_6828,N_6378);
xor U7494 (N_7494,N_6590,N_6332);
or U7495 (N_7495,N_6293,N_6685);
nor U7496 (N_7496,N_6845,N_6705);
nor U7497 (N_7497,N_6590,N_6637);
and U7498 (N_7498,N_6401,N_6366);
and U7499 (N_7499,N_6382,N_6735);
and U7500 (N_7500,N_7273,N_7148);
nand U7501 (N_7501,N_7410,N_7145);
and U7502 (N_7502,N_7332,N_7258);
xnor U7503 (N_7503,N_6976,N_6981);
nand U7504 (N_7504,N_7463,N_7132);
and U7505 (N_7505,N_7337,N_7253);
or U7506 (N_7506,N_7076,N_7450);
and U7507 (N_7507,N_7413,N_7162);
nor U7508 (N_7508,N_7391,N_7173);
and U7509 (N_7509,N_7180,N_7026);
and U7510 (N_7510,N_7248,N_6945);
nor U7511 (N_7511,N_7384,N_7215);
xnor U7512 (N_7512,N_6977,N_7019);
xor U7513 (N_7513,N_7157,N_7404);
or U7514 (N_7514,N_7046,N_7231);
and U7515 (N_7515,N_7269,N_6912);
and U7516 (N_7516,N_6980,N_6999);
nand U7517 (N_7517,N_7047,N_7119);
xor U7518 (N_7518,N_7419,N_7270);
xnor U7519 (N_7519,N_7010,N_6950);
and U7520 (N_7520,N_7444,N_7149);
xnor U7521 (N_7521,N_7007,N_7295);
and U7522 (N_7522,N_7060,N_7000);
nor U7523 (N_7523,N_7255,N_7333);
xnor U7524 (N_7524,N_7197,N_7219);
nor U7525 (N_7525,N_6951,N_7227);
and U7526 (N_7526,N_6926,N_6938);
nor U7527 (N_7527,N_7317,N_7210);
xor U7528 (N_7528,N_6901,N_7266);
xnor U7529 (N_7529,N_6896,N_7446);
nor U7530 (N_7530,N_7044,N_7318);
or U7531 (N_7531,N_7361,N_7238);
xnor U7532 (N_7532,N_7335,N_6965);
nand U7533 (N_7533,N_7191,N_7403);
nand U7534 (N_7534,N_7177,N_6986);
xor U7535 (N_7535,N_7349,N_6947);
and U7536 (N_7536,N_7206,N_7497);
or U7537 (N_7537,N_7251,N_7017);
xor U7538 (N_7538,N_7471,N_7375);
or U7539 (N_7539,N_7345,N_7062);
or U7540 (N_7540,N_7376,N_7240);
nor U7541 (N_7541,N_7336,N_7179);
or U7542 (N_7542,N_7196,N_7280);
nor U7543 (N_7543,N_7261,N_7291);
nor U7544 (N_7544,N_7071,N_7042);
nor U7545 (N_7545,N_6998,N_7385);
xor U7546 (N_7546,N_7469,N_6913);
nor U7547 (N_7547,N_7285,N_7299);
nor U7548 (N_7548,N_7265,N_7095);
or U7549 (N_7549,N_6928,N_7038);
or U7550 (N_7550,N_7088,N_7014);
or U7551 (N_7551,N_7058,N_7478);
or U7552 (N_7552,N_7292,N_6970);
nand U7553 (N_7553,N_7066,N_7396);
nor U7554 (N_7554,N_7399,N_6930);
and U7555 (N_7555,N_6968,N_7004);
nor U7556 (N_7556,N_6987,N_7358);
nand U7557 (N_7557,N_7051,N_7131);
nand U7558 (N_7558,N_7432,N_7288);
and U7559 (N_7559,N_7204,N_6971);
or U7560 (N_7560,N_7302,N_7040);
xnor U7561 (N_7561,N_7479,N_7303);
xor U7562 (N_7562,N_7315,N_6927);
and U7563 (N_7563,N_7327,N_7170);
nor U7564 (N_7564,N_7232,N_6989);
or U7565 (N_7565,N_7125,N_7141);
or U7566 (N_7566,N_7077,N_7343);
and U7567 (N_7567,N_7369,N_6948);
nand U7568 (N_7568,N_7468,N_7439);
nand U7569 (N_7569,N_6904,N_7424);
nand U7570 (N_7570,N_7434,N_6939);
nand U7571 (N_7571,N_7389,N_7164);
or U7572 (N_7572,N_7362,N_7172);
xor U7573 (N_7573,N_7146,N_7277);
nor U7574 (N_7574,N_7281,N_7250);
nor U7575 (N_7575,N_7247,N_6929);
xor U7576 (N_7576,N_6886,N_7454);
and U7577 (N_7577,N_7313,N_6899);
nand U7578 (N_7578,N_6979,N_7344);
or U7579 (N_7579,N_7453,N_6918);
nand U7580 (N_7580,N_6898,N_6982);
or U7581 (N_7581,N_6969,N_7153);
or U7582 (N_7582,N_6889,N_6933);
nor U7583 (N_7583,N_7340,N_7234);
nor U7584 (N_7584,N_7381,N_7449);
nor U7585 (N_7585,N_7049,N_7334);
or U7586 (N_7586,N_7166,N_7118);
and U7587 (N_7587,N_7305,N_7256);
nor U7588 (N_7588,N_7475,N_7325);
or U7589 (N_7589,N_7428,N_6887);
nor U7590 (N_7590,N_7390,N_7368);
and U7591 (N_7591,N_7402,N_7242);
nand U7592 (N_7592,N_7174,N_6924);
xor U7593 (N_7593,N_7211,N_6975);
nor U7594 (N_7594,N_6879,N_7466);
and U7595 (N_7595,N_7121,N_6935);
nor U7596 (N_7596,N_6931,N_7455);
xnor U7597 (N_7597,N_7456,N_7012);
and U7598 (N_7598,N_7073,N_7353);
and U7599 (N_7599,N_7063,N_6902);
nand U7600 (N_7600,N_7161,N_7268);
or U7601 (N_7601,N_7027,N_7300);
and U7602 (N_7602,N_7189,N_7374);
nor U7603 (N_7603,N_7380,N_7018);
xnor U7604 (N_7604,N_7423,N_6900);
or U7605 (N_7605,N_7142,N_7176);
and U7606 (N_7606,N_7022,N_6909);
nor U7607 (N_7607,N_6996,N_7160);
nor U7608 (N_7608,N_7495,N_7101);
or U7609 (N_7609,N_6941,N_7094);
xnor U7610 (N_7610,N_6997,N_7208);
xor U7611 (N_7611,N_7113,N_7346);
xor U7612 (N_7612,N_7339,N_6884);
xor U7613 (N_7613,N_6885,N_7167);
xnor U7614 (N_7614,N_6910,N_7416);
or U7615 (N_7615,N_7430,N_7243);
xnor U7616 (N_7616,N_7275,N_7043);
or U7617 (N_7617,N_7059,N_7457);
xor U7618 (N_7618,N_7401,N_6917);
nor U7619 (N_7619,N_7129,N_7100);
nand U7620 (N_7620,N_7322,N_7233);
and U7621 (N_7621,N_7283,N_7476);
nor U7622 (N_7622,N_7482,N_7356);
nand U7623 (N_7623,N_6934,N_7003);
nand U7624 (N_7624,N_7392,N_6920);
nor U7625 (N_7625,N_7331,N_7351);
and U7626 (N_7626,N_7134,N_6990);
or U7627 (N_7627,N_7214,N_7330);
xnor U7628 (N_7628,N_7110,N_7140);
xor U7629 (N_7629,N_7224,N_7383);
nand U7630 (N_7630,N_6959,N_7225);
and U7631 (N_7631,N_7421,N_7407);
xor U7632 (N_7632,N_7090,N_7105);
nand U7633 (N_7633,N_7481,N_7467);
nor U7634 (N_7634,N_7382,N_7309);
nand U7635 (N_7635,N_7267,N_7154);
or U7636 (N_7636,N_7218,N_7130);
or U7637 (N_7637,N_7326,N_6978);
or U7638 (N_7638,N_7108,N_7279);
nor U7639 (N_7639,N_6890,N_7460);
and U7640 (N_7640,N_6916,N_7257);
and U7641 (N_7641,N_6952,N_7087);
or U7642 (N_7642,N_7143,N_7494);
xnor U7643 (N_7643,N_7035,N_6993);
or U7644 (N_7644,N_6949,N_7239);
nand U7645 (N_7645,N_7459,N_7081);
xnor U7646 (N_7646,N_7338,N_7477);
xor U7647 (N_7647,N_7308,N_7365);
or U7648 (N_7648,N_7122,N_7438);
and U7649 (N_7649,N_7237,N_6907);
xor U7650 (N_7650,N_6966,N_7249);
xor U7651 (N_7651,N_7103,N_7433);
nor U7652 (N_7652,N_7072,N_7386);
xor U7653 (N_7653,N_7021,N_7470);
and U7654 (N_7654,N_6925,N_7098);
and U7655 (N_7655,N_7414,N_6992);
and U7656 (N_7656,N_7229,N_7395);
xnor U7657 (N_7657,N_7425,N_7363);
and U7658 (N_7658,N_7418,N_7074);
nor U7659 (N_7659,N_7067,N_7082);
and U7660 (N_7660,N_7093,N_7397);
nor U7661 (N_7661,N_7039,N_7441);
nand U7662 (N_7662,N_7111,N_7024);
nor U7663 (N_7663,N_7474,N_6943);
and U7664 (N_7664,N_7075,N_7178);
xnor U7665 (N_7665,N_7289,N_7379);
nor U7666 (N_7666,N_6876,N_7055);
nand U7667 (N_7667,N_6946,N_7230);
nor U7668 (N_7668,N_7272,N_7394);
nand U7669 (N_7669,N_6983,N_7321);
xor U7670 (N_7670,N_7411,N_7451);
and U7671 (N_7671,N_6963,N_7084);
or U7672 (N_7672,N_7053,N_7310);
nor U7673 (N_7673,N_7306,N_7246);
nor U7674 (N_7674,N_7184,N_6881);
xor U7675 (N_7675,N_7028,N_7034);
or U7676 (N_7676,N_7106,N_6967);
or U7677 (N_7677,N_6960,N_7284);
nand U7678 (N_7678,N_6937,N_7168);
nand U7679 (N_7679,N_7083,N_6894);
nand U7680 (N_7680,N_7480,N_7462);
and U7681 (N_7681,N_7092,N_7473);
nand U7682 (N_7682,N_7169,N_7221);
xor U7683 (N_7683,N_7190,N_6908);
nor U7684 (N_7684,N_6954,N_7437);
or U7685 (N_7685,N_7228,N_7415);
nor U7686 (N_7686,N_7187,N_7427);
nor U7687 (N_7687,N_7276,N_7205);
and U7688 (N_7688,N_7117,N_7278);
xor U7689 (N_7689,N_7138,N_7316);
nor U7690 (N_7690,N_7194,N_7127);
nand U7691 (N_7691,N_7274,N_7156);
and U7692 (N_7692,N_7136,N_7492);
and U7693 (N_7693,N_7175,N_6914);
or U7694 (N_7694,N_7364,N_7484);
nor U7695 (N_7695,N_6984,N_7171);
nor U7696 (N_7696,N_7264,N_7448);
and U7697 (N_7697,N_7398,N_7135);
and U7698 (N_7698,N_7199,N_6932);
and U7699 (N_7699,N_6974,N_7298);
or U7700 (N_7700,N_6923,N_7252);
xnor U7701 (N_7701,N_7400,N_7220);
nand U7702 (N_7702,N_7236,N_7151);
nor U7703 (N_7703,N_7420,N_7186);
nor U7704 (N_7704,N_6962,N_7036);
xnor U7705 (N_7705,N_7352,N_6955);
or U7706 (N_7706,N_7417,N_7133);
and U7707 (N_7707,N_7263,N_7045);
or U7708 (N_7708,N_7002,N_7096);
nand U7709 (N_7709,N_7183,N_7112);
or U7710 (N_7710,N_6961,N_7254);
xor U7711 (N_7711,N_7314,N_6972);
xnor U7712 (N_7712,N_7408,N_7486);
xor U7713 (N_7713,N_7294,N_7202);
nand U7714 (N_7714,N_7097,N_7282);
nor U7715 (N_7715,N_7359,N_7354);
and U7716 (N_7716,N_6892,N_7104);
nor U7717 (N_7717,N_7393,N_7188);
xnor U7718 (N_7718,N_7465,N_7445);
nor U7719 (N_7719,N_7209,N_6877);
or U7720 (N_7720,N_7241,N_7442);
xor U7721 (N_7721,N_7086,N_7217);
nand U7722 (N_7722,N_7472,N_6880);
nand U7723 (N_7723,N_7013,N_7213);
and U7724 (N_7724,N_7159,N_7371);
and U7725 (N_7725,N_7052,N_7037);
xnor U7726 (N_7726,N_6903,N_6958);
or U7727 (N_7727,N_6919,N_7378);
or U7728 (N_7728,N_7311,N_7426);
and U7729 (N_7729,N_7496,N_7422);
or U7730 (N_7730,N_6883,N_7005);
or U7731 (N_7731,N_7015,N_7009);
nor U7732 (N_7732,N_6897,N_7091);
xor U7733 (N_7733,N_7079,N_7025);
nor U7734 (N_7734,N_7259,N_7489);
xor U7735 (N_7735,N_7226,N_7262);
or U7736 (N_7736,N_7447,N_6953);
or U7737 (N_7737,N_6891,N_7355);
and U7738 (N_7738,N_7078,N_7297);
and U7739 (N_7739,N_7409,N_7350);
nand U7740 (N_7740,N_6956,N_7307);
nand U7741 (N_7741,N_7287,N_7499);
and U7742 (N_7742,N_7452,N_7114);
nand U7743 (N_7743,N_7023,N_7011);
xnor U7744 (N_7744,N_7443,N_6994);
nand U7745 (N_7745,N_7296,N_7057);
nand U7746 (N_7746,N_7271,N_7286);
nor U7747 (N_7747,N_7431,N_7487);
nand U7748 (N_7748,N_7033,N_7373);
nand U7749 (N_7749,N_7367,N_7244);
nand U7750 (N_7750,N_7464,N_6921);
xnor U7751 (N_7751,N_7323,N_6888);
nor U7752 (N_7752,N_7069,N_6944);
xnor U7753 (N_7753,N_7319,N_7498);
or U7754 (N_7754,N_7128,N_7320);
xnor U7755 (N_7755,N_7341,N_6922);
or U7756 (N_7756,N_7366,N_7152);
nor U7757 (N_7757,N_6936,N_7245);
or U7758 (N_7758,N_6911,N_7031);
nand U7759 (N_7759,N_6942,N_7436);
xor U7760 (N_7760,N_6895,N_7137);
xor U7761 (N_7761,N_7068,N_7109);
or U7762 (N_7762,N_7328,N_7372);
xnor U7763 (N_7763,N_6985,N_7201);
or U7764 (N_7764,N_7488,N_7008);
nand U7765 (N_7765,N_7064,N_7029);
nor U7766 (N_7766,N_7405,N_7020);
and U7767 (N_7767,N_7120,N_7387);
or U7768 (N_7768,N_7099,N_7493);
xor U7769 (N_7769,N_7032,N_7357);
nor U7770 (N_7770,N_7491,N_7185);
nand U7771 (N_7771,N_7126,N_7198);
and U7772 (N_7772,N_7412,N_6875);
nand U7773 (N_7773,N_6964,N_7192);
nor U7774 (N_7774,N_7216,N_7144);
or U7775 (N_7775,N_7070,N_7016);
or U7776 (N_7776,N_6995,N_7429);
and U7777 (N_7777,N_6906,N_7054);
nand U7778 (N_7778,N_7203,N_6915);
and U7779 (N_7779,N_7163,N_7085);
nor U7780 (N_7780,N_6882,N_7006);
nor U7781 (N_7781,N_7388,N_6893);
nor U7782 (N_7782,N_6988,N_7195);
nand U7783 (N_7783,N_7080,N_7342);
nor U7784 (N_7784,N_7158,N_6905);
or U7785 (N_7785,N_7182,N_7139);
nand U7786 (N_7786,N_7123,N_7360);
xnor U7787 (N_7787,N_7347,N_7200);
nand U7788 (N_7788,N_7001,N_7193);
and U7789 (N_7789,N_7223,N_7293);
xnor U7790 (N_7790,N_7107,N_7458);
xor U7791 (N_7791,N_7102,N_7370);
or U7792 (N_7792,N_7124,N_7048);
nand U7793 (N_7793,N_7312,N_7324);
nand U7794 (N_7794,N_7061,N_7165);
nand U7795 (N_7795,N_7377,N_7212);
nor U7796 (N_7796,N_7116,N_7301);
xor U7797 (N_7797,N_7147,N_7406);
and U7798 (N_7798,N_7440,N_7235);
xnor U7799 (N_7799,N_7222,N_7329);
xnor U7800 (N_7800,N_6973,N_7490);
nor U7801 (N_7801,N_6957,N_7304);
or U7802 (N_7802,N_7115,N_7155);
nand U7803 (N_7803,N_7435,N_7056);
xnor U7804 (N_7804,N_7150,N_7207);
nor U7805 (N_7805,N_6991,N_7260);
xnor U7806 (N_7806,N_7461,N_7485);
and U7807 (N_7807,N_7181,N_7348);
nand U7808 (N_7808,N_7483,N_6878);
nand U7809 (N_7809,N_7065,N_7290);
nand U7810 (N_7810,N_7089,N_7050);
nor U7811 (N_7811,N_7041,N_6940);
nor U7812 (N_7812,N_7030,N_7165);
nand U7813 (N_7813,N_7178,N_7313);
nor U7814 (N_7814,N_7012,N_7204);
and U7815 (N_7815,N_7457,N_7038);
xor U7816 (N_7816,N_7275,N_6900);
nand U7817 (N_7817,N_6926,N_7320);
nor U7818 (N_7818,N_6915,N_7153);
and U7819 (N_7819,N_6965,N_7459);
or U7820 (N_7820,N_7469,N_7357);
nor U7821 (N_7821,N_7012,N_7158);
xnor U7822 (N_7822,N_7437,N_7325);
nor U7823 (N_7823,N_7274,N_7348);
and U7824 (N_7824,N_7050,N_7154);
nor U7825 (N_7825,N_7127,N_7341);
or U7826 (N_7826,N_7345,N_7250);
and U7827 (N_7827,N_7185,N_7177);
xor U7828 (N_7828,N_7473,N_6903);
nand U7829 (N_7829,N_6977,N_7093);
xor U7830 (N_7830,N_7110,N_6910);
nand U7831 (N_7831,N_7194,N_7486);
nand U7832 (N_7832,N_7083,N_6904);
nor U7833 (N_7833,N_7314,N_7123);
nor U7834 (N_7834,N_6886,N_7394);
or U7835 (N_7835,N_7300,N_7382);
and U7836 (N_7836,N_7147,N_7129);
nand U7837 (N_7837,N_7441,N_6964);
nor U7838 (N_7838,N_7345,N_7158);
xnor U7839 (N_7839,N_7044,N_7423);
xnor U7840 (N_7840,N_7210,N_7078);
nand U7841 (N_7841,N_7484,N_7121);
nor U7842 (N_7842,N_7236,N_7470);
xnor U7843 (N_7843,N_6900,N_7082);
and U7844 (N_7844,N_6997,N_7267);
xnor U7845 (N_7845,N_7431,N_6943);
or U7846 (N_7846,N_7380,N_7320);
or U7847 (N_7847,N_7201,N_6972);
nor U7848 (N_7848,N_7083,N_7110);
xor U7849 (N_7849,N_7132,N_7300);
nor U7850 (N_7850,N_7481,N_7049);
xor U7851 (N_7851,N_7192,N_7444);
and U7852 (N_7852,N_7337,N_7247);
nand U7853 (N_7853,N_7076,N_6946);
nor U7854 (N_7854,N_6939,N_7482);
nand U7855 (N_7855,N_6912,N_7212);
and U7856 (N_7856,N_7117,N_7127);
nand U7857 (N_7857,N_7421,N_7413);
and U7858 (N_7858,N_7451,N_7321);
and U7859 (N_7859,N_7102,N_6950);
xor U7860 (N_7860,N_6932,N_6936);
nor U7861 (N_7861,N_7013,N_7427);
xnor U7862 (N_7862,N_7008,N_7215);
and U7863 (N_7863,N_7495,N_7366);
nand U7864 (N_7864,N_7246,N_6954);
xor U7865 (N_7865,N_7051,N_7070);
nand U7866 (N_7866,N_7202,N_7110);
or U7867 (N_7867,N_7463,N_7394);
xnor U7868 (N_7868,N_6891,N_7453);
or U7869 (N_7869,N_7126,N_7354);
nand U7870 (N_7870,N_7445,N_6913);
and U7871 (N_7871,N_7066,N_7145);
or U7872 (N_7872,N_6981,N_7364);
nor U7873 (N_7873,N_7339,N_7248);
or U7874 (N_7874,N_7277,N_7427);
xor U7875 (N_7875,N_6908,N_7342);
and U7876 (N_7876,N_7153,N_7064);
nand U7877 (N_7877,N_7025,N_6897);
nor U7878 (N_7878,N_7382,N_7438);
xor U7879 (N_7879,N_7235,N_7323);
or U7880 (N_7880,N_7197,N_7464);
nor U7881 (N_7881,N_7146,N_7025);
or U7882 (N_7882,N_6932,N_6940);
nand U7883 (N_7883,N_7193,N_6899);
xor U7884 (N_7884,N_6910,N_7447);
xor U7885 (N_7885,N_7468,N_7236);
or U7886 (N_7886,N_6914,N_7131);
or U7887 (N_7887,N_7228,N_7031);
and U7888 (N_7888,N_7317,N_7156);
nor U7889 (N_7889,N_6949,N_7085);
or U7890 (N_7890,N_7437,N_7129);
and U7891 (N_7891,N_7185,N_7490);
and U7892 (N_7892,N_7083,N_7314);
nor U7893 (N_7893,N_7410,N_6886);
or U7894 (N_7894,N_7244,N_6959);
or U7895 (N_7895,N_7476,N_7305);
and U7896 (N_7896,N_7179,N_6912);
or U7897 (N_7897,N_7315,N_7436);
xnor U7898 (N_7898,N_7426,N_6934);
xor U7899 (N_7899,N_6940,N_7464);
and U7900 (N_7900,N_7163,N_7364);
and U7901 (N_7901,N_6943,N_7311);
or U7902 (N_7902,N_6977,N_7409);
xor U7903 (N_7903,N_6886,N_7212);
or U7904 (N_7904,N_7110,N_7482);
and U7905 (N_7905,N_6975,N_7279);
or U7906 (N_7906,N_7229,N_7172);
nand U7907 (N_7907,N_7224,N_7115);
or U7908 (N_7908,N_6956,N_7115);
nor U7909 (N_7909,N_7425,N_7085);
xor U7910 (N_7910,N_7314,N_7487);
nor U7911 (N_7911,N_6980,N_7434);
xnor U7912 (N_7912,N_7387,N_6919);
xnor U7913 (N_7913,N_7302,N_7418);
or U7914 (N_7914,N_7454,N_7298);
nor U7915 (N_7915,N_7131,N_6887);
nor U7916 (N_7916,N_7424,N_7461);
nor U7917 (N_7917,N_6890,N_6895);
xor U7918 (N_7918,N_7313,N_7317);
nor U7919 (N_7919,N_7108,N_7342);
nor U7920 (N_7920,N_7461,N_7177);
xor U7921 (N_7921,N_7000,N_7186);
or U7922 (N_7922,N_7357,N_6934);
or U7923 (N_7923,N_7004,N_7071);
or U7924 (N_7924,N_7248,N_7312);
xor U7925 (N_7925,N_6889,N_7262);
or U7926 (N_7926,N_7272,N_7342);
xor U7927 (N_7927,N_6984,N_7178);
nor U7928 (N_7928,N_7148,N_6916);
and U7929 (N_7929,N_7302,N_7492);
nor U7930 (N_7930,N_7309,N_7067);
nor U7931 (N_7931,N_7031,N_7044);
nand U7932 (N_7932,N_7104,N_7008);
and U7933 (N_7933,N_7040,N_7208);
and U7934 (N_7934,N_7158,N_7023);
nor U7935 (N_7935,N_7061,N_7125);
xor U7936 (N_7936,N_6914,N_6975);
xnor U7937 (N_7937,N_7079,N_6880);
nand U7938 (N_7938,N_6932,N_6963);
and U7939 (N_7939,N_7107,N_7299);
nor U7940 (N_7940,N_6937,N_7220);
or U7941 (N_7941,N_7098,N_7070);
and U7942 (N_7942,N_7046,N_7182);
or U7943 (N_7943,N_6962,N_7279);
or U7944 (N_7944,N_7225,N_7443);
and U7945 (N_7945,N_7245,N_7220);
xor U7946 (N_7946,N_7151,N_7277);
nand U7947 (N_7947,N_7383,N_7093);
nand U7948 (N_7948,N_7245,N_7230);
xnor U7949 (N_7949,N_7318,N_6884);
or U7950 (N_7950,N_7240,N_6915);
nand U7951 (N_7951,N_7484,N_6941);
nor U7952 (N_7952,N_7272,N_7087);
xor U7953 (N_7953,N_7204,N_7441);
or U7954 (N_7954,N_7404,N_6919);
or U7955 (N_7955,N_7105,N_7356);
xor U7956 (N_7956,N_6967,N_7374);
and U7957 (N_7957,N_7296,N_7140);
nand U7958 (N_7958,N_7011,N_7384);
and U7959 (N_7959,N_7095,N_7106);
or U7960 (N_7960,N_6940,N_7390);
xnor U7961 (N_7961,N_7432,N_7374);
and U7962 (N_7962,N_7100,N_7217);
nand U7963 (N_7963,N_7175,N_7168);
nor U7964 (N_7964,N_7048,N_7492);
nand U7965 (N_7965,N_7231,N_7117);
xnor U7966 (N_7966,N_7088,N_7409);
xor U7967 (N_7967,N_7359,N_7448);
or U7968 (N_7968,N_7247,N_7400);
nor U7969 (N_7969,N_7001,N_7434);
or U7970 (N_7970,N_7377,N_7266);
nand U7971 (N_7971,N_7188,N_7366);
or U7972 (N_7972,N_7302,N_7092);
nor U7973 (N_7973,N_7211,N_7146);
and U7974 (N_7974,N_7431,N_7033);
nor U7975 (N_7975,N_7426,N_7348);
nor U7976 (N_7976,N_7446,N_6936);
and U7977 (N_7977,N_7186,N_6984);
nor U7978 (N_7978,N_7351,N_7219);
nor U7979 (N_7979,N_7468,N_7315);
nand U7980 (N_7980,N_7285,N_7270);
or U7981 (N_7981,N_7299,N_7255);
or U7982 (N_7982,N_7233,N_6881);
xnor U7983 (N_7983,N_7243,N_7362);
or U7984 (N_7984,N_6881,N_7310);
xnor U7985 (N_7985,N_7301,N_7106);
nand U7986 (N_7986,N_7114,N_7137);
or U7987 (N_7987,N_7070,N_7258);
and U7988 (N_7988,N_7005,N_7245);
nand U7989 (N_7989,N_6925,N_7311);
xor U7990 (N_7990,N_7194,N_7109);
nand U7991 (N_7991,N_7431,N_7133);
xnor U7992 (N_7992,N_7009,N_7294);
nor U7993 (N_7993,N_7261,N_7486);
nor U7994 (N_7994,N_6982,N_7200);
or U7995 (N_7995,N_7347,N_6895);
nor U7996 (N_7996,N_7444,N_7418);
or U7997 (N_7997,N_7448,N_7207);
xor U7998 (N_7998,N_6900,N_7016);
and U7999 (N_7999,N_7145,N_7298);
and U8000 (N_8000,N_7118,N_7010);
or U8001 (N_8001,N_7368,N_7042);
nand U8002 (N_8002,N_7187,N_7374);
or U8003 (N_8003,N_6967,N_7089);
or U8004 (N_8004,N_6886,N_7492);
and U8005 (N_8005,N_7320,N_7140);
nand U8006 (N_8006,N_6918,N_7416);
xnor U8007 (N_8007,N_7020,N_7053);
xor U8008 (N_8008,N_7291,N_7119);
nor U8009 (N_8009,N_6916,N_7008);
nand U8010 (N_8010,N_7249,N_6923);
xor U8011 (N_8011,N_7277,N_7102);
nor U8012 (N_8012,N_6936,N_6970);
nor U8013 (N_8013,N_7345,N_7301);
xnor U8014 (N_8014,N_7475,N_7007);
nor U8015 (N_8015,N_6970,N_7001);
or U8016 (N_8016,N_7293,N_7086);
nand U8017 (N_8017,N_7467,N_7235);
nand U8018 (N_8018,N_7000,N_6997);
xor U8019 (N_8019,N_7197,N_7467);
and U8020 (N_8020,N_6889,N_7265);
or U8021 (N_8021,N_7281,N_6996);
and U8022 (N_8022,N_7252,N_7128);
nand U8023 (N_8023,N_7393,N_7047);
and U8024 (N_8024,N_7145,N_6927);
nor U8025 (N_8025,N_7317,N_7088);
or U8026 (N_8026,N_7242,N_7284);
and U8027 (N_8027,N_7413,N_6887);
nor U8028 (N_8028,N_7072,N_7423);
nor U8029 (N_8029,N_6940,N_7158);
nand U8030 (N_8030,N_7376,N_7418);
xor U8031 (N_8031,N_6887,N_7344);
nor U8032 (N_8032,N_7296,N_7391);
or U8033 (N_8033,N_6953,N_7152);
xnor U8034 (N_8034,N_7309,N_7400);
or U8035 (N_8035,N_7411,N_7079);
nand U8036 (N_8036,N_7380,N_7021);
and U8037 (N_8037,N_6927,N_7234);
and U8038 (N_8038,N_6907,N_7337);
nand U8039 (N_8039,N_7464,N_7118);
nand U8040 (N_8040,N_7148,N_6897);
and U8041 (N_8041,N_7246,N_7310);
or U8042 (N_8042,N_6885,N_7220);
and U8043 (N_8043,N_6890,N_7477);
and U8044 (N_8044,N_7271,N_6952);
or U8045 (N_8045,N_6997,N_6968);
and U8046 (N_8046,N_6970,N_7467);
and U8047 (N_8047,N_7189,N_7444);
nor U8048 (N_8048,N_7169,N_6892);
xnor U8049 (N_8049,N_7251,N_7429);
nand U8050 (N_8050,N_7160,N_7078);
or U8051 (N_8051,N_7320,N_7431);
or U8052 (N_8052,N_6959,N_7138);
nor U8053 (N_8053,N_7043,N_7187);
nand U8054 (N_8054,N_7233,N_7147);
nand U8055 (N_8055,N_7369,N_6950);
nor U8056 (N_8056,N_7488,N_7199);
nor U8057 (N_8057,N_7344,N_7050);
or U8058 (N_8058,N_6948,N_7432);
xor U8059 (N_8059,N_7377,N_7311);
or U8060 (N_8060,N_6897,N_7340);
nand U8061 (N_8061,N_6983,N_6942);
and U8062 (N_8062,N_7402,N_7435);
and U8063 (N_8063,N_7040,N_7119);
nand U8064 (N_8064,N_7126,N_7495);
and U8065 (N_8065,N_6936,N_7064);
nor U8066 (N_8066,N_7436,N_7270);
nor U8067 (N_8067,N_7114,N_7310);
or U8068 (N_8068,N_7371,N_7092);
and U8069 (N_8069,N_7432,N_7208);
and U8070 (N_8070,N_7313,N_6966);
xor U8071 (N_8071,N_7145,N_7339);
and U8072 (N_8072,N_7466,N_6931);
or U8073 (N_8073,N_7433,N_7095);
nor U8074 (N_8074,N_6958,N_7015);
nor U8075 (N_8075,N_7156,N_6890);
nor U8076 (N_8076,N_7255,N_7254);
nor U8077 (N_8077,N_6897,N_6904);
xnor U8078 (N_8078,N_6943,N_6983);
nand U8079 (N_8079,N_7217,N_7453);
and U8080 (N_8080,N_7172,N_7214);
and U8081 (N_8081,N_7160,N_7341);
or U8082 (N_8082,N_6951,N_7487);
and U8083 (N_8083,N_7111,N_7108);
xnor U8084 (N_8084,N_7490,N_7012);
nor U8085 (N_8085,N_7375,N_6906);
or U8086 (N_8086,N_7098,N_7018);
nand U8087 (N_8087,N_7449,N_7334);
or U8088 (N_8088,N_7410,N_7272);
and U8089 (N_8089,N_6982,N_7142);
and U8090 (N_8090,N_7325,N_7071);
or U8091 (N_8091,N_6951,N_7307);
and U8092 (N_8092,N_7489,N_6988);
or U8093 (N_8093,N_7207,N_7233);
nand U8094 (N_8094,N_7176,N_7417);
and U8095 (N_8095,N_7459,N_7287);
nor U8096 (N_8096,N_7080,N_6934);
nand U8097 (N_8097,N_7208,N_6891);
xor U8098 (N_8098,N_6994,N_7076);
nor U8099 (N_8099,N_7344,N_7275);
nand U8100 (N_8100,N_7176,N_7311);
nor U8101 (N_8101,N_7358,N_6925);
or U8102 (N_8102,N_7347,N_7442);
nor U8103 (N_8103,N_7006,N_6978);
or U8104 (N_8104,N_6910,N_7326);
nand U8105 (N_8105,N_7480,N_7270);
nand U8106 (N_8106,N_7243,N_7057);
nor U8107 (N_8107,N_7269,N_6911);
xor U8108 (N_8108,N_7153,N_7409);
nor U8109 (N_8109,N_7003,N_7113);
nor U8110 (N_8110,N_7378,N_7239);
nor U8111 (N_8111,N_6877,N_7464);
and U8112 (N_8112,N_7203,N_7405);
nand U8113 (N_8113,N_6954,N_7187);
nand U8114 (N_8114,N_7093,N_7442);
xnor U8115 (N_8115,N_6926,N_7105);
or U8116 (N_8116,N_7458,N_7488);
and U8117 (N_8117,N_7046,N_7127);
nor U8118 (N_8118,N_7032,N_7141);
nand U8119 (N_8119,N_7274,N_7201);
nor U8120 (N_8120,N_7378,N_7253);
xnor U8121 (N_8121,N_6936,N_7363);
and U8122 (N_8122,N_7255,N_7397);
and U8123 (N_8123,N_7262,N_7100);
nand U8124 (N_8124,N_7326,N_7099);
and U8125 (N_8125,N_7540,N_7801);
nor U8126 (N_8126,N_7525,N_7637);
nor U8127 (N_8127,N_7994,N_7656);
nor U8128 (N_8128,N_8075,N_8008);
xor U8129 (N_8129,N_7545,N_7918);
nor U8130 (N_8130,N_7975,N_7507);
nand U8131 (N_8131,N_7935,N_7881);
and U8132 (N_8132,N_7817,N_7627);
or U8133 (N_8133,N_8067,N_7800);
and U8134 (N_8134,N_7899,N_7731);
and U8135 (N_8135,N_7745,N_7527);
nor U8136 (N_8136,N_7551,N_8070);
or U8137 (N_8137,N_7596,N_8032);
or U8138 (N_8138,N_7886,N_7981);
nand U8139 (N_8139,N_7968,N_7699);
or U8140 (N_8140,N_7766,N_7575);
nand U8141 (N_8141,N_7970,N_7837);
xor U8142 (N_8142,N_7520,N_8011);
nand U8143 (N_8143,N_7997,N_7664);
nor U8144 (N_8144,N_7762,N_7868);
nand U8145 (N_8145,N_7541,N_8046);
nand U8146 (N_8146,N_7585,N_7707);
nor U8147 (N_8147,N_7717,N_7539);
nor U8148 (N_8148,N_8002,N_8082);
and U8149 (N_8149,N_7849,N_7647);
nor U8150 (N_8150,N_7865,N_7802);
and U8151 (N_8151,N_7770,N_7963);
and U8152 (N_8152,N_8071,N_7913);
and U8153 (N_8153,N_8050,N_7526);
nor U8154 (N_8154,N_7660,N_7738);
or U8155 (N_8155,N_7673,N_7787);
xor U8156 (N_8156,N_7680,N_8051);
xnor U8157 (N_8157,N_7819,N_7923);
and U8158 (N_8158,N_7916,N_8117);
nor U8159 (N_8159,N_7677,N_8030);
nor U8160 (N_8160,N_8012,N_7531);
nor U8161 (N_8161,N_7910,N_7911);
or U8162 (N_8162,N_7879,N_7948);
and U8163 (N_8163,N_7934,N_7518);
nand U8164 (N_8164,N_7659,N_7511);
nand U8165 (N_8165,N_8119,N_8007);
nand U8166 (N_8166,N_7562,N_7654);
nor U8167 (N_8167,N_7907,N_7856);
nor U8168 (N_8168,N_8102,N_7998);
nand U8169 (N_8169,N_8110,N_7603);
xnor U8170 (N_8170,N_7506,N_7846);
nand U8171 (N_8171,N_8076,N_7550);
nand U8172 (N_8172,N_7564,N_7676);
xor U8173 (N_8173,N_7712,N_7876);
and U8174 (N_8174,N_7862,N_7776);
nor U8175 (N_8175,N_7920,N_7696);
xor U8176 (N_8176,N_7548,N_7845);
nor U8177 (N_8177,N_7620,N_7769);
or U8178 (N_8178,N_8006,N_8014);
nor U8179 (N_8179,N_7915,N_7552);
nor U8180 (N_8180,N_8044,N_7543);
xnor U8181 (N_8181,N_7852,N_7653);
or U8182 (N_8182,N_7591,N_7804);
and U8183 (N_8183,N_7624,N_7874);
and U8184 (N_8184,N_7588,N_7625);
nand U8185 (N_8185,N_7622,N_7686);
and U8186 (N_8186,N_7718,N_7985);
xnor U8187 (N_8187,N_7533,N_8057);
nand U8188 (N_8188,N_8037,N_7888);
xnor U8189 (N_8189,N_7767,N_7955);
xor U8190 (N_8190,N_7748,N_8062);
and U8191 (N_8191,N_7559,N_7754);
and U8192 (N_8192,N_7840,N_7880);
nor U8193 (N_8193,N_8040,N_7989);
xor U8194 (N_8194,N_8053,N_7882);
and U8195 (N_8195,N_7508,N_7959);
nor U8196 (N_8196,N_7872,N_7792);
xnor U8197 (N_8197,N_7752,N_7519);
xnor U8198 (N_8198,N_8020,N_7662);
or U8199 (N_8199,N_7853,N_7690);
xnor U8200 (N_8200,N_7965,N_7933);
or U8201 (N_8201,N_7813,N_7958);
or U8202 (N_8202,N_8120,N_8003);
and U8203 (N_8203,N_7595,N_7655);
and U8204 (N_8204,N_7553,N_8028);
nand U8205 (N_8205,N_7904,N_7715);
and U8206 (N_8206,N_7729,N_7877);
xnor U8207 (N_8207,N_7902,N_7809);
and U8208 (N_8208,N_7784,N_7777);
xnor U8209 (N_8209,N_7972,N_8108);
nand U8210 (N_8210,N_7799,N_7889);
and U8211 (N_8211,N_7633,N_7821);
nor U8212 (N_8212,N_7836,N_7612);
and U8213 (N_8213,N_7786,N_7600);
nand U8214 (N_8214,N_8096,N_8038);
and U8215 (N_8215,N_8042,N_7570);
xor U8216 (N_8216,N_8078,N_7844);
or U8217 (N_8217,N_8095,N_7943);
or U8218 (N_8218,N_7890,N_8063);
or U8219 (N_8219,N_7950,N_7829);
xor U8220 (N_8220,N_7896,N_7884);
or U8221 (N_8221,N_8036,N_8034);
xnor U8222 (N_8222,N_7919,N_7650);
nand U8223 (N_8223,N_7513,N_7720);
xnor U8224 (N_8224,N_8039,N_7628);
and U8225 (N_8225,N_7665,N_7700);
xnor U8226 (N_8226,N_7960,N_7940);
nand U8227 (N_8227,N_7832,N_7798);
or U8228 (N_8228,N_7536,N_8086);
nor U8229 (N_8229,N_8066,N_8004);
and U8230 (N_8230,N_7768,N_7667);
xor U8231 (N_8231,N_8087,N_7704);
xor U8232 (N_8232,N_7638,N_7936);
nor U8233 (N_8233,N_8043,N_7901);
xnor U8234 (N_8234,N_7679,N_7636);
or U8235 (N_8235,N_8103,N_7557);
and U8236 (N_8236,N_7558,N_8085);
xnor U8237 (N_8237,N_7791,N_7706);
and U8238 (N_8238,N_7996,N_8097);
nor U8239 (N_8239,N_8045,N_7579);
and U8240 (N_8240,N_7775,N_8015);
xnor U8241 (N_8241,N_7645,N_8101);
nor U8242 (N_8242,N_7944,N_7721);
or U8243 (N_8243,N_7534,N_7573);
nand U8244 (N_8244,N_8060,N_8111);
xnor U8245 (N_8245,N_7723,N_8059);
xnor U8246 (N_8246,N_7737,N_7713);
or U8247 (N_8247,N_8116,N_7582);
or U8248 (N_8248,N_7567,N_7735);
or U8249 (N_8249,N_7993,N_8022);
nor U8250 (N_8250,N_8080,N_7951);
or U8251 (N_8251,N_7709,N_7510);
or U8252 (N_8252,N_7857,N_7986);
or U8253 (N_8253,N_7546,N_7692);
nand U8254 (N_8254,N_7961,N_7578);
nand U8255 (N_8255,N_7561,N_7749);
and U8256 (N_8256,N_7693,N_8124);
xor U8257 (N_8257,N_8093,N_7885);
nor U8258 (N_8258,N_7708,N_7866);
xor U8259 (N_8259,N_7974,N_7730);
nor U8260 (N_8260,N_7580,N_7710);
or U8261 (N_8261,N_7756,N_8035);
xnor U8262 (N_8262,N_7682,N_7987);
xor U8263 (N_8263,N_7672,N_7674);
and U8264 (N_8264,N_7571,N_8069);
and U8265 (N_8265,N_7788,N_8054);
xor U8266 (N_8266,N_7663,N_7932);
nor U8267 (N_8267,N_7535,N_7529);
or U8268 (N_8268,N_8065,N_7938);
or U8269 (N_8269,N_7605,N_7629);
or U8270 (N_8270,N_7823,N_8048);
xor U8271 (N_8271,N_7893,N_7931);
or U8272 (N_8272,N_7725,N_7668);
or U8273 (N_8273,N_7842,N_8061);
xnor U8274 (N_8274,N_7939,N_7812);
or U8275 (N_8275,N_7678,N_7517);
nor U8276 (N_8276,N_7966,N_7554);
nand U8277 (N_8277,N_7599,N_7694);
or U8278 (N_8278,N_7538,N_8029);
or U8279 (N_8279,N_8094,N_7773);
nand U8280 (N_8280,N_7758,N_8092);
or U8281 (N_8281,N_8041,N_7779);
nor U8282 (N_8282,N_7983,N_7547);
xor U8283 (N_8283,N_8089,N_7514);
nand U8284 (N_8284,N_7670,N_7781);
and U8285 (N_8285,N_7875,N_7666);
or U8286 (N_8286,N_7500,N_7967);
nor U8287 (N_8287,N_7691,N_8001);
xor U8288 (N_8288,N_7626,N_7922);
or U8289 (N_8289,N_7592,N_7505);
xnor U8290 (N_8290,N_7615,N_7765);
xnor U8291 (N_8291,N_7521,N_7905);
and U8292 (N_8292,N_7891,N_7604);
nand U8293 (N_8293,N_8084,N_7528);
xor U8294 (N_8294,N_7532,N_7563);
nor U8295 (N_8295,N_7623,N_8056);
xnor U8296 (N_8296,N_7740,N_8047);
nor U8297 (N_8297,N_7759,N_7681);
and U8298 (N_8298,N_7621,N_7942);
xnor U8299 (N_8299,N_7808,N_7838);
and U8300 (N_8300,N_7785,N_7727);
nor U8301 (N_8301,N_8019,N_7711);
xnor U8302 (N_8302,N_7887,N_8068);
or U8303 (N_8303,N_7794,N_7810);
nor U8304 (N_8304,N_7761,N_7747);
xnor U8305 (N_8305,N_7978,N_8105);
and U8306 (N_8306,N_7930,N_7515);
nor U8307 (N_8307,N_7831,N_7912);
nand U8308 (N_8308,N_7695,N_7607);
nor U8309 (N_8309,N_8115,N_7999);
nand U8310 (N_8310,N_7524,N_7698);
nor U8311 (N_8311,N_7632,N_8017);
nor U8312 (N_8312,N_7892,N_7504);
nand U8313 (N_8313,N_7635,N_8081);
and U8314 (N_8314,N_7805,N_7992);
and U8315 (N_8315,N_7646,N_7598);
nand U8316 (N_8316,N_7764,N_7643);
or U8317 (N_8317,N_8100,N_7614);
xnor U8318 (N_8318,N_8031,N_7608);
or U8319 (N_8319,N_8072,N_7962);
and U8320 (N_8320,N_7512,N_7522);
nor U8321 (N_8321,N_7669,N_7954);
nand U8322 (N_8322,N_8064,N_8026);
nand U8323 (N_8323,N_7976,N_8010);
nand U8324 (N_8324,N_7732,N_8122);
and U8325 (N_8325,N_7991,N_7979);
xor U8326 (N_8326,N_7908,N_7826);
or U8327 (N_8327,N_7878,N_8106);
nor U8328 (N_8328,N_7565,N_7897);
nor U8329 (N_8329,N_7530,N_8112);
nand U8330 (N_8330,N_7658,N_8098);
nand U8331 (N_8331,N_7854,N_7914);
xnor U8332 (N_8332,N_7883,N_7924);
or U8333 (N_8333,N_8118,N_8005);
nand U8334 (N_8334,N_7705,N_8013);
nor U8335 (N_8335,N_7587,N_7611);
nor U8336 (N_8336,N_7793,N_7675);
nand U8337 (N_8337,N_7815,N_7859);
and U8338 (N_8338,N_7824,N_7855);
nor U8339 (N_8339,N_7733,N_7909);
and U8340 (N_8340,N_7661,N_7728);
xnor U8341 (N_8341,N_7778,N_7701);
xor U8342 (N_8342,N_7926,N_7929);
nand U8343 (N_8343,N_7606,N_7617);
or U8344 (N_8344,N_7555,N_7825);
nand U8345 (N_8345,N_7850,N_7689);
and U8346 (N_8346,N_7618,N_7742);
and U8347 (N_8347,N_7927,N_7871);
nand U8348 (N_8348,N_7807,N_7744);
nor U8349 (N_8349,N_7956,N_7542);
and U8350 (N_8350,N_7848,N_7806);
or U8351 (N_8351,N_7895,N_7581);
nand U8352 (N_8352,N_8083,N_7990);
xor U8353 (N_8353,N_7726,N_7640);
nor U8354 (N_8354,N_7988,N_7610);
nor U8355 (N_8355,N_7750,N_7843);
or U8356 (N_8356,N_7949,N_7818);
nand U8357 (N_8357,N_7739,N_8025);
xnor U8358 (N_8358,N_8074,N_8099);
nor U8359 (N_8359,N_7716,N_7964);
and U8360 (N_8360,N_7751,N_7873);
or U8361 (N_8361,N_7577,N_7957);
xor U8362 (N_8362,N_7969,N_7851);
or U8363 (N_8363,N_8090,N_7734);
xor U8364 (N_8364,N_7746,N_7652);
nand U8365 (N_8365,N_7774,N_7523);
and U8366 (N_8366,N_7839,N_8023);
xnor U8367 (N_8367,N_7906,N_7590);
nor U8368 (N_8368,N_7946,N_7569);
and U8369 (N_8369,N_7644,N_7803);
nand U8370 (N_8370,N_7772,N_8073);
nor U8371 (N_8371,N_8009,N_7566);
or U8372 (N_8372,N_7743,N_8113);
xnor U8373 (N_8373,N_7771,N_7811);
and U8374 (N_8374,N_7688,N_7816);
or U8375 (N_8375,N_7619,N_7516);
or U8376 (N_8376,N_8107,N_8123);
xor U8377 (N_8377,N_8055,N_7649);
nor U8378 (N_8378,N_7589,N_7574);
nor U8379 (N_8379,N_7502,N_7642);
nor U8380 (N_8380,N_7861,N_7834);
and U8381 (N_8381,N_8077,N_7789);
and U8382 (N_8382,N_7602,N_7860);
xor U8383 (N_8383,N_7763,N_8052);
xor U8384 (N_8384,N_8033,N_7945);
or U8385 (N_8385,N_7953,N_7741);
or U8386 (N_8386,N_7941,N_7828);
xor U8387 (N_8387,N_7900,N_7830);
and U8388 (N_8388,N_7753,N_7947);
nor U8389 (N_8389,N_7572,N_7984);
xnor U8390 (N_8390,N_7864,N_8018);
xnor U8391 (N_8391,N_8088,N_7714);
or U8392 (N_8392,N_7917,N_7783);
xor U8393 (N_8393,N_7651,N_7835);
or U8394 (N_8394,N_7971,N_7613);
nand U8395 (N_8395,N_8024,N_7833);
and U8396 (N_8396,N_7827,N_7797);
nor U8397 (N_8397,N_7869,N_7544);
xnor U8398 (N_8398,N_7995,N_7980);
nand U8399 (N_8399,N_8104,N_7820);
nor U8400 (N_8400,N_7549,N_7790);
or U8401 (N_8401,N_8049,N_7501);
nor U8402 (N_8402,N_8058,N_7687);
nor U8403 (N_8403,N_7703,N_8079);
and U8404 (N_8404,N_7977,N_7952);
and U8405 (N_8405,N_7657,N_8000);
and U8406 (N_8406,N_7584,N_7641);
or U8407 (N_8407,N_7736,N_8027);
nand U8408 (N_8408,N_7928,N_7583);
nor U8409 (N_8409,N_7867,N_7863);
nand U8410 (N_8410,N_7796,N_7648);
and U8411 (N_8411,N_7782,N_7601);
nand U8412 (N_8412,N_7925,N_7537);
or U8413 (N_8413,N_7858,N_7973);
and U8414 (N_8414,N_8021,N_7671);
nor U8415 (N_8415,N_8121,N_7556);
xnor U8416 (N_8416,N_7780,N_7795);
nor U8417 (N_8417,N_8114,N_7593);
and U8418 (N_8418,N_7503,N_7702);
or U8419 (N_8419,N_7509,N_7841);
nand U8420 (N_8420,N_7685,N_7639);
nor U8421 (N_8421,N_7616,N_7684);
nor U8422 (N_8422,N_7814,N_7937);
xor U8423 (N_8423,N_7568,N_7822);
xnor U8424 (N_8424,N_7982,N_7724);
nor U8425 (N_8425,N_7560,N_7586);
and U8426 (N_8426,N_7683,N_8016);
nor U8427 (N_8427,N_7697,N_8091);
nand U8428 (N_8428,N_7719,N_7594);
nor U8429 (N_8429,N_7631,N_7870);
xnor U8430 (N_8430,N_7921,N_7894);
and U8431 (N_8431,N_8109,N_7576);
nand U8432 (N_8432,N_7847,N_7609);
xnor U8433 (N_8433,N_7760,N_7630);
or U8434 (N_8434,N_7757,N_7634);
xnor U8435 (N_8435,N_7903,N_7597);
nand U8436 (N_8436,N_7722,N_7755);
and U8437 (N_8437,N_7898,N_7593);
or U8438 (N_8438,N_7803,N_7646);
and U8439 (N_8439,N_7685,N_7605);
nand U8440 (N_8440,N_7566,N_7600);
nand U8441 (N_8441,N_7707,N_7595);
or U8442 (N_8442,N_7619,N_7997);
nand U8443 (N_8443,N_7932,N_7736);
xor U8444 (N_8444,N_7737,N_7554);
nand U8445 (N_8445,N_7943,N_7740);
nand U8446 (N_8446,N_7853,N_7738);
xnor U8447 (N_8447,N_7943,N_8119);
xnor U8448 (N_8448,N_8039,N_7850);
xor U8449 (N_8449,N_7794,N_7984);
nor U8450 (N_8450,N_7663,N_7598);
nand U8451 (N_8451,N_8032,N_8040);
or U8452 (N_8452,N_8002,N_8092);
nand U8453 (N_8453,N_7839,N_7543);
and U8454 (N_8454,N_8121,N_8096);
or U8455 (N_8455,N_8115,N_7596);
and U8456 (N_8456,N_8031,N_7604);
and U8457 (N_8457,N_8035,N_7687);
nor U8458 (N_8458,N_8087,N_7594);
or U8459 (N_8459,N_7956,N_7877);
nor U8460 (N_8460,N_7702,N_7767);
xnor U8461 (N_8461,N_7724,N_7744);
and U8462 (N_8462,N_7644,N_7553);
and U8463 (N_8463,N_7908,N_8052);
nand U8464 (N_8464,N_7771,N_7546);
nand U8465 (N_8465,N_7522,N_8102);
and U8466 (N_8466,N_7903,N_7882);
and U8467 (N_8467,N_7636,N_7832);
and U8468 (N_8468,N_7820,N_7960);
xor U8469 (N_8469,N_7849,N_7993);
xnor U8470 (N_8470,N_7928,N_8034);
and U8471 (N_8471,N_7955,N_7740);
and U8472 (N_8472,N_7561,N_7794);
nand U8473 (N_8473,N_7882,N_7864);
nor U8474 (N_8474,N_7815,N_7995);
and U8475 (N_8475,N_7799,N_7941);
nand U8476 (N_8476,N_7938,N_7995);
nor U8477 (N_8477,N_7597,N_7507);
nand U8478 (N_8478,N_7653,N_8087);
or U8479 (N_8479,N_7555,N_8066);
xnor U8480 (N_8480,N_7989,N_7610);
nand U8481 (N_8481,N_7921,N_7796);
xnor U8482 (N_8482,N_7996,N_8098);
or U8483 (N_8483,N_7632,N_7610);
nor U8484 (N_8484,N_7660,N_7899);
or U8485 (N_8485,N_7714,N_7687);
or U8486 (N_8486,N_8099,N_8092);
or U8487 (N_8487,N_7503,N_8118);
nor U8488 (N_8488,N_8015,N_7569);
xor U8489 (N_8489,N_7981,N_7876);
nand U8490 (N_8490,N_7771,N_8099);
nand U8491 (N_8491,N_7537,N_7774);
nor U8492 (N_8492,N_7631,N_7996);
and U8493 (N_8493,N_7524,N_7706);
nand U8494 (N_8494,N_8109,N_7871);
nor U8495 (N_8495,N_7960,N_7691);
xor U8496 (N_8496,N_7727,N_8004);
and U8497 (N_8497,N_7810,N_7859);
nor U8498 (N_8498,N_8098,N_7696);
xor U8499 (N_8499,N_7994,N_8040);
or U8500 (N_8500,N_7567,N_7846);
nor U8501 (N_8501,N_7607,N_7565);
nor U8502 (N_8502,N_7957,N_7803);
xnor U8503 (N_8503,N_7558,N_8088);
and U8504 (N_8504,N_8119,N_7526);
or U8505 (N_8505,N_7601,N_7599);
and U8506 (N_8506,N_8093,N_8052);
nor U8507 (N_8507,N_8007,N_8096);
nand U8508 (N_8508,N_7539,N_7831);
and U8509 (N_8509,N_7865,N_7679);
or U8510 (N_8510,N_7949,N_8037);
and U8511 (N_8511,N_8005,N_7931);
and U8512 (N_8512,N_7669,N_7886);
and U8513 (N_8513,N_7890,N_8051);
xor U8514 (N_8514,N_7519,N_7564);
and U8515 (N_8515,N_7662,N_7666);
and U8516 (N_8516,N_7712,N_7595);
nand U8517 (N_8517,N_8015,N_7930);
and U8518 (N_8518,N_7718,N_7896);
and U8519 (N_8519,N_7709,N_7964);
xnor U8520 (N_8520,N_8037,N_7998);
nand U8521 (N_8521,N_7736,N_7586);
nor U8522 (N_8522,N_8049,N_7868);
and U8523 (N_8523,N_7680,N_7583);
and U8524 (N_8524,N_7856,N_7913);
or U8525 (N_8525,N_7650,N_7516);
xnor U8526 (N_8526,N_7933,N_7907);
xor U8527 (N_8527,N_7591,N_7619);
nor U8528 (N_8528,N_7686,N_7714);
and U8529 (N_8529,N_7562,N_7592);
and U8530 (N_8530,N_7882,N_7697);
and U8531 (N_8531,N_7832,N_8112);
and U8532 (N_8532,N_8087,N_7607);
nand U8533 (N_8533,N_7898,N_7513);
xnor U8534 (N_8534,N_7875,N_7625);
xnor U8535 (N_8535,N_7864,N_7740);
or U8536 (N_8536,N_8101,N_7976);
nor U8537 (N_8537,N_8102,N_7547);
or U8538 (N_8538,N_8043,N_7701);
nor U8539 (N_8539,N_7753,N_7928);
nand U8540 (N_8540,N_7944,N_7985);
or U8541 (N_8541,N_7509,N_7792);
nor U8542 (N_8542,N_7591,N_7882);
xor U8543 (N_8543,N_7890,N_7971);
or U8544 (N_8544,N_8121,N_8117);
xor U8545 (N_8545,N_7659,N_7826);
nand U8546 (N_8546,N_7771,N_8001);
nor U8547 (N_8547,N_8037,N_8107);
and U8548 (N_8548,N_7931,N_8104);
xnor U8549 (N_8549,N_7861,N_7972);
or U8550 (N_8550,N_7824,N_8013);
or U8551 (N_8551,N_7669,N_7692);
nor U8552 (N_8552,N_8069,N_7783);
xor U8553 (N_8553,N_7760,N_7815);
and U8554 (N_8554,N_7981,N_7746);
nand U8555 (N_8555,N_8118,N_7674);
xor U8556 (N_8556,N_7815,N_7912);
or U8557 (N_8557,N_7845,N_8012);
or U8558 (N_8558,N_7549,N_7576);
nand U8559 (N_8559,N_8067,N_8034);
xor U8560 (N_8560,N_7732,N_7809);
nor U8561 (N_8561,N_7520,N_8003);
and U8562 (N_8562,N_7734,N_8096);
or U8563 (N_8563,N_7581,N_7921);
nand U8564 (N_8564,N_7692,N_7507);
nor U8565 (N_8565,N_7694,N_7907);
or U8566 (N_8566,N_7550,N_8124);
and U8567 (N_8567,N_7552,N_7820);
or U8568 (N_8568,N_7840,N_7763);
and U8569 (N_8569,N_7719,N_7870);
nand U8570 (N_8570,N_8038,N_7998);
nor U8571 (N_8571,N_7712,N_7814);
and U8572 (N_8572,N_7974,N_7812);
nor U8573 (N_8573,N_7646,N_7992);
and U8574 (N_8574,N_8037,N_7762);
nand U8575 (N_8575,N_7580,N_8121);
nor U8576 (N_8576,N_7970,N_8123);
nor U8577 (N_8577,N_7768,N_8116);
nor U8578 (N_8578,N_7959,N_7996);
and U8579 (N_8579,N_8124,N_8121);
xnor U8580 (N_8580,N_7797,N_8100);
nand U8581 (N_8581,N_7947,N_7779);
and U8582 (N_8582,N_7758,N_7989);
or U8583 (N_8583,N_7787,N_7994);
nand U8584 (N_8584,N_7696,N_7771);
nand U8585 (N_8585,N_8038,N_7777);
nor U8586 (N_8586,N_7713,N_7820);
nor U8587 (N_8587,N_7776,N_8076);
xnor U8588 (N_8588,N_7661,N_7662);
nand U8589 (N_8589,N_8085,N_7905);
or U8590 (N_8590,N_7839,N_8104);
nand U8591 (N_8591,N_8098,N_7919);
nand U8592 (N_8592,N_7603,N_7645);
or U8593 (N_8593,N_7627,N_7748);
or U8594 (N_8594,N_8112,N_7682);
nand U8595 (N_8595,N_8069,N_7674);
nand U8596 (N_8596,N_7678,N_8007);
xnor U8597 (N_8597,N_8033,N_7862);
or U8598 (N_8598,N_7757,N_8042);
xor U8599 (N_8599,N_7706,N_7848);
and U8600 (N_8600,N_7848,N_7822);
nor U8601 (N_8601,N_7649,N_7988);
xnor U8602 (N_8602,N_7575,N_7911);
nor U8603 (N_8603,N_7605,N_7949);
and U8604 (N_8604,N_8093,N_7685);
nor U8605 (N_8605,N_7996,N_7727);
xnor U8606 (N_8606,N_7810,N_7616);
nor U8607 (N_8607,N_7682,N_7886);
nor U8608 (N_8608,N_7604,N_8019);
nand U8609 (N_8609,N_8122,N_7984);
xnor U8610 (N_8610,N_7602,N_7706);
nor U8611 (N_8611,N_8077,N_7847);
nor U8612 (N_8612,N_7870,N_8045);
xor U8613 (N_8613,N_7550,N_7788);
nand U8614 (N_8614,N_8083,N_7952);
or U8615 (N_8615,N_7948,N_7705);
xor U8616 (N_8616,N_8037,N_7632);
nor U8617 (N_8617,N_7799,N_8100);
xor U8618 (N_8618,N_7785,N_8027);
nand U8619 (N_8619,N_7600,N_7519);
nand U8620 (N_8620,N_8086,N_7617);
nor U8621 (N_8621,N_7944,N_7924);
or U8622 (N_8622,N_7938,N_8036);
and U8623 (N_8623,N_7691,N_7755);
and U8624 (N_8624,N_7655,N_7513);
nor U8625 (N_8625,N_7999,N_7637);
xor U8626 (N_8626,N_7729,N_8107);
and U8627 (N_8627,N_7841,N_8016);
and U8628 (N_8628,N_7939,N_7732);
and U8629 (N_8629,N_7509,N_7899);
or U8630 (N_8630,N_7601,N_8064);
nor U8631 (N_8631,N_8123,N_7720);
and U8632 (N_8632,N_7931,N_7690);
and U8633 (N_8633,N_7745,N_7746);
or U8634 (N_8634,N_7634,N_7857);
or U8635 (N_8635,N_7943,N_8045);
xor U8636 (N_8636,N_7541,N_7668);
and U8637 (N_8637,N_7879,N_7988);
nor U8638 (N_8638,N_8102,N_7835);
xnor U8639 (N_8639,N_7543,N_8093);
nor U8640 (N_8640,N_7640,N_7772);
xnor U8641 (N_8641,N_7893,N_8022);
nand U8642 (N_8642,N_7782,N_7516);
xor U8643 (N_8643,N_8078,N_7853);
xnor U8644 (N_8644,N_7698,N_7558);
xor U8645 (N_8645,N_7788,N_7938);
and U8646 (N_8646,N_8091,N_7676);
and U8647 (N_8647,N_8056,N_7507);
xnor U8648 (N_8648,N_8027,N_7636);
nor U8649 (N_8649,N_7678,N_7584);
nand U8650 (N_8650,N_7879,N_7955);
nor U8651 (N_8651,N_8018,N_8045);
and U8652 (N_8652,N_7911,N_7720);
or U8653 (N_8653,N_7687,N_7647);
nor U8654 (N_8654,N_7949,N_8013);
nand U8655 (N_8655,N_7575,N_7841);
and U8656 (N_8656,N_7971,N_7821);
or U8657 (N_8657,N_8092,N_7749);
and U8658 (N_8658,N_7706,N_7588);
nand U8659 (N_8659,N_7859,N_7786);
and U8660 (N_8660,N_7502,N_7780);
or U8661 (N_8661,N_7628,N_7638);
xnor U8662 (N_8662,N_7565,N_7567);
and U8663 (N_8663,N_7974,N_7734);
and U8664 (N_8664,N_8056,N_8000);
or U8665 (N_8665,N_7950,N_7729);
and U8666 (N_8666,N_7932,N_7593);
and U8667 (N_8667,N_7725,N_7709);
nand U8668 (N_8668,N_8007,N_7971);
or U8669 (N_8669,N_7997,N_7551);
nor U8670 (N_8670,N_7832,N_7569);
xnor U8671 (N_8671,N_7545,N_8013);
and U8672 (N_8672,N_8028,N_7902);
and U8673 (N_8673,N_8100,N_8088);
nor U8674 (N_8674,N_7577,N_8046);
nand U8675 (N_8675,N_7778,N_7804);
nand U8676 (N_8676,N_8045,N_7917);
or U8677 (N_8677,N_8093,N_7618);
nand U8678 (N_8678,N_7539,N_7650);
nand U8679 (N_8679,N_7629,N_7874);
nor U8680 (N_8680,N_8014,N_7695);
nand U8681 (N_8681,N_7861,N_7540);
xor U8682 (N_8682,N_7779,N_7544);
and U8683 (N_8683,N_7939,N_7971);
and U8684 (N_8684,N_7655,N_7772);
or U8685 (N_8685,N_7671,N_7670);
or U8686 (N_8686,N_7875,N_7605);
or U8687 (N_8687,N_8056,N_7804);
nand U8688 (N_8688,N_7966,N_8121);
nand U8689 (N_8689,N_7908,N_7989);
nand U8690 (N_8690,N_7649,N_7762);
xor U8691 (N_8691,N_8042,N_7733);
or U8692 (N_8692,N_7619,N_7777);
or U8693 (N_8693,N_7814,N_8040);
xnor U8694 (N_8694,N_7998,N_8028);
nor U8695 (N_8695,N_7533,N_8076);
or U8696 (N_8696,N_7774,N_7722);
xnor U8697 (N_8697,N_7747,N_7661);
nor U8698 (N_8698,N_7969,N_7866);
xnor U8699 (N_8699,N_7874,N_7860);
nor U8700 (N_8700,N_7864,N_7970);
nor U8701 (N_8701,N_7606,N_8088);
xnor U8702 (N_8702,N_7918,N_7963);
xor U8703 (N_8703,N_7845,N_7607);
and U8704 (N_8704,N_7640,N_7908);
and U8705 (N_8705,N_7702,N_8005);
and U8706 (N_8706,N_7547,N_7651);
and U8707 (N_8707,N_8105,N_7668);
and U8708 (N_8708,N_7699,N_7651);
nor U8709 (N_8709,N_7900,N_7742);
or U8710 (N_8710,N_8012,N_7731);
or U8711 (N_8711,N_7503,N_7901);
xnor U8712 (N_8712,N_7701,N_7716);
xnor U8713 (N_8713,N_7547,N_7618);
and U8714 (N_8714,N_8076,N_7617);
nor U8715 (N_8715,N_8102,N_7903);
nand U8716 (N_8716,N_7935,N_7534);
or U8717 (N_8717,N_8040,N_8002);
nand U8718 (N_8718,N_7586,N_7679);
nor U8719 (N_8719,N_7597,N_7761);
and U8720 (N_8720,N_7601,N_7648);
or U8721 (N_8721,N_7583,N_8025);
xnor U8722 (N_8722,N_8010,N_7985);
nor U8723 (N_8723,N_7502,N_7625);
and U8724 (N_8724,N_8056,N_7559);
nand U8725 (N_8725,N_7580,N_7926);
or U8726 (N_8726,N_8000,N_7589);
nor U8727 (N_8727,N_7537,N_7834);
and U8728 (N_8728,N_8020,N_7545);
and U8729 (N_8729,N_7760,N_7673);
nand U8730 (N_8730,N_7501,N_7656);
nand U8731 (N_8731,N_7848,N_7712);
and U8732 (N_8732,N_7558,N_8123);
and U8733 (N_8733,N_7948,N_7696);
xor U8734 (N_8734,N_7829,N_8123);
xor U8735 (N_8735,N_7641,N_7674);
nand U8736 (N_8736,N_7828,N_8017);
or U8737 (N_8737,N_7698,N_8018);
nor U8738 (N_8738,N_7795,N_7748);
xnor U8739 (N_8739,N_8076,N_7908);
xnor U8740 (N_8740,N_7597,N_7527);
xor U8741 (N_8741,N_7716,N_7656);
or U8742 (N_8742,N_8092,N_8048);
nand U8743 (N_8743,N_8013,N_7700);
or U8744 (N_8744,N_7680,N_7556);
or U8745 (N_8745,N_7955,N_7851);
or U8746 (N_8746,N_7873,N_7976);
or U8747 (N_8747,N_7914,N_8041);
and U8748 (N_8748,N_7706,N_8050);
and U8749 (N_8749,N_7534,N_7647);
or U8750 (N_8750,N_8536,N_8404);
xor U8751 (N_8751,N_8410,N_8181);
or U8752 (N_8752,N_8196,N_8491);
nand U8753 (N_8753,N_8293,N_8364);
and U8754 (N_8754,N_8529,N_8263);
nor U8755 (N_8755,N_8260,N_8299);
or U8756 (N_8756,N_8723,N_8488);
and U8757 (N_8757,N_8317,N_8200);
nand U8758 (N_8758,N_8414,N_8581);
or U8759 (N_8759,N_8674,N_8272);
or U8760 (N_8760,N_8378,N_8199);
nand U8761 (N_8761,N_8172,N_8653);
nor U8762 (N_8762,N_8733,N_8138);
nand U8763 (N_8763,N_8694,N_8238);
nand U8764 (N_8764,N_8718,N_8435);
and U8765 (N_8765,N_8541,N_8441);
nor U8766 (N_8766,N_8585,N_8338);
nand U8767 (N_8767,N_8737,N_8713);
xor U8768 (N_8768,N_8325,N_8192);
or U8769 (N_8769,N_8143,N_8277);
nor U8770 (N_8770,N_8603,N_8337);
nor U8771 (N_8771,N_8382,N_8709);
and U8772 (N_8772,N_8605,N_8542);
xor U8773 (N_8773,N_8180,N_8567);
nor U8774 (N_8774,N_8344,N_8207);
nand U8775 (N_8775,N_8455,N_8463);
and U8776 (N_8776,N_8399,N_8712);
nand U8777 (N_8777,N_8500,N_8150);
xor U8778 (N_8778,N_8482,N_8547);
nand U8779 (N_8779,N_8682,N_8292);
and U8780 (N_8780,N_8310,N_8251);
nor U8781 (N_8781,N_8217,N_8554);
xor U8782 (N_8782,N_8738,N_8628);
nand U8783 (N_8783,N_8162,N_8619);
and U8784 (N_8784,N_8356,N_8522);
nor U8785 (N_8785,N_8357,N_8175);
nor U8786 (N_8786,N_8168,N_8249);
nor U8787 (N_8787,N_8649,N_8692);
nand U8788 (N_8788,N_8584,N_8431);
nor U8789 (N_8789,N_8328,N_8205);
or U8790 (N_8790,N_8691,N_8517);
nand U8791 (N_8791,N_8747,N_8507);
or U8792 (N_8792,N_8160,N_8306);
nor U8793 (N_8793,N_8257,N_8198);
or U8794 (N_8794,N_8373,N_8508);
nand U8795 (N_8795,N_8322,N_8426);
nand U8796 (N_8796,N_8142,N_8631);
or U8797 (N_8797,N_8498,N_8440);
and U8798 (N_8798,N_8565,N_8134);
or U8799 (N_8799,N_8144,N_8155);
or U8800 (N_8800,N_8701,N_8453);
nand U8801 (N_8801,N_8472,N_8475);
xnor U8802 (N_8802,N_8496,N_8719);
and U8803 (N_8803,N_8450,N_8502);
xor U8804 (N_8804,N_8130,N_8485);
nor U8805 (N_8805,N_8135,N_8208);
nand U8806 (N_8806,N_8259,N_8646);
nor U8807 (N_8807,N_8253,N_8244);
nor U8808 (N_8808,N_8185,N_8630);
nand U8809 (N_8809,N_8690,N_8533);
xnor U8810 (N_8810,N_8169,N_8424);
nor U8811 (N_8811,N_8369,N_8609);
xor U8812 (N_8812,N_8131,N_8158);
and U8813 (N_8813,N_8275,N_8477);
nand U8814 (N_8814,N_8710,N_8526);
nand U8815 (N_8815,N_8673,N_8157);
nor U8816 (N_8816,N_8334,N_8367);
and U8817 (N_8817,N_8589,N_8736);
or U8818 (N_8818,N_8599,N_8288);
nor U8819 (N_8819,N_8360,N_8281);
or U8820 (N_8820,N_8551,N_8569);
nand U8821 (N_8821,N_8165,N_8156);
xor U8822 (N_8822,N_8248,N_8315);
or U8823 (N_8823,N_8413,N_8278);
nor U8824 (N_8824,N_8722,N_8643);
nand U8825 (N_8825,N_8451,N_8206);
and U8826 (N_8826,N_8741,N_8375);
and U8827 (N_8827,N_8283,N_8326);
or U8828 (N_8828,N_8678,N_8335);
xnor U8829 (N_8829,N_8311,N_8697);
xor U8830 (N_8830,N_8210,N_8420);
xor U8831 (N_8831,N_8540,N_8389);
nand U8832 (N_8832,N_8327,N_8429);
or U8833 (N_8833,N_8125,N_8647);
xor U8834 (N_8834,N_8242,N_8481);
nand U8835 (N_8835,N_8528,N_8629);
nand U8836 (N_8836,N_8476,N_8298);
nor U8837 (N_8837,N_8724,N_8195);
xor U8838 (N_8838,N_8607,N_8748);
nor U8839 (N_8839,N_8381,N_8717);
and U8840 (N_8840,N_8405,N_8663);
xor U8841 (N_8841,N_8197,N_8323);
or U8842 (N_8842,N_8672,N_8408);
or U8843 (N_8843,N_8398,N_8376);
nand U8844 (N_8844,N_8146,N_8573);
and U8845 (N_8845,N_8139,N_8341);
xnor U8846 (N_8846,N_8417,N_8279);
nand U8847 (N_8847,N_8739,N_8515);
or U8848 (N_8848,N_8560,N_8174);
or U8849 (N_8849,N_8677,N_8329);
nor U8850 (N_8850,N_8368,N_8163);
or U8851 (N_8851,N_8286,N_8432);
or U8852 (N_8852,N_8596,N_8636);
or U8853 (N_8853,N_8583,N_8255);
nand U8854 (N_8854,N_8383,N_8655);
or U8855 (N_8855,N_8610,N_8484);
xor U8856 (N_8856,N_8220,N_8639);
xor U8857 (N_8857,N_8332,N_8204);
or U8858 (N_8858,N_8240,N_8236);
xor U8859 (N_8859,N_8262,N_8266);
and U8860 (N_8860,N_8705,N_8706);
nor U8861 (N_8861,N_8556,N_8428);
nand U8862 (N_8862,N_8421,N_8228);
nor U8863 (N_8863,N_8521,N_8695);
or U8864 (N_8864,N_8203,N_8419);
nand U8865 (N_8865,N_8676,N_8258);
and U8866 (N_8866,N_8330,N_8187);
nor U8867 (N_8867,N_8137,N_8176);
nand U8868 (N_8868,N_8704,N_8557);
and U8869 (N_8869,N_8347,N_8177);
and U8870 (N_8870,N_8478,N_8470);
nor U8871 (N_8871,N_8400,N_8390);
or U8872 (N_8872,N_8633,N_8224);
nand U8873 (N_8873,N_8611,N_8189);
or U8874 (N_8874,N_8422,N_8640);
nand U8875 (N_8875,N_8680,N_8295);
nor U8876 (N_8876,N_8285,N_8297);
nor U8877 (N_8877,N_8708,N_8650);
and U8878 (N_8878,N_8430,N_8675);
nand U8879 (N_8879,N_8743,N_8444);
nand U8880 (N_8880,N_8568,N_8361);
nor U8881 (N_8881,N_8129,N_8576);
nand U8882 (N_8882,N_8634,N_8387);
nor U8883 (N_8883,N_8237,N_8728);
xnor U8884 (N_8884,N_8336,N_8161);
nor U8885 (N_8885,N_8686,N_8648);
nand U8886 (N_8886,N_8303,N_8524);
or U8887 (N_8887,N_8574,N_8553);
nor U8888 (N_8888,N_8726,N_8183);
or U8889 (N_8889,N_8366,N_8469);
xor U8890 (N_8890,N_8651,N_8614);
nand U8891 (N_8891,N_8638,N_8456);
nor U8892 (N_8892,N_8495,N_8664);
nor U8893 (N_8893,N_8370,N_8149);
or U8894 (N_8894,N_8222,N_8182);
xnor U8895 (N_8895,N_8627,N_8462);
nor U8896 (N_8896,N_8159,N_8213);
nor U8897 (N_8897,N_8164,N_8570);
xnor U8898 (N_8898,N_8740,N_8714);
xor U8899 (N_8899,N_8284,N_8537);
nand U8900 (N_8900,N_8391,N_8550);
or U8901 (N_8901,N_8403,N_8667);
xor U8902 (N_8902,N_8394,N_8267);
xor U8903 (N_8903,N_8296,N_8720);
nand U8904 (N_8904,N_8152,N_8438);
or U8905 (N_8905,N_8645,N_8351);
xor U8906 (N_8906,N_8393,N_8269);
and U8907 (N_8907,N_8386,N_8490);
or U8908 (N_8908,N_8506,N_8660);
nor U8909 (N_8909,N_8384,N_8345);
nand U8910 (N_8910,N_8613,N_8186);
xor U8911 (N_8911,N_8302,N_8623);
nand U8912 (N_8912,N_8270,N_8305);
or U8913 (N_8913,N_8577,N_8353);
nand U8914 (N_8914,N_8331,N_8612);
and U8915 (N_8915,N_8178,N_8412);
or U8916 (N_8916,N_8241,N_8621);
or U8917 (N_8917,N_8173,N_8148);
nor U8918 (N_8918,N_8211,N_8590);
or U8919 (N_8919,N_8308,N_8264);
nand U8920 (N_8920,N_8592,N_8730);
nand U8921 (N_8921,N_8616,N_8534);
nor U8922 (N_8922,N_8597,N_8716);
xor U8923 (N_8923,N_8578,N_8601);
nand U8924 (N_8924,N_8711,N_8735);
nand U8925 (N_8925,N_8231,N_8434);
nor U8926 (N_8926,N_8501,N_8666);
or U8927 (N_8927,N_8209,N_8504);
or U8928 (N_8928,N_8497,N_8349);
nand U8929 (N_8929,N_8392,N_8535);
nand U8930 (N_8930,N_8214,N_8698);
or U8931 (N_8931,N_8406,N_8343);
and U8932 (N_8932,N_8519,N_8234);
nand U8933 (N_8933,N_8617,N_8604);
and U8934 (N_8934,N_8523,N_8742);
xnor U8935 (N_8935,N_8509,N_8512);
and U8936 (N_8936,N_8465,N_8564);
and U8937 (N_8937,N_8274,N_8471);
nand U8938 (N_8938,N_8538,N_8670);
nand U8939 (N_8939,N_8731,N_8493);
nor U8940 (N_8940,N_8622,N_8363);
xor U8941 (N_8941,N_8513,N_8586);
nor U8942 (N_8942,N_8215,N_8598);
or U8943 (N_8943,N_8350,N_8447);
and U8944 (N_8944,N_8700,N_8219);
nand U8945 (N_8945,N_8397,N_8665);
or U8946 (N_8946,N_8657,N_8388);
or U8947 (N_8947,N_8626,N_8734);
nand U8948 (N_8948,N_8247,N_8503);
and U8949 (N_8949,N_8683,N_8530);
xnor U8950 (N_8950,N_8184,N_8333);
and U8951 (N_8951,N_8658,N_8532);
and U8952 (N_8952,N_8442,N_8212);
and U8953 (N_8953,N_8562,N_8575);
or U8954 (N_8954,N_8290,N_8494);
and U8955 (N_8955,N_8304,N_8127);
nor U8956 (N_8956,N_8749,N_8687);
and U8957 (N_8957,N_8729,N_8549);
or U8958 (N_8958,N_8246,N_8489);
or U8959 (N_8959,N_8320,N_8457);
nand U8960 (N_8960,N_8216,N_8289);
nor U8961 (N_8961,N_8377,N_8745);
xnor U8962 (N_8962,N_8602,N_8656);
nor U8963 (N_8963,N_8688,N_8443);
or U8964 (N_8964,N_8153,N_8151);
or U8965 (N_8965,N_8715,N_8448);
and U8966 (N_8966,N_8468,N_8167);
nand U8967 (N_8967,N_8136,N_8239);
nor U8968 (N_8968,N_8652,N_8318);
nand U8969 (N_8969,N_8379,N_8202);
xor U8970 (N_8970,N_8354,N_8511);
and U8971 (N_8971,N_8141,N_8510);
and U8972 (N_8972,N_8133,N_8371);
nand U8973 (N_8973,N_8684,N_8271);
nand U8974 (N_8974,N_8254,N_8461);
or U8975 (N_8975,N_8128,N_8637);
xnor U8976 (N_8976,N_8294,N_8746);
or U8977 (N_8977,N_8571,N_8221);
nor U8978 (N_8978,N_8669,N_8473);
and U8979 (N_8979,N_8190,N_8348);
nor U8980 (N_8980,N_8454,N_8486);
or U8981 (N_8981,N_8309,N_8339);
nand U8982 (N_8982,N_8300,N_8668);
or U8983 (N_8983,N_8437,N_8250);
or U8984 (N_8984,N_8395,N_8572);
nand U8985 (N_8985,N_8446,N_8407);
and U8986 (N_8986,N_8411,N_8685);
xor U8987 (N_8987,N_8409,N_8166);
or U8988 (N_8988,N_8595,N_8699);
xor U8989 (N_8989,N_8232,N_8555);
xor U8990 (N_8990,N_8312,N_8268);
nand U8991 (N_8991,N_8233,N_8615);
or U8992 (N_8992,N_8632,N_8702);
xor U8993 (N_8993,N_8539,N_8467);
xnor U8994 (N_8994,N_8452,N_8689);
nor U8995 (N_8995,N_8480,N_8516);
nor U8996 (N_8996,N_8662,N_8544);
and U8997 (N_8997,N_8527,N_8703);
nor U8998 (N_8998,N_8321,N_8641);
or U8999 (N_8999,N_8449,N_8546);
nor U9000 (N_9000,N_8226,N_8126);
xor U9001 (N_9001,N_8342,N_8492);
nand U9002 (N_9002,N_8548,N_8261);
and U9003 (N_9003,N_8280,N_8225);
nor U9004 (N_9004,N_8245,N_8727);
nor U9005 (N_9005,N_8644,N_8433);
xnor U9006 (N_9006,N_8525,N_8307);
nand U9007 (N_9007,N_8732,N_8372);
and U9008 (N_9008,N_8552,N_8252);
xnor U9009 (N_9009,N_8154,N_8600);
or U9010 (N_9010,N_8558,N_8499);
or U9011 (N_9011,N_8721,N_8230);
and U9012 (N_9012,N_8314,N_8561);
nand U9013 (N_9013,N_8460,N_8194);
xor U9014 (N_9014,N_8282,N_8474);
nand U9015 (N_9015,N_8618,N_8380);
nor U9016 (N_9016,N_8579,N_8374);
and U9017 (N_9017,N_8179,N_8520);
nor U9018 (N_9018,N_8436,N_8582);
nand U9019 (N_9019,N_8681,N_8543);
or U9020 (N_9020,N_8188,N_8679);
xor U9021 (N_9021,N_8505,N_8193);
and U9022 (N_9022,N_8243,N_8464);
nor U9023 (N_9023,N_8580,N_8518);
xnor U9024 (N_9024,N_8416,N_8147);
nor U9025 (N_9025,N_8479,N_8223);
and U9026 (N_9026,N_8218,N_8287);
xnor U9027 (N_9027,N_8439,N_8744);
nor U9028 (N_9028,N_8608,N_8587);
nand U9029 (N_9029,N_8362,N_8346);
nor U9030 (N_9030,N_8301,N_8624);
and U9031 (N_9031,N_8593,N_8340);
and U9032 (N_9032,N_8425,N_8171);
nor U9033 (N_9033,N_8466,N_8276);
xnor U9034 (N_9034,N_8358,N_8291);
nor U9035 (N_9035,N_8559,N_8693);
nand U9036 (N_9036,N_8132,N_8707);
nand U9037 (N_9037,N_8659,N_8402);
nor U9038 (N_9038,N_8256,N_8145);
or U9039 (N_9039,N_8313,N_8316);
xor U9040 (N_9040,N_8324,N_8273);
or U9041 (N_9041,N_8642,N_8563);
and U9042 (N_9042,N_8594,N_8227);
nor U9043 (N_9043,N_8396,N_8170);
and U9044 (N_9044,N_8235,N_8696);
and U9045 (N_9045,N_8401,N_8661);
or U9046 (N_9046,N_8427,N_8265);
xnor U9047 (N_9047,N_8365,N_8514);
xor U9048 (N_9048,N_8635,N_8591);
xnor U9049 (N_9049,N_8319,N_8625);
or U9050 (N_9050,N_8352,N_8531);
xor U9051 (N_9051,N_8487,N_8415);
nor U9052 (N_9052,N_8566,N_8671);
xnor U9053 (N_9053,N_8588,N_8355);
or U9054 (N_9054,N_8191,N_8385);
or U9055 (N_9055,N_8620,N_8201);
nor U9056 (N_9056,N_8483,N_8654);
or U9057 (N_9057,N_8445,N_8606);
nor U9058 (N_9058,N_8545,N_8459);
and U9059 (N_9059,N_8418,N_8458);
and U9060 (N_9060,N_8140,N_8229);
or U9061 (N_9061,N_8725,N_8359);
and U9062 (N_9062,N_8423,N_8701);
or U9063 (N_9063,N_8622,N_8721);
nor U9064 (N_9064,N_8340,N_8192);
xnor U9065 (N_9065,N_8425,N_8609);
or U9066 (N_9066,N_8474,N_8736);
nand U9067 (N_9067,N_8567,N_8401);
and U9068 (N_9068,N_8258,N_8177);
and U9069 (N_9069,N_8626,N_8243);
or U9070 (N_9070,N_8708,N_8435);
xnor U9071 (N_9071,N_8136,N_8734);
and U9072 (N_9072,N_8698,N_8341);
or U9073 (N_9073,N_8285,N_8417);
nand U9074 (N_9074,N_8489,N_8717);
nand U9075 (N_9075,N_8463,N_8349);
and U9076 (N_9076,N_8644,N_8556);
xor U9077 (N_9077,N_8592,N_8285);
and U9078 (N_9078,N_8393,N_8675);
and U9079 (N_9079,N_8460,N_8629);
and U9080 (N_9080,N_8430,N_8674);
xnor U9081 (N_9081,N_8499,N_8648);
and U9082 (N_9082,N_8212,N_8491);
xor U9083 (N_9083,N_8641,N_8476);
or U9084 (N_9084,N_8361,N_8424);
or U9085 (N_9085,N_8349,N_8313);
xnor U9086 (N_9086,N_8127,N_8402);
or U9087 (N_9087,N_8349,N_8242);
and U9088 (N_9088,N_8501,N_8137);
xor U9089 (N_9089,N_8607,N_8449);
or U9090 (N_9090,N_8664,N_8423);
xnor U9091 (N_9091,N_8342,N_8506);
nor U9092 (N_9092,N_8528,N_8393);
nor U9093 (N_9093,N_8470,N_8401);
and U9094 (N_9094,N_8270,N_8195);
nand U9095 (N_9095,N_8482,N_8590);
and U9096 (N_9096,N_8415,N_8653);
or U9097 (N_9097,N_8461,N_8449);
nor U9098 (N_9098,N_8205,N_8447);
or U9099 (N_9099,N_8671,N_8409);
nand U9100 (N_9100,N_8355,N_8721);
xnor U9101 (N_9101,N_8347,N_8144);
xor U9102 (N_9102,N_8323,N_8156);
or U9103 (N_9103,N_8394,N_8549);
and U9104 (N_9104,N_8198,N_8457);
nor U9105 (N_9105,N_8461,N_8564);
and U9106 (N_9106,N_8590,N_8688);
nor U9107 (N_9107,N_8195,N_8670);
and U9108 (N_9108,N_8216,N_8721);
nor U9109 (N_9109,N_8238,N_8151);
and U9110 (N_9110,N_8226,N_8616);
nand U9111 (N_9111,N_8333,N_8443);
xnor U9112 (N_9112,N_8211,N_8429);
nand U9113 (N_9113,N_8147,N_8274);
xor U9114 (N_9114,N_8727,N_8633);
nand U9115 (N_9115,N_8277,N_8161);
nand U9116 (N_9116,N_8567,N_8730);
nor U9117 (N_9117,N_8290,N_8150);
nor U9118 (N_9118,N_8610,N_8247);
nor U9119 (N_9119,N_8380,N_8337);
and U9120 (N_9120,N_8414,N_8159);
or U9121 (N_9121,N_8309,N_8576);
nand U9122 (N_9122,N_8338,N_8214);
or U9123 (N_9123,N_8620,N_8268);
nand U9124 (N_9124,N_8513,N_8387);
nor U9125 (N_9125,N_8252,N_8445);
nand U9126 (N_9126,N_8131,N_8428);
and U9127 (N_9127,N_8545,N_8322);
or U9128 (N_9128,N_8438,N_8403);
or U9129 (N_9129,N_8275,N_8614);
nor U9130 (N_9130,N_8271,N_8494);
or U9131 (N_9131,N_8352,N_8610);
and U9132 (N_9132,N_8703,N_8677);
nor U9133 (N_9133,N_8538,N_8706);
or U9134 (N_9134,N_8537,N_8670);
xnor U9135 (N_9135,N_8228,N_8393);
nor U9136 (N_9136,N_8492,N_8670);
nor U9137 (N_9137,N_8217,N_8580);
or U9138 (N_9138,N_8300,N_8596);
xnor U9139 (N_9139,N_8272,N_8140);
or U9140 (N_9140,N_8138,N_8575);
xnor U9141 (N_9141,N_8462,N_8368);
or U9142 (N_9142,N_8227,N_8257);
and U9143 (N_9143,N_8406,N_8259);
nand U9144 (N_9144,N_8372,N_8245);
xnor U9145 (N_9145,N_8598,N_8481);
and U9146 (N_9146,N_8548,N_8435);
nand U9147 (N_9147,N_8685,N_8620);
or U9148 (N_9148,N_8346,N_8593);
nor U9149 (N_9149,N_8629,N_8649);
nand U9150 (N_9150,N_8519,N_8440);
or U9151 (N_9151,N_8637,N_8224);
nor U9152 (N_9152,N_8213,N_8431);
and U9153 (N_9153,N_8500,N_8480);
xor U9154 (N_9154,N_8359,N_8164);
nor U9155 (N_9155,N_8620,N_8295);
xor U9156 (N_9156,N_8446,N_8494);
nor U9157 (N_9157,N_8550,N_8483);
or U9158 (N_9158,N_8532,N_8273);
nor U9159 (N_9159,N_8192,N_8675);
or U9160 (N_9160,N_8142,N_8353);
xnor U9161 (N_9161,N_8179,N_8420);
xnor U9162 (N_9162,N_8258,N_8203);
or U9163 (N_9163,N_8495,N_8463);
and U9164 (N_9164,N_8396,N_8548);
nand U9165 (N_9165,N_8571,N_8268);
and U9166 (N_9166,N_8390,N_8310);
xor U9167 (N_9167,N_8524,N_8481);
xor U9168 (N_9168,N_8745,N_8730);
nand U9169 (N_9169,N_8218,N_8449);
or U9170 (N_9170,N_8697,N_8578);
nand U9171 (N_9171,N_8428,N_8703);
and U9172 (N_9172,N_8598,N_8385);
xor U9173 (N_9173,N_8651,N_8477);
or U9174 (N_9174,N_8709,N_8290);
and U9175 (N_9175,N_8590,N_8410);
or U9176 (N_9176,N_8301,N_8188);
nand U9177 (N_9177,N_8460,N_8310);
or U9178 (N_9178,N_8364,N_8386);
and U9179 (N_9179,N_8735,N_8292);
or U9180 (N_9180,N_8605,N_8652);
xnor U9181 (N_9181,N_8243,N_8376);
nand U9182 (N_9182,N_8405,N_8511);
and U9183 (N_9183,N_8364,N_8216);
and U9184 (N_9184,N_8509,N_8412);
nor U9185 (N_9185,N_8476,N_8740);
nor U9186 (N_9186,N_8173,N_8417);
and U9187 (N_9187,N_8430,N_8152);
nor U9188 (N_9188,N_8357,N_8698);
nor U9189 (N_9189,N_8699,N_8176);
nor U9190 (N_9190,N_8315,N_8301);
or U9191 (N_9191,N_8154,N_8183);
and U9192 (N_9192,N_8179,N_8489);
nor U9193 (N_9193,N_8440,N_8647);
xor U9194 (N_9194,N_8380,N_8666);
and U9195 (N_9195,N_8488,N_8653);
nor U9196 (N_9196,N_8574,N_8558);
nand U9197 (N_9197,N_8332,N_8555);
nor U9198 (N_9198,N_8193,N_8339);
or U9199 (N_9199,N_8675,N_8172);
nor U9200 (N_9200,N_8486,N_8498);
and U9201 (N_9201,N_8280,N_8282);
nand U9202 (N_9202,N_8559,N_8288);
or U9203 (N_9203,N_8519,N_8668);
and U9204 (N_9204,N_8244,N_8582);
and U9205 (N_9205,N_8492,N_8332);
and U9206 (N_9206,N_8485,N_8327);
nor U9207 (N_9207,N_8167,N_8637);
nand U9208 (N_9208,N_8373,N_8258);
and U9209 (N_9209,N_8611,N_8704);
nor U9210 (N_9210,N_8433,N_8710);
xnor U9211 (N_9211,N_8679,N_8213);
nor U9212 (N_9212,N_8550,N_8590);
nand U9213 (N_9213,N_8127,N_8395);
nor U9214 (N_9214,N_8408,N_8478);
and U9215 (N_9215,N_8447,N_8630);
xnor U9216 (N_9216,N_8315,N_8226);
and U9217 (N_9217,N_8266,N_8160);
nand U9218 (N_9218,N_8181,N_8742);
and U9219 (N_9219,N_8387,N_8126);
nand U9220 (N_9220,N_8582,N_8152);
and U9221 (N_9221,N_8455,N_8470);
nand U9222 (N_9222,N_8328,N_8345);
and U9223 (N_9223,N_8690,N_8592);
or U9224 (N_9224,N_8547,N_8306);
nor U9225 (N_9225,N_8507,N_8520);
nand U9226 (N_9226,N_8286,N_8648);
xnor U9227 (N_9227,N_8526,N_8503);
nor U9228 (N_9228,N_8253,N_8575);
and U9229 (N_9229,N_8282,N_8659);
nor U9230 (N_9230,N_8725,N_8334);
nor U9231 (N_9231,N_8258,N_8498);
xnor U9232 (N_9232,N_8676,N_8320);
xnor U9233 (N_9233,N_8675,N_8520);
nand U9234 (N_9234,N_8223,N_8536);
nand U9235 (N_9235,N_8616,N_8637);
nor U9236 (N_9236,N_8466,N_8294);
xor U9237 (N_9237,N_8689,N_8161);
nand U9238 (N_9238,N_8324,N_8177);
nor U9239 (N_9239,N_8649,N_8227);
nor U9240 (N_9240,N_8632,N_8676);
nand U9241 (N_9241,N_8611,N_8352);
nand U9242 (N_9242,N_8493,N_8431);
nor U9243 (N_9243,N_8625,N_8156);
nand U9244 (N_9244,N_8496,N_8422);
xnor U9245 (N_9245,N_8621,N_8399);
or U9246 (N_9246,N_8129,N_8231);
nor U9247 (N_9247,N_8516,N_8156);
xnor U9248 (N_9248,N_8345,N_8645);
nand U9249 (N_9249,N_8153,N_8634);
nor U9250 (N_9250,N_8703,N_8722);
xnor U9251 (N_9251,N_8452,N_8467);
nor U9252 (N_9252,N_8356,N_8709);
xor U9253 (N_9253,N_8442,N_8624);
and U9254 (N_9254,N_8282,N_8157);
and U9255 (N_9255,N_8347,N_8594);
nand U9256 (N_9256,N_8378,N_8666);
nand U9257 (N_9257,N_8450,N_8166);
or U9258 (N_9258,N_8446,N_8677);
nand U9259 (N_9259,N_8485,N_8577);
nand U9260 (N_9260,N_8685,N_8512);
xor U9261 (N_9261,N_8342,N_8397);
xor U9262 (N_9262,N_8507,N_8191);
xnor U9263 (N_9263,N_8704,N_8601);
and U9264 (N_9264,N_8638,N_8214);
or U9265 (N_9265,N_8300,N_8505);
and U9266 (N_9266,N_8324,N_8199);
xor U9267 (N_9267,N_8312,N_8487);
nand U9268 (N_9268,N_8699,N_8653);
xor U9269 (N_9269,N_8552,N_8432);
or U9270 (N_9270,N_8508,N_8532);
xnor U9271 (N_9271,N_8613,N_8340);
or U9272 (N_9272,N_8605,N_8215);
nand U9273 (N_9273,N_8194,N_8739);
xnor U9274 (N_9274,N_8399,N_8216);
or U9275 (N_9275,N_8701,N_8671);
nor U9276 (N_9276,N_8614,N_8372);
xnor U9277 (N_9277,N_8322,N_8148);
nand U9278 (N_9278,N_8492,N_8641);
xnor U9279 (N_9279,N_8483,N_8281);
nand U9280 (N_9280,N_8521,N_8509);
and U9281 (N_9281,N_8714,N_8135);
nor U9282 (N_9282,N_8203,N_8644);
xnor U9283 (N_9283,N_8340,N_8171);
xor U9284 (N_9284,N_8605,N_8536);
nand U9285 (N_9285,N_8331,N_8262);
or U9286 (N_9286,N_8505,N_8576);
or U9287 (N_9287,N_8526,N_8443);
xnor U9288 (N_9288,N_8347,N_8161);
nand U9289 (N_9289,N_8396,N_8359);
and U9290 (N_9290,N_8714,N_8323);
and U9291 (N_9291,N_8513,N_8348);
xor U9292 (N_9292,N_8358,N_8158);
xnor U9293 (N_9293,N_8731,N_8351);
nand U9294 (N_9294,N_8371,N_8295);
or U9295 (N_9295,N_8711,N_8434);
xor U9296 (N_9296,N_8464,N_8282);
xnor U9297 (N_9297,N_8630,N_8694);
xnor U9298 (N_9298,N_8233,N_8141);
or U9299 (N_9299,N_8558,N_8336);
xnor U9300 (N_9300,N_8454,N_8378);
xnor U9301 (N_9301,N_8693,N_8499);
and U9302 (N_9302,N_8669,N_8320);
and U9303 (N_9303,N_8732,N_8670);
or U9304 (N_9304,N_8453,N_8740);
or U9305 (N_9305,N_8609,N_8453);
nor U9306 (N_9306,N_8514,N_8579);
and U9307 (N_9307,N_8517,N_8251);
or U9308 (N_9308,N_8647,N_8354);
nor U9309 (N_9309,N_8213,N_8412);
or U9310 (N_9310,N_8539,N_8544);
nor U9311 (N_9311,N_8446,N_8666);
and U9312 (N_9312,N_8460,N_8381);
or U9313 (N_9313,N_8633,N_8477);
nor U9314 (N_9314,N_8703,N_8384);
or U9315 (N_9315,N_8163,N_8205);
or U9316 (N_9316,N_8207,N_8415);
nand U9317 (N_9317,N_8656,N_8134);
and U9318 (N_9318,N_8529,N_8741);
and U9319 (N_9319,N_8645,N_8379);
nand U9320 (N_9320,N_8368,N_8281);
nor U9321 (N_9321,N_8295,N_8553);
nand U9322 (N_9322,N_8676,N_8721);
xor U9323 (N_9323,N_8232,N_8155);
nand U9324 (N_9324,N_8734,N_8325);
nand U9325 (N_9325,N_8433,N_8604);
xor U9326 (N_9326,N_8178,N_8537);
and U9327 (N_9327,N_8709,N_8598);
xnor U9328 (N_9328,N_8589,N_8161);
nand U9329 (N_9329,N_8655,N_8712);
nor U9330 (N_9330,N_8630,N_8679);
nor U9331 (N_9331,N_8271,N_8707);
nand U9332 (N_9332,N_8489,N_8279);
xor U9333 (N_9333,N_8433,N_8298);
nor U9334 (N_9334,N_8463,N_8297);
or U9335 (N_9335,N_8462,N_8535);
or U9336 (N_9336,N_8582,N_8161);
xnor U9337 (N_9337,N_8341,N_8538);
or U9338 (N_9338,N_8520,N_8213);
nand U9339 (N_9339,N_8534,N_8705);
and U9340 (N_9340,N_8641,N_8621);
and U9341 (N_9341,N_8325,N_8234);
or U9342 (N_9342,N_8441,N_8405);
xnor U9343 (N_9343,N_8714,N_8672);
xor U9344 (N_9344,N_8138,N_8477);
or U9345 (N_9345,N_8521,N_8157);
xor U9346 (N_9346,N_8539,N_8729);
nor U9347 (N_9347,N_8270,N_8400);
and U9348 (N_9348,N_8579,N_8441);
and U9349 (N_9349,N_8726,N_8462);
nor U9350 (N_9350,N_8705,N_8531);
and U9351 (N_9351,N_8338,N_8705);
nor U9352 (N_9352,N_8248,N_8519);
nor U9353 (N_9353,N_8717,N_8169);
or U9354 (N_9354,N_8425,N_8602);
and U9355 (N_9355,N_8436,N_8345);
and U9356 (N_9356,N_8613,N_8701);
nor U9357 (N_9357,N_8260,N_8589);
nand U9358 (N_9358,N_8129,N_8193);
nor U9359 (N_9359,N_8493,N_8720);
or U9360 (N_9360,N_8588,N_8143);
or U9361 (N_9361,N_8173,N_8286);
nor U9362 (N_9362,N_8501,N_8512);
nand U9363 (N_9363,N_8618,N_8644);
xnor U9364 (N_9364,N_8690,N_8229);
and U9365 (N_9365,N_8613,N_8732);
nor U9366 (N_9366,N_8620,N_8173);
nand U9367 (N_9367,N_8658,N_8461);
and U9368 (N_9368,N_8512,N_8137);
xnor U9369 (N_9369,N_8730,N_8235);
nand U9370 (N_9370,N_8522,N_8336);
and U9371 (N_9371,N_8197,N_8706);
and U9372 (N_9372,N_8639,N_8412);
or U9373 (N_9373,N_8650,N_8701);
nand U9374 (N_9374,N_8254,N_8420);
and U9375 (N_9375,N_8750,N_9335);
or U9376 (N_9376,N_8804,N_9372);
or U9377 (N_9377,N_8798,N_9340);
nand U9378 (N_9378,N_8987,N_8825);
and U9379 (N_9379,N_9319,N_9235);
xnor U9380 (N_9380,N_9238,N_8945);
or U9381 (N_9381,N_9345,N_9178);
and U9382 (N_9382,N_9118,N_8778);
and U9383 (N_9383,N_9143,N_8848);
and U9384 (N_9384,N_9146,N_9069);
or U9385 (N_9385,N_8950,N_9149);
xnor U9386 (N_9386,N_8972,N_9274);
nor U9387 (N_9387,N_8874,N_8787);
nand U9388 (N_9388,N_9236,N_8940);
and U9389 (N_9389,N_9194,N_9242);
and U9390 (N_9390,N_8948,N_9239);
and U9391 (N_9391,N_8754,N_8819);
nor U9392 (N_9392,N_8762,N_9190);
xor U9393 (N_9393,N_8860,N_9021);
and U9394 (N_9394,N_9344,N_9222);
or U9395 (N_9395,N_9036,N_8790);
or U9396 (N_9396,N_9187,N_8974);
and U9397 (N_9397,N_9373,N_9042);
or U9398 (N_9398,N_9070,N_9191);
nand U9399 (N_9399,N_9096,N_8780);
or U9400 (N_9400,N_8980,N_8912);
xnor U9401 (N_9401,N_8801,N_8997);
nand U9402 (N_9402,N_8908,N_8800);
and U9403 (N_9403,N_8993,N_9362);
xor U9404 (N_9404,N_8865,N_9005);
nor U9405 (N_9405,N_8952,N_9243);
and U9406 (N_9406,N_8872,N_8766);
nand U9407 (N_9407,N_9025,N_9010);
or U9408 (N_9408,N_9234,N_8994);
xnor U9409 (N_9409,N_9091,N_9278);
nor U9410 (N_9410,N_9293,N_9034);
xnor U9411 (N_9411,N_8978,N_9364);
or U9412 (N_9412,N_9229,N_8861);
or U9413 (N_9413,N_8836,N_8967);
nand U9414 (N_9414,N_8870,N_9333);
nand U9415 (N_9415,N_9285,N_9150);
or U9416 (N_9416,N_9246,N_9268);
nand U9417 (N_9417,N_8965,N_9189);
and U9418 (N_9418,N_8977,N_9126);
nor U9419 (N_9419,N_9291,N_9078);
nand U9420 (N_9420,N_9352,N_9286);
or U9421 (N_9421,N_9108,N_9103);
and U9422 (N_9422,N_8853,N_8964);
and U9423 (N_9423,N_9053,N_8768);
nand U9424 (N_9424,N_9316,N_8898);
or U9425 (N_9425,N_9113,N_8820);
and U9426 (N_9426,N_9253,N_9092);
and U9427 (N_9427,N_8923,N_9047);
or U9428 (N_9428,N_8802,N_8845);
nor U9429 (N_9429,N_8827,N_9035);
or U9430 (N_9430,N_9098,N_9301);
nand U9431 (N_9431,N_8932,N_8863);
xor U9432 (N_9432,N_9367,N_8990);
nor U9433 (N_9433,N_8953,N_9244);
and U9434 (N_9434,N_8823,N_9199);
xnor U9435 (N_9435,N_9241,N_8770);
nand U9436 (N_9436,N_9101,N_8777);
or U9437 (N_9437,N_9240,N_8811);
and U9438 (N_9438,N_9084,N_9130);
nor U9439 (N_9439,N_9022,N_9365);
or U9440 (N_9440,N_8913,N_9224);
or U9441 (N_9441,N_9266,N_9120);
or U9442 (N_9442,N_9007,N_9267);
nor U9443 (N_9443,N_8869,N_9147);
xor U9444 (N_9444,N_9115,N_8864);
nand U9445 (N_9445,N_8946,N_9009);
and U9446 (N_9446,N_8979,N_9139);
nand U9447 (N_9447,N_8831,N_8951);
nand U9448 (N_9448,N_8833,N_9183);
nor U9449 (N_9449,N_9024,N_8917);
nand U9450 (N_9450,N_9000,N_9250);
nor U9451 (N_9451,N_9262,N_9251);
nor U9452 (N_9452,N_8854,N_8789);
and U9453 (N_9453,N_9175,N_8909);
or U9454 (N_9454,N_9231,N_8839);
or U9455 (N_9455,N_9326,N_9029);
xnor U9456 (N_9456,N_9075,N_9201);
or U9457 (N_9457,N_9046,N_9044);
nor U9458 (N_9458,N_9245,N_8887);
nor U9459 (N_9459,N_9325,N_8984);
or U9460 (N_9460,N_9346,N_9052);
nand U9461 (N_9461,N_8807,N_9309);
and U9462 (N_9462,N_9014,N_8813);
or U9463 (N_9463,N_9017,N_8973);
xnor U9464 (N_9464,N_8910,N_8935);
and U9465 (N_9465,N_9343,N_9271);
nor U9466 (N_9466,N_8775,N_9356);
nor U9467 (N_9467,N_9225,N_8764);
nand U9468 (N_9468,N_8796,N_9060);
nor U9469 (N_9469,N_9073,N_9077);
or U9470 (N_9470,N_8779,N_8765);
nand U9471 (N_9471,N_9003,N_9230);
nor U9472 (N_9472,N_9002,N_8834);
xnor U9473 (N_9473,N_9166,N_8934);
xor U9474 (N_9474,N_8937,N_8850);
nand U9475 (N_9475,N_9181,N_9314);
and U9476 (N_9476,N_9083,N_8999);
nor U9477 (N_9477,N_8817,N_8877);
nor U9478 (N_9478,N_9051,N_8954);
xor U9479 (N_9479,N_9311,N_9121);
or U9480 (N_9480,N_9031,N_9127);
and U9481 (N_9481,N_9341,N_9111);
or U9482 (N_9482,N_9237,N_8989);
xnor U9483 (N_9483,N_9257,N_8982);
or U9484 (N_9484,N_8772,N_9059);
or U9485 (N_9485,N_9369,N_9023);
or U9486 (N_9486,N_8806,N_9152);
and U9487 (N_9487,N_8992,N_9159);
xnor U9488 (N_9488,N_8856,N_9217);
or U9489 (N_9489,N_8810,N_9287);
nand U9490 (N_9490,N_8962,N_9303);
and U9491 (N_9491,N_9158,N_9312);
xnor U9492 (N_9492,N_8891,N_8929);
xor U9493 (N_9493,N_8838,N_9028);
nand U9494 (N_9494,N_8963,N_9049);
nor U9495 (N_9495,N_9330,N_9221);
and U9496 (N_9496,N_9161,N_8767);
or U9497 (N_9497,N_9012,N_8896);
nand U9498 (N_9498,N_9145,N_9097);
and U9499 (N_9499,N_8842,N_9058);
xor U9500 (N_9500,N_8921,N_8981);
xnor U9501 (N_9501,N_9013,N_9361);
or U9502 (N_9502,N_8835,N_9085);
nor U9503 (N_9503,N_8915,N_8995);
nand U9504 (N_9504,N_9313,N_9180);
or U9505 (N_9505,N_9131,N_9068);
nor U9506 (N_9506,N_8841,N_9354);
nand U9507 (N_9507,N_9299,N_8895);
xnor U9508 (N_9508,N_9144,N_8941);
xor U9509 (N_9509,N_8924,N_8855);
or U9510 (N_9510,N_9305,N_8957);
nand U9511 (N_9511,N_8983,N_8824);
nor U9512 (N_9512,N_9254,N_8873);
or U9513 (N_9513,N_8881,N_9102);
nor U9514 (N_9514,N_8914,N_9055);
and U9515 (N_9515,N_9184,N_9197);
nand U9516 (N_9516,N_9215,N_8866);
nand U9517 (N_9517,N_8821,N_8944);
nor U9518 (N_9518,N_9104,N_8829);
or U9519 (N_9519,N_9290,N_9050);
nand U9520 (N_9520,N_9202,N_9196);
xor U9521 (N_9521,N_9247,N_8828);
nor U9522 (N_9522,N_8816,N_9348);
or U9523 (N_9523,N_9106,N_9258);
or U9524 (N_9524,N_9216,N_8927);
xor U9525 (N_9525,N_8903,N_8902);
or U9526 (N_9526,N_8851,N_8920);
nand U9527 (N_9527,N_9327,N_9289);
xor U9528 (N_9528,N_9032,N_8774);
and U9529 (N_9529,N_8793,N_9255);
and U9530 (N_9530,N_9094,N_8961);
xnor U9531 (N_9531,N_8959,N_9037);
and U9532 (N_9532,N_8846,N_8878);
nand U9533 (N_9533,N_8859,N_9163);
xnor U9534 (N_9534,N_8760,N_9043);
xnor U9535 (N_9535,N_8947,N_9192);
and U9536 (N_9536,N_9208,N_9125);
nand U9537 (N_9537,N_9321,N_8773);
xor U9538 (N_9538,N_9228,N_8892);
and U9539 (N_9539,N_8875,N_9347);
xnor U9540 (N_9540,N_9071,N_8968);
and U9541 (N_9541,N_8784,N_9209);
nor U9542 (N_9542,N_8938,N_9095);
and U9543 (N_9543,N_9318,N_9363);
xnor U9544 (N_9544,N_8782,N_9156);
nor U9545 (N_9545,N_8985,N_8925);
nand U9546 (N_9546,N_8847,N_9076);
nand U9547 (N_9547,N_8751,N_9038);
nand U9548 (N_9548,N_9116,N_9086);
nand U9549 (N_9549,N_9020,N_9162);
nand U9550 (N_9550,N_9370,N_9026);
or U9551 (N_9551,N_8966,N_9105);
or U9552 (N_9552,N_8971,N_9066);
nor U9553 (N_9553,N_9054,N_9355);
xor U9554 (N_9554,N_9089,N_8876);
nand U9555 (N_9555,N_9294,N_9336);
nor U9556 (N_9556,N_8969,N_9160);
nand U9557 (N_9557,N_9317,N_9357);
or U9558 (N_9558,N_9117,N_9211);
or U9559 (N_9559,N_9315,N_9082);
xor U9560 (N_9560,N_9272,N_9207);
or U9561 (N_9561,N_8803,N_8857);
and U9562 (N_9562,N_9114,N_9081);
and U9563 (N_9563,N_9174,N_9329);
nor U9564 (N_9564,N_9323,N_8926);
and U9565 (N_9565,N_9281,N_9273);
xnor U9566 (N_9566,N_9223,N_9310);
or U9567 (N_9567,N_9334,N_9008);
or U9568 (N_9568,N_9136,N_9132);
xor U9569 (N_9569,N_8832,N_8757);
nand U9570 (N_9570,N_9033,N_9172);
nand U9571 (N_9571,N_8988,N_9109);
nor U9572 (N_9572,N_9128,N_8852);
nor U9573 (N_9573,N_8931,N_8970);
nand U9574 (N_9574,N_8919,N_9358);
and U9575 (N_9575,N_9320,N_9260);
nand U9576 (N_9576,N_8916,N_8905);
or U9577 (N_9577,N_9133,N_8840);
nand U9578 (N_9578,N_9001,N_9041);
and U9579 (N_9579,N_9203,N_9186);
and U9580 (N_9580,N_8867,N_9107);
xor U9581 (N_9581,N_9185,N_8880);
nor U9582 (N_9582,N_9135,N_9252);
nand U9583 (N_9583,N_8911,N_8830);
xnor U9584 (N_9584,N_9212,N_9045);
nand U9585 (N_9585,N_9308,N_8862);
and U9586 (N_9586,N_8928,N_8960);
xor U9587 (N_9587,N_9368,N_9337);
nand U9588 (N_9588,N_9018,N_9100);
xnor U9589 (N_9589,N_8756,N_9112);
or U9590 (N_9590,N_8794,N_9155);
xnor U9591 (N_9591,N_9366,N_8771);
nand U9592 (N_9592,N_9302,N_9263);
and U9593 (N_9593,N_8888,N_9173);
or U9594 (N_9594,N_9322,N_9176);
nor U9595 (N_9595,N_9204,N_9332);
nand U9596 (N_9596,N_8890,N_9064);
nor U9597 (N_9597,N_8998,N_9195);
nand U9598 (N_9598,N_8792,N_9342);
or U9599 (N_9599,N_9275,N_9062);
xnor U9600 (N_9600,N_9205,N_9137);
nor U9601 (N_9601,N_8955,N_9259);
nand U9602 (N_9602,N_9122,N_9295);
or U9603 (N_9603,N_9298,N_8812);
nand U9604 (N_9604,N_9288,N_9016);
xor U9605 (N_9605,N_9218,N_8844);
or U9606 (N_9606,N_9048,N_9349);
nor U9607 (N_9607,N_9165,N_8930);
and U9608 (N_9608,N_9249,N_8759);
and U9609 (N_9609,N_8904,N_9350);
xor U9610 (N_9610,N_8882,N_9256);
nor U9611 (N_9611,N_8879,N_9072);
and U9612 (N_9612,N_9200,N_8939);
xor U9613 (N_9613,N_9093,N_9277);
xnor U9614 (N_9614,N_9276,N_9219);
nand U9615 (N_9615,N_8906,N_8885);
xnor U9616 (N_9616,N_9129,N_9269);
xnor U9617 (N_9617,N_8752,N_9088);
xnor U9618 (N_9618,N_9142,N_9039);
or U9619 (N_9619,N_8991,N_9119);
xnor U9620 (N_9620,N_9099,N_9074);
or U9621 (N_9621,N_9168,N_8897);
and U9622 (N_9622,N_9063,N_8818);
nor U9623 (N_9623,N_8901,N_9040);
or U9624 (N_9624,N_9374,N_9177);
xnor U9625 (N_9625,N_8769,N_8858);
and U9626 (N_9626,N_8849,N_8871);
nor U9627 (N_9627,N_8797,N_9154);
and U9628 (N_9628,N_9011,N_8884);
or U9629 (N_9629,N_9124,N_8761);
nand U9630 (N_9630,N_9198,N_9304);
nand U9631 (N_9631,N_9331,N_9151);
nor U9632 (N_9632,N_9153,N_9090);
and U9633 (N_9633,N_9261,N_9280);
nor U9634 (N_9634,N_8758,N_8889);
nor U9635 (N_9635,N_8837,N_9351);
and U9636 (N_9636,N_8763,N_9164);
nor U9637 (N_9637,N_9087,N_8907);
xor U9638 (N_9638,N_9169,N_8814);
and U9639 (N_9639,N_9080,N_9179);
or U9640 (N_9640,N_9248,N_9265);
nand U9641 (N_9641,N_8788,N_8868);
xnor U9642 (N_9642,N_9193,N_8799);
and U9643 (N_9643,N_8976,N_8886);
or U9644 (N_9644,N_8996,N_8781);
nor U9645 (N_9645,N_8791,N_8894);
and U9646 (N_9646,N_9210,N_9338);
nand U9647 (N_9647,N_9353,N_9171);
xor U9648 (N_9648,N_8942,N_8805);
and U9649 (N_9649,N_8822,N_9057);
nand U9650 (N_9650,N_9027,N_8786);
or U9651 (N_9651,N_9188,N_8776);
nor U9652 (N_9652,N_8808,N_9270);
nor U9653 (N_9653,N_8949,N_9015);
nand U9654 (N_9654,N_8943,N_9170);
nor U9655 (N_9655,N_9232,N_8893);
and U9656 (N_9656,N_9056,N_9157);
xor U9657 (N_9657,N_8986,N_9148);
nor U9658 (N_9658,N_8783,N_9371);
and U9659 (N_9659,N_9226,N_9138);
or U9660 (N_9660,N_8899,N_8815);
and U9661 (N_9661,N_9067,N_9339);
and U9662 (N_9662,N_9182,N_9030);
nor U9663 (N_9663,N_8753,N_9360);
nand U9664 (N_9664,N_9167,N_9227);
and U9665 (N_9665,N_9282,N_9019);
nor U9666 (N_9666,N_9359,N_9213);
nand U9667 (N_9667,N_9297,N_9283);
or U9668 (N_9668,N_9134,N_9061);
nor U9669 (N_9669,N_8975,N_9110);
or U9670 (N_9670,N_9065,N_9220);
nor U9671 (N_9671,N_9300,N_9123);
and U9672 (N_9672,N_9214,N_8826);
and U9673 (N_9673,N_9324,N_9264);
nand U9674 (N_9674,N_9140,N_8755);
xor U9675 (N_9675,N_9306,N_8883);
and U9676 (N_9676,N_8843,N_8956);
xor U9677 (N_9677,N_8809,N_9006);
nand U9678 (N_9678,N_9307,N_9284);
nand U9679 (N_9679,N_9233,N_8795);
nand U9680 (N_9680,N_9279,N_9296);
nor U9681 (N_9681,N_9004,N_9328);
nor U9682 (N_9682,N_8900,N_8933);
nand U9683 (N_9683,N_9079,N_9141);
xor U9684 (N_9684,N_8918,N_9206);
and U9685 (N_9685,N_9292,N_8785);
and U9686 (N_9686,N_8922,N_8958);
nand U9687 (N_9687,N_8936,N_8811);
nand U9688 (N_9688,N_9134,N_9211);
or U9689 (N_9689,N_9108,N_9244);
nor U9690 (N_9690,N_9037,N_8765);
nand U9691 (N_9691,N_8760,N_9022);
nor U9692 (N_9692,N_8846,N_9044);
nor U9693 (N_9693,N_9026,N_8903);
and U9694 (N_9694,N_8945,N_8965);
xor U9695 (N_9695,N_9072,N_8935);
and U9696 (N_9696,N_9374,N_8866);
or U9697 (N_9697,N_8848,N_8922);
nand U9698 (N_9698,N_8914,N_9044);
nor U9699 (N_9699,N_9196,N_9045);
nand U9700 (N_9700,N_9019,N_8939);
or U9701 (N_9701,N_9185,N_9173);
or U9702 (N_9702,N_9040,N_8911);
or U9703 (N_9703,N_8881,N_9099);
and U9704 (N_9704,N_8942,N_9184);
or U9705 (N_9705,N_9208,N_9340);
nor U9706 (N_9706,N_9341,N_9373);
and U9707 (N_9707,N_9000,N_8759);
nor U9708 (N_9708,N_9211,N_9270);
and U9709 (N_9709,N_9001,N_9303);
nor U9710 (N_9710,N_9126,N_9145);
nor U9711 (N_9711,N_8991,N_9342);
nand U9712 (N_9712,N_8912,N_9323);
or U9713 (N_9713,N_9153,N_8999);
or U9714 (N_9714,N_9372,N_8759);
xor U9715 (N_9715,N_8865,N_9058);
nor U9716 (N_9716,N_9275,N_9329);
xor U9717 (N_9717,N_8925,N_9219);
or U9718 (N_9718,N_9182,N_8768);
nor U9719 (N_9719,N_9228,N_8839);
or U9720 (N_9720,N_9296,N_8955);
nor U9721 (N_9721,N_8770,N_8915);
and U9722 (N_9722,N_9324,N_8801);
or U9723 (N_9723,N_9038,N_9049);
nand U9724 (N_9724,N_8799,N_8864);
nand U9725 (N_9725,N_9176,N_9224);
and U9726 (N_9726,N_9080,N_9324);
or U9727 (N_9727,N_8880,N_8761);
and U9728 (N_9728,N_8887,N_8974);
or U9729 (N_9729,N_8934,N_8994);
or U9730 (N_9730,N_9097,N_9176);
nand U9731 (N_9731,N_9162,N_9103);
nand U9732 (N_9732,N_9301,N_9189);
and U9733 (N_9733,N_8764,N_9200);
and U9734 (N_9734,N_9188,N_8848);
nand U9735 (N_9735,N_9007,N_8911);
nor U9736 (N_9736,N_9055,N_9138);
xor U9737 (N_9737,N_9165,N_9273);
or U9738 (N_9738,N_8857,N_9038);
and U9739 (N_9739,N_8875,N_8958);
and U9740 (N_9740,N_8868,N_9349);
nor U9741 (N_9741,N_9268,N_9016);
nor U9742 (N_9742,N_9140,N_9171);
xor U9743 (N_9743,N_8865,N_8790);
nand U9744 (N_9744,N_8856,N_9350);
xor U9745 (N_9745,N_9037,N_9235);
and U9746 (N_9746,N_9013,N_8852);
nand U9747 (N_9747,N_9161,N_9309);
or U9748 (N_9748,N_8847,N_9246);
or U9749 (N_9749,N_8996,N_8883);
xor U9750 (N_9750,N_8976,N_9327);
xnor U9751 (N_9751,N_8869,N_9207);
nor U9752 (N_9752,N_9058,N_9029);
nand U9753 (N_9753,N_8768,N_9003);
and U9754 (N_9754,N_8959,N_8812);
and U9755 (N_9755,N_9296,N_9167);
and U9756 (N_9756,N_8858,N_8916);
or U9757 (N_9757,N_9164,N_9350);
xor U9758 (N_9758,N_9202,N_8946);
and U9759 (N_9759,N_8811,N_8891);
and U9760 (N_9760,N_9305,N_8876);
and U9761 (N_9761,N_9117,N_9076);
nand U9762 (N_9762,N_8813,N_8909);
and U9763 (N_9763,N_8865,N_9133);
and U9764 (N_9764,N_9104,N_8910);
nor U9765 (N_9765,N_9093,N_9260);
and U9766 (N_9766,N_9172,N_8997);
xor U9767 (N_9767,N_8755,N_9175);
nand U9768 (N_9768,N_9188,N_8984);
xor U9769 (N_9769,N_9125,N_8859);
xnor U9770 (N_9770,N_8914,N_8752);
and U9771 (N_9771,N_9020,N_9073);
or U9772 (N_9772,N_9346,N_9015);
or U9773 (N_9773,N_9129,N_8978);
and U9774 (N_9774,N_9128,N_9218);
or U9775 (N_9775,N_9047,N_8815);
or U9776 (N_9776,N_8833,N_9257);
and U9777 (N_9777,N_9298,N_8939);
and U9778 (N_9778,N_8881,N_9274);
nand U9779 (N_9779,N_9103,N_8799);
and U9780 (N_9780,N_9076,N_9180);
nand U9781 (N_9781,N_9101,N_9029);
and U9782 (N_9782,N_9367,N_8960);
xnor U9783 (N_9783,N_8871,N_9135);
xor U9784 (N_9784,N_9302,N_9112);
and U9785 (N_9785,N_9242,N_9243);
nor U9786 (N_9786,N_8756,N_9272);
and U9787 (N_9787,N_9215,N_9248);
nor U9788 (N_9788,N_8917,N_8914);
nand U9789 (N_9789,N_8969,N_8909);
or U9790 (N_9790,N_9315,N_9026);
xnor U9791 (N_9791,N_9131,N_8923);
or U9792 (N_9792,N_8790,N_8998);
or U9793 (N_9793,N_9045,N_8755);
xnor U9794 (N_9794,N_9285,N_9340);
nor U9795 (N_9795,N_9060,N_9234);
nor U9796 (N_9796,N_9289,N_9315);
nor U9797 (N_9797,N_9245,N_9221);
and U9798 (N_9798,N_9192,N_9109);
xor U9799 (N_9799,N_9258,N_8778);
nor U9800 (N_9800,N_8839,N_9202);
and U9801 (N_9801,N_8828,N_9313);
nor U9802 (N_9802,N_9019,N_8965);
and U9803 (N_9803,N_9013,N_9149);
xor U9804 (N_9804,N_9286,N_9081);
and U9805 (N_9805,N_8753,N_8938);
nor U9806 (N_9806,N_8870,N_8779);
nand U9807 (N_9807,N_9076,N_8785);
or U9808 (N_9808,N_8999,N_9349);
xnor U9809 (N_9809,N_8796,N_8920);
nor U9810 (N_9810,N_9298,N_8752);
and U9811 (N_9811,N_9331,N_8929);
nand U9812 (N_9812,N_9293,N_9187);
nor U9813 (N_9813,N_8963,N_8913);
or U9814 (N_9814,N_9076,N_9208);
xor U9815 (N_9815,N_8751,N_8774);
and U9816 (N_9816,N_8896,N_9072);
and U9817 (N_9817,N_9056,N_9081);
nand U9818 (N_9818,N_8926,N_8970);
or U9819 (N_9819,N_9238,N_9373);
nand U9820 (N_9820,N_9358,N_9328);
or U9821 (N_9821,N_9295,N_9300);
nand U9822 (N_9822,N_8853,N_8956);
nor U9823 (N_9823,N_9162,N_8894);
and U9824 (N_9824,N_8962,N_9168);
nand U9825 (N_9825,N_8797,N_9027);
nand U9826 (N_9826,N_8871,N_9213);
or U9827 (N_9827,N_9111,N_9055);
xor U9828 (N_9828,N_9092,N_9358);
or U9829 (N_9829,N_8980,N_9239);
nor U9830 (N_9830,N_8917,N_8782);
nor U9831 (N_9831,N_8841,N_8885);
nand U9832 (N_9832,N_8976,N_8798);
xor U9833 (N_9833,N_9183,N_8904);
nand U9834 (N_9834,N_9099,N_8965);
and U9835 (N_9835,N_9025,N_8891);
nand U9836 (N_9836,N_9026,N_8800);
xor U9837 (N_9837,N_9184,N_9019);
nor U9838 (N_9838,N_9251,N_9090);
nand U9839 (N_9839,N_9024,N_9105);
nor U9840 (N_9840,N_9024,N_9225);
xnor U9841 (N_9841,N_9264,N_9195);
and U9842 (N_9842,N_8912,N_9284);
or U9843 (N_9843,N_8984,N_9305);
or U9844 (N_9844,N_9079,N_8839);
nand U9845 (N_9845,N_8992,N_8966);
xor U9846 (N_9846,N_9208,N_9269);
and U9847 (N_9847,N_9193,N_9096);
and U9848 (N_9848,N_8986,N_8818);
nor U9849 (N_9849,N_9355,N_8930);
nor U9850 (N_9850,N_9063,N_9090);
nand U9851 (N_9851,N_8791,N_9278);
or U9852 (N_9852,N_8860,N_9361);
xor U9853 (N_9853,N_8998,N_8757);
or U9854 (N_9854,N_8843,N_8996);
and U9855 (N_9855,N_9051,N_8931);
or U9856 (N_9856,N_9261,N_8950);
and U9857 (N_9857,N_8790,N_9003);
nor U9858 (N_9858,N_8883,N_8760);
nor U9859 (N_9859,N_9015,N_8973);
nand U9860 (N_9860,N_9225,N_8975);
xnor U9861 (N_9861,N_9039,N_9310);
or U9862 (N_9862,N_9003,N_8878);
or U9863 (N_9863,N_8903,N_9296);
and U9864 (N_9864,N_9295,N_9250);
nor U9865 (N_9865,N_9096,N_9181);
xor U9866 (N_9866,N_9225,N_9109);
nor U9867 (N_9867,N_9179,N_8889);
nand U9868 (N_9868,N_9238,N_9240);
nor U9869 (N_9869,N_9048,N_8983);
nand U9870 (N_9870,N_9275,N_8755);
and U9871 (N_9871,N_9150,N_9034);
nand U9872 (N_9872,N_8860,N_9345);
and U9873 (N_9873,N_9251,N_9228);
nand U9874 (N_9874,N_9063,N_8964);
and U9875 (N_9875,N_8899,N_8962);
and U9876 (N_9876,N_9020,N_9220);
nand U9877 (N_9877,N_8976,N_8797);
nand U9878 (N_9878,N_9076,N_9203);
and U9879 (N_9879,N_8765,N_9051);
or U9880 (N_9880,N_9156,N_8753);
and U9881 (N_9881,N_8789,N_9310);
or U9882 (N_9882,N_9367,N_8943);
or U9883 (N_9883,N_9173,N_8779);
nand U9884 (N_9884,N_8806,N_8890);
or U9885 (N_9885,N_9302,N_8802);
nor U9886 (N_9886,N_9297,N_9262);
and U9887 (N_9887,N_8779,N_9213);
or U9888 (N_9888,N_8955,N_8813);
nand U9889 (N_9889,N_9295,N_9294);
or U9890 (N_9890,N_8779,N_9358);
nor U9891 (N_9891,N_9357,N_9194);
nor U9892 (N_9892,N_9204,N_9106);
nor U9893 (N_9893,N_9296,N_9068);
xor U9894 (N_9894,N_9087,N_9156);
nor U9895 (N_9895,N_9153,N_8864);
xnor U9896 (N_9896,N_9223,N_9346);
nor U9897 (N_9897,N_9324,N_9223);
xor U9898 (N_9898,N_9251,N_9048);
xor U9899 (N_9899,N_9069,N_9361);
and U9900 (N_9900,N_8998,N_9056);
nand U9901 (N_9901,N_9221,N_8853);
and U9902 (N_9902,N_8896,N_9299);
nand U9903 (N_9903,N_8862,N_8996);
xor U9904 (N_9904,N_9291,N_9262);
and U9905 (N_9905,N_9121,N_9137);
and U9906 (N_9906,N_9058,N_8891);
or U9907 (N_9907,N_9116,N_9343);
nand U9908 (N_9908,N_9066,N_9277);
nor U9909 (N_9909,N_8901,N_9178);
and U9910 (N_9910,N_9269,N_8836);
and U9911 (N_9911,N_8866,N_8964);
nor U9912 (N_9912,N_8844,N_9361);
xor U9913 (N_9913,N_8991,N_9367);
xnor U9914 (N_9914,N_9025,N_9177);
nor U9915 (N_9915,N_9010,N_8896);
and U9916 (N_9916,N_8903,N_8970);
nand U9917 (N_9917,N_8861,N_9066);
or U9918 (N_9918,N_9196,N_9233);
or U9919 (N_9919,N_9045,N_9039);
or U9920 (N_9920,N_9243,N_9035);
nand U9921 (N_9921,N_9120,N_8908);
xor U9922 (N_9922,N_9128,N_8869);
and U9923 (N_9923,N_9348,N_9040);
xor U9924 (N_9924,N_9100,N_8905);
xor U9925 (N_9925,N_9070,N_8958);
xnor U9926 (N_9926,N_9060,N_8994);
xor U9927 (N_9927,N_8942,N_8994);
nor U9928 (N_9928,N_9176,N_8831);
xor U9929 (N_9929,N_8753,N_9062);
or U9930 (N_9930,N_8795,N_8985);
nor U9931 (N_9931,N_9283,N_8836);
nand U9932 (N_9932,N_9058,N_8765);
and U9933 (N_9933,N_8971,N_8863);
nor U9934 (N_9934,N_9142,N_9093);
xor U9935 (N_9935,N_9283,N_8969);
or U9936 (N_9936,N_8917,N_9141);
nor U9937 (N_9937,N_9128,N_9041);
xnor U9938 (N_9938,N_9356,N_8760);
nor U9939 (N_9939,N_9039,N_8840);
xor U9940 (N_9940,N_9243,N_9006);
and U9941 (N_9941,N_8806,N_8798);
xnor U9942 (N_9942,N_9175,N_8838);
nand U9943 (N_9943,N_8896,N_8885);
nand U9944 (N_9944,N_9323,N_8913);
and U9945 (N_9945,N_8956,N_9363);
nor U9946 (N_9946,N_9096,N_9167);
or U9947 (N_9947,N_8861,N_8771);
xnor U9948 (N_9948,N_8823,N_9174);
or U9949 (N_9949,N_8900,N_9013);
nand U9950 (N_9950,N_8982,N_8843);
nor U9951 (N_9951,N_9201,N_9223);
and U9952 (N_9952,N_9035,N_9055);
and U9953 (N_9953,N_9127,N_8929);
or U9954 (N_9954,N_8931,N_9255);
or U9955 (N_9955,N_9095,N_8754);
and U9956 (N_9956,N_9173,N_9305);
and U9957 (N_9957,N_9325,N_8816);
and U9958 (N_9958,N_8781,N_8900);
nor U9959 (N_9959,N_8774,N_9205);
xor U9960 (N_9960,N_8942,N_9149);
xnor U9961 (N_9961,N_9258,N_8863);
and U9962 (N_9962,N_8911,N_9236);
and U9963 (N_9963,N_9229,N_8881);
nand U9964 (N_9964,N_8914,N_8842);
nor U9965 (N_9965,N_8962,N_9260);
nor U9966 (N_9966,N_8896,N_9285);
nand U9967 (N_9967,N_9321,N_8944);
and U9968 (N_9968,N_9085,N_9231);
and U9969 (N_9969,N_9295,N_9111);
xnor U9970 (N_9970,N_9360,N_9355);
or U9971 (N_9971,N_9061,N_9198);
nand U9972 (N_9972,N_9103,N_9026);
nand U9973 (N_9973,N_8954,N_9273);
xnor U9974 (N_9974,N_9230,N_9300);
nand U9975 (N_9975,N_9182,N_9293);
nor U9976 (N_9976,N_9228,N_9248);
nand U9977 (N_9977,N_9342,N_8883);
nor U9978 (N_9978,N_9213,N_9186);
nor U9979 (N_9979,N_9079,N_9065);
nor U9980 (N_9980,N_8798,N_9227);
or U9981 (N_9981,N_8972,N_9031);
nand U9982 (N_9982,N_8890,N_9374);
and U9983 (N_9983,N_9092,N_9032);
or U9984 (N_9984,N_9361,N_9348);
xor U9985 (N_9985,N_9026,N_9292);
xnor U9986 (N_9986,N_9194,N_9273);
xor U9987 (N_9987,N_8893,N_9196);
nor U9988 (N_9988,N_8764,N_8797);
nand U9989 (N_9989,N_8797,N_9165);
nand U9990 (N_9990,N_8856,N_8865);
and U9991 (N_9991,N_8881,N_9115);
nor U9992 (N_9992,N_8836,N_9042);
xor U9993 (N_9993,N_8959,N_8913);
and U9994 (N_9994,N_9336,N_8970);
nor U9995 (N_9995,N_8905,N_8899);
nand U9996 (N_9996,N_8988,N_9089);
xor U9997 (N_9997,N_9043,N_9218);
nor U9998 (N_9998,N_8864,N_8842);
xor U9999 (N_9999,N_8818,N_9208);
and U10000 (N_10000,N_9781,N_9874);
nor U10001 (N_10001,N_9977,N_9898);
xnor U10002 (N_10002,N_9394,N_9725);
xor U10003 (N_10003,N_9695,N_9544);
nor U10004 (N_10004,N_9410,N_9663);
and U10005 (N_10005,N_9859,N_9403);
xor U10006 (N_10006,N_9624,N_9887);
xor U10007 (N_10007,N_9979,N_9831);
and U10008 (N_10008,N_9949,N_9908);
xnor U10009 (N_10009,N_9390,N_9751);
nand U10010 (N_10010,N_9958,N_9416);
or U10011 (N_10011,N_9535,N_9760);
nand U10012 (N_10012,N_9407,N_9658);
nor U10013 (N_10013,N_9467,N_9952);
xnor U10014 (N_10014,N_9820,N_9758);
nor U10015 (N_10015,N_9505,N_9918);
nand U10016 (N_10016,N_9912,N_9702);
nor U10017 (N_10017,N_9682,N_9630);
nand U10018 (N_10018,N_9449,N_9805);
nand U10019 (N_10019,N_9989,N_9896);
or U10020 (N_10020,N_9925,N_9627);
and U10021 (N_10021,N_9384,N_9381);
nand U10022 (N_10022,N_9901,N_9812);
nor U10023 (N_10023,N_9691,N_9744);
or U10024 (N_10024,N_9891,N_9755);
nor U10025 (N_10025,N_9763,N_9617);
nand U10026 (N_10026,N_9964,N_9404);
and U10027 (N_10027,N_9440,N_9558);
nand U10028 (N_10028,N_9612,N_9562);
xnor U10029 (N_10029,N_9942,N_9444);
xnor U10030 (N_10030,N_9645,N_9459);
xnor U10031 (N_10031,N_9936,N_9965);
nand U10032 (N_10032,N_9460,N_9547);
or U10033 (N_10033,N_9772,N_9427);
or U10034 (N_10034,N_9511,N_9639);
nand U10035 (N_10035,N_9869,N_9548);
xor U10036 (N_10036,N_9894,N_9959);
and U10037 (N_10037,N_9411,N_9516);
and U10038 (N_10038,N_9610,N_9872);
nand U10039 (N_10039,N_9541,N_9793);
nand U10040 (N_10040,N_9988,N_9454);
nand U10041 (N_10041,N_9470,N_9423);
and U10042 (N_10042,N_9521,N_9580);
xor U10043 (N_10043,N_9937,N_9383);
and U10044 (N_10044,N_9604,N_9774);
and U10045 (N_10045,N_9824,N_9780);
and U10046 (N_10046,N_9704,N_9506);
and U10047 (N_10047,N_9591,N_9689);
nand U10048 (N_10048,N_9480,N_9865);
nor U10049 (N_10049,N_9552,N_9892);
nor U10050 (N_10050,N_9884,N_9858);
and U10051 (N_10051,N_9752,N_9439);
and U10052 (N_10052,N_9487,N_9736);
and U10053 (N_10053,N_9756,N_9995);
or U10054 (N_10054,N_9693,N_9587);
and U10055 (N_10055,N_9750,N_9815);
and U10056 (N_10056,N_9779,N_9400);
nand U10057 (N_10057,N_9500,N_9644);
xnor U10058 (N_10058,N_9985,N_9453);
xor U10059 (N_10059,N_9714,N_9839);
and U10060 (N_10060,N_9983,N_9712);
nor U10061 (N_10061,N_9987,N_9569);
and U10062 (N_10062,N_9385,N_9462);
nor U10063 (N_10063,N_9741,N_9635);
nand U10064 (N_10064,N_9661,N_9943);
and U10065 (N_10065,N_9451,N_9852);
xor U10066 (N_10066,N_9534,N_9897);
xnor U10067 (N_10067,N_9655,N_9817);
xor U10068 (N_10068,N_9659,N_9559);
nor U10069 (N_10069,N_9856,N_9463);
or U10070 (N_10070,N_9398,N_9537);
or U10071 (N_10071,N_9543,N_9503);
or U10072 (N_10072,N_9709,N_9507);
and U10073 (N_10073,N_9576,N_9414);
or U10074 (N_10074,N_9531,N_9420);
xor U10075 (N_10075,N_9938,N_9551);
xnor U10076 (N_10076,N_9790,N_9546);
and U10077 (N_10077,N_9766,N_9915);
and U10078 (N_10078,N_9792,N_9926);
and U10079 (N_10079,N_9711,N_9406);
nand U10080 (N_10080,N_9388,N_9759);
and U10081 (N_10081,N_9450,N_9795);
xnor U10082 (N_10082,N_9436,N_9731);
and U10083 (N_10083,N_9803,N_9382);
xor U10084 (N_10084,N_9694,N_9701);
xnor U10085 (N_10085,N_9881,N_9556);
or U10086 (N_10086,N_9726,N_9706);
and U10087 (N_10087,N_9745,N_9491);
nand U10088 (N_10088,N_9483,N_9412);
nand U10089 (N_10089,N_9944,N_9889);
or U10090 (N_10090,N_9961,N_9703);
nand U10091 (N_10091,N_9434,N_9561);
and U10092 (N_10092,N_9818,N_9677);
or U10093 (N_10093,N_9642,N_9652);
and U10094 (N_10094,N_9939,N_9636);
or U10095 (N_10095,N_9800,N_9907);
nor U10096 (N_10096,N_9418,N_9900);
nor U10097 (N_10097,N_9433,N_9575);
nor U10098 (N_10098,N_9718,N_9466);
nand U10099 (N_10099,N_9523,N_9623);
and U10100 (N_10100,N_9667,N_9929);
nand U10101 (N_10101,N_9729,N_9681);
or U10102 (N_10102,N_9565,N_9861);
nand U10103 (N_10103,N_9847,N_9654);
nor U10104 (N_10104,N_9475,N_9796);
nand U10105 (N_10105,N_9499,N_9860);
xnor U10106 (N_10106,N_9494,N_9842);
nor U10107 (N_10107,N_9885,N_9598);
or U10108 (N_10108,N_9947,N_9857);
nor U10109 (N_10109,N_9910,N_9621);
and U10110 (N_10110,N_9783,N_9474);
nor U10111 (N_10111,N_9679,N_9422);
xor U10112 (N_10112,N_9733,N_9431);
xor U10113 (N_10113,N_9571,N_9829);
xnor U10114 (N_10114,N_9637,N_9504);
and U10115 (N_10115,N_9683,N_9764);
and U10116 (N_10116,N_9582,N_9528);
nor U10117 (N_10117,N_9438,N_9441);
xor U10118 (N_10118,N_9782,N_9395);
or U10119 (N_10119,N_9375,N_9904);
xor U10120 (N_10120,N_9909,N_9799);
nand U10121 (N_10121,N_9396,N_9666);
and U10122 (N_10122,N_9473,N_9953);
xnor U10123 (N_10123,N_9927,N_9919);
nand U10124 (N_10124,N_9950,N_9670);
xnor U10125 (N_10125,N_9513,N_9854);
xor U10126 (N_10126,N_9844,N_9622);
and U10127 (N_10127,N_9848,N_9809);
nand U10128 (N_10128,N_9498,N_9788);
xor U10129 (N_10129,N_9966,N_9605);
or U10130 (N_10130,N_9456,N_9732);
nor U10131 (N_10131,N_9674,N_9720);
nand U10132 (N_10132,N_9941,N_9485);
or U10133 (N_10133,N_9962,N_9584);
nor U10134 (N_10134,N_9607,N_9785);
or U10135 (N_10135,N_9443,N_9377);
or U10136 (N_10136,N_9405,N_9409);
or U10137 (N_10137,N_9867,N_9588);
xnor U10138 (N_10138,N_9975,N_9515);
or U10139 (N_10139,N_9748,N_9747);
nand U10140 (N_10140,N_9452,N_9963);
xnor U10141 (N_10141,N_9540,N_9845);
or U10142 (N_10142,N_9471,N_9833);
and U10143 (N_10143,N_9616,N_9802);
nor U10144 (N_10144,N_9819,N_9994);
nand U10145 (N_10145,N_9754,N_9933);
xnor U10146 (N_10146,N_9493,N_9868);
nor U10147 (N_10147,N_9469,N_9419);
or U10148 (N_10148,N_9628,N_9734);
or U10149 (N_10149,N_9830,N_9922);
xor U10150 (N_10150,N_9972,N_9986);
nand U10151 (N_10151,N_9606,N_9742);
nand U10152 (N_10152,N_9457,N_9501);
nor U10153 (N_10153,N_9735,N_9960);
and U10154 (N_10154,N_9533,N_9692);
and U10155 (N_10155,N_9631,N_9435);
nand U10156 (N_10156,N_9837,N_9461);
or U10157 (N_10157,N_9794,N_9698);
xnor U10158 (N_10158,N_9951,N_9827);
nand U10159 (N_10159,N_9722,N_9710);
nand U10160 (N_10160,N_9804,N_9832);
nor U10161 (N_10161,N_9512,N_9634);
nor U10162 (N_10162,N_9775,N_9902);
nor U10163 (N_10163,N_9386,N_9492);
xnor U10164 (N_10164,N_9554,N_9862);
nand U10165 (N_10165,N_9532,N_9539);
nor U10166 (N_10166,N_9520,N_9583);
nor U10167 (N_10167,N_9413,N_9846);
nand U10168 (N_10168,N_9821,N_9397);
and U10169 (N_10169,N_9660,N_9825);
or U10170 (N_10170,N_9905,N_9510);
xor U10171 (N_10171,N_9640,N_9651);
xnor U10172 (N_10172,N_9619,N_9990);
nand U10173 (N_10173,N_9719,N_9458);
xnor U10174 (N_10174,N_9529,N_9526);
nand U10175 (N_10175,N_9776,N_9389);
or U10176 (N_10176,N_9579,N_9527);
nand U10177 (N_10177,N_9590,N_9468);
nand U10178 (N_10178,N_9669,N_9849);
xnor U10179 (N_10179,N_9743,N_9585);
xnor U10180 (N_10180,N_9835,N_9613);
and U10181 (N_10181,N_9870,N_9968);
nor U10182 (N_10182,N_9629,N_9429);
and U10183 (N_10183,N_9808,N_9596);
and U10184 (N_10184,N_9903,N_9810);
or U10185 (N_10185,N_9864,N_9762);
nor U10186 (N_10186,N_9999,N_9424);
nor U10187 (N_10187,N_9982,N_9415);
xor U10188 (N_10188,N_9773,N_9866);
and U10189 (N_10189,N_9813,N_9542);
or U10190 (N_10190,N_9488,N_9597);
nor U10191 (N_10191,N_9997,N_9784);
nor U10192 (N_10192,N_9970,N_9768);
nand U10193 (N_10193,N_9478,N_9948);
nor U10194 (N_10194,N_9777,N_9391);
and U10195 (N_10195,N_9954,N_9538);
xnor U10196 (N_10196,N_9967,N_9574);
xnor U10197 (N_10197,N_9464,N_9568);
and U10198 (N_10198,N_9448,N_9567);
nor U10199 (N_10199,N_9921,N_9816);
xnor U10200 (N_10200,N_9611,N_9586);
xor U10201 (N_10201,N_9886,N_9671);
and U10202 (N_10202,N_9717,N_9633);
or U10203 (N_10203,N_9978,N_9871);
nor U10204 (N_10204,N_9757,N_9417);
nand U10205 (N_10205,N_9662,N_9888);
and U10206 (N_10206,N_9992,N_9680);
or U10207 (N_10207,N_9955,N_9738);
or U10208 (N_10208,N_9822,N_9545);
nor U10209 (N_10209,N_9497,N_9855);
or U10210 (N_10210,N_9724,N_9570);
nand U10211 (N_10211,N_9566,N_9653);
and U10212 (N_10212,N_9932,N_9996);
xor U10213 (N_10213,N_9798,N_9826);
nor U10214 (N_10214,N_9530,N_9749);
or U10215 (N_10215,N_9899,N_9442);
nor U10216 (N_10216,N_9601,N_9518);
nand U10217 (N_10217,N_9836,N_9879);
xor U10218 (N_10218,N_9626,N_9646);
nor U10219 (N_10219,N_9550,N_9700);
or U10220 (N_10220,N_9770,N_9421);
and U10221 (N_10221,N_9761,N_9913);
and U10222 (N_10222,N_9519,N_9916);
nor U10223 (N_10223,N_9957,N_9882);
and U10224 (N_10224,N_9946,N_9924);
nand U10225 (N_10225,N_9876,N_9873);
xor U10226 (N_10226,N_9625,N_9524);
and U10227 (N_10227,N_9509,N_9850);
or U10228 (N_10228,N_9578,N_9676);
nor U10229 (N_10229,N_9618,N_9664);
or U10230 (N_10230,N_9895,N_9739);
xnor U10231 (N_10231,N_9589,N_9976);
and U10232 (N_10232,N_9806,N_9684);
or U10233 (N_10233,N_9984,N_9811);
xnor U10234 (N_10234,N_9807,N_9956);
and U10235 (N_10235,N_9974,N_9593);
xor U10236 (N_10236,N_9599,N_9797);
nand U10237 (N_10237,N_9697,N_9594);
xor U10238 (N_10238,N_9823,N_9981);
xnor U10239 (N_10239,N_9609,N_9934);
xnor U10240 (N_10240,N_9437,N_9393);
and U10241 (N_10241,N_9392,N_9786);
nand U10242 (N_10242,N_9746,N_9880);
or U10243 (N_10243,N_9484,N_9557);
xor U10244 (N_10244,N_9878,N_9841);
nor U10245 (N_10245,N_9787,N_9705);
xnor U10246 (N_10246,N_9665,N_9928);
nand U10247 (N_10247,N_9998,N_9685);
nor U10248 (N_10248,N_9477,N_9971);
xnor U10249 (N_10249,N_9638,N_9863);
and U10250 (N_10250,N_9708,N_9696);
or U10251 (N_10251,N_9911,N_9602);
nor U10252 (N_10252,N_9707,N_9426);
nand U10253 (N_10253,N_9716,N_9379);
and U10254 (N_10254,N_9486,N_9490);
nor U10255 (N_10255,N_9522,N_9840);
and U10256 (N_10256,N_9430,N_9673);
nand U10257 (N_10257,N_9647,N_9791);
nor U10258 (N_10258,N_9893,N_9428);
and U10259 (N_10259,N_9920,N_9801);
nand U10260 (N_10260,N_9380,N_9940);
nand U10261 (N_10261,N_9581,N_9969);
nand U10262 (N_10262,N_9945,N_9387);
and U10263 (N_10263,N_9432,N_9657);
or U10264 (N_10264,N_9402,N_9650);
or U10265 (N_10265,N_9401,N_9476);
nor U10266 (N_10266,N_9495,N_9648);
or U10267 (N_10267,N_9479,N_9721);
nor U10268 (N_10268,N_9672,N_9489);
nand U10269 (N_10269,N_9875,N_9536);
nor U10270 (N_10270,N_9834,N_9771);
and U10271 (N_10271,N_9603,N_9686);
nor U10272 (N_10272,N_9668,N_9767);
or U10273 (N_10273,N_9641,N_9917);
and U10274 (N_10274,N_9560,N_9525);
nor U10275 (N_10275,N_9715,N_9572);
nor U10276 (N_10276,N_9973,N_9789);
nand U10277 (N_10277,N_9455,N_9980);
and U10278 (N_10278,N_9713,N_9906);
and U10279 (N_10279,N_9502,N_9555);
nand U10280 (N_10280,N_9482,N_9378);
nand U10281 (N_10281,N_9496,N_9408);
nand U10282 (N_10282,N_9553,N_9914);
xnor U10283 (N_10283,N_9399,N_9993);
xnor U10284 (N_10284,N_9425,N_9481);
or U10285 (N_10285,N_9577,N_9472);
nand U10286 (N_10286,N_9890,N_9643);
nand U10287 (N_10287,N_9446,N_9930);
and U10288 (N_10288,N_9730,N_9935);
xor U10289 (N_10289,N_9549,N_9675);
nor U10290 (N_10290,N_9563,N_9931);
xor U10291 (N_10291,N_9465,N_9728);
xor U10292 (N_10292,N_9608,N_9649);
and U10293 (N_10293,N_9564,N_9615);
nor U10294 (N_10294,N_9517,N_9877);
nand U10295 (N_10295,N_9600,N_9620);
and U10296 (N_10296,N_9851,N_9778);
nor U10297 (N_10297,N_9508,N_9592);
or U10298 (N_10298,N_9883,N_9690);
or U10299 (N_10299,N_9828,N_9699);
xnor U10300 (N_10300,N_9656,N_9753);
nor U10301 (N_10301,N_9687,N_9853);
nor U10302 (N_10302,N_9814,N_9514);
and U10303 (N_10303,N_9688,N_9447);
or U10304 (N_10304,N_9737,N_9769);
xor U10305 (N_10305,N_9740,N_9632);
xor U10306 (N_10306,N_9445,N_9727);
nand U10307 (N_10307,N_9765,N_9595);
nand U10308 (N_10308,N_9376,N_9723);
xnor U10309 (N_10309,N_9838,N_9614);
nand U10310 (N_10310,N_9991,N_9843);
xor U10311 (N_10311,N_9573,N_9923);
and U10312 (N_10312,N_9678,N_9453);
or U10313 (N_10313,N_9868,N_9684);
xnor U10314 (N_10314,N_9851,N_9931);
nand U10315 (N_10315,N_9457,N_9515);
nand U10316 (N_10316,N_9378,N_9540);
and U10317 (N_10317,N_9540,N_9674);
xnor U10318 (N_10318,N_9927,N_9502);
or U10319 (N_10319,N_9975,N_9731);
nor U10320 (N_10320,N_9738,N_9852);
nand U10321 (N_10321,N_9395,N_9528);
nor U10322 (N_10322,N_9851,N_9448);
and U10323 (N_10323,N_9941,N_9884);
and U10324 (N_10324,N_9750,N_9411);
nor U10325 (N_10325,N_9443,N_9384);
and U10326 (N_10326,N_9780,N_9627);
xnor U10327 (N_10327,N_9458,N_9727);
or U10328 (N_10328,N_9950,N_9396);
and U10329 (N_10329,N_9800,N_9962);
or U10330 (N_10330,N_9865,N_9422);
nor U10331 (N_10331,N_9536,N_9491);
xnor U10332 (N_10332,N_9792,N_9995);
and U10333 (N_10333,N_9386,N_9862);
nand U10334 (N_10334,N_9601,N_9925);
or U10335 (N_10335,N_9891,N_9798);
xnor U10336 (N_10336,N_9642,N_9934);
xor U10337 (N_10337,N_9864,N_9586);
and U10338 (N_10338,N_9928,N_9841);
or U10339 (N_10339,N_9681,N_9888);
nor U10340 (N_10340,N_9877,N_9459);
nand U10341 (N_10341,N_9699,N_9960);
nand U10342 (N_10342,N_9656,N_9566);
or U10343 (N_10343,N_9732,N_9687);
nand U10344 (N_10344,N_9515,N_9700);
xnor U10345 (N_10345,N_9736,N_9630);
and U10346 (N_10346,N_9962,N_9382);
xor U10347 (N_10347,N_9580,N_9577);
nand U10348 (N_10348,N_9915,N_9985);
nor U10349 (N_10349,N_9902,N_9498);
and U10350 (N_10350,N_9825,N_9819);
nand U10351 (N_10351,N_9968,N_9985);
nand U10352 (N_10352,N_9893,N_9613);
and U10353 (N_10353,N_9777,N_9560);
or U10354 (N_10354,N_9882,N_9799);
or U10355 (N_10355,N_9828,N_9854);
nand U10356 (N_10356,N_9862,N_9756);
nand U10357 (N_10357,N_9623,N_9701);
nand U10358 (N_10358,N_9784,N_9760);
nand U10359 (N_10359,N_9586,N_9408);
nor U10360 (N_10360,N_9596,N_9782);
or U10361 (N_10361,N_9666,N_9383);
xnor U10362 (N_10362,N_9776,N_9543);
nand U10363 (N_10363,N_9975,N_9634);
or U10364 (N_10364,N_9608,N_9585);
xnor U10365 (N_10365,N_9630,N_9508);
or U10366 (N_10366,N_9459,N_9780);
and U10367 (N_10367,N_9478,N_9782);
and U10368 (N_10368,N_9417,N_9760);
nand U10369 (N_10369,N_9567,N_9692);
nand U10370 (N_10370,N_9588,N_9875);
xnor U10371 (N_10371,N_9770,N_9531);
or U10372 (N_10372,N_9709,N_9915);
and U10373 (N_10373,N_9482,N_9768);
nand U10374 (N_10374,N_9939,N_9606);
or U10375 (N_10375,N_9527,N_9439);
nand U10376 (N_10376,N_9536,N_9813);
and U10377 (N_10377,N_9597,N_9476);
and U10378 (N_10378,N_9965,N_9844);
and U10379 (N_10379,N_9939,N_9963);
nand U10380 (N_10380,N_9980,N_9526);
and U10381 (N_10381,N_9812,N_9999);
xnor U10382 (N_10382,N_9606,N_9502);
xnor U10383 (N_10383,N_9823,N_9772);
nand U10384 (N_10384,N_9476,N_9770);
or U10385 (N_10385,N_9460,N_9467);
nand U10386 (N_10386,N_9387,N_9471);
xor U10387 (N_10387,N_9659,N_9649);
nand U10388 (N_10388,N_9396,N_9554);
or U10389 (N_10389,N_9733,N_9833);
xnor U10390 (N_10390,N_9453,N_9751);
and U10391 (N_10391,N_9793,N_9479);
xor U10392 (N_10392,N_9711,N_9474);
nor U10393 (N_10393,N_9407,N_9529);
or U10394 (N_10394,N_9453,N_9980);
xor U10395 (N_10395,N_9655,N_9875);
xor U10396 (N_10396,N_9427,N_9786);
xnor U10397 (N_10397,N_9828,N_9791);
xor U10398 (N_10398,N_9866,N_9573);
nand U10399 (N_10399,N_9694,N_9752);
or U10400 (N_10400,N_9862,N_9906);
xnor U10401 (N_10401,N_9715,N_9491);
and U10402 (N_10402,N_9481,N_9855);
and U10403 (N_10403,N_9889,N_9447);
or U10404 (N_10404,N_9728,N_9959);
xor U10405 (N_10405,N_9923,N_9819);
or U10406 (N_10406,N_9459,N_9430);
xnor U10407 (N_10407,N_9401,N_9759);
and U10408 (N_10408,N_9859,N_9703);
xor U10409 (N_10409,N_9501,N_9740);
and U10410 (N_10410,N_9450,N_9541);
xor U10411 (N_10411,N_9467,N_9816);
and U10412 (N_10412,N_9825,N_9850);
xor U10413 (N_10413,N_9556,N_9570);
or U10414 (N_10414,N_9712,N_9925);
and U10415 (N_10415,N_9544,N_9404);
xor U10416 (N_10416,N_9390,N_9890);
or U10417 (N_10417,N_9651,N_9687);
nand U10418 (N_10418,N_9579,N_9952);
xnor U10419 (N_10419,N_9446,N_9912);
and U10420 (N_10420,N_9574,N_9633);
and U10421 (N_10421,N_9894,N_9484);
nand U10422 (N_10422,N_9848,N_9741);
nor U10423 (N_10423,N_9621,N_9613);
nor U10424 (N_10424,N_9448,N_9467);
or U10425 (N_10425,N_9883,N_9773);
or U10426 (N_10426,N_9740,N_9863);
or U10427 (N_10427,N_9687,N_9618);
and U10428 (N_10428,N_9606,N_9801);
and U10429 (N_10429,N_9942,N_9732);
xnor U10430 (N_10430,N_9594,N_9977);
nand U10431 (N_10431,N_9604,N_9663);
nor U10432 (N_10432,N_9751,N_9907);
nand U10433 (N_10433,N_9527,N_9653);
and U10434 (N_10434,N_9412,N_9384);
and U10435 (N_10435,N_9710,N_9596);
xor U10436 (N_10436,N_9946,N_9509);
and U10437 (N_10437,N_9474,N_9861);
nor U10438 (N_10438,N_9953,N_9532);
and U10439 (N_10439,N_9843,N_9591);
nor U10440 (N_10440,N_9773,N_9899);
xnor U10441 (N_10441,N_9819,N_9406);
xnor U10442 (N_10442,N_9605,N_9910);
and U10443 (N_10443,N_9469,N_9665);
or U10444 (N_10444,N_9478,N_9530);
xnor U10445 (N_10445,N_9723,N_9447);
xnor U10446 (N_10446,N_9947,N_9378);
or U10447 (N_10447,N_9964,N_9901);
or U10448 (N_10448,N_9727,N_9922);
or U10449 (N_10449,N_9527,N_9675);
or U10450 (N_10450,N_9399,N_9795);
or U10451 (N_10451,N_9768,N_9542);
nor U10452 (N_10452,N_9413,N_9679);
or U10453 (N_10453,N_9860,N_9383);
nor U10454 (N_10454,N_9412,N_9602);
nor U10455 (N_10455,N_9878,N_9761);
xnor U10456 (N_10456,N_9546,N_9395);
nand U10457 (N_10457,N_9996,N_9891);
xnor U10458 (N_10458,N_9746,N_9918);
xnor U10459 (N_10459,N_9467,N_9723);
xnor U10460 (N_10460,N_9526,N_9582);
and U10461 (N_10461,N_9951,N_9761);
or U10462 (N_10462,N_9384,N_9657);
nand U10463 (N_10463,N_9944,N_9476);
nor U10464 (N_10464,N_9666,N_9522);
and U10465 (N_10465,N_9881,N_9521);
nor U10466 (N_10466,N_9447,N_9458);
or U10467 (N_10467,N_9744,N_9433);
xnor U10468 (N_10468,N_9836,N_9388);
or U10469 (N_10469,N_9528,N_9617);
nand U10470 (N_10470,N_9962,N_9818);
nand U10471 (N_10471,N_9926,N_9598);
or U10472 (N_10472,N_9904,N_9422);
nor U10473 (N_10473,N_9422,N_9971);
and U10474 (N_10474,N_9820,N_9565);
xnor U10475 (N_10475,N_9774,N_9928);
nor U10476 (N_10476,N_9808,N_9959);
or U10477 (N_10477,N_9545,N_9699);
nand U10478 (N_10478,N_9392,N_9708);
nor U10479 (N_10479,N_9550,N_9950);
or U10480 (N_10480,N_9433,N_9893);
or U10481 (N_10481,N_9698,N_9968);
xor U10482 (N_10482,N_9698,N_9694);
nand U10483 (N_10483,N_9593,N_9434);
nor U10484 (N_10484,N_9845,N_9687);
nor U10485 (N_10485,N_9568,N_9826);
or U10486 (N_10486,N_9683,N_9563);
and U10487 (N_10487,N_9487,N_9918);
and U10488 (N_10488,N_9950,N_9930);
xnor U10489 (N_10489,N_9571,N_9979);
and U10490 (N_10490,N_9816,N_9486);
nand U10491 (N_10491,N_9463,N_9929);
nor U10492 (N_10492,N_9600,N_9675);
or U10493 (N_10493,N_9660,N_9553);
and U10494 (N_10494,N_9719,N_9700);
nand U10495 (N_10495,N_9777,N_9909);
xor U10496 (N_10496,N_9407,N_9749);
xor U10497 (N_10497,N_9538,N_9802);
and U10498 (N_10498,N_9410,N_9744);
nand U10499 (N_10499,N_9979,N_9924);
nor U10500 (N_10500,N_9871,N_9601);
nor U10501 (N_10501,N_9937,N_9432);
xor U10502 (N_10502,N_9987,N_9889);
or U10503 (N_10503,N_9599,N_9758);
nand U10504 (N_10504,N_9748,N_9985);
and U10505 (N_10505,N_9765,N_9486);
and U10506 (N_10506,N_9987,N_9836);
or U10507 (N_10507,N_9965,N_9930);
or U10508 (N_10508,N_9804,N_9525);
or U10509 (N_10509,N_9966,N_9540);
and U10510 (N_10510,N_9686,N_9571);
nand U10511 (N_10511,N_9727,N_9764);
nand U10512 (N_10512,N_9474,N_9538);
nand U10513 (N_10513,N_9470,N_9677);
xor U10514 (N_10514,N_9690,N_9918);
xor U10515 (N_10515,N_9405,N_9934);
nor U10516 (N_10516,N_9460,N_9801);
and U10517 (N_10517,N_9989,N_9955);
nand U10518 (N_10518,N_9871,N_9955);
xnor U10519 (N_10519,N_9690,N_9873);
nand U10520 (N_10520,N_9685,N_9452);
nor U10521 (N_10521,N_9626,N_9729);
nand U10522 (N_10522,N_9655,N_9465);
xor U10523 (N_10523,N_9474,N_9389);
or U10524 (N_10524,N_9898,N_9410);
xor U10525 (N_10525,N_9710,N_9614);
nand U10526 (N_10526,N_9643,N_9579);
nand U10527 (N_10527,N_9959,N_9706);
xnor U10528 (N_10528,N_9947,N_9636);
xor U10529 (N_10529,N_9741,N_9856);
nor U10530 (N_10530,N_9802,N_9857);
and U10531 (N_10531,N_9872,N_9755);
or U10532 (N_10532,N_9915,N_9635);
and U10533 (N_10533,N_9496,N_9460);
nand U10534 (N_10534,N_9688,N_9411);
or U10535 (N_10535,N_9535,N_9531);
or U10536 (N_10536,N_9491,N_9946);
xor U10537 (N_10537,N_9971,N_9808);
or U10538 (N_10538,N_9695,N_9733);
or U10539 (N_10539,N_9393,N_9436);
or U10540 (N_10540,N_9498,N_9681);
nor U10541 (N_10541,N_9764,N_9595);
nand U10542 (N_10542,N_9629,N_9649);
and U10543 (N_10543,N_9868,N_9598);
xor U10544 (N_10544,N_9673,N_9799);
xor U10545 (N_10545,N_9951,N_9993);
or U10546 (N_10546,N_9655,N_9400);
xor U10547 (N_10547,N_9809,N_9441);
and U10548 (N_10548,N_9500,N_9977);
xnor U10549 (N_10549,N_9705,N_9957);
and U10550 (N_10550,N_9846,N_9420);
nand U10551 (N_10551,N_9711,N_9573);
xnor U10552 (N_10552,N_9620,N_9803);
and U10553 (N_10553,N_9493,N_9744);
xnor U10554 (N_10554,N_9649,N_9617);
or U10555 (N_10555,N_9492,N_9867);
xor U10556 (N_10556,N_9389,N_9479);
nand U10557 (N_10557,N_9526,N_9757);
nor U10558 (N_10558,N_9405,N_9617);
nand U10559 (N_10559,N_9801,N_9601);
and U10560 (N_10560,N_9393,N_9620);
nand U10561 (N_10561,N_9381,N_9830);
nor U10562 (N_10562,N_9619,N_9822);
or U10563 (N_10563,N_9705,N_9833);
or U10564 (N_10564,N_9747,N_9507);
nor U10565 (N_10565,N_9982,N_9523);
and U10566 (N_10566,N_9491,N_9621);
or U10567 (N_10567,N_9999,N_9612);
nor U10568 (N_10568,N_9930,N_9466);
nor U10569 (N_10569,N_9442,N_9498);
or U10570 (N_10570,N_9632,N_9813);
nor U10571 (N_10571,N_9561,N_9815);
and U10572 (N_10572,N_9462,N_9410);
or U10573 (N_10573,N_9958,N_9624);
xnor U10574 (N_10574,N_9691,N_9380);
or U10575 (N_10575,N_9679,N_9629);
or U10576 (N_10576,N_9508,N_9947);
nand U10577 (N_10577,N_9627,N_9577);
or U10578 (N_10578,N_9968,N_9902);
xnor U10579 (N_10579,N_9652,N_9684);
and U10580 (N_10580,N_9833,N_9781);
and U10581 (N_10581,N_9846,N_9582);
and U10582 (N_10582,N_9814,N_9625);
nand U10583 (N_10583,N_9716,N_9638);
nor U10584 (N_10584,N_9817,N_9380);
or U10585 (N_10585,N_9698,N_9906);
and U10586 (N_10586,N_9399,N_9821);
xnor U10587 (N_10587,N_9639,N_9666);
xnor U10588 (N_10588,N_9376,N_9765);
nand U10589 (N_10589,N_9789,N_9936);
nor U10590 (N_10590,N_9894,N_9835);
and U10591 (N_10591,N_9702,N_9541);
xor U10592 (N_10592,N_9784,N_9605);
xnor U10593 (N_10593,N_9622,N_9953);
xnor U10594 (N_10594,N_9756,N_9506);
xnor U10595 (N_10595,N_9928,N_9767);
or U10596 (N_10596,N_9436,N_9596);
or U10597 (N_10597,N_9503,N_9554);
nor U10598 (N_10598,N_9527,N_9896);
and U10599 (N_10599,N_9707,N_9816);
and U10600 (N_10600,N_9904,N_9459);
nor U10601 (N_10601,N_9918,N_9757);
xnor U10602 (N_10602,N_9849,N_9591);
xnor U10603 (N_10603,N_9651,N_9711);
xor U10604 (N_10604,N_9447,N_9460);
xnor U10605 (N_10605,N_9634,N_9712);
nand U10606 (N_10606,N_9687,N_9431);
xnor U10607 (N_10607,N_9922,N_9612);
and U10608 (N_10608,N_9825,N_9403);
or U10609 (N_10609,N_9496,N_9391);
xnor U10610 (N_10610,N_9474,N_9717);
nor U10611 (N_10611,N_9850,N_9845);
nor U10612 (N_10612,N_9595,N_9458);
nand U10613 (N_10613,N_9619,N_9722);
nor U10614 (N_10614,N_9912,N_9709);
xnor U10615 (N_10615,N_9715,N_9868);
and U10616 (N_10616,N_9911,N_9833);
nand U10617 (N_10617,N_9634,N_9570);
nand U10618 (N_10618,N_9861,N_9763);
nand U10619 (N_10619,N_9762,N_9958);
nand U10620 (N_10620,N_9824,N_9986);
xor U10621 (N_10621,N_9738,N_9985);
or U10622 (N_10622,N_9599,N_9458);
or U10623 (N_10623,N_9852,N_9483);
or U10624 (N_10624,N_9934,N_9821);
nand U10625 (N_10625,N_10129,N_10033);
and U10626 (N_10626,N_10378,N_10456);
and U10627 (N_10627,N_10581,N_10293);
xor U10628 (N_10628,N_10253,N_10319);
xor U10629 (N_10629,N_10026,N_10406);
nor U10630 (N_10630,N_10149,N_10452);
xor U10631 (N_10631,N_10298,N_10186);
xor U10632 (N_10632,N_10175,N_10619);
xor U10633 (N_10633,N_10357,N_10037);
xnor U10634 (N_10634,N_10524,N_10522);
xnor U10635 (N_10635,N_10296,N_10562);
nand U10636 (N_10636,N_10084,N_10220);
or U10637 (N_10637,N_10019,N_10170);
xnor U10638 (N_10638,N_10481,N_10178);
and U10639 (N_10639,N_10153,N_10394);
nor U10640 (N_10640,N_10287,N_10521);
xor U10641 (N_10641,N_10317,N_10001);
nor U10642 (N_10642,N_10448,N_10372);
xor U10643 (N_10643,N_10229,N_10135);
or U10644 (N_10644,N_10161,N_10071);
or U10645 (N_10645,N_10155,N_10416);
xnor U10646 (N_10646,N_10530,N_10586);
xor U10647 (N_10647,N_10484,N_10017);
and U10648 (N_10648,N_10100,N_10344);
nor U10649 (N_10649,N_10348,N_10483);
nor U10650 (N_10650,N_10476,N_10563);
and U10651 (N_10651,N_10313,N_10486);
or U10652 (N_10652,N_10151,N_10127);
nor U10653 (N_10653,N_10393,N_10021);
xor U10654 (N_10654,N_10396,N_10463);
xor U10655 (N_10655,N_10095,N_10116);
xnor U10656 (N_10656,N_10526,N_10173);
or U10657 (N_10657,N_10035,N_10402);
nor U10658 (N_10658,N_10320,N_10600);
nand U10659 (N_10659,N_10371,N_10027);
and U10660 (N_10660,N_10460,N_10340);
and U10661 (N_10661,N_10141,N_10308);
or U10662 (N_10662,N_10236,N_10596);
nor U10663 (N_10663,N_10609,N_10454);
nor U10664 (N_10664,N_10086,N_10509);
or U10665 (N_10665,N_10098,N_10252);
nand U10666 (N_10666,N_10089,N_10176);
nand U10667 (N_10667,N_10496,N_10039);
nor U10668 (N_10668,N_10488,N_10603);
and U10669 (N_10669,N_10497,N_10615);
xnor U10670 (N_10670,N_10223,N_10144);
and U10671 (N_10671,N_10540,N_10601);
nand U10672 (N_10672,N_10025,N_10589);
nand U10673 (N_10673,N_10459,N_10218);
or U10674 (N_10674,N_10267,N_10554);
nor U10675 (N_10675,N_10381,N_10042);
or U10676 (N_10676,N_10111,N_10584);
and U10677 (N_10677,N_10262,N_10499);
nand U10678 (N_10678,N_10230,N_10567);
xnor U10679 (N_10679,N_10281,N_10269);
or U10680 (N_10680,N_10582,N_10055);
xor U10681 (N_10681,N_10527,N_10342);
and U10682 (N_10682,N_10446,N_10438);
and U10683 (N_10683,N_10002,N_10558);
nor U10684 (N_10684,N_10171,N_10383);
and U10685 (N_10685,N_10442,N_10215);
nand U10686 (N_10686,N_10045,N_10096);
nand U10687 (N_10687,N_10079,N_10246);
and U10688 (N_10688,N_10489,N_10386);
xor U10689 (N_10689,N_10485,N_10400);
xnor U10690 (N_10690,N_10380,N_10066);
or U10691 (N_10691,N_10228,N_10598);
xor U10692 (N_10692,N_10290,N_10472);
nor U10693 (N_10693,N_10180,N_10477);
nand U10694 (N_10694,N_10196,N_10292);
or U10695 (N_10695,N_10610,N_10323);
or U10696 (N_10696,N_10411,N_10005);
nor U10697 (N_10697,N_10106,N_10117);
nand U10698 (N_10698,N_10085,N_10605);
and U10699 (N_10699,N_10191,N_10058);
nor U10700 (N_10700,N_10611,N_10076);
and U10701 (N_10701,N_10133,N_10044);
and U10702 (N_10702,N_10368,N_10195);
nor U10703 (N_10703,N_10333,N_10213);
and U10704 (N_10704,N_10205,N_10245);
and U10705 (N_10705,N_10103,N_10599);
nor U10706 (N_10706,N_10053,N_10054);
nand U10707 (N_10707,N_10546,N_10192);
nor U10708 (N_10708,N_10221,N_10336);
nand U10709 (N_10709,N_10209,N_10064);
nor U10710 (N_10710,N_10107,N_10061);
nor U10711 (N_10711,N_10250,N_10181);
or U10712 (N_10712,N_10238,N_10617);
and U10713 (N_10713,N_10295,N_10108);
xor U10714 (N_10714,N_10036,N_10128);
nand U10715 (N_10715,N_10275,N_10571);
xnor U10716 (N_10716,N_10138,N_10011);
or U10717 (N_10717,N_10373,N_10360);
xnor U10718 (N_10718,N_10356,N_10326);
nand U10719 (N_10719,N_10556,N_10322);
and U10720 (N_10720,N_10088,N_10003);
nand U10721 (N_10721,N_10427,N_10550);
xnor U10722 (N_10722,N_10305,N_10234);
nand U10723 (N_10723,N_10034,N_10444);
xor U10724 (N_10724,N_10056,N_10227);
and U10725 (N_10725,N_10078,N_10219);
or U10726 (N_10726,N_10433,N_10552);
or U10727 (N_10727,N_10212,N_10043);
xnor U10728 (N_10728,N_10490,N_10614);
nand U10729 (N_10729,N_10453,N_10255);
nor U10730 (N_10730,N_10118,N_10410);
nand U10731 (N_10731,N_10000,N_10504);
nor U10732 (N_10732,N_10572,N_10137);
or U10733 (N_10733,N_10211,N_10346);
xor U10734 (N_10734,N_10533,N_10478);
nand U10735 (N_10735,N_10082,N_10125);
and U10736 (N_10736,N_10193,N_10154);
xor U10737 (N_10737,N_10102,N_10101);
or U10738 (N_10738,N_10624,N_10506);
nor U10739 (N_10739,N_10266,N_10502);
nor U10740 (N_10740,N_10491,N_10471);
xnor U10741 (N_10741,N_10508,N_10534);
xor U10742 (N_10742,N_10315,N_10022);
nand U10743 (N_10743,N_10143,N_10131);
nand U10744 (N_10744,N_10505,N_10525);
nor U10745 (N_10745,N_10539,N_10353);
nor U10746 (N_10746,N_10382,N_10465);
and U10747 (N_10747,N_10294,N_10300);
or U10748 (N_10748,N_10408,N_10029);
or U10749 (N_10749,N_10473,N_10240);
nand U10750 (N_10750,N_10561,N_10543);
nand U10751 (N_10751,N_10265,N_10520);
nand U10752 (N_10752,N_10097,N_10146);
and U10753 (N_10753,N_10041,N_10541);
and U10754 (N_10754,N_10060,N_10006);
nand U10755 (N_10755,N_10349,N_10403);
nor U10756 (N_10756,N_10457,N_10425);
or U10757 (N_10757,N_10415,N_10009);
or U10758 (N_10758,N_10426,N_10545);
nor U10759 (N_10759,N_10578,N_10474);
xnor U10760 (N_10760,N_10350,N_10487);
or U10761 (N_10761,N_10225,N_10007);
and U10762 (N_10762,N_10094,N_10222);
xnor U10763 (N_10763,N_10283,N_10551);
and U10764 (N_10764,N_10560,N_10437);
and U10765 (N_10765,N_10395,N_10413);
and U10766 (N_10766,N_10420,N_10365);
nand U10767 (N_10767,N_10592,N_10169);
and U10768 (N_10768,N_10419,N_10038);
nand U10769 (N_10769,N_10286,N_10436);
or U10770 (N_10770,N_10503,N_10165);
and U10771 (N_10771,N_10580,N_10316);
nand U10772 (N_10772,N_10384,N_10608);
or U10773 (N_10773,N_10004,N_10148);
or U10774 (N_10774,N_10203,N_10341);
or U10775 (N_10775,N_10087,N_10324);
nor U10776 (N_10776,N_10105,N_10210);
or U10777 (N_10777,N_10013,N_10397);
or U10778 (N_10778,N_10335,N_10217);
and U10779 (N_10779,N_10355,N_10516);
nand U10780 (N_10780,N_10115,N_10070);
nand U10781 (N_10781,N_10432,N_10142);
nor U10782 (N_10782,N_10440,N_10303);
nand U10783 (N_10783,N_10622,N_10276);
nand U10784 (N_10784,N_10214,N_10553);
nand U10785 (N_10785,N_10259,N_10405);
nand U10786 (N_10786,N_10260,N_10233);
and U10787 (N_10787,N_10069,N_10291);
xor U10788 (N_10788,N_10535,N_10075);
and U10789 (N_10789,N_10168,N_10174);
and U10790 (N_10790,N_10401,N_10242);
xor U10791 (N_10791,N_10249,N_10239);
and U10792 (N_10792,N_10469,N_10574);
nand U10793 (N_10793,N_10126,N_10409);
or U10794 (N_10794,N_10159,N_10197);
nor U10795 (N_10795,N_10555,N_10590);
nand U10796 (N_10796,N_10351,N_10237);
and U10797 (N_10797,N_10597,N_10422);
or U10798 (N_10798,N_10428,N_10354);
nand U10799 (N_10799,N_10424,N_10362);
xor U10800 (N_10800,N_10157,N_10270);
xor U10801 (N_10801,N_10059,N_10049);
xnor U10802 (N_10802,N_10235,N_10389);
nand U10803 (N_10803,N_10492,N_10309);
and U10804 (N_10804,N_10528,N_10542);
nor U10805 (N_10805,N_10156,N_10172);
nor U10806 (N_10806,N_10304,N_10529);
and U10807 (N_10807,N_10392,N_10136);
nand U10808 (N_10808,N_10390,N_10374);
xor U10809 (N_10809,N_10498,N_10455);
and U10810 (N_10810,N_10421,N_10470);
or U10811 (N_10811,N_10514,N_10570);
nand U10812 (N_10812,N_10251,N_10429);
xnor U10813 (N_10813,N_10065,N_10271);
nor U10814 (N_10814,N_10032,N_10339);
xor U10815 (N_10815,N_10583,N_10407);
xor U10816 (N_10816,N_10081,N_10519);
nor U10817 (N_10817,N_10050,N_10536);
xor U10818 (N_10818,N_10189,N_10202);
xnor U10819 (N_10819,N_10361,N_10312);
nor U10820 (N_10820,N_10591,N_10207);
nor U10821 (N_10821,N_10417,N_10152);
or U10822 (N_10822,N_10538,N_10122);
nor U10823 (N_10823,N_10014,N_10020);
xnor U10824 (N_10824,N_10160,N_10162);
and U10825 (N_10825,N_10307,N_10187);
nand U10826 (N_10826,N_10375,N_10537);
and U10827 (N_10827,N_10548,N_10338);
nand U10828 (N_10828,N_10464,N_10123);
nor U10829 (N_10829,N_10364,N_10493);
xor U10830 (N_10830,N_10461,N_10208);
or U10831 (N_10831,N_10347,N_10145);
nor U10832 (N_10832,N_10345,N_10593);
nor U10833 (N_10833,N_10216,N_10099);
or U10834 (N_10834,N_10274,N_10564);
nor U10835 (N_10835,N_10080,N_10363);
and U10836 (N_10836,N_10048,N_10370);
or U10837 (N_10837,N_10412,N_10575);
or U10838 (N_10838,N_10258,N_10376);
nor U10839 (N_10839,N_10450,N_10458);
or U10840 (N_10840,N_10447,N_10434);
or U10841 (N_10841,N_10404,N_10623);
xor U10842 (N_10842,N_10494,N_10254);
nand U10843 (N_10843,N_10482,N_10147);
xnor U10844 (N_10844,N_10532,N_10012);
nand U10845 (N_10845,N_10515,N_10579);
xnor U10846 (N_10846,N_10329,N_10243);
or U10847 (N_10847,N_10139,N_10198);
nand U10848 (N_10848,N_10423,N_10414);
or U10849 (N_10849,N_10366,N_10057);
and U10850 (N_10850,N_10587,N_10388);
nand U10851 (N_10851,N_10311,N_10051);
and U10852 (N_10852,N_10273,N_10507);
xnor U10853 (N_10853,N_10285,N_10475);
nor U10854 (N_10854,N_10387,N_10566);
nor U10855 (N_10855,N_10248,N_10369);
xor U10856 (N_10856,N_10167,N_10093);
xor U10857 (N_10857,N_10468,N_10263);
and U10858 (N_10858,N_10268,N_10439);
xnor U10859 (N_10859,N_10569,N_10431);
nand U10860 (N_10860,N_10279,N_10606);
or U10861 (N_10861,N_10164,N_10449);
or U10862 (N_10862,N_10337,N_10030);
xnor U10863 (N_10863,N_10299,N_10612);
nor U10864 (N_10864,N_10008,N_10090);
xor U10865 (N_10865,N_10278,N_10501);
and U10866 (N_10866,N_10015,N_10616);
nor U10867 (N_10867,N_10018,N_10512);
or U10868 (N_10868,N_10301,N_10379);
or U10869 (N_10869,N_10231,N_10523);
nand U10870 (N_10870,N_10023,N_10352);
or U10871 (N_10871,N_10334,N_10188);
nand U10872 (N_10872,N_10330,N_10264);
and U10873 (N_10873,N_10310,N_10120);
nor U10874 (N_10874,N_10067,N_10028);
nor U10875 (N_10875,N_10130,N_10547);
and U10876 (N_10876,N_10083,N_10518);
and U10877 (N_10877,N_10114,N_10140);
nand U10878 (N_10878,N_10201,N_10288);
xor U10879 (N_10879,N_10511,N_10435);
and U10880 (N_10880,N_10358,N_10092);
nor U10881 (N_10881,N_10559,N_10289);
nor U10882 (N_10882,N_10185,N_10620);
nor U10883 (N_10883,N_10166,N_10072);
xnor U10884 (N_10884,N_10328,N_10479);
xor U10885 (N_10885,N_10595,N_10112);
nand U10886 (N_10886,N_10531,N_10576);
or U10887 (N_10887,N_10302,N_10613);
xnor U10888 (N_10888,N_10343,N_10241);
and U10889 (N_10889,N_10047,N_10391);
nand U10890 (N_10890,N_10282,N_10052);
or U10891 (N_10891,N_10510,N_10573);
or U10892 (N_10892,N_10318,N_10297);
xnor U10893 (N_10893,N_10332,N_10577);
xnor U10894 (N_10894,N_10104,N_10158);
or U10895 (N_10895,N_10091,N_10077);
xor U10896 (N_10896,N_10256,N_10445);
nand U10897 (N_10897,N_10602,N_10257);
xnor U10898 (N_10898,N_10321,N_10132);
and U10899 (N_10899,N_10177,N_10031);
nand U10900 (N_10900,N_10443,N_10441);
and U10901 (N_10901,N_10124,N_10277);
nand U10902 (N_10902,N_10010,N_10607);
xor U10903 (N_10903,N_10232,N_10544);
xnor U10904 (N_10904,N_10466,N_10063);
xnor U10905 (N_10905,N_10306,N_10451);
or U10906 (N_10906,N_10430,N_10113);
or U10907 (N_10907,N_10024,N_10109);
or U10908 (N_10908,N_10224,N_10183);
xnor U10909 (N_10909,N_10557,N_10480);
nand U10910 (N_10910,N_10467,N_10068);
nand U10911 (N_10911,N_10062,N_10226);
xor U10912 (N_10912,N_10621,N_10073);
nand U10913 (N_10913,N_10331,N_10399);
or U10914 (N_10914,N_10204,N_10604);
nor U10915 (N_10915,N_10549,N_10134);
nand U10916 (N_10916,N_10199,N_10182);
and U10917 (N_10917,N_10040,N_10074);
nand U10918 (N_10918,N_10618,N_10119);
xor U10919 (N_10919,N_10517,N_10568);
and U10920 (N_10920,N_10163,N_10325);
or U10921 (N_10921,N_10261,N_10588);
xor U10922 (N_10922,N_10327,N_10206);
nand U10923 (N_10923,N_10513,N_10495);
and U10924 (N_10924,N_10462,N_10046);
and U10925 (N_10925,N_10194,N_10280);
and U10926 (N_10926,N_10272,N_10418);
or U10927 (N_10927,N_10377,N_10247);
nand U10928 (N_10928,N_10016,N_10184);
xor U10929 (N_10929,N_10314,N_10150);
and U10930 (N_10930,N_10585,N_10359);
xor U10931 (N_10931,N_10565,N_10594);
or U10932 (N_10932,N_10367,N_10385);
xor U10933 (N_10933,N_10190,N_10500);
xor U10934 (N_10934,N_10244,N_10110);
xor U10935 (N_10935,N_10179,N_10284);
nor U10936 (N_10936,N_10121,N_10398);
nor U10937 (N_10937,N_10200,N_10134);
xor U10938 (N_10938,N_10233,N_10022);
xor U10939 (N_10939,N_10288,N_10027);
xor U10940 (N_10940,N_10179,N_10595);
nand U10941 (N_10941,N_10210,N_10265);
xnor U10942 (N_10942,N_10327,N_10205);
and U10943 (N_10943,N_10415,N_10031);
nand U10944 (N_10944,N_10621,N_10615);
or U10945 (N_10945,N_10623,N_10102);
or U10946 (N_10946,N_10510,N_10412);
or U10947 (N_10947,N_10231,N_10053);
and U10948 (N_10948,N_10280,N_10325);
xor U10949 (N_10949,N_10168,N_10208);
nand U10950 (N_10950,N_10002,N_10358);
nor U10951 (N_10951,N_10210,N_10445);
xor U10952 (N_10952,N_10208,N_10419);
nand U10953 (N_10953,N_10579,N_10282);
nor U10954 (N_10954,N_10507,N_10153);
and U10955 (N_10955,N_10282,N_10292);
and U10956 (N_10956,N_10164,N_10095);
nand U10957 (N_10957,N_10498,N_10596);
nand U10958 (N_10958,N_10428,N_10119);
nand U10959 (N_10959,N_10577,N_10074);
or U10960 (N_10960,N_10387,N_10206);
or U10961 (N_10961,N_10122,N_10356);
xor U10962 (N_10962,N_10464,N_10231);
nor U10963 (N_10963,N_10398,N_10268);
or U10964 (N_10964,N_10468,N_10451);
xor U10965 (N_10965,N_10188,N_10214);
and U10966 (N_10966,N_10088,N_10438);
xnor U10967 (N_10967,N_10068,N_10097);
nand U10968 (N_10968,N_10060,N_10258);
nand U10969 (N_10969,N_10215,N_10152);
and U10970 (N_10970,N_10422,N_10444);
or U10971 (N_10971,N_10301,N_10428);
nand U10972 (N_10972,N_10409,N_10515);
nand U10973 (N_10973,N_10436,N_10115);
nor U10974 (N_10974,N_10032,N_10517);
nor U10975 (N_10975,N_10607,N_10203);
nand U10976 (N_10976,N_10599,N_10569);
nor U10977 (N_10977,N_10108,N_10168);
and U10978 (N_10978,N_10624,N_10108);
and U10979 (N_10979,N_10524,N_10515);
nor U10980 (N_10980,N_10593,N_10004);
and U10981 (N_10981,N_10282,N_10387);
and U10982 (N_10982,N_10482,N_10384);
xor U10983 (N_10983,N_10109,N_10167);
nor U10984 (N_10984,N_10485,N_10577);
or U10985 (N_10985,N_10019,N_10232);
or U10986 (N_10986,N_10052,N_10554);
nor U10987 (N_10987,N_10095,N_10243);
or U10988 (N_10988,N_10564,N_10246);
or U10989 (N_10989,N_10083,N_10134);
xor U10990 (N_10990,N_10169,N_10281);
and U10991 (N_10991,N_10602,N_10045);
nor U10992 (N_10992,N_10194,N_10152);
xnor U10993 (N_10993,N_10273,N_10379);
nand U10994 (N_10994,N_10455,N_10077);
nor U10995 (N_10995,N_10595,N_10447);
xnor U10996 (N_10996,N_10012,N_10400);
xnor U10997 (N_10997,N_10469,N_10480);
nand U10998 (N_10998,N_10394,N_10543);
and U10999 (N_10999,N_10433,N_10478);
and U11000 (N_11000,N_10463,N_10156);
nor U11001 (N_11001,N_10597,N_10285);
or U11002 (N_11002,N_10568,N_10223);
xor U11003 (N_11003,N_10365,N_10205);
or U11004 (N_11004,N_10514,N_10100);
xor U11005 (N_11005,N_10535,N_10609);
nor U11006 (N_11006,N_10452,N_10366);
xor U11007 (N_11007,N_10434,N_10451);
or U11008 (N_11008,N_10342,N_10291);
and U11009 (N_11009,N_10566,N_10445);
nor U11010 (N_11010,N_10441,N_10125);
nand U11011 (N_11011,N_10196,N_10074);
nand U11012 (N_11012,N_10000,N_10226);
nand U11013 (N_11013,N_10194,N_10133);
and U11014 (N_11014,N_10239,N_10039);
nor U11015 (N_11015,N_10334,N_10597);
xor U11016 (N_11016,N_10624,N_10608);
nand U11017 (N_11017,N_10552,N_10042);
nand U11018 (N_11018,N_10056,N_10259);
nand U11019 (N_11019,N_10065,N_10500);
nor U11020 (N_11020,N_10491,N_10282);
nor U11021 (N_11021,N_10084,N_10521);
or U11022 (N_11022,N_10392,N_10480);
xnor U11023 (N_11023,N_10086,N_10014);
and U11024 (N_11024,N_10281,N_10143);
and U11025 (N_11025,N_10193,N_10265);
nand U11026 (N_11026,N_10187,N_10236);
and U11027 (N_11027,N_10389,N_10027);
nor U11028 (N_11028,N_10081,N_10335);
or U11029 (N_11029,N_10357,N_10389);
or U11030 (N_11030,N_10177,N_10005);
nor U11031 (N_11031,N_10594,N_10524);
nand U11032 (N_11032,N_10270,N_10318);
nand U11033 (N_11033,N_10057,N_10196);
and U11034 (N_11034,N_10064,N_10046);
nor U11035 (N_11035,N_10419,N_10179);
nor U11036 (N_11036,N_10171,N_10172);
and U11037 (N_11037,N_10091,N_10384);
xor U11038 (N_11038,N_10226,N_10283);
and U11039 (N_11039,N_10407,N_10209);
and U11040 (N_11040,N_10410,N_10144);
xor U11041 (N_11041,N_10220,N_10355);
nor U11042 (N_11042,N_10011,N_10565);
nor U11043 (N_11043,N_10191,N_10135);
nor U11044 (N_11044,N_10161,N_10486);
nand U11045 (N_11045,N_10237,N_10532);
or U11046 (N_11046,N_10267,N_10591);
and U11047 (N_11047,N_10034,N_10176);
nand U11048 (N_11048,N_10558,N_10018);
and U11049 (N_11049,N_10537,N_10135);
nand U11050 (N_11050,N_10543,N_10446);
nor U11051 (N_11051,N_10110,N_10188);
nor U11052 (N_11052,N_10177,N_10089);
xor U11053 (N_11053,N_10573,N_10576);
nor U11054 (N_11054,N_10577,N_10039);
nor U11055 (N_11055,N_10256,N_10077);
and U11056 (N_11056,N_10380,N_10477);
nand U11057 (N_11057,N_10606,N_10136);
and U11058 (N_11058,N_10447,N_10405);
and U11059 (N_11059,N_10100,N_10536);
nand U11060 (N_11060,N_10270,N_10286);
nor U11061 (N_11061,N_10364,N_10309);
and U11062 (N_11062,N_10621,N_10081);
nand U11063 (N_11063,N_10565,N_10408);
or U11064 (N_11064,N_10501,N_10131);
xor U11065 (N_11065,N_10407,N_10011);
nand U11066 (N_11066,N_10274,N_10187);
nand U11067 (N_11067,N_10560,N_10039);
nand U11068 (N_11068,N_10013,N_10435);
nor U11069 (N_11069,N_10215,N_10523);
and U11070 (N_11070,N_10268,N_10115);
and U11071 (N_11071,N_10156,N_10528);
and U11072 (N_11072,N_10151,N_10139);
or U11073 (N_11073,N_10243,N_10088);
nor U11074 (N_11074,N_10613,N_10075);
nor U11075 (N_11075,N_10315,N_10498);
nand U11076 (N_11076,N_10443,N_10494);
or U11077 (N_11077,N_10546,N_10621);
xnor U11078 (N_11078,N_10205,N_10520);
nor U11079 (N_11079,N_10450,N_10084);
nor U11080 (N_11080,N_10437,N_10031);
nand U11081 (N_11081,N_10275,N_10021);
nand U11082 (N_11082,N_10355,N_10285);
or U11083 (N_11083,N_10467,N_10285);
xor U11084 (N_11084,N_10414,N_10506);
or U11085 (N_11085,N_10026,N_10294);
or U11086 (N_11086,N_10025,N_10540);
nor U11087 (N_11087,N_10384,N_10310);
nand U11088 (N_11088,N_10105,N_10624);
xor U11089 (N_11089,N_10329,N_10366);
nand U11090 (N_11090,N_10112,N_10373);
xor U11091 (N_11091,N_10492,N_10541);
and U11092 (N_11092,N_10446,N_10518);
nor U11093 (N_11093,N_10427,N_10502);
or U11094 (N_11094,N_10490,N_10447);
and U11095 (N_11095,N_10534,N_10530);
and U11096 (N_11096,N_10291,N_10124);
or U11097 (N_11097,N_10574,N_10458);
nor U11098 (N_11098,N_10065,N_10188);
nor U11099 (N_11099,N_10028,N_10090);
and U11100 (N_11100,N_10192,N_10161);
nand U11101 (N_11101,N_10307,N_10081);
and U11102 (N_11102,N_10066,N_10183);
and U11103 (N_11103,N_10104,N_10045);
nand U11104 (N_11104,N_10419,N_10171);
xor U11105 (N_11105,N_10091,N_10106);
xor U11106 (N_11106,N_10265,N_10573);
xnor U11107 (N_11107,N_10024,N_10364);
xor U11108 (N_11108,N_10385,N_10504);
or U11109 (N_11109,N_10229,N_10268);
nor U11110 (N_11110,N_10182,N_10559);
nor U11111 (N_11111,N_10138,N_10534);
nor U11112 (N_11112,N_10328,N_10519);
and U11113 (N_11113,N_10200,N_10250);
nand U11114 (N_11114,N_10538,N_10581);
and U11115 (N_11115,N_10186,N_10437);
or U11116 (N_11116,N_10131,N_10479);
or U11117 (N_11117,N_10496,N_10452);
or U11118 (N_11118,N_10258,N_10287);
or U11119 (N_11119,N_10511,N_10524);
and U11120 (N_11120,N_10406,N_10400);
and U11121 (N_11121,N_10406,N_10568);
xnor U11122 (N_11122,N_10262,N_10596);
nand U11123 (N_11123,N_10259,N_10174);
nor U11124 (N_11124,N_10123,N_10579);
or U11125 (N_11125,N_10159,N_10461);
nand U11126 (N_11126,N_10417,N_10573);
and U11127 (N_11127,N_10583,N_10269);
or U11128 (N_11128,N_10234,N_10451);
and U11129 (N_11129,N_10475,N_10038);
or U11130 (N_11130,N_10021,N_10078);
nor U11131 (N_11131,N_10341,N_10265);
nor U11132 (N_11132,N_10548,N_10174);
nor U11133 (N_11133,N_10431,N_10014);
nor U11134 (N_11134,N_10535,N_10073);
nor U11135 (N_11135,N_10380,N_10053);
xor U11136 (N_11136,N_10035,N_10102);
and U11137 (N_11137,N_10311,N_10009);
nor U11138 (N_11138,N_10336,N_10353);
or U11139 (N_11139,N_10225,N_10430);
nor U11140 (N_11140,N_10473,N_10263);
nand U11141 (N_11141,N_10206,N_10557);
nor U11142 (N_11142,N_10090,N_10510);
or U11143 (N_11143,N_10291,N_10174);
and U11144 (N_11144,N_10014,N_10622);
xnor U11145 (N_11145,N_10124,N_10352);
xnor U11146 (N_11146,N_10000,N_10558);
and U11147 (N_11147,N_10624,N_10190);
nand U11148 (N_11148,N_10324,N_10437);
or U11149 (N_11149,N_10326,N_10008);
nand U11150 (N_11150,N_10318,N_10145);
nand U11151 (N_11151,N_10259,N_10210);
and U11152 (N_11152,N_10127,N_10508);
or U11153 (N_11153,N_10145,N_10293);
nor U11154 (N_11154,N_10593,N_10179);
xor U11155 (N_11155,N_10567,N_10004);
xnor U11156 (N_11156,N_10441,N_10452);
or U11157 (N_11157,N_10172,N_10511);
nor U11158 (N_11158,N_10252,N_10232);
xor U11159 (N_11159,N_10153,N_10296);
and U11160 (N_11160,N_10407,N_10346);
nand U11161 (N_11161,N_10318,N_10083);
xor U11162 (N_11162,N_10234,N_10379);
xor U11163 (N_11163,N_10083,N_10220);
nor U11164 (N_11164,N_10512,N_10040);
or U11165 (N_11165,N_10589,N_10040);
and U11166 (N_11166,N_10258,N_10137);
or U11167 (N_11167,N_10216,N_10298);
xor U11168 (N_11168,N_10532,N_10399);
or U11169 (N_11169,N_10281,N_10004);
xnor U11170 (N_11170,N_10089,N_10155);
and U11171 (N_11171,N_10407,N_10531);
xor U11172 (N_11172,N_10207,N_10123);
or U11173 (N_11173,N_10024,N_10239);
or U11174 (N_11174,N_10427,N_10210);
and U11175 (N_11175,N_10097,N_10508);
and U11176 (N_11176,N_10223,N_10460);
nor U11177 (N_11177,N_10302,N_10179);
nand U11178 (N_11178,N_10525,N_10297);
xnor U11179 (N_11179,N_10109,N_10014);
nand U11180 (N_11180,N_10073,N_10056);
and U11181 (N_11181,N_10205,N_10302);
and U11182 (N_11182,N_10583,N_10053);
nor U11183 (N_11183,N_10196,N_10003);
nand U11184 (N_11184,N_10593,N_10497);
nand U11185 (N_11185,N_10585,N_10590);
or U11186 (N_11186,N_10063,N_10088);
or U11187 (N_11187,N_10079,N_10439);
or U11188 (N_11188,N_10296,N_10602);
or U11189 (N_11189,N_10259,N_10180);
xnor U11190 (N_11190,N_10562,N_10535);
nor U11191 (N_11191,N_10178,N_10010);
nor U11192 (N_11192,N_10161,N_10360);
and U11193 (N_11193,N_10337,N_10589);
xor U11194 (N_11194,N_10069,N_10355);
nand U11195 (N_11195,N_10434,N_10074);
and U11196 (N_11196,N_10518,N_10130);
nand U11197 (N_11197,N_10510,N_10624);
and U11198 (N_11198,N_10009,N_10095);
or U11199 (N_11199,N_10239,N_10555);
xor U11200 (N_11200,N_10254,N_10605);
nand U11201 (N_11201,N_10125,N_10130);
and U11202 (N_11202,N_10376,N_10593);
nor U11203 (N_11203,N_10390,N_10218);
or U11204 (N_11204,N_10481,N_10168);
xnor U11205 (N_11205,N_10101,N_10466);
and U11206 (N_11206,N_10248,N_10299);
xnor U11207 (N_11207,N_10566,N_10412);
xnor U11208 (N_11208,N_10154,N_10061);
and U11209 (N_11209,N_10404,N_10104);
xor U11210 (N_11210,N_10274,N_10201);
nor U11211 (N_11211,N_10366,N_10498);
and U11212 (N_11212,N_10247,N_10138);
and U11213 (N_11213,N_10053,N_10619);
nor U11214 (N_11214,N_10031,N_10401);
xnor U11215 (N_11215,N_10087,N_10292);
xnor U11216 (N_11216,N_10337,N_10102);
and U11217 (N_11217,N_10373,N_10377);
xor U11218 (N_11218,N_10137,N_10078);
nand U11219 (N_11219,N_10519,N_10583);
and U11220 (N_11220,N_10374,N_10036);
nand U11221 (N_11221,N_10573,N_10059);
or U11222 (N_11222,N_10287,N_10336);
nor U11223 (N_11223,N_10476,N_10095);
and U11224 (N_11224,N_10433,N_10029);
or U11225 (N_11225,N_10049,N_10561);
xor U11226 (N_11226,N_10122,N_10310);
xnor U11227 (N_11227,N_10151,N_10087);
and U11228 (N_11228,N_10243,N_10429);
nand U11229 (N_11229,N_10152,N_10134);
nand U11230 (N_11230,N_10146,N_10114);
nor U11231 (N_11231,N_10235,N_10339);
nor U11232 (N_11232,N_10046,N_10364);
nor U11233 (N_11233,N_10338,N_10525);
and U11234 (N_11234,N_10370,N_10126);
xor U11235 (N_11235,N_10536,N_10371);
xnor U11236 (N_11236,N_10110,N_10438);
and U11237 (N_11237,N_10492,N_10445);
nor U11238 (N_11238,N_10524,N_10508);
and U11239 (N_11239,N_10142,N_10153);
or U11240 (N_11240,N_10481,N_10286);
xnor U11241 (N_11241,N_10208,N_10145);
nand U11242 (N_11242,N_10200,N_10207);
and U11243 (N_11243,N_10368,N_10219);
or U11244 (N_11244,N_10032,N_10037);
or U11245 (N_11245,N_10328,N_10212);
or U11246 (N_11246,N_10452,N_10612);
xor U11247 (N_11247,N_10026,N_10327);
xor U11248 (N_11248,N_10134,N_10196);
nor U11249 (N_11249,N_10374,N_10211);
xnor U11250 (N_11250,N_10766,N_10896);
or U11251 (N_11251,N_11096,N_11115);
nor U11252 (N_11252,N_10952,N_10734);
and U11253 (N_11253,N_11105,N_10872);
or U11254 (N_11254,N_10651,N_11237);
nand U11255 (N_11255,N_10824,N_11076);
nand U11256 (N_11256,N_11019,N_10640);
and U11257 (N_11257,N_10750,N_10695);
and U11258 (N_11258,N_11007,N_11229);
nand U11259 (N_11259,N_11062,N_11089);
and U11260 (N_11260,N_10764,N_10806);
or U11261 (N_11261,N_10926,N_11038);
nand U11262 (N_11262,N_11234,N_10707);
xor U11263 (N_11263,N_10888,N_10979);
nor U11264 (N_11264,N_10785,N_10756);
nand U11265 (N_11265,N_10646,N_10835);
and U11266 (N_11266,N_10794,N_10757);
nand U11267 (N_11267,N_10712,N_11092);
nand U11268 (N_11268,N_10967,N_10660);
or U11269 (N_11269,N_11233,N_10983);
xor U11270 (N_11270,N_11131,N_11039);
and U11271 (N_11271,N_10997,N_11168);
and U11272 (N_11272,N_11130,N_10724);
xor U11273 (N_11273,N_10694,N_11203);
and U11274 (N_11274,N_10716,N_11159);
xnor U11275 (N_11275,N_10783,N_11023);
xor U11276 (N_11276,N_11249,N_11008);
xor U11277 (N_11277,N_11172,N_11107);
nor U11278 (N_11278,N_10637,N_10927);
xor U11279 (N_11279,N_10991,N_11033);
nand U11280 (N_11280,N_10720,N_10976);
or U11281 (N_11281,N_10752,N_11171);
or U11282 (N_11282,N_11197,N_11167);
nor U11283 (N_11283,N_10698,N_10971);
nor U11284 (N_11284,N_10930,N_10986);
nor U11285 (N_11285,N_11065,N_10892);
or U11286 (N_11286,N_10700,N_10643);
and U11287 (N_11287,N_10679,N_11148);
nand U11288 (N_11288,N_11202,N_10995);
nor U11289 (N_11289,N_10788,N_10918);
nor U11290 (N_11290,N_11052,N_11022);
xnor U11291 (N_11291,N_10726,N_10733);
nor U11292 (N_11292,N_11177,N_11060);
or U11293 (N_11293,N_11059,N_11143);
and U11294 (N_11294,N_10838,N_11078);
nand U11295 (N_11295,N_10663,N_10741);
nor U11296 (N_11296,N_10877,N_11009);
and U11297 (N_11297,N_11054,N_10960);
xor U11298 (N_11298,N_10682,N_10987);
nor U11299 (N_11299,N_11098,N_11160);
and U11300 (N_11300,N_10933,N_11137);
and U11301 (N_11301,N_10938,N_11138);
and U11302 (N_11302,N_11163,N_10642);
nor U11303 (N_11303,N_10721,N_10902);
and U11304 (N_11304,N_10943,N_10895);
nand U11305 (N_11305,N_10920,N_11086);
or U11306 (N_11306,N_11087,N_11174);
nand U11307 (N_11307,N_11027,N_10941);
and U11308 (N_11308,N_10740,N_10836);
nand U11309 (N_11309,N_11020,N_10846);
nand U11310 (N_11310,N_10645,N_11241);
or U11311 (N_11311,N_11194,N_11067);
nand U11312 (N_11312,N_11013,N_11072);
xor U11313 (N_11313,N_10865,N_10944);
xnor U11314 (N_11314,N_11166,N_10728);
nor U11315 (N_11315,N_11176,N_11201);
xor U11316 (N_11316,N_10860,N_11103);
or U11317 (N_11317,N_11217,N_10963);
nand U11318 (N_11318,N_10826,N_10666);
nor U11319 (N_11319,N_11097,N_11232);
nand U11320 (N_11320,N_10980,N_11040);
xor U11321 (N_11321,N_10650,N_11212);
nand U11322 (N_11322,N_10706,N_10774);
and U11323 (N_11323,N_10777,N_11073);
nor U11324 (N_11324,N_10825,N_10885);
and U11325 (N_11325,N_11046,N_10684);
xnor U11326 (N_11326,N_10714,N_10989);
or U11327 (N_11327,N_11108,N_10935);
nand U11328 (N_11328,N_10688,N_11026);
xor U11329 (N_11329,N_11122,N_11156);
and U11330 (N_11330,N_11061,N_11180);
xnor U11331 (N_11331,N_11014,N_10665);
nand U11332 (N_11332,N_11200,N_10680);
and U11333 (N_11333,N_10880,N_11124);
xnor U11334 (N_11334,N_10898,N_11185);
nand U11335 (N_11335,N_10855,N_10932);
or U11336 (N_11336,N_10951,N_10917);
nand U11337 (N_11337,N_10737,N_11225);
nor U11338 (N_11338,N_10809,N_11074);
or U11339 (N_11339,N_11015,N_10644);
nor U11340 (N_11340,N_10886,N_10953);
nor U11341 (N_11341,N_10656,N_10715);
nor U11342 (N_11342,N_10866,N_11002);
nand U11343 (N_11343,N_11178,N_10819);
nor U11344 (N_11344,N_10845,N_11001);
xnor U11345 (N_11345,N_10831,N_11081);
xnor U11346 (N_11346,N_11181,N_10730);
or U11347 (N_11347,N_11042,N_10914);
nand U11348 (N_11348,N_10638,N_10887);
xor U11349 (N_11349,N_11104,N_11184);
or U11350 (N_11350,N_10924,N_11169);
and U11351 (N_11351,N_11085,N_11221);
nor U11352 (N_11352,N_11247,N_10863);
nor U11353 (N_11353,N_10678,N_10994);
nor U11354 (N_11354,N_10973,N_10767);
and U11355 (N_11355,N_11133,N_10889);
nand U11356 (N_11356,N_11165,N_10697);
nor U11357 (N_11357,N_10760,N_11035);
xor U11358 (N_11358,N_11183,N_10870);
xnor U11359 (N_11359,N_11179,N_10790);
xor U11360 (N_11360,N_11211,N_11208);
xor U11361 (N_11361,N_10744,N_10956);
or U11362 (N_11362,N_10659,N_10894);
nand U11363 (N_11363,N_11210,N_11209);
or U11364 (N_11364,N_11069,N_11017);
nor U11365 (N_11365,N_10999,N_10811);
nor U11366 (N_11366,N_10843,N_10667);
or U11367 (N_11367,N_10639,N_10862);
nand U11368 (N_11368,N_11031,N_10751);
and U11369 (N_11369,N_10881,N_11173);
or U11370 (N_11370,N_10735,N_10796);
xor U11371 (N_11371,N_10670,N_11094);
xor U11372 (N_11372,N_11029,N_11125);
or U11373 (N_11373,N_10805,N_11034);
nand U11374 (N_11374,N_10725,N_10627);
xnor U11375 (N_11375,N_10940,N_11110);
xnor U11376 (N_11376,N_10975,N_11196);
xor U11377 (N_11377,N_11158,N_11117);
or U11378 (N_11378,N_10792,N_10647);
or U11379 (N_11379,N_10769,N_10625);
xor U11380 (N_11380,N_11030,N_10736);
nand U11381 (N_11381,N_10801,N_10799);
or U11382 (N_11382,N_10984,N_10633);
or U11383 (N_11383,N_10705,N_10683);
xor U11384 (N_11384,N_11175,N_10701);
or U11385 (N_11385,N_11090,N_11000);
or U11386 (N_11386,N_11161,N_10906);
or U11387 (N_11387,N_10878,N_10823);
and U11388 (N_11388,N_10711,N_11239);
nand U11389 (N_11389,N_10985,N_11248);
or U11390 (N_11390,N_10753,N_10628);
nand U11391 (N_11391,N_10791,N_11219);
nand U11392 (N_11392,N_10754,N_11136);
nor U11393 (N_11393,N_10850,N_11222);
or U11394 (N_11394,N_10818,N_10832);
or U11395 (N_11395,N_10709,N_10739);
or U11396 (N_11396,N_10847,N_10890);
nor U11397 (N_11397,N_10871,N_11224);
xnor U11398 (N_11398,N_11189,N_10844);
xor U11399 (N_11399,N_11246,N_10936);
or U11400 (N_11400,N_11135,N_10852);
nor U11401 (N_11401,N_10648,N_11231);
xor U11402 (N_11402,N_10814,N_10743);
nand U11403 (N_11403,N_11213,N_11106);
nor U11404 (N_11404,N_11113,N_11240);
nor U11405 (N_11405,N_11063,N_11091);
nor U11406 (N_11406,N_11064,N_10817);
or U11407 (N_11407,N_10770,N_10830);
nand U11408 (N_11408,N_10797,N_11121);
nor U11409 (N_11409,N_10954,N_11041);
or U11410 (N_11410,N_10626,N_11226);
nand U11411 (N_11411,N_10849,N_11101);
nor U11412 (N_11412,N_10910,N_10854);
xnor U11413 (N_11413,N_11170,N_10840);
and U11414 (N_11414,N_10658,N_11223);
xor U11415 (N_11415,N_10717,N_11036);
xor U11416 (N_11416,N_11099,N_11032);
or U11417 (N_11417,N_10718,N_10929);
xnor U11418 (N_11418,N_10758,N_11126);
and U11419 (N_11419,N_10691,N_11195);
xnor U11420 (N_11420,N_10900,N_10765);
nor U11421 (N_11421,N_10681,N_10807);
nor U11422 (N_11422,N_10674,N_11244);
and U11423 (N_11423,N_10867,N_11164);
or U11424 (N_11424,N_11018,N_11070);
and U11425 (N_11425,N_11193,N_10781);
nor U11426 (N_11426,N_11095,N_10653);
and U11427 (N_11427,N_10861,N_10812);
xor U11428 (N_11428,N_11152,N_10687);
and U11429 (N_11429,N_10925,N_11218);
and U11430 (N_11430,N_10719,N_11047);
nand U11431 (N_11431,N_10988,N_11192);
xnor U11432 (N_11432,N_10978,N_11116);
nand U11433 (N_11433,N_11088,N_10897);
nand U11434 (N_11434,N_11214,N_10820);
or U11435 (N_11435,N_10652,N_10772);
nor U11436 (N_11436,N_10636,N_11003);
nor U11437 (N_11437,N_10876,N_10841);
xnor U11438 (N_11438,N_10798,N_10710);
nor U11439 (N_11439,N_11128,N_10629);
nand U11440 (N_11440,N_10907,N_10789);
nor U11441 (N_11441,N_11146,N_11140);
nor U11442 (N_11442,N_11083,N_11245);
or U11443 (N_11443,N_10673,N_11227);
or U11444 (N_11444,N_11057,N_10827);
nand U11445 (N_11445,N_10996,N_10928);
nor U11446 (N_11446,N_11187,N_10795);
and U11447 (N_11447,N_11111,N_10748);
and U11448 (N_11448,N_10749,N_10822);
or U11449 (N_11449,N_10990,N_10787);
xor U11450 (N_11450,N_10873,N_10837);
nor U11451 (N_11451,N_11228,N_10632);
xnor U11452 (N_11452,N_10833,N_10962);
and U11453 (N_11453,N_11051,N_10704);
xnor U11454 (N_11454,N_10780,N_10968);
or U11455 (N_11455,N_10759,N_10955);
xor U11456 (N_11456,N_10634,N_10828);
or U11457 (N_11457,N_10675,N_10803);
xnor U11458 (N_11458,N_10786,N_10768);
nand U11459 (N_11459,N_10703,N_10690);
or U11460 (N_11460,N_11045,N_10713);
nand U11461 (N_11461,N_10696,N_10972);
or U11462 (N_11462,N_10908,N_10883);
or U11463 (N_11463,N_10661,N_10631);
nand U11464 (N_11464,N_11006,N_11075);
nor U11465 (N_11465,N_10722,N_10856);
nand U11466 (N_11466,N_10993,N_11093);
xor U11467 (N_11467,N_10692,N_11132);
xnor U11468 (N_11468,N_10905,N_10912);
or U11469 (N_11469,N_11186,N_10964);
and U11470 (N_11470,N_11120,N_11118);
nor U11471 (N_11471,N_11190,N_11114);
xor U11472 (N_11472,N_10657,N_11109);
nor U11473 (N_11473,N_10738,N_11084);
nand U11474 (N_11474,N_10949,N_10958);
nor U11475 (N_11475,N_11157,N_10884);
or U11476 (N_11476,N_10868,N_10702);
and U11477 (N_11477,N_10946,N_10649);
nor U11478 (N_11478,N_10974,N_11139);
nor U11479 (N_11479,N_10911,N_11100);
nor U11480 (N_11480,N_11058,N_11056);
nor U11481 (N_11481,N_10755,N_10810);
nor U11482 (N_11482,N_11149,N_10934);
xor U11483 (N_11483,N_10899,N_10879);
xor U11484 (N_11484,N_10793,N_11150);
xnor U11485 (N_11485,N_10784,N_10723);
nor U11486 (N_11486,N_10668,N_11021);
xor U11487 (N_11487,N_11010,N_10654);
nand U11488 (N_11488,N_11080,N_11153);
or U11489 (N_11489,N_11242,N_10800);
xnor U11490 (N_11490,N_10808,N_10708);
or U11491 (N_11491,N_11071,N_11123);
xnor U11492 (N_11492,N_10761,N_10662);
nor U11493 (N_11493,N_10630,N_11220);
nand U11494 (N_11494,N_10950,N_10815);
xnor U11495 (N_11495,N_11005,N_10913);
and U11496 (N_11496,N_11024,N_11141);
or U11497 (N_11497,N_11236,N_10763);
and U11498 (N_11498,N_11216,N_10677);
xor U11499 (N_11499,N_10776,N_10998);
and U11500 (N_11500,N_10893,N_11199);
xnor U11501 (N_11501,N_11144,N_10961);
or U11502 (N_11502,N_10802,N_10909);
nand U11503 (N_11503,N_11053,N_11049);
or U11504 (N_11504,N_11188,N_11151);
xor U11505 (N_11505,N_11154,N_10982);
xnor U11506 (N_11506,N_10945,N_10672);
nor U11507 (N_11507,N_11238,N_11147);
nand U11508 (N_11508,N_10947,N_11145);
nor U11509 (N_11509,N_10731,N_10859);
xnor U11510 (N_11510,N_11028,N_10966);
nand U11511 (N_11511,N_10641,N_10957);
nand U11512 (N_11512,N_11044,N_11205);
or U11513 (N_11513,N_11068,N_10775);
nor U11514 (N_11514,N_11079,N_11043);
nand U11515 (N_11515,N_10858,N_11082);
xor U11516 (N_11516,N_11182,N_11142);
xnor U11517 (N_11517,N_10729,N_10903);
nand U11518 (N_11518,N_10851,N_10782);
nand U11519 (N_11519,N_11011,N_10857);
nand U11520 (N_11520,N_11207,N_10919);
and U11521 (N_11521,N_11191,N_10816);
nor U11522 (N_11522,N_10977,N_11155);
xor U11523 (N_11523,N_10992,N_10671);
nor U11524 (N_11524,N_11004,N_10746);
nor U11525 (N_11525,N_10939,N_11127);
and U11526 (N_11526,N_10693,N_11129);
nor U11527 (N_11527,N_10875,N_10931);
and U11528 (N_11528,N_11243,N_10773);
and U11529 (N_11529,N_11025,N_11077);
or U11530 (N_11530,N_10969,N_10742);
and U11531 (N_11531,N_10689,N_10874);
xnor U11532 (N_11532,N_10834,N_10655);
nand U11533 (N_11533,N_10981,N_10959);
xor U11534 (N_11534,N_11048,N_10771);
and U11535 (N_11535,N_10747,N_10821);
and U11536 (N_11536,N_10699,N_10664);
or U11537 (N_11537,N_10732,N_10778);
xnor U11538 (N_11538,N_10915,N_11012);
xor U11539 (N_11539,N_11119,N_10942);
and U11540 (N_11540,N_10635,N_11235);
or U11541 (N_11541,N_10922,N_10762);
nand U11542 (N_11542,N_11204,N_11230);
nor U11543 (N_11543,N_10948,N_10685);
nor U11544 (N_11544,N_10937,N_10842);
or U11545 (N_11545,N_10965,N_11162);
xnor U11546 (N_11546,N_11112,N_10882);
nor U11547 (N_11547,N_11066,N_11134);
or U11548 (N_11548,N_11206,N_10864);
or U11549 (N_11549,N_10970,N_10869);
xnor U11550 (N_11550,N_10848,N_10839);
and U11551 (N_11551,N_10923,N_10891);
and U11552 (N_11552,N_10686,N_10829);
or U11553 (N_11553,N_11055,N_11050);
and U11554 (N_11554,N_10904,N_10901);
nand U11555 (N_11555,N_11037,N_11198);
and U11556 (N_11556,N_10779,N_11102);
nor U11557 (N_11557,N_10853,N_10727);
and U11558 (N_11558,N_10676,N_10916);
xnor U11559 (N_11559,N_10745,N_10921);
and U11560 (N_11560,N_11215,N_10813);
xnor U11561 (N_11561,N_10669,N_11016);
nand U11562 (N_11562,N_10804,N_11125);
and U11563 (N_11563,N_11100,N_11224);
and U11564 (N_11564,N_11030,N_10635);
nand U11565 (N_11565,N_10852,N_11078);
and U11566 (N_11566,N_10904,N_11232);
nand U11567 (N_11567,N_11154,N_10678);
nand U11568 (N_11568,N_10936,N_10795);
nor U11569 (N_11569,N_10682,N_11054);
and U11570 (N_11570,N_11036,N_10628);
nor U11571 (N_11571,N_10897,N_11007);
or U11572 (N_11572,N_10704,N_11003);
nor U11573 (N_11573,N_10878,N_11231);
and U11574 (N_11574,N_11094,N_10667);
and U11575 (N_11575,N_10625,N_11039);
nand U11576 (N_11576,N_10876,N_10758);
nand U11577 (N_11577,N_10977,N_11004);
nand U11578 (N_11578,N_10943,N_10633);
nand U11579 (N_11579,N_11249,N_10985);
xor U11580 (N_11580,N_10875,N_11155);
or U11581 (N_11581,N_11162,N_11192);
nand U11582 (N_11582,N_11015,N_11132);
or U11583 (N_11583,N_10864,N_10754);
nor U11584 (N_11584,N_11105,N_10982);
nor U11585 (N_11585,N_11235,N_10974);
nand U11586 (N_11586,N_11160,N_11143);
nand U11587 (N_11587,N_11221,N_10646);
and U11588 (N_11588,N_11160,N_11102);
nor U11589 (N_11589,N_10962,N_10678);
and U11590 (N_11590,N_10751,N_10885);
xnor U11591 (N_11591,N_10875,N_11086);
or U11592 (N_11592,N_11122,N_10950);
nand U11593 (N_11593,N_10887,N_10870);
nand U11594 (N_11594,N_10670,N_10931);
or U11595 (N_11595,N_10886,N_10892);
or U11596 (N_11596,N_10631,N_10989);
nand U11597 (N_11597,N_11037,N_10811);
nand U11598 (N_11598,N_10982,N_10801);
or U11599 (N_11599,N_10968,N_11125);
nand U11600 (N_11600,N_11188,N_10862);
xnor U11601 (N_11601,N_10833,N_10736);
xor U11602 (N_11602,N_11101,N_10734);
or U11603 (N_11603,N_10920,N_10957);
and U11604 (N_11604,N_11093,N_11213);
xor U11605 (N_11605,N_10828,N_10930);
nor U11606 (N_11606,N_11221,N_11209);
or U11607 (N_11607,N_10715,N_11226);
or U11608 (N_11608,N_10781,N_10997);
nor U11609 (N_11609,N_10853,N_11198);
and U11610 (N_11610,N_11235,N_10835);
nor U11611 (N_11611,N_11100,N_10635);
and U11612 (N_11612,N_10788,N_11169);
or U11613 (N_11613,N_11024,N_10824);
xor U11614 (N_11614,N_10764,N_10628);
xnor U11615 (N_11615,N_10898,N_10730);
nor U11616 (N_11616,N_10676,N_11100);
xnor U11617 (N_11617,N_10787,N_10703);
and U11618 (N_11618,N_10861,N_11125);
xnor U11619 (N_11619,N_11136,N_10800);
nand U11620 (N_11620,N_10768,N_11058);
nor U11621 (N_11621,N_10926,N_10938);
and U11622 (N_11622,N_10947,N_11099);
nand U11623 (N_11623,N_10646,N_10917);
nor U11624 (N_11624,N_11120,N_10852);
nor U11625 (N_11625,N_10813,N_10938);
xnor U11626 (N_11626,N_10727,N_11080);
nor U11627 (N_11627,N_10993,N_10654);
or U11628 (N_11628,N_10744,N_10670);
nand U11629 (N_11629,N_11052,N_11042);
and U11630 (N_11630,N_11021,N_10895);
and U11631 (N_11631,N_10633,N_11066);
and U11632 (N_11632,N_11020,N_11111);
nand U11633 (N_11633,N_11063,N_11055);
xor U11634 (N_11634,N_10630,N_11159);
nand U11635 (N_11635,N_11057,N_11246);
or U11636 (N_11636,N_11091,N_11022);
or U11637 (N_11637,N_11165,N_10816);
nand U11638 (N_11638,N_11149,N_10847);
or U11639 (N_11639,N_10809,N_10651);
nand U11640 (N_11640,N_10855,N_10640);
nand U11641 (N_11641,N_10697,N_11221);
xor U11642 (N_11642,N_10986,N_10682);
nand U11643 (N_11643,N_10682,N_11112);
and U11644 (N_11644,N_10885,N_11189);
and U11645 (N_11645,N_11016,N_11055);
and U11646 (N_11646,N_10964,N_10856);
nor U11647 (N_11647,N_10977,N_10759);
xor U11648 (N_11648,N_10645,N_10885);
nor U11649 (N_11649,N_11051,N_10750);
nand U11650 (N_11650,N_10862,N_10775);
nor U11651 (N_11651,N_11233,N_10999);
or U11652 (N_11652,N_11007,N_10786);
nand U11653 (N_11653,N_11114,N_11161);
and U11654 (N_11654,N_11145,N_10707);
or U11655 (N_11655,N_11102,N_11027);
or U11656 (N_11656,N_11158,N_11116);
nor U11657 (N_11657,N_10810,N_10847);
xor U11658 (N_11658,N_11201,N_10811);
nand U11659 (N_11659,N_11096,N_11196);
nor U11660 (N_11660,N_10990,N_10882);
and U11661 (N_11661,N_11062,N_10697);
xor U11662 (N_11662,N_10850,N_11064);
nand U11663 (N_11663,N_10887,N_10880);
nand U11664 (N_11664,N_10815,N_11086);
xnor U11665 (N_11665,N_11239,N_10802);
or U11666 (N_11666,N_10799,N_11044);
and U11667 (N_11667,N_10858,N_10668);
and U11668 (N_11668,N_10645,N_10816);
xor U11669 (N_11669,N_11235,N_10984);
nor U11670 (N_11670,N_11124,N_11109);
xor U11671 (N_11671,N_11185,N_10777);
or U11672 (N_11672,N_10657,N_10840);
and U11673 (N_11673,N_11079,N_11183);
or U11674 (N_11674,N_10886,N_11185);
nor U11675 (N_11675,N_10893,N_10659);
xnor U11676 (N_11676,N_11215,N_10862);
or U11677 (N_11677,N_11180,N_10922);
or U11678 (N_11678,N_11030,N_10970);
xnor U11679 (N_11679,N_11079,N_10906);
and U11680 (N_11680,N_10842,N_11012);
or U11681 (N_11681,N_11246,N_10809);
nand U11682 (N_11682,N_11107,N_10739);
or U11683 (N_11683,N_10981,N_11222);
nand U11684 (N_11684,N_10936,N_11211);
xnor U11685 (N_11685,N_11100,N_11038);
nor U11686 (N_11686,N_10702,N_11244);
xnor U11687 (N_11687,N_10731,N_10928);
nand U11688 (N_11688,N_10870,N_11074);
or U11689 (N_11689,N_10692,N_11128);
nand U11690 (N_11690,N_10924,N_10823);
nor U11691 (N_11691,N_11193,N_10961);
xor U11692 (N_11692,N_10891,N_11008);
and U11693 (N_11693,N_11196,N_11204);
xor U11694 (N_11694,N_10968,N_11017);
xnor U11695 (N_11695,N_10689,N_10926);
or U11696 (N_11696,N_11192,N_11157);
or U11697 (N_11697,N_10812,N_10882);
xor U11698 (N_11698,N_10687,N_10954);
nor U11699 (N_11699,N_10740,N_10922);
xnor U11700 (N_11700,N_10780,N_10826);
and U11701 (N_11701,N_10784,N_11198);
xor U11702 (N_11702,N_10674,N_10886);
xor U11703 (N_11703,N_11123,N_10774);
nor U11704 (N_11704,N_11163,N_11118);
or U11705 (N_11705,N_10994,N_10776);
nor U11706 (N_11706,N_10936,N_10764);
or U11707 (N_11707,N_10996,N_10802);
nor U11708 (N_11708,N_10820,N_10677);
or U11709 (N_11709,N_10990,N_10651);
nand U11710 (N_11710,N_10660,N_10708);
or U11711 (N_11711,N_11002,N_10990);
and U11712 (N_11712,N_10630,N_10940);
nand U11713 (N_11713,N_11022,N_10716);
nor U11714 (N_11714,N_10814,N_10898);
and U11715 (N_11715,N_10829,N_11028);
xnor U11716 (N_11716,N_10637,N_10691);
xor U11717 (N_11717,N_10951,N_10625);
xnor U11718 (N_11718,N_10753,N_11021);
xor U11719 (N_11719,N_10813,N_11180);
nand U11720 (N_11720,N_10777,N_10860);
or U11721 (N_11721,N_10783,N_10625);
and U11722 (N_11722,N_11025,N_11222);
and U11723 (N_11723,N_11138,N_11148);
or U11724 (N_11724,N_11128,N_11245);
xnor U11725 (N_11725,N_10994,N_11032);
and U11726 (N_11726,N_11135,N_11238);
and U11727 (N_11727,N_10882,N_11001);
or U11728 (N_11728,N_10632,N_10821);
xnor U11729 (N_11729,N_11071,N_10953);
nor U11730 (N_11730,N_10737,N_10987);
nor U11731 (N_11731,N_10925,N_10692);
nand U11732 (N_11732,N_10907,N_10830);
or U11733 (N_11733,N_10790,N_10845);
xor U11734 (N_11734,N_10699,N_10655);
nor U11735 (N_11735,N_10905,N_11099);
or U11736 (N_11736,N_10765,N_10903);
or U11737 (N_11737,N_10917,N_11184);
and U11738 (N_11738,N_10782,N_10628);
or U11739 (N_11739,N_10662,N_11042);
and U11740 (N_11740,N_11247,N_10808);
nand U11741 (N_11741,N_11225,N_10853);
nor U11742 (N_11742,N_10784,N_11052);
nor U11743 (N_11743,N_11119,N_11146);
or U11744 (N_11744,N_10771,N_10898);
nand U11745 (N_11745,N_10927,N_11227);
xor U11746 (N_11746,N_11103,N_10789);
or U11747 (N_11747,N_10976,N_10791);
xnor U11748 (N_11748,N_10813,N_11201);
or U11749 (N_11749,N_10748,N_11136);
nand U11750 (N_11750,N_10874,N_10992);
xor U11751 (N_11751,N_10959,N_11181);
or U11752 (N_11752,N_11162,N_10710);
nand U11753 (N_11753,N_10832,N_10931);
xnor U11754 (N_11754,N_10807,N_11014);
nand U11755 (N_11755,N_11043,N_10997);
nand U11756 (N_11756,N_10924,N_11129);
or U11757 (N_11757,N_10827,N_10958);
or U11758 (N_11758,N_11002,N_11086);
nor U11759 (N_11759,N_11082,N_11227);
nor U11760 (N_11760,N_10990,N_11096);
nand U11761 (N_11761,N_10701,N_11248);
nand U11762 (N_11762,N_11099,N_10695);
nand U11763 (N_11763,N_11015,N_11221);
nor U11764 (N_11764,N_10703,N_11120);
nor U11765 (N_11765,N_10988,N_11059);
nor U11766 (N_11766,N_10677,N_10662);
nor U11767 (N_11767,N_11224,N_10635);
or U11768 (N_11768,N_10930,N_10996);
nor U11769 (N_11769,N_11021,N_10928);
nand U11770 (N_11770,N_10736,N_10874);
and U11771 (N_11771,N_10781,N_10838);
and U11772 (N_11772,N_11181,N_11002);
nand U11773 (N_11773,N_11120,N_10922);
xnor U11774 (N_11774,N_10889,N_10684);
nor U11775 (N_11775,N_10904,N_10747);
or U11776 (N_11776,N_11018,N_10959);
nand U11777 (N_11777,N_10919,N_11166);
or U11778 (N_11778,N_11120,N_11150);
nor U11779 (N_11779,N_10918,N_10960);
nor U11780 (N_11780,N_11232,N_10793);
nand U11781 (N_11781,N_11212,N_10999);
xnor U11782 (N_11782,N_10881,N_10763);
nor U11783 (N_11783,N_11232,N_10990);
nand U11784 (N_11784,N_11165,N_10678);
and U11785 (N_11785,N_10785,N_11208);
nand U11786 (N_11786,N_10719,N_10869);
and U11787 (N_11787,N_10677,N_10737);
xnor U11788 (N_11788,N_10864,N_10742);
or U11789 (N_11789,N_10889,N_10932);
xnor U11790 (N_11790,N_11220,N_10887);
xnor U11791 (N_11791,N_10754,N_10979);
nand U11792 (N_11792,N_10943,N_10828);
or U11793 (N_11793,N_10934,N_10808);
or U11794 (N_11794,N_10773,N_10812);
nor U11795 (N_11795,N_10855,N_10839);
or U11796 (N_11796,N_11049,N_11077);
or U11797 (N_11797,N_10962,N_11018);
and U11798 (N_11798,N_11158,N_10770);
nor U11799 (N_11799,N_11001,N_10867);
nor U11800 (N_11800,N_11236,N_11043);
or U11801 (N_11801,N_11177,N_11006);
nand U11802 (N_11802,N_11069,N_11111);
nor U11803 (N_11803,N_11030,N_11085);
xor U11804 (N_11804,N_10754,N_10896);
or U11805 (N_11805,N_10940,N_11015);
nor U11806 (N_11806,N_10948,N_10716);
nor U11807 (N_11807,N_11200,N_10796);
and U11808 (N_11808,N_10833,N_11083);
or U11809 (N_11809,N_10862,N_10962);
nand U11810 (N_11810,N_11126,N_11001);
or U11811 (N_11811,N_10827,N_10984);
xor U11812 (N_11812,N_11075,N_10627);
and U11813 (N_11813,N_10737,N_11224);
nor U11814 (N_11814,N_10698,N_10808);
nand U11815 (N_11815,N_11202,N_10635);
and U11816 (N_11816,N_10679,N_10790);
nor U11817 (N_11817,N_10998,N_10753);
nor U11818 (N_11818,N_10706,N_10936);
or U11819 (N_11819,N_10956,N_11098);
nor U11820 (N_11820,N_11083,N_10642);
nor U11821 (N_11821,N_11037,N_10669);
nor U11822 (N_11822,N_11102,N_10642);
or U11823 (N_11823,N_11114,N_11223);
nor U11824 (N_11824,N_10662,N_10923);
nand U11825 (N_11825,N_10780,N_11188);
or U11826 (N_11826,N_10768,N_10673);
or U11827 (N_11827,N_10952,N_10759);
or U11828 (N_11828,N_10664,N_10872);
and U11829 (N_11829,N_10890,N_11142);
nand U11830 (N_11830,N_10692,N_10721);
nand U11831 (N_11831,N_10887,N_10735);
nand U11832 (N_11832,N_10887,N_10995);
nor U11833 (N_11833,N_10938,N_10706);
nor U11834 (N_11834,N_10998,N_11067);
and U11835 (N_11835,N_11111,N_10766);
nor U11836 (N_11836,N_10786,N_10962);
or U11837 (N_11837,N_11197,N_10963);
or U11838 (N_11838,N_11186,N_10934);
and U11839 (N_11839,N_10795,N_11180);
or U11840 (N_11840,N_10680,N_11009);
and U11841 (N_11841,N_10901,N_10819);
and U11842 (N_11842,N_10717,N_11183);
xnor U11843 (N_11843,N_10874,N_10965);
xnor U11844 (N_11844,N_10651,N_11035);
nor U11845 (N_11845,N_11118,N_10835);
nor U11846 (N_11846,N_10796,N_11098);
nand U11847 (N_11847,N_10767,N_10837);
xnor U11848 (N_11848,N_10737,N_10641);
nand U11849 (N_11849,N_10638,N_11144);
or U11850 (N_11850,N_11004,N_11182);
nand U11851 (N_11851,N_11008,N_11015);
nor U11852 (N_11852,N_10880,N_11248);
nand U11853 (N_11853,N_11035,N_10823);
xor U11854 (N_11854,N_10752,N_10760);
nand U11855 (N_11855,N_10972,N_10772);
nand U11856 (N_11856,N_10911,N_10888);
nor U11857 (N_11857,N_11141,N_10628);
xor U11858 (N_11858,N_10656,N_10696);
or U11859 (N_11859,N_11126,N_10887);
or U11860 (N_11860,N_10994,N_10756);
xnor U11861 (N_11861,N_10778,N_10932);
and U11862 (N_11862,N_11176,N_10629);
nor U11863 (N_11863,N_10824,N_10685);
xor U11864 (N_11864,N_11117,N_11056);
and U11865 (N_11865,N_11139,N_11239);
or U11866 (N_11866,N_10718,N_11115);
nor U11867 (N_11867,N_10818,N_11243);
and U11868 (N_11868,N_10795,N_11039);
xnor U11869 (N_11869,N_10840,N_11143);
xnor U11870 (N_11870,N_11169,N_10851);
and U11871 (N_11871,N_10786,N_10918);
nor U11872 (N_11872,N_11040,N_11203);
nor U11873 (N_11873,N_10768,N_10882);
or U11874 (N_11874,N_11173,N_11130);
nand U11875 (N_11875,N_11583,N_11785);
xor U11876 (N_11876,N_11674,N_11362);
nand U11877 (N_11877,N_11816,N_11410);
nor U11878 (N_11878,N_11778,N_11868);
xnor U11879 (N_11879,N_11408,N_11495);
or U11880 (N_11880,N_11597,N_11861);
and U11881 (N_11881,N_11568,N_11694);
nor U11882 (N_11882,N_11565,N_11270);
nand U11883 (N_11883,N_11775,N_11588);
and U11884 (N_11884,N_11442,N_11275);
nor U11885 (N_11885,N_11279,N_11557);
or U11886 (N_11886,N_11676,N_11625);
nand U11887 (N_11887,N_11691,N_11782);
nand U11888 (N_11888,N_11379,N_11686);
nor U11889 (N_11889,N_11830,N_11504);
nand U11890 (N_11890,N_11373,N_11315);
nor U11891 (N_11891,N_11759,N_11751);
or U11892 (N_11892,N_11455,N_11754);
nand U11893 (N_11893,N_11327,N_11571);
nor U11894 (N_11894,N_11470,N_11548);
xnor U11895 (N_11895,N_11267,N_11652);
and U11896 (N_11896,N_11735,N_11556);
and U11897 (N_11897,N_11731,N_11789);
nor U11898 (N_11898,N_11726,N_11558);
and U11899 (N_11899,N_11609,N_11390);
xor U11900 (N_11900,N_11532,N_11632);
nor U11901 (N_11901,N_11836,N_11675);
or U11902 (N_11902,N_11607,N_11377);
xor U11903 (N_11903,N_11357,N_11440);
and U11904 (N_11904,N_11699,N_11400);
and U11905 (N_11905,N_11630,N_11765);
nor U11906 (N_11906,N_11288,N_11569);
xor U11907 (N_11907,N_11320,N_11596);
or U11908 (N_11908,N_11446,N_11344);
nor U11909 (N_11909,N_11684,N_11473);
or U11910 (N_11910,N_11781,N_11866);
nor U11911 (N_11911,N_11807,N_11303);
nand U11912 (N_11912,N_11843,N_11654);
and U11913 (N_11913,N_11516,N_11394);
and U11914 (N_11914,N_11281,N_11380);
and U11915 (N_11915,N_11813,N_11773);
nand U11916 (N_11916,N_11546,N_11544);
and U11917 (N_11917,N_11323,N_11734);
and U11918 (N_11918,N_11697,N_11559);
nor U11919 (N_11919,N_11431,N_11859);
and U11920 (N_11920,N_11517,N_11856);
nor U11921 (N_11921,N_11586,N_11295);
nand U11922 (N_11922,N_11852,N_11550);
or U11923 (N_11923,N_11587,N_11450);
nor U11924 (N_11924,N_11695,N_11405);
and U11925 (N_11925,N_11439,N_11633);
or U11926 (N_11926,N_11515,N_11724);
xnor U11927 (N_11927,N_11808,N_11743);
and U11928 (N_11928,N_11522,N_11461);
nor U11929 (N_11929,N_11414,N_11257);
xnor U11930 (N_11930,N_11776,N_11612);
nand U11931 (N_11931,N_11613,N_11831);
or U11932 (N_11932,N_11576,N_11733);
nand U11933 (N_11933,N_11825,N_11398);
or U11934 (N_11934,N_11783,N_11779);
nand U11935 (N_11935,N_11619,N_11462);
nor U11936 (N_11936,N_11551,N_11269);
and U11937 (N_11937,N_11812,N_11356);
nand U11938 (N_11938,N_11667,N_11611);
xor U11939 (N_11939,N_11304,N_11449);
and U11940 (N_11940,N_11709,N_11512);
xnor U11941 (N_11941,N_11715,N_11797);
nand U11942 (N_11942,N_11575,N_11484);
and U11943 (N_11943,N_11845,N_11372);
or U11944 (N_11944,N_11313,N_11435);
or U11945 (N_11945,N_11767,N_11665);
xnor U11946 (N_11946,N_11501,N_11722);
xor U11947 (N_11947,N_11293,N_11788);
and U11948 (N_11948,N_11475,N_11423);
xnor U11949 (N_11949,N_11755,N_11650);
and U11950 (N_11950,N_11786,N_11780);
xnor U11951 (N_11951,N_11840,N_11605);
and U11952 (N_11952,N_11753,N_11865);
xnor U11953 (N_11953,N_11407,N_11381);
nor U11954 (N_11954,N_11530,N_11794);
and U11955 (N_11955,N_11302,N_11520);
nand U11956 (N_11956,N_11509,N_11508);
or U11957 (N_11957,N_11309,N_11490);
and U11958 (N_11958,N_11480,N_11749);
nand U11959 (N_11959,N_11680,N_11326);
nand U11960 (N_11960,N_11430,N_11272);
nand U11961 (N_11961,N_11614,N_11260);
nor U11962 (N_11962,N_11453,N_11713);
and U11963 (N_11963,N_11454,N_11447);
and U11964 (N_11964,N_11796,N_11493);
xnor U11965 (N_11965,N_11581,N_11488);
xnor U11966 (N_11966,N_11312,N_11354);
nor U11967 (N_11967,N_11396,N_11636);
xnor U11968 (N_11968,N_11818,N_11294);
or U11969 (N_11969,N_11547,N_11672);
nor U11970 (N_11970,N_11485,N_11253);
nor U11971 (N_11971,N_11671,N_11760);
nand U11972 (N_11972,N_11638,N_11815);
nor U11973 (N_11973,N_11496,N_11723);
nand U11974 (N_11974,N_11688,N_11701);
or U11975 (N_11975,N_11535,N_11523);
nand U11976 (N_11976,N_11339,N_11623);
nor U11977 (N_11977,N_11573,N_11385);
nor U11978 (N_11978,N_11710,N_11404);
nand U11979 (N_11979,N_11582,N_11376);
and U11980 (N_11980,N_11719,N_11335);
or U11981 (N_11981,N_11444,N_11841);
xnor U11982 (N_11982,N_11441,N_11629);
nand U11983 (N_11983,N_11682,N_11443);
or U11984 (N_11984,N_11764,N_11791);
or U11985 (N_11985,N_11799,N_11527);
or U11986 (N_11986,N_11858,N_11664);
nand U11987 (N_11987,N_11353,N_11562);
nand U11988 (N_11988,N_11746,N_11502);
or U11989 (N_11989,N_11748,N_11298);
nand U11990 (N_11990,N_11591,N_11805);
nand U11991 (N_11991,N_11685,N_11615);
xor U11992 (N_11992,N_11850,N_11716);
nand U11993 (N_11993,N_11345,N_11598);
nand U11994 (N_11994,N_11463,N_11622);
or U11995 (N_11995,N_11601,N_11540);
xnor U11996 (N_11996,N_11666,N_11563);
and U11997 (N_11997,N_11683,N_11677);
nor U11998 (N_11998,N_11262,N_11321);
nor U11999 (N_11999,N_11482,N_11857);
nor U12000 (N_12000,N_11590,N_11403);
xnor U12001 (N_12001,N_11624,N_11459);
nor U12002 (N_12002,N_11338,N_11521);
and U12003 (N_12003,N_11437,N_11310);
and U12004 (N_12004,N_11740,N_11471);
and U12005 (N_12005,N_11584,N_11707);
and U12006 (N_12006,N_11538,N_11367);
and U12007 (N_12007,N_11763,N_11698);
nor U12008 (N_12008,N_11874,N_11341);
nor U12009 (N_12009,N_11314,N_11739);
xor U12010 (N_12010,N_11851,N_11416);
or U12011 (N_12011,N_11474,N_11600);
nand U12012 (N_12012,N_11280,N_11478);
or U12013 (N_12013,N_11771,N_11700);
nand U12014 (N_12014,N_11711,N_11351);
and U12015 (N_12015,N_11616,N_11670);
and U12016 (N_12016,N_11458,N_11424);
nand U12017 (N_12017,N_11251,N_11640);
nand U12018 (N_12018,N_11549,N_11593);
and U12019 (N_12019,N_11567,N_11278);
or U12020 (N_12020,N_11814,N_11503);
and U12021 (N_12021,N_11266,N_11769);
or U12022 (N_12022,N_11827,N_11727);
nand U12023 (N_12023,N_11784,N_11330);
or U12024 (N_12024,N_11369,N_11660);
nor U12025 (N_12025,N_11290,N_11511);
nor U12026 (N_12026,N_11637,N_11445);
xor U12027 (N_12027,N_11752,N_11491);
nor U12028 (N_12028,N_11645,N_11787);
and U12029 (N_12029,N_11679,N_11661);
nand U12030 (N_12030,N_11655,N_11854);
and U12031 (N_12031,N_11274,N_11250);
nor U12032 (N_12032,N_11301,N_11420);
nor U12033 (N_12033,N_11844,N_11292);
nor U12034 (N_12034,N_11595,N_11456);
xor U12035 (N_12035,N_11428,N_11276);
or U12036 (N_12036,N_11870,N_11331);
or U12037 (N_12037,N_11286,N_11536);
nor U12038 (N_12038,N_11252,N_11777);
nor U12039 (N_12039,N_11687,N_11651);
nor U12040 (N_12040,N_11525,N_11417);
nor U12041 (N_12041,N_11421,N_11631);
nand U12042 (N_12042,N_11757,N_11307);
and U12043 (N_12043,N_11318,N_11533);
nor U12044 (N_12044,N_11737,N_11627);
and U12045 (N_12045,N_11368,N_11359);
or U12046 (N_12046,N_11564,N_11506);
or U12047 (N_12047,N_11678,N_11849);
or U12048 (N_12048,N_11519,N_11610);
nand U12049 (N_12049,N_11297,N_11452);
or U12050 (N_12050,N_11669,N_11529);
xnor U12051 (N_12051,N_11388,N_11834);
or U12052 (N_12052,N_11510,N_11822);
and U12053 (N_12053,N_11277,N_11617);
nand U12054 (N_12054,N_11641,N_11347);
and U12055 (N_12055,N_11486,N_11299);
xnor U12056 (N_12056,N_11729,N_11690);
and U12057 (N_12057,N_11864,N_11702);
or U12058 (N_12058,N_11255,N_11693);
nand U12059 (N_12059,N_11393,N_11324);
nor U12060 (N_12060,N_11489,N_11392);
nand U12061 (N_12061,N_11464,N_11422);
xnor U12062 (N_12062,N_11360,N_11378);
and U12063 (N_12063,N_11258,N_11770);
nor U12064 (N_12064,N_11725,N_11528);
xnor U12065 (N_12065,N_11663,N_11662);
xor U12066 (N_12066,N_11837,N_11507);
or U12067 (N_12067,N_11448,N_11264);
and U12068 (N_12068,N_11653,N_11839);
and U12069 (N_12069,N_11804,N_11429);
and U12070 (N_12070,N_11518,N_11658);
xnor U12071 (N_12071,N_11853,N_11401);
xor U12072 (N_12072,N_11479,N_11855);
xor U12073 (N_12073,N_11657,N_11499);
or U12074 (N_12074,N_11412,N_11720);
and U12075 (N_12075,N_11761,N_11513);
nor U12076 (N_12076,N_11333,N_11524);
xor U12077 (N_12077,N_11766,N_11537);
or U12078 (N_12078,N_11863,N_11768);
and U12079 (N_12079,N_11329,N_11375);
nand U12080 (N_12080,N_11644,N_11539);
xnor U12081 (N_12081,N_11626,N_11284);
nor U12082 (N_12082,N_11409,N_11306);
nor U12083 (N_12083,N_11289,N_11265);
nor U12084 (N_12084,N_11311,N_11634);
nor U12085 (N_12085,N_11317,N_11319);
and U12086 (N_12086,N_11566,N_11316);
xnor U12087 (N_12087,N_11366,N_11871);
nand U12088 (N_12088,N_11860,N_11296);
nand U12089 (N_12089,N_11334,N_11714);
and U12090 (N_12090,N_11426,N_11824);
nor U12091 (N_12091,N_11828,N_11476);
xnor U12092 (N_12092,N_11842,N_11427);
nor U12093 (N_12093,N_11494,N_11340);
or U12094 (N_12094,N_11806,N_11732);
nor U12095 (N_12095,N_11343,N_11425);
xnor U12096 (N_12096,N_11432,N_11656);
nor U12097 (N_12097,N_11618,N_11820);
xnor U12098 (N_12098,N_11742,N_11692);
and U12099 (N_12099,N_11497,N_11673);
nand U12100 (N_12100,N_11399,N_11332);
or U12101 (N_12101,N_11741,N_11337);
nand U12102 (N_12102,N_11589,N_11552);
xor U12103 (N_12103,N_11592,N_11395);
nor U12104 (N_12104,N_11358,N_11603);
xor U12105 (N_12105,N_11873,N_11460);
xor U12106 (N_12106,N_11371,N_11554);
nor U12107 (N_12107,N_11261,N_11717);
xnor U12108 (N_12108,N_11580,N_11469);
xor U12109 (N_12109,N_11635,N_11689);
xor U12110 (N_12110,N_11457,N_11553);
nor U12111 (N_12111,N_11604,N_11728);
nor U12112 (N_12112,N_11659,N_11826);
or U12113 (N_12113,N_11704,N_11649);
and U12114 (N_12114,N_11492,N_11397);
nand U12115 (N_12115,N_11572,N_11418);
or U12116 (N_12116,N_11336,N_11772);
or U12117 (N_12117,N_11829,N_11833);
and U12118 (N_12118,N_11570,N_11795);
xnor U12119 (N_12119,N_11481,N_11413);
nor U12120 (N_12120,N_11706,N_11747);
or U12121 (N_12121,N_11545,N_11579);
and U12122 (N_12122,N_11594,N_11703);
nand U12123 (N_12123,N_11736,N_11792);
nor U12124 (N_12124,N_11467,N_11578);
nand U12125 (N_12125,N_11500,N_11477);
nor U12126 (N_12126,N_11483,N_11468);
nand U12127 (N_12127,N_11531,N_11869);
nor U12128 (N_12128,N_11273,N_11346);
or U12129 (N_12129,N_11823,N_11415);
nor U12130 (N_12130,N_11387,N_11821);
xor U12131 (N_12131,N_11639,N_11465);
nand U12132 (N_12132,N_11608,N_11526);
xor U12133 (N_12133,N_11803,N_11790);
and U12134 (N_12134,N_11451,N_11308);
and U12135 (N_12135,N_11287,N_11819);
nand U12136 (N_12136,N_11758,N_11348);
nor U12137 (N_12137,N_11560,N_11648);
or U12138 (N_12138,N_11411,N_11291);
nand U12139 (N_12139,N_11389,N_11718);
nor U12140 (N_12140,N_11283,N_11832);
and U12141 (N_12141,N_11466,N_11774);
nand U12142 (N_12142,N_11433,N_11542);
nand U12143 (N_12143,N_11364,N_11342);
nand U12144 (N_12144,N_11352,N_11300);
xnor U12145 (N_12145,N_11708,N_11374);
nor U12146 (N_12146,N_11434,N_11259);
xnor U12147 (N_12147,N_11721,N_11862);
or U12148 (N_12148,N_11577,N_11505);
nand U12149 (N_12149,N_11534,N_11802);
nor U12150 (N_12150,N_11472,N_11282);
xnor U12151 (N_12151,N_11256,N_11744);
or U12152 (N_12152,N_11599,N_11487);
or U12153 (N_12153,N_11800,N_11681);
xnor U12154 (N_12154,N_11574,N_11705);
or U12155 (N_12155,N_11730,N_11406);
and U12156 (N_12156,N_11514,N_11541);
xor U12157 (N_12157,N_11322,N_11436);
nor U12158 (N_12158,N_11254,N_11809);
or U12159 (N_12159,N_11355,N_11391);
nand U12160 (N_12160,N_11384,N_11263);
nand U12161 (N_12161,N_11848,N_11647);
xnor U12162 (N_12162,N_11543,N_11756);
nand U12163 (N_12163,N_11555,N_11419);
or U12164 (N_12164,N_11602,N_11643);
xnor U12165 (N_12165,N_11646,N_11606);
xnor U12166 (N_12166,N_11383,N_11585);
nand U12167 (N_12167,N_11402,N_11872);
and U12168 (N_12168,N_11811,N_11365);
and U12169 (N_12169,N_11642,N_11350);
and U12170 (N_12170,N_11798,N_11498);
nor U12171 (N_12171,N_11382,N_11285);
xor U12172 (N_12172,N_11668,N_11328);
xor U12173 (N_12173,N_11271,N_11846);
nor U12174 (N_12174,N_11835,N_11325);
xor U12175 (N_12175,N_11712,N_11438);
xor U12176 (N_12176,N_11349,N_11838);
nor U12177 (N_12177,N_11847,N_11305);
nand U12178 (N_12178,N_11620,N_11801);
nor U12179 (N_12179,N_11745,N_11793);
and U12180 (N_12180,N_11361,N_11363);
or U12181 (N_12181,N_11810,N_11370);
xnor U12182 (N_12182,N_11738,N_11817);
nor U12183 (N_12183,N_11628,N_11561);
or U12184 (N_12184,N_11621,N_11268);
xnor U12185 (N_12185,N_11386,N_11750);
xor U12186 (N_12186,N_11762,N_11696);
and U12187 (N_12187,N_11867,N_11813);
and U12188 (N_12188,N_11362,N_11353);
and U12189 (N_12189,N_11349,N_11328);
nor U12190 (N_12190,N_11781,N_11519);
xnor U12191 (N_12191,N_11720,N_11609);
or U12192 (N_12192,N_11552,N_11831);
and U12193 (N_12193,N_11360,N_11437);
nor U12194 (N_12194,N_11760,N_11502);
and U12195 (N_12195,N_11413,N_11819);
xnor U12196 (N_12196,N_11547,N_11322);
or U12197 (N_12197,N_11648,N_11827);
xnor U12198 (N_12198,N_11439,N_11459);
and U12199 (N_12199,N_11392,N_11300);
nand U12200 (N_12200,N_11593,N_11449);
or U12201 (N_12201,N_11482,N_11349);
or U12202 (N_12202,N_11553,N_11779);
nand U12203 (N_12203,N_11603,N_11460);
nor U12204 (N_12204,N_11401,N_11474);
and U12205 (N_12205,N_11596,N_11563);
and U12206 (N_12206,N_11446,N_11260);
xnor U12207 (N_12207,N_11330,N_11615);
nor U12208 (N_12208,N_11747,N_11286);
or U12209 (N_12209,N_11473,N_11511);
nor U12210 (N_12210,N_11313,N_11326);
nand U12211 (N_12211,N_11737,N_11549);
or U12212 (N_12212,N_11731,N_11294);
xnor U12213 (N_12213,N_11847,N_11584);
xor U12214 (N_12214,N_11740,N_11434);
nand U12215 (N_12215,N_11524,N_11719);
and U12216 (N_12216,N_11596,N_11491);
nand U12217 (N_12217,N_11599,N_11859);
and U12218 (N_12218,N_11695,N_11592);
nor U12219 (N_12219,N_11614,N_11600);
xor U12220 (N_12220,N_11548,N_11482);
or U12221 (N_12221,N_11587,N_11805);
nor U12222 (N_12222,N_11482,N_11822);
xnor U12223 (N_12223,N_11439,N_11741);
xnor U12224 (N_12224,N_11754,N_11449);
and U12225 (N_12225,N_11616,N_11258);
and U12226 (N_12226,N_11333,N_11307);
nand U12227 (N_12227,N_11273,N_11309);
nand U12228 (N_12228,N_11316,N_11616);
and U12229 (N_12229,N_11719,N_11379);
and U12230 (N_12230,N_11606,N_11321);
or U12231 (N_12231,N_11780,N_11714);
and U12232 (N_12232,N_11547,N_11819);
or U12233 (N_12233,N_11352,N_11366);
nand U12234 (N_12234,N_11617,N_11565);
nand U12235 (N_12235,N_11382,N_11843);
nor U12236 (N_12236,N_11661,N_11416);
nand U12237 (N_12237,N_11777,N_11505);
and U12238 (N_12238,N_11413,N_11595);
and U12239 (N_12239,N_11723,N_11609);
nand U12240 (N_12240,N_11669,N_11374);
nand U12241 (N_12241,N_11580,N_11411);
xor U12242 (N_12242,N_11703,N_11802);
nand U12243 (N_12243,N_11581,N_11348);
nor U12244 (N_12244,N_11341,N_11473);
xor U12245 (N_12245,N_11535,N_11344);
nand U12246 (N_12246,N_11775,N_11735);
nand U12247 (N_12247,N_11723,N_11866);
nor U12248 (N_12248,N_11448,N_11386);
nand U12249 (N_12249,N_11850,N_11335);
nand U12250 (N_12250,N_11794,N_11338);
xnor U12251 (N_12251,N_11505,N_11723);
nor U12252 (N_12252,N_11735,N_11305);
xnor U12253 (N_12253,N_11850,N_11573);
and U12254 (N_12254,N_11729,N_11635);
xnor U12255 (N_12255,N_11306,N_11340);
and U12256 (N_12256,N_11317,N_11373);
and U12257 (N_12257,N_11824,N_11740);
or U12258 (N_12258,N_11746,N_11495);
nand U12259 (N_12259,N_11637,N_11811);
xnor U12260 (N_12260,N_11534,N_11719);
nor U12261 (N_12261,N_11523,N_11428);
or U12262 (N_12262,N_11630,N_11671);
and U12263 (N_12263,N_11580,N_11386);
and U12264 (N_12264,N_11463,N_11438);
and U12265 (N_12265,N_11540,N_11861);
and U12266 (N_12266,N_11464,N_11761);
nor U12267 (N_12267,N_11865,N_11293);
nand U12268 (N_12268,N_11845,N_11403);
and U12269 (N_12269,N_11803,N_11657);
and U12270 (N_12270,N_11663,N_11378);
or U12271 (N_12271,N_11333,N_11758);
or U12272 (N_12272,N_11501,N_11618);
nand U12273 (N_12273,N_11768,N_11615);
and U12274 (N_12274,N_11547,N_11298);
nand U12275 (N_12275,N_11529,N_11731);
and U12276 (N_12276,N_11384,N_11535);
and U12277 (N_12277,N_11531,N_11496);
or U12278 (N_12278,N_11556,N_11501);
or U12279 (N_12279,N_11336,N_11735);
and U12280 (N_12280,N_11691,N_11724);
nor U12281 (N_12281,N_11424,N_11267);
or U12282 (N_12282,N_11461,N_11502);
nand U12283 (N_12283,N_11301,N_11804);
nor U12284 (N_12284,N_11507,N_11627);
nand U12285 (N_12285,N_11338,N_11801);
nand U12286 (N_12286,N_11614,N_11557);
nand U12287 (N_12287,N_11478,N_11591);
nor U12288 (N_12288,N_11625,N_11559);
and U12289 (N_12289,N_11266,N_11639);
xor U12290 (N_12290,N_11746,N_11402);
or U12291 (N_12291,N_11749,N_11389);
and U12292 (N_12292,N_11848,N_11601);
or U12293 (N_12293,N_11567,N_11533);
or U12294 (N_12294,N_11563,N_11753);
nor U12295 (N_12295,N_11601,N_11419);
and U12296 (N_12296,N_11621,N_11545);
xor U12297 (N_12297,N_11294,N_11667);
xor U12298 (N_12298,N_11280,N_11442);
and U12299 (N_12299,N_11751,N_11481);
nand U12300 (N_12300,N_11506,N_11780);
or U12301 (N_12301,N_11778,N_11328);
or U12302 (N_12302,N_11261,N_11570);
nor U12303 (N_12303,N_11646,N_11512);
or U12304 (N_12304,N_11253,N_11439);
nor U12305 (N_12305,N_11642,N_11666);
nand U12306 (N_12306,N_11259,N_11436);
nor U12307 (N_12307,N_11789,N_11302);
nor U12308 (N_12308,N_11301,N_11593);
xnor U12309 (N_12309,N_11599,N_11763);
and U12310 (N_12310,N_11773,N_11747);
nand U12311 (N_12311,N_11593,N_11259);
nor U12312 (N_12312,N_11313,N_11668);
xor U12313 (N_12313,N_11855,N_11285);
xnor U12314 (N_12314,N_11595,N_11478);
nand U12315 (N_12315,N_11550,N_11406);
or U12316 (N_12316,N_11541,N_11842);
nor U12317 (N_12317,N_11329,N_11341);
and U12318 (N_12318,N_11252,N_11284);
xnor U12319 (N_12319,N_11663,N_11326);
and U12320 (N_12320,N_11434,N_11557);
xnor U12321 (N_12321,N_11803,N_11532);
xor U12322 (N_12322,N_11567,N_11765);
and U12323 (N_12323,N_11609,N_11794);
or U12324 (N_12324,N_11506,N_11320);
xnor U12325 (N_12325,N_11417,N_11632);
nand U12326 (N_12326,N_11442,N_11481);
xor U12327 (N_12327,N_11795,N_11294);
or U12328 (N_12328,N_11384,N_11469);
nand U12329 (N_12329,N_11776,N_11407);
or U12330 (N_12330,N_11389,N_11377);
and U12331 (N_12331,N_11677,N_11846);
xor U12332 (N_12332,N_11604,N_11703);
nand U12333 (N_12333,N_11373,N_11744);
nor U12334 (N_12334,N_11296,N_11538);
nor U12335 (N_12335,N_11509,N_11588);
or U12336 (N_12336,N_11418,N_11610);
and U12337 (N_12337,N_11653,N_11290);
and U12338 (N_12338,N_11372,N_11360);
nor U12339 (N_12339,N_11532,N_11664);
nand U12340 (N_12340,N_11517,N_11616);
xor U12341 (N_12341,N_11641,N_11264);
nand U12342 (N_12342,N_11332,N_11338);
nor U12343 (N_12343,N_11743,N_11795);
nand U12344 (N_12344,N_11250,N_11484);
or U12345 (N_12345,N_11672,N_11539);
and U12346 (N_12346,N_11589,N_11548);
nor U12347 (N_12347,N_11825,N_11779);
and U12348 (N_12348,N_11475,N_11768);
nor U12349 (N_12349,N_11468,N_11607);
nand U12350 (N_12350,N_11594,N_11324);
xnor U12351 (N_12351,N_11298,N_11468);
or U12352 (N_12352,N_11509,N_11356);
and U12353 (N_12353,N_11822,N_11628);
xnor U12354 (N_12354,N_11818,N_11404);
and U12355 (N_12355,N_11464,N_11868);
and U12356 (N_12356,N_11479,N_11418);
nand U12357 (N_12357,N_11567,N_11613);
nor U12358 (N_12358,N_11448,N_11733);
xnor U12359 (N_12359,N_11367,N_11832);
nor U12360 (N_12360,N_11649,N_11660);
nor U12361 (N_12361,N_11766,N_11320);
or U12362 (N_12362,N_11434,N_11340);
and U12363 (N_12363,N_11818,N_11500);
nor U12364 (N_12364,N_11368,N_11828);
or U12365 (N_12365,N_11759,N_11740);
xor U12366 (N_12366,N_11397,N_11490);
xor U12367 (N_12367,N_11796,N_11802);
and U12368 (N_12368,N_11619,N_11376);
nor U12369 (N_12369,N_11264,N_11822);
or U12370 (N_12370,N_11258,N_11301);
and U12371 (N_12371,N_11555,N_11667);
xnor U12372 (N_12372,N_11541,N_11755);
nand U12373 (N_12373,N_11383,N_11483);
or U12374 (N_12374,N_11484,N_11266);
nand U12375 (N_12375,N_11829,N_11834);
and U12376 (N_12376,N_11308,N_11582);
nand U12377 (N_12377,N_11769,N_11357);
nor U12378 (N_12378,N_11582,N_11862);
xnor U12379 (N_12379,N_11313,N_11741);
nor U12380 (N_12380,N_11269,N_11778);
or U12381 (N_12381,N_11603,N_11523);
nor U12382 (N_12382,N_11659,N_11375);
nor U12383 (N_12383,N_11673,N_11594);
or U12384 (N_12384,N_11405,N_11529);
and U12385 (N_12385,N_11614,N_11386);
nand U12386 (N_12386,N_11548,N_11855);
xnor U12387 (N_12387,N_11301,N_11470);
and U12388 (N_12388,N_11639,N_11461);
nand U12389 (N_12389,N_11564,N_11764);
nand U12390 (N_12390,N_11857,N_11500);
nand U12391 (N_12391,N_11311,N_11612);
nand U12392 (N_12392,N_11826,N_11572);
xor U12393 (N_12393,N_11530,N_11451);
xor U12394 (N_12394,N_11286,N_11752);
nand U12395 (N_12395,N_11677,N_11699);
or U12396 (N_12396,N_11809,N_11304);
nand U12397 (N_12397,N_11700,N_11366);
or U12398 (N_12398,N_11417,N_11291);
nor U12399 (N_12399,N_11769,N_11378);
nand U12400 (N_12400,N_11697,N_11809);
xnor U12401 (N_12401,N_11326,N_11852);
and U12402 (N_12402,N_11710,N_11658);
nor U12403 (N_12403,N_11735,N_11759);
or U12404 (N_12404,N_11740,N_11726);
or U12405 (N_12405,N_11862,N_11595);
and U12406 (N_12406,N_11692,N_11349);
nor U12407 (N_12407,N_11746,N_11672);
nor U12408 (N_12408,N_11551,N_11360);
and U12409 (N_12409,N_11667,N_11609);
nor U12410 (N_12410,N_11863,N_11705);
or U12411 (N_12411,N_11618,N_11601);
nor U12412 (N_12412,N_11557,N_11369);
or U12413 (N_12413,N_11473,N_11693);
xnor U12414 (N_12414,N_11314,N_11749);
and U12415 (N_12415,N_11622,N_11633);
or U12416 (N_12416,N_11423,N_11539);
and U12417 (N_12417,N_11701,N_11287);
or U12418 (N_12418,N_11310,N_11260);
or U12419 (N_12419,N_11804,N_11738);
xor U12420 (N_12420,N_11564,N_11250);
xnor U12421 (N_12421,N_11299,N_11356);
xnor U12422 (N_12422,N_11266,N_11715);
nor U12423 (N_12423,N_11701,N_11566);
or U12424 (N_12424,N_11727,N_11443);
xnor U12425 (N_12425,N_11441,N_11785);
or U12426 (N_12426,N_11843,N_11833);
and U12427 (N_12427,N_11531,N_11753);
xnor U12428 (N_12428,N_11319,N_11619);
or U12429 (N_12429,N_11469,N_11739);
nor U12430 (N_12430,N_11424,N_11381);
nand U12431 (N_12431,N_11298,N_11264);
or U12432 (N_12432,N_11669,N_11831);
and U12433 (N_12433,N_11538,N_11588);
xnor U12434 (N_12434,N_11737,N_11508);
xnor U12435 (N_12435,N_11305,N_11272);
xor U12436 (N_12436,N_11354,N_11557);
and U12437 (N_12437,N_11657,N_11592);
and U12438 (N_12438,N_11285,N_11583);
nand U12439 (N_12439,N_11327,N_11645);
nand U12440 (N_12440,N_11371,N_11643);
and U12441 (N_12441,N_11434,N_11281);
xnor U12442 (N_12442,N_11580,N_11538);
or U12443 (N_12443,N_11548,N_11662);
nand U12444 (N_12444,N_11424,N_11620);
and U12445 (N_12445,N_11573,N_11858);
or U12446 (N_12446,N_11718,N_11471);
and U12447 (N_12447,N_11610,N_11688);
nand U12448 (N_12448,N_11486,N_11322);
nand U12449 (N_12449,N_11668,N_11351);
xnor U12450 (N_12450,N_11768,N_11477);
xnor U12451 (N_12451,N_11528,N_11312);
and U12452 (N_12452,N_11805,N_11633);
xor U12453 (N_12453,N_11868,N_11451);
xnor U12454 (N_12454,N_11556,N_11871);
nand U12455 (N_12455,N_11708,N_11348);
xnor U12456 (N_12456,N_11717,N_11832);
nor U12457 (N_12457,N_11514,N_11436);
xor U12458 (N_12458,N_11344,N_11514);
nor U12459 (N_12459,N_11729,N_11574);
nor U12460 (N_12460,N_11312,N_11755);
nor U12461 (N_12461,N_11834,N_11729);
nand U12462 (N_12462,N_11646,N_11674);
or U12463 (N_12463,N_11454,N_11865);
and U12464 (N_12464,N_11785,N_11598);
xor U12465 (N_12465,N_11258,N_11668);
or U12466 (N_12466,N_11860,N_11385);
nor U12467 (N_12467,N_11543,N_11290);
nor U12468 (N_12468,N_11264,N_11554);
or U12469 (N_12469,N_11608,N_11458);
and U12470 (N_12470,N_11551,N_11404);
xnor U12471 (N_12471,N_11275,N_11729);
and U12472 (N_12472,N_11642,N_11572);
nand U12473 (N_12473,N_11350,N_11724);
or U12474 (N_12474,N_11806,N_11252);
xor U12475 (N_12475,N_11292,N_11735);
or U12476 (N_12476,N_11851,N_11592);
or U12477 (N_12477,N_11741,N_11841);
xor U12478 (N_12478,N_11475,N_11670);
nand U12479 (N_12479,N_11503,N_11604);
and U12480 (N_12480,N_11784,N_11495);
nor U12481 (N_12481,N_11760,N_11687);
nand U12482 (N_12482,N_11578,N_11735);
or U12483 (N_12483,N_11854,N_11558);
or U12484 (N_12484,N_11700,N_11660);
nor U12485 (N_12485,N_11758,N_11396);
nor U12486 (N_12486,N_11459,N_11849);
nor U12487 (N_12487,N_11408,N_11646);
and U12488 (N_12488,N_11655,N_11475);
nand U12489 (N_12489,N_11850,N_11611);
and U12490 (N_12490,N_11297,N_11739);
nand U12491 (N_12491,N_11265,N_11725);
and U12492 (N_12492,N_11277,N_11681);
or U12493 (N_12493,N_11730,N_11621);
and U12494 (N_12494,N_11743,N_11494);
or U12495 (N_12495,N_11264,N_11344);
xor U12496 (N_12496,N_11535,N_11513);
and U12497 (N_12497,N_11585,N_11836);
nand U12498 (N_12498,N_11444,N_11443);
nor U12499 (N_12499,N_11571,N_11660);
nand U12500 (N_12500,N_12242,N_12474);
xor U12501 (N_12501,N_12140,N_12068);
xnor U12502 (N_12502,N_12454,N_12138);
and U12503 (N_12503,N_11946,N_12208);
and U12504 (N_12504,N_12216,N_11902);
and U12505 (N_12505,N_11951,N_12088);
xnor U12506 (N_12506,N_11958,N_12086);
nor U12507 (N_12507,N_11997,N_12002);
or U12508 (N_12508,N_11883,N_12286);
and U12509 (N_12509,N_12029,N_12435);
nand U12510 (N_12510,N_12410,N_12425);
nand U12511 (N_12511,N_12494,N_12129);
or U12512 (N_12512,N_12337,N_12482);
or U12513 (N_12513,N_12241,N_12119);
nand U12514 (N_12514,N_11921,N_12195);
and U12515 (N_12515,N_12205,N_12288);
nor U12516 (N_12516,N_11929,N_12020);
nor U12517 (N_12517,N_12325,N_11894);
xor U12518 (N_12518,N_11897,N_12308);
and U12519 (N_12519,N_12420,N_12437);
nand U12520 (N_12520,N_12063,N_12496);
and U12521 (N_12521,N_11896,N_12274);
or U12522 (N_12522,N_12409,N_12266);
nand U12523 (N_12523,N_12073,N_12185);
and U12524 (N_12524,N_12219,N_12051);
nor U12525 (N_12525,N_11887,N_12270);
nor U12526 (N_12526,N_12180,N_12207);
or U12527 (N_12527,N_12317,N_12191);
xor U12528 (N_12528,N_11910,N_12391);
and U12529 (N_12529,N_11957,N_12400);
nor U12530 (N_12530,N_11924,N_12309);
or U12531 (N_12531,N_12121,N_11901);
and U12532 (N_12532,N_12285,N_12457);
or U12533 (N_12533,N_12374,N_12467);
xor U12534 (N_12534,N_12444,N_12030);
and U12535 (N_12535,N_11944,N_12247);
xnor U12536 (N_12536,N_12061,N_11956);
nor U12537 (N_12537,N_12214,N_12228);
and U12538 (N_12538,N_12303,N_12415);
nor U12539 (N_12539,N_12259,N_12289);
and U12540 (N_12540,N_11967,N_11983);
xor U12541 (N_12541,N_12294,N_12157);
and U12542 (N_12542,N_11959,N_12243);
nor U12543 (N_12543,N_12047,N_12336);
nand U12544 (N_12544,N_12442,N_11985);
or U12545 (N_12545,N_11936,N_12393);
nor U12546 (N_12546,N_12299,N_12472);
and U12547 (N_12547,N_12440,N_12025);
and U12548 (N_12548,N_12024,N_12137);
nand U12549 (N_12549,N_12232,N_12463);
nor U12550 (N_12550,N_12231,N_12417);
nor U12551 (N_12551,N_12104,N_12396);
nand U12552 (N_12552,N_12124,N_12324);
nor U12553 (N_12553,N_11892,N_12182);
or U12554 (N_12554,N_11934,N_12136);
xnor U12555 (N_12555,N_12212,N_12036);
nand U12556 (N_12556,N_12326,N_12392);
nand U12557 (N_12557,N_12009,N_12049);
nand U12558 (N_12558,N_12403,N_11988);
nand U12559 (N_12559,N_12443,N_12023);
xnor U12560 (N_12560,N_11970,N_11881);
nand U12561 (N_12561,N_12387,N_11882);
or U12562 (N_12562,N_12075,N_12322);
and U12563 (N_12563,N_12125,N_12433);
nor U12564 (N_12564,N_12007,N_12162);
nand U12565 (N_12565,N_12370,N_12082);
xor U12566 (N_12566,N_12421,N_11912);
nor U12567 (N_12567,N_12430,N_12188);
or U12568 (N_12568,N_12152,N_12488);
or U12569 (N_12569,N_11980,N_11884);
nand U12570 (N_12570,N_12071,N_12161);
xor U12571 (N_12571,N_12077,N_12215);
nand U12572 (N_12572,N_12462,N_12209);
nor U12573 (N_12573,N_12445,N_11914);
or U12574 (N_12574,N_12422,N_12016);
xnor U12575 (N_12575,N_12290,N_11926);
and U12576 (N_12576,N_12103,N_12250);
xnor U12577 (N_12577,N_12166,N_11994);
and U12578 (N_12578,N_12495,N_12134);
nor U12579 (N_12579,N_12210,N_12343);
and U12580 (N_12580,N_11984,N_12144);
and U12581 (N_12581,N_12223,N_12383);
xnor U12582 (N_12582,N_12480,N_12240);
nand U12583 (N_12583,N_12473,N_12107);
xor U12584 (N_12584,N_12055,N_12203);
and U12585 (N_12585,N_12112,N_12269);
nand U12586 (N_12586,N_12318,N_12168);
nor U12587 (N_12587,N_12174,N_12089);
nand U12588 (N_12588,N_12220,N_12375);
or U12589 (N_12589,N_11922,N_12311);
or U12590 (N_12590,N_11990,N_12260);
and U12591 (N_12591,N_12395,N_12117);
or U12592 (N_12592,N_12281,N_11947);
nand U12593 (N_12593,N_12352,N_12096);
nand U12594 (N_12594,N_11918,N_12331);
or U12595 (N_12595,N_12006,N_12486);
nor U12596 (N_12596,N_12287,N_12476);
nor U12597 (N_12597,N_12001,N_12187);
and U12598 (N_12598,N_12426,N_12262);
or U12599 (N_12599,N_12019,N_12327);
or U12600 (N_12600,N_11886,N_12159);
xnor U12601 (N_12601,N_12199,N_12005);
xnor U12602 (N_12602,N_12147,N_11974);
xnor U12603 (N_12603,N_12349,N_12320);
or U12604 (N_12604,N_12306,N_12227);
and U12605 (N_12605,N_12377,N_11898);
xnor U12606 (N_12606,N_12236,N_12074);
and U12607 (N_12607,N_12492,N_12423);
nor U12608 (N_12608,N_12164,N_12366);
and U12609 (N_12609,N_12255,N_12062);
nor U12610 (N_12610,N_12487,N_12438);
nor U12611 (N_12611,N_12499,N_12135);
nand U12612 (N_12612,N_12084,N_11941);
or U12613 (N_12613,N_11908,N_12113);
nor U12614 (N_12614,N_12371,N_12453);
nor U12615 (N_12615,N_12000,N_12334);
or U12616 (N_12616,N_12280,N_11923);
nor U12617 (N_12617,N_12278,N_12095);
xnor U12618 (N_12618,N_12043,N_12046);
nor U12619 (N_12619,N_12276,N_12356);
xor U12620 (N_12620,N_11930,N_12221);
or U12621 (N_12621,N_11925,N_12233);
and U12622 (N_12622,N_11999,N_12106);
nand U12623 (N_12623,N_11966,N_12466);
xor U12624 (N_12624,N_12382,N_12246);
nor U12625 (N_12625,N_12183,N_12319);
nor U12626 (N_12626,N_12235,N_12003);
xor U12627 (N_12627,N_11876,N_12268);
or U12628 (N_12628,N_12339,N_12059);
nand U12629 (N_12629,N_12363,N_12470);
and U12630 (N_12630,N_11998,N_12155);
xnor U12631 (N_12631,N_12175,N_12156);
xnor U12632 (N_12632,N_11919,N_11991);
xor U12633 (N_12633,N_12257,N_12066);
and U12634 (N_12634,N_12039,N_12158);
xor U12635 (N_12635,N_11975,N_12398);
nor U12636 (N_12636,N_12018,N_12305);
nor U12637 (N_12637,N_12427,N_12347);
nand U12638 (N_12638,N_12411,N_11909);
nand U12639 (N_12639,N_12146,N_12279);
and U12640 (N_12640,N_12298,N_12404);
and U12641 (N_12641,N_12297,N_12419);
nand U12642 (N_12642,N_12110,N_11937);
and U12643 (N_12643,N_11950,N_12154);
or U12644 (N_12644,N_12132,N_12361);
and U12645 (N_12645,N_12072,N_12459);
nand U12646 (N_12646,N_12116,N_12458);
nor U12647 (N_12647,N_12332,N_12340);
or U12648 (N_12648,N_11900,N_11893);
nor U12649 (N_12649,N_12364,N_12170);
or U12650 (N_12650,N_12378,N_12042);
nor U12651 (N_12651,N_12081,N_12198);
nor U12652 (N_12652,N_12252,N_12050);
nor U12653 (N_12653,N_11964,N_12338);
nor U12654 (N_12654,N_12054,N_12441);
xor U12655 (N_12655,N_12217,N_12384);
xnor U12656 (N_12656,N_11949,N_11889);
nor U12657 (N_12657,N_12078,N_12429);
or U12658 (N_12658,N_12315,N_12031);
and U12659 (N_12659,N_12165,N_12224);
nor U12660 (N_12660,N_12004,N_12434);
nand U12661 (N_12661,N_12330,N_12301);
nand U12662 (N_12662,N_12035,N_12368);
or U12663 (N_12663,N_12380,N_12069);
and U12664 (N_12664,N_12150,N_12148);
nand U12665 (N_12665,N_12076,N_11891);
nand U12666 (N_12666,N_12131,N_12376);
nand U12667 (N_12667,N_12407,N_12090);
nor U12668 (N_12668,N_11961,N_11972);
nor U12669 (N_12669,N_12328,N_12449);
or U12670 (N_12670,N_11973,N_12133);
or U12671 (N_12671,N_11938,N_12254);
nor U12672 (N_12672,N_12416,N_12012);
nor U12673 (N_12673,N_12479,N_12193);
nor U12674 (N_12674,N_12105,N_12184);
xor U12675 (N_12675,N_12093,N_11945);
nor U12676 (N_12676,N_12114,N_12027);
xnor U12677 (N_12677,N_11878,N_12481);
or U12678 (N_12678,N_12013,N_11903);
nand U12679 (N_12679,N_12310,N_12357);
or U12680 (N_12680,N_12283,N_12098);
nand U12681 (N_12681,N_12355,N_12028);
nand U12682 (N_12682,N_12413,N_12037);
xor U12683 (N_12683,N_12354,N_12056);
or U12684 (N_12684,N_12094,N_12484);
nand U12685 (N_12685,N_12275,N_11981);
nand U12686 (N_12686,N_12362,N_11954);
xnor U12687 (N_12687,N_12360,N_12109);
or U12688 (N_12688,N_12021,N_12141);
xor U12689 (N_12689,N_12222,N_12258);
nand U12690 (N_12690,N_12389,N_11978);
and U12691 (N_12691,N_12173,N_11955);
xor U12692 (N_12692,N_12225,N_12044);
xnor U12693 (N_12693,N_12153,N_12065);
nor U12694 (N_12694,N_12314,N_12204);
xnor U12695 (N_12695,N_12261,N_12351);
and U12696 (N_12696,N_11880,N_12014);
and U12697 (N_12697,N_12333,N_12026);
xor U12698 (N_12698,N_11913,N_12265);
nor U12699 (N_12699,N_12118,N_11943);
nor U12700 (N_12700,N_11916,N_12249);
or U12701 (N_12701,N_11904,N_12253);
nand U12702 (N_12702,N_12211,N_12431);
and U12703 (N_12703,N_12277,N_11935);
or U12704 (N_12704,N_11940,N_12379);
or U12705 (N_12705,N_12149,N_12060);
and U12706 (N_12706,N_12201,N_12358);
nand U12707 (N_12707,N_12475,N_12451);
nand U12708 (N_12708,N_12083,N_12034);
or U12709 (N_12709,N_12127,N_12091);
and U12710 (N_12710,N_12196,N_12238);
nor U12711 (N_12711,N_11939,N_11915);
or U12712 (N_12712,N_12372,N_12032);
xor U12713 (N_12713,N_12386,N_12267);
and U12714 (N_12714,N_12057,N_11977);
xnor U12715 (N_12715,N_12239,N_12367);
nor U12716 (N_12716,N_12181,N_12424);
and U12717 (N_12717,N_12229,N_12452);
nand U12718 (N_12718,N_12111,N_12100);
xor U12719 (N_12719,N_12040,N_12300);
or U12720 (N_12720,N_12350,N_11906);
nand U12721 (N_12721,N_11979,N_12329);
and U12722 (N_12722,N_12213,N_12151);
or U12723 (N_12723,N_11969,N_12369);
xnor U12724 (N_12724,N_12293,N_11976);
nor U12725 (N_12725,N_12450,N_12230);
nor U12726 (N_12726,N_12010,N_12045);
nor U12727 (N_12727,N_12169,N_12033);
and U12728 (N_12728,N_12291,N_12038);
xnor U12729 (N_12729,N_12058,N_12418);
xnor U12730 (N_12730,N_12070,N_12085);
and U12731 (N_12731,N_12359,N_12385);
nand U12732 (N_12732,N_11987,N_12064);
xor U12733 (N_12733,N_11952,N_12272);
nand U12734 (N_12734,N_12471,N_12405);
nand U12735 (N_12735,N_11933,N_12200);
nand U12736 (N_12736,N_12335,N_12456);
nand U12737 (N_12737,N_12296,N_12087);
or U12738 (N_12738,N_12263,N_12478);
nand U12739 (N_12739,N_12053,N_12142);
nand U12740 (N_12740,N_12353,N_11942);
nand U12741 (N_12741,N_12316,N_12365);
nand U12742 (N_12742,N_12176,N_11948);
nand U12743 (N_12743,N_12115,N_12295);
nor U12744 (N_12744,N_12145,N_12079);
or U12745 (N_12745,N_12312,N_11962);
xnor U12746 (N_12746,N_12122,N_11993);
or U12747 (N_12747,N_12489,N_12432);
and U12748 (N_12748,N_12344,N_12381);
xnor U12749 (N_12749,N_11953,N_12226);
nor U12750 (N_12750,N_12206,N_12202);
xor U12751 (N_12751,N_11877,N_12041);
and U12752 (N_12752,N_12439,N_12497);
or U12753 (N_12753,N_11927,N_12015);
xor U12754 (N_12754,N_12498,N_12271);
nor U12755 (N_12755,N_12313,N_11907);
and U12756 (N_12756,N_11989,N_12128);
nor U12757 (N_12757,N_12446,N_11995);
nor U12758 (N_12758,N_12388,N_12292);
xnor U12759 (N_12759,N_12244,N_11968);
nand U12760 (N_12760,N_12067,N_12304);
or U12761 (N_12761,N_12189,N_12469);
or U12762 (N_12762,N_12408,N_12342);
nor U12763 (N_12763,N_12092,N_12436);
nor U12764 (N_12764,N_12179,N_11895);
nand U12765 (N_12765,N_12108,N_12017);
nand U12766 (N_12766,N_12302,N_12390);
and U12767 (N_12767,N_12406,N_12493);
xnor U12768 (N_12768,N_12307,N_12218);
xor U12769 (N_12769,N_12163,N_11992);
or U12770 (N_12770,N_12256,N_12101);
and U12771 (N_12771,N_12485,N_12126);
and U12772 (N_12772,N_12123,N_12477);
or U12773 (N_12773,N_11965,N_12282);
or U12774 (N_12774,N_12346,N_12102);
nand U12775 (N_12775,N_11971,N_11960);
xnor U12776 (N_12776,N_12234,N_11986);
or U12777 (N_12777,N_12251,N_12099);
and U12778 (N_12778,N_12186,N_12461);
or U12779 (N_12779,N_12345,N_12245);
xor U12780 (N_12780,N_12048,N_11885);
or U12781 (N_12781,N_12399,N_12190);
and U12782 (N_12782,N_11911,N_12160);
nand U12783 (N_12783,N_12448,N_12120);
and U12784 (N_12784,N_12237,N_11879);
nand U12785 (N_12785,N_11920,N_12248);
xor U12786 (N_12786,N_12273,N_11875);
nor U12787 (N_12787,N_12321,N_12412);
and U12788 (N_12788,N_11890,N_12483);
nand U12789 (N_12789,N_12468,N_11996);
nor U12790 (N_12790,N_12491,N_12394);
and U12791 (N_12791,N_12139,N_11963);
nor U12792 (N_12792,N_12401,N_11917);
nand U12793 (N_12793,N_12460,N_12455);
nand U12794 (N_12794,N_12397,N_12011);
and U12795 (N_12795,N_12447,N_12097);
nor U12796 (N_12796,N_12373,N_11888);
and U12797 (N_12797,N_11931,N_12008);
nand U12798 (N_12798,N_12428,N_12465);
nand U12799 (N_12799,N_12080,N_12052);
nor U12800 (N_12800,N_11899,N_11982);
nor U12801 (N_12801,N_12172,N_11905);
xor U12802 (N_12802,N_12402,N_12130);
nor U12803 (N_12803,N_12194,N_12167);
and U12804 (N_12804,N_12171,N_12464);
nor U12805 (N_12805,N_12490,N_12197);
and U12806 (N_12806,N_12414,N_12264);
xor U12807 (N_12807,N_12323,N_12022);
and U12808 (N_12808,N_12177,N_11928);
xnor U12809 (N_12809,N_11932,N_12341);
nor U12810 (N_12810,N_12348,N_12143);
and U12811 (N_12811,N_12192,N_12178);
and U12812 (N_12812,N_12284,N_12445);
or U12813 (N_12813,N_11928,N_12289);
xnor U12814 (N_12814,N_12112,N_12154);
xnor U12815 (N_12815,N_12205,N_11948);
nand U12816 (N_12816,N_11893,N_12154);
nor U12817 (N_12817,N_11883,N_12482);
nand U12818 (N_12818,N_12264,N_12213);
nor U12819 (N_12819,N_11875,N_12334);
xnor U12820 (N_12820,N_12315,N_11946);
and U12821 (N_12821,N_12068,N_12120);
xnor U12822 (N_12822,N_12143,N_12284);
nand U12823 (N_12823,N_12228,N_12119);
and U12824 (N_12824,N_12034,N_12256);
nor U12825 (N_12825,N_12369,N_12153);
nor U12826 (N_12826,N_12037,N_12252);
or U12827 (N_12827,N_12419,N_12341);
nor U12828 (N_12828,N_11900,N_12018);
nand U12829 (N_12829,N_12462,N_11983);
and U12830 (N_12830,N_12307,N_12170);
and U12831 (N_12831,N_11991,N_11968);
and U12832 (N_12832,N_11894,N_12043);
xnor U12833 (N_12833,N_12027,N_12107);
nor U12834 (N_12834,N_12348,N_12053);
xnor U12835 (N_12835,N_12324,N_12335);
xnor U12836 (N_12836,N_11912,N_12357);
and U12837 (N_12837,N_12179,N_11986);
and U12838 (N_12838,N_12432,N_12208);
or U12839 (N_12839,N_12338,N_11900);
xnor U12840 (N_12840,N_12299,N_12204);
or U12841 (N_12841,N_12313,N_12276);
and U12842 (N_12842,N_12432,N_11970);
or U12843 (N_12843,N_12447,N_12353);
nand U12844 (N_12844,N_12059,N_11899);
nor U12845 (N_12845,N_12209,N_12436);
nor U12846 (N_12846,N_12360,N_12156);
xnor U12847 (N_12847,N_11876,N_12486);
or U12848 (N_12848,N_11971,N_12382);
or U12849 (N_12849,N_12391,N_11966);
and U12850 (N_12850,N_12365,N_12143);
or U12851 (N_12851,N_12392,N_12113);
nand U12852 (N_12852,N_12192,N_12006);
nand U12853 (N_12853,N_11993,N_12163);
nand U12854 (N_12854,N_12282,N_11937);
xnor U12855 (N_12855,N_12068,N_12252);
or U12856 (N_12856,N_12051,N_12282);
or U12857 (N_12857,N_12432,N_12251);
nor U12858 (N_12858,N_12093,N_12013);
or U12859 (N_12859,N_12278,N_12363);
or U12860 (N_12860,N_12347,N_11946);
nand U12861 (N_12861,N_12200,N_11923);
xor U12862 (N_12862,N_12023,N_12215);
nor U12863 (N_12863,N_12148,N_12081);
and U12864 (N_12864,N_12065,N_12134);
xnor U12865 (N_12865,N_12281,N_12472);
xnor U12866 (N_12866,N_12107,N_11963);
nor U12867 (N_12867,N_12052,N_12392);
or U12868 (N_12868,N_11927,N_11993);
xnor U12869 (N_12869,N_12065,N_12315);
nand U12870 (N_12870,N_11929,N_12011);
nor U12871 (N_12871,N_12416,N_12379);
xor U12872 (N_12872,N_12032,N_11976);
nor U12873 (N_12873,N_12401,N_12003);
or U12874 (N_12874,N_12069,N_12473);
xor U12875 (N_12875,N_11909,N_12116);
nand U12876 (N_12876,N_11976,N_11879);
nor U12877 (N_12877,N_12427,N_12277);
and U12878 (N_12878,N_11886,N_12414);
xnor U12879 (N_12879,N_12140,N_12247);
nor U12880 (N_12880,N_11907,N_12419);
xor U12881 (N_12881,N_12017,N_12164);
or U12882 (N_12882,N_12430,N_12183);
and U12883 (N_12883,N_11909,N_12210);
xnor U12884 (N_12884,N_12151,N_12251);
or U12885 (N_12885,N_12350,N_12386);
or U12886 (N_12886,N_12058,N_11922);
and U12887 (N_12887,N_12440,N_12388);
nor U12888 (N_12888,N_11918,N_12156);
or U12889 (N_12889,N_11933,N_12444);
xnor U12890 (N_12890,N_12201,N_11892);
or U12891 (N_12891,N_12430,N_12308);
or U12892 (N_12892,N_12302,N_11954);
xnor U12893 (N_12893,N_12466,N_12103);
xor U12894 (N_12894,N_11936,N_12395);
or U12895 (N_12895,N_12040,N_12288);
or U12896 (N_12896,N_12018,N_11988);
or U12897 (N_12897,N_11909,N_11879);
nor U12898 (N_12898,N_12103,N_12485);
and U12899 (N_12899,N_12288,N_12339);
xor U12900 (N_12900,N_12456,N_12312);
nand U12901 (N_12901,N_12065,N_12458);
nand U12902 (N_12902,N_11967,N_11999);
xor U12903 (N_12903,N_11901,N_12248);
xor U12904 (N_12904,N_12247,N_11910);
nand U12905 (N_12905,N_11885,N_12204);
nand U12906 (N_12906,N_12022,N_12236);
and U12907 (N_12907,N_12191,N_11956);
or U12908 (N_12908,N_12362,N_12404);
and U12909 (N_12909,N_12474,N_11878);
or U12910 (N_12910,N_12134,N_12338);
xor U12911 (N_12911,N_12010,N_12247);
or U12912 (N_12912,N_12038,N_12481);
nand U12913 (N_12913,N_11972,N_12472);
or U12914 (N_12914,N_12233,N_12061);
or U12915 (N_12915,N_12334,N_12391);
xor U12916 (N_12916,N_11890,N_11896);
xor U12917 (N_12917,N_11954,N_12152);
xor U12918 (N_12918,N_12366,N_11997);
xnor U12919 (N_12919,N_12157,N_12326);
nand U12920 (N_12920,N_12082,N_12498);
nand U12921 (N_12921,N_12297,N_11876);
nor U12922 (N_12922,N_12209,N_12229);
nand U12923 (N_12923,N_12222,N_12126);
nor U12924 (N_12924,N_12269,N_11949);
and U12925 (N_12925,N_12162,N_12419);
xor U12926 (N_12926,N_12064,N_12254);
nand U12927 (N_12927,N_12155,N_12400);
or U12928 (N_12928,N_12203,N_12140);
xnor U12929 (N_12929,N_12140,N_12102);
xor U12930 (N_12930,N_12243,N_12261);
and U12931 (N_12931,N_12367,N_12105);
or U12932 (N_12932,N_12049,N_12003);
and U12933 (N_12933,N_12060,N_11882);
and U12934 (N_12934,N_12153,N_12496);
nor U12935 (N_12935,N_12441,N_12181);
xor U12936 (N_12936,N_12410,N_11919);
nand U12937 (N_12937,N_11885,N_11977);
nand U12938 (N_12938,N_12014,N_12060);
or U12939 (N_12939,N_12460,N_12158);
and U12940 (N_12940,N_12036,N_12088);
and U12941 (N_12941,N_12304,N_12241);
or U12942 (N_12942,N_12462,N_12441);
or U12943 (N_12943,N_12152,N_12270);
nand U12944 (N_12944,N_12347,N_12159);
or U12945 (N_12945,N_12131,N_12386);
nor U12946 (N_12946,N_12091,N_12276);
nand U12947 (N_12947,N_11993,N_12062);
and U12948 (N_12948,N_12327,N_12081);
or U12949 (N_12949,N_12068,N_12034);
xor U12950 (N_12950,N_12195,N_12337);
nor U12951 (N_12951,N_12405,N_12438);
and U12952 (N_12952,N_12181,N_12104);
nor U12953 (N_12953,N_12256,N_11998);
nand U12954 (N_12954,N_12104,N_12463);
nor U12955 (N_12955,N_12189,N_12161);
nor U12956 (N_12956,N_11963,N_12219);
nor U12957 (N_12957,N_12472,N_12054);
or U12958 (N_12958,N_12312,N_12305);
nand U12959 (N_12959,N_11950,N_12392);
nand U12960 (N_12960,N_11936,N_12268);
xor U12961 (N_12961,N_12228,N_12288);
or U12962 (N_12962,N_11984,N_12008);
nand U12963 (N_12963,N_12355,N_11990);
xor U12964 (N_12964,N_11900,N_11919);
xor U12965 (N_12965,N_12165,N_12009);
nor U12966 (N_12966,N_12423,N_12123);
xnor U12967 (N_12967,N_12060,N_12391);
and U12968 (N_12968,N_12305,N_12042);
and U12969 (N_12969,N_12332,N_12182);
nand U12970 (N_12970,N_12315,N_12400);
and U12971 (N_12971,N_12160,N_12479);
and U12972 (N_12972,N_11985,N_11947);
nor U12973 (N_12973,N_12036,N_12446);
nor U12974 (N_12974,N_12044,N_12121);
or U12975 (N_12975,N_11878,N_11982);
and U12976 (N_12976,N_12382,N_12237);
xnor U12977 (N_12977,N_12484,N_12325);
or U12978 (N_12978,N_11982,N_12308);
and U12979 (N_12979,N_12476,N_12197);
nand U12980 (N_12980,N_12020,N_12468);
nor U12981 (N_12981,N_11893,N_12470);
and U12982 (N_12982,N_12282,N_11973);
xor U12983 (N_12983,N_12157,N_12447);
and U12984 (N_12984,N_12188,N_11996);
or U12985 (N_12985,N_12249,N_12266);
nor U12986 (N_12986,N_12357,N_12322);
or U12987 (N_12987,N_11898,N_12293);
or U12988 (N_12988,N_12442,N_12486);
nor U12989 (N_12989,N_12050,N_12017);
or U12990 (N_12990,N_12250,N_12453);
and U12991 (N_12991,N_12071,N_12465);
xor U12992 (N_12992,N_12038,N_11925);
nor U12993 (N_12993,N_12056,N_12457);
and U12994 (N_12994,N_11936,N_12214);
nand U12995 (N_12995,N_12280,N_12100);
nand U12996 (N_12996,N_12039,N_12272);
nor U12997 (N_12997,N_11879,N_12493);
xnor U12998 (N_12998,N_12107,N_12311);
xnor U12999 (N_12999,N_12140,N_12421);
nor U13000 (N_13000,N_12021,N_12423);
nor U13001 (N_13001,N_12168,N_12288);
nor U13002 (N_13002,N_12096,N_12274);
xnor U13003 (N_13003,N_12431,N_12268);
nand U13004 (N_13004,N_12483,N_12347);
xnor U13005 (N_13005,N_12252,N_12243);
nand U13006 (N_13006,N_11965,N_11944);
and U13007 (N_13007,N_12410,N_12237);
or U13008 (N_13008,N_12332,N_12296);
nand U13009 (N_13009,N_12368,N_12133);
nand U13010 (N_13010,N_11881,N_12301);
nor U13011 (N_13011,N_12485,N_12397);
and U13012 (N_13012,N_12084,N_12030);
nor U13013 (N_13013,N_12120,N_12000);
or U13014 (N_13014,N_12354,N_12165);
nor U13015 (N_13015,N_12069,N_12063);
or U13016 (N_13016,N_12354,N_12374);
nor U13017 (N_13017,N_11884,N_11906);
xor U13018 (N_13018,N_12032,N_12370);
nand U13019 (N_13019,N_12490,N_12475);
xnor U13020 (N_13020,N_12132,N_12477);
xor U13021 (N_13021,N_12207,N_12274);
nor U13022 (N_13022,N_12243,N_12027);
nor U13023 (N_13023,N_12366,N_11900);
and U13024 (N_13024,N_12173,N_12203);
and U13025 (N_13025,N_11980,N_12059);
xor U13026 (N_13026,N_12381,N_11970);
and U13027 (N_13027,N_12092,N_12051);
nand U13028 (N_13028,N_12456,N_12285);
xor U13029 (N_13029,N_12169,N_12093);
and U13030 (N_13030,N_11894,N_12142);
and U13031 (N_13031,N_12086,N_12478);
xnor U13032 (N_13032,N_11928,N_11947);
nand U13033 (N_13033,N_12248,N_12007);
nor U13034 (N_13034,N_12245,N_12321);
nor U13035 (N_13035,N_12228,N_12246);
nand U13036 (N_13036,N_12412,N_11905);
and U13037 (N_13037,N_11887,N_12156);
nor U13038 (N_13038,N_12083,N_12438);
and U13039 (N_13039,N_11986,N_12358);
and U13040 (N_13040,N_12258,N_12202);
or U13041 (N_13041,N_12300,N_12181);
nand U13042 (N_13042,N_12012,N_12063);
or U13043 (N_13043,N_12451,N_12357);
nor U13044 (N_13044,N_11982,N_12284);
xnor U13045 (N_13045,N_11949,N_12256);
nor U13046 (N_13046,N_11878,N_11934);
nand U13047 (N_13047,N_12380,N_12113);
nand U13048 (N_13048,N_12141,N_12232);
or U13049 (N_13049,N_11943,N_12023);
or U13050 (N_13050,N_12188,N_11898);
nor U13051 (N_13051,N_12333,N_12464);
xor U13052 (N_13052,N_11905,N_11885);
nand U13053 (N_13053,N_11919,N_12428);
nor U13054 (N_13054,N_12439,N_12317);
or U13055 (N_13055,N_12073,N_12046);
and U13056 (N_13056,N_12435,N_12318);
xor U13057 (N_13057,N_12416,N_12403);
nor U13058 (N_13058,N_12468,N_12436);
xnor U13059 (N_13059,N_12472,N_11983);
nand U13060 (N_13060,N_12205,N_12109);
or U13061 (N_13061,N_11963,N_12003);
and U13062 (N_13062,N_12216,N_12204);
nand U13063 (N_13063,N_12179,N_12151);
and U13064 (N_13064,N_11978,N_12027);
and U13065 (N_13065,N_11911,N_11912);
and U13066 (N_13066,N_11971,N_12052);
and U13067 (N_13067,N_12452,N_11933);
nand U13068 (N_13068,N_11892,N_11994);
and U13069 (N_13069,N_11922,N_12002);
nor U13070 (N_13070,N_12264,N_12334);
and U13071 (N_13071,N_12223,N_12111);
xor U13072 (N_13072,N_12498,N_12085);
nand U13073 (N_13073,N_12345,N_11904);
and U13074 (N_13074,N_12022,N_12424);
nor U13075 (N_13075,N_12189,N_12128);
nor U13076 (N_13076,N_12426,N_12222);
or U13077 (N_13077,N_11965,N_12245);
and U13078 (N_13078,N_12061,N_12041);
and U13079 (N_13079,N_12425,N_12075);
and U13080 (N_13080,N_12245,N_12415);
nor U13081 (N_13081,N_11911,N_12209);
xnor U13082 (N_13082,N_12417,N_12059);
nand U13083 (N_13083,N_12216,N_11974);
nand U13084 (N_13084,N_12383,N_12065);
or U13085 (N_13085,N_12228,N_12083);
or U13086 (N_13086,N_11991,N_12479);
and U13087 (N_13087,N_12378,N_12428);
xnor U13088 (N_13088,N_11884,N_12413);
or U13089 (N_13089,N_12344,N_11890);
and U13090 (N_13090,N_12489,N_12289);
nor U13091 (N_13091,N_12242,N_12480);
and U13092 (N_13092,N_12421,N_12280);
nor U13093 (N_13093,N_12124,N_12284);
or U13094 (N_13094,N_12437,N_12395);
nand U13095 (N_13095,N_12490,N_12218);
or U13096 (N_13096,N_12131,N_12310);
nor U13097 (N_13097,N_12098,N_12206);
xor U13098 (N_13098,N_12448,N_12481);
and U13099 (N_13099,N_12486,N_12386);
xor U13100 (N_13100,N_12268,N_12403);
nor U13101 (N_13101,N_12132,N_12110);
or U13102 (N_13102,N_12285,N_12442);
nand U13103 (N_13103,N_11981,N_12206);
or U13104 (N_13104,N_12319,N_12069);
and U13105 (N_13105,N_12340,N_12344);
xnor U13106 (N_13106,N_12395,N_11966);
nor U13107 (N_13107,N_12420,N_11932);
and U13108 (N_13108,N_12105,N_12422);
and U13109 (N_13109,N_12190,N_12174);
xor U13110 (N_13110,N_12176,N_12374);
or U13111 (N_13111,N_12432,N_12156);
xor U13112 (N_13112,N_11963,N_12465);
nand U13113 (N_13113,N_12350,N_12365);
or U13114 (N_13114,N_12318,N_12220);
nor U13115 (N_13115,N_12360,N_12170);
and U13116 (N_13116,N_11958,N_12486);
xnor U13117 (N_13117,N_12208,N_12093);
xor U13118 (N_13118,N_11927,N_12485);
xor U13119 (N_13119,N_11878,N_12003);
nand U13120 (N_13120,N_11978,N_11877);
or U13121 (N_13121,N_11999,N_12020);
or U13122 (N_13122,N_12100,N_12327);
xor U13123 (N_13123,N_12492,N_11953);
nand U13124 (N_13124,N_12298,N_12398);
and U13125 (N_13125,N_12549,N_12718);
xnor U13126 (N_13126,N_12777,N_12710);
and U13127 (N_13127,N_12552,N_12558);
and U13128 (N_13128,N_12940,N_12507);
or U13129 (N_13129,N_13007,N_12951);
nor U13130 (N_13130,N_13048,N_13121);
or U13131 (N_13131,N_12743,N_13092);
and U13132 (N_13132,N_12663,N_12837);
nor U13133 (N_13133,N_12791,N_12541);
or U13134 (N_13134,N_13119,N_12809);
or U13135 (N_13135,N_12853,N_13067);
or U13136 (N_13136,N_12588,N_13046);
xor U13137 (N_13137,N_13036,N_12828);
and U13138 (N_13138,N_12999,N_13052);
nand U13139 (N_13139,N_13094,N_13068);
nand U13140 (N_13140,N_12759,N_12754);
nor U13141 (N_13141,N_12536,N_12736);
nor U13142 (N_13142,N_12638,N_12907);
xnor U13143 (N_13143,N_12964,N_12734);
and U13144 (N_13144,N_13047,N_12904);
and U13145 (N_13145,N_12591,N_12617);
or U13146 (N_13146,N_13101,N_12740);
and U13147 (N_13147,N_12953,N_12962);
nor U13148 (N_13148,N_12513,N_12739);
nor U13149 (N_13149,N_12988,N_12858);
nor U13150 (N_13150,N_12755,N_12578);
nor U13151 (N_13151,N_12772,N_12646);
xnor U13152 (N_13152,N_12846,N_13014);
xnor U13153 (N_13153,N_13085,N_12579);
nand U13154 (N_13154,N_12587,N_12593);
xor U13155 (N_13155,N_13102,N_12997);
or U13156 (N_13156,N_12527,N_12938);
and U13157 (N_13157,N_12872,N_12935);
nor U13158 (N_13158,N_12672,N_12876);
nand U13159 (N_13159,N_13008,N_12529);
nor U13160 (N_13160,N_12577,N_13069);
nand U13161 (N_13161,N_12655,N_12670);
nand U13162 (N_13162,N_12891,N_12781);
nand U13163 (N_13163,N_12598,N_12715);
and U13164 (N_13164,N_12893,N_12773);
xor U13165 (N_13165,N_12787,N_12647);
nand U13166 (N_13166,N_13090,N_12628);
and U13167 (N_13167,N_12918,N_12512);
nand U13168 (N_13168,N_12794,N_13064);
xnor U13169 (N_13169,N_12599,N_12697);
nand U13170 (N_13170,N_13003,N_12738);
nor U13171 (N_13171,N_13105,N_12745);
or U13172 (N_13172,N_12835,N_12987);
nor U13173 (N_13173,N_12609,N_12685);
or U13174 (N_13174,N_12566,N_12774);
xor U13175 (N_13175,N_12836,N_13022);
nor U13176 (N_13176,N_12542,N_12582);
or U13177 (N_13177,N_13072,N_12568);
or U13178 (N_13178,N_12871,N_12636);
or U13179 (N_13179,N_12623,N_12900);
or U13180 (N_13180,N_12922,N_12669);
xnor U13181 (N_13181,N_12981,N_12839);
nand U13182 (N_13182,N_13021,N_12695);
and U13183 (N_13183,N_12892,N_12696);
xor U13184 (N_13184,N_12852,N_13099);
and U13185 (N_13185,N_12522,N_13097);
or U13186 (N_13186,N_12996,N_12866);
nand U13187 (N_13187,N_12899,N_13096);
nand U13188 (N_13188,N_12789,N_12925);
nand U13189 (N_13189,N_12505,N_12965);
nand U13190 (N_13190,N_12750,N_12571);
and U13191 (N_13191,N_12650,N_12915);
xnor U13192 (N_13192,N_12929,N_12676);
nor U13193 (N_13193,N_12592,N_12909);
and U13194 (N_13194,N_12887,N_12714);
nand U13195 (N_13195,N_12500,N_12863);
nand U13196 (N_13196,N_12680,N_12991);
nor U13197 (N_13197,N_12882,N_12573);
nor U13198 (N_13198,N_12844,N_12562);
nor U13199 (N_13199,N_12632,N_12749);
or U13200 (N_13200,N_12662,N_12911);
nor U13201 (N_13201,N_12805,N_12679);
nor U13202 (N_13202,N_12614,N_12833);
or U13203 (N_13203,N_12842,N_12501);
xor U13204 (N_13204,N_12825,N_12810);
nor U13205 (N_13205,N_13104,N_12945);
nand U13206 (N_13206,N_12531,N_12888);
nor U13207 (N_13207,N_12544,N_12982);
nand U13208 (N_13208,N_12684,N_13054);
nand U13209 (N_13209,N_12741,N_12709);
or U13210 (N_13210,N_12631,N_12782);
xnor U13211 (N_13211,N_12534,N_12503);
xnor U13212 (N_13212,N_12790,N_13044);
nand U13213 (N_13213,N_12776,N_13088);
nor U13214 (N_13214,N_12744,N_13042);
nand U13215 (N_13215,N_12622,N_12801);
xnor U13216 (N_13216,N_12737,N_12916);
nand U13217 (N_13217,N_12873,N_12702);
xnor U13218 (N_13218,N_12509,N_12731);
nor U13219 (N_13219,N_12701,N_12808);
nand U13220 (N_13220,N_12619,N_12765);
nand U13221 (N_13221,N_12616,N_12796);
xor U13222 (N_13222,N_12517,N_12937);
xor U13223 (N_13223,N_12797,N_12611);
nor U13224 (N_13224,N_12926,N_12747);
or U13225 (N_13225,N_12860,N_12589);
and U13226 (N_13226,N_12594,N_12763);
nand U13227 (N_13227,N_13040,N_12526);
or U13228 (N_13228,N_13106,N_12989);
nand U13229 (N_13229,N_12625,N_12969);
or U13230 (N_13230,N_12978,N_12976);
or U13231 (N_13231,N_12923,N_12800);
nor U13232 (N_13232,N_12713,N_12519);
or U13233 (N_13233,N_12766,N_12977);
and U13234 (N_13234,N_12525,N_12620);
nand U13235 (N_13235,N_12597,N_13058);
or U13236 (N_13236,N_12548,N_13049);
nand U13237 (N_13237,N_12574,N_12950);
nor U13238 (N_13238,N_12653,N_12807);
xor U13239 (N_13239,N_12851,N_13061);
xor U13240 (N_13240,N_12752,N_12683);
nor U13241 (N_13241,N_13029,N_12979);
xnor U13242 (N_13242,N_12716,N_12586);
and U13243 (N_13243,N_12533,N_12931);
xor U13244 (N_13244,N_12581,N_13111);
or U13245 (N_13245,N_12719,N_13118);
or U13246 (N_13246,N_12504,N_12986);
xnor U13247 (N_13247,N_12829,N_13077);
nand U13248 (N_13248,N_12564,N_12726);
nor U13249 (N_13249,N_12648,N_12895);
nor U13250 (N_13250,N_13009,N_12910);
or U13251 (N_13251,N_12799,N_13084);
or U13252 (N_13252,N_12700,N_12643);
xor U13253 (N_13253,N_12818,N_12771);
and U13254 (N_13254,N_12990,N_12847);
and U13255 (N_13255,N_12855,N_12711);
xor U13256 (N_13256,N_12658,N_12613);
xor U13257 (N_13257,N_13082,N_12928);
xor U13258 (N_13258,N_12841,N_12880);
xnor U13259 (N_13259,N_12681,N_12724);
xnor U13260 (N_13260,N_12601,N_12948);
or U13261 (N_13261,N_13083,N_12874);
or U13262 (N_13262,N_13065,N_12814);
and U13263 (N_13263,N_12551,N_12843);
and U13264 (N_13264,N_12823,N_12932);
xnor U13265 (N_13265,N_13030,N_12570);
nand U13266 (N_13266,N_12758,N_12793);
xnor U13267 (N_13267,N_12603,N_12565);
xor U13268 (N_13268,N_12877,N_12727);
and U13269 (N_13269,N_12768,N_12687);
xor U13270 (N_13270,N_12831,N_13098);
nand U13271 (N_13271,N_12621,N_12634);
xnor U13272 (N_13272,N_12971,N_12967);
and U13273 (N_13273,N_13053,N_12933);
or U13274 (N_13274,N_12703,N_12686);
nor U13275 (N_13275,N_12820,N_12612);
or U13276 (N_13276,N_12678,N_12973);
and U13277 (N_13277,N_12816,N_13062);
nor U13278 (N_13278,N_12659,N_12970);
and U13279 (N_13279,N_12756,N_13034);
and U13280 (N_13280,N_12942,N_13113);
and U13281 (N_13281,N_13023,N_12626);
and U13282 (N_13282,N_12567,N_12920);
or U13283 (N_13283,N_12606,N_12633);
or U13284 (N_13284,N_12879,N_12707);
nor U13285 (N_13285,N_12889,N_12682);
nor U13286 (N_13286,N_12532,N_12575);
nand U13287 (N_13287,N_12753,N_12939);
xnor U13288 (N_13288,N_12824,N_12917);
or U13289 (N_13289,N_12886,N_12723);
and U13290 (N_13290,N_12983,N_13031);
nor U13291 (N_13291,N_12733,N_12795);
or U13292 (N_13292,N_12884,N_13073);
nand U13293 (N_13293,N_12821,N_12784);
xor U13294 (N_13294,N_13078,N_12607);
xnor U13295 (N_13295,N_12604,N_12595);
nand U13296 (N_13296,N_12959,N_12518);
nor U13297 (N_13297,N_12720,N_13001);
or U13298 (N_13298,N_12767,N_12732);
xor U13299 (N_13299,N_12864,N_12946);
and U13300 (N_13300,N_13025,N_12660);
and U13301 (N_13301,N_12764,N_12694);
xnor U13302 (N_13302,N_12848,N_13107);
nor U13303 (N_13303,N_12742,N_12778);
xor U13304 (N_13304,N_12610,N_12537);
or U13305 (N_13305,N_12651,N_12735);
xnor U13306 (N_13306,N_12897,N_13024);
or U13307 (N_13307,N_12572,N_12870);
or U13308 (N_13308,N_13081,N_12602);
or U13309 (N_13309,N_12802,N_12652);
nor U13310 (N_13310,N_12803,N_12661);
xnor U13311 (N_13311,N_12941,N_12914);
nand U13312 (N_13312,N_13100,N_12867);
and U13313 (N_13313,N_12665,N_13089);
nor U13314 (N_13314,N_12639,N_13115);
and U13315 (N_13315,N_12538,N_12783);
or U13316 (N_13316,N_12975,N_12806);
nand U13317 (N_13317,N_12554,N_12792);
and U13318 (N_13318,N_12528,N_12540);
and U13319 (N_13319,N_13116,N_12569);
xnor U13320 (N_13320,N_12798,N_13056);
or U13321 (N_13321,N_13050,N_12974);
nand U13322 (N_13322,N_12717,N_12691);
nor U13323 (N_13323,N_12510,N_13028);
xor U13324 (N_13324,N_12520,N_13027);
xnor U13325 (N_13325,N_12675,N_12712);
xnor U13326 (N_13326,N_12952,N_13123);
nor U13327 (N_13327,N_12868,N_12561);
or U13328 (N_13328,N_13016,N_12748);
or U13329 (N_13329,N_13095,N_12644);
nor U13330 (N_13330,N_12690,N_13051);
xor U13331 (N_13331,N_12913,N_13110);
or U13332 (N_13332,N_12698,N_13086);
nand U13333 (N_13333,N_12608,N_13074);
or U13334 (N_13334,N_12629,N_12961);
xor U13335 (N_13335,N_12968,N_12725);
xnor U13336 (N_13336,N_12908,N_12838);
and U13337 (N_13337,N_12530,N_12666);
xor U13338 (N_13338,N_12630,N_13045);
xnor U13339 (N_13339,N_12786,N_12506);
and U13340 (N_13340,N_12822,N_12769);
or U13341 (N_13341,N_12642,N_12692);
nor U13342 (N_13342,N_12555,N_13000);
and U13343 (N_13343,N_13017,N_12854);
nor U13344 (N_13344,N_13079,N_13039);
xnor U13345 (N_13345,N_12780,N_12688);
and U13346 (N_13346,N_12722,N_12963);
xor U13347 (N_13347,N_12779,N_12869);
or U13348 (N_13348,N_12514,N_12905);
or U13349 (N_13349,N_12934,N_12955);
or U13350 (N_13350,N_13109,N_13004);
and U13351 (N_13351,N_13124,N_12956);
or U13352 (N_13352,N_12985,N_12811);
or U13353 (N_13353,N_12834,N_12708);
and U13354 (N_13354,N_13032,N_13002);
nand U13355 (N_13355,N_12775,N_13075);
nand U13356 (N_13356,N_12585,N_12762);
and U13357 (N_13357,N_13071,N_12543);
nor U13358 (N_13358,N_12830,N_12890);
nand U13359 (N_13359,N_12995,N_12645);
xnor U13360 (N_13360,N_13019,N_12556);
or U13361 (N_13361,N_12674,N_12857);
xnor U13362 (N_13362,N_12673,N_13013);
xnor U13363 (N_13363,N_12635,N_13122);
nor U13364 (N_13364,N_13093,N_12521);
xnor U13365 (N_13365,N_12998,N_12550);
nor U13366 (N_13366,N_12580,N_12912);
and U13367 (N_13367,N_12947,N_12760);
and U13368 (N_13368,N_12511,N_13091);
xor U13369 (N_13369,N_12817,N_13012);
nor U13370 (N_13370,N_12859,N_12832);
xnor U13371 (N_13371,N_12804,N_12721);
xor U13372 (N_13372,N_13038,N_12746);
nand U13373 (N_13373,N_12654,N_13018);
and U13374 (N_13374,N_12667,N_12576);
nor U13375 (N_13375,N_12902,N_12557);
or U13376 (N_13376,N_13066,N_12657);
or U13377 (N_13377,N_13063,N_12896);
xor U13378 (N_13378,N_12546,N_12705);
nor U13379 (N_13379,N_12865,N_13103);
nand U13380 (N_13380,N_12980,N_12845);
nand U13381 (N_13381,N_12924,N_13035);
xor U13382 (N_13382,N_12770,N_12689);
and U13383 (N_13383,N_12668,N_12757);
xnor U13384 (N_13384,N_12957,N_13120);
and U13385 (N_13385,N_12584,N_13020);
xnor U13386 (N_13386,N_12883,N_12815);
or U13387 (N_13387,N_12788,N_12856);
nor U13388 (N_13388,N_12559,N_12553);
and U13389 (N_13389,N_13060,N_12728);
or U13390 (N_13390,N_12994,N_13114);
xnor U13391 (N_13391,N_12761,N_12966);
and U13392 (N_13392,N_12943,N_12901);
xnor U13393 (N_13393,N_12993,N_13011);
xor U13394 (N_13394,N_13070,N_12618);
and U13395 (N_13395,N_12903,N_13055);
nand U13396 (N_13396,N_13117,N_12878);
or U13397 (N_13397,N_12649,N_12704);
nor U13398 (N_13398,N_13010,N_13087);
or U13399 (N_13399,N_12515,N_13108);
nand U13400 (N_13400,N_13041,N_12640);
and U13401 (N_13401,N_12671,N_12624);
and U13402 (N_13402,N_12751,N_12992);
or U13403 (N_13403,N_12523,N_12919);
nand U13404 (N_13404,N_12930,N_13037);
xor U13405 (N_13405,N_13112,N_12590);
and U13406 (N_13406,N_12596,N_12547);
and U13407 (N_13407,N_12921,N_12583);
xor U13408 (N_13408,N_12677,N_12972);
and U13409 (N_13409,N_12693,N_12861);
nand U13410 (N_13410,N_12885,N_12927);
nor U13411 (N_13411,N_12949,N_13080);
xor U13412 (N_13412,N_12627,N_12958);
xnor U13413 (N_13413,N_12524,N_12960);
nand U13414 (N_13414,N_12508,N_12827);
nor U13415 (N_13415,N_12637,N_12560);
nand U13416 (N_13416,N_12881,N_12875);
nor U13417 (N_13417,N_13076,N_13043);
or U13418 (N_13418,N_12944,N_12615);
nand U13419 (N_13419,N_12936,N_12906);
xnor U13420 (N_13420,N_12812,N_12699);
xnor U13421 (N_13421,N_12894,N_13005);
or U13422 (N_13422,N_13059,N_12730);
xor U13423 (N_13423,N_12850,N_12656);
xnor U13424 (N_13424,N_12516,N_13057);
nor U13425 (N_13425,N_12605,N_12502);
nand U13426 (N_13426,N_13026,N_12819);
nor U13427 (N_13427,N_13033,N_13015);
and U13428 (N_13428,N_12898,N_12954);
nand U13429 (N_13429,N_12785,N_12535);
or U13430 (N_13430,N_12641,N_12539);
nand U13431 (N_13431,N_12729,N_12563);
xor U13432 (N_13432,N_12984,N_12664);
xnor U13433 (N_13433,N_12813,N_12849);
and U13434 (N_13434,N_12706,N_12600);
or U13435 (N_13435,N_12826,N_12862);
or U13436 (N_13436,N_12545,N_13006);
xor U13437 (N_13437,N_12840,N_12750);
nand U13438 (N_13438,N_12753,N_13005);
xnor U13439 (N_13439,N_12601,N_12698);
nand U13440 (N_13440,N_12631,N_12673);
xnor U13441 (N_13441,N_12834,N_12658);
and U13442 (N_13442,N_12946,N_12895);
nand U13443 (N_13443,N_12635,N_12553);
xor U13444 (N_13444,N_12594,N_12657);
or U13445 (N_13445,N_12814,N_12712);
or U13446 (N_13446,N_12924,N_12963);
nor U13447 (N_13447,N_12974,N_12947);
and U13448 (N_13448,N_13061,N_12937);
nand U13449 (N_13449,N_12721,N_13025);
and U13450 (N_13450,N_12699,N_13053);
and U13451 (N_13451,N_12806,N_12581);
and U13452 (N_13452,N_13008,N_12887);
nand U13453 (N_13453,N_12580,N_13028);
nor U13454 (N_13454,N_12781,N_12836);
or U13455 (N_13455,N_13118,N_13081);
xnor U13456 (N_13456,N_12958,N_12758);
xor U13457 (N_13457,N_12638,N_12847);
nand U13458 (N_13458,N_12806,N_12697);
nand U13459 (N_13459,N_13085,N_12971);
or U13460 (N_13460,N_12597,N_13060);
nand U13461 (N_13461,N_12749,N_12752);
xor U13462 (N_13462,N_12559,N_12710);
and U13463 (N_13463,N_12797,N_12903);
or U13464 (N_13464,N_12740,N_13003);
xnor U13465 (N_13465,N_12941,N_13006);
nand U13466 (N_13466,N_12662,N_12673);
or U13467 (N_13467,N_12836,N_12700);
or U13468 (N_13468,N_12533,N_12511);
xor U13469 (N_13469,N_13079,N_12555);
and U13470 (N_13470,N_12838,N_12670);
nor U13471 (N_13471,N_12964,N_13038);
or U13472 (N_13472,N_12856,N_12771);
or U13473 (N_13473,N_12502,N_12893);
xor U13474 (N_13474,N_13006,N_12888);
or U13475 (N_13475,N_12691,N_12726);
or U13476 (N_13476,N_13019,N_12786);
nand U13477 (N_13477,N_13035,N_13053);
and U13478 (N_13478,N_13113,N_12792);
or U13479 (N_13479,N_12934,N_12817);
or U13480 (N_13480,N_12513,N_12946);
xnor U13481 (N_13481,N_13067,N_12943);
nor U13482 (N_13482,N_12774,N_13075);
nor U13483 (N_13483,N_12738,N_12945);
nor U13484 (N_13484,N_12701,N_12820);
nand U13485 (N_13485,N_12983,N_12869);
and U13486 (N_13486,N_13070,N_12932);
nand U13487 (N_13487,N_12622,N_12839);
xnor U13488 (N_13488,N_12954,N_12510);
or U13489 (N_13489,N_12593,N_12831);
nor U13490 (N_13490,N_13030,N_12891);
and U13491 (N_13491,N_13103,N_12790);
nor U13492 (N_13492,N_12748,N_12873);
nand U13493 (N_13493,N_12553,N_12833);
or U13494 (N_13494,N_12611,N_12643);
and U13495 (N_13495,N_12671,N_12801);
and U13496 (N_13496,N_12850,N_12503);
or U13497 (N_13497,N_13121,N_12978);
nor U13498 (N_13498,N_12912,N_12819);
xnor U13499 (N_13499,N_12574,N_12716);
xnor U13500 (N_13500,N_13112,N_12945);
nand U13501 (N_13501,N_12885,N_12813);
and U13502 (N_13502,N_13096,N_12868);
and U13503 (N_13503,N_13091,N_13031);
xnor U13504 (N_13504,N_12703,N_12913);
xor U13505 (N_13505,N_12647,N_13114);
and U13506 (N_13506,N_13079,N_12660);
and U13507 (N_13507,N_12990,N_12962);
or U13508 (N_13508,N_13016,N_12723);
xnor U13509 (N_13509,N_12783,N_13011);
xnor U13510 (N_13510,N_12880,N_12514);
nand U13511 (N_13511,N_12809,N_12975);
and U13512 (N_13512,N_12736,N_13109);
nor U13513 (N_13513,N_12888,N_12845);
and U13514 (N_13514,N_12884,N_12530);
nand U13515 (N_13515,N_12597,N_13038);
or U13516 (N_13516,N_13036,N_12673);
nor U13517 (N_13517,N_13044,N_12872);
xor U13518 (N_13518,N_12781,N_12693);
or U13519 (N_13519,N_12514,N_12525);
or U13520 (N_13520,N_13093,N_12792);
xor U13521 (N_13521,N_12662,N_12598);
nor U13522 (N_13522,N_12673,N_13099);
or U13523 (N_13523,N_12973,N_12879);
and U13524 (N_13524,N_12722,N_12735);
or U13525 (N_13525,N_12961,N_12638);
xnor U13526 (N_13526,N_12786,N_12716);
and U13527 (N_13527,N_12603,N_12661);
xor U13528 (N_13528,N_12741,N_12569);
nand U13529 (N_13529,N_13074,N_12773);
nor U13530 (N_13530,N_12590,N_12837);
nor U13531 (N_13531,N_12727,N_12743);
nor U13532 (N_13532,N_12711,N_13101);
nor U13533 (N_13533,N_13041,N_12656);
nor U13534 (N_13534,N_12849,N_13118);
nor U13535 (N_13535,N_13072,N_13120);
or U13536 (N_13536,N_12734,N_12706);
and U13537 (N_13537,N_13064,N_13082);
xor U13538 (N_13538,N_12894,N_12813);
or U13539 (N_13539,N_12620,N_13040);
or U13540 (N_13540,N_12622,N_12553);
xor U13541 (N_13541,N_13043,N_12694);
xnor U13542 (N_13542,N_13043,N_13091);
or U13543 (N_13543,N_12591,N_12858);
nor U13544 (N_13544,N_12695,N_12807);
nor U13545 (N_13545,N_12887,N_12671);
nor U13546 (N_13546,N_12632,N_12790);
and U13547 (N_13547,N_12512,N_12528);
nor U13548 (N_13548,N_13082,N_12619);
nor U13549 (N_13549,N_12935,N_12836);
nand U13550 (N_13550,N_12555,N_12770);
and U13551 (N_13551,N_12829,N_12567);
nand U13552 (N_13552,N_13004,N_12541);
xor U13553 (N_13553,N_12781,N_12641);
and U13554 (N_13554,N_12832,N_13052);
xnor U13555 (N_13555,N_12525,N_12773);
nor U13556 (N_13556,N_12519,N_12952);
nand U13557 (N_13557,N_12595,N_12895);
and U13558 (N_13558,N_12675,N_13043);
nor U13559 (N_13559,N_13011,N_12591);
xnor U13560 (N_13560,N_12724,N_12974);
nand U13561 (N_13561,N_12841,N_12916);
and U13562 (N_13562,N_12734,N_12984);
nand U13563 (N_13563,N_12579,N_13016);
xor U13564 (N_13564,N_13047,N_12653);
nor U13565 (N_13565,N_12962,N_12625);
and U13566 (N_13566,N_12630,N_12950);
nor U13567 (N_13567,N_12806,N_12962);
and U13568 (N_13568,N_12747,N_12961);
or U13569 (N_13569,N_12755,N_12627);
xor U13570 (N_13570,N_12567,N_12875);
xor U13571 (N_13571,N_12779,N_12599);
xnor U13572 (N_13572,N_12994,N_12602);
nand U13573 (N_13573,N_12574,N_12900);
xor U13574 (N_13574,N_12541,N_12809);
or U13575 (N_13575,N_12647,N_12729);
and U13576 (N_13576,N_12508,N_12822);
or U13577 (N_13577,N_12914,N_13058);
nand U13578 (N_13578,N_12960,N_12645);
nand U13579 (N_13579,N_12747,N_12850);
xnor U13580 (N_13580,N_12508,N_12510);
or U13581 (N_13581,N_12636,N_12880);
nor U13582 (N_13582,N_13055,N_13065);
or U13583 (N_13583,N_12781,N_12730);
nand U13584 (N_13584,N_12745,N_12567);
and U13585 (N_13585,N_12896,N_12714);
and U13586 (N_13586,N_12761,N_12677);
xor U13587 (N_13587,N_12916,N_12977);
xor U13588 (N_13588,N_13095,N_12988);
xor U13589 (N_13589,N_12528,N_13071);
nand U13590 (N_13590,N_12915,N_12970);
and U13591 (N_13591,N_12587,N_12841);
nor U13592 (N_13592,N_12671,N_13101);
xnor U13593 (N_13593,N_13081,N_12966);
or U13594 (N_13594,N_13009,N_13007);
nand U13595 (N_13595,N_12659,N_12868);
and U13596 (N_13596,N_12961,N_12521);
nor U13597 (N_13597,N_12913,N_13071);
nand U13598 (N_13598,N_12747,N_12939);
and U13599 (N_13599,N_13002,N_12814);
nand U13600 (N_13600,N_12899,N_12813);
nor U13601 (N_13601,N_13074,N_13101);
nand U13602 (N_13602,N_12913,N_12826);
nor U13603 (N_13603,N_12825,N_12785);
xor U13604 (N_13604,N_12826,N_13090);
nor U13605 (N_13605,N_12924,N_12554);
or U13606 (N_13606,N_13006,N_12960);
or U13607 (N_13607,N_12608,N_12872);
and U13608 (N_13608,N_12798,N_13089);
xnor U13609 (N_13609,N_12806,N_12886);
or U13610 (N_13610,N_12750,N_12852);
xnor U13611 (N_13611,N_12981,N_12843);
nor U13612 (N_13612,N_13102,N_12509);
nand U13613 (N_13613,N_12868,N_13025);
and U13614 (N_13614,N_12742,N_12982);
or U13615 (N_13615,N_12897,N_12989);
nand U13616 (N_13616,N_12785,N_12695);
and U13617 (N_13617,N_12764,N_12881);
or U13618 (N_13618,N_12671,N_12807);
nor U13619 (N_13619,N_12598,N_13047);
nor U13620 (N_13620,N_13043,N_12818);
or U13621 (N_13621,N_12521,N_12646);
xnor U13622 (N_13622,N_12505,N_12746);
or U13623 (N_13623,N_12835,N_13073);
nor U13624 (N_13624,N_12910,N_12615);
and U13625 (N_13625,N_12992,N_12746);
nor U13626 (N_13626,N_13098,N_13099);
nand U13627 (N_13627,N_12995,N_12915);
and U13628 (N_13628,N_12843,N_13038);
nor U13629 (N_13629,N_12674,N_12888);
or U13630 (N_13630,N_13068,N_12503);
and U13631 (N_13631,N_12734,N_12934);
and U13632 (N_13632,N_12699,N_12766);
nor U13633 (N_13633,N_12871,N_12519);
nand U13634 (N_13634,N_12794,N_12858);
xnor U13635 (N_13635,N_12681,N_12703);
or U13636 (N_13636,N_12565,N_12845);
nor U13637 (N_13637,N_12679,N_12795);
xnor U13638 (N_13638,N_12953,N_12522);
and U13639 (N_13639,N_12527,N_12673);
xnor U13640 (N_13640,N_12657,N_12560);
and U13641 (N_13641,N_12755,N_12925);
or U13642 (N_13642,N_12728,N_12517);
xnor U13643 (N_13643,N_12748,N_12999);
or U13644 (N_13644,N_12931,N_13007);
and U13645 (N_13645,N_12568,N_12638);
or U13646 (N_13646,N_12714,N_12515);
nor U13647 (N_13647,N_12881,N_12725);
xnor U13648 (N_13648,N_13101,N_12501);
or U13649 (N_13649,N_12702,N_12595);
nor U13650 (N_13650,N_12793,N_12795);
nand U13651 (N_13651,N_12955,N_13084);
nand U13652 (N_13652,N_12984,N_12830);
xnor U13653 (N_13653,N_12889,N_12915);
nor U13654 (N_13654,N_12561,N_13052);
or U13655 (N_13655,N_12769,N_12549);
and U13656 (N_13656,N_12715,N_13095);
nor U13657 (N_13657,N_12669,N_12833);
xnor U13658 (N_13658,N_12988,N_12517);
or U13659 (N_13659,N_12927,N_12836);
and U13660 (N_13660,N_12749,N_12809);
nand U13661 (N_13661,N_12966,N_12595);
nor U13662 (N_13662,N_12959,N_12947);
and U13663 (N_13663,N_12654,N_12946);
nand U13664 (N_13664,N_12556,N_13089);
nor U13665 (N_13665,N_13013,N_13019);
nand U13666 (N_13666,N_12924,N_12964);
or U13667 (N_13667,N_12618,N_12804);
and U13668 (N_13668,N_12548,N_12799);
xor U13669 (N_13669,N_13043,N_13059);
or U13670 (N_13670,N_13032,N_12714);
and U13671 (N_13671,N_12619,N_12894);
or U13672 (N_13672,N_12634,N_12656);
xnor U13673 (N_13673,N_12560,N_13072);
nor U13674 (N_13674,N_12554,N_12953);
or U13675 (N_13675,N_12650,N_12524);
nand U13676 (N_13676,N_12688,N_13107);
nand U13677 (N_13677,N_12726,N_12575);
xor U13678 (N_13678,N_12922,N_12602);
nor U13679 (N_13679,N_13099,N_13005);
or U13680 (N_13680,N_12819,N_13109);
and U13681 (N_13681,N_13108,N_12625);
nand U13682 (N_13682,N_12955,N_13116);
xor U13683 (N_13683,N_13076,N_12745);
nand U13684 (N_13684,N_12770,N_12749);
nand U13685 (N_13685,N_12586,N_13066);
nand U13686 (N_13686,N_12803,N_12574);
or U13687 (N_13687,N_12799,N_12832);
xnor U13688 (N_13688,N_12997,N_12702);
or U13689 (N_13689,N_12628,N_12995);
and U13690 (N_13690,N_12718,N_12565);
nand U13691 (N_13691,N_12536,N_13006);
nor U13692 (N_13692,N_12739,N_13087);
and U13693 (N_13693,N_12550,N_12710);
nor U13694 (N_13694,N_13020,N_12779);
xor U13695 (N_13695,N_13031,N_12936);
xnor U13696 (N_13696,N_12721,N_12527);
nor U13697 (N_13697,N_12651,N_12622);
nor U13698 (N_13698,N_13118,N_12904);
nor U13699 (N_13699,N_12603,N_12629);
xnor U13700 (N_13700,N_13112,N_12729);
nor U13701 (N_13701,N_12643,N_12538);
and U13702 (N_13702,N_12509,N_13114);
or U13703 (N_13703,N_12666,N_12601);
nor U13704 (N_13704,N_12896,N_12894);
or U13705 (N_13705,N_12873,N_12814);
nor U13706 (N_13706,N_12507,N_13067);
nor U13707 (N_13707,N_12917,N_13099);
nor U13708 (N_13708,N_12628,N_12624);
nor U13709 (N_13709,N_12604,N_12708);
and U13710 (N_13710,N_12825,N_12559);
nor U13711 (N_13711,N_13102,N_12566);
and U13712 (N_13712,N_12842,N_12587);
and U13713 (N_13713,N_13039,N_13027);
xor U13714 (N_13714,N_12610,N_13077);
nor U13715 (N_13715,N_12727,N_12945);
or U13716 (N_13716,N_13094,N_13086);
nand U13717 (N_13717,N_12594,N_12563);
nand U13718 (N_13718,N_12999,N_12976);
or U13719 (N_13719,N_12656,N_12751);
nor U13720 (N_13720,N_12625,N_12523);
and U13721 (N_13721,N_12924,N_12921);
xnor U13722 (N_13722,N_12715,N_12569);
nor U13723 (N_13723,N_12535,N_12818);
nand U13724 (N_13724,N_12775,N_12502);
xnor U13725 (N_13725,N_13046,N_12709);
xor U13726 (N_13726,N_12618,N_13030);
nand U13727 (N_13727,N_12901,N_12683);
or U13728 (N_13728,N_12580,N_12544);
nand U13729 (N_13729,N_13009,N_12952);
nor U13730 (N_13730,N_12672,N_12783);
and U13731 (N_13731,N_12591,N_12715);
xor U13732 (N_13732,N_13035,N_12741);
nor U13733 (N_13733,N_12553,N_13017);
nor U13734 (N_13734,N_12629,N_12986);
nand U13735 (N_13735,N_12810,N_12828);
and U13736 (N_13736,N_12678,N_13054);
nor U13737 (N_13737,N_12789,N_13035);
nand U13738 (N_13738,N_12713,N_12924);
or U13739 (N_13739,N_12940,N_12679);
and U13740 (N_13740,N_12896,N_12835);
and U13741 (N_13741,N_13063,N_12740);
xor U13742 (N_13742,N_12637,N_12644);
and U13743 (N_13743,N_12949,N_12967);
nand U13744 (N_13744,N_12546,N_12596);
or U13745 (N_13745,N_12532,N_12655);
xor U13746 (N_13746,N_13018,N_12676);
nor U13747 (N_13747,N_12738,N_12773);
nand U13748 (N_13748,N_12978,N_12629);
and U13749 (N_13749,N_12675,N_12973);
nor U13750 (N_13750,N_13594,N_13542);
or U13751 (N_13751,N_13605,N_13578);
nand U13752 (N_13752,N_13144,N_13279);
nand U13753 (N_13753,N_13725,N_13507);
nand U13754 (N_13754,N_13417,N_13565);
or U13755 (N_13755,N_13681,N_13700);
or U13756 (N_13756,N_13159,N_13195);
nor U13757 (N_13757,N_13416,N_13495);
nor U13758 (N_13758,N_13713,N_13561);
xnor U13759 (N_13759,N_13459,N_13454);
nor U13760 (N_13760,N_13723,N_13566);
xor U13761 (N_13761,N_13170,N_13320);
nor U13762 (N_13762,N_13656,N_13240);
nor U13763 (N_13763,N_13152,N_13145);
or U13764 (N_13764,N_13233,N_13692);
xor U13765 (N_13765,N_13512,N_13601);
xnor U13766 (N_13766,N_13284,N_13138);
and U13767 (N_13767,N_13410,N_13552);
xor U13768 (N_13768,N_13608,N_13161);
and U13769 (N_13769,N_13401,N_13160);
xor U13770 (N_13770,N_13272,N_13215);
and U13771 (N_13771,N_13529,N_13588);
or U13772 (N_13772,N_13423,N_13206);
xor U13773 (N_13773,N_13386,N_13438);
and U13774 (N_13774,N_13217,N_13576);
and U13775 (N_13775,N_13388,N_13347);
nor U13776 (N_13776,N_13475,N_13245);
nand U13777 (N_13777,N_13338,N_13319);
nor U13778 (N_13778,N_13327,N_13406);
nand U13779 (N_13779,N_13137,N_13352);
nand U13780 (N_13780,N_13573,N_13719);
or U13781 (N_13781,N_13168,N_13526);
and U13782 (N_13782,N_13182,N_13505);
xnor U13783 (N_13783,N_13627,N_13707);
nand U13784 (N_13784,N_13645,N_13664);
nand U13785 (N_13785,N_13580,N_13239);
nor U13786 (N_13786,N_13612,N_13361);
nor U13787 (N_13787,N_13541,N_13421);
or U13788 (N_13788,N_13194,N_13235);
xnor U13789 (N_13789,N_13722,N_13395);
nor U13790 (N_13790,N_13596,N_13616);
nand U13791 (N_13791,N_13367,N_13282);
or U13792 (N_13792,N_13589,N_13355);
and U13793 (N_13793,N_13130,N_13344);
nand U13794 (N_13794,N_13415,N_13521);
or U13795 (N_13795,N_13516,N_13639);
or U13796 (N_13796,N_13356,N_13610);
xor U13797 (N_13797,N_13362,N_13726);
nand U13798 (N_13798,N_13568,N_13582);
or U13799 (N_13799,N_13398,N_13702);
and U13800 (N_13800,N_13525,N_13301);
nand U13801 (N_13801,N_13624,N_13285);
or U13802 (N_13802,N_13326,N_13538);
nand U13803 (N_13803,N_13293,N_13557);
xor U13804 (N_13804,N_13228,N_13729);
nand U13805 (N_13805,N_13522,N_13597);
nor U13806 (N_13806,N_13489,N_13611);
nand U13807 (N_13807,N_13308,N_13218);
or U13808 (N_13808,N_13405,N_13185);
and U13809 (N_13809,N_13317,N_13188);
nor U13810 (N_13810,N_13126,N_13671);
nand U13811 (N_13811,N_13314,N_13472);
nand U13812 (N_13812,N_13389,N_13141);
and U13813 (N_13813,N_13404,N_13211);
xor U13814 (N_13814,N_13368,N_13618);
or U13815 (N_13815,N_13278,N_13135);
nor U13816 (N_13816,N_13704,N_13458);
and U13817 (N_13817,N_13520,N_13174);
or U13818 (N_13818,N_13148,N_13519);
xor U13819 (N_13819,N_13378,N_13440);
xor U13820 (N_13820,N_13237,N_13654);
nor U13821 (N_13821,N_13457,N_13387);
or U13822 (N_13822,N_13246,N_13657);
xnor U13823 (N_13823,N_13331,N_13393);
nor U13824 (N_13824,N_13658,N_13465);
nand U13825 (N_13825,N_13744,N_13470);
nor U13826 (N_13826,N_13383,N_13321);
or U13827 (N_13827,N_13251,N_13176);
and U13828 (N_13828,N_13517,N_13456);
or U13829 (N_13829,N_13603,N_13305);
and U13830 (N_13830,N_13180,N_13644);
nand U13831 (N_13831,N_13183,N_13379);
xor U13832 (N_13832,N_13660,N_13701);
or U13833 (N_13833,N_13675,N_13679);
and U13834 (N_13834,N_13150,N_13452);
nor U13835 (N_13835,N_13167,N_13162);
and U13836 (N_13836,N_13382,N_13419);
or U13837 (N_13837,N_13665,N_13689);
and U13838 (N_13838,N_13477,N_13177);
and U13839 (N_13839,N_13436,N_13297);
nor U13840 (N_13840,N_13740,N_13376);
nand U13841 (N_13841,N_13418,N_13289);
nand U13842 (N_13842,N_13346,N_13207);
or U13843 (N_13843,N_13351,N_13636);
and U13844 (N_13844,N_13254,N_13492);
nand U13845 (N_13845,N_13553,N_13370);
xor U13846 (N_13846,N_13306,N_13140);
or U13847 (N_13847,N_13128,N_13513);
xor U13848 (N_13848,N_13545,N_13485);
and U13849 (N_13849,N_13337,N_13621);
xor U13850 (N_13850,N_13163,N_13455);
and U13851 (N_13851,N_13313,N_13201);
xnor U13852 (N_13852,N_13697,N_13662);
nor U13853 (N_13853,N_13742,N_13585);
and U13854 (N_13854,N_13154,N_13486);
nor U13855 (N_13855,N_13695,N_13350);
and U13856 (N_13856,N_13175,N_13699);
nor U13857 (N_13857,N_13508,N_13435);
nand U13858 (N_13858,N_13609,N_13734);
nand U13859 (N_13859,N_13502,N_13478);
nand U13860 (N_13860,N_13631,N_13226);
or U13861 (N_13861,N_13515,N_13666);
and U13862 (N_13862,N_13592,N_13225);
nand U13863 (N_13863,N_13655,N_13493);
xnor U13864 (N_13864,N_13374,N_13295);
or U13865 (N_13865,N_13728,N_13528);
nand U13866 (N_13866,N_13205,N_13504);
nor U13867 (N_13867,N_13748,N_13577);
or U13868 (N_13868,N_13550,N_13635);
and U13869 (N_13869,N_13506,N_13271);
nor U13870 (N_13870,N_13646,N_13222);
and U13871 (N_13871,N_13381,N_13567);
xor U13872 (N_13872,N_13511,N_13446);
or U13873 (N_13873,N_13524,N_13433);
nor U13874 (N_13874,N_13281,N_13358);
and U13875 (N_13875,N_13709,N_13287);
nand U13876 (N_13876,N_13536,N_13718);
nand U13877 (N_13877,N_13659,N_13441);
nor U13878 (N_13878,N_13310,N_13746);
xor U13879 (N_13879,N_13261,N_13743);
or U13880 (N_13880,N_13309,N_13210);
xnor U13881 (N_13881,N_13431,N_13745);
and U13882 (N_13882,N_13187,N_13330);
nand U13883 (N_13883,N_13533,N_13628);
nor U13884 (N_13884,N_13149,N_13684);
nor U13885 (N_13885,N_13706,N_13527);
nand U13886 (N_13886,N_13680,N_13498);
xor U13887 (N_13887,N_13333,N_13257);
and U13888 (N_13888,N_13633,N_13230);
and U13889 (N_13889,N_13357,N_13209);
xnor U13890 (N_13890,N_13291,N_13643);
nand U13891 (N_13891,N_13461,N_13208);
and U13892 (N_13892,N_13348,N_13220);
or U13893 (N_13893,N_13641,N_13572);
xor U13894 (N_13894,N_13721,N_13501);
or U13895 (N_13895,N_13634,N_13638);
or U13896 (N_13896,N_13280,N_13464);
xor U13897 (N_13897,N_13453,N_13584);
nor U13898 (N_13898,N_13411,N_13685);
nand U13899 (N_13899,N_13693,N_13364);
or U13900 (N_13900,N_13648,N_13642);
nand U13901 (N_13901,N_13676,N_13476);
xnor U13902 (N_13902,N_13224,N_13328);
xnor U13903 (N_13903,N_13617,N_13575);
nor U13904 (N_13904,N_13630,N_13715);
or U13905 (N_13905,N_13397,N_13593);
nand U13906 (N_13906,N_13683,N_13143);
nor U13907 (N_13907,N_13467,N_13710);
and U13908 (N_13908,N_13165,N_13409);
xnor U13909 (N_13909,N_13727,N_13275);
and U13910 (N_13910,N_13136,N_13652);
nor U13911 (N_13911,N_13298,N_13329);
nor U13912 (N_13912,N_13733,N_13559);
nor U13913 (N_13913,N_13324,N_13653);
xnor U13914 (N_13914,N_13200,N_13428);
or U13915 (N_13915,N_13549,N_13178);
and U13916 (N_13916,N_13236,N_13626);
nor U13917 (N_13917,N_13345,N_13434);
xnor U13918 (N_13918,N_13266,N_13544);
and U13919 (N_13919,N_13373,N_13640);
and U13920 (N_13920,N_13496,N_13142);
xor U13921 (N_13921,N_13663,N_13164);
or U13922 (N_13922,N_13340,N_13420);
nor U13923 (N_13923,N_13335,N_13602);
xnor U13924 (N_13924,N_13203,N_13259);
nand U13925 (N_13925,N_13392,N_13372);
nand U13926 (N_13926,N_13412,N_13248);
or U13927 (N_13927,N_13385,N_13131);
xor U13928 (N_13928,N_13290,N_13625);
or U13929 (N_13929,N_13484,N_13294);
or U13930 (N_13930,N_13427,N_13384);
xnor U13931 (N_13931,N_13125,N_13546);
nor U13932 (N_13932,N_13463,N_13682);
nand U13933 (N_13933,N_13623,N_13479);
xnor U13934 (N_13934,N_13686,N_13637);
xnor U13935 (N_13935,N_13468,N_13619);
xor U13936 (N_13936,N_13336,N_13363);
nand U13937 (N_13937,N_13413,N_13668);
and U13938 (N_13938,N_13156,N_13252);
and U13939 (N_13939,N_13667,N_13717);
nand U13940 (N_13940,N_13179,N_13139);
and U13941 (N_13941,N_13547,N_13322);
nor U13942 (N_13942,N_13551,N_13450);
or U13943 (N_13943,N_13651,N_13229);
and U13944 (N_13944,N_13243,N_13570);
xor U13945 (N_13945,N_13724,N_13469);
or U13946 (N_13946,N_13255,N_13197);
nand U13947 (N_13947,N_13445,N_13391);
nand U13948 (N_13948,N_13134,N_13661);
xor U13949 (N_13949,N_13543,N_13482);
xor U13950 (N_13950,N_13554,N_13292);
and U13951 (N_13951,N_13583,N_13153);
nor U13952 (N_13952,N_13598,N_13615);
and U13953 (N_13953,N_13678,N_13253);
or U13954 (N_13954,N_13151,N_13696);
nor U13955 (N_13955,N_13443,N_13171);
xnor U13956 (N_13956,N_13447,N_13672);
or U13957 (N_13957,N_13739,N_13562);
xor U13958 (N_13958,N_13269,N_13741);
nor U13959 (N_13959,N_13155,N_13198);
and U13960 (N_13960,N_13720,N_13560);
or U13961 (N_13961,N_13451,N_13747);
nor U13962 (N_13962,N_13614,N_13586);
and U13963 (N_13963,N_13196,N_13369);
nand U13964 (N_13964,N_13181,N_13703);
or U13965 (N_13965,N_13343,N_13669);
xor U13966 (N_13966,N_13147,N_13189);
nand U13967 (N_13967,N_13673,N_13303);
and U13968 (N_13968,N_13341,N_13213);
xnor U13969 (N_13969,N_13166,N_13539);
xor U13970 (N_13970,N_13499,N_13234);
or U13971 (N_13971,N_13339,N_13315);
nor U13972 (N_13972,N_13256,N_13221);
xnor U13973 (N_13973,N_13714,N_13349);
xnor U13974 (N_13974,N_13371,N_13318);
and U13975 (N_13975,N_13587,N_13311);
nand U13976 (N_13976,N_13555,N_13563);
nand U13977 (N_13977,N_13242,N_13494);
nor U13978 (N_13978,N_13227,N_13705);
xnor U13979 (N_13979,N_13591,N_13283);
nor U13980 (N_13980,N_13247,N_13731);
nand U13981 (N_13981,N_13432,N_13241);
and U13982 (N_13982,N_13414,N_13487);
or U13983 (N_13983,N_13500,N_13223);
or U13984 (N_13984,N_13250,N_13408);
xnor U13985 (N_13985,N_13523,N_13425);
and U13986 (N_13986,N_13647,N_13273);
nand U13987 (N_13987,N_13390,N_13690);
nand U13988 (N_13988,N_13249,N_13574);
or U13989 (N_13989,N_13300,N_13540);
and U13990 (N_13990,N_13444,N_13579);
xor U13991 (N_13991,N_13202,N_13606);
nand U13992 (N_13992,N_13276,N_13730);
nand U13993 (N_13993,N_13629,N_13490);
nor U13994 (N_13994,N_13691,N_13407);
nor U13995 (N_13995,N_13716,N_13564);
nand U13996 (N_13996,N_13262,N_13263);
xor U13997 (N_13997,N_13510,N_13732);
xnor U13998 (N_13998,N_13437,N_13749);
or U13999 (N_13999,N_13286,N_13158);
xnor U14000 (N_14000,N_13342,N_13480);
and U14001 (N_14001,N_13632,N_13622);
and U14002 (N_14002,N_13172,N_13191);
xor U14003 (N_14003,N_13360,N_13497);
xor U14004 (N_14004,N_13366,N_13534);
and U14005 (N_14005,N_13238,N_13535);
and U14006 (N_14006,N_13571,N_13449);
nor U14007 (N_14007,N_13190,N_13132);
or U14008 (N_14008,N_13157,N_13698);
nor U14009 (N_14009,N_13354,N_13649);
or U14010 (N_14010,N_13316,N_13424);
or U14011 (N_14011,N_13442,N_13460);
and U14012 (N_14012,N_13670,N_13556);
nand U14013 (N_14013,N_13264,N_13377);
or U14014 (N_14014,N_13288,N_13270);
or U14015 (N_14015,N_13595,N_13323);
nor U14016 (N_14016,N_13491,N_13129);
xnor U14017 (N_14017,N_13509,N_13334);
nand U14018 (N_14018,N_13604,N_13481);
and U14019 (N_14019,N_13192,N_13466);
and U14020 (N_14020,N_13268,N_13199);
and U14021 (N_14021,N_13133,N_13711);
xnor U14022 (N_14022,N_13503,N_13274);
xor U14023 (N_14023,N_13312,N_13712);
nor U14024 (N_14024,N_13216,N_13267);
xor U14025 (N_14025,N_13402,N_13400);
or U14026 (N_14026,N_13173,N_13325);
nor U14027 (N_14027,N_13394,N_13212);
and U14028 (N_14028,N_13296,N_13375);
or U14029 (N_14029,N_13204,N_13687);
or U14030 (N_14030,N_13214,N_13530);
nor U14031 (N_14031,N_13403,N_13677);
nand U14032 (N_14032,N_13548,N_13532);
or U14033 (N_14033,N_13558,N_13429);
xnor U14034 (N_14034,N_13302,N_13694);
nor U14035 (N_14035,N_13736,N_13537);
nand U14036 (N_14036,N_13353,N_13307);
nor U14037 (N_14037,N_13399,N_13674);
and U14038 (N_14038,N_13514,N_13483);
and U14039 (N_14039,N_13193,N_13332);
and U14040 (N_14040,N_13708,N_13299);
nand U14041 (N_14041,N_13184,N_13232);
or U14042 (N_14042,N_13569,N_13439);
xor U14043 (N_14043,N_13737,N_13581);
nor U14044 (N_14044,N_13258,N_13359);
nor U14045 (N_14045,N_13650,N_13396);
and U14046 (N_14046,N_13471,N_13474);
nand U14047 (N_14047,N_13473,N_13607);
nand U14048 (N_14048,N_13277,N_13365);
or U14049 (N_14049,N_13620,N_13304);
xnor U14050 (N_14050,N_13688,N_13146);
xnor U14051 (N_14051,N_13426,N_13590);
xor U14052 (N_14052,N_13231,N_13422);
nand U14053 (N_14053,N_13735,N_13462);
and U14054 (N_14054,N_13518,N_13738);
nand U14055 (N_14055,N_13219,N_13265);
xnor U14056 (N_14056,N_13244,N_13448);
or U14057 (N_14057,N_13531,N_13169);
or U14058 (N_14058,N_13260,N_13488);
xnor U14059 (N_14059,N_13127,N_13613);
xnor U14060 (N_14060,N_13380,N_13186);
and U14061 (N_14061,N_13599,N_13600);
or U14062 (N_14062,N_13430,N_13385);
and U14063 (N_14063,N_13644,N_13550);
or U14064 (N_14064,N_13290,N_13244);
xnor U14065 (N_14065,N_13710,N_13317);
nor U14066 (N_14066,N_13654,N_13552);
nand U14067 (N_14067,N_13688,N_13647);
nor U14068 (N_14068,N_13608,N_13514);
or U14069 (N_14069,N_13132,N_13413);
xnor U14070 (N_14070,N_13573,N_13241);
or U14071 (N_14071,N_13383,N_13433);
and U14072 (N_14072,N_13539,N_13153);
nand U14073 (N_14073,N_13163,N_13504);
and U14074 (N_14074,N_13291,N_13295);
nor U14075 (N_14075,N_13638,N_13661);
nor U14076 (N_14076,N_13563,N_13564);
xnor U14077 (N_14077,N_13579,N_13391);
or U14078 (N_14078,N_13520,N_13425);
nor U14079 (N_14079,N_13158,N_13527);
xnor U14080 (N_14080,N_13169,N_13667);
or U14081 (N_14081,N_13550,N_13456);
nand U14082 (N_14082,N_13291,N_13692);
and U14083 (N_14083,N_13467,N_13132);
nor U14084 (N_14084,N_13498,N_13474);
and U14085 (N_14085,N_13610,N_13603);
nand U14086 (N_14086,N_13637,N_13432);
xnor U14087 (N_14087,N_13708,N_13696);
nand U14088 (N_14088,N_13208,N_13714);
xnor U14089 (N_14089,N_13286,N_13714);
and U14090 (N_14090,N_13572,N_13128);
or U14091 (N_14091,N_13252,N_13657);
or U14092 (N_14092,N_13275,N_13367);
nand U14093 (N_14093,N_13702,N_13164);
nand U14094 (N_14094,N_13200,N_13258);
and U14095 (N_14095,N_13243,N_13554);
xor U14096 (N_14096,N_13444,N_13536);
or U14097 (N_14097,N_13369,N_13749);
xor U14098 (N_14098,N_13450,N_13387);
nor U14099 (N_14099,N_13579,N_13455);
nand U14100 (N_14100,N_13237,N_13129);
xnor U14101 (N_14101,N_13224,N_13269);
xnor U14102 (N_14102,N_13552,N_13251);
nor U14103 (N_14103,N_13399,N_13167);
and U14104 (N_14104,N_13610,N_13459);
nor U14105 (N_14105,N_13550,N_13489);
nor U14106 (N_14106,N_13718,N_13326);
xnor U14107 (N_14107,N_13563,N_13206);
nand U14108 (N_14108,N_13482,N_13318);
or U14109 (N_14109,N_13475,N_13556);
nor U14110 (N_14110,N_13547,N_13689);
xnor U14111 (N_14111,N_13596,N_13496);
xor U14112 (N_14112,N_13435,N_13329);
xnor U14113 (N_14113,N_13171,N_13745);
nand U14114 (N_14114,N_13584,N_13489);
xnor U14115 (N_14115,N_13388,N_13340);
nand U14116 (N_14116,N_13440,N_13354);
nor U14117 (N_14117,N_13378,N_13688);
or U14118 (N_14118,N_13196,N_13642);
nand U14119 (N_14119,N_13131,N_13628);
nand U14120 (N_14120,N_13298,N_13461);
or U14121 (N_14121,N_13344,N_13235);
and U14122 (N_14122,N_13314,N_13175);
and U14123 (N_14123,N_13528,N_13144);
xnor U14124 (N_14124,N_13567,N_13593);
nand U14125 (N_14125,N_13503,N_13421);
and U14126 (N_14126,N_13583,N_13376);
nand U14127 (N_14127,N_13314,N_13231);
xnor U14128 (N_14128,N_13732,N_13255);
or U14129 (N_14129,N_13164,N_13374);
and U14130 (N_14130,N_13555,N_13581);
nand U14131 (N_14131,N_13339,N_13560);
or U14132 (N_14132,N_13673,N_13618);
or U14133 (N_14133,N_13385,N_13721);
and U14134 (N_14134,N_13667,N_13274);
or U14135 (N_14135,N_13194,N_13206);
or U14136 (N_14136,N_13428,N_13218);
or U14137 (N_14137,N_13182,N_13177);
and U14138 (N_14138,N_13254,N_13276);
or U14139 (N_14139,N_13194,N_13541);
and U14140 (N_14140,N_13180,N_13468);
nand U14141 (N_14141,N_13472,N_13399);
xor U14142 (N_14142,N_13146,N_13571);
or U14143 (N_14143,N_13130,N_13477);
or U14144 (N_14144,N_13730,N_13556);
nor U14145 (N_14145,N_13324,N_13358);
and U14146 (N_14146,N_13476,N_13289);
or U14147 (N_14147,N_13616,N_13250);
nand U14148 (N_14148,N_13616,N_13299);
nor U14149 (N_14149,N_13186,N_13632);
xor U14150 (N_14150,N_13465,N_13401);
xnor U14151 (N_14151,N_13625,N_13227);
or U14152 (N_14152,N_13192,N_13150);
nand U14153 (N_14153,N_13488,N_13657);
nor U14154 (N_14154,N_13581,N_13394);
or U14155 (N_14155,N_13220,N_13487);
nand U14156 (N_14156,N_13470,N_13154);
nor U14157 (N_14157,N_13521,N_13311);
nor U14158 (N_14158,N_13177,N_13279);
nor U14159 (N_14159,N_13571,N_13717);
nand U14160 (N_14160,N_13288,N_13491);
nand U14161 (N_14161,N_13428,N_13582);
nand U14162 (N_14162,N_13451,N_13161);
nor U14163 (N_14163,N_13192,N_13431);
xnor U14164 (N_14164,N_13280,N_13626);
xor U14165 (N_14165,N_13300,N_13285);
and U14166 (N_14166,N_13526,N_13233);
or U14167 (N_14167,N_13708,N_13304);
nand U14168 (N_14168,N_13551,N_13303);
or U14169 (N_14169,N_13313,N_13637);
xor U14170 (N_14170,N_13179,N_13248);
nor U14171 (N_14171,N_13482,N_13308);
nand U14172 (N_14172,N_13348,N_13439);
nand U14173 (N_14173,N_13486,N_13249);
nand U14174 (N_14174,N_13494,N_13287);
nor U14175 (N_14175,N_13214,N_13682);
nor U14176 (N_14176,N_13362,N_13582);
nand U14177 (N_14177,N_13645,N_13466);
xnor U14178 (N_14178,N_13616,N_13544);
nor U14179 (N_14179,N_13598,N_13218);
nor U14180 (N_14180,N_13626,N_13494);
and U14181 (N_14181,N_13631,N_13196);
and U14182 (N_14182,N_13274,N_13473);
nand U14183 (N_14183,N_13494,N_13261);
or U14184 (N_14184,N_13141,N_13340);
nor U14185 (N_14185,N_13469,N_13648);
nor U14186 (N_14186,N_13583,N_13220);
and U14187 (N_14187,N_13698,N_13452);
and U14188 (N_14188,N_13277,N_13490);
nor U14189 (N_14189,N_13573,N_13609);
and U14190 (N_14190,N_13700,N_13470);
and U14191 (N_14191,N_13676,N_13380);
nor U14192 (N_14192,N_13527,N_13500);
xnor U14193 (N_14193,N_13264,N_13125);
nor U14194 (N_14194,N_13701,N_13494);
xnor U14195 (N_14195,N_13341,N_13602);
or U14196 (N_14196,N_13260,N_13216);
nor U14197 (N_14197,N_13388,N_13265);
or U14198 (N_14198,N_13296,N_13609);
and U14199 (N_14199,N_13624,N_13660);
nand U14200 (N_14200,N_13445,N_13201);
and U14201 (N_14201,N_13308,N_13523);
nand U14202 (N_14202,N_13666,N_13335);
nand U14203 (N_14203,N_13125,N_13297);
nand U14204 (N_14204,N_13700,N_13482);
nor U14205 (N_14205,N_13629,N_13209);
or U14206 (N_14206,N_13692,N_13718);
or U14207 (N_14207,N_13595,N_13163);
or U14208 (N_14208,N_13255,N_13666);
or U14209 (N_14209,N_13131,N_13725);
or U14210 (N_14210,N_13419,N_13576);
nor U14211 (N_14211,N_13224,N_13717);
and U14212 (N_14212,N_13607,N_13175);
and U14213 (N_14213,N_13449,N_13209);
nand U14214 (N_14214,N_13688,N_13282);
nor U14215 (N_14215,N_13321,N_13510);
nand U14216 (N_14216,N_13637,N_13565);
and U14217 (N_14217,N_13484,N_13586);
nand U14218 (N_14218,N_13470,N_13632);
xor U14219 (N_14219,N_13379,N_13411);
and U14220 (N_14220,N_13201,N_13521);
or U14221 (N_14221,N_13389,N_13125);
nand U14222 (N_14222,N_13369,N_13653);
and U14223 (N_14223,N_13563,N_13389);
and U14224 (N_14224,N_13289,N_13272);
xor U14225 (N_14225,N_13469,N_13307);
nor U14226 (N_14226,N_13278,N_13691);
or U14227 (N_14227,N_13654,N_13432);
xor U14228 (N_14228,N_13465,N_13335);
nand U14229 (N_14229,N_13411,N_13538);
or U14230 (N_14230,N_13346,N_13394);
or U14231 (N_14231,N_13317,N_13426);
xnor U14232 (N_14232,N_13199,N_13304);
and U14233 (N_14233,N_13574,N_13626);
nor U14234 (N_14234,N_13279,N_13357);
nand U14235 (N_14235,N_13421,N_13706);
nor U14236 (N_14236,N_13534,N_13399);
nor U14237 (N_14237,N_13473,N_13404);
nand U14238 (N_14238,N_13304,N_13562);
nor U14239 (N_14239,N_13720,N_13219);
xor U14240 (N_14240,N_13447,N_13621);
or U14241 (N_14241,N_13415,N_13313);
nor U14242 (N_14242,N_13694,N_13298);
or U14243 (N_14243,N_13363,N_13200);
nand U14244 (N_14244,N_13472,N_13565);
nor U14245 (N_14245,N_13446,N_13259);
nor U14246 (N_14246,N_13185,N_13221);
nor U14247 (N_14247,N_13628,N_13359);
or U14248 (N_14248,N_13465,N_13184);
xnor U14249 (N_14249,N_13369,N_13654);
nor U14250 (N_14250,N_13552,N_13725);
and U14251 (N_14251,N_13304,N_13591);
nand U14252 (N_14252,N_13435,N_13658);
and U14253 (N_14253,N_13323,N_13724);
nand U14254 (N_14254,N_13643,N_13390);
nor U14255 (N_14255,N_13587,N_13432);
nor U14256 (N_14256,N_13444,N_13368);
nand U14257 (N_14257,N_13615,N_13335);
nand U14258 (N_14258,N_13602,N_13139);
xor U14259 (N_14259,N_13614,N_13308);
or U14260 (N_14260,N_13484,N_13475);
nor U14261 (N_14261,N_13422,N_13665);
or U14262 (N_14262,N_13669,N_13396);
or U14263 (N_14263,N_13137,N_13305);
nor U14264 (N_14264,N_13558,N_13353);
nor U14265 (N_14265,N_13179,N_13173);
and U14266 (N_14266,N_13499,N_13468);
nand U14267 (N_14267,N_13421,N_13469);
and U14268 (N_14268,N_13599,N_13530);
or U14269 (N_14269,N_13633,N_13656);
xor U14270 (N_14270,N_13740,N_13735);
nand U14271 (N_14271,N_13284,N_13609);
and U14272 (N_14272,N_13513,N_13185);
and U14273 (N_14273,N_13705,N_13129);
xnor U14274 (N_14274,N_13444,N_13624);
nand U14275 (N_14275,N_13690,N_13176);
xnor U14276 (N_14276,N_13576,N_13593);
nand U14277 (N_14277,N_13546,N_13748);
xnor U14278 (N_14278,N_13289,N_13125);
nor U14279 (N_14279,N_13521,N_13550);
nor U14280 (N_14280,N_13551,N_13732);
or U14281 (N_14281,N_13229,N_13470);
and U14282 (N_14282,N_13558,N_13221);
nor U14283 (N_14283,N_13428,N_13182);
xor U14284 (N_14284,N_13749,N_13196);
and U14285 (N_14285,N_13547,N_13193);
or U14286 (N_14286,N_13460,N_13147);
or U14287 (N_14287,N_13699,N_13683);
or U14288 (N_14288,N_13293,N_13740);
nand U14289 (N_14289,N_13145,N_13194);
nor U14290 (N_14290,N_13747,N_13257);
nor U14291 (N_14291,N_13181,N_13256);
nor U14292 (N_14292,N_13636,N_13384);
nor U14293 (N_14293,N_13533,N_13668);
nand U14294 (N_14294,N_13382,N_13614);
nand U14295 (N_14295,N_13628,N_13388);
xnor U14296 (N_14296,N_13405,N_13473);
or U14297 (N_14297,N_13480,N_13357);
and U14298 (N_14298,N_13348,N_13340);
nand U14299 (N_14299,N_13402,N_13321);
and U14300 (N_14300,N_13662,N_13239);
and U14301 (N_14301,N_13308,N_13262);
nor U14302 (N_14302,N_13545,N_13372);
and U14303 (N_14303,N_13547,N_13555);
xnor U14304 (N_14304,N_13146,N_13496);
xor U14305 (N_14305,N_13633,N_13415);
or U14306 (N_14306,N_13522,N_13287);
xor U14307 (N_14307,N_13543,N_13531);
and U14308 (N_14308,N_13537,N_13215);
or U14309 (N_14309,N_13386,N_13540);
nand U14310 (N_14310,N_13350,N_13540);
xor U14311 (N_14311,N_13344,N_13746);
nand U14312 (N_14312,N_13568,N_13579);
nand U14313 (N_14313,N_13129,N_13221);
and U14314 (N_14314,N_13199,N_13314);
xor U14315 (N_14315,N_13494,N_13483);
nand U14316 (N_14316,N_13171,N_13615);
and U14317 (N_14317,N_13619,N_13301);
or U14318 (N_14318,N_13687,N_13294);
nor U14319 (N_14319,N_13432,N_13176);
and U14320 (N_14320,N_13459,N_13282);
xor U14321 (N_14321,N_13555,N_13177);
nor U14322 (N_14322,N_13323,N_13265);
or U14323 (N_14323,N_13684,N_13733);
nor U14324 (N_14324,N_13491,N_13502);
xnor U14325 (N_14325,N_13617,N_13646);
or U14326 (N_14326,N_13282,N_13749);
nand U14327 (N_14327,N_13552,N_13306);
xor U14328 (N_14328,N_13668,N_13435);
nor U14329 (N_14329,N_13648,N_13278);
or U14330 (N_14330,N_13589,N_13721);
nand U14331 (N_14331,N_13742,N_13646);
nand U14332 (N_14332,N_13700,N_13452);
xnor U14333 (N_14333,N_13179,N_13374);
nand U14334 (N_14334,N_13247,N_13445);
and U14335 (N_14335,N_13135,N_13443);
nand U14336 (N_14336,N_13729,N_13150);
and U14337 (N_14337,N_13577,N_13685);
nor U14338 (N_14338,N_13557,N_13625);
nor U14339 (N_14339,N_13488,N_13555);
nand U14340 (N_14340,N_13422,N_13287);
xor U14341 (N_14341,N_13669,N_13197);
nor U14342 (N_14342,N_13274,N_13670);
or U14343 (N_14343,N_13138,N_13161);
or U14344 (N_14344,N_13329,N_13586);
nand U14345 (N_14345,N_13596,N_13178);
nor U14346 (N_14346,N_13170,N_13587);
xor U14347 (N_14347,N_13463,N_13604);
nor U14348 (N_14348,N_13144,N_13445);
nor U14349 (N_14349,N_13397,N_13157);
nor U14350 (N_14350,N_13269,N_13276);
nor U14351 (N_14351,N_13376,N_13459);
or U14352 (N_14352,N_13596,N_13153);
or U14353 (N_14353,N_13131,N_13448);
nor U14354 (N_14354,N_13266,N_13713);
xor U14355 (N_14355,N_13427,N_13385);
and U14356 (N_14356,N_13390,N_13488);
xor U14357 (N_14357,N_13424,N_13488);
nor U14358 (N_14358,N_13492,N_13138);
xnor U14359 (N_14359,N_13241,N_13204);
xnor U14360 (N_14360,N_13670,N_13492);
xnor U14361 (N_14361,N_13515,N_13133);
nand U14362 (N_14362,N_13672,N_13652);
nand U14363 (N_14363,N_13133,N_13265);
and U14364 (N_14364,N_13620,N_13417);
nor U14365 (N_14365,N_13526,N_13455);
nand U14366 (N_14366,N_13649,N_13464);
nor U14367 (N_14367,N_13708,N_13662);
or U14368 (N_14368,N_13265,N_13736);
nor U14369 (N_14369,N_13171,N_13153);
nand U14370 (N_14370,N_13698,N_13630);
and U14371 (N_14371,N_13479,N_13734);
or U14372 (N_14372,N_13652,N_13573);
or U14373 (N_14373,N_13720,N_13582);
and U14374 (N_14374,N_13164,N_13185);
and U14375 (N_14375,N_14194,N_14333);
nor U14376 (N_14376,N_14061,N_14321);
and U14377 (N_14377,N_14329,N_14224);
nor U14378 (N_14378,N_14093,N_14356);
xnor U14379 (N_14379,N_13774,N_14341);
nor U14380 (N_14380,N_13933,N_13794);
and U14381 (N_14381,N_13989,N_13752);
nand U14382 (N_14382,N_14002,N_14016);
xor U14383 (N_14383,N_13833,N_13859);
xnor U14384 (N_14384,N_13764,N_13891);
or U14385 (N_14385,N_13909,N_14334);
or U14386 (N_14386,N_13876,N_14342);
nand U14387 (N_14387,N_14137,N_14105);
nand U14388 (N_14388,N_14279,N_14115);
nor U14389 (N_14389,N_14070,N_13816);
xnor U14390 (N_14390,N_13791,N_14065);
nor U14391 (N_14391,N_13836,N_13968);
nor U14392 (N_14392,N_13982,N_13939);
xor U14393 (N_14393,N_13799,N_13849);
nand U14394 (N_14394,N_14191,N_14271);
nor U14395 (N_14395,N_13823,N_13879);
xor U14396 (N_14396,N_14017,N_14108);
nor U14397 (N_14397,N_14063,N_13838);
xnor U14398 (N_14398,N_14074,N_13922);
and U14399 (N_14399,N_13938,N_14230);
nor U14400 (N_14400,N_14192,N_13897);
nand U14401 (N_14401,N_14285,N_14216);
and U14402 (N_14402,N_13906,N_14261);
nand U14403 (N_14403,N_14225,N_14210);
xor U14404 (N_14404,N_13918,N_14220);
nand U14405 (N_14405,N_14046,N_13796);
nand U14406 (N_14406,N_14033,N_14109);
nor U14407 (N_14407,N_14123,N_13821);
or U14408 (N_14408,N_14095,N_14305);
nor U14409 (N_14409,N_14255,N_14055);
nand U14410 (N_14410,N_14314,N_13957);
nor U14411 (N_14411,N_13948,N_14252);
nand U14412 (N_14412,N_13777,N_14098);
nand U14413 (N_14413,N_14096,N_14136);
nor U14414 (N_14414,N_14286,N_13868);
and U14415 (N_14415,N_14080,N_13901);
or U14416 (N_14416,N_13924,N_14039);
xor U14417 (N_14417,N_14086,N_14323);
xnor U14418 (N_14418,N_14274,N_13929);
xnor U14419 (N_14419,N_14048,N_14228);
nand U14420 (N_14420,N_14332,N_14142);
nand U14421 (N_14421,N_13881,N_14138);
and U14422 (N_14422,N_14062,N_13975);
nor U14423 (N_14423,N_13803,N_13788);
or U14424 (N_14424,N_14134,N_14180);
xor U14425 (N_14425,N_14248,N_14207);
nor U14426 (N_14426,N_14037,N_13870);
or U14427 (N_14427,N_13770,N_14031);
nand U14428 (N_14428,N_13984,N_14087);
or U14429 (N_14429,N_14263,N_14362);
or U14430 (N_14430,N_13978,N_13830);
nor U14431 (N_14431,N_13977,N_13793);
nand U14432 (N_14432,N_14245,N_13807);
or U14433 (N_14433,N_14316,N_14367);
xor U14434 (N_14434,N_14139,N_14283);
or U14435 (N_14435,N_14164,N_13923);
and U14436 (N_14436,N_13899,N_14116);
xor U14437 (N_14437,N_14097,N_13778);
xor U14438 (N_14438,N_14311,N_13877);
nor U14439 (N_14439,N_13920,N_14102);
xnor U14440 (N_14440,N_14290,N_14050);
nor U14441 (N_14441,N_13753,N_14235);
and U14442 (N_14442,N_14158,N_14111);
and U14443 (N_14443,N_14336,N_13907);
nand U14444 (N_14444,N_13857,N_13851);
or U14445 (N_14445,N_14347,N_14145);
nand U14446 (N_14446,N_13852,N_13902);
xnor U14447 (N_14447,N_13875,N_14160);
and U14448 (N_14448,N_14232,N_13979);
nor U14449 (N_14449,N_14067,N_14029);
or U14450 (N_14450,N_14217,N_14124);
nand U14451 (N_14451,N_13750,N_13790);
nor U14452 (N_14452,N_14349,N_14227);
or U14453 (N_14453,N_14094,N_13860);
nand U14454 (N_14454,N_14103,N_13892);
and U14455 (N_14455,N_14154,N_13758);
or U14456 (N_14456,N_14231,N_14173);
nor U14457 (N_14457,N_14068,N_14135);
or U14458 (N_14458,N_13954,N_14038);
and U14459 (N_14459,N_13962,N_14112);
xnor U14460 (N_14460,N_14035,N_13964);
or U14461 (N_14461,N_13776,N_13782);
and U14462 (N_14462,N_14335,N_14358);
nor U14463 (N_14463,N_14253,N_14200);
and U14464 (N_14464,N_14309,N_13900);
nor U14465 (N_14465,N_13898,N_14306);
xor U14466 (N_14466,N_14076,N_13767);
nand U14467 (N_14467,N_13878,N_14299);
or U14468 (N_14468,N_14260,N_13812);
nor U14469 (N_14469,N_14148,N_14268);
and U14470 (N_14470,N_14012,N_14167);
and U14471 (N_14471,N_14045,N_14298);
or U14472 (N_14472,N_14113,N_13798);
xnor U14473 (N_14473,N_14132,N_14014);
nand U14474 (N_14474,N_14163,N_13944);
xnor U14475 (N_14475,N_13926,N_13890);
or U14476 (N_14476,N_13932,N_14205);
nand U14477 (N_14477,N_14292,N_14089);
nand U14478 (N_14478,N_14275,N_14190);
or U14479 (N_14479,N_14237,N_14100);
nand U14480 (N_14480,N_14373,N_14133);
nand U14481 (N_14481,N_14131,N_14247);
xnor U14482 (N_14482,N_13806,N_14310);
xor U14483 (N_14483,N_13916,N_14318);
xnor U14484 (N_14484,N_13912,N_13955);
nand U14485 (N_14485,N_13751,N_13950);
or U14486 (N_14486,N_14184,N_14325);
nand U14487 (N_14487,N_14301,N_13971);
and U14488 (N_14488,N_14120,N_14312);
and U14489 (N_14489,N_14288,N_14345);
xnor U14490 (N_14490,N_13969,N_14084);
or U14491 (N_14491,N_13905,N_14064);
nand U14492 (N_14492,N_13809,N_14078);
nand U14493 (N_14493,N_13949,N_14175);
and U14494 (N_14494,N_13840,N_13917);
and U14495 (N_14495,N_14223,N_14011);
nor U14496 (N_14496,N_14088,N_13886);
xnor U14497 (N_14497,N_13853,N_13822);
or U14498 (N_14498,N_14110,N_14250);
or U14499 (N_14499,N_13802,N_13831);
nor U14500 (N_14500,N_13835,N_14229);
or U14501 (N_14501,N_13894,N_14319);
nand U14502 (N_14502,N_14256,N_14077);
nand U14503 (N_14503,N_14010,N_13756);
and U14504 (N_14504,N_14042,N_14032);
nor U14505 (N_14505,N_14213,N_14215);
or U14506 (N_14506,N_14370,N_13828);
nand U14507 (N_14507,N_14289,N_13829);
and U14508 (N_14508,N_14313,N_14056);
nand U14509 (N_14509,N_14083,N_13862);
and U14510 (N_14510,N_13762,N_14206);
nor U14511 (N_14511,N_13826,N_14197);
and U14512 (N_14512,N_14143,N_13874);
nand U14513 (N_14513,N_13936,N_14172);
and U14514 (N_14514,N_14251,N_14331);
nand U14515 (N_14515,N_14041,N_13783);
and U14516 (N_14516,N_13771,N_14106);
xor U14517 (N_14517,N_14085,N_14308);
nor U14518 (N_14518,N_13827,N_13808);
or U14519 (N_14519,N_14337,N_13994);
and U14520 (N_14520,N_14182,N_14262);
and U14521 (N_14521,N_14198,N_13987);
nor U14522 (N_14522,N_13795,N_13972);
and U14523 (N_14523,N_14144,N_14202);
nor U14524 (N_14524,N_14125,N_14179);
xor U14525 (N_14525,N_14155,N_13847);
nand U14526 (N_14526,N_14277,N_14185);
nand U14527 (N_14527,N_14027,N_14241);
nand U14528 (N_14528,N_13887,N_13843);
and U14529 (N_14529,N_13786,N_14340);
xor U14530 (N_14530,N_14302,N_13910);
and U14531 (N_14531,N_13873,N_13904);
xnor U14532 (N_14532,N_14361,N_14019);
nor U14533 (N_14533,N_14270,N_14303);
or U14534 (N_14534,N_13991,N_14130);
or U14535 (N_14535,N_13925,N_14254);
nor U14536 (N_14536,N_13820,N_13946);
nand U14537 (N_14537,N_13844,N_14058);
or U14538 (N_14538,N_14304,N_14181);
nand U14539 (N_14539,N_13961,N_13911);
or U14540 (N_14540,N_13882,N_14147);
or U14541 (N_14541,N_14278,N_14051);
nor U14542 (N_14542,N_13866,N_13841);
xor U14543 (N_14543,N_14365,N_14296);
nand U14544 (N_14544,N_14249,N_14343);
xnor U14545 (N_14545,N_13985,N_13930);
and U14546 (N_14546,N_14141,N_14233);
xnor U14547 (N_14547,N_14327,N_13934);
or U14548 (N_14548,N_14267,N_14276);
nand U14549 (N_14549,N_13825,N_14069);
nand U14550 (N_14550,N_14236,N_14282);
or U14551 (N_14551,N_13811,N_14360);
and U14552 (N_14552,N_13872,N_14307);
and U14553 (N_14553,N_14259,N_14118);
xor U14554 (N_14554,N_14350,N_14280);
nand U14555 (N_14555,N_14122,N_14006);
or U14556 (N_14556,N_13931,N_14211);
nor U14557 (N_14557,N_14346,N_14161);
nor U14558 (N_14558,N_13974,N_13766);
nand U14559 (N_14559,N_14153,N_13837);
or U14560 (N_14560,N_13880,N_14040);
nand U14561 (N_14561,N_14072,N_13959);
and U14562 (N_14562,N_14242,N_14363);
nor U14563 (N_14563,N_14025,N_13965);
or U14564 (N_14564,N_14183,N_14000);
nor U14565 (N_14565,N_14091,N_14157);
nand U14566 (N_14566,N_13773,N_14057);
and U14567 (N_14567,N_14047,N_14090);
xnor U14568 (N_14568,N_13960,N_14008);
nand U14569 (N_14569,N_14364,N_14293);
xor U14570 (N_14570,N_13998,N_13858);
or U14571 (N_14571,N_13981,N_14060);
and U14572 (N_14572,N_13824,N_14328);
or U14573 (N_14573,N_14005,N_14352);
or U14574 (N_14574,N_14193,N_13915);
nand U14575 (N_14575,N_13792,N_13754);
xnor U14576 (N_14576,N_14151,N_14127);
and U14577 (N_14577,N_13993,N_14369);
nand U14578 (N_14578,N_14099,N_14003);
xor U14579 (N_14579,N_14082,N_13980);
nand U14580 (N_14580,N_13848,N_14300);
nand U14581 (N_14581,N_14009,N_13990);
xor U14582 (N_14582,N_13885,N_14126);
or U14583 (N_14583,N_13819,N_14114);
or U14584 (N_14584,N_14001,N_14152);
or U14585 (N_14585,N_13956,N_14265);
nand U14586 (N_14586,N_13787,N_13913);
nand U14587 (N_14587,N_14066,N_13769);
or U14588 (N_14588,N_14052,N_14214);
xnor U14589 (N_14589,N_14272,N_13893);
nor U14590 (N_14590,N_13856,N_14344);
xor U14591 (N_14591,N_14297,N_14156);
and U14592 (N_14592,N_14195,N_14353);
nand U14593 (N_14593,N_13953,N_14140);
or U14594 (N_14594,N_14257,N_14372);
or U14595 (N_14595,N_14013,N_13800);
xnor U14596 (N_14596,N_14357,N_14169);
xnor U14597 (N_14597,N_13884,N_13761);
and U14598 (N_14598,N_14053,N_14294);
and U14599 (N_14599,N_14188,N_14044);
nor U14600 (N_14600,N_13888,N_14326);
and U14601 (N_14601,N_13760,N_14121);
xnor U14602 (N_14602,N_13850,N_14287);
and U14603 (N_14603,N_14119,N_14004);
and U14604 (N_14604,N_13845,N_13976);
or U14605 (N_14605,N_13864,N_13967);
nor U14606 (N_14606,N_14176,N_14269);
and U14607 (N_14607,N_13988,N_13883);
xor U14608 (N_14608,N_14209,N_14178);
or U14609 (N_14609,N_14324,N_14150);
or U14610 (N_14610,N_14036,N_14273);
or U14611 (N_14611,N_13755,N_14238);
nor U14612 (N_14612,N_13801,N_14015);
nand U14613 (N_14613,N_14243,N_14049);
xor U14614 (N_14614,N_14117,N_14054);
nor U14615 (N_14615,N_14339,N_13903);
xor U14616 (N_14616,N_13818,N_13865);
xor U14617 (N_14617,N_14166,N_14244);
nor U14618 (N_14618,N_13759,N_14030);
xor U14619 (N_14619,N_13804,N_14320);
or U14620 (N_14620,N_14351,N_13935);
and U14621 (N_14621,N_14021,N_14258);
nand U14622 (N_14622,N_13810,N_14149);
xnor U14623 (N_14623,N_13966,N_13772);
nand U14624 (N_14624,N_14081,N_14196);
and U14625 (N_14625,N_13846,N_13999);
and U14626 (N_14626,N_13785,N_14170);
or U14627 (N_14627,N_14338,N_14359);
or U14628 (N_14628,N_14240,N_14317);
xnor U14629 (N_14629,N_13941,N_14330);
nor U14630 (N_14630,N_14023,N_14348);
or U14631 (N_14631,N_13832,N_13963);
and U14632 (N_14632,N_14007,N_14159);
xor U14633 (N_14633,N_13861,N_14168);
nand U14634 (N_14634,N_13871,N_14366);
xnor U14635 (N_14635,N_14024,N_14355);
or U14636 (N_14636,N_14221,N_13908);
xnor U14637 (N_14637,N_13997,N_14204);
xnor U14638 (N_14638,N_13863,N_13780);
nand U14639 (N_14639,N_14368,N_14177);
xor U14640 (N_14640,N_14234,N_14146);
xnor U14641 (N_14641,N_14208,N_13834);
and U14642 (N_14642,N_13895,N_13896);
nand U14643 (N_14643,N_13789,N_13869);
xnor U14644 (N_14644,N_13940,N_14174);
or U14645 (N_14645,N_14075,N_14128);
and U14646 (N_14646,N_13952,N_14186);
and U14647 (N_14647,N_13805,N_14291);
xor U14648 (N_14648,N_14104,N_13797);
nor U14649 (N_14649,N_13839,N_13855);
nand U14650 (N_14650,N_14187,N_13973);
or U14651 (N_14651,N_13815,N_14264);
and U14652 (N_14652,N_14322,N_13996);
nor U14653 (N_14653,N_14222,N_14374);
nand U14654 (N_14654,N_14079,N_14028);
xnor U14655 (N_14655,N_13784,N_13781);
nand U14656 (N_14656,N_14071,N_13814);
or U14657 (N_14657,N_14199,N_13842);
nor U14658 (N_14658,N_14020,N_13951);
xor U14659 (N_14659,N_14203,N_13937);
nand U14660 (N_14660,N_14092,N_14129);
and U14661 (N_14661,N_13943,N_14171);
xnor U14662 (N_14662,N_13757,N_14043);
nor U14663 (N_14663,N_13765,N_14034);
nor U14664 (N_14664,N_13945,N_13942);
xnor U14665 (N_14665,N_13970,N_14189);
nand U14666 (N_14666,N_14073,N_14212);
and U14667 (N_14667,N_13813,N_14281);
and U14668 (N_14668,N_14284,N_14315);
nand U14669 (N_14669,N_14246,N_13927);
or U14670 (N_14670,N_13763,N_14022);
or U14671 (N_14671,N_13889,N_13867);
and U14672 (N_14672,N_14239,N_14026);
nand U14673 (N_14673,N_14018,N_14218);
xor U14674 (N_14674,N_14219,N_13947);
nor U14675 (N_14675,N_13779,N_14201);
nor U14676 (N_14676,N_13995,N_14354);
nor U14677 (N_14677,N_14162,N_14107);
xnor U14678 (N_14678,N_13854,N_14165);
nand U14679 (N_14679,N_13919,N_13983);
nor U14680 (N_14680,N_13921,N_13817);
and U14681 (N_14681,N_13986,N_13958);
nor U14682 (N_14682,N_13992,N_14266);
and U14683 (N_14683,N_14295,N_13768);
and U14684 (N_14684,N_14371,N_14101);
xnor U14685 (N_14685,N_13775,N_14226);
nand U14686 (N_14686,N_13914,N_13928);
nor U14687 (N_14687,N_14059,N_13898);
xnor U14688 (N_14688,N_13832,N_14047);
nand U14689 (N_14689,N_13930,N_14137);
nor U14690 (N_14690,N_13966,N_14218);
and U14691 (N_14691,N_13858,N_13925);
nor U14692 (N_14692,N_14216,N_13953);
nor U14693 (N_14693,N_14286,N_14233);
and U14694 (N_14694,N_14126,N_13942);
or U14695 (N_14695,N_14035,N_13966);
nor U14696 (N_14696,N_13761,N_13893);
or U14697 (N_14697,N_14176,N_14060);
nor U14698 (N_14698,N_13934,N_14251);
or U14699 (N_14699,N_14222,N_13888);
or U14700 (N_14700,N_14313,N_14035);
or U14701 (N_14701,N_14344,N_14249);
xor U14702 (N_14702,N_13833,N_14300);
and U14703 (N_14703,N_14152,N_14084);
nand U14704 (N_14704,N_13916,N_14079);
xor U14705 (N_14705,N_13789,N_13932);
and U14706 (N_14706,N_14286,N_13940);
or U14707 (N_14707,N_13880,N_14223);
xor U14708 (N_14708,N_14224,N_13750);
or U14709 (N_14709,N_14218,N_14310);
nand U14710 (N_14710,N_14075,N_13996);
or U14711 (N_14711,N_14137,N_13834);
nand U14712 (N_14712,N_13817,N_13960);
nor U14713 (N_14713,N_13821,N_14368);
or U14714 (N_14714,N_13924,N_13878);
xnor U14715 (N_14715,N_14333,N_13973);
nand U14716 (N_14716,N_14127,N_13762);
xnor U14717 (N_14717,N_14260,N_14023);
or U14718 (N_14718,N_14300,N_14330);
or U14719 (N_14719,N_14081,N_14106);
nor U14720 (N_14720,N_14365,N_14336);
and U14721 (N_14721,N_13784,N_13881);
nand U14722 (N_14722,N_14343,N_13971);
and U14723 (N_14723,N_14064,N_13966);
and U14724 (N_14724,N_13973,N_13947);
and U14725 (N_14725,N_14329,N_13854);
xnor U14726 (N_14726,N_14038,N_14335);
or U14727 (N_14727,N_14083,N_14115);
nor U14728 (N_14728,N_13878,N_14349);
xor U14729 (N_14729,N_14351,N_14275);
and U14730 (N_14730,N_14127,N_14009);
nor U14731 (N_14731,N_14269,N_14085);
or U14732 (N_14732,N_14361,N_13969);
xor U14733 (N_14733,N_13769,N_14269);
nand U14734 (N_14734,N_13907,N_13776);
nor U14735 (N_14735,N_14016,N_14084);
or U14736 (N_14736,N_14215,N_13824);
and U14737 (N_14737,N_14157,N_13926);
nand U14738 (N_14738,N_13973,N_13949);
nor U14739 (N_14739,N_14132,N_13851);
xor U14740 (N_14740,N_14287,N_13978);
xor U14741 (N_14741,N_13843,N_14132);
nor U14742 (N_14742,N_13966,N_13904);
xor U14743 (N_14743,N_14042,N_14136);
or U14744 (N_14744,N_14035,N_14344);
and U14745 (N_14745,N_13833,N_13939);
nor U14746 (N_14746,N_14234,N_14160);
xor U14747 (N_14747,N_13986,N_13809);
xnor U14748 (N_14748,N_13837,N_14038);
and U14749 (N_14749,N_14332,N_13750);
xor U14750 (N_14750,N_13756,N_14197);
or U14751 (N_14751,N_14221,N_14044);
nor U14752 (N_14752,N_13920,N_13865);
xor U14753 (N_14753,N_13831,N_14198);
or U14754 (N_14754,N_14092,N_13908);
xnor U14755 (N_14755,N_14241,N_14213);
and U14756 (N_14756,N_13781,N_13763);
xnor U14757 (N_14757,N_14095,N_14016);
nand U14758 (N_14758,N_14362,N_14055);
nor U14759 (N_14759,N_14173,N_14351);
nor U14760 (N_14760,N_14091,N_14327);
or U14761 (N_14761,N_13919,N_13776);
nor U14762 (N_14762,N_13822,N_14237);
nand U14763 (N_14763,N_14067,N_14060);
or U14764 (N_14764,N_13923,N_14047);
xnor U14765 (N_14765,N_13899,N_14147);
xor U14766 (N_14766,N_13892,N_13993);
or U14767 (N_14767,N_14261,N_13996);
nand U14768 (N_14768,N_14038,N_14260);
or U14769 (N_14769,N_14091,N_14006);
and U14770 (N_14770,N_13966,N_13995);
nor U14771 (N_14771,N_14051,N_13923);
or U14772 (N_14772,N_14045,N_13754);
nand U14773 (N_14773,N_14148,N_14120);
and U14774 (N_14774,N_13980,N_13953);
or U14775 (N_14775,N_13902,N_13818);
nor U14776 (N_14776,N_14107,N_13869);
xnor U14777 (N_14777,N_13806,N_13944);
and U14778 (N_14778,N_14179,N_14083);
nand U14779 (N_14779,N_14120,N_13791);
nand U14780 (N_14780,N_14001,N_13802);
nand U14781 (N_14781,N_13861,N_14265);
xnor U14782 (N_14782,N_14227,N_14102);
or U14783 (N_14783,N_14056,N_14057);
nand U14784 (N_14784,N_13930,N_13857);
and U14785 (N_14785,N_14317,N_13887);
and U14786 (N_14786,N_14023,N_13832);
and U14787 (N_14787,N_14016,N_14080);
and U14788 (N_14788,N_14327,N_14215);
and U14789 (N_14789,N_14321,N_14350);
and U14790 (N_14790,N_14129,N_14226);
and U14791 (N_14791,N_14231,N_13955);
nand U14792 (N_14792,N_13874,N_14092);
and U14793 (N_14793,N_14349,N_14246);
nand U14794 (N_14794,N_13773,N_13755);
or U14795 (N_14795,N_14092,N_13997);
and U14796 (N_14796,N_14141,N_13800);
and U14797 (N_14797,N_13751,N_13780);
nand U14798 (N_14798,N_14321,N_14291);
nor U14799 (N_14799,N_14222,N_14187);
nor U14800 (N_14800,N_14218,N_13855);
and U14801 (N_14801,N_14361,N_14294);
and U14802 (N_14802,N_14264,N_14171);
and U14803 (N_14803,N_14293,N_14300);
xor U14804 (N_14804,N_14289,N_13920);
and U14805 (N_14805,N_13906,N_13792);
or U14806 (N_14806,N_14009,N_14090);
nand U14807 (N_14807,N_13945,N_13954);
and U14808 (N_14808,N_14310,N_14017);
nor U14809 (N_14809,N_14010,N_13912);
nor U14810 (N_14810,N_14010,N_13847);
or U14811 (N_14811,N_14056,N_14333);
nand U14812 (N_14812,N_13774,N_14049);
nor U14813 (N_14813,N_14124,N_14242);
nand U14814 (N_14814,N_13984,N_14107);
nand U14815 (N_14815,N_14026,N_14151);
xor U14816 (N_14816,N_14083,N_13956);
or U14817 (N_14817,N_14335,N_14295);
and U14818 (N_14818,N_14060,N_14025);
and U14819 (N_14819,N_14309,N_14167);
or U14820 (N_14820,N_13954,N_14082);
or U14821 (N_14821,N_14371,N_13929);
nand U14822 (N_14822,N_14056,N_13781);
and U14823 (N_14823,N_13959,N_13857);
and U14824 (N_14824,N_14358,N_14180);
xnor U14825 (N_14825,N_14303,N_13888);
or U14826 (N_14826,N_14088,N_13945);
xor U14827 (N_14827,N_14269,N_13921);
nor U14828 (N_14828,N_14076,N_14361);
or U14829 (N_14829,N_14342,N_13905);
and U14830 (N_14830,N_13897,N_14211);
xnor U14831 (N_14831,N_14331,N_14218);
nor U14832 (N_14832,N_13769,N_13781);
nand U14833 (N_14833,N_13839,N_14342);
or U14834 (N_14834,N_13979,N_13755);
and U14835 (N_14835,N_14337,N_13957);
and U14836 (N_14836,N_13764,N_14334);
and U14837 (N_14837,N_14158,N_14128);
and U14838 (N_14838,N_14008,N_14299);
nand U14839 (N_14839,N_14248,N_13994);
and U14840 (N_14840,N_13945,N_13768);
and U14841 (N_14841,N_14307,N_13825);
or U14842 (N_14842,N_14297,N_13849);
or U14843 (N_14843,N_14119,N_14211);
or U14844 (N_14844,N_14297,N_14057);
or U14845 (N_14845,N_14148,N_13814);
and U14846 (N_14846,N_14291,N_14205);
nor U14847 (N_14847,N_14137,N_14170);
or U14848 (N_14848,N_14351,N_14238);
or U14849 (N_14849,N_14209,N_13896);
nand U14850 (N_14850,N_13811,N_13921);
or U14851 (N_14851,N_14318,N_14115);
or U14852 (N_14852,N_14181,N_13921);
nand U14853 (N_14853,N_14198,N_14232);
nor U14854 (N_14854,N_13914,N_13766);
nand U14855 (N_14855,N_14339,N_14296);
nor U14856 (N_14856,N_14306,N_13842);
or U14857 (N_14857,N_13785,N_14336);
or U14858 (N_14858,N_14011,N_13831);
or U14859 (N_14859,N_14192,N_14223);
nor U14860 (N_14860,N_14319,N_14063);
nand U14861 (N_14861,N_13800,N_14190);
xnor U14862 (N_14862,N_13811,N_14126);
and U14863 (N_14863,N_14150,N_14047);
nand U14864 (N_14864,N_13858,N_14236);
nand U14865 (N_14865,N_14184,N_14164);
nand U14866 (N_14866,N_14164,N_13786);
xnor U14867 (N_14867,N_14054,N_14309);
nor U14868 (N_14868,N_14365,N_13800);
nor U14869 (N_14869,N_14263,N_14215);
nor U14870 (N_14870,N_14250,N_13872);
nor U14871 (N_14871,N_14006,N_14033);
nand U14872 (N_14872,N_14132,N_13954);
nand U14873 (N_14873,N_13753,N_14113);
or U14874 (N_14874,N_14348,N_14259);
or U14875 (N_14875,N_13897,N_14214);
nand U14876 (N_14876,N_13783,N_13961);
xor U14877 (N_14877,N_13926,N_13760);
or U14878 (N_14878,N_13863,N_14226);
nand U14879 (N_14879,N_14372,N_14340);
and U14880 (N_14880,N_14349,N_14313);
xnor U14881 (N_14881,N_13905,N_13948);
and U14882 (N_14882,N_13786,N_13921);
or U14883 (N_14883,N_14337,N_13896);
xnor U14884 (N_14884,N_14012,N_13974);
and U14885 (N_14885,N_14267,N_14091);
xor U14886 (N_14886,N_14059,N_14272);
or U14887 (N_14887,N_14233,N_14197);
or U14888 (N_14888,N_13939,N_14350);
or U14889 (N_14889,N_14207,N_14281);
or U14890 (N_14890,N_14024,N_14112);
and U14891 (N_14891,N_13860,N_13977);
or U14892 (N_14892,N_13828,N_13842);
or U14893 (N_14893,N_14143,N_13896);
nand U14894 (N_14894,N_13976,N_14328);
xnor U14895 (N_14895,N_14007,N_14138);
nand U14896 (N_14896,N_13815,N_14081);
xnor U14897 (N_14897,N_14203,N_13773);
nand U14898 (N_14898,N_14296,N_14127);
or U14899 (N_14899,N_13761,N_13891);
or U14900 (N_14900,N_13928,N_14254);
or U14901 (N_14901,N_14017,N_13935);
nand U14902 (N_14902,N_14206,N_13933);
xor U14903 (N_14903,N_14061,N_13923);
and U14904 (N_14904,N_14346,N_14171);
nand U14905 (N_14905,N_14188,N_14109);
nand U14906 (N_14906,N_13950,N_14253);
or U14907 (N_14907,N_14050,N_13987);
nor U14908 (N_14908,N_14045,N_14148);
and U14909 (N_14909,N_14166,N_14330);
nand U14910 (N_14910,N_14077,N_14350);
or U14911 (N_14911,N_14157,N_14272);
and U14912 (N_14912,N_13833,N_13830);
or U14913 (N_14913,N_14175,N_13990);
xnor U14914 (N_14914,N_14025,N_14167);
or U14915 (N_14915,N_13875,N_13941);
nor U14916 (N_14916,N_14320,N_13821);
nand U14917 (N_14917,N_14098,N_14192);
nor U14918 (N_14918,N_13895,N_14078);
xnor U14919 (N_14919,N_14282,N_14124);
or U14920 (N_14920,N_14048,N_13838);
and U14921 (N_14921,N_14139,N_14312);
nor U14922 (N_14922,N_14027,N_14348);
and U14923 (N_14923,N_14227,N_14104);
or U14924 (N_14924,N_14139,N_13897);
xnor U14925 (N_14925,N_14041,N_13931);
nand U14926 (N_14926,N_13972,N_14300);
or U14927 (N_14927,N_14193,N_14171);
or U14928 (N_14928,N_14076,N_13755);
xor U14929 (N_14929,N_14191,N_14078);
nand U14930 (N_14930,N_14110,N_14282);
and U14931 (N_14931,N_14039,N_13789);
or U14932 (N_14932,N_13775,N_13949);
xnor U14933 (N_14933,N_14110,N_14189);
nand U14934 (N_14934,N_14332,N_13835);
xnor U14935 (N_14935,N_13759,N_13906);
xnor U14936 (N_14936,N_14178,N_13759);
nand U14937 (N_14937,N_14166,N_14215);
nand U14938 (N_14938,N_14291,N_14209);
and U14939 (N_14939,N_14277,N_14176);
or U14940 (N_14940,N_14118,N_13866);
nand U14941 (N_14941,N_14174,N_14230);
or U14942 (N_14942,N_14043,N_14126);
xnor U14943 (N_14943,N_14062,N_13994);
nor U14944 (N_14944,N_14248,N_14349);
and U14945 (N_14945,N_13961,N_14258);
and U14946 (N_14946,N_14107,N_14269);
nand U14947 (N_14947,N_13814,N_14229);
xor U14948 (N_14948,N_13911,N_13879);
or U14949 (N_14949,N_14075,N_14032);
nor U14950 (N_14950,N_14125,N_13856);
or U14951 (N_14951,N_13991,N_14308);
and U14952 (N_14952,N_14289,N_14314);
xor U14953 (N_14953,N_14309,N_14229);
or U14954 (N_14954,N_13850,N_14064);
nand U14955 (N_14955,N_13796,N_14329);
nand U14956 (N_14956,N_13751,N_14122);
or U14957 (N_14957,N_13863,N_14075);
xor U14958 (N_14958,N_14286,N_14240);
xor U14959 (N_14959,N_14025,N_14087);
or U14960 (N_14960,N_14342,N_13855);
xnor U14961 (N_14961,N_14204,N_13920);
nor U14962 (N_14962,N_14244,N_13756);
nand U14963 (N_14963,N_14124,N_13784);
or U14964 (N_14964,N_14278,N_14057);
and U14965 (N_14965,N_14146,N_13866);
xor U14966 (N_14966,N_14021,N_14214);
and U14967 (N_14967,N_14334,N_13860);
nand U14968 (N_14968,N_13927,N_13998);
or U14969 (N_14969,N_13955,N_13881);
nor U14970 (N_14970,N_14244,N_14206);
xnor U14971 (N_14971,N_14091,N_13784);
nand U14972 (N_14972,N_14007,N_13801);
nor U14973 (N_14973,N_13868,N_14318);
nand U14974 (N_14974,N_14371,N_14073);
and U14975 (N_14975,N_14230,N_13939);
and U14976 (N_14976,N_14214,N_13847);
and U14977 (N_14977,N_13816,N_14039);
and U14978 (N_14978,N_14323,N_13768);
or U14979 (N_14979,N_13963,N_13792);
or U14980 (N_14980,N_13890,N_13891);
nor U14981 (N_14981,N_14114,N_14151);
nor U14982 (N_14982,N_13778,N_13795);
xor U14983 (N_14983,N_14143,N_13856);
xnor U14984 (N_14984,N_13763,N_14337);
and U14985 (N_14985,N_13885,N_13815);
nor U14986 (N_14986,N_14164,N_14185);
or U14987 (N_14987,N_14149,N_13878);
nor U14988 (N_14988,N_14282,N_13949);
nand U14989 (N_14989,N_13877,N_14254);
xor U14990 (N_14990,N_14240,N_13856);
and U14991 (N_14991,N_13884,N_14199);
nand U14992 (N_14992,N_14306,N_13784);
nor U14993 (N_14993,N_14040,N_13806);
or U14994 (N_14994,N_13794,N_13766);
nor U14995 (N_14995,N_14164,N_13965);
xnor U14996 (N_14996,N_14227,N_14295);
or U14997 (N_14997,N_14370,N_13837);
or U14998 (N_14998,N_13930,N_14206);
nor U14999 (N_14999,N_14240,N_13957);
xor U15000 (N_15000,N_14754,N_14879);
nand U15001 (N_15001,N_14761,N_14756);
xnor U15002 (N_15002,N_14418,N_14758);
xor U15003 (N_15003,N_14613,N_14741);
xor U15004 (N_15004,N_14672,N_14687);
nor U15005 (N_15005,N_14956,N_14597);
or U15006 (N_15006,N_14883,N_14710);
nor U15007 (N_15007,N_14656,N_14443);
or U15008 (N_15008,N_14950,N_14641);
nand U15009 (N_15009,N_14826,N_14383);
nor U15010 (N_15010,N_14704,N_14606);
nand U15011 (N_15011,N_14564,N_14622);
nor U15012 (N_15012,N_14457,N_14954);
or U15013 (N_15013,N_14814,N_14948);
nand U15014 (N_15014,N_14554,N_14744);
nand U15015 (N_15015,N_14655,N_14451);
and U15016 (N_15016,N_14771,N_14737);
nor U15017 (N_15017,N_14742,N_14893);
xnor U15018 (N_15018,N_14422,N_14843);
xor U15019 (N_15019,N_14612,N_14567);
and U15020 (N_15020,N_14963,N_14575);
or U15021 (N_15021,N_14726,N_14568);
nor U15022 (N_15022,N_14976,N_14671);
and U15023 (N_15023,N_14732,N_14524);
nor U15024 (N_15024,N_14553,N_14456);
nand U15025 (N_15025,N_14619,N_14962);
nor U15026 (N_15026,N_14694,N_14510);
xor U15027 (N_15027,N_14839,N_14856);
or U15028 (N_15028,N_14447,N_14590);
nand U15029 (N_15029,N_14495,N_14667);
xor U15030 (N_15030,N_14609,N_14511);
nor U15031 (N_15031,N_14435,N_14740);
nand U15032 (N_15032,N_14616,N_14965);
and U15033 (N_15033,N_14934,N_14611);
and U15034 (N_15034,N_14483,N_14604);
or U15035 (N_15035,N_14469,N_14503);
nor U15036 (N_15036,N_14395,N_14891);
or U15037 (N_15037,N_14413,N_14900);
and U15038 (N_15038,N_14561,N_14866);
xor U15039 (N_15039,N_14584,N_14514);
nor U15040 (N_15040,N_14804,N_14479);
xor U15041 (N_15041,N_14513,N_14907);
nand U15042 (N_15042,N_14781,N_14795);
and U15043 (N_15043,N_14541,N_14724);
nand U15044 (N_15044,N_14684,N_14995);
or U15045 (N_15045,N_14660,N_14802);
or U15046 (N_15046,N_14428,N_14733);
nor U15047 (N_15047,N_14708,N_14512);
nor U15048 (N_15048,N_14790,N_14788);
xor U15049 (N_15049,N_14381,N_14662);
or U15050 (N_15050,N_14565,N_14959);
or U15051 (N_15051,N_14916,N_14751);
nand U15052 (N_15052,N_14940,N_14657);
and U15053 (N_15053,N_14952,N_14625);
nand U15054 (N_15054,N_14621,N_14562);
nand U15055 (N_15055,N_14600,N_14643);
or U15056 (N_15056,N_14401,N_14496);
xnor U15057 (N_15057,N_14727,N_14847);
xor U15058 (N_15058,N_14881,N_14982);
or U15059 (N_15059,N_14407,N_14650);
nand U15060 (N_15060,N_14617,N_14777);
and U15061 (N_15061,N_14644,N_14887);
or U15062 (N_15062,N_14715,N_14983);
nor U15063 (N_15063,N_14698,N_14791);
or U15064 (N_15064,N_14391,N_14477);
nor U15065 (N_15065,N_14666,N_14505);
nor U15066 (N_15066,N_14515,N_14527);
nand U15067 (N_15067,N_14652,N_14996);
nand U15068 (N_15068,N_14593,N_14569);
or U15069 (N_15069,N_14803,N_14476);
or U15070 (N_15070,N_14844,N_14389);
xnor U15071 (N_15071,N_14624,N_14419);
or U15072 (N_15072,N_14416,N_14734);
and U15073 (N_15073,N_14425,N_14805);
nor U15074 (N_15074,N_14653,N_14836);
nor U15075 (N_15075,N_14472,N_14592);
or U15076 (N_15076,N_14819,N_14430);
and U15077 (N_15077,N_14988,N_14536);
nor U15078 (N_15078,N_14785,N_14432);
and U15079 (N_15079,N_14431,N_14608);
nor U15080 (N_15080,N_14542,N_14936);
nor U15081 (N_15081,N_14858,N_14471);
and U15082 (N_15082,N_14718,N_14961);
and U15083 (N_15083,N_14434,N_14668);
nand U15084 (N_15084,N_14522,N_14498);
or U15085 (N_15085,N_14500,N_14448);
xnor U15086 (N_15086,N_14830,N_14999);
nor U15087 (N_15087,N_14598,N_14967);
nor U15088 (N_15088,N_14827,N_14379);
nand U15089 (N_15089,N_14626,N_14499);
nor U15090 (N_15090,N_14701,N_14405);
nand U15091 (N_15091,N_14882,N_14922);
xnor U15092 (N_15092,N_14695,N_14378);
nand U15093 (N_15093,N_14974,N_14696);
and U15094 (N_15094,N_14441,N_14993);
and U15095 (N_15095,N_14601,N_14540);
nor U15096 (N_15096,N_14851,N_14556);
and U15097 (N_15097,N_14870,N_14411);
or U15098 (N_15098,N_14753,N_14945);
nor U15099 (N_15099,N_14423,N_14786);
xor U15100 (N_15100,N_14943,N_14829);
nand U15101 (N_15101,N_14571,N_14485);
nor U15102 (N_15102,N_14645,N_14837);
xnor U15103 (N_15103,N_14835,N_14816);
and U15104 (N_15104,N_14627,N_14989);
or U15105 (N_15105,N_14638,N_14923);
xnor U15106 (N_15106,N_14991,N_14482);
nor U15107 (N_15107,N_14973,N_14654);
nand U15108 (N_15108,N_14459,N_14525);
or U15109 (N_15109,N_14720,N_14426);
nand U15110 (N_15110,N_14594,N_14393);
xor U15111 (N_15111,N_14587,N_14550);
or U15112 (N_15112,N_14449,N_14583);
or U15113 (N_15113,N_14665,N_14917);
nor U15114 (N_15114,N_14581,N_14812);
nor U15115 (N_15115,N_14647,N_14534);
xor U15116 (N_15116,N_14926,N_14690);
and U15117 (N_15117,N_14857,N_14658);
xnor U15118 (N_15118,N_14840,N_14390);
and U15119 (N_15119,N_14800,N_14942);
xor U15120 (N_15120,N_14558,N_14927);
nand U15121 (N_15121,N_14719,N_14406);
nor U15122 (N_15122,N_14994,N_14670);
nand U15123 (N_15123,N_14530,N_14637);
and U15124 (N_15124,N_14886,N_14394);
nor U15125 (N_15125,N_14484,N_14639);
xor U15126 (N_15126,N_14822,N_14415);
nor U15127 (N_15127,N_14738,N_14605);
xnor U15128 (N_15128,N_14833,N_14576);
xnor U15129 (N_15129,N_14473,N_14507);
xnor U15130 (N_15130,N_14466,N_14478);
or U15131 (N_15131,N_14746,N_14453);
and U15132 (N_15132,N_14664,N_14966);
xor U15133 (N_15133,N_14642,N_14545);
nor U15134 (N_15134,N_14944,N_14424);
or U15135 (N_15135,N_14398,N_14725);
xor U15136 (N_15136,N_14997,N_14832);
nand U15137 (N_15137,N_14544,N_14560);
or U15138 (N_15138,N_14912,N_14508);
xor U15139 (N_15139,N_14504,N_14770);
xnor U15140 (N_15140,N_14794,N_14888);
or U15141 (N_15141,N_14410,N_14969);
xor U15142 (N_15142,N_14610,N_14980);
xor U15143 (N_15143,N_14949,N_14728);
nor U15144 (N_15144,N_14636,N_14535);
and U15145 (N_15145,N_14552,N_14585);
or U15146 (N_15146,N_14702,N_14489);
xnor U15147 (N_15147,N_14661,N_14528);
and U15148 (N_15148,N_14834,N_14905);
nand U15149 (N_15149,N_14382,N_14772);
xor U15150 (N_15150,N_14615,N_14409);
xor U15151 (N_15151,N_14686,N_14517);
xor U15152 (N_15152,N_14951,N_14890);
xnor U15153 (N_15153,N_14818,N_14436);
and U15154 (N_15154,N_14480,N_14981);
xor U15155 (N_15155,N_14501,N_14823);
xnor U15156 (N_15156,N_14909,N_14376);
or U15157 (N_15157,N_14978,N_14789);
nor U15158 (N_15158,N_14537,N_14828);
xor U15159 (N_15159,N_14439,N_14846);
or U15160 (N_15160,N_14730,N_14555);
xor U15161 (N_15161,N_14779,N_14502);
xnor U15162 (N_15162,N_14903,N_14745);
nor U15163 (N_15163,N_14864,N_14375);
nand U15164 (N_15164,N_14557,N_14723);
and U15165 (N_15165,N_14780,N_14572);
and U15166 (N_15166,N_14902,N_14885);
and U15167 (N_15167,N_14403,N_14855);
nor U15168 (N_15168,N_14955,N_14599);
and U15169 (N_15169,N_14607,N_14678);
nand U15170 (N_15170,N_14464,N_14938);
nor U15171 (N_15171,N_14468,N_14736);
and U15172 (N_15172,N_14752,N_14697);
nand U15173 (N_15173,N_14928,N_14768);
and U15174 (N_15174,N_14824,N_14404);
xor U15175 (N_15175,N_14747,N_14749);
nor U15176 (N_15176,N_14968,N_14918);
nand U15177 (N_15177,N_14578,N_14461);
and U15178 (N_15178,N_14769,N_14792);
xnor U15179 (N_15179,N_14591,N_14860);
xor U15180 (N_15180,N_14458,N_14573);
xor U15181 (N_15181,N_14586,N_14546);
nor U15182 (N_15182,N_14392,N_14631);
and U15183 (N_15183,N_14577,N_14596);
or U15184 (N_15184,N_14767,N_14801);
xnor U15185 (N_15185,N_14778,N_14445);
nand U15186 (N_15186,N_14825,N_14709);
nor U15187 (N_15187,N_14743,N_14990);
or U15188 (N_15188,N_14437,N_14632);
nor U15189 (N_15189,N_14813,N_14659);
nor U15190 (N_15190,N_14623,N_14915);
and U15191 (N_15191,N_14739,N_14529);
and U15192 (N_15192,N_14821,N_14531);
and U15193 (N_15193,N_14614,N_14396);
nand U15194 (N_15194,N_14998,N_14676);
nor U15195 (N_15195,N_14486,N_14925);
nand U15196 (N_15196,N_14589,N_14474);
nor U15197 (N_15197,N_14455,N_14603);
or U15198 (N_15198,N_14979,N_14904);
or U15199 (N_15199,N_14845,N_14475);
or U15200 (N_15200,N_14932,N_14452);
nor U15201 (N_15201,N_14811,N_14675);
nand U15202 (N_15202,N_14869,N_14992);
xor U15203 (N_15203,N_14493,N_14681);
nand U15204 (N_15204,N_14892,N_14692);
or U15205 (N_15205,N_14871,N_14735);
nor U15206 (N_15206,N_14729,N_14651);
nor U15207 (N_15207,N_14387,N_14438);
xor U15208 (N_15208,N_14539,N_14633);
nor U15209 (N_15209,N_14798,N_14750);
or U15210 (N_15210,N_14958,N_14731);
nor U15211 (N_15211,N_14763,N_14721);
and U15212 (N_15212,N_14532,N_14908);
and U15213 (N_15213,N_14931,N_14850);
and U15214 (N_15214,N_14933,N_14852);
and U15215 (N_15215,N_14526,N_14463);
and U15216 (N_15216,N_14516,N_14783);
nor U15217 (N_15217,N_14875,N_14867);
nand U15218 (N_15218,N_14716,N_14865);
xnor U15219 (N_15219,N_14972,N_14714);
nand U15220 (N_15220,N_14674,N_14700);
xnor U15221 (N_15221,N_14450,N_14548);
nor U15222 (N_15222,N_14899,N_14774);
xor U15223 (N_15223,N_14929,N_14838);
and U15224 (N_15224,N_14854,N_14760);
or U15225 (N_15225,N_14682,N_14914);
nor U15226 (N_15226,N_14699,N_14635);
nand U15227 (N_15227,N_14853,N_14467);
nand U15228 (N_15228,N_14859,N_14685);
xor U15229 (N_15229,N_14683,N_14971);
or U15230 (N_15230,N_14941,N_14764);
xnor U15231 (N_15231,N_14399,N_14533);
nor U15232 (N_15232,N_14796,N_14759);
nor U15233 (N_15233,N_14487,N_14566);
nand U15234 (N_15234,N_14970,N_14820);
xnor U15235 (N_15235,N_14693,N_14519);
or U15236 (N_15236,N_14784,N_14717);
nand U15237 (N_15237,N_14986,N_14862);
xor U15238 (N_15238,N_14861,N_14397);
and U15239 (N_15239,N_14388,N_14549);
or U15240 (N_15240,N_14620,N_14547);
nand U15241 (N_15241,N_14712,N_14806);
or U15242 (N_15242,N_14629,N_14414);
and U15243 (N_15243,N_14648,N_14679);
or U15244 (N_15244,N_14618,N_14628);
nand U15245 (N_15245,N_14874,N_14582);
and U15246 (N_15246,N_14680,N_14446);
nor U15247 (N_15247,N_14570,N_14543);
or U15248 (N_15248,N_14497,N_14402);
nor U15249 (N_15249,N_14490,N_14521);
nor U15250 (N_15250,N_14946,N_14462);
xor U15251 (N_15251,N_14831,N_14776);
or U15252 (N_15252,N_14960,N_14444);
nor U15253 (N_15253,N_14884,N_14574);
or U15254 (N_15254,N_14848,N_14705);
and U15255 (N_15255,N_14787,N_14509);
nand U15256 (N_15256,N_14649,N_14677);
or U15257 (N_15257,N_14817,N_14880);
or U15258 (N_15258,N_14876,N_14460);
nand U15259 (N_15259,N_14377,N_14551);
xnor U15260 (N_15260,N_14957,N_14722);
xor U15261 (N_15261,N_14663,N_14935);
nand U15262 (N_15262,N_14877,N_14580);
and U15263 (N_15263,N_14559,N_14384);
or U15264 (N_15264,N_14913,N_14984);
nand U15265 (N_15265,N_14470,N_14762);
nand U15266 (N_15266,N_14689,N_14906);
nand U15267 (N_15267,N_14815,N_14757);
or U15268 (N_15268,N_14793,N_14894);
nand U15269 (N_15269,N_14454,N_14417);
nor U15270 (N_15270,N_14868,N_14440);
and U15271 (N_15271,N_14939,N_14380);
or U15272 (N_15272,N_14506,N_14579);
or U15273 (N_15273,N_14773,N_14412);
nand U15274 (N_15274,N_14385,N_14518);
nor U15275 (N_15275,N_14588,N_14429);
xor U15276 (N_15276,N_14707,N_14889);
and U15277 (N_15277,N_14520,N_14433);
nor U15278 (N_15278,N_14713,N_14523);
or U15279 (N_15279,N_14673,N_14987);
or U15280 (N_15280,N_14841,N_14634);
nand U15281 (N_15281,N_14895,N_14873);
nand U15282 (N_15282,N_14897,N_14386);
or U15283 (N_15283,N_14863,N_14400);
nor U15284 (N_15284,N_14538,N_14494);
or U15285 (N_15285,N_14782,N_14809);
nand U15286 (N_15286,N_14755,N_14492);
xor U15287 (N_15287,N_14878,N_14849);
or U15288 (N_15288,N_14977,N_14691);
nor U15289 (N_15289,N_14810,N_14765);
nand U15290 (N_15290,N_14703,N_14901);
xnor U15291 (N_15291,N_14898,N_14442);
nor U15292 (N_15292,N_14937,N_14930);
xnor U15293 (N_15293,N_14920,N_14910);
xor U15294 (N_15294,N_14872,N_14640);
xnor U15295 (N_15295,N_14985,N_14964);
or U15296 (N_15296,N_14706,N_14896);
nor U15297 (N_15297,N_14921,N_14427);
and U15298 (N_15298,N_14491,N_14711);
nand U15299 (N_15299,N_14688,N_14797);
nor U15300 (N_15300,N_14924,N_14465);
nor U15301 (N_15301,N_14842,N_14488);
nor U15302 (N_15302,N_14911,N_14630);
xnor U15303 (N_15303,N_14602,N_14775);
nand U15304 (N_15304,N_14947,N_14481);
nor U15305 (N_15305,N_14766,N_14807);
xnor U15306 (N_15306,N_14975,N_14646);
and U15307 (N_15307,N_14953,N_14919);
xor U15308 (N_15308,N_14669,N_14595);
and U15309 (N_15309,N_14421,N_14799);
xnor U15310 (N_15310,N_14420,N_14748);
and U15311 (N_15311,N_14408,N_14563);
nor U15312 (N_15312,N_14808,N_14403);
nand U15313 (N_15313,N_14575,N_14669);
xor U15314 (N_15314,N_14906,N_14889);
or U15315 (N_15315,N_14604,N_14678);
and U15316 (N_15316,N_14398,N_14796);
or U15317 (N_15317,N_14937,N_14940);
nand U15318 (N_15318,N_14412,N_14703);
nand U15319 (N_15319,N_14453,N_14931);
and U15320 (N_15320,N_14449,N_14751);
nor U15321 (N_15321,N_14485,N_14760);
or U15322 (N_15322,N_14582,N_14774);
nand U15323 (N_15323,N_14815,N_14396);
nor U15324 (N_15324,N_14757,N_14905);
or U15325 (N_15325,N_14516,N_14562);
and U15326 (N_15326,N_14791,N_14968);
xor U15327 (N_15327,N_14547,N_14473);
xnor U15328 (N_15328,N_14821,N_14936);
or U15329 (N_15329,N_14853,N_14465);
and U15330 (N_15330,N_14957,N_14615);
or U15331 (N_15331,N_14863,N_14403);
nor U15332 (N_15332,N_14545,N_14822);
or U15333 (N_15333,N_14804,N_14699);
and U15334 (N_15334,N_14780,N_14805);
and U15335 (N_15335,N_14961,N_14483);
nand U15336 (N_15336,N_14617,N_14922);
nand U15337 (N_15337,N_14601,N_14991);
nor U15338 (N_15338,N_14892,N_14842);
or U15339 (N_15339,N_14556,N_14764);
xor U15340 (N_15340,N_14706,N_14508);
xor U15341 (N_15341,N_14444,N_14515);
and U15342 (N_15342,N_14552,N_14638);
xor U15343 (N_15343,N_14664,N_14456);
or U15344 (N_15344,N_14538,N_14696);
xnor U15345 (N_15345,N_14577,N_14450);
nor U15346 (N_15346,N_14472,N_14932);
and U15347 (N_15347,N_14732,N_14644);
nand U15348 (N_15348,N_14546,N_14527);
nor U15349 (N_15349,N_14906,N_14965);
xnor U15350 (N_15350,N_14470,N_14728);
nand U15351 (N_15351,N_14879,N_14606);
nand U15352 (N_15352,N_14395,N_14775);
nor U15353 (N_15353,N_14479,N_14739);
nand U15354 (N_15354,N_14775,N_14578);
or U15355 (N_15355,N_14811,N_14455);
or U15356 (N_15356,N_14646,N_14515);
nor U15357 (N_15357,N_14766,N_14581);
or U15358 (N_15358,N_14818,N_14733);
nand U15359 (N_15359,N_14876,N_14407);
nand U15360 (N_15360,N_14703,N_14759);
and U15361 (N_15361,N_14972,N_14526);
or U15362 (N_15362,N_14987,N_14649);
nand U15363 (N_15363,N_14428,N_14656);
nand U15364 (N_15364,N_14766,N_14926);
or U15365 (N_15365,N_14927,N_14530);
nor U15366 (N_15366,N_14530,N_14730);
and U15367 (N_15367,N_14904,N_14397);
nand U15368 (N_15368,N_14722,N_14386);
or U15369 (N_15369,N_14703,N_14777);
or U15370 (N_15370,N_14946,N_14459);
xnor U15371 (N_15371,N_14482,N_14820);
nand U15372 (N_15372,N_14692,N_14961);
and U15373 (N_15373,N_14602,N_14556);
and U15374 (N_15374,N_14940,N_14562);
nor U15375 (N_15375,N_14746,N_14415);
or U15376 (N_15376,N_14978,N_14516);
nor U15377 (N_15377,N_14434,N_14980);
and U15378 (N_15378,N_14691,N_14874);
nor U15379 (N_15379,N_14695,N_14986);
nand U15380 (N_15380,N_14547,N_14833);
nand U15381 (N_15381,N_14977,N_14557);
and U15382 (N_15382,N_14565,N_14806);
nand U15383 (N_15383,N_14785,N_14520);
nand U15384 (N_15384,N_14508,N_14517);
nand U15385 (N_15385,N_14512,N_14481);
nand U15386 (N_15386,N_14495,N_14447);
and U15387 (N_15387,N_14491,N_14872);
nor U15388 (N_15388,N_14419,N_14716);
nor U15389 (N_15389,N_14767,N_14449);
nor U15390 (N_15390,N_14527,N_14419);
or U15391 (N_15391,N_14674,N_14978);
nand U15392 (N_15392,N_14462,N_14576);
xor U15393 (N_15393,N_14737,N_14545);
xor U15394 (N_15394,N_14766,N_14674);
nand U15395 (N_15395,N_14989,N_14829);
and U15396 (N_15396,N_14581,N_14920);
xnor U15397 (N_15397,N_14552,N_14635);
xnor U15398 (N_15398,N_14735,N_14625);
or U15399 (N_15399,N_14579,N_14520);
xnor U15400 (N_15400,N_14845,N_14600);
and U15401 (N_15401,N_14861,N_14561);
nand U15402 (N_15402,N_14533,N_14549);
nor U15403 (N_15403,N_14501,N_14691);
or U15404 (N_15404,N_14401,N_14893);
xnor U15405 (N_15405,N_14705,N_14746);
xnor U15406 (N_15406,N_14745,N_14918);
and U15407 (N_15407,N_14804,N_14694);
nor U15408 (N_15408,N_14767,N_14752);
or U15409 (N_15409,N_14383,N_14773);
or U15410 (N_15410,N_14543,N_14911);
and U15411 (N_15411,N_14435,N_14977);
xor U15412 (N_15412,N_14991,N_14731);
nand U15413 (N_15413,N_14399,N_14952);
nand U15414 (N_15414,N_14592,N_14636);
xnor U15415 (N_15415,N_14444,N_14824);
and U15416 (N_15416,N_14444,N_14919);
and U15417 (N_15417,N_14796,N_14858);
xor U15418 (N_15418,N_14464,N_14892);
nor U15419 (N_15419,N_14820,N_14728);
nor U15420 (N_15420,N_14839,N_14432);
xor U15421 (N_15421,N_14663,N_14775);
xnor U15422 (N_15422,N_14432,N_14712);
xnor U15423 (N_15423,N_14804,N_14508);
nand U15424 (N_15424,N_14763,N_14480);
xor U15425 (N_15425,N_14636,N_14580);
or U15426 (N_15426,N_14804,N_14790);
and U15427 (N_15427,N_14471,N_14678);
nand U15428 (N_15428,N_14941,N_14401);
xor U15429 (N_15429,N_14816,N_14880);
or U15430 (N_15430,N_14643,N_14739);
or U15431 (N_15431,N_14961,N_14496);
or U15432 (N_15432,N_14684,N_14500);
nor U15433 (N_15433,N_14803,N_14865);
nand U15434 (N_15434,N_14882,N_14738);
nor U15435 (N_15435,N_14789,N_14753);
or U15436 (N_15436,N_14838,N_14502);
or U15437 (N_15437,N_14709,N_14962);
xor U15438 (N_15438,N_14908,N_14491);
and U15439 (N_15439,N_14590,N_14888);
nor U15440 (N_15440,N_14681,N_14879);
or U15441 (N_15441,N_14903,N_14376);
nor U15442 (N_15442,N_14673,N_14455);
xor U15443 (N_15443,N_14481,N_14957);
xor U15444 (N_15444,N_14649,N_14936);
xor U15445 (N_15445,N_14491,N_14564);
or U15446 (N_15446,N_14918,N_14843);
or U15447 (N_15447,N_14477,N_14613);
nor U15448 (N_15448,N_14878,N_14696);
nand U15449 (N_15449,N_14657,N_14447);
and U15450 (N_15450,N_14756,N_14683);
nand U15451 (N_15451,N_14527,N_14785);
nor U15452 (N_15452,N_14960,N_14379);
xnor U15453 (N_15453,N_14789,N_14567);
nor U15454 (N_15454,N_14474,N_14681);
nand U15455 (N_15455,N_14546,N_14791);
nand U15456 (N_15456,N_14939,N_14648);
xnor U15457 (N_15457,N_14643,N_14557);
nor U15458 (N_15458,N_14515,N_14947);
xor U15459 (N_15459,N_14775,N_14951);
nor U15460 (N_15460,N_14776,N_14445);
nand U15461 (N_15461,N_14861,N_14699);
and U15462 (N_15462,N_14421,N_14604);
nand U15463 (N_15463,N_14539,N_14807);
or U15464 (N_15464,N_14923,N_14490);
or U15465 (N_15465,N_14712,N_14639);
nor U15466 (N_15466,N_14454,N_14984);
xor U15467 (N_15467,N_14855,N_14630);
xor U15468 (N_15468,N_14552,N_14914);
or U15469 (N_15469,N_14518,N_14640);
or U15470 (N_15470,N_14747,N_14861);
or U15471 (N_15471,N_14986,N_14953);
xnor U15472 (N_15472,N_14712,N_14701);
xor U15473 (N_15473,N_14569,N_14408);
nor U15474 (N_15474,N_14659,N_14447);
nor U15475 (N_15475,N_14918,N_14672);
and U15476 (N_15476,N_14871,N_14705);
and U15477 (N_15477,N_14723,N_14753);
nor U15478 (N_15478,N_14450,N_14864);
and U15479 (N_15479,N_14636,N_14694);
nand U15480 (N_15480,N_14412,N_14829);
and U15481 (N_15481,N_14804,N_14613);
xnor U15482 (N_15482,N_14463,N_14778);
or U15483 (N_15483,N_14803,N_14809);
nor U15484 (N_15484,N_14951,N_14828);
nand U15485 (N_15485,N_14868,N_14446);
nand U15486 (N_15486,N_14764,N_14754);
nor U15487 (N_15487,N_14492,N_14811);
nand U15488 (N_15488,N_14607,N_14758);
or U15489 (N_15489,N_14573,N_14788);
xnor U15490 (N_15490,N_14643,N_14444);
nor U15491 (N_15491,N_14963,N_14908);
nand U15492 (N_15492,N_14622,N_14810);
and U15493 (N_15493,N_14683,N_14554);
and U15494 (N_15494,N_14454,N_14712);
nand U15495 (N_15495,N_14941,N_14741);
nand U15496 (N_15496,N_14802,N_14969);
and U15497 (N_15497,N_14634,N_14402);
nand U15498 (N_15498,N_14378,N_14876);
nor U15499 (N_15499,N_14682,N_14977);
and U15500 (N_15500,N_14909,N_14936);
nor U15501 (N_15501,N_14841,N_14568);
nor U15502 (N_15502,N_14610,N_14915);
or U15503 (N_15503,N_14975,N_14833);
or U15504 (N_15504,N_14646,N_14720);
and U15505 (N_15505,N_14944,N_14652);
or U15506 (N_15506,N_14785,N_14996);
and U15507 (N_15507,N_14766,N_14618);
and U15508 (N_15508,N_14722,N_14440);
nor U15509 (N_15509,N_14924,N_14792);
nand U15510 (N_15510,N_14405,N_14821);
nor U15511 (N_15511,N_14437,N_14540);
nand U15512 (N_15512,N_14958,N_14475);
xor U15513 (N_15513,N_14549,N_14981);
nand U15514 (N_15514,N_14934,N_14509);
xor U15515 (N_15515,N_14443,N_14516);
xnor U15516 (N_15516,N_14765,N_14523);
xor U15517 (N_15517,N_14646,N_14900);
nor U15518 (N_15518,N_14629,N_14586);
nor U15519 (N_15519,N_14972,N_14922);
or U15520 (N_15520,N_14502,N_14393);
xor U15521 (N_15521,N_14423,N_14984);
or U15522 (N_15522,N_14416,N_14772);
xor U15523 (N_15523,N_14703,N_14812);
and U15524 (N_15524,N_14410,N_14981);
and U15525 (N_15525,N_14848,N_14854);
and U15526 (N_15526,N_14903,N_14521);
or U15527 (N_15527,N_14520,N_14875);
nand U15528 (N_15528,N_14608,N_14392);
nor U15529 (N_15529,N_14406,N_14522);
nor U15530 (N_15530,N_14480,N_14650);
xor U15531 (N_15531,N_14625,N_14763);
or U15532 (N_15532,N_14566,N_14893);
or U15533 (N_15533,N_14471,N_14550);
or U15534 (N_15534,N_14470,N_14765);
xor U15535 (N_15535,N_14734,N_14414);
nor U15536 (N_15536,N_14736,N_14599);
nor U15537 (N_15537,N_14910,N_14437);
xnor U15538 (N_15538,N_14702,N_14950);
and U15539 (N_15539,N_14739,N_14547);
xor U15540 (N_15540,N_14862,N_14849);
nor U15541 (N_15541,N_14831,N_14984);
and U15542 (N_15542,N_14457,N_14507);
xnor U15543 (N_15543,N_14854,N_14920);
or U15544 (N_15544,N_14608,N_14558);
nor U15545 (N_15545,N_14583,N_14523);
nand U15546 (N_15546,N_14799,N_14906);
or U15547 (N_15547,N_14909,N_14590);
xor U15548 (N_15548,N_14642,N_14946);
xor U15549 (N_15549,N_14530,N_14549);
and U15550 (N_15550,N_14452,N_14789);
nand U15551 (N_15551,N_14660,N_14456);
or U15552 (N_15552,N_14632,N_14641);
nand U15553 (N_15553,N_14519,N_14383);
xor U15554 (N_15554,N_14928,N_14953);
xor U15555 (N_15555,N_14816,N_14488);
or U15556 (N_15556,N_14395,N_14485);
or U15557 (N_15557,N_14739,N_14597);
or U15558 (N_15558,N_14659,N_14734);
or U15559 (N_15559,N_14645,N_14868);
nand U15560 (N_15560,N_14740,N_14960);
nor U15561 (N_15561,N_14568,N_14627);
xor U15562 (N_15562,N_14717,N_14929);
nand U15563 (N_15563,N_14937,N_14945);
or U15564 (N_15564,N_14872,N_14545);
or U15565 (N_15565,N_14878,N_14692);
and U15566 (N_15566,N_14388,N_14712);
nand U15567 (N_15567,N_14554,N_14821);
or U15568 (N_15568,N_14798,N_14643);
or U15569 (N_15569,N_14890,N_14557);
or U15570 (N_15570,N_14517,N_14506);
xnor U15571 (N_15571,N_14960,N_14412);
or U15572 (N_15572,N_14698,N_14433);
and U15573 (N_15573,N_14805,N_14813);
xor U15574 (N_15574,N_14638,N_14626);
nand U15575 (N_15575,N_14415,N_14933);
xnor U15576 (N_15576,N_14559,N_14865);
nand U15577 (N_15577,N_14810,N_14758);
nor U15578 (N_15578,N_14967,N_14495);
xor U15579 (N_15579,N_14879,N_14705);
or U15580 (N_15580,N_14573,N_14963);
nor U15581 (N_15581,N_14490,N_14869);
nor U15582 (N_15582,N_14419,N_14393);
nor U15583 (N_15583,N_14463,N_14921);
xor U15584 (N_15584,N_14834,N_14407);
and U15585 (N_15585,N_14510,N_14979);
xnor U15586 (N_15586,N_14904,N_14474);
xnor U15587 (N_15587,N_14860,N_14953);
nand U15588 (N_15588,N_14811,N_14505);
xnor U15589 (N_15589,N_14539,N_14696);
or U15590 (N_15590,N_14557,N_14883);
xor U15591 (N_15591,N_14944,N_14798);
nand U15592 (N_15592,N_14984,N_14493);
xor U15593 (N_15593,N_14997,N_14549);
xnor U15594 (N_15594,N_14549,N_14675);
nand U15595 (N_15595,N_14435,N_14841);
nand U15596 (N_15596,N_14921,N_14941);
nor U15597 (N_15597,N_14490,N_14932);
nor U15598 (N_15598,N_14657,N_14547);
nand U15599 (N_15599,N_14556,N_14511);
or U15600 (N_15600,N_14509,N_14552);
nor U15601 (N_15601,N_14700,N_14772);
nor U15602 (N_15602,N_14663,N_14898);
nor U15603 (N_15603,N_14504,N_14718);
and U15604 (N_15604,N_14555,N_14868);
and U15605 (N_15605,N_14593,N_14937);
or U15606 (N_15606,N_14641,N_14603);
and U15607 (N_15607,N_14861,N_14698);
nor U15608 (N_15608,N_14909,N_14828);
nor U15609 (N_15609,N_14575,N_14629);
nand U15610 (N_15610,N_14821,N_14998);
or U15611 (N_15611,N_14634,N_14471);
xor U15612 (N_15612,N_14602,N_14534);
xnor U15613 (N_15613,N_14662,N_14478);
or U15614 (N_15614,N_14376,N_14928);
or U15615 (N_15615,N_14683,N_14973);
and U15616 (N_15616,N_14907,N_14773);
xnor U15617 (N_15617,N_14504,N_14494);
nor U15618 (N_15618,N_14382,N_14542);
nand U15619 (N_15619,N_14432,N_14535);
nand U15620 (N_15620,N_14457,N_14875);
nand U15621 (N_15621,N_14969,N_14665);
nand U15622 (N_15622,N_14555,N_14778);
or U15623 (N_15623,N_14641,N_14697);
or U15624 (N_15624,N_14756,N_14744);
nand U15625 (N_15625,N_15372,N_15303);
xor U15626 (N_15626,N_15555,N_15212);
nor U15627 (N_15627,N_15005,N_15050);
or U15628 (N_15628,N_15165,N_15217);
and U15629 (N_15629,N_15047,N_15409);
nor U15630 (N_15630,N_15166,N_15490);
xnor U15631 (N_15631,N_15171,N_15355);
or U15632 (N_15632,N_15525,N_15234);
nand U15633 (N_15633,N_15444,N_15553);
nand U15634 (N_15634,N_15317,N_15346);
and U15635 (N_15635,N_15397,N_15055);
and U15636 (N_15636,N_15455,N_15602);
and U15637 (N_15637,N_15264,N_15144);
nand U15638 (N_15638,N_15349,N_15118);
nand U15639 (N_15639,N_15445,N_15468);
nor U15640 (N_15640,N_15247,N_15186);
nor U15641 (N_15641,N_15597,N_15147);
or U15642 (N_15642,N_15379,N_15156);
and U15643 (N_15643,N_15466,N_15133);
nor U15644 (N_15644,N_15495,N_15266);
and U15645 (N_15645,N_15319,N_15290);
nand U15646 (N_15646,N_15322,N_15457);
or U15647 (N_15647,N_15185,N_15188);
or U15648 (N_15648,N_15439,N_15369);
nand U15649 (N_15649,N_15207,N_15310);
nand U15650 (N_15650,N_15599,N_15391);
xnor U15651 (N_15651,N_15568,N_15586);
or U15652 (N_15652,N_15235,N_15281);
and U15653 (N_15653,N_15014,N_15128);
nand U15654 (N_15654,N_15110,N_15620);
xor U15655 (N_15655,N_15535,N_15549);
xnor U15656 (N_15656,N_15079,N_15243);
xnor U15657 (N_15657,N_15565,N_15563);
xnor U15658 (N_15658,N_15526,N_15167);
and U15659 (N_15659,N_15263,N_15226);
xnor U15660 (N_15660,N_15280,N_15206);
or U15661 (N_15661,N_15363,N_15410);
and U15662 (N_15662,N_15276,N_15508);
nand U15663 (N_15663,N_15371,N_15056);
xor U15664 (N_15664,N_15403,N_15145);
and U15665 (N_15665,N_15275,N_15010);
xor U15666 (N_15666,N_15125,N_15245);
and U15667 (N_15667,N_15170,N_15139);
and U15668 (N_15668,N_15137,N_15127);
and U15669 (N_15669,N_15399,N_15378);
and U15670 (N_15670,N_15447,N_15540);
xnor U15671 (N_15671,N_15499,N_15215);
and U15672 (N_15672,N_15108,N_15130);
or U15673 (N_15673,N_15046,N_15161);
nor U15674 (N_15674,N_15590,N_15094);
and U15675 (N_15675,N_15509,N_15283);
xnor U15676 (N_15676,N_15614,N_15175);
xor U15677 (N_15677,N_15465,N_15313);
nor U15678 (N_15678,N_15566,N_15204);
nor U15679 (N_15679,N_15438,N_15429);
nor U15680 (N_15680,N_15442,N_15287);
and U15681 (N_15681,N_15398,N_15343);
or U15682 (N_15682,N_15311,N_15520);
and U15683 (N_15683,N_15591,N_15471);
or U15684 (N_15684,N_15558,N_15262);
and U15685 (N_15685,N_15102,N_15511);
and U15686 (N_15686,N_15123,N_15277);
xor U15687 (N_15687,N_15446,N_15009);
nand U15688 (N_15688,N_15463,N_15416);
or U15689 (N_15689,N_15464,N_15522);
xor U15690 (N_15690,N_15023,N_15286);
nor U15691 (N_15691,N_15220,N_15202);
nand U15692 (N_15692,N_15260,N_15358);
and U15693 (N_15693,N_15273,N_15049);
xor U15694 (N_15694,N_15306,N_15577);
or U15695 (N_15695,N_15299,N_15103);
nor U15696 (N_15696,N_15270,N_15381);
nand U15697 (N_15697,N_15078,N_15539);
or U15698 (N_15698,N_15435,N_15300);
or U15699 (N_15699,N_15564,N_15594);
or U15700 (N_15700,N_15489,N_15459);
nand U15701 (N_15701,N_15155,N_15182);
nand U15702 (N_15702,N_15084,N_15451);
nor U15703 (N_15703,N_15026,N_15148);
nand U15704 (N_15704,N_15031,N_15183);
nor U15705 (N_15705,N_15248,N_15475);
and U15706 (N_15706,N_15037,N_15480);
nand U15707 (N_15707,N_15562,N_15146);
and U15708 (N_15708,N_15058,N_15592);
and U15709 (N_15709,N_15282,N_15051);
nor U15710 (N_15710,N_15087,N_15428);
nand U15711 (N_15711,N_15241,N_15407);
nand U15712 (N_15712,N_15353,N_15033);
or U15713 (N_15713,N_15417,N_15066);
xor U15714 (N_15714,N_15570,N_15261);
nand U15715 (N_15715,N_15007,N_15593);
or U15716 (N_15716,N_15140,N_15232);
and U15717 (N_15717,N_15612,N_15560);
xor U15718 (N_15718,N_15221,N_15519);
xnor U15719 (N_15719,N_15431,N_15199);
xnor U15720 (N_15720,N_15240,N_15479);
or U15721 (N_15721,N_15502,N_15227);
and U15722 (N_15722,N_15491,N_15169);
and U15723 (N_15723,N_15362,N_15605);
xor U15724 (N_15724,N_15019,N_15482);
nand U15725 (N_15725,N_15542,N_15041);
or U15726 (N_15726,N_15470,N_15160);
xor U15727 (N_15727,N_15496,N_15030);
or U15728 (N_15728,N_15422,N_15003);
xnor U15729 (N_15729,N_15143,N_15029);
nand U15730 (N_15730,N_15345,N_15423);
xnor U15731 (N_15731,N_15205,N_15134);
xor U15732 (N_15732,N_15406,N_15301);
nand U15733 (N_15733,N_15507,N_15331);
xor U15734 (N_15734,N_15149,N_15173);
or U15735 (N_15735,N_15623,N_15357);
nand U15736 (N_15736,N_15392,N_15082);
nand U15737 (N_15737,N_15330,N_15505);
nor U15738 (N_15738,N_15559,N_15556);
and U15739 (N_15739,N_15308,N_15585);
or U15740 (N_15740,N_15124,N_15462);
nand U15741 (N_15741,N_15316,N_15579);
nand U15742 (N_15742,N_15622,N_15070);
and U15743 (N_15743,N_15052,N_15601);
xor U15744 (N_15744,N_15158,N_15208);
or U15745 (N_15745,N_15059,N_15352);
nor U15746 (N_15746,N_15191,N_15150);
nor U15747 (N_15747,N_15068,N_15016);
or U15748 (N_15748,N_15126,N_15515);
and U15749 (N_15749,N_15524,N_15472);
or U15750 (N_15750,N_15119,N_15044);
nand U15751 (N_15751,N_15440,N_15481);
and U15752 (N_15752,N_15254,N_15116);
and U15753 (N_15753,N_15021,N_15596);
nand U15754 (N_15754,N_15418,N_15365);
nor U15755 (N_15755,N_15424,N_15450);
nor U15756 (N_15756,N_15174,N_15436);
or U15757 (N_15757,N_15527,N_15427);
nor U15758 (N_15758,N_15334,N_15192);
or U15759 (N_15759,N_15008,N_15546);
xor U15760 (N_15760,N_15583,N_15223);
or U15761 (N_15761,N_15255,N_15394);
nand U15762 (N_15762,N_15176,N_15159);
or U15763 (N_15763,N_15387,N_15541);
or U15764 (N_15764,N_15053,N_15615);
and U15765 (N_15765,N_15484,N_15244);
nor U15766 (N_15766,N_15588,N_15101);
and U15767 (N_15767,N_15333,N_15064);
and U15768 (N_15768,N_15218,N_15298);
and U15769 (N_15769,N_15257,N_15004);
and U15770 (N_15770,N_15621,N_15483);
xnor U15771 (N_15771,N_15210,N_15396);
or U15772 (N_15772,N_15411,N_15497);
and U15773 (N_15773,N_15587,N_15315);
and U15774 (N_15774,N_15214,N_15239);
nand U15775 (N_15775,N_15097,N_15374);
and U15776 (N_15776,N_15104,N_15598);
or U15777 (N_15777,N_15380,N_15121);
nor U15778 (N_15778,N_15342,N_15012);
xor U15779 (N_15779,N_15400,N_15237);
and U15780 (N_15780,N_15285,N_15504);
nand U15781 (N_15781,N_15448,N_15500);
nand U15782 (N_15782,N_15350,N_15164);
nor U15783 (N_15783,N_15571,N_15370);
and U15784 (N_15784,N_15487,N_15194);
nand U15785 (N_15785,N_15545,N_15610);
nor U15786 (N_15786,N_15368,N_15375);
nor U15787 (N_15787,N_15426,N_15554);
and U15788 (N_15788,N_15619,N_15032);
nand U15789 (N_15789,N_15187,N_15328);
or U15790 (N_15790,N_15383,N_15531);
and U15791 (N_15791,N_15474,N_15268);
or U15792 (N_15792,N_15314,N_15521);
and U15793 (N_15793,N_15271,N_15573);
nor U15794 (N_15794,N_15272,N_15576);
xnor U15795 (N_15795,N_15312,N_15180);
and U15796 (N_15796,N_15179,N_15112);
xnor U15797 (N_15797,N_15252,N_15025);
or U15798 (N_15798,N_15338,N_15584);
nor U15799 (N_15799,N_15393,N_15512);
nand U15800 (N_15800,N_15061,N_15421);
or U15801 (N_15801,N_15109,N_15335);
nor U15802 (N_15802,N_15246,N_15224);
nand U15803 (N_15803,N_15274,N_15142);
xor U15804 (N_15804,N_15390,N_15074);
or U15805 (N_15805,N_15193,N_15537);
xnor U15806 (N_15806,N_15093,N_15578);
or U15807 (N_15807,N_15547,N_15324);
or U15808 (N_15808,N_15360,N_15203);
and U15809 (N_15809,N_15096,N_15113);
xor U15810 (N_15810,N_15318,N_15098);
nor U15811 (N_15811,N_15415,N_15561);
xnor U15812 (N_15812,N_15543,N_15388);
or U15813 (N_15813,N_15361,N_15307);
nand U15814 (N_15814,N_15073,N_15136);
and U15815 (N_15815,N_15550,N_15434);
nand U15816 (N_15816,N_15200,N_15493);
and U15817 (N_15817,N_15006,N_15075);
and U15818 (N_15818,N_15544,N_15154);
xnor U15819 (N_15819,N_15107,N_15100);
nand U15820 (N_15820,N_15057,N_15514);
xor U15821 (N_15821,N_15453,N_15296);
or U15822 (N_15822,N_15595,N_15501);
or U15823 (N_15823,N_15105,N_15233);
nor U15824 (N_15824,N_15117,N_15213);
nor U15825 (N_15825,N_15469,N_15503);
nor U15826 (N_15826,N_15092,N_15606);
nor U15827 (N_15827,N_15076,N_15534);
and U15828 (N_15828,N_15384,N_15419);
xor U15829 (N_15829,N_15609,N_15538);
nand U15830 (N_15830,N_15336,N_15405);
or U15831 (N_15831,N_15111,N_15477);
and U15832 (N_15832,N_15086,N_15532);
and U15833 (N_15833,N_15321,N_15091);
nor U15834 (N_15834,N_15048,N_15359);
nand U15835 (N_15835,N_15251,N_15242);
nor U15836 (N_15836,N_15138,N_15265);
or U15837 (N_15837,N_15413,N_15581);
nor U15838 (N_15838,N_15485,N_15395);
nor U15839 (N_15839,N_15367,N_15326);
and U15840 (N_15840,N_15184,N_15486);
nor U15841 (N_15841,N_15060,N_15231);
and U15842 (N_15842,N_15425,N_15467);
xnor U15843 (N_15843,N_15256,N_15219);
and U15844 (N_15844,N_15552,N_15077);
nand U15845 (N_15845,N_15035,N_15258);
nor U15846 (N_15846,N_15197,N_15302);
nand U15847 (N_15847,N_15449,N_15510);
nor U15848 (N_15848,N_15209,N_15284);
nand U15849 (N_15849,N_15373,N_15611);
or U15850 (N_15850,N_15607,N_15190);
nor U15851 (N_15851,N_15291,N_15339);
nor U15852 (N_15852,N_15325,N_15329);
or U15853 (N_15853,N_15132,N_15414);
nand U15854 (N_15854,N_15305,N_15178);
nor U15855 (N_15855,N_15529,N_15250);
nand U15856 (N_15856,N_15292,N_15011);
and U15857 (N_15857,N_15054,N_15377);
xnor U15858 (N_15858,N_15114,N_15473);
nand U15859 (N_15859,N_15095,N_15071);
nor U15860 (N_15860,N_15344,N_15351);
or U15861 (N_15861,N_15616,N_15153);
nor U15862 (N_15862,N_15518,N_15106);
and U15863 (N_15863,N_15580,N_15603);
nor U15864 (N_15864,N_15476,N_15404);
or U15865 (N_15865,N_15618,N_15279);
nor U15866 (N_15866,N_15617,N_15177);
xor U15867 (N_15867,N_15013,N_15201);
and U15868 (N_15868,N_15230,N_15382);
nor U15869 (N_15869,N_15020,N_15080);
nand U15870 (N_15870,N_15458,N_15015);
nor U15871 (N_15871,N_15412,N_15548);
and U15872 (N_15872,N_15402,N_15433);
and U15873 (N_15873,N_15135,N_15420);
nand U15874 (N_15874,N_15181,N_15028);
or U15875 (N_15875,N_15249,N_15065);
nand U15876 (N_15876,N_15567,N_15081);
nand U15877 (N_15877,N_15498,N_15062);
xnor U15878 (N_15878,N_15040,N_15027);
nand U15879 (N_15879,N_15533,N_15253);
or U15880 (N_15880,N_15225,N_15323);
nor U15881 (N_15881,N_15189,N_15385);
and U15882 (N_15882,N_15000,N_15072);
or U15883 (N_15883,N_15354,N_15452);
nor U15884 (N_15884,N_15327,N_15288);
nand U15885 (N_15885,N_15386,N_15088);
xor U15886 (N_15886,N_15120,N_15557);
xnor U15887 (N_15887,N_15454,N_15608);
nor U15888 (N_15888,N_15168,N_15297);
nand U15889 (N_15889,N_15528,N_15613);
or U15890 (N_15890,N_15478,N_15582);
or U15891 (N_15891,N_15067,N_15295);
nor U15892 (N_15892,N_15228,N_15460);
xnor U15893 (N_15893,N_15017,N_15151);
or U15894 (N_15894,N_15034,N_15002);
and U15895 (N_15895,N_15341,N_15001);
nand U15896 (N_15896,N_15309,N_15461);
xor U15897 (N_15897,N_15195,N_15122);
nor U15898 (N_15898,N_15604,N_15401);
and U15899 (N_15899,N_15293,N_15569);
or U15900 (N_15900,N_15348,N_15523);
and U15901 (N_15901,N_15043,N_15198);
nand U15902 (N_15902,N_15574,N_15236);
nand U15903 (N_15903,N_15456,N_15024);
and U15904 (N_15904,N_15172,N_15443);
or U15905 (N_15905,N_15551,N_15432);
or U15906 (N_15906,N_15356,N_15229);
and U15907 (N_15907,N_15115,N_15022);
xnor U15908 (N_15908,N_15269,N_15131);
and U15909 (N_15909,N_15129,N_15085);
and U15910 (N_15910,N_15042,N_15408);
xor U15911 (N_15911,N_15216,N_15600);
nand U15912 (N_15912,N_15304,N_15441);
nor U15913 (N_15913,N_15238,N_15437);
nor U15914 (N_15914,N_15069,N_15152);
xor U15915 (N_15915,N_15430,N_15036);
or U15916 (N_15916,N_15513,N_15389);
and U15917 (N_15917,N_15063,N_15589);
nor U15918 (N_15918,N_15278,N_15506);
xor U15919 (N_15919,N_15157,N_15572);
or U15920 (N_15920,N_15366,N_15083);
xor U15921 (N_15921,N_15141,N_15163);
or U15922 (N_15922,N_15289,N_15320);
nor U15923 (N_15923,N_15376,N_15099);
xor U15924 (N_15924,N_15090,N_15162);
nor U15925 (N_15925,N_15332,N_15492);
or U15926 (N_15926,N_15039,N_15494);
and U15927 (N_15927,N_15347,N_15267);
and U15928 (N_15928,N_15018,N_15196);
nor U15929 (N_15929,N_15294,N_15089);
or U15930 (N_15930,N_15488,N_15045);
xnor U15931 (N_15931,N_15516,N_15337);
and U15932 (N_15932,N_15211,N_15624);
xor U15933 (N_15933,N_15340,N_15222);
nor U15934 (N_15934,N_15517,N_15038);
nand U15935 (N_15935,N_15364,N_15259);
xnor U15936 (N_15936,N_15536,N_15575);
nor U15937 (N_15937,N_15530,N_15021);
xnor U15938 (N_15938,N_15170,N_15319);
or U15939 (N_15939,N_15579,N_15352);
or U15940 (N_15940,N_15545,N_15366);
nand U15941 (N_15941,N_15563,N_15175);
nand U15942 (N_15942,N_15219,N_15542);
and U15943 (N_15943,N_15316,N_15587);
or U15944 (N_15944,N_15553,N_15251);
xor U15945 (N_15945,N_15613,N_15275);
xnor U15946 (N_15946,N_15291,N_15201);
or U15947 (N_15947,N_15003,N_15209);
and U15948 (N_15948,N_15623,N_15511);
nor U15949 (N_15949,N_15443,N_15187);
nand U15950 (N_15950,N_15417,N_15256);
nor U15951 (N_15951,N_15178,N_15454);
or U15952 (N_15952,N_15375,N_15149);
xnor U15953 (N_15953,N_15246,N_15534);
xor U15954 (N_15954,N_15408,N_15445);
and U15955 (N_15955,N_15205,N_15186);
xnor U15956 (N_15956,N_15167,N_15135);
xnor U15957 (N_15957,N_15551,N_15030);
xor U15958 (N_15958,N_15028,N_15532);
or U15959 (N_15959,N_15446,N_15255);
or U15960 (N_15960,N_15399,N_15526);
nor U15961 (N_15961,N_15325,N_15509);
nand U15962 (N_15962,N_15459,N_15464);
nand U15963 (N_15963,N_15322,N_15583);
nor U15964 (N_15964,N_15059,N_15427);
nor U15965 (N_15965,N_15354,N_15581);
xor U15966 (N_15966,N_15602,N_15561);
and U15967 (N_15967,N_15062,N_15107);
or U15968 (N_15968,N_15167,N_15372);
xor U15969 (N_15969,N_15609,N_15314);
xor U15970 (N_15970,N_15187,N_15058);
nor U15971 (N_15971,N_15393,N_15421);
xnor U15972 (N_15972,N_15291,N_15482);
xor U15973 (N_15973,N_15004,N_15593);
nor U15974 (N_15974,N_15319,N_15435);
xnor U15975 (N_15975,N_15136,N_15306);
xnor U15976 (N_15976,N_15196,N_15457);
and U15977 (N_15977,N_15535,N_15181);
nor U15978 (N_15978,N_15325,N_15566);
nand U15979 (N_15979,N_15529,N_15348);
xnor U15980 (N_15980,N_15095,N_15218);
and U15981 (N_15981,N_15521,N_15397);
xnor U15982 (N_15982,N_15581,N_15082);
nand U15983 (N_15983,N_15031,N_15184);
or U15984 (N_15984,N_15484,N_15495);
nand U15985 (N_15985,N_15061,N_15588);
xnor U15986 (N_15986,N_15573,N_15103);
nor U15987 (N_15987,N_15573,N_15447);
xnor U15988 (N_15988,N_15540,N_15513);
or U15989 (N_15989,N_15009,N_15071);
xor U15990 (N_15990,N_15358,N_15445);
nor U15991 (N_15991,N_15286,N_15150);
nand U15992 (N_15992,N_15615,N_15521);
or U15993 (N_15993,N_15600,N_15072);
or U15994 (N_15994,N_15263,N_15219);
nand U15995 (N_15995,N_15596,N_15559);
nor U15996 (N_15996,N_15090,N_15454);
nand U15997 (N_15997,N_15516,N_15271);
and U15998 (N_15998,N_15622,N_15150);
xor U15999 (N_15999,N_15434,N_15285);
xor U16000 (N_16000,N_15502,N_15600);
nor U16001 (N_16001,N_15080,N_15452);
and U16002 (N_16002,N_15624,N_15081);
nor U16003 (N_16003,N_15190,N_15179);
or U16004 (N_16004,N_15087,N_15263);
xor U16005 (N_16005,N_15464,N_15126);
xnor U16006 (N_16006,N_15326,N_15002);
or U16007 (N_16007,N_15143,N_15192);
and U16008 (N_16008,N_15596,N_15454);
and U16009 (N_16009,N_15258,N_15254);
nor U16010 (N_16010,N_15272,N_15446);
nor U16011 (N_16011,N_15480,N_15011);
nand U16012 (N_16012,N_15192,N_15076);
nor U16013 (N_16013,N_15073,N_15030);
and U16014 (N_16014,N_15388,N_15173);
and U16015 (N_16015,N_15619,N_15042);
and U16016 (N_16016,N_15496,N_15377);
nand U16017 (N_16017,N_15586,N_15481);
nand U16018 (N_16018,N_15166,N_15376);
and U16019 (N_16019,N_15560,N_15486);
and U16020 (N_16020,N_15015,N_15319);
or U16021 (N_16021,N_15155,N_15003);
and U16022 (N_16022,N_15225,N_15266);
xor U16023 (N_16023,N_15237,N_15456);
and U16024 (N_16024,N_15485,N_15198);
nand U16025 (N_16025,N_15025,N_15607);
xor U16026 (N_16026,N_15068,N_15004);
xnor U16027 (N_16027,N_15359,N_15112);
nand U16028 (N_16028,N_15095,N_15363);
and U16029 (N_16029,N_15007,N_15380);
and U16030 (N_16030,N_15571,N_15599);
nor U16031 (N_16031,N_15590,N_15005);
and U16032 (N_16032,N_15416,N_15231);
or U16033 (N_16033,N_15326,N_15398);
and U16034 (N_16034,N_15151,N_15229);
or U16035 (N_16035,N_15505,N_15234);
nor U16036 (N_16036,N_15435,N_15004);
and U16037 (N_16037,N_15175,N_15125);
nor U16038 (N_16038,N_15032,N_15077);
or U16039 (N_16039,N_15191,N_15472);
xor U16040 (N_16040,N_15171,N_15106);
and U16041 (N_16041,N_15217,N_15430);
or U16042 (N_16042,N_15134,N_15543);
or U16043 (N_16043,N_15098,N_15471);
nor U16044 (N_16044,N_15376,N_15537);
xnor U16045 (N_16045,N_15137,N_15035);
and U16046 (N_16046,N_15517,N_15577);
or U16047 (N_16047,N_15104,N_15142);
nand U16048 (N_16048,N_15613,N_15470);
or U16049 (N_16049,N_15522,N_15311);
nand U16050 (N_16050,N_15281,N_15078);
xnor U16051 (N_16051,N_15065,N_15503);
and U16052 (N_16052,N_15619,N_15476);
nand U16053 (N_16053,N_15027,N_15524);
nand U16054 (N_16054,N_15118,N_15114);
nand U16055 (N_16055,N_15426,N_15425);
and U16056 (N_16056,N_15054,N_15180);
and U16057 (N_16057,N_15050,N_15608);
or U16058 (N_16058,N_15194,N_15209);
or U16059 (N_16059,N_15122,N_15359);
and U16060 (N_16060,N_15544,N_15433);
and U16061 (N_16061,N_15551,N_15244);
or U16062 (N_16062,N_15389,N_15037);
nor U16063 (N_16063,N_15056,N_15256);
nand U16064 (N_16064,N_15336,N_15611);
nor U16065 (N_16065,N_15176,N_15624);
nand U16066 (N_16066,N_15110,N_15403);
xnor U16067 (N_16067,N_15064,N_15253);
or U16068 (N_16068,N_15560,N_15515);
xnor U16069 (N_16069,N_15094,N_15262);
nor U16070 (N_16070,N_15168,N_15086);
or U16071 (N_16071,N_15352,N_15208);
and U16072 (N_16072,N_15254,N_15107);
nand U16073 (N_16073,N_15293,N_15487);
xnor U16074 (N_16074,N_15595,N_15327);
and U16075 (N_16075,N_15236,N_15026);
or U16076 (N_16076,N_15410,N_15578);
or U16077 (N_16077,N_15569,N_15287);
nand U16078 (N_16078,N_15531,N_15427);
or U16079 (N_16079,N_15158,N_15397);
xor U16080 (N_16080,N_15131,N_15537);
nor U16081 (N_16081,N_15176,N_15286);
nor U16082 (N_16082,N_15350,N_15407);
nor U16083 (N_16083,N_15513,N_15281);
nand U16084 (N_16084,N_15599,N_15135);
and U16085 (N_16085,N_15284,N_15182);
nand U16086 (N_16086,N_15099,N_15591);
nand U16087 (N_16087,N_15344,N_15273);
nor U16088 (N_16088,N_15289,N_15315);
nand U16089 (N_16089,N_15198,N_15182);
nor U16090 (N_16090,N_15570,N_15586);
and U16091 (N_16091,N_15208,N_15395);
nor U16092 (N_16092,N_15037,N_15345);
nor U16093 (N_16093,N_15095,N_15467);
nor U16094 (N_16094,N_15158,N_15069);
nand U16095 (N_16095,N_15612,N_15076);
xor U16096 (N_16096,N_15168,N_15089);
nor U16097 (N_16097,N_15257,N_15041);
nand U16098 (N_16098,N_15101,N_15152);
xnor U16099 (N_16099,N_15473,N_15562);
and U16100 (N_16100,N_15110,N_15385);
and U16101 (N_16101,N_15481,N_15433);
or U16102 (N_16102,N_15322,N_15573);
or U16103 (N_16103,N_15361,N_15013);
or U16104 (N_16104,N_15097,N_15235);
and U16105 (N_16105,N_15379,N_15451);
xor U16106 (N_16106,N_15219,N_15436);
or U16107 (N_16107,N_15131,N_15505);
nand U16108 (N_16108,N_15045,N_15432);
nand U16109 (N_16109,N_15164,N_15348);
and U16110 (N_16110,N_15222,N_15180);
or U16111 (N_16111,N_15471,N_15131);
xnor U16112 (N_16112,N_15602,N_15425);
xor U16113 (N_16113,N_15337,N_15198);
nor U16114 (N_16114,N_15252,N_15247);
nor U16115 (N_16115,N_15361,N_15049);
nand U16116 (N_16116,N_15187,N_15371);
and U16117 (N_16117,N_15227,N_15555);
xnor U16118 (N_16118,N_15029,N_15582);
xnor U16119 (N_16119,N_15482,N_15602);
xor U16120 (N_16120,N_15244,N_15436);
nor U16121 (N_16121,N_15112,N_15345);
nand U16122 (N_16122,N_15385,N_15037);
nand U16123 (N_16123,N_15226,N_15481);
or U16124 (N_16124,N_15087,N_15109);
nor U16125 (N_16125,N_15585,N_15217);
or U16126 (N_16126,N_15618,N_15156);
and U16127 (N_16127,N_15409,N_15169);
nand U16128 (N_16128,N_15052,N_15410);
nand U16129 (N_16129,N_15296,N_15369);
xor U16130 (N_16130,N_15093,N_15127);
xnor U16131 (N_16131,N_15581,N_15461);
nand U16132 (N_16132,N_15550,N_15321);
nand U16133 (N_16133,N_15069,N_15511);
or U16134 (N_16134,N_15015,N_15368);
nand U16135 (N_16135,N_15019,N_15146);
nor U16136 (N_16136,N_15129,N_15446);
xor U16137 (N_16137,N_15211,N_15114);
xnor U16138 (N_16138,N_15375,N_15492);
nor U16139 (N_16139,N_15121,N_15234);
nor U16140 (N_16140,N_15166,N_15200);
nor U16141 (N_16141,N_15151,N_15242);
and U16142 (N_16142,N_15604,N_15167);
xnor U16143 (N_16143,N_15272,N_15024);
and U16144 (N_16144,N_15556,N_15124);
nor U16145 (N_16145,N_15531,N_15601);
xnor U16146 (N_16146,N_15133,N_15423);
nor U16147 (N_16147,N_15020,N_15207);
xor U16148 (N_16148,N_15384,N_15084);
nand U16149 (N_16149,N_15479,N_15200);
or U16150 (N_16150,N_15385,N_15244);
nor U16151 (N_16151,N_15479,N_15502);
nor U16152 (N_16152,N_15572,N_15520);
nand U16153 (N_16153,N_15132,N_15182);
nand U16154 (N_16154,N_15208,N_15020);
nor U16155 (N_16155,N_15582,N_15090);
nor U16156 (N_16156,N_15587,N_15021);
nor U16157 (N_16157,N_15548,N_15583);
and U16158 (N_16158,N_15511,N_15331);
nand U16159 (N_16159,N_15385,N_15446);
or U16160 (N_16160,N_15579,N_15207);
nand U16161 (N_16161,N_15597,N_15383);
or U16162 (N_16162,N_15401,N_15018);
nor U16163 (N_16163,N_15001,N_15461);
nor U16164 (N_16164,N_15218,N_15118);
or U16165 (N_16165,N_15127,N_15593);
xnor U16166 (N_16166,N_15198,N_15086);
nor U16167 (N_16167,N_15555,N_15359);
and U16168 (N_16168,N_15364,N_15564);
nand U16169 (N_16169,N_15250,N_15469);
and U16170 (N_16170,N_15067,N_15031);
and U16171 (N_16171,N_15217,N_15138);
and U16172 (N_16172,N_15475,N_15225);
or U16173 (N_16173,N_15576,N_15144);
nand U16174 (N_16174,N_15157,N_15352);
xnor U16175 (N_16175,N_15596,N_15452);
nor U16176 (N_16176,N_15101,N_15606);
nor U16177 (N_16177,N_15200,N_15548);
or U16178 (N_16178,N_15254,N_15597);
xor U16179 (N_16179,N_15449,N_15468);
nor U16180 (N_16180,N_15160,N_15468);
xor U16181 (N_16181,N_15461,N_15443);
nor U16182 (N_16182,N_15025,N_15085);
nor U16183 (N_16183,N_15377,N_15094);
nand U16184 (N_16184,N_15417,N_15389);
nand U16185 (N_16185,N_15335,N_15540);
nor U16186 (N_16186,N_15232,N_15574);
xnor U16187 (N_16187,N_15318,N_15545);
nand U16188 (N_16188,N_15038,N_15356);
and U16189 (N_16189,N_15096,N_15585);
nor U16190 (N_16190,N_15603,N_15177);
xnor U16191 (N_16191,N_15202,N_15262);
xnor U16192 (N_16192,N_15343,N_15230);
or U16193 (N_16193,N_15406,N_15038);
nor U16194 (N_16194,N_15289,N_15514);
nand U16195 (N_16195,N_15293,N_15426);
nor U16196 (N_16196,N_15483,N_15076);
or U16197 (N_16197,N_15182,N_15445);
or U16198 (N_16198,N_15078,N_15063);
nand U16199 (N_16199,N_15188,N_15542);
and U16200 (N_16200,N_15473,N_15614);
nand U16201 (N_16201,N_15272,N_15497);
nand U16202 (N_16202,N_15176,N_15462);
nand U16203 (N_16203,N_15527,N_15036);
xnor U16204 (N_16204,N_15406,N_15581);
and U16205 (N_16205,N_15149,N_15452);
and U16206 (N_16206,N_15522,N_15258);
xnor U16207 (N_16207,N_15040,N_15268);
or U16208 (N_16208,N_15543,N_15171);
or U16209 (N_16209,N_15559,N_15140);
or U16210 (N_16210,N_15479,N_15375);
xnor U16211 (N_16211,N_15283,N_15613);
and U16212 (N_16212,N_15264,N_15330);
nor U16213 (N_16213,N_15114,N_15090);
and U16214 (N_16214,N_15347,N_15106);
nor U16215 (N_16215,N_15602,N_15284);
xnor U16216 (N_16216,N_15459,N_15204);
nand U16217 (N_16217,N_15501,N_15398);
nand U16218 (N_16218,N_15423,N_15212);
and U16219 (N_16219,N_15312,N_15186);
or U16220 (N_16220,N_15109,N_15003);
xnor U16221 (N_16221,N_15180,N_15457);
and U16222 (N_16222,N_15204,N_15084);
nor U16223 (N_16223,N_15605,N_15622);
and U16224 (N_16224,N_15434,N_15344);
nor U16225 (N_16225,N_15534,N_15416);
nor U16226 (N_16226,N_15297,N_15624);
or U16227 (N_16227,N_15461,N_15624);
nor U16228 (N_16228,N_15167,N_15286);
and U16229 (N_16229,N_15352,N_15167);
xor U16230 (N_16230,N_15043,N_15051);
and U16231 (N_16231,N_15181,N_15269);
nor U16232 (N_16232,N_15336,N_15122);
or U16233 (N_16233,N_15328,N_15524);
nor U16234 (N_16234,N_15526,N_15133);
or U16235 (N_16235,N_15465,N_15348);
or U16236 (N_16236,N_15072,N_15430);
or U16237 (N_16237,N_15429,N_15285);
nand U16238 (N_16238,N_15376,N_15130);
or U16239 (N_16239,N_15357,N_15294);
or U16240 (N_16240,N_15357,N_15168);
nand U16241 (N_16241,N_15229,N_15075);
and U16242 (N_16242,N_15199,N_15460);
xor U16243 (N_16243,N_15529,N_15180);
and U16244 (N_16244,N_15228,N_15069);
xnor U16245 (N_16245,N_15165,N_15566);
xor U16246 (N_16246,N_15471,N_15509);
nor U16247 (N_16247,N_15469,N_15520);
xor U16248 (N_16248,N_15089,N_15108);
and U16249 (N_16249,N_15067,N_15137);
and U16250 (N_16250,N_16136,N_15713);
and U16251 (N_16251,N_15655,N_15892);
and U16252 (N_16252,N_15946,N_16092);
xor U16253 (N_16253,N_16204,N_15684);
and U16254 (N_16254,N_15945,N_15634);
or U16255 (N_16255,N_15727,N_15660);
nand U16256 (N_16256,N_16030,N_15954);
or U16257 (N_16257,N_15978,N_16071);
or U16258 (N_16258,N_15707,N_16165);
and U16259 (N_16259,N_16208,N_16052);
nand U16260 (N_16260,N_15724,N_15725);
nor U16261 (N_16261,N_15692,N_16176);
nand U16262 (N_16262,N_16227,N_15959);
or U16263 (N_16263,N_15890,N_15891);
or U16264 (N_16264,N_15794,N_16199);
nand U16265 (N_16265,N_15714,N_16170);
nor U16266 (N_16266,N_15759,N_16110);
nor U16267 (N_16267,N_16184,N_15732);
nor U16268 (N_16268,N_16181,N_15632);
nor U16269 (N_16269,N_15793,N_16230);
or U16270 (N_16270,N_15960,N_15918);
nand U16271 (N_16271,N_15821,N_15803);
nor U16272 (N_16272,N_15653,N_15943);
and U16273 (N_16273,N_16241,N_16049);
nor U16274 (N_16274,N_15916,N_16141);
and U16275 (N_16275,N_16025,N_15845);
or U16276 (N_16276,N_15770,N_16143);
or U16277 (N_16277,N_16095,N_15736);
xnor U16278 (N_16278,N_15630,N_15764);
nand U16279 (N_16279,N_16187,N_15828);
nor U16280 (N_16280,N_15756,N_15863);
or U16281 (N_16281,N_15932,N_15939);
nand U16282 (N_16282,N_16157,N_15651);
and U16283 (N_16283,N_16166,N_15846);
and U16284 (N_16284,N_16015,N_16216);
nor U16285 (N_16285,N_15919,N_16192);
nand U16286 (N_16286,N_15799,N_16103);
nor U16287 (N_16287,N_15710,N_16243);
nor U16288 (N_16288,N_15666,N_16068);
and U16289 (N_16289,N_15875,N_15685);
nand U16290 (N_16290,N_16084,N_16182);
and U16291 (N_16291,N_15762,N_15995);
nor U16292 (N_16292,N_15831,N_15937);
nor U16293 (N_16293,N_16116,N_16244);
nand U16294 (N_16294,N_15789,N_16145);
xor U16295 (N_16295,N_16212,N_15984);
nor U16296 (N_16296,N_15872,N_16233);
nand U16297 (N_16297,N_15838,N_16123);
and U16298 (N_16298,N_16220,N_15687);
xor U16299 (N_16299,N_15869,N_15849);
nand U16300 (N_16300,N_15865,N_15885);
xnor U16301 (N_16301,N_16022,N_15740);
nand U16302 (N_16302,N_15683,N_16113);
xnor U16303 (N_16303,N_16105,N_15656);
and U16304 (N_16304,N_15867,N_15766);
and U16305 (N_16305,N_15862,N_16101);
nor U16306 (N_16306,N_15800,N_15807);
nor U16307 (N_16307,N_15626,N_15640);
nor U16308 (N_16308,N_16053,N_16147);
and U16309 (N_16309,N_16032,N_16185);
nor U16310 (N_16310,N_15778,N_15851);
and U16311 (N_16311,N_15933,N_16169);
nor U16312 (N_16312,N_15850,N_15643);
nand U16313 (N_16313,N_15680,N_16222);
nand U16314 (N_16314,N_15681,N_16081);
and U16315 (N_16315,N_15952,N_16029);
xnor U16316 (N_16316,N_16074,N_15797);
and U16317 (N_16317,N_16193,N_16137);
nor U16318 (N_16318,N_15925,N_15990);
nor U16319 (N_16319,N_15819,N_16229);
or U16320 (N_16320,N_15716,N_16205);
and U16321 (N_16321,N_16154,N_16044);
and U16322 (N_16322,N_16142,N_15809);
xor U16323 (N_16323,N_15813,N_15888);
nand U16324 (N_16324,N_15922,N_15751);
and U16325 (N_16325,N_15864,N_16162);
and U16326 (N_16326,N_15992,N_16221);
or U16327 (N_16327,N_15674,N_15745);
or U16328 (N_16328,N_15972,N_16000);
nor U16329 (N_16329,N_16218,N_15915);
nor U16330 (N_16330,N_15773,N_16094);
nand U16331 (N_16331,N_16002,N_16115);
xnor U16332 (N_16332,N_15742,N_15836);
and U16333 (N_16333,N_16106,N_16102);
nand U16334 (N_16334,N_16083,N_16189);
nand U16335 (N_16335,N_16001,N_16100);
and U16336 (N_16336,N_15844,N_15926);
xnor U16337 (N_16337,N_16086,N_16056);
nor U16338 (N_16338,N_15859,N_15798);
xor U16339 (N_16339,N_15883,N_15991);
and U16340 (N_16340,N_15782,N_16163);
or U16341 (N_16341,N_15839,N_16202);
or U16342 (N_16342,N_15750,N_15901);
and U16343 (N_16343,N_16159,N_15711);
or U16344 (N_16344,N_15763,N_15715);
xor U16345 (N_16345,N_15868,N_15955);
xor U16346 (N_16346,N_15893,N_15953);
nor U16347 (N_16347,N_16121,N_15729);
xor U16348 (N_16348,N_15835,N_15889);
nand U16349 (N_16349,N_15748,N_15934);
or U16350 (N_16350,N_15689,N_15823);
or U16351 (N_16351,N_16213,N_16235);
nand U16352 (N_16352,N_15817,N_15822);
nand U16353 (N_16353,N_15784,N_15895);
and U16354 (N_16354,N_15769,N_16160);
nor U16355 (N_16355,N_16042,N_15629);
nor U16356 (N_16356,N_15744,N_15765);
or U16357 (N_16357,N_16158,N_15987);
or U16358 (N_16358,N_15921,N_16190);
nor U16359 (N_16359,N_15733,N_15814);
nand U16360 (N_16360,N_16201,N_15967);
nor U16361 (N_16361,N_15975,N_15854);
and U16362 (N_16362,N_15699,N_16139);
nand U16363 (N_16363,N_16073,N_15738);
or U16364 (N_16364,N_15627,N_15876);
nor U16365 (N_16365,N_15974,N_15658);
or U16366 (N_16366,N_15812,N_15887);
nand U16367 (N_16367,N_16246,N_15996);
nand U16368 (N_16368,N_16174,N_15776);
nor U16369 (N_16369,N_15625,N_15777);
xnor U16370 (N_16370,N_15741,N_16003);
xor U16371 (N_16371,N_16228,N_15718);
and U16372 (N_16372,N_16172,N_16043);
and U16373 (N_16373,N_15944,N_16041);
nor U16374 (N_16374,N_16067,N_15752);
nand U16375 (N_16375,N_15785,N_15826);
nor U16376 (N_16376,N_15648,N_16045);
nand U16377 (N_16377,N_16186,N_16148);
and U16378 (N_16378,N_15962,N_16156);
nand U16379 (N_16379,N_15663,N_16206);
and U16380 (N_16380,N_16080,N_15772);
xnor U16381 (N_16381,N_15871,N_15897);
or U16382 (N_16382,N_16130,N_15841);
xnor U16383 (N_16383,N_16183,N_15870);
nand U16384 (N_16384,N_15982,N_16017);
xnor U16385 (N_16385,N_15726,N_16033);
xor U16386 (N_16386,N_16180,N_16076);
or U16387 (N_16387,N_15679,N_15788);
nand U16388 (N_16388,N_15855,N_15896);
nand U16389 (N_16389,N_15950,N_15914);
xor U16390 (N_16390,N_15673,N_15903);
nor U16391 (N_16391,N_16104,N_16098);
or U16392 (N_16392,N_15644,N_15938);
nor U16393 (N_16393,N_16027,N_15816);
nand U16394 (N_16394,N_15697,N_15979);
xor U16395 (N_16395,N_16038,N_16082);
xor U16396 (N_16396,N_16050,N_15804);
nand U16397 (N_16397,N_15912,N_16062);
and U16398 (N_16398,N_16236,N_15830);
nand U16399 (N_16399,N_15675,N_15677);
xor U16400 (N_16400,N_16088,N_15704);
or U16401 (N_16401,N_15913,N_16069);
xor U16402 (N_16402,N_15881,N_15811);
or U16403 (N_16403,N_15693,N_15678);
nor U16404 (N_16404,N_15635,N_16061);
xor U16405 (N_16405,N_15909,N_16217);
or U16406 (N_16406,N_16198,N_16087);
nand U16407 (N_16407,N_15976,N_15873);
or U16408 (N_16408,N_15723,N_15927);
xnor U16409 (N_16409,N_16168,N_15721);
or U16410 (N_16410,N_16125,N_15637);
and U16411 (N_16411,N_15880,N_16231);
nand U16412 (N_16412,N_15942,N_16135);
nand U16413 (N_16413,N_15998,N_15902);
or U16414 (N_16414,N_16091,N_15791);
and U16415 (N_16415,N_16239,N_15825);
and U16416 (N_16416,N_15661,N_15815);
or U16417 (N_16417,N_15667,N_16023);
and U16418 (N_16418,N_16026,N_16014);
nand U16419 (N_16419,N_15801,N_15917);
nand U16420 (N_16420,N_16112,N_15747);
or U16421 (N_16421,N_15795,N_15786);
or U16422 (N_16422,N_16240,N_15861);
nor U16423 (N_16423,N_15818,N_16215);
or U16424 (N_16424,N_16118,N_16065);
nand U16425 (N_16425,N_16099,N_15884);
nand U16426 (N_16426,N_15698,N_15796);
or U16427 (N_16427,N_16191,N_15717);
xor U16428 (N_16428,N_15860,N_15771);
or U16429 (N_16429,N_16072,N_15672);
and U16430 (N_16430,N_16119,N_15628);
or U16431 (N_16431,N_16128,N_16093);
or U16432 (N_16432,N_15709,N_16150);
nand U16433 (N_16433,N_16097,N_15970);
xnor U16434 (N_16434,N_15965,N_15702);
and U16435 (N_16435,N_16047,N_15877);
nand U16436 (N_16436,N_15806,N_16005);
xor U16437 (N_16437,N_16211,N_16196);
nand U16438 (N_16438,N_15905,N_15706);
and U16439 (N_16439,N_15690,N_15827);
or U16440 (N_16440,N_16109,N_16161);
or U16441 (N_16441,N_15935,N_15688);
and U16442 (N_16442,N_15805,N_15908);
xor U16443 (N_16443,N_15966,N_15758);
nand U16444 (N_16444,N_15951,N_15856);
xnor U16445 (N_16445,N_16124,N_16127);
nor U16446 (N_16446,N_15981,N_15654);
and U16447 (N_16447,N_15924,N_15829);
nor U16448 (N_16448,N_15923,N_15842);
nand U16449 (N_16449,N_15963,N_16085);
nand U16450 (N_16450,N_16167,N_16096);
or U16451 (N_16451,N_16070,N_16077);
nand U16452 (N_16452,N_15936,N_16010);
nor U16453 (N_16453,N_15997,N_15941);
and U16454 (N_16454,N_15650,N_16089);
or U16455 (N_16455,N_15852,N_15719);
or U16456 (N_16456,N_16090,N_15768);
and U16457 (N_16457,N_15969,N_16059);
or U16458 (N_16458,N_15695,N_15682);
or U16459 (N_16459,N_15755,N_16200);
nor U16460 (N_16460,N_16203,N_16058);
nor U16461 (N_16461,N_15767,N_16179);
and U16462 (N_16462,N_15958,N_16232);
nand U16463 (N_16463,N_16131,N_15947);
nand U16464 (N_16464,N_15961,N_15708);
nand U16465 (N_16465,N_15730,N_15848);
xnor U16466 (N_16466,N_15670,N_16012);
xnor U16467 (N_16467,N_15761,N_15808);
nand U16468 (N_16468,N_16210,N_16018);
or U16469 (N_16469,N_15980,N_16078);
nor U16470 (N_16470,N_16075,N_16144);
and U16471 (N_16471,N_15712,N_15734);
nand U16472 (N_16472,N_16079,N_16060);
nand U16473 (N_16473,N_16152,N_15878);
nand U16474 (N_16474,N_15671,N_15832);
nor U16475 (N_16475,N_16138,N_15728);
or U16476 (N_16476,N_15900,N_15930);
and U16477 (N_16477,N_16237,N_15886);
nand U16478 (N_16478,N_16048,N_15874);
nand U16479 (N_16479,N_15866,N_16155);
and U16480 (N_16480,N_16146,N_15940);
nand U16481 (N_16481,N_16063,N_15701);
or U16482 (N_16482,N_15911,N_15781);
nor U16483 (N_16483,N_15657,N_15731);
nand U16484 (N_16484,N_15668,N_16016);
and U16485 (N_16485,N_16248,N_16126);
xnor U16486 (N_16486,N_16225,N_15647);
or U16487 (N_16487,N_15686,N_15920);
and U16488 (N_16488,N_16234,N_16140);
and U16489 (N_16489,N_15746,N_15760);
or U16490 (N_16490,N_15783,N_15971);
xor U16491 (N_16491,N_15847,N_16031);
nor U16492 (N_16492,N_16178,N_16209);
xnor U16493 (N_16493,N_16175,N_16207);
nand U16494 (N_16494,N_15691,N_16066);
nand U16495 (N_16495,N_15720,N_15705);
nor U16496 (N_16496,N_16013,N_15735);
xor U16497 (N_16497,N_16008,N_16224);
xor U16498 (N_16498,N_15993,N_16035);
or U16499 (N_16499,N_15994,N_15929);
or U16500 (N_16500,N_16219,N_15743);
xnor U16501 (N_16501,N_15931,N_15662);
nor U16502 (N_16502,N_15857,N_16108);
xor U16503 (N_16503,N_15739,N_15879);
or U16504 (N_16504,N_16021,N_16009);
or U16505 (N_16505,N_15638,N_15757);
or U16506 (N_16506,N_15986,N_15858);
and U16507 (N_16507,N_15833,N_16034);
nand U16508 (N_16508,N_16223,N_16197);
and U16509 (N_16509,N_16054,N_16214);
nand U16510 (N_16510,N_16046,N_16194);
nand U16511 (N_16511,N_15780,N_15753);
or U16512 (N_16512,N_15834,N_16249);
or U16513 (N_16513,N_16151,N_16164);
xnor U16514 (N_16514,N_15973,N_16134);
nand U16515 (N_16515,N_15641,N_16020);
nor U16516 (N_16516,N_15956,N_15636);
nand U16517 (N_16517,N_15703,N_15999);
or U16518 (N_16518,N_15906,N_15894);
and U16519 (N_16519,N_15988,N_15840);
and U16520 (N_16520,N_15843,N_16149);
and U16521 (N_16521,N_16004,N_16024);
nor U16522 (N_16522,N_15968,N_15722);
nor U16523 (N_16523,N_15949,N_15737);
nor U16524 (N_16524,N_15649,N_15899);
nand U16525 (N_16525,N_15790,N_15633);
nand U16526 (N_16526,N_15659,N_16133);
or U16527 (N_16527,N_16064,N_15957);
nor U16528 (N_16528,N_15837,N_16111);
or U16529 (N_16529,N_15792,N_16039);
nand U16530 (N_16530,N_15977,N_15669);
or U16531 (N_16531,N_15787,N_15882);
nor U16532 (N_16532,N_16117,N_15664);
or U16533 (N_16533,N_16037,N_15639);
or U16534 (N_16534,N_16120,N_15676);
and U16535 (N_16535,N_15824,N_16153);
and U16536 (N_16536,N_15802,N_16055);
nor U16537 (N_16537,N_16238,N_15779);
nor U16538 (N_16538,N_15853,N_15700);
or U16539 (N_16539,N_15646,N_16114);
or U16540 (N_16540,N_15820,N_16006);
nand U16541 (N_16541,N_15749,N_16132);
xnor U16542 (N_16542,N_16173,N_16129);
and U16543 (N_16543,N_16040,N_15910);
or U16544 (N_16544,N_15989,N_15948);
xnor U16545 (N_16545,N_15696,N_16188);
or U16546 (N_16546,N_15694,N_16036);
nand U16547 (N_16547,N_16011,N_15631);
nand U16548 (N_16548,N_15985,N_15642);
or U16549 (N_16549,N_15904,N_16007);
nor U16550 (N_16550,N_16028,N_15645);
and U16551 (N_16551,N_15754,N_16177);
or U16552 (N_16552,N_16242,N_15652);
or U16553 (N_16553,N_15665,N_16171);
and U16554 (N_16554,N_15775,N_16245);
nand U16555 (N_16555,N_16019,N_15907);
or U16556 (N_16556,N_16051,N_15983);
nor U16557 (N_16557,N_15810,N_16226);
nor U16558 (N_16558,N_15898,N_16107);
nor U16559 (N_16559,N_16247,N_16057);
nand U16560 (N_16560,N_16122,N_15928);
xor U16561 (N_16561,N_16195,N_15964);
nand U16562 (N_16562,N_15774,N_15631);
nand U16563 (N_16563,N_16058,N_16239);
nor U16564 (N_16564,N_16018,N_15699);
xnor U16565 (N_16565,N_15985,N_15807);
xor U16566 (N_16566,N_15672,N_15856);
nand U16567 (N_16567,N_15752,N_15952);
nor U16568 (N_16568,N_16120,N_15641);
nand U16569 (N_16569,N_15884,N_16012);
and U16570 (N_16570,N_15661,N_16118);
nor U16571 (N_16571,N_16125,N_15713);
or U16572 (N_16572,N_15937,N_15866);
or U16573 (N_16573,N_15787,N_16164);
xor U16574 (N_16574,N_15688,N_15806);
nor U16575 (N_16575,N_15849,N_16147);
nor U16576 (N_16576,N_15753,N_16184);
xnor U16577 (N_16577,N_15638,N_15654);
or U16578 (N_16578,N_16121,N_15989);
nor U16579 (N_16579,N_15702,N_15769);
or U16580 (N_16580,N_15714,N_15729);
and U16581 (N_16581,N_15636,N_15628);
or U16582 (N_16582,N_16200,N_15688);
and U16583 (N_16583,N_16055,N_15719);
and U16584 (N_16584,N_16082,N_15889);
nand U16585 (N_16585,N_16073,N_15666);
nor U16586 (N_16586,N_16090,N_16092);
or U16587 (N_16587,N_15845,N_15633);
nor U16588 (N_16588,N_16191,N_15940);
and U16589 (N_16589,N_16229,N_15677);
nor U16590 (N_16590,N_15758,N_16136);
or U16591 (N_16591,N_16022,N_15657);
nand U16592 (N_16592,N_15959,N_15832);
or U16593 (N_16593,N_15757,N_16101);
nand U16594 (N_16594,N_16036,N_15688);
nand U16595 (N_16595,N_16125,N_15631);
nand U16596 (N_16596,N_16247,N_15757);
nor U16597 (N_16597,N_15817,N_16047);
and U16598 (N_16598,N_16137,N_16148);
xnor U16599 (N_16599,N_16049,N_15637);
nor U16600 (N_16600,N_16202,N_15814);
and U16601 (N_16601,N_16245,N_15708);
nand U16602 (N_16602,N_15881,N_16208);
xnor U16603 (N_16603,N_16003,N_16073);
nor U16604 (N_16604,N_16128,N_16170);
nor U16605 (N_16605,N_16121,N_16012);
nand U16606 (N_16606,N_15662,N_16018);
xor U16607 (N_16607,N_15863,N_16137);
nand U16608 (N_16608,N_16112,N_15952);
nand U16609 (N_16609,N_15988,N_16044);
nand U16610 (N_16610,N_15998,N_15875);
nand U16611 (N_16611,N_16184,N_16049);
and U16612 (N_16612,N_15728,N_15925);
nor U16613 (N_16613,N_15950,N_15960);
xor U16614 (N_16614,N_16045,N_16171);
and U16615 (N_16615,N_16126,N_16034);
xnor U16616 (N_16616,N_15874,N_16061);
or U16617 (N_16617,N_16130,N_15827);
or U16618 (N_16618,N_15775,N_16033);
nand U16619 (N_16619,N_15634,N_15931);
and U16620 (N_16620,N_16198,N_15667);
nand U16621 (N_16621,N_15782,N_15874);
nand U16622 (N_16622,N_16052,N_15680);
xor U16623 (N_16623,N_16156,N_15687);
nand U16624 (N_16624,N_16085,N_15895);
xor U16625 (N_16625,N_15920,N_15774);
nor U16626 (N_16626,N_16006,N_15891);
nand U16627 (N_16627,N_15970,N_15813);
nand U16628 (N_16628,N_16124,N_16043);
and U16629 (N_16629,N_15962,N_15696);
xnor U16630 (N_16630,N_15745,N_15830);
nor U16631 (N_16631,N_15631,N_15825);
or U16632 (N_16632,N_16031,N_15661);
xnor U16633 (N_16633,N_15728,N_15779);
and U16634 (N_16634,N_16045,N_16158);
or U16635 (N_16635,N_16014,N_15710);
xnor U16636 (N_16636,N_15981,N_15694);
and U16637 (N_16637,N_16118,N_15742);
nand U16638 (N_16638,N_15801,N_16006);
nand U16639 (N_16639,N_15745,N_15638);
nand U16640 (N_16640,N_16150,N_15891);
and U16641 (N_16641,N_16064,N_15741);
nor U16642 (N_16642,N_15775,N_16005);
nand U16643 (N_16643,N_16035,N_16242);
xnor U16644 (N_16644,N_15706,N_15929);
xnor U16645 (N_16645,N_15628,N_16146);
or U16646 (N_16646,N_15791,N_15658);
xnor U16647 (N_16647,N_16194,N_15665);
xnor U16648 (N_16648,N_15791,N_15857);
nor U16649 (N_16649,N_16028,N_15708);
nand U16650 (N_16650,N_15689,N_15758);
and U16651 (N_16651,N_16151,N_16190);
xor U16652 (N_16652,N_16154,N_15716);
nand U16653 (N_16653,N_15957,N_16145);
nor U16654 (N_16654,N_16218,N_16031);
nand U16655 (N_16655,N_15737,N_15701);
nand U16656 (N_16656,N_15966,N_16220);
and U16657 (N_16657,N_16027,N_15797);
nand U16658 (N_16658,N_15965,N_15784);
nand U16659 (N_16659,N_16098,N_15636);
or U16660 (N_16660,N_16120,N_16234);
and U16661 (N_16661,N_15726,N_16193);
xor U16662 (N_16662,N_15800,N_15732);
nor U16663 (N_16663,N_15640,N_16010);
nor U16664 (N_16664,N_16231,N_15783);
nand U16665 (N_16665,N_16029,N_16077);
xnor U16666 (N_16666,N_15774,N_15883);
xor U16667 (N_16667,N_16059,N_15799);
or U16668 (N_16668,N_16032,N_15979);
nor U16669 (N_16669,N_16013,N_15922);
xor U16670 (N_16670,N_16157,N_16090);
nor U16671 (N_16671,N_16183,N_15683);
nand U16672 (N_16672,N_15787,N_16149);
nand U16673 (N_16673,N_16109,N_15645);
nand U16674 (N_16674,N_15625,N_15860);
nor U16675 (N_16675,N_15688,N_15864);
nand U16676 (N_16676,N_15766,N_16136);
nand U16677 (N_16677,N_16235,N_15787);
and U16678 (N_16678,N_15913,N_16225);
and U16679 (N_16679,N_15633,N_16235);
or U16680 (N_16680,N_15686,N_15974);
and U16681 (N_16681,N_15667,N_15951);
nor U16682 (N_16682,N_15736,N_15648);
or U16683 (N_16683,N_15793,N_16099);
xnor U16684 (N_16684,N_16227,N_15655);
and U16685 (N_16685,N_16147,N_15636);
xor U16686 (N_16686,N_15946,N_16203);
nand U16687 (N_16687,N_15792,N_15852);
and U16688 (N_16688,N_15822,N_15921);
nand U16689 (N_16689,N_15642,N_15737);
nand U16690 (N_16690,N_16088,N_15933);
and U16691 (N_16691,N_15783,N_15791);
xor U16692 (N_16692,N_15780,N_15895);
xnor U16693 (N_16693,N_15833,N_16001);
and U16694 (N_16694,N_15769,N_16071);
and U16695 (N_16695,N_16095,N_15822);
nor U16696 (N_16696,N_15993,N_15946);
and U16697 (N_16697,N_16224,N_15924);
or U16698 (N_16698,N_15798,N_15893);
or U16699 (N_16699,N_16152,N_16224);
nand U16700 (N_16700,N_16185,N_15970);
nand U16701 (N_16701,N_16142,N_16178);
and U16702 (N_16702,N_15923,N_16147);
or U16703 (N_16703,N_15813,N_15625);
nor U16704 (N_16704,N_15949,N_15638);
xor U16705 (N_16705,N_15712,N_16041);
nand U16706 (N_16706,N_15948,N_15954);
and U16707 (N_16707,N_15644,N_16218);
nand U16708 (N_16708,N_15796,N_15805);
nand U16709 (N_16709,N_15798,N_16035);
nand U16710 (N_16710,N_15842,N_16170);
xnor U16711 (N_16711,N_16121,N_15946);
xnor U16712 (N_16712,N_15692,N_15709);
or U16713 (N_16713,N_15652,N_15811);
xor U16714 (N_16714,N_16216,N_15731);
or U16715 (N_16715,N_15752,N_15973);
nand U16716 (N_16716,N_16188,N_15976);
xnor U16717 (N_16717,N_15895,N_16133);
nor U16718 (N_16718,N_16210,N_16026);
xor U16719 (N_16719,N_15676,N_15864);
nand U16720 (N_16720,N_15642,N_15848);
nand U16721 (N_16721,N_16222,N_15737);
nand U16722 (N_16722,N_15888,N_15630);
and U16723 (N_16723,N_15654,N_16083);
xnor U16724 (N_16724,N_16125,N_16054);
nor U16725 (N_16725,N_15918,N_15646);
nor U16726 (N_16726,N_15958,N_16130);
or U16727 (N_16727,N_15809,N_15906);
xnor U16728 (N_16728,N_15970,N_15748);
xor U16729 (N_16729,N_16131,N_15701);
or U16730 (N_16730,N_15626,N_16206);
or U16731 (N_16731,N_16009,N_16080);
nand U16732 (N_16732,N_16011,N_15679);
and U16733 (N_16733,N_16192,N_16141);
or U16734 (N_16734,N_16126,N_16199);
nand U16735 (N_16735,N_15808,N_15946);
nor U16736 (N_16736,N_16186,N_15726);
nand U16737 (N_16737,N_16150,N_15808);
xor U16738 (N_16738,N_16083,N_16105);
nor U16739 (N_16739,N_15866,N_15846);
nor U16740 (N_16740,N_15949,N_15734);
xnor U16741 (N_16741,N_15862,N_16006);
and U16742 (N_16742,N_15666,N_15862);
nor U16743 (N_16743,N_16152,N_15988);
nor U16744 (N_16744,N_16002,N_15868);
xor U16745 (N_16745,N_16134,N_16078);
xnor U16746 (N_16746,N_16230,N_15674);
xor U16747 (N_16747,N_16082,N_16110);
nor U16748 (N_16748,N_15777,N_15994);
or U16749 (N_16749,N_15959,N_15990);
nor U16750 (N_16750,N_16111,N_16199);
xnor U16751 (N_16751,N_15962,N_15990);
nor U16752 (N_16752,N_16220,N_15872);
nor U16753 (N_16753,N_15867,N_15921);
or U16754 (N_16754,N_16065,N_15641);
nand U16755 (N_16755,N_15716,N_15625);
nand U16756 (N_16756,N_15868,N_15645);
xor U16757 (N_16757,N_15681,N_15923);
and U16758 (N_16758,N_16183,N_15823);
and U16759 (N_16759,N_16083,N_15773);
xor U16760 (N_16760,N_15789,N_15878);
nand U16761 (N_16761,N_16040,N_16071);
nor U16762 (N_16762,N_15846,N_16147);
and U16763 (N_16763,N_16138,N_15843);
xnor U16764 (N_16764,N_16203,N_16132);
xor U16765 (N_16765,N_15857,N_15676);
or U16766 (N_16766,N_15931,N_16053);
nand U16767 (N_16767,N_15957,N_15779);
nand U16768 (N_16768,N_16075,N_16091);
or U16769 (N_16769,N_15989,N_15687);
nand U16770 (N_16770,N_15635,N_16238);
xnor U16771 (N_16771,N_15920,N_15982);
or U16772 (N_16772,N_15846,N_15923);
or U16773 (N_16773,N_16135,N_15772);
nor U16774 (N_16774,N_15728,N_15796);
and U16775 (N_16775,N_16198,N_15984);
nor U16776 (N_16776,N_16129,N_15828);
nor U16777 (N_16777,N_15962,N_15743);
nand U16778 (N_16778,N_16104,N_15951);
xor U16779 (N_16779,N_15973,N_15635);
xnor U16780 (N_16780,N_15994,N_15883);
nor U16781 (N_16781,N_15909,N_16129);
or U16782 (N_16782,N_16242,N_15918);
and U16783 (N_16783,N_15858,N_16045);
nor U16784 (N_16784,N_15791,N_15836);
xnor U16785 (N_16785,N_16002,N_15668);
or U16786 (N_16786,N_16195,N_15648);
or U16787 (N_16787,N_16018,N_15957);
and U16788 (N_16788,N_15774,N_15800);
xnor U16789 (N_16789,N_15813,N_15993);
xnor U16790 (N_16790,N_16026,N_15967);
nand U16791 (N_16791,N_16018,N_16183);
and U16792 (N_16792,N_15888,N_16058);
nor U16793 (N_16793,N_15788,N_15647);
xor U16794 (N_16794,N_16225,N_15836);
xnor U16795 (N_16795,N_16019,N_15748);
xor U16796 (N_16796,N_15642,N_15901);
nand U16797 (N_16797,N_16248,N_15628);
or U16798 (N_16798,N_15757,N_16225);
or U16799 (N_16799,N_16015,N_16150);
or U16800 (N_16800,N_15738,N_16024);
and U16801 (N_16801,N_16086,N_16127);
nand U16802 (N_16802,N_15974,N_16231);
nand U16803 (N_16803,N_15781,N_16204);
xnor U16804 (N_16804,N_15916,N_16007);
xor U16805 (N_16805,N_16095,N_15954);
nand U16806 (N_16806,N_15678,N_16008);
and U16807 (N_16807,N_15936,N_15814);
or U16808 (N_16808,N_16070,N_16212);
nor U16809 (N_16809,N_16082,N_16034);
and U16810 (N_16810,N_16174,N_16185);
or U16811 (N_16811,N_15765,N_16206);
nand U16812 (N_16812,N_15629,N_15914);
and U16813 (N_16813,N_15991,N_16036);
and U16814 (N_16814,N_16035,N_15992);
nand U16815 (N_16815,N_15798,N_15873);
xnor U16816 (N_16816,N_16100,N_16085);
nand U16817 (N_16817,N_15673,N_15976);
nand U16818 (N_16818,N_16249,N_16085);
and U16819 (N_16819,N_16178,N_15842);
or U16820 (N_16820,N_16186,N_16085);
or U16821 (N_16821,N_16106,N_16233);
nor U16822 (N_16822,N_15641,N_16190);
and U16823 (N_16823,N_16247,N_15990);
or U16824 (N_16824,N_16097,N_15846);
and U16825 (N_16825,N_16087,N_16033);
or U16826 (N_16826,N_15713,N_15660);
and U16827 (N_16827,N_16179,N_15968);
or U16828 (N_16828,N_15748,N_15847);
xor U16829 (N_16829,N_15933,N_16224);
nor U16830 (N_16830,N_15845,N_15911);
and U16831 (N_16831,N_15698,N_16167);
xor U16832 (N_16832,N_16056,N_15785);
xnor U16833 (N_16833,N_15920,N_15640);
xnor U16834 (N_16834,N_16115,N_15631);
nand U16835 (N_16835,N_16092,N_15627);
or U16836 (N_16836,N_15940,N_15794);
nand U16837 (N_16837,N_15828,N_15991);
or U16838 (N_16838,N_15853,N_15830);
or U16839 (N_16839,N_15957,N_16159);
xnor U16840 (N_16840,N_15711,N_15644);
nand U16841 (N_16841,N_15907,N_15888);
and U16842 (N_16842,N_15785,N_16009);
xnor U16843 (N_16843,N_15640,N_16235);
and U16844 (N_16844,N_15709,N_16104);
nand U16845 (N_16845,N_15915,N_16196);
nor U16846 (N_16846,N_15814,N_15963);
or U16847 (N_16847,N_15808,N_16211);
nor U16848 (N_16848,N_16217,N_16174);
nand U16849 (N_16849,N_15678,N_16021);
nand U16850 (N_16850,N_15811,N_16236);
nand U16851 (N_16851,N_16012,N_15651);
nand U16852 (N_16852,N_15742,N_15669);
and U16853 (N_16853,N_16095,N_15757);
xnor U16854 (N_16854,N_15949,N_15926);
xnor U16855 (N_16855,N_15959,N_15674);
or U16856 (N_16856,N_16224,N_15956);
nand U16857 (N_16857,N_16031,N_15794);
or U16858 (N_16858,N_15999,N_15859);
xnor U16859 (N_16859,N_15937,N_15683);
or U16860 (N_16860,N_16207,N_16249);
nand U16861 (N_16861,N_15684,N_15794);
xnor U16862 (N_16862,N_16076,N_15669);
xnor U16863 (N_16863,N_16228,N_16072);
nor U16864 (N_16864,N_15759,N_15665);
xor U16865 (N_16865,N_15933,N_16115);
xor U16866 (N_16866,N_15656,N_15807);
nor U16867 (N_16867,N_15730,N_16231);
nor U16868 (N_16868,N_15749,N_15732);
and U16869 (N_16869,N_15821,N_15699);
and U16870 (N_16870,N_16204,N_15820);
or U16871 (N_16871,N_15638,N_16210);
nor U16872 (N_16872,N_15965,N_16197);
and U16873 (N_16873,N_15815,N_15951);
or U16874 (N_16874,N_16248,N_15900);
xor U16875 (N_16875,N_16849,N_16692);
and U16876 (N_16876,N_16771,N_16669);
or U16877 (N_16877,N_16678,N_16674);
xnor U16878 (N_16878,N_16699,N_16368);
xor U16879 (N_16879,N_16333,N_16540);
and U16880 (N_16880,N_16837,N_16461);
and U16881 (N_16881,N_16677,N_16450);
and U16882 (N_16882,N_16797,N_16606);
or U16883 (N_16883,N_16836,N_16256);
and U16884 (N_16884,N_16719,N_16639);
nand U16885 (N_16885,N_16277,N_16658);
and U16886 (N_16886,N_16703,N_16482);
xor U16887 (N_16887,N_16613,N_16300);
and U16888 (N_16888,N_16637,N_16360);
and U16889 (N_16889,N_16352,N_16727);
nand U16890 (N_16890,N_16321,N_16496);
or U16891 (N_16891,N_16254,N_16251);
nand U16892 (N_16892,N_16303,N_16745);
and U16893 (N_16893,N_16460,N_16549);
nand U16894 (N_16894,N_16769,N_16710);
and U16895 (N_16895,N_16817,N_16630);
and U16896 (N_16896,N_16825,N_16681);
xnor U16897 (N_16897,N_16497,N_16708);
and U16898 (N_16898,N_16426,N_16605);
and U16899 (N_16899,N_16400,N_16591);
nand U16900 (N_16900,N_16583,N_16468);
xnor U16901 (N_16901,N_16868,N_16272);
or U16902 (N_16902,N_16279,N_16622);
or U16903 (N_16903,N_16255,N_16419);
and U16904 (N_16904,N_16379,N_16484);
xor U16905 (N_16905,N_16268,N_16447);
and U16906 (N_16906,N_16594,N_16494);
xnor U16907 (N_16907,N_16388,N_16705);
or U16908 (N_16908,N_16507,N_16476);
nand U16909 (N_16909,N_16404,N_16690);
and U16910 (N_16910,N_16571,N_16487);
nor U16911 (N_16911,N_16269,N_16773);
or U16912 (N_16912,N_16418,N_16713);
nor U16913 (N_16913,N_16304,N_16676);
nand U16914 (N_16914,N_16364,N_16357);
or U16915 (N_16915,N_16252,N_16545);
or U16916 (N_16916,N_16414,N_16626);
or U16917 (N_16917,N_16832,N_16638);
nor U16918 (N_16918,N_16307,N_16532);
xor U16919 (N_16919,N_16409,N_16642);
or U16920 (N_16920,N_16790,N_16467);
xor U16921 (N_16921,N_16804,N_16577);
xor U16922 (N_16922,N_16818,N_16266);
and U16923 (N_16923,N_16310,N_16761);
or U16924 (N_16924,N_16471,N_16595);
xor U16925 (N_16925,N_16442,N_16617);
or U16926 (N_16926,N_16864,N_16709);
xor U16927 (N_16927,N_16643,N_16263);
and U16928 (N_16928,N_16866,N_16353);
xnor U16929 (N_16929,N_16558,N_16556);
and U16930 (N_16930,N_16776,N_16566);
or U16931 (N_16931,N_16351,N_16329);
or U16932 (N_16932,N_16589,N_16309);
and U16933 (N_16933,N_16679,N_16371);
or U16934 (N_16934,N_16750,N_16423);
nor U16935 (N_16935,N_16367,N_16632);
nor U16936 (N_16936,N_16501,N_16311);
nand U16937 (N_16937,N_16616,N_16520);
or U16938 (N_16938,N_16809,N_16847);
or U16939 (N_16939,N_16446,N_16281);
or U16940 (N_16940,N_16671,N_16253);
nand U16941 (N_16941,N_16607,N_16573);
nor U16942 (N_16942,N_16402,N_16539);
nor U16943 (N_16943,N_16493,N_16298);
nand U16944 (N_16944,N_16738,N_16387);
nand U16945 (N_16945,N_16465,N_16728);
and U16946 (N_16946,N_16601,N_16778);
or U16947 (N_16947,N_16814,N_16726);
xnor U16948 (N_16948,N_16722,N_16801);
xor U16949 (N_16949,N_16731,N_16555);
xnor U16950 (N_16950,N_16609,N_16410);
and U16951 (N_16951,N_16844,N_16324);
and U16952 (N_16952,N_16634,N_16546);
xor U16953 (N_16953,N_16748,N_16313);
nor U16954 (N_16954,N_16628,N_16625);
nor U16955 (N_16955,N_16859,N_16752);
nand U16956 (N_16956,N_16853,N_16820);
nor U16957 (N_16957,N_16373,N_16541);
xor U16958 (N_16958,N_16598,N_16720);
nand U16959 (N_16959,N_16537,N_16342);
xor U16960 (N_16960,N_16302,N_16506);
and U16961 (N_16961,N_16308,N_16448);
or U16962 (N_16962,N_16723,N_16327);
xnor U16963 (N_16963,N_16798,N_16624);
nand U16964 (N_16964,N_16502,N_16840);
and U16965 (N_16965,N_16438,N_16366);
nand U16966 (N_16966,N_16258,N_16375);
nor U16967 (N_16967,N_16664,N_16764);
or U16968 (N_16968,N_16547,N_16629);
nor U16969 (N_16969,N_16276,N_16821);
xor U16970 (N_16970,N_16829,N_16401);
and U16971 (N_16971,N_16271,N_16680);
nand U16972 (N_16972,N_16384,N_16485);
xnor U16973 (N_16973,N_16785,N_16359);
and U16974 (N_16974,N_16376,N_16759);
and U16975 (N_16975,N_16667,N_16766);
nand U16976 (N_16976,N_16570,N_16662);
and U16977 (N_16977,N_16744,N_16619);
and U16978 (N_16978,N_16633,N_16848);
nand U16979 (N_16979,N_16348,N_16683);
nor U16980 (N_16980,N_16795,N_16312);
nand U16981 (N_16981,N_16441,N_16445);
nand U16982 (N_16982,N_16433,N_16466);
or U16983 (N_16983,N_16623,N_16783);
and U16984 (N_16984,N_16697,N_16597);
or U16985 (N_16985,N_16620,N_16429);
nor U16986 (N_16986,N_16526,N_16346);
and U16987 (N_16987,N_16582,N_16542);
nor U16988 (N_16988,N_16294,N_16530);
xnor U16989 (N_16989,N_16655,N_16415);
nand U16990 (N_16990,N_16645,N_16479);
nor U16991 (N_16991,N_16337,N_16296);
nand U16992 (N_16992,N_16464,N_16574);
nor U16993 (N_16993,N_16686,N_16650);
nor U16994 (N_16994,N_16335,N_16666);
xnor U16995 (N_16995,N_16627,N_16865);
and U16996 (N_16996,N_16757,N_16792);
nor U16997 (N_16997,N_16845,N_16751);
xnor U16998 (N_16998,N_16872,N_16284);
and U16999 (N_16999,N_16793,N_16331);
and U17000 (N_17000,N_16397,N_16406);
nand U17001 (N_17001,N_16320,N_16405);
or U17002 (N_17002,N_16382,N_16819);
or U17003 (N_17003,N_16283,N_16280);
xnor U17004 (N_17004,N_16481,N_16578);
xor U17005 (N_17005,N_16521,N_16693);
xor U17006 (N_17006,N_16610,N_16259);
or U17007 (N_17007,N_16552,N_16668);
and U17008 (N_17008,N_16857,N_16670);
nand U17009 (N_17009,N_16694,N_16575);
nand U17010 (N_17010,N_16843,N_16512);
nor U17011 (N_17011,N_16444,N_16528);
nor U17012 (N_17012,N_16338,N_16685);
or U17013 (N_17013,N_16398,N_16740);
xnor U17014 (N_17014,N_16553,N_16816);
xnor U17015 (N_17015,N_16656,N_16343);
nor U17016 (N_17016,N_16863,N_16381);
xor U17017 (N_17017,N_16858,N_16636);
xnor U17018 (N_17018,N_16784,N_16569);
nor U17019 (N_17019,N_16470,N_16873);
xor U17020 (N_17020,N_16608,N_16808);
or U17021 (N_17021,N_16392,N_16399);
xnor U17022 (N_17022,N_16260,N_16615);
and U17023 (N_17023,N_16533,N_16449);
nor U17024 (N_17024,N_16370,N_16391);
xor U17025 (N_17025,N_16250,N_16531);
and U17026 (N_17026,N_16417,N_16475);
or U17027 (N_17027,N_16285,N_16517);
and U17028 (N_17028,N_16275,N_16377);
xor U17029 (N_17029,N_16644,N_16319);
nor U17030 (N_17030,N_16695,N_16839);
nor U17031 (N_17031,N_16505,N_16649);
nor U17032 (N_17032,N_16647,N_16716);
or U17033 (N_17033,N_16763,N_16805);
and U17034 (N_17034,N_16557,N_16600);
and U17035 (N_17035,N_16653,N_16301);
nor U17036 (N_17036,N_16860,N_16767);
and U17037 (N_17037,N_16344,N_16499);
and U17038 (N_17038,N_16869,N_16780);
xnor U17039 (N_17039,N_16704,N_16336);
xnor U17040 (N_17040,N_16513,N_16394);
or U17041 (N_17041,N_16463,N_16349);
and U17042 (N_17042,N_16721,N_16328);
nand U17043 (N_17043,N_16456,N_16746);
or U17044 (N_17044,N_16599,N_16440);
nor U17045 (N_17045,N_16715,N_16584);
nand U17046 (N_17046,N_16295,N_16424);
nand U17047 (N_17047,N_16282,N_16604);
nand U17048 (N_17048,N_16459,N_16831);
and U17049 (N_17049,N_16455,N_16529);
nor U17050 (N_17050,N_16407,N_16551);
or U17051 (N_17051,N_16462,N_16828);
nand U17052 (N_17052,N_16374,N_16563);
xor U17053 (N_17053,N_16457,N_16714);
and U17054 (N_17054,N_16453,N_16325);
nor U17055 (N_17055,N_16305,N_16706);
xnor U17056 (N_17056,N_16510,N_16492);
nand U17057 (N_17057,N_16389,N_16372);
or U17058 (N_17058,N_16742,N_16754);
or U17059 (N_17059,N_16514,N_16518);
nand U17060 (N_17060,N_16810,N_16472);
xor U17061 (N_17061,N_16432,N_16561);
nor U17062 (N_17062,N_16454,N_16293);
or U17063 (N_17063,N_16593,N_16490);
and U17064 (N_17064,N_16538,N_16807);
and U17065 (N_17065,N_16760,N_16508);
or U17066 (N_17066,N_16729,N_16422);
nand U17067 (N_17067,N_16425,N_16576);
and U17068 (N_17068,N_16408,N_16443);
nor U17069 (N_17069,N_16824,N_16675);
nand U17070 (N_17070,N_16846,N_16567);
or U17071 (N_17071,N_16564,N_16291);
nor U17072 (N_17072,N_16548,N_16356);
xor U17073 (N_17073,N_16856,N_16306);
and U17074 (N_17074,N_16473,N_16646);
nor U17075 (N_17075,N_16842,N_16749);
and U17076 (N_17076,N_16559,N_16395);
and U17077 (N_17077,N_16786,N_16322);
nand U17078 (N_17078,N_16581,N_16725);
xnor U17079 (N_17079,N_16830,N_16289);
nand U17080 (N_17080,N_16736,N_16550);
nor U17081 (N_17081,N_16660,N_16318);
xnor U17082 (N_17082,N_16635,N_16515);
xor U17083 (N_17083,N_16522,N_16823);
nand U17084 (N_17084,N_16469,N_16451);
nand U17085 (N_17085,N_16815,N_16516);
nor U17086 (N_17086,N_16486,N_16700);
or U17087 (N_17087,N_16698,N_16588);
nand U17088 (N_17088,N_16596,N_16874);
or U17089 (N_17089,N_16592,N_16796);
and U17090 (N_17090,N_16527,N_16534);
xnor U17091 (N_17091,N_16621,N_16772);
xnor U17092 (N_17092,N_16315,N_16524);
and U17093 (N_17093,N_16264,N_16437);
nor U17094 (N_17094,N_16436,N_16354);
xnor U17095 (N_17095,N_16385,N_16568);
or U17096 (N_17096,N_16416,N_16488);
or U17097 (N_17097,N_16519,N_16758);
nand U17098 (N_17098,N_16412,N_16452);
and U17099 (N_17099,N_16345,N_16383);
xor U17100 (N_17100,N_16386,N_16587);
and U17101 (N_17101,N_16687,N_16743);
and U17102 (N_17102,N_16411,N_16503);
xnor U17103 (N_17103,N_16586,N_16270);
xor U17104 (N_17104,N_16737,N_16314);
nor U17105 (N_17105,N_16332,N_16317);
nand U17106 (N_17106,N_16560,N_16782);
xor U17107 (N_17107,N_16326,N_16851);
xor U17108 (N_17108,N_16340,N_16612);
or U17109 (N_17109,N_16525,N_16811);
or U17110 (N_17110,N_16862,N_16702);
or U17111 (N_17111,N_16717,N_16286);
nor U17112 (N_17112,N_16711,N_16355);
xnor U17113 (N_17113,N_16396,N_16585);
nor U17114 (N_17114,N_16835,N_16491);
or U17115 (N_17115,N_16822,N_16762);
and U17116 (N_17116,N_16287,N_16421);
xor U17117 (N_17117,N_16659,N_16274);
nor U17118 (N_17118,N_16739,N_16565);
or U17119 (N_17119,N_16439,N_16362);
or U17120 (N_17120,N_16339,N_16813);
or U17121 (N_17121,N_16834,N_16267);
nand U17122 (N_17122,N_16509,N_16614);
xnor U17123 (N_17123,N_16273,N_16827);
and U17124 (N_17124,N_16265,N_16673);
nand U17125 (N_17125,N_16435,N_16779);
nand U17126 (N_17126,N_16631,N_16755);
nor U17127 (N_17127,N_16707,N_16734);
or U17128 (N_17128,N_16572,N_16768);
and U17129 (N_17129,N_16350,N_16618);
and U17130 (N_17130,N_16543,N_16718);
and U17131 (N_17131,N_16536,N_16870);
nor U17132 (N_17132,N_16765,N_16806);
and U17133 (N_17133,N_16652,N_16641);
nand U17134 (N_17134,N_16257,N_16458);
nand U17135 (N_17135,N_16500,N_16347);
or U17136 (N_17136,N_16489,N_16504);
xor U17137 (N_17137,N_16661,N_16741);
and U17138 (N_17138,N_16278,N_16365);
nand U17139 (N_17139,N_16420,N_16403);
xor U17140 (N_17140,N_16774,N_16833);
or U17141 (N_17141,N_16554,N_16781);
nand U17142 (N_17142,N_16800,N_16602);
and U17143 (N_17143,N_16477,N_16361);
xor U17144 (N_17144,N_16334,N_16724);
nor U17145 (N_17145,N_16299,N_16871);
or U17146 (N_17146,N_16495,N_16611);
or U17147 (N_17147,N_16434,N_16789);
or U17148 (N_17148,N_16640,N_16735);
xnor U17149 (N_17149,N_16483,N_16380);
and U17150 (N_17150,N_16787,N_16867);
xor U17151 (N_17151,N_16684,N_16288);
nand U17152 (N_17152,N_16297,N_16733);
or U17153 (N_17153,N_16430,N_16788);
and U17154 (N_17154,N_16369,N_16657);
and U17155 (N_17155,N_16753,N_16855);
nor U17156 (N_17156,N_16544,N_16651);
and U17157 (N_17157,N_16648,N_16791);
nor U17158 (N_17158,N_16672,N_16850);
nand U17159 (N_17159,N_16691,N_16794);
nor U17160 (N_17160,N_16330,N_16696);
or U17161 (N_17161,N_16654,N_16802);
nor U17162 (N_17162,N_16730,N_16701);
xor U17163 (N_17163,N_16262,N_16590);
nand U17164 (N_17164,N_16363,N_16812);
nand U17165 (N_17165,N_16854,N_16290);
and U17166 (N_17166,N_16838,N_16562);
nand U17167 (N_17167,N_16480,N_16603);
and U17168 (N_17168,N_16682,N_16841);
or U17169 (N_17169,N_16523,N_16535);
or U17170 (N_17170,N_16474,N_16292);
or U17171 (N_17171,N_16358,N_16393);
and U17172 (N_17172,N_16323,N_16478);
nor U17173 (N_17173,N_16428,N_16511);
or U17174 (N_17174,N_16390,N_16777);
xor U17175 (N_17175,N_16861,N_16579);
nor U17176 (N_17176,N_16663,N_16770);
xor U17177 (N_17177,N_16427,N_16413);
or U17178 (N_17178,N_16756,N_16826);
and U17179 (N_17179,N_16378,N_16747);
and U17180 (N_17180,N_16431,N_16852);
xnor U17181 (N_17181,N_16580,N_16316);
nor U17182 (N_17182,N_16665,N_16775);
xor U17183 (N_17183,N_16803,N_16799);
or U17184 (N_17184,N_16689,N_16341);
nor U17185 (N_17185,N_16688,N_16498);
nand U17186 (N_17186,N_16712,N_16261);
and U17187 (N_17187,N_16732,N_16532);
nand U17188 (N_17188,N_16766,N_16852);
nor U17189 (N_17189,N_16516,N_16751);
nand U17190 (N_17190,N_16626,N_16465);
or U17191 (N_17191,N_16536,N_16813);
nor U17192 (N_17192,N_16794,N_16476);
and U17193 (N_17193,N_16345,N_16627);
or U17194 (N_17194,N_16616,N_16409);
or U17195 (N_17195,N_16870,N_16689);
xor U17196 (N_17196,N_16330,N_16784);
and U17197 (N_17197,N_16558,N_16304);
nand U17198 (N_17198,N_16830,N_16622);
or U17199 (N_17199,N_16341,N_16776);
xor U17200 (N_17200,N_16727,N_16759);
xor U17201 (N_17201,N_16426,N_16656);
nor U17202 (N_17202,N_16403,N_16615);
and U17203 (N_17203,N_16508,N_16654);
xor U17204 (N_17204,N_16741,N_16292);
and U17205 (N_17205,N_16533,N_16334);
or U17206 (N_17206,N_16462,N_16408);
nor U17207 (N_17207,N_16512,N_16742);
nand U17208 (N_17208,N_16361,N_16835);
xnor U17209 (N_17209,N_16744,N_16282);
and U17210 (N_17210,N_16874,N_16409);
xor U17211 (N_17211,N_16628,N_16296);
and U17212 (N_17212,N_16479,N_16405);
nand U17213 (N_17213,N_16271,N_16436);
nand U17214 (N_17214,N_16840,N_16825);
and U17215 (N_17215,N_16775,N_16291);
xnor U17216 (N_17216,N_16361,N_16471);
xor U17217 (N_17217,N_16504,N_16556);
and U17218 (N_17218,N_16263,N_16461);
nand U17219 (N_17219,N_16483,N_16682);
nand U17220 (N_17220,N_16738,N_16841);
nor U17221 (N_17221,N_16594,N_16530);
xor U17222 (N_17222,N_16771,N_16706);
and U17223 (N_17223,N_16844,N_16834);
nor U17224 (N_17224,N_16819,N_16514);
or U17225 (N_17225,N_16321,N_16444);
nor U17226 (N_17226,N_16710,N_16295);
nand U17227 (N_17227,N_16356,N_16271);
and U17228 (N_17228,N_16429,N_16411);
nor U17229 (N_17229,N_16687,N_16322);
and U17230 (N_17230,N_16556,N_16300);
nor U17231 (N_17231,N_16556,N_16365);
or U17232 (N_17232,N_16680,N_16610);
or U17233 (N_17233,N_16624,N_16303);
nand U17234 (N_17234,N_16609,N_16456);
xor U17235 (N_17235,N_16447,N_16789);
nand U17236 (N_17236,N_16712,N_16476);
and U17237 (N_17237,N_16804,N_16433);
nor U17238 (N_17238,N_16376,N_16256);
or U17239 (N_17239,N_16619,N_16323);
nor U17240 (N_17240,N_16440,N_16278);
and U17241 (N_17241,N_16690,N_16693);
nand U17242 (N_17242,N_16264,N_16520);
nand U17243 (N_17243,N_16607,N_16278);
nand U17244 (N_17244,N_16652,N_16284);
and U17245 (N_17245,N_16322,N_16774);
xnor U17246 (N_17246,N_16715,N_16717);
and U17247 (N_17247,N_16413,N_16865);
and U17248 (N_17248,N_16422,N_16255);
or U17249 (N_17249,N_16534,N_16817);
or U17250 (N_17250,N_16851,N_16353);
and U17251 (N_17251,N_16301,N_16472);
or U17252 (N_17252,N_16303,N_16361);
or U17253 (N_17253,N_16497,N_16326);
nand U17254 (N_17254,N_16781,N_16448);
and U17255 (N_17255,N_16417,N_16368);
nand U17256 (N_17256,N_16269,N_16842);
xor U17257 (N_17257,N_16865,N_16319);
and U17258 (N_17258,N_16466,N_16711);
or U17259 (N_17259,N_16491,N_16599);
or U17260 (N_17260,N_16635,N_16311);
nor U17261 (N_17261,N_16764,N_16573);
nand U17262 (N_17262,N_16758,N_16656);
and U17263 (N_17263,N_16428,N_16707);
nor U17264 (N_17264,N_16702,N_16651);
nor U17265 (N_17265,N_16346,N_16590);
xor U17266 (N_17266,N_16273,N_16744);
nand U17267 (N_17267,N_16524,N_16357);
nand U17268 (N_17268,N_16315,N_16534);
nor U17269 (N_17269,N_16852,N_16270);
and U17270 (N_17270,N_16770,N_16640);
nand U17271 (N_17271,N_16422,N_16786);
nor U17272 (N_17272,N_16658,N_16300);
or U17273 (N_17273,N_16654,N_16753);
and U17274 (N_17274,N_16274,N_16806);
or U17275 (N_17275,N_16305,N_16264);
nand U17276 (N_17276,N_16290,N_16664);
xor U17277 (N_17277,N_16532,N_16865);
nor U17278 (N_17278,N_16328,N_16377);
nor U17279 (N_17279,N_16724,N_16483);
nor U17280 (N_17280,N_16665,N_16376);
nor U17281 (N_17281,N_16748,N_16467);
and U17282 (N_17282,N_16814,N_16282);
nor U17283 (N_17283,N_16625,N_16785);
nand U17284 (N_17284,N_16594,N_16689);
nor U17285 (N_17285,N_16798,N_16722);
xnor U17286 (N_17286,N_16531,N_16327);
xnor U17287 (N_17287,N_16745,N_16701);
or U17288 (N_17288,N_16431,N_16853);
or U17289 (N_17289,N_16275,N_16784);
nor U17290 (N_17290,N_16284,N_16735);
or U17291 (N_17291,N_16570,N_16791);
nor U17292 (N_17292,N_16783,N_16724);
nor U17293 (N_17293,N_16311,N_16866);
and U17294 (N_17294,N_16705,N_16435);
nor U17295 (N_17295,N_16555,N_16680);
xnor U17296 (N_17296,N_16391,N_16831);
and U17297 (N_17297,N_16486,N_16676);
or U17298 (N_17298,N_16498,N_16796);
and U17299 (N_17299,N_16729,N_16308);
or U17300 (N_17300,N_16672,N_16607);
nor U17301 (N_17301,N_16773,N_16432);
nor U17302 (N_17302,N_16821,N_16777);
nand U17303 (N_17303,N_16523,N_16768);
nand U17304 (N_17304,N_16725,N_16682);
nor U17305 (N_17305,N_16645,N_16625);
xnor U17306 (N_17306,N_16441,N_16594);
and U17307 (N_17307,N_16535,N_16310);
or U17308 (N_17308,N_16287,N_16471);
nor U17309 (N_17309,N_16338,N_16766);
nand U17310 (N_17310,N_16381,N_16516);
and U17311 (N_17311,N_16287,N_16725);
xor U17312 (N_17312,N_16578,N_16670);
xnor U17313 (N_17313,N_16562,N_16369);
or U17314 (N_17314,N_16628,N_16680);
nor U17315 (N_17315,N_16821,N_16689);
xor U17316 (N_17316,N_16558,N_16780);
nor U17317 (N_17317,N_16657,N_16822);
xor U17318 (N_17318,N_16350,N_16756);
or U17319 (N_17319,N_16648,N_16578);
and U17320 (N_17320,N_16374,N_16368);
or U17321 (N_17321,N_16703,N_16347);
or U17322 (N_17322,N_16457,N_16849);
nand U17323 (N_17323,N_16776,N_16522);
or U17324 (N_17324,N_16545,N_16526);
or U17325 (N_17325,N_16316,N_16638);
or U17326 (N_17326,N_16605,N_16811);
or U17327 (N_17327,N_16481,N_16572);
nand U17328 (N_17328,N_16460,N_16714);
or U17329 (N_17329,N_16427,N_16335);
and U17330 (N_17330,N_16421,N_16609);
nor U17331 (N_17331,N_16699,N_16267);
nand U17332 (N_17332,N_16262,N_16664);
xnor U17333 (N_17333,N_16334,N_16457);
nor U17334 (N_17334,N_16664,N_16763);
or U17335 (N_17335,N_16280,N_16321);
nor U17336 (N_17336,N_16821,N_16671);
xnor U17337 (N_17337,N_16421,N_16747);
xnor U17338 (N_17338,N_16733,N_16870);
nor U17339 (N_17339,N_16564,N_16422);
or U17340 (N_17340,N_16731,N_16420);
xnor U17341 (N_17341,N_16733,N_16455);
nand U17342 (N_17342,N_16368,N_16777);
xor U17343 (N_17343,N_16665,N_16536);
nor U17344 (N_17344,N_16472,N_16706);
nand U17345 (N_17345,N_16838,N_16640);
or U17346 (N_17346,N_16365,N_16371);
and U17347 (N_17347,N_16668,N_16276);
nand U17348 (N_17348,N_16454,N_16703);
nor U17349 (N_17349,N_16265,N_16300);
or U17350 (N_17350,N_16587,N_16394);
and U17351 (N_17351,N_16340,N_16643);
and U17352 (N_17352,N_16723,N_16268);
nand U17353 (N_17353,N_16831,N_16657);
nand U17354 (N_17354,N_16572,N_16403);
nand U17355 (N_17355,N_16584,N_16347);
or U17356 (N_17356,N_16870,N_16863);
nor U17357 (N_17357,N_16568,N_16744);
and U17358 (N_17358,N_16383,N_16446);
nor U17359 (N_17359,N_16401,N_16734);
nor U17360 (N_17360,N_16434,N_16689);
or U17361 (N_17361,N_16269,N_16445);
xor U17362 (N_17362,N_16566,N_16419);
and U17363 (N_17363,N_16467,N_16609);
nor U17364 (N_17364,N_16375,N_16607);
nor U17365 (N_17365,N_16710,N_16453);
or U17366 (N_17366,N_16537,N_16633);
nand U17367 (N_17367,N_16347,N_16553);
nor U17368 (N_17368,N_16587,N_16465);
or U17369 (N_17369,N_16376,N_16443);
or U17370 (N_17370,N_16531,N_16361);
or U17371 (N_17371,N_16393,N_16611);
xnor U17372 (N_17372,N_16816,N_16289);
nor U17373 (N_17373,N_16561,N_16534);
xnor U17374 (N_17374,N_16395,N_16625);
and U17375 (N_17375,N_16870,N_16706);
nand U17376 (N_17376,N_16719,N_16366);
nand U17377 (N_17377,N_16431,N_16543);
nand U17378 (N_17378,N_16551,N_16338);
xor U17379 (N_17379,N_16848,N_16838);
or U17380 (N_17380,N_16785,N_16763);
nand U17381 (N_17381,N_16655,N_16783);
xnor U17382 (N_17382,N_16287,N_16502);
xnor U17383 (N_17383,N_16597,N_16630);
nand U17384 (N_17384,N_16664,N_16311);
xor U17385 (N_17385,N_16604,N_16779);
or U17386 (N_17386,N_16467,N_16824);
nand U17387 (N_17387,N_16785,N_16566);
nor U17388 (N_17388,N_16387,N_16328);
nand U17389 (N_17389,N_16252,N_16278);
xnor U17390 (N_17390,N_16434,N_16748);
or U17391 (N_17391,N_16775,N_16633);
and U17392 (N_17392,N_16494,N_16402);
and U17393 (N_17393,N_16515,N_16820);
nor U17394 (N_17394,N_16264,N_16409);
and U17395 (N_17395,N_16704,N_16307);
and U17396 (N_17396,N_16802,N_16861);
and U17397 (N_17397,N_16751,N_16816);
xor U17398 (N_17398,N_16447,N_16563);
nor U17399 (N_17399,N_16364,N_16407);
and U17400 (N_17400,N_16401,N_16717);
and U17401 (N_17401,N_16813,N_16312);
and U17402 (N_17402,N_16560,N_16419);
and U17403 (N_17403,N_16307,N_16769);
nand U17404 (N_17404,N_16758,N_16612);
xnor U17405 (N_17405,N_16269,N_16319);
xor U17406 (N_17406,N_16554,N_16569);
nor U17407 (N_17407,N_16511,N_16672);
and U17408 (N_17408,N_16387,N_16310);
and U17409 (N_17409,N_16621,N_16551);
or U17410 (N_17410,N_16727,N_16635);
xnor U17411 (N_17411,N_16271,N_16833);
nand U17412 (N_17412,N_16599,N_16612);
nor U17413 (N_17413,N_16673,N_16264);
nand U17414 (N_17414,N_16873,N_16493);
nor U17415 (N_17415,N_16311,N_16781);
xnor U17416 (N_17416,N_16428,N_16496);
xnor U17417 (N_17417,N_16454,N_16570);
nand U17418 (N_17418,N_16396,N_16615);
or U17419 (N_17419,N_16452,N_16415);
nand U17420 (N_17420,N_16535,N_16580);
or U17421 (N_17421,N_16387,N_16659);
xnor U17422 (N_17422,N_16826,N_16693);
nand U17423 (N_17423,N_16554,N_16324);
or U17424 (N_17424,N_16354,N_16542);
or U17425 (N_17425,N_16556,N_16873);
nand U17426 (N_17426,N_16787,N_16763);
or U17427 (N_17427,N_16439,N_16711);
nor U17428 (N_17428,N_16510,N_16301);
or U17429 (N_17429,N_16525,N_16504);
or U17430 (N_17430,N_16368,N_16756);
nor U17431 (N_17431,N_16448,N_16327);
xor U17432 (N_17432,N_16467,N_16481);
nor U17433 (N_17433,N_16396,N_16484);
nor U17434 (N_17434,N_16598,N_16336);
nand U17435 (N_17435,N_16704,N_16832);
xor U17436 (N_17436,N_16527,N_16325);
nor U17437 (N_17437,N_16323,N_16540);
xnor U17438 (N_17438,N_16334,N_16698);
and U17439 (N_17439,N_16420,N_16683);
nor U17440 (N_17440,N_16314,N_16759);
and U17441 (N_17441,N_16799,N_16437);
or U17442 (N_17442,N_16270,N_16525);
or U17443 (N_17443,N_16424,N_16420);
nand U17444 (N_17444,N_16347,N_16515);
nand U17445 (N_17445,N_16833,N_16691);
and U17446 (N_17446,N_16502,N_16750);
nor U17447 (N_17447,N_16395,N_16619);
and U17448 (N_17448,N_16832,N_16700);
nor U17449 (N_17449,N_16480,N_16756);
nor U17450 (N_17450,N_16702,N_16640);
or U17451 (N_17451,N_16636,N_16798);
nand U17452 (N_17452,N_16767,N_16662);
nand U17453 (N_17453,N_16857,N_16580);
xnor U17454 (N_17454,N_16656,N_16654);
and U17455 (N_17455,N_16578,N_16405);
nand U17456 (N_17456,N_16317,N_16584);
and U17457 (N_17457,N_16275,N_16762);
and U17458 (N_17458,N_16818,N_16323);
and U17459 (N_17459,N_16286,N_16825);
nor U17460 (N_17460,N_16503,N_16507);
xor U17461 (N_17461,N_16535,N_16819);
nor U17462 (N_17462,N_16852,N_16470);
xnor U17463 (N_17463,N_16746,N_16255);
and U17464 (N_17464,N_16578,N_16599);
and U17465 (N_17465,N_16657,N_16753);
and U17466 (N_17466,N_16638,N_16592);
nand U17467 (N_17467,N_16326,N_16304);
nand U17468 (N_17468,N_16667,N_16839);
and U17469 (N_17469,N_16260,N_16768);
nand U17470 (N_17470,N_16351,N_16620);
nor U17471 (N_17471,N_16650,N_16489);
nand U17472 (N_17472,N_16546,N_16859);
nor U17473 (N_17473,N_16874,N_16804);
nor U17474 (N_17474,N_16378,N_16356);
nor U17475 (N_17475,N_16510,N_16593);
nor U17476 (N_17476,N_16490,N_16401);
nand U17477 (N_17477,N_16498,N_16341);
and U17478 (N_17478,N_16694,N_16351);
or U17479 (N_17479,N_16675,N_16834);
and U17480 (N_17480,N_16406,N_16431);
or U17481 (N_17481,N_16709,N_16620);
and U17482 (N_17482,N_16418,N_16807);
and U17483 (N_17483,N_16755,N_16622);
or U17484 (N_17484,N_16310,N_16302);
nand U17485 (N_17485,N_16397,N_16795);
nor U17486 (N_17486,N_16444,N_16350);
and U17487 (N_17487,N_16616,N_16552);
xor U17488 (N_17488,N_16505,N_16531);
nor U17489 (N_17489,N_16720,N_16686);
nor U17490 (N_17490,N_16301,N_16855);
and U17491 (N_17491,N_16549,N_16530);
nor U17492 (N_17492,N_16561,N_16314);
nand U17493 (N_17493,N_16511,N_16367);
xor U17494 (N_17494,N_16557,N_16307);
and U17495 (N_17495,N_16534,N_16361);
nor U17496 (N_17496,N_16681,N_16283);
nand U17497 (N_17497,N_16574,N_16843);
nand U17498 (N_17498,N_16821,N_16395);
nor U17499 (N_17499,N_16657,N_16862);
nor U17500 (N_17500,N_16920,N_17201);
nor U17501 (N_17501,N_17022,N_17460);
nor U17502 (N_17502,N_17457,N_17048);
nand U17503 (N_17503,N_16955,N_17134);
nand U17504 (N_17504,N_17086,N_17316);
xor U17505 (N_17505,N_17055,N_17449);
nand U17506 (N_17506,N_17492,N_16974);
and U17507 (N_17507,N_17325,N_17049);
nor U17508 (N_17508,N_17102,N_17481);
and U17509 (N_17509,N_17373,N_17437);
nand U17510 (N_17510,N_16888,N_16892);
and U17511 (N_17511,N_17295,N_17137);
and U17512 (N_17512,N_17181,N_17307);
or U17513 (N_17513,N_17385,N_16942);
nor U17514 (N_17514,N_17497,N_17461);
nor U17515 (N_17515,N_17262,N_16970);
nor U17516 (N_17516,N_17265,N_16972);
nor U17517 (N_17517,N_17237,N_17165);
xnor U17518 (N_17518,N_17225,N_17231);
or U17519 (N_17519,N_17032,N_17442);
and U17520 (N_17520,N_17164,N_17254);
xnor U17521 (N_17521,N_17104,N_17489);
and U17522 (N_17522,N_16975,N_16880);
nor U17523 (N_17523,N_17339,N_17269);
or U17524 (N_17524,N_17112,N_16895);
and U17525 (N_17525,N_17259,N_16982);
xnor U17526 (N_17526,N_17235,N_16935);
xnor U17527 (N_17527,N_17143,N_17093);
nor U17528 (N_17528,N_17219,N_17127);
nand U17529 (N_17529,N_16945,N_17072);
and U17530 (N_17530,N_17266,N_17340);
and U17531 (N_17531,N_17178,N_17400);
and U17532 (N_17532,N_17308,N_17029);
xor U17533 (N_17533,N_16997,N_16907);
nor U17534 (N_17534,N_17183,N_17313);
and U17535 (N_17535,N_17470,N_17162);
or U17536 (N_17536,N_16959,N_17263);
xor U17537 (N_17537,N_16924,N_16979);
xnor U17538 (N_17538,N_16969,N_17484);
nand U17539 (N_17539,N_17478,N_17116);
nor U17540 (N_17540,N_16897,N_16887);
nand U17541 (N_17541,N_17364,N_17474);
nand U17542 (N_17542,N_16931,N_17079);
nand U17543 (N_17543,N_17311,N_17078);
nor U17544 (N_17544,N_17033,N_17320);
nor U17545 (N_17545,N_17499,N_17106);
or U17546 (N_17546,N_17190,N_16981);
nor U17547 (N_17547,N_17006,N_17180);
nand U17548 (N_17548,N_16909,N_16911);
or U17549 (N_17549,N_17192,N_17230);
nor U17550 (N_17550,N_17346,N_16906);
xor U17551 (N_17551,N_17184,N_17261);
or U17552 (N_17552,N_16899,N_17117);
and U17553 (N_17553,N_17063,N_17153);
nor U17554 (N_17554,N_17439,N_17351);
nand U17555 (N_17555,N_17448,N_17074);
and U17556 (N_17556,N_16923,N_17288);
or U17557 (N_17557,N_17120,N_17228);
and U17558 (N_17558,N_17089,N_17349);
and U17559 (N_17559,N_17473,N_17047);
xnor U17560 (N_17560,N_17174,N_17455);
nand U17561 (N_17561,N_17493,N_16876);
nor U17562 (N_17562,N_16886,N_17271);
xor U17563 (N_17563,N_17329,N_17430);
xor U17564 (N_17564,N_16990,N_17166);
nor U17565 (N_17565,N_17217,N_17186);
xor U17566 (N_17566,N_16878,N_17103);
nor U17567 (N_17567,N_17378,N_17065);
nor U17568 (N_17568,N_16958,N_17101);
and U17569 (N_17569,N_16904,N_17283);
xnor U17570 (N_17570,N_17030,N_17002);
nor U17571 (N_17571,N_17468,N_17393);
nand U17572 (N_17572,N_17368,N_17221);
xor U17573 (N_17573,N_17383,N_17163);
or U17574 (N_17574,N_16950,N_17429);
xor U17575 (N_17575,N_16996,N_17064);
or U17576 (N_17576,N_17399,N_16966);
or U17577 (N_17577,N_17396,N_17294);
xnor U17578 (N_17578,N_17077,N_17012);
nand U17579 (N_17579,N_17009,N_16929);
or U17580 (N_17580,N_16896,N_16927);
nor U17581 (N_17581,N_17130,N_17182);
and U17582 (N_17582,N_16949,N_17491);
xor U17583 (N_17583,N_17345,N_16995);
and U17584 (N_17584,N_17305,N_17110);
nor U17585 (N_17585,N_17152,N_17249);
nand U17586 (N_17586,N_17224,N_17234);
and U17587 (N_17587,N_17053,N_17046);
nand U17588 (N_17588,N_17148,N_17397);
or U17589 (N_17589,N_17095,N_17291);
nand U17590 (N_17590,N_17081,N_17125);
nand U17591 (N_17591,N_17350,N_16980);
or U17592 (N_17592,N_17475,N_17045);
nor U17593 (N_17593,N_17394,N_16940);
or U17594 (N_17594,N_16914,N_17435);
and U17595 (N_17595,N_17194,N_17222);
xor U17596 (N_17596,N_17278,N_17171);
nor U17597 (N_17597,N_17494,N_17140);
nand U17598 (N_17598,N_17352,N_17302);
nor U17599 (N_17599,N_16879,N_17310);
and U17600 (N_17600,N_17293,N_17466);
nor U17601 (N_17601,N_17415,N_17292);
and U17602 (N_17602,N_17070,N_17129);
or U17603 (N_17603,N_17014,N_17482);
or U17604 (N_17604,N_16918,N_17010);
and U17605 (N_17605,N_16994,N_17196);
or U17606 (N_17606,N_17142,N_17007);
and U17607 (N_17607,N_16960,N_16991);
nor U17608 (N_17608,N_17253,N_17264);
nor U17609 (N_17609,N_17428,N_16919);
xor U17610 (N_17610,N_17318,N_16956);
nand U17611 (N_17611,N_17179,N_17131);
xnor U17612 (N_17612,N_17213,N_17337);
or U17613 (N_17613,N_17068,N_17066);
or U17614 (N_17614,N_17158,N_17139);
and U17615 (N_17615,N_17365,N_17467);
xnor U17616 (N_17616,N_17232,N_17214);
nand U17617 (N_17617,N_17144,N_17317);
or U17618 (N_17618,N_16973,N_17042);
nand U17619 (N_17619,N_17456,N_17091);
or U17620 (N_17620,N_17105,N_17187);
xnor U17621 (N_17621,N_17098,N_17114);
or U17622 (N_17622,N_17398,N_17245);
nand U17623 (N_17623,N_16971,N_17075);
xor U17624 (N_17624,N_17191,N_17464);
and U17625 (N_17625,N_17150,N_17040);
or U17626 (N_17626,N_17013,N_17335);
and U17627 (N_17627,N_16921,N_17326);
nand U17628 (N_17628,N_17369,N_16985);
nor U17629 (N_17629,N_17207,N_17087);
and U17630 (N_17630,N_17301,N_17490);
nand U17631 (N_17631,N_17004,N_17479);
or U17632 (N_17632,N_17388,N_17353);
nor U17633 (N_17633,N_17107,N_17356);
xnor U17634 (N_17634,N_17359,N_16947);
or U17635 (N_17635,N_16984,N_16963);
nand U17636 (N_17636,N_16910,N_17324);
nand U17637 (N_17637,N_17362,N_17067);
and U17638 (N_17638,N_17003,N_17204);
xor U17639 (N_17639,N_16925,N_16999);
and U17640 (N_17640,N_17472,N_17239);
and U17641 (N_17641,N_16946,N_17108);
xor U17642 (N_17642,N_17019,N_17433);
and U17643 (N_17643,N_17347,N_16987);
nor U17644 (N_17644,N_17005,N_17247);
or U17645 (N_17645,N_17136,N_17412);
or U17646 (N_17646,N_17306,N_17242);
nor U17647 (N_17647,N_17371,N_17476);
xnor U17648 (N_17648,N_17149,N_16988);
xor U17649 (N_17649,N_17200,N_17360);
nand U17650 (N_17650,N_17281,N_17197);
nor U17651 (N_17651,N_16941,N_17000);
and U17652 (N_17652,N_17280,N_17372);
xnor U17653 (N_17653,N_17252,N_17043);
nor U17654 (N_17654,N_17109,N_17319);
and U17655 (N_17655,N_16898,N_17205);
xnor U17656 (N_17656,N_17272,N_17173);
or U17657 (N_17657,N_16891,N_17290);
and U17658 (N_17658,N_17297,N_17099);
and U17659 (N_17659,N_16917,N_17405);
nand U17660 (N_17660,N_17469,N_17277);
or U17661 (N_17661,N_17025,N_17157);
xor U17662 (N_17662,N_17409,N_17315);
and U17663 (N_17663,N_17374,N_17327);
xor U17664 (N_17664,N_17008,N_17097);
xnor U17665 (N_17665,N_17020,N_17168);
and U17666 (N_17666,N_16938,N_17298);
nand U17667 (N_17667,N_17251,N_16889);
nand U17668 (N_17668,N_17026,N_17241);
and U17669 (N_17669,N_17496,N_17121);
and U17670 (N_17670,N_17023,N_17260);
nand U17671 (N_17671,N_16986,N_17051);
and U17672 (N_17672,N_17471,N_16939);
and U17673 (N_17673,N_17155,N_17216);
xnor U17674 (N_17674,N_16937,N_17274);
nand U17675 (N_17675,N_17386,N_17331);
nor U17676 (N_17676,N_17419,N_17395);
nand U17677 (N_17677,N_16912,N_17227);
and U17678 (N_17678,N_17041,N_17255);
xnor U17679 (N_17679,N_17403,N_17275);
or U17680 (N_17680,N_16968,N_17463);
or U17681 (N_17681,N_17343,N_17411);
nand U17682 (N_17682,N_17058,N_17024);
nand U17683 (N_17683,N_17060,N_17250);
and U17684 (N_17684,N_17085,N_17389);
nand U17685 (N_17685,N_16932,N_17309);
nor U17686 (N_17686,N_16894,N_17156);
or U17687 (N_17687,N_17240,N_17407);
and U17688 (N_17688,N_17154,N_17314);
nand U17689 (N_17689,N_17417,N_17233);
or U17690 (N_17690,N_17487,N_17418);
nor U17691 (N_17691,N_17034,N_17248);
xnor U17692 (N_17692,N_17044,N_17027);
and U17693 (N_17693,N_17159,N_17458);
and U17694 (N_17694,N_17050,N_17416);
nand U17695 (N_17695,N_17289,N_17328);
nor U17696 (N_17696,N_17172,N_16951);
or U17697 (N_17697,N_16908,N_17270);
or U17698 (N_17698,N_16903,N_17211);
nor U17699 (N_17699,N_16993,N_17321);
or U17700 (N_17700,N_17332,N_17446);
or U17701 (N_17701,N_17312,N_17377);
nand U17702 (N_17702,N_16875,N_17447);
or U17703 (N_17703,N_17483,N_17284);
nor U17704 (N_17704,N_16928,N_17342);
and U17705 (N_17705,N_17486,N_17257);
nor U17706 (N_17706,N_16893,N_17193);
xor U17707 (N_17707,N_17229,N_17322);
or U17708 (N_17708,N_17018,N_17119);
nor U17709 (N_17709,N_17056,N_16998);
nor U17710 (N_17710,N_17236,N_17052);
and U17711 (N_17711,N_17355,N_17276);
nor U17712 (N_17712,N_17036,N_17423);
and U17713 (N_17713,N_17054,N_17035);
xnor U17714 (N_17714,N_17015,N_16953);
nand U17715 (N_17715,N_17210,N_17083);
xor U17716 (N_17716,N_16934,N_16890);
nor U17717 (N_17717,N_17113,N_17188);
and U17718 (N_17718,N_17246,N_17176);
nor U17719 (N_17719,N_17438,N_16965);
and U17720 (N_17720,N_16916,N_16881);
xnor U17721 (N_17721,N_17189,N_17096);
nor U17722 (N_17722,N_17432,N_16944);
and U17723 (N_17723,N_17118,N_17132);
or U17724 (N_17724,N_17244,N_16882);
and U17725 (N_17725,N_16948,N_17256);
or U17726 (N_17726,N_17146,N_17223);
and U17727 (N_17727,N_16954,N_16883);
xnor U17728 (N_17728,N_17382,N_16877);
nand U17729 (N_17729,N_17169,N_17141);
and U17730 (N_17730,N_17425,N_16978);
nor U17731 (N_17731,N_17031,N_16884);
xnor U17732 (N_17732,N_17406,N_17238);
or U17733 (N_17733,N_17122,N_17126);
or U17734 (N_17734,N_17123,N_17401);
nor U17735 (N_17735,N_17021,N_16900);
and U17736 (N_17736,N_17443,N_17195);
nand U17737 (N_17737,N_17358,N_17088);
nand U17738 (N_17738,N_17167,N_17444);
and U17739 (N_17739,N_17062,N_17424);
nand U17740 (N_17740,N_17381,N_17175);
nand U17741 (N_17741,N_17287,N_17390);
xor U17742 (N_17742,N_17160,N_17380);
xor U17743 (N_17743,N_17300,N_17094);
nor U17744 (N_17744,N_17414,N_17080);
xor U17745 (N_17745,N_17084,N_17303);
nand U17746 (N_17746,N_17151,N_17334);
nand U17747 (N_17747,N_16957,N_16885);
xor U17748 (N_17748,N_17434,N_17498);
and U17749 (N_17749,N_17391,N_16915);
nor U17750 (N_17750,N_17422,N_17038);
nand U17751 (N_17751,N_17402,N_17124);
and U17752 (N_17752,N_17299,N_17459);
or U17753 (N_17753,N_17285,N_17017);
nand U17754 (N_17754,N_17488,N_17453);
nor U17755 (N_17755,N_17037,N_17115);
nand U17756 (N_17756,N_17440,N_17100);
xor U17757 (N_17757,N_17177,N_17243);
or U17758 (N_17758,N_16977,N_17338);
and U17759 (N_17759,N_17296,N_17413);
xnor U17760 (N_17760,N_16943,N_16902);
or U17761 (N_17761,N_17011,N_17092);
nand U17762 (N_17762,N_17408,N_17450);
and U17763 (N_17763,N_17427,N_17028);
xor U17764 (N_17764,N_17354,N_17363);
or U17765 (N_17765,N_16905,N_17039);
nor U17766 (N_17766,N_17384,N_17421);
and U17767 (N_17767,N_17082,N_17001);
nor U17768 (N_17768,N_17128,N_16964);
or U17769 (N_17769,N_17344,N_17073);
nand U17770 (N_17770,N_16976,N_17203);
nand U17771 (N_17771,N_17323,N_17061);
xnor U17772 (N_17772,N_16926,N_17273);
or U17773 (N_17773,N_17258,N_17336);
xor U17774 (N_17774,N_17218,N_17451);
or U17775 (N_17775,N_17436,N_17220);
nor U17776 (N_17776,N_16962,N_16952);
and U17777 (N_17777,N_17212,N_17286);
or U17778 (N_17778,N_17366,N_17333);
or U17779 (N_17779,N_17392,N_17135);
xor U17780 (N_17780,N_17485,N_17090);
nand U17781 (N_17781,N_17138,N_17330);
and U17782 (N_17782,N_17057,N_17431);
nand U17783 (N_17783,N_17404,N_17069);
nand U17784 (N_17784,N_17161,N_16936);
and U17785 (N_17785,N_17076,N_17208);
or U17786 (N_17786,N_17387,N_17454);
nor U17787 (N_17787,N_17198,N_17375);
xor U17788 (N_17788,N_16930,N_17304);
nand U17789 (N_17789,N_17477,N_17379);
or U17790 (N_17790,N_16989,N_17361);
xnor U17791 (N_17791,N_17348,N_17341);
and U17792 (N_17792,N_17267,N_17480);
or U17793 (N_17793,N_17202,N_17145);
xor U17794 (N_17794,N_17370,N_17452);
nand U17795 (N_17795,N_17147,N_16913);
or U17796 (N_17796,N_17133,N_17367);
or U17797 (N_17797,N_17282,N_17445);
xnor U17798 (N_17798,N_17059,N_17215);
nor U17799 (N_17799,N_17206,N_16922);
xnor U17800 (N_17800,N_17268,N_17465);
and U17801 (N_17801,N_16933,N_17226);
nand U17802 (N_17802,N_17185,N_17199);
xor U17803 (N_17803,N_16901,N_16961);
nand U17804 (N_17804,N_17441,N_17170);
nor U17805 (N_17805,N_17209,N_16967);
xor U17806 (N_17806,N_16992,N_17495);
xor U17807 (N_17807,N_17420,N_17426);
nand U17808 (N_17808,N_17111,N_17462);
nor U17809 (N_17809,N_17410,N_17279);
nand U17810 (N_17810,N_16983,N_17357);
and U17811 (N_17811,N_17071,N_17016);
or U17812 (N_17812,N_17376,N_17204);
or U17813 (N_17813,N_17420,N_17332);
or U17814 (N_17814,N_17391,N_17222);
nand U17815 (N_17815,N_16934,N_17391);
xor U17816 (N_17816,N_17231,N_16899);
nor U17817 (N_17817,N_17473,N_17053);
or U17818 (N_17818,N_17321,N_17332);
and U17819 (N_17819,N_16891,N_17409);
nor U17820 (N_17820,N_17405,N_16934);
xor U17821 (N_17821,N_16979,N_17242);
nand U17822 (N_17822,N_17017,N_16891);
nor U17823 (N_17823,N_17336,N_17123);
nand U17824 (N_17824,N_17476,N_17254);
xnor U17825 (N_17825,N_17404,N_17151);
and U17826 (N_17826,N_17336,N_16890);
xor U17827 (N_17827,N_17184,N_16986);
or U17828 (N_17828,N_17168,N_17268);
nor U17829 (N_17829,N_16907,N_16914);
nand U17830 (N_17830,N_16988,N_17376);
nand U17831 (N_17831,N_17343,N_17425);
and U17832 (N_17832,N_17423,N_17273);
nand U17833 (N_17833,N_17274,N_17078);
or U17834 (N_17834,N_17268,N_17124);
and U17835 (N_17835,N_17192,N_16986);
xnor U17836 (N_17836,N_16890,N_17132);
and U17837 (N_17837,N_16912,N_17337);
or U17838 (N_17838,N_17309,N_16991);
xor U17839 (N_17839,N_17243,N_17195);
nand U17840 (N_17840,N_17260,N_17345);
xnor U17841 (N_17841,N_17409,N_17151);
and U17842 (N_17842,N_17226,N_17127);
and U17843 (N_17843,N_17294,N_16901);
nor U17844 (N_17844,N_17338,N_17132);
or U17845 (N_17845,N_17490,N_17397);
xnor U17846 (N_17846,N_17126,N_17478);
nand U17847 (N_17847,N_17153,N_17442);
or U17848 (N_17848,N_17087,N_17164);
and U17849 (N_17849,N_17262,N_16951);
nand U17850 (N_17850,N_17017,N_17442);
xor U17851 (N_17851,N_17211,N_17038);
nand U17852 (N_17852,N_17133,N_17032);
nand U17853 (N_17853,N_17438,N_16962);
and U17854 (N_17854,N_17326,N_17347);
nand U17855 (N_17855,N_16917,N_17484);
nor U17856 (N_17856,N_17359,N_17122);
or U17857 (N_17857,N_17483,N_17296);
and U17858 (N_17858,N_17460,N_17317);
nor U17859 (N_17859,N_17044,N_17119);
or U17860 (N_17860,N_17001,N_17494);
or U17861 (N_17861,N_17247,N_17295);
xnor U17862 (N_17862,N_17445,N_17153);
nor U17863 (N_17863,N_17231,N_16893);
or U17864 (N_17864,N_17166,N_17095);
nand U17865 (N_17865,N_17051,N_16908);
xor U17866 (N_17866,N_17271,N_17275);
nand U17867 (N_17867,N_17359,N_17195);
or U17868 (N_17868,N_17454,N_16964);
nor U17869 (N_17869,N_17139,N_16946);
xnor U17870 (N_17870,N_17475,N_17040);
nor U17871 (N_17871,N_17252,N_16887);
xor U17872 (N_17872,N_16907,N_17463);
and U17873 (N_17873,N_17346,N_17473);
nand U17874 (N_17874,N_17264,N_17154);
xor U17875 (N_17875,N_16966,N_17122);
xor U17876 (N_17876,N_17225,N_16964);
and U17877 (N_17877,N_17429,N_17338);
xnor U17878 (N_17878,N_17223,N_17234);
nand U17879 (N_17879,N_16902,N_17282);
xor U17880 (N_17880,N_17011,N_17289);
nand U17881 (N_17881,N_17231,N_17478);
or U17882 (N_17882,N_16967,N_17308);
nor U17883 (N_17883,N_16884,N_17422);
nor U17884 (N_17884,N_17207,N_17221);
and U17885 (N_17885,N_16945,N_17396);
and U17886 (N_17886,N_17300,N_16972);
nor U17887 (N_17887,N_17478,N_17467);
or U17888 (N_17888,N_17021,N_17003);
nor U17889 (N_17889,N_17351,N_17125);
or U17890 (N_17890,N_17092,N_17165);
and U17891 (N_17891,N_17298,N_17146);
and U17892 (N_17892,N_17309,N_16984);
or U17893 (N_17893,N_17191,N_17487);
or U17894 (N_17894,N_17170,N_17404);
nand U17895 (N_17895,N_17030,N_17138);
or U17896 (N_17896,N_17320,N_17138);
and U17897 (N_17897,N_17261,N_17058);
nor U17898 (N_17898,N_17112,N_17265);
and U17899 (N_17899,N_16973,N_16906);
or U17900 (N_17900,N_17302,N_17306);
or U17901 (N_17901,N_17133,N_17211);
xor U17902 (N_17902,N_17244,N_17125);
xnor U17903 (N_17903,N_17451,N_17021);
and U17904 (N_17904,N_17239,N_16950);
and U17905 (N_17905,N_17212,N_17061);
nor U17906 (N_17906,N_17093,N_16993);
nand U17907 (N_17907,N_17339,N_17343);
and U17908 (N_17908,N_16920,N_17411);
or U17909 (N_17909,N_17495,N_16995);
nand U17910 (N_17910,N_16968,N_17037);
xnor U17911 (N_17911,N_17282,N_17215);
or U17912 (N_17912,N_17353,N_17467);
nor U17913 (N_17913,N_17274,N_17087);
nor U17914 (N_17914,N_17453,N_17058);
nor U17915 (N_17915,N_17362,N_16966);
and U17916 (N_17916,N_17126,N_17247);
nand U17917 (N_17917,N_17172,N_16927);
nand U17918 (N_17918,N_17417,N_17325);
nor U17919 (N_17919,N_17181,N_16940);
and U17920 (N_17920,N_17406,N_17404);
and U17921 (N_17921,N_16927,N_16987);
and U17922 (N_17922,N_17258,N_17338);
and U17923 (N_17923,N_17214,N_16971);
nor U17924 (N_17924,N_17468,N_17059);
xnor U17925 (N_17925,N_17011,N_17433);
xnor U17926 (N_17926,N_16891,N_17284);
nand U17927 (N_17927,N_17078,N_17213);
or U17928 (N_17928,N_17049,N_17363);
nand U17929 (N_17929,N_17427,N_17440);
and U17930 (N_17930,N_16876,N_16880);
or U17931 (N_17931,N_17134,N_17432);
or U17932 (N_17932,N_17072,N_17142);
and U17933 (N_17933,N_17041,N_17206);
or U17934 (N_17934,N_17300,N_16876);
xor U17935 (N_17935,N_16979,N_17043);
and U17936 (N_17936,N_16938,N_17021);
nand U17937 (N_17937,N_16957,N_16996);
or U17938 (N_17938,N_17181,N_16953);
nand U17939 (N_17939,N_17331,N_17039);
xnor U17940 (N_17940,N_17456,N_17000);
and U17941 (N_17941,N_16930,N_17035);
nor U17942 (N_17942,N_17170,N_17444);
nand U17943 (N_17943,N_17213,N_17108);
nor U17944 (N_17944,N_17129,N_17140);
xor U17945 (N_17945,N_17423,N_17271);
nor U17946 (N_17946,N_17337,N_17439);
nor U17947 (N_17947,N_16995,N_17414);
nand U17948 (N_17948,N_17498,N_17229);
or U17949 (N_17949,N_17374,N_17312);
nand U17950 (N_17950,N_17048,N_17252);
or U17951 (N_17951,N_17128,N_17226);
or U17952 (N_17952,N_16944,N_17008);
or U17953 (N_17953,N_16990,N_17037);
xnor U17954 (N_17954,N_17201,N_17238);
nor U17955 (N_17955,N_17265,N_17178);
xnor U17956 (N_17956,N_17166,N_16950);
and U17957 (N_17957,N_16885,N_17145);
and U17958 (N_17958,N_17202,N_17034);
xnor U17959 (N_17959,N_17135,N_17356);
or U17960 (N_17960,N_17264,N_17066);
or U17961 (N_17961,N_17029,N_17361);
nor U17962 (N_17962,N_16970,N_17450);
xnor U17963 (N_17963,N_17049,N_17106);
nor U17964 (N_17964,N_16975,N_16976);
nand U17965 (N_17965,N_17011,N_17194);
nor U17966 (N_17966,N_17370,N_16928);
and U17967 (N_17967,N_17384,N_17287);
nor U17968 (N_17968,N_17199,N_17134);
and U17969 (N_17969,N_17284,N_17336);
nand U17970 (N_17970,N_17015,N_17354);
xor U17971 (N_17971,N_16967,N_17185);
nand U17972 (N_17972,N_17150,N_17397);
or U17973 (N_17973,N_17230,N_17017);
nor U17974 (N_17974,N_17228,N_17106);
or U17975 (N_17975,N_17484,N_17332);
nor U17976 (N_17976,N_17239,N_17129);
or U17977 (N_17977,N_17460,N_17396);
xor U17978 (N_17978,N_17400,N_17451);
nand U17979 (N_17979,N_16993,N_17162);
xnor U17980 (N_17980,N_17266,N_17301);
or U17981 (N_17981,N_17454,N_17134);
xor U17982 (N_17982,N_17239,N_16882);
or U17983 (N_17983,N_16966,N_17001);
or U17984 (N_17984,N_16918,N_17148);
nor U17985 (N_17985,N_16935,N_16984);
xnor U17986 (N_17986,N_16952,N_17412);
nor U17987 (N_17987,N_17311,N_16999);
nor U17988 (N_17988,N_17195,N_17393);
nand U17989 (N_17989,N_17021,N_17226);
nor U17990 (N_17990,N_17210,N_17049);
nand U17991 (N_17991,N_17171,N_17316);
nand U17992 (N_17992,N_17273,N_16954);
nand U17993 (N_17993,N_17307,N_17333);
nor U17994 (N_17994,N_17104,N_17382);
or U17995 (N_17995,N_17032,N_17409);
and U17996 (N_17996,N_16905,N_17402);
and U17997 (N_17997,N_17441,N_17010);
xor U17998 (N_17998,N_17149,N_16887);
xor U17999 (N_17999,N_17185,N_17161);
and U18000 (N_18000,N_16960,N_17145);
or U18001 (N_18001,N_17301,N_17190);
nor U18002 (N_18002,N_17279,N_16975);
xor U18003 (N_18003,N_17338,N_17471);
nor U18004 (N_18004,N_17050,N_17260);
or U18005 (N_18005,N_16991,N_17386);
and U18006 (N_18006,N_17254,N_17459);
nand U18007 (N_18007,N_17093,N_17112);
xnor U18008 (N_18008,N_17162,N_17269);
xnor U18009 (N_18009,N_17321,N_17126);
and U18010 (N_18010,N_17436,N_17219);
xnor U18011 (N_18011,N_17378,N_17399);
and U18012 (N_18012,N_17433,N_17471);
or U18013 (N_18013,N_17226,N_17389);
xnor U18014 (N_18014,N_17483,N_16913);
or U18015 (N_18015,N_17232,N_17361);
and U18016 (N_18016,N_17315,N_16984);
and U18017 (N_18017,N_17492,N_17477);
or U18018 (N_18018,N_17341,N_17034);
nor U18019 (N_18019,N_17361,N_17307);
xor U18020 (N_18020,N_16929,N_16899);
nand U18021 (N_18021,N_17255,N_17131);
nor U18022 (N_18022,N_17313,N_17059);
or U18023 (N_18023,N_17160,N_17350);
and U18024 (N_18024,N_17223,N_17161);
and U18025 (N_18025,N_16932,N_17473);
nor U18026 (N_18026,N_17035,N_17262);
xor U18027 (N_18027,N_17086,N_16892);
and U18028 (N_18028,N_17119,N_17302);
xor U18029 (N_18029,N_17136,N_17012);
nand U18030 (N_18030,N_17391,N_17341);
or U18031 (N_18031,N_17312,N_17135);
nand U18032 (N_18032,N_17390,N_17422);
and U18033 (N_18033,N_17446,N_17192);
nand U18034 (N_18034,N_17103,N_17282);
xor U18035 (N_18035,N_17294,N_17073);
and U18036 (N_18036,N_16954,N_17046);
nand U18037 (N_18037,N_17487,N_17378);
nand U18038 (N_18038,N_16902,N_17074);
xor U18039 (N_18039,N_17294,N_17066);
or U18040 (N_18040,N_17243,N_17098);
nand U18041 (N_18041,N_17209,N_16948);
xnor U18042 (N_18042,N_17220,N_17176);
and U18043 (N_18043,N_17266,N_17128);
nor U18044 (N_18044,N_17492,N_17310);
and U18045 (N_18045,N_16879,N_17264);
nor U18046 (N_18046,N_17185,N_17402);
nor U18047 (N_18047,N_16994,N_17402);
or U18048 (N_18048,N_17051,N_16895);
nor U18049 (N_18049,N_17265,N_16976);
or U18050 (N_18050,N_16946,N_17411);
nand U18051 (N_18051,N_17487,N_17436);
xor U18052 (N_18052,N_17471,N_17105);
nor U18053 (N_18053,N_17159,N_17436);
nor U18054 (N_18054,N_17235,N_16961);
or U18055 (N_18055,N_17180,N_17459);
or U18056 (N_18056,N_17377,N_17319);
or U18057 (N_18057,N_17201,N_16952);
xnor U18058 (N_18058,N_17388,N_17070);
nor U18059 (N_18059,N_17253,N_17098);
nor U18060 (N_18060,N_17406,N_17331);
or U18061 (N_18061,N_17258,N_17402);
nand U18062 (N_18062,N_16993,N_16997);
nand U18063 (N_18063,N_17301,N_17007);
and U18064 (N_18064,N_17380,N_17061);
nor U18065 (N_18065,N_17421,N_17292);
or U18066 (N_18066,N_17380,N_17093);
nor U18067 (N_18067,N_16930,N_16944);
xnor U18068 (N_18068,N_16985,N_17394);
nor U18069 (N_18069,N_17491,N_17010);
and U18070 (N_18070,N_17403,N_17352);
nor U18071 (N_18071,N_17038,N_17349);
xor U18072 (N_18072,N_17034,N_17430);
nand U18073 (N_18073,N_17026,N_17104);
or U18074 (N_18074,N_17201,N_17065);
or U18075 (N_18075,N_17128,N_17136);
or U18076 (N_18076,N_17117,N_16930);
nor U18077 (N_18077,N_16895,N_17196);
xnor U18078 (N_18078,N_17246,N_17097);
nand U18079 (N_18079,N_17280,N_17249);
xor U18080 (N_18080,N_16897,N_16932);
or U18081 (N_18081,N_17344,N_17128);
and U18082 (N_18082,N_16974,N_16945);
nand U18083 (N_18083,N_17471,N_17328);
and U18084 (N_18084,N_17419,N_17207);
and U18085 (N_18085,N_16892,N_17201);
or U18086 (N_18086,N_17112,N_17289);
nor U18087 (N_18087,N_17452,N_17173);
nor U18088 (N_18088,N_17081,N_17244);
xor U18089 (N_18089,N_17418,N_17245);
nor U18090 (N_18090,N_17443,N_17160);
and U18091 (N_18091,N_16977,N_16913);
nor U18092 (N_18092,N_17374,N_17226);
xor U18093 (N_18093,N_17206,N_17434);
and U18094 (N_18094,N_17146,N_17130);
or U18095 (N_18095,N_17135,N_16877);
or U18096 (N_18096,N_17400,N_17163);
xor U18097 (N_18097,N_17205,N_17433);
nand U18098 (N_18098,N_16904,N_16946);
nor U18099 (N_18099,N_17492,N_16918);
nor U18100 (N_18100,N_16982,N_17263);
xnor U18101 (N_18101,N_17337,N_17040);
xor U18102 (N_18102,N_17330,N_17332);
nor U18103 (N_18103,N_17115,N_17444);
and U18104 (N_18104,N_17157,N_17370);
and U18105 (N_18105,N_17402,N_16983);
or U18106 (N_18106,N_17163,N_17440);
or U18107 (N_18107,N_16914,N_17406);
nor U18108 (N_18108,N_16934,N_17388);
and U18109 (N_18109,N_17178,N_17209);
or U18110 (N_18110,N_17248,N_17187);
and U18111 (N_18111,N_17383,N_17327);
nand U18112 (N_18112,N_16991,N_17087);
xnor U18113 (N_18113,N_17461,N_17274);
or U18114 (N_18114,N_17471,N_17499);
and U18115 (N_18115,N_16879,N_17105);
nand U18116 (N_18116,N_17324,N_17430);
or U18117 (N_18117,N_17102,N_17044);
and U18118 (N_18118,N_17014,N_17175);
or U18119 (N_18119,N_17087,N_17069);
nor U18120 (N_18120,N_17016,N_17125);
or U18121 (N_18121,N_16969,N_17420);
nor U18122 (N_18122,N_17040,N_17027);
and U18123 (N_18123,N_17070,N_17203);
nor U18124 (N_18124,N_17350,N_17196);
nand U18125 (N_18125,N_17790,N_17741);
or U18126 (N_18126,N_17869,N_17724);
or U18127 (N_18127,N_17873,N_17917);
xor U18128 (N_18128,N_17574,N_17987);
or U18129 (N_18129,N_17820,N_17984);
nand U18130 (N_18130,N_18061,N_17688);
nand U18131 (N_18131,N_18099,N_18054);
xnor U18132 (N_18132,N_17512,N_17890);
xor U18133 (N_18133,N_17960,N_17847);
nor U18134 (N_18134,N_17630,N_17739);
nand U18135 (N_18135,N_17562,N_17850);
xor U18136 (N_18136,N_18079,N_17657);
or U18137 (N_18137,N_17931,N_17924);
and U18138 (N_18138,N_17798,N_17545);
xor U18139 (N_18139,N_17505,N_17811);
xor U18140 (N_18140,N_17944,N_18119);
xnor U18141 (N_18141,N_17668,N_17882);
xnor U18142 (N_18142,N_17637,N_17620);
or U18143 (N_18143,N_18027,N_17902);
and U18144 (N_18144,N_17569,N_17615);
nor U18145 (N_18145,N_17778,N_18007);
and U18146 (N_18146,N_18009,N_18102);
xor U18147 (N_18147,N_17504,N_17952);
xnor U18148 (N_18148,N_17521,N_17743);
or U18149 (N_18149,N_17605,N_17550);
and U18150 (N_18150,N_17868,N_17571);
nor U18151 (N_18151,N_17855,N_17888);
and U18152 (N_18152,N_18074,N_17883);
nand U18153 (N_18153,N_17655,N_17553);
xnor U18154 (N_18154,N_18075,N_17649);
or U18155 (N_18155,N_17700,N_17996);
nor U18156 (N_18156,N_17968,N_17541);
nor U18157 (N_18157,N_17841,N_17794);
nand U18158 (N_18158,N_17993,N_18066);
xnor U18159 (N_18159,N_17886,N_18076);
nand U18160 (N_18160,N_17681,N_17740);
nand U18161 (N_18161,N_17835,N_17815);
nand U18162 (N_18162,N_17826,N_17747);
nand U18163 (N_18163,N_17540,N_17971);
or U18164 (N_18164,N_17704,N_17723);
xnor U18165 (N_18165,N_17706,N_17654);
or U18166 (N_18166,N_18060,N_17542);
and U18167 (N_18167,N_17889,N_18080);
and U18168 (N_18168,N_17807,N_17581);
nand U18169 (N_18169,N_17726,N_17638);
nand U18170 (N_18170,N_18063,N_17988);
and U18171 (N_18171,N_17619,N_18035);
nand U18172 (N_18172,N_18016,N_17604);
or U18173 (N_18173,N_17840,N_17774);
xnor U18174 (N_18174,N_17560,N_18124);
or U18175 (N_18175,N_17548,N_17782);
nand U18176 (N_18176,N_17733,N_18015);
nand U18177 (N_18177,N_17634,N_17893);
or U18178 (N_18178,N_17641,N_18034);
nor U18179 (N_18179,N_17920,N_17858);
and U18180 (N_18180,N_17628,N_18103);
nor U18181 (N_18181,N_18040,N_17861);
nand U18182 (N_18182,N_18083,N_17537);
or U18183 (N_18183,N_17769,N_17750);
or U18184 (N_18184,N_18020,N_17972);
xnor U18185 (N_18185,N_17701,N_17508);
or U18186 (N_18186,N_17770,N_17953);
nand U18187 (N_18187,N_18085,N_17923);
nand U18188 (N_18188,N_17853,N_17863);
nor U18189 (N_18189,N_17925,N_17880);
and U18190 (N_18190,N_17839,N_17516);
xor U18191 (N_18191,N_17608,N_17500);
or U18192 (N_18192,N_17691,N_17720);
or U18193 (N_18193,N_17866,N_17831);
nor U18194 (N_18194,N_18008,N_18114);
nor U18195 (N_18195,N_17609,N_17989);
xnor U18196 (N_18196,N_17591,N_17843);
xor U18197 (N_18197,N_18037,N_17990);
nand U18198 (N_18198,N_18047,N_17897);
nand U18199 (N_18199,N_18056,N_17502);
and U18200 (N_18200,N_17833,N_17728);
nor U18201 (N_18201,N_18070,N_17819);
xnor U18202 (N_18202,N_18123,N_17799);
nor U18203 (N_18203,N_18052,N_17879);
and U18204 (N_18204,N_17584,N_18071);
and U18205 (N_18205,N_17683,N_17506);
or U18206 (N_18206,N_17690,N_17570);
or U18207 (N_18207,N_18068,N_17806);
nand U18208 (N_18208,N_17875,N_18098);
nand U18209 (N_18209,N_17527,N_17905);
xnor U18210 (N_18210,N_18033,N_17896);
nor U18211 (N_18211,N_17519,N_18097);
xor U18212 (N_18212,N_17695,N_17525);
nand U18213 (N_18213,N_17640,N_17597);
nor U18214 (N_18214,N_17556,N_17746);
xnor U18215 (N_18215,N_17791,N_18118);
xnor U18216 (N_18216,N_18117,N_18105);
xor U18217 (N_18217,N_17535,N_17809);
nor U18218 (N_18218,N_18030,N_17891);
or U18219 (N_18219,N_17689,N_17767);
or U18220 (N_18220,N_17760,N_17511);
or U18221 (N_18221,N_18055,N_17563);
xnor U18222 (N_18222,N_17670,N_17577);
xor U18223 (N_18223,N_17965,N_17981);
and U18224 (N_18224,N_17633,N_17587);
xnor U18225 (N_18225,N_17599,N_17732);
nand U18226 (N_18226,N_17844,N_18110);
nor U18227 (N_18227,N_17694,N_17651);
nand U18228 (N_18228,N_17552,N_17696);
and U18229 (N_18229,N_18023,N_17955);
nor U18230 (N_18230,N_17729,N_17629);
nand U18231 (N_18231,N_17606,N_17699);
nand U18232 (N_18232,N_18108,N_17864);
nor U18233 (N_18233,N_17539,N_17588);
nor U18234 (N_18234,N_18053,N_17718);
nor U18235 (N_18235,N_17503,N_17939);
nand U18236 (N_18236,N_17713,N_18045);
nor U18237 (N_18237,N_17773,N_17959);
nand U18238 (N_18238,N_17942,N_17983);
nand U18239 (N_18239,N_17846,N_17594);
nand U18240 (N_18240,N_17618,N_17738);
nand U18241 (N_18241,N_17632,N_17582);
and U18242 (N_18242,N_17602,N_17522);
and U18243 (N_18243,N_18042,N_17513);
xnor U18244 (N_18244,N_18006,N_17867);
or U18245 (N_18245,N_18028,N_17758);
nand U18246 (N_18246,N_17737,N_17832);
xnor U18247 (N_18247,N_17803,N_17899);
and U18248 (N_18248,N_17631,N_17967);
nor U18249 (N_18249,N_17781,N_18089);
or U18250 (N_18250,N_18014,N_17837);
xor U18251 (N_18251,N_17966,N_17666);
nor U18252 (N_18252,N_17617,N_17580);
nor U18253 (N_18253,N_18101,N_17636);
or U18254 (N_18254,N_17593,N_17936);
nor U18255 (N_18255,N_17823,N_17792);
or U18256 (N_18256,N_17671,N_17995);
nand U18257 (N_18257,N_17528,N_18010);
or U18258 (N_18258,N_17812,N_17674);
nand U18259 (N_18259,N_17547,N_17711);
xor U18260 (N_18260,N_17786,N_17979);
nor U18261 (N_18261,N_18073,N_17946);
or U18262 (N_18262,N_17661,N_17538);
or U18263 (N_18263,N_17603,N_17531);
and U18264 (N_18264,N_17533,N_17518);
nand U18265 (N_18265,N_17607,N_18081);
or U18266 (N_18266,N_17783,N_17887);
xor U18267 (N_18267,N_17561,N_17785);
or U18268 (N_18268,N_17682,N_17777);
xor U18269 (N_18269,N_18093,N_17693);
xor U18270 (N_18270,N_17793,N_17816);
and U18271 (N_18271,N_18090,N_17677);
and U18272 (N_18272,N_17572,N_17749);
nand U18273 (N_18273,N_17878,N_18072);
xor U18274 (N_18274,N_17915,N_18065);
or U18275 (N_18275,N_17529,N_17913);
nand U18276 (N_18276,N_17994,N_17635);
or U18277 (N_18277,N_17517,N_17788);
xnor U18278 (N_18278,N_17731,N_18082);
xnor U18279 (N_18279,N_17849,N_17980);
nor U18280 (N_18280,N_17872,N_18112);
and U18281 (N_18281,N_17940,N_17828);
and U18282 (N_18282,N_17950,N_17565);
or U18283 (N_18283,N_17757,N_17817);
or U18284 (N_18284,N_17575,N_17626);
nor U18285 (N_18285,N_17780,N_17999);
xnor U18286 (N_18286,N_17717,N_17546);
nor U18287 (N_18287,N_17627,N_18029);
nor U18288 (N_18288,N_17851,N_17754);
nand U18289 (N_18289,N_17943,N_17705);
nand U18290 (N_18290,N_17800,N_18012);
and U18291 (N_18291,N_17797,N_18013);
xor U18292 (N_18292,N_17862,N_17702);
or U18293 (N_18293,N_17663,N_17895);
and U18294 (N_18294,N_17600,N_17892);
and U18295 (N_18295,N_17558,N_17721);
xnor U18296 (N_18296,N_17650,N_17673);
or U18297 (N_18297,N_17991,N_17997);
nor U18298 (N_18298,N_17611,N_17568);
xnor U18299 (N_18299,N_17712,N_17669);
and U18300 (N_18300,N_17659,N_17830);
nor U18301 (N_18301,N_17596,N_17910);
nor U18302 (N_18302,N_17762,N_17524);
nor U18303 (N_18303,N_17544,N_17933);
or U18304 (N_18304,N_17859,N_17687);
and U18305 (N_18305,N_18001,N_17860);
xor U18306 (N_18306,N_17822,N_17643);
nand U18307 (N_18307,N_17874,N_17814);
nor U18308 (N_18308,N_17871,N_17672);
xnor U18309 (N_18309,N_17926,N_18057);
and U18310 (N_18310,N_17736,N_18087);
and U18311 (N_18311,N_18019,N_18046);
xnor U18312 (N_18312,N_17573,N_17813);
nand U18313 (N_18313,N_17958,N_17845);
and U18314 (N_18314,N_17795,N_17616);
nor U18315 (N_18315,N_17595,N_17821);
nand U18316 (N_18316,N_17555,N_17507);
nand U18317 (N_18317,N_17623,N_17675);
nor U18318 (N_18318,N_17789,N_17919);
or U18319 (N_18319,N_17656,N_17719);
xnor U18320 (N_18320,N_18018,N_17510);
nor U18321 (N_18321,N_17658,N_17679);
or U18322 (N_18322,N_18064,N_17802);
xnor U18323 (N_18323,N_17804,N_17963);
nor U18324 (N_18324,N_17557,N_17709);
and U18325 (N_18325,N_17536,N_17934);
nand U18326 (N_18326,N_17992,N_17898);
and U18327 (N_18327,N_18111,N_17610);
and U18328 (N_18328,N_17652,N_18106);
nand U18329 (N_18329,N_17856,N_17906);
xor U18330 (N_18330,N_17900,N_17526);
and U18331 (N_18331,N_17928,N_18043);
or U18332 (N_18332,N_17956,N_17775);
nor U18333 (N_18333,N_18025,N_17614);
nand U18334 (N_18334,N_17827,N_17578);
nor U18335 (N_18335,N_17753,N_18088);
or U18336 (N_18336,N_17664,N_17771);
xnor U18337 (N_18337,N_17876,N_17685);
nand U18338 (N_18338,N_18084,N_18078);
xor U18339 (N_18339,N_17662,N_18058);
nand U18340 (N_18340,N_17697,N_17766);
nand U18341 (N_18341,N_17509,N_17865);
xor U18342 (N_18342,N_17918,N_17715);
nand U18343 (N_18343,N_18026,N_17586);
or U18344 (N_18344,N_18095,N_17838);
or U18345 (N_18345,N_18115,N_17549);
or U18346 (N_18346,N_17639,N_17514);
and U18347 (N_18347,N_17707,N_17751);
or U18348 (N_18348,N_17722,N_17911);
xor U18349 (N_18349,N_18094,N_17857);
and U18350 (N_18350,N_18109,N_17885);
and U18351 (N_18351,N_18059,N_17559);
nor U18352 (N_18352,N_17929,N_17554);
nand U18353 (N_18353,N_17759,N_17667);
nand U18354 (N_18354,N_17796,N_17684);
nand U18355 (N_18355,N_17937,N_17824);
and U18356 (N_18356,N_18041,N_18036);
and U18357 (N_18357,N_17982,N_17744);
and U18358 (N_18358,N_17612,N_18122);
xor U18359 (N_18359,N_17613,N_18096);
and U18360 (N_18360,N_17515,N_17938);
nor U18361 (N_18361,N_18086,N_18039);
and U18362 (N_18362,N_17648,N_17752);
or U18363 (N_18363,N_17973,N_17703);
or U18364 (N_18364,N_17948,N_17692);
xnor U18365 (N_18365,N_17742,N_18031);
and U18366 (N_18366,N_17625,N_17801);
and U18367 (N_18367,N_17761,N_17909);
nand U18368 (N_18368,N_17852,N_17589);
nand U18369 (N_18369,N_17622,N_17825);
and U18370 (N_18370,N_17585,N_17908);
and U18371 (N_18371,N_17818,N_17765);
nor U18372 (N_18372,N_18021,N_17921);
xnor U18373 (N_18373,N_17583,N_17564);
xnor U18374 (N_18374,N_17748,N_18104);
nand U18375 (N_18375,N_17930,N_18077);
nor U18376 (N_18376,N_18004,N_17710);
xnor U18377 (N_18377,N_18049,N_17579);
xor U18378 (N_18378,N_17970,N_17543);
xnor U18379 (N_18379,N_17601,N_17949);
and U18380 (N_18380,N_17986,N_17842);
or U18381 (N_18381,N_17954,N_17566);
and U18382 (N_18382,N_18044,N_18032);
nand U18383 (N_18383,N_17784,N_18107);
xnor U18384 (N_18384,N_17964,N_17776);
or U18385 (N_18385,N_17714,N_17922);
and U18386 (N_18386,N_18017,N_18091);
and U18387 (N_18387,N_17534,N_17877);
and U18388 (N_18388,N_17532,N_17810);
and U18389 (N_18389,N_17698,N_18050);
or U18390 (N_18390,N_17894,N_17763);
and U18391 (N_18391,N_17624,N_17947);
and U18392 (N_18392,N_17977,N_18005);
or U18393 (N_18393,N_17551,N_17621);
nand U18394 (N_18394,N_18113,N_17567);
and U18395 (N_18395,N_17756,N_17907);
nand U18396 (N_18396,N_17716,N_17592);
or U18397 (N_18397,N_17975,N_17884);
or U18398 (N_18398,N_17598,N_17881);
and U18399 (N_18399,N_17523,N_17642);
nand U18400 (N_18400,N_17735,N_17725);
nand U18401 (N_18401,N_17914,N_18092);
xor U18402 (N_18402,N_17644,N_18120);
or U18403 (N_18403,N_18011,N_17985);
xnor U18404 (N_18404,N_18116,N_17520);
nand U18405 (N_18405,N_17962,N_17834);
and U18406 (N_18406,N_17647,N_17808);
or U18407 (N_18407,N_17951,N_17957);
nand U18408 (N_18408,N_17927,N_17904);
and U18409 (N_18409,N_17590,N_17708);
nand U18410 (N_18410,N_17755,N_18100);
nor U18411 (N_18411,N_18121,N_17870);
nor U18412 (N_18412,N_17686,N_17680);
nand U18413 (N_18413,N_17501,N_17530);
and U18414 (N_18414,N_17978,N_17660);
nand U18415 (N_18415,N_18002,N_17745);
nor U18416 (N_18416,N_17653,N_18051);
nand U18417 (N_18417,N_17645,N_18024);
or U18418 (N_18418,N_17805,N_17961);
nor U18419 (N_18419,N_17848,N_17976);
xor U18420 (N_18420,N_17916,N_18067);
xor U18421 (N_18421,N_18069,N_17969);
and U18422 (N_18422,N_17676,N_17730);
xnor U18423 (N_18423,N_17901,N_17974);
nor U18424 (N_18424,N_18038,N_17768);
or U18425 (N_18425,N_18022,N_17764);
or U18426 (N_18426,N_18048,N_17935);
or U18427 (N_18427,N_17772,N_17836);
nor U18428 (N_18428,N_17787,N_18000);
nor U18429 (N_18429,N_17665,N_17903);
and U18430 (N_18430,N_17854,N_17678);
nor U18431 (N_18431,N_17727,N_18062);
and U18432 (N_18432,N_17998,N_17912);
or U18433 (N_18433,N_17576,N_17779);
or U18434 (N_18434,N_17941,N_17646);
nor U18435 (N_18435,N_17829,N_17932);
nor U18436 (N_18436,N_17945,N_18003);
nand U18437 (N_18437,N_17734,N_17772);
nor U18438 (N_18438,N_17715,N_17543);
nor U18439 (N_18439,N_17987,N_17646);
and U18440 (N_18440,N_17834,N_17503);
or U18441 (N_18441,N_17777,N_18072);
nor U18442 (N_18442,N_17937,N_17883);
or U18443 (N_18443,N_17912,N_17781);
or U18444 (N_18444,N_17592,N_18093);
nand U18445 (N_18445,N_17932,N_17860);
nor U18446 (N_18446,N_17588,N_17684);
nand U18447 (N_18447,N_17634,N_18001);
or U18448 (N_18448,N_17983,N_18004);
nor U18449 (N_18449,N_17951,N_18020);
nor U18450 (N_18450,N_17841,N_17941);
xnor U18451 (N_18451,N_18072,N_17964);
xnor U18452 (N_18452,N_17688,N_17802);
nor U18453 (N_18453,N_17609,N_17582);
nor U18454 (N_18454,N_18003,N_17644);
nand U18455 (N_18455,N_17718,N_17853);
nor U18456 (N_18456,N_17608,N_17996);
and U18457 (N_18457,N_18053,N_17945);
nand U18458 (N_18458,N_17847,N_17652);
or U18459 (N_18459,N_17693,N_18100);
nor U18460 (N_18460,N_17547,N_17848);
nand U18461 (N_18461,N_17844,N_17674);
nand U18462 (N_18462,N_17977,N_17591);
xor U18463 (N_18463,N_18063,N_18065);
or U18464 (N_18464,N_18043,N_17942);
nand U18465 (N_18465,N_17687,N_18049);
and U18466 (N_18466,N_17902,N_17548);
nand U18467 (N_18467,N_17513,N_17777);
or U18468 (N_18468,N_17504,N_17852);
nor U18469 (N_18469,N_18074,N_18043);
nand U18470 (N_18470,N_18103,N_17809);
and U18471 (N_18471,N_17888,N_17924);
or U18472 (N_18472,N_17874,N_17936);
nand U18473 (N_18473,N_17634,N_18040);
and U18474 (N_18474,N_18033,N_17727);
nand U18475 (N_18475,N_17874,N_18056);
nor U18476 (N_18476,N_17855,N_17984);
and U18477 (N_18477,N_18054,N_17643);
or U18478 (N_18478,N_17543,N_17821);
nand U18479 (N_18479,N_17605,N_17607);
nand U18480 (N_18480,N_17741,N_17523);
xnor U18481 (N_18481,N_18069,N_17568);
and U18482 (N_18482,N_17510,N_18043);
and U18483 (N_18483,N_17961,N_17855);
or U18484 (N_18484,N_17940,N_17568);
xor U18485 (N_18485,N_17506,N_17742);
or U18486 (N_18486,N_17866,N_17964);
xor U18487 (N_18487,N_17726,N_17804);
nand U18488 (N_18488,N_18083,N_18039);
nor U18489 (N_18489,N_17943,N_17561);
nor U18490 (N_18490,N_17693,N_17885);
and U18491 (N_18491,N_17811,N_17778);
xor U18492 (N_18492,N_18116,N_18048);
xnor U18493 (N_18493,N_17868,N_17551);
and U18494 (N_18494,N_17837,N_18075);
nor U18495 (N_18495,N_17985,N_17632);
nor U18496 (N_18496,N_18019,N_18043);
and U18497 (N_18497,N_17775,N_17715);
or U18498 (N_18498,N_17831,N_18096);
and U18499 (N_18499,N_17633,N_18049);
nor U18500 (N_18500,N_17576,N_17855);
and U18501 (N_18501,N_18053,N_17953);
and U18502 (N_18502,N_18124,N_17844);
nand U18503 (N_18503,N_17998,N_17837);
nor U18504 (N_18504,N_17799,N_17642);
nand U18505 (N_18505,N_17740,N_18040);
or U18506 (N_18506,N_18046,N_17758);
nor U18507 (N_18507,N_17977,N_17835);
or U18508 (N_18508,N_18016,N_17566);
nor U18509 (N_18509,N_17687,N_17647);
xnor U18510 (N_18510,N_17782,N_17952);
nor U18511 (N_18511,N_17639,N_17538);
nand U18512 (N_18512,N_17805,N_17503);
or U18513 (N_18513,N_18117,N_17554);
xor U18514 (N_18514,N_18089,N_17780);
nor U18515 (N_18515,N_18021,N_17780);
and U18516 (N_18516,N_17557,N_18065);
nand U18517 (N_18517,N_17631,N_17954);
and U18518 (N_18518,N_17610,N_17895);
xnor U18519 (N_18519,N_17727,N_17742);
nor U18520 (N_18520,N_17855,N_17546);
or U18521 (N_18521,N_17764,N_17771);
nor U18522 (N_18522,N_17781,N_17693);
xor U18523 (N_18523,N_17608,N_17641);
nor U18524 (N_18524,N_17674,N_17842);
and U18525 (N_18525,N_18026,N_18073);
and U18526 (N_18526,N_18073,N_17856);
nand U18527 (N_18527,N_17557,N_17738);
nand U18528 (N_18528,N_17556,N_17581);
or U18529 (N_18529,N_17644,N_18043);
or U18530 (N_18530,N_18006,N_17655);
nor U18531 (N_18531,N_17817,N_17698);
or U18532 (N_18532,N_17803,N_17801);
nor U18533 (N_18533,N_17849,N_18090);
or U18534 (N_18534,N_17756,N_17706);
or U18535 (N_18535,N_17772,N_17777);
and U18536 (N_18536,N_18122,N_17786);
xor U18537 (N_18537,N_18044,N_17613);
xnor U18538 (N_18538,N_17918,N_17512);
nor U18539 (N_18539,N_18053,N_18004);
xnor U18540 (N_18540,N_18049,N_17606);
xnor U18541 (N_18541,N_17646,N_17594);
and U18542 (N_18542,N_17715,N_17757);
nor U18543 (N_18543,N_17916,N_18010);
xor U18544 (N_18544,N_17674,N_18101);
nor U18545 (N_18545,N_18000,N_17562);
nand U18546 (N_18546,N_17785,N_18084);
nand U18547 (N_18547,N_17806,N_17589);
and U18548 (N_18548,N_17710,N_17870);
nor U18549 (N_18549,N_17506,N_18076);
nand U18550 (N_18550,N_18036,N_17899);
nand U18551 (N_18551,N_17880,N_18046);
or U18552 (N_18552,N_17553,N_17594);
nand U18553 (N_18553,N_17629,N_17619);
or U18554 (N_18554,N_17947,N_17657);
and U18555 (N_18555,N_17813,N_18040);
nand U18556 (N_18556,N_17680,N_17582);
xor U18557 (N_18557,N_18007,N_17764);
or U18558 (N_18558,N_17735,N_17835);
or U18559 (N_18559,N_18019,N_17509);
xnor U18560 (N_18560,N_17832,N_17918);
nand U18561 (N_18561,N_17870,N_17647);
nand U18562 (N_18562,N_17677,N_17663);
nand U18563 (N_18563,N_17767,N_17698);
or U18564 (N_18564,N_17549,N_18094);
xor U18565 (N_18565,N_17784,N_18084);
xnor U18566 (N_18566,N_17804,N_17694);
nor U18567 (N_18567,N_17689,N_17500);
xnor U18568 (N_18568,N_17760,N_17609);
xnor U18569 (N_18569,N_18121,N_17535);
nand U18570 (N_18570,N_17773,N_17904);
xnor U18571 (N_18571,N_18006,N_17809);
or U18572 (N_18572,N_17759,N_17732);
nor U18573 (N_18573,N_17973,N_17807);
and U18574 (N_18574,N_17503,N_17913);
and U18575 (N_18575,N_17692,N_18117);
xnor U18576 (N_18576,N_17681,N_17996);
nor U18577 (N_18577,N_17591,N_17913);
nor U18578 (N_18578,N_17869,N_18009);
xor U18579 (N_18579,N_17806,N_17603);
nor U18580 (N_18580,N_17651,N_17718);
nor U18581 (N_18581,N_18107,N_17971);
or U18582 (N_18582,N_17690,N_17842);
and U18583 (N_18583,N_17772,N_17655);
or U18584 (N_18584,N_17613,N_18040);
nor U18585 (N_18585,N_17986,N_17724);
xnor U18586 (N_18586,N_17751,N_17576);
nor U18587 (N_18587,N_17895,N_17750);
nand U18588 (N_18588,N_17884,N_17880);
or U18589 (N_18589,N_17617,N_18026);
or U18590 (N_18590,N_17599,N_17603);
nor U18591 (N_18591,N_17632,N_17659);
xor U18592 (N_18592,N_17512,N_17728);
nand U18593 (N_18593,N_17667,N_17701);
and U18594 (N_18594,N_18123,N_17696);
nor U18595 (N_18595,N_17802,N_17719);
nor U18596 (N_18596,N_17956,N_17760);
and U18597 (N_18597,N_17746,N_17739);
and U18598 (N_18598,N_17502,N_17648);
and U18599 (N_18599,N_17622,N_17737);
nor U18600 (N_18600,N_17744,N_17793);
nand U18601 (N_18601,N_17650,N_18115);
nor U18602 (N_18602,N_18005,N_17695);
or U18603 (N_18603,N_17596,N_17903);
xor U18604 (N_18604,N_17994,N_18066);
nand U18605 (N_18605,N_18079,N_17571);
and U18606 (N_18606,N_17795,N_17931);
nor U18607 (N_18607,N_17807,N_17766);
xor U18608 (N_18608,N_17882,N_17510);
and U18609 (N_18609,N_17555,N_18080);
or U18610 (N_18610,N_17720,N_17623);
xnor U18611 (N_18611,N_17809,N_17510);
or U18612 (N_18612,N_17547,N_17888);
nor U18613 (N_18613,N_18051,N_17543);
or U18614 (N_18614,N_17787,N_17594);
xnor U18615 (N_18615,N_17893,N_17850);
nor U18616 (N_18616,N_18086,N_17638);
and U18617 (N_18617,N_17894,N_18071);
nor U18618 (N_18618,N_17583,N_17946);
nand U18619 (N_18619,N_17652,N_17803);
or U18620 (N_18620,N_17651,N_17537);
or U18621 (N_18621,N_17957,N_17510);
nor U18622 (N_18622,N_17620,N_17833);
and U18623 (N_18623,N_17503,N_17827);
nor U18624 (N_18624,N_17888,N_17751);
nand U18625 (N_18625,N_17816,N_17927);
or U18626 (N_18626,N_17691,N_17673);
nand U18627 (N_18627,N_17701,N_17623);
and U18628 (N_18628,N_18059,N_17874);
nor U18629 (N_18629,N_17950,N_17660);
or U18630 (N_18630,N_17695,N_17969);
nor U18631 (N_18631,N_17846,N_17665);
xnor U18632 (N_18632,N_17573,N_17594);
xnor U18633 (N_18633,N_18056,N_17815);
xnor U18634 (N_18634,N_17907,N_17536);
nor U18635 (N_18635,N_18047,N_17838);
nor U18636 (N_18636,N_17703,N_17897);
nand U18637 (N_18637,N_18038,N_17641);
xnor U18638 (N_18638,N_17546,N_17944);
nor U18639 (N_18639,N_17821,N_17593);
xnor U18640 (N_18640,N_18112,N_17955);
nor U18641 (N_18641,N_17826,N_17644);
xor U18642 (N_18642,N_18005,N_17588);
and U18643 (N_18643,N_17831,N_17667);
or U18644 (N_18644,N_18018,N_17719);
and U18645 (N_18645,N_17708,N_17692);
or U18646 (N_18646,N_17783,N_17836);
nand U18647 (N_18647,N_17995,N_17745);
and U18648 (N_18648,N_17571,N_17926);
xnor U18649 (N_18649,N_17838,N_17689);
nand U18650 (N_18650,N_17927,N_17762);
or U18651 (N_18651,N_17978,N_18078);
nand U18652 (N_18652,N_17953,N_17829);
and U18653 (N_18653,N_17511,N_18032);
and U18654 (N_18654,N_17756,N_17843);
nor U18655 (N_18655,N_17852,N_17793);
nor U18656 (N_18656,N_18104,N_18003);
nand U18657 (N_18657,N_18071,N_17603);
xnor U18658 (N_18658,N_17921,N_17820);
nor U18659 (N_18659,N_17738,N_17703);
nand U18660 (N_18660,N_17869,N_17726);
and U18661 (N_18661,N_18119,N_17778);
xor U18662 (N_18662,N_17591,N_17666);
and U18663 (N_18663,N_17540,N_17764);
nand U18664 (N_18664,N_17757,N_17727);
or U18665 (N_18665,N_18082,N_17857);
and U18666 (N_18666,N_17599,N_17770);
xor U18667 (N_18667,N_17737,N_18083);
nor U18668 (N_18668,N_17512,N_17759);
xor U18669 (N_18669,N_17750,N_17985);
xnor U18670 (N_18670,N_17735,N_17546);
nand U18671 (N_18671,N_17805,N_17922);
nor U18672 (N_18672,N_17500,N_17929);
nor U18673 (N_18673,N_17836,N_18031);
and U18674 (N_18674,N_17677,N_17753);
nor U18675 (N_18675,N_17632,N_17539);
or U18676 (N_18676,N_17612,N_17687);
nand U18677 (N_18677,N_17937,N_17688);
nor U18678 (N_18678,N_17533,N_17847);
xor U18679 (N_18679,N_17547,N_18058);
xnor U18680 (N_18680,N_17721,N_17704);
nor U18681 (N_18681,N_17605,N_17583);
or U18682 (N_18682,N_17920,N_17796);
and U18683 (N_18683,N_17761,N_18106);
or U18684 (N_18684,N_18050,N_17649);
nor U18685 (N_18685,N_17809,N_17500);
nor U18686 (N_18686,N_17657,N_18060);
xnor U18687 (N_18687,N_17669,N_17569);
nand U18688 (N_18688,N_18042,N_17717);
nand U18689 (N_18689,N_17520,N_17516);
and U18690 (N_18690,N_17923,N_17965);
nand U18691 (N_18691,N_17672,N_18017);
nor U18692 (N_18692,N_17621,N_18062);
nor U18693 (N_18693,N_17897,N_17771);
nor U18694 (N_18694,N_17739,N_17905);
xnor U18695 (N_18695,N_18047,N_17854);
or U18696 (N_18696,N_17642,N_17806);
and U18697 (N_18697,N_17653,N_18063);
nor U18698 (N_18698,N_17891,N_17776);
and U18699 (N_18699,N_18048,N_17938);
nand U18700 (N_18700,N_17539,N_17606);
or U18701 (N_18701,N_17952,N_17727);
or U18702 (N_18702,N_17612,N_17651);
nand U18703 (N_18703,N_18066,N_17987);
or U18704 (N_18704,N_17718,N_18122);
and U18705 (N_18705,N_17946,N_18022);
xnor U18706 (N_18706,N_17815,N_17669);
nor U18707 (N_18707,N_17896,N_17550);
nor U18708 (N_18708,N_18009,N_17767);
nand U18709 (N_18709,N_18117,N_17885);
or U18710 (N_18710,N_17782,N_18037);
and U18711 (N_18711,N_17910,N_17574);
and U18712 (N_18712,N_18016,N_17528);
nand U18713 (N_18713,N_17696,N_18071);
nand U18714 (N_18714,N_17832,N_17660);
and U18715 (N_18715,N_17958,N_18067);
or U18716 (N_18716,N_17783,N_17879);
nor U18717 (N_18717,N_17709,N_18014);
xor U18718 (N_18718,N_18052,N_17859);
nor U18719 (N_18719,N_18051,N_18017);
nand U18720 (N_18720,N_17993,N_17705);
nand U18721 (N_18721,N_17923,N_17865);
and U18722 (N_18722,N_17672,N_18057);
and U18723 (N_18723,N_17888,N_17613);
and U18724 (N_18724,N_18081,N_18100);
or U18725 (N_18725,N_17665,N_18049);
nor U18726 (N_18726,N_17630,N_18061);
or U18727 (N_18727,N_18025,N_17860);
xor U18728 (N_18728,N_17890,N_17723);
or U18729 (N_18729,N_18037,N_17515);
or U18730 (N_18730,N_17562,N_17830);
or U18731 (N_18731,N_17613,N_17679);
or U18732 (N_18732,N_18071,N_17977);
or U18733 (N_18733,N_18091,N_18119);
nand U18734 (N_18734,N_17800,N_17621);
nor U18735 (N_18735,N_17507,N_17586);
xor U18736 (N_18736,N_17522,N_17931);
xnor U18737 (N_18737,N_17575,N_17667);
nand U18738 (N_18738,N_17976,N_18039);
xnor U18739 (N_18739,N_17712,N_18048);
xnor U18740 (N_18740,N_17841,N_17510);
or U18741 (N_18741,N_17895,N_18046);
nor U18742 (N_18742,N_17551,N_17668);
and U18743 (N_18743,N_17544,N_17803);
and U18744 (N_18744,N_17624,N_17796);
nand U18745 (N_18745,N_17785,N_17899);
xor U18746 (N_18746,N_17699,N_17955);
nor U18747 (N_18747,N_17871,N_17991);
nor U18748 (N_18748,N_17807,N_17859);
nor U18749 (N_18749,N_17935,N_17624);
xnor U18750 (N_18750,N_18621,N_18262);
or U18751 (N_18751,N_18428,N_18593);
xnor U18752 (N_18752,N_18178,N_18689);
nor U18753 (N_18753,N_18380,N_18278);
nor U18754 (N_18754,N_18470,N_18498);
xnor U18755 (N_18755,N_18196,N_18711);
nor U18756 (N_18756,N_18436,N_18194);
or U18757 (N_18757,N_18740,N_18395);
or U18758 (N_18758,N_18410,N_18149);
and U18759 (N_18759,N_18336,N_18722);
or U18760 (N_18760,N_18360,N_18468);
nand U18761 (N_18761,N_18630,N_18346);
nand U18762 (N_18762,N_18710,N_18610);
nor U18763 (N_18763,N_18382,N_18501);
xor U18764 (N_18764,N_18606,N_18729);
nor U18765 (N_18765,N_18686,N_18153);
xor U18766 (N_18766,N_18645,N_18670);
or U18767 (N_18767,N_18644,N_18411);
xnor U18768 (N_18768,N_18728,N_18313);
nor U18769 (N_18769,N_18130,N_18446);
nor U18770 (N_18770,N_18700,N_18224);
nand U18771 (N_18771,N_18212,N_18595);
and U18772 (N_18772,N_18325,N_18643);
xor U18773 (N_18773,N_18189,N_18459);
xnor U18774 (N_18774,N_18698,N_18443);
or U18775 (N_18775,N_18569,N_18444);
or U18776 (N_18776,N_18682,N_18421);
nor U18777 (N_18777,N_18640,N_18604);
and U18778 (N_18778,N_18423,N_18519);
nor U18779 (N_18779,N_18537,N_18612);
or U18780 (N_18780,N_18478,N_18633);
or U18781 (N_18781,N_18495,N_18575);
and U18782 (N_18782,N_18546,N_18291);
nand U18783 (N_18783,N_18581,N_18496);
nor U18784 (N_18784,N_18182,N_18745);
and U18785 (N_18785,N_18426,N_18329);
xor U18786 (N_18786,N_18678,N_18422);
nand U18787 (N_18787,N_18551,N_18587);
nor U18788 (N_18788,N_18339,N_18237);
xor U18789 (N_18789,N_18260,N_18383);
nor U18790 (N_18790,N_18191,N_18174);
nor U18791 (N_18791,N_18173,N_18417);
nor U18792 (N_18792,N_18431,N_18736);
and U18793 (N_18793,N_18284,N_18205);
nor U18794 (N_18794,N_18139,N_18467);
xor U18795 (N_18795,N_18500,N_18208);
or U18796 (N_18796,N_18374,N_18254);
nand U18797 (N_18797,N_18386,N_18331);
nand U18798 (N_18798,N_18227,N_18337);
nor U18799 (N_18799,N_18508,N_18330);
nor U18800 (N_18800,N_18517,N_18165);
xnor U18801 (N_18801,N_18602,N_18735);
nand U18802 (N_18802,N_18529,N_18287);
nor U18803 (N_18803,N_18715,N_18151);
and U18804 (N_18804,N_18457,N_18163);
nor U18805 (N_18805,N_18349,N_18355);
or U18806 (N_18806,N_18691,N_18415);
or U18807 (N_18807,N_18437,N_18717);
nor U18808 (N_18808,N_18680,N_18694);
nor U18809 (N_18809,N_18352,N_18162);
nor U18810 (N_18810,N_18474,N_18513);
or U18811 (N_18811,N_18128,N_18371);
or U18812 (N_18812,N_18219,N_18539);
and U18813 (N_18813,N_18536,N_18220);
nand U18814 (N_18814,N_18504,N_18193);
and U18815 (N_18815,N_18268,N_18699);
nand U18816 (N_18816,N_18512,N_18659);
nand U18817 (N_18817,N_18358,N_18127);
and U18818 (N_18818,N_18565,N_18541);
nor U18819 (N_18819,N_18323,N_18449);
and U18820 (N_18820,N_18579,N_18140);
nor U18821 (N_18821,N_18239,N_18527);
nor U18822 (N_18822,N_18402,N_18363);
or U18823 (N_18823,N_18530,N_18332);
nor U18824 (N_18824,N_18607,N_18660);
or U18825 (N_18825,N_18738,N_18390);
xnor U18826 (N_18826,N_18248,N_18540);
xnor U18827 (N_18827,N_18142,N_18552);
xnor U18828 (N_18828,N_18672,N_18535);
nand U18829 (N_18829,N_18509,N_18697);
nand U18830 (N_18830,N_18282,N_18350);
xnor U18831 (N_18831,N_18261,N_18186);
nor U18832 (N_18832,N_18458,N_18412);
nor U18833 (N_18833,N_18147,N_18150);
xnor U18834 (N_18834,N_18211,N_18524);
nor U18835 (N_18835,N_18742,N_18472);
xnor U18836 (N_18836,N_18195,N_18401);
and U18837 (N_18837,N_18302,N_18634);
nor U18838 (N_18838,N_18272,N_18746);
nor U18839 (N_18839,N_18393,N_18286);
xor U18840 (N_18840,N_18187,N_18463);
and U18841 (N_18841,N_18560,N_18280);
or U18842 (N_18842,N_18281,N_18143);
nor U18843 (N_18843,N_18623,N_18420);
nand U18844 (N_18844,N_18669,N_18418);
and U18845 (N_18845,N_18319,N_18202);
nor U18846 (N_18846,N_18703,N_18161);
nor U18847 (N_18847,N_18376,N_18741);
nand U18848 (N_18848,N_18279,N_18730);
or U18849 (N_18849,N_18131,N_18615);
or U18850 (N_18850,N_18218,N_18157);
and U18851 (N_18851,N_18304,N_18609);
nor U18852 (N_18852,N_18599,N_18274);
nand U18853 (N_18853,N_18413,N_18583);
and U18854 (N_18854,N_18723,N_18432);
and U18855 (N_18855,N_18335,N_18309);
or U18856 (N_18856,N_18333,N_18226);
or U18857 (N_18857,N_18663,N_18164);
xnor U18858 (N_18858,N_18695,N_18259);
nor U18859 (N_18859,N_18362,N_18392);
or U18860 (N_18860,N_18314,N_18480);
nand U18861 (N_18861,N_18617,N_18430);
nor U18862 (N_18862,N_18559,N_18405);
nand U18863 (N_18863,N_18398,N_18525);
nor U18864 (N_18864,N_18505,N_18315);
and U18865 (N_18865,N_18515,N_18601);
or U18866 (N_18866,N_18377,N_18298);
xnor U18867 (N_18867,N_18733,N_18154);
or U18868 (N_18868,N_18347,N_18448);
xnor U18869 (N_18869,N_18526,N_18646);
nand U18870 (N_18870,N_18485,N_18450);
nor U18871 (N_18871,N_18658,N_18176);
nand U18872 (N_18872,N_18255,N_18198);
or U18873 (N_18873,N_18605,N_18667);
or U18874 (N_18874,N_18693,N_18499);
and U18875 (N_18875,N_18600,N_18132);
nor U18876 (N_18876,N_18493,N_18217);
and U18877 (N_18877,N_18673,N_18241);
nand U18878 (N_18878,N_18522,N_18635);
nor U18879 (N_18879,N_18580,N_18148);
and U18880 (N_18880,N_18242,N_18543);
and U18881 (N_18881,N_18234,N_18531);
nand U18882 (N_18882,N_18396,N_18308);
nand U18883 (N_18883,N_18275,N_18622);
and U18884 (N_18884,N_18385,N_18688);
or U18885 (N_18885,N_18481,N_18231);
nor U18886 (N_18886,N_18483,N_18747);
xor U18887 (N_18887,N_18225,N_18632);
nor U18888 (N_18888,N_18271,N_18320);
nor U18889 (N_18889,N_18144,N_18343);
nor U18890 (N_18890,N_18650,N_18190);
or U18891 (N_18891,N_18582,N_18188);
xnor U18892 (N_18892,N_18408,N_18707);
nor U18893 (N_18893,N_18642,N_18351);
nor U18894 (N_18894,N_18460,N_18136);
nor U18895 (N_18895,N_18183,N_18438);
nor U18896 (N_18896,N_18125,N_18381);
or U18897 (N_18897,N_18613,N_18353);
or U18898 (N_18898,N_18564,N_18326);
xnor U18899 (N_18899,N_18288,N_18263);
and U18900 (N_18900,N_18433,N_18427);
nand U18901 (N_18901,N_18676,N_18591);
nand U18902 (N_18902,N_18236,N_18192);
nor U18903 (N_18903,N_18168,N_18435);
or U18904 (N_18904,N_18283,N_18338);
nor U18905 (N_18905,N_18434,N_18324);
nor U18906 (N_18906,N_18441,N_18316);
or U18907 (N_18907,N_18520,N_18589);
or U18908 (N_18908,N_18618,N_18506);
and U18909 (N_18909,N_18514,N_18230);
xor U18910 (N_18910,N_18684,N_18661);
nor U18911 (N_18911,N_18614,N_18486);
nor U18912 (N_18912,N_18368,N_18456);
nor U18913 (N_18913,N_18429,N_18451);
xor U18914 (N_18914,N_18709,N_18258);
xnor U18915 (N_18915,N_18222,N_18155);
or U18916 (N_18916,N_18584,N_18229);
and U18917 (N_18917,N_18373,N_18243);
or U18918 (N_18918,N_18516,N_18175);
xor U18919 (N_18919,N_18475,N_18488);
or U18920 (N_18920,N_18354,N_18454);
nor U18921 (N_18921,N_18292,N_18538);
and U18922 (N_18922,N_18199,N_18273);
or U18923 (N_18923,N_18487,N_18732);
and U18924 (N_18924,N_18573,N_18716);
nand U18925 (N_18925,N_18249,N_18647);
nand U18926 (N_18926,N_18521,N_18361);
and U18927 (N_18927,N_18177,N_18727);
xnor U18928 (N_18928,N_18636,N_18206);
nor U18929 (N_18929,N_18549,N_18494);
and U18930 (N_18930,N_18654,N_18322);
nand U18931 (N_18931,N_18317,N_18648);
or U18932 (N_18932,N_18370,N_18553);
xor U18933 (N_18933,N_18397,N_18141);
nor U18934 (N_18934,N_18657,N_18510);
and U18935 (N_18935,N_18611,N_18681);
and U18936 (N_18936,N_18653,N_18616);
and U18937 (N_18937,N_18586,N_18312);
xnor U18938 (N_18938,N_18184,N_18562);
and U18939 (N_18939,N_18156,N_18492);
and U18940 (N_18940,N_18384,N_18712);
and U18941 (N_18941,N_18713,N_18718);
xor U18942 (N_18942,N_18447,N_18389);
or U18943 (N_18943,N_18706,N_18200);
xnor U18944 (N_18944,N_18238,N_18185);
xnor U18945 (N_18945,N_18507,N_18749);
nor U18946 (N_18946,N_18692,N_18656);
nand U18947 (N_18947,N_18476,N_18534);
nor U18948 (N_18948,N_18743,N_18369);
or U18949 (N_18949,N_18596,N_18625);
nand U18950 (N_18950,N_18639,N_18251);
and U18951 (N_18951,N_18570,N_18327);
or U18952 (N_18952,N_18482,N_18318);
and U18953 (N_18953,N_18477,N_18419);
xnor U18954 (N_18954,N_18708,N_18590);
xnor U18955 (N_18955,N_18620,N_18266);
and U18956 (N_18956,N_18379,N_18484);
nor U18957 (N_18957,N_18145,N_18264);
nand U18958 (N_18958,N_18558,N_18250);
nand U18959 (N_18959,N_18270,N_18677);
and U18960 (N_18960,N_18424,N_18726);
xnor U18961 (N_18961,N_18294,N_18167);
or U18962 (N_18962,N_18364,N_18702);
or U18963 (N_18963,N_18719,N_18652);
nand U18964 (N_18964,N_18301,N_18341);
xnor U18965 (N_18965,N_18245,N_18440);
nand U18966 (N_18966,N_18567,N_18403);
nand U18967 (N_18967,N_18497,N_18300);
or U18968 (N_18968,N_18137,N_18597);
xor U18969 (N_18969,N_18138,N_18394);
nand U18970 (N_18970,N_18638,N_18399);
or U18971 (N_18971,N_18734,N_18674);
xor U18972 (N_18972,N_18503,N_18626);
and U18973 (N_18973,N_18671,N_18289);
nand U18974 (N_18974,N_18704,N_18223);
or U18975 (N_18975,N_18532,N_18252);
nand U18976 (N_18976,N_18407,N_18391);
and U18977 (N_18977,N_18244,N_18598);
or U18978 (N_18978,N_18213,N_18357);
and U18979 (N_18979,N_18221,N_18629);
nor U18980 (N_18980,N_18180,N_18701);
nand U18981 (N_18981,N_18297,N_18303);
and U18982 (N_18982,N_18561,N_18209);
or U18983 (N_18983,N_18267,N_18572);
nor U18984 (N_18984,N_18511,N_18179);
or U18985 (N_18985,N_18152,N_18170);
nor U18986 (N_18986,N_18556,N_18299);
xnor U18987 (N_18987,N_18310,N_18628);
xnor U18988 (N_18988,N_18345,N_18471);
nor U18989 (N_18989,N_18359,N_18631);
nand U18990 (N_18990,N_18547,N_18690);
and U18991 (N_18991,N_18135,N_18181);
nor U18992 (N_18992,N_18464,N_18683);
xnor U18993 (N_18993,N_18666,N_18554);
and U18994 (N_18994,N_18585,N_18296);
or U18995 (N_18995,N_18207,N_18664);
or U18996 (N_18996,N_18528,N_18406);
and U18997 (N_18997,N_18603,N_18714);
nor U18998 (N_18998,N_18233,N_18473);
xor U18999 (N_18999,N_18276,N_18328);
or U19000 (N_19000,N_18159,N_18721);
and U19001 (N_19001,N_18568,N_18133);
and U19002 (N_19002,N_18518,N_18356);
xnor U19003 (N_19003,N_18348,N_18172);
or U19004 (N_19004,N_18367,N_18344);
or U19005 (N_19005,N_18388,N_18146);
nand U19006 (N_19006,N_18588,N_18204);
and U19007 (N_19007,N_18557,N_18624);
xnor U19008 (N_19008,N_18295,N_18169);
nor U19009 (N_19009,N_18387,N_18240);
or U19010 (N_19010,N_18340,N_18679);
nor U19011 (N_19011,N_18563,N_18416);
and U19012 (N_19012,N_18739,N_18134);
xor U19013 (N_19013,N_18409,N_18725);
nand U19014 (N_19014,N_18290,N_18649);
nor U19015 (N_19015,N_18203,N_18269);
xnor U19016 (N_19016,N_18544,N_18197);
nor U19017 (N_19017,N_18465,N_18453);
nand U19018 (N_19018,N_18491,N_18461);
and U19019 (N_19019,N_18334,N_18414);
xnor U19020 (N_19020,N_18129,N_18574);
or U19021 (N_19021,N_18523,N_18235);
xor U19022 (N_19022,N_18375,N_18651);
nor U19023 (N_19023,N_18228,N_18439);
nor U19024 (N_19024,N_18293,N_18365);
and U19025 (N_19025,N_18533,N_18342);
xnor U19026 (N_19026,N_18724,N_18366);
or U19027 (N_19027,N_18425,N_18201);
xnor U19028 (N_19028,N_18257,N_18305);
nor U19029 (N_19029,N_18247,N_18696);
and U19030 (N_19030,N_18321,N_18214);
and U19031 (N_19031,N_18641,N_18372);
or U19032 (N_19032,N_18489,N_18378);
and U19033 (N_19033,N_18577,N_18479);
xnor U19034 (N_19034,N_18246,N_18166);
nor U19035 (N_19035,N_18490,N_18311);
nor U19036 (N_19036,N_18668,N_18285);
or U19037 (N_19037,N_18215,N_18608);
and U19038 (N_19038,N_18555,N_18256);
nor U19039 (N_19039,N_18744,N_18578);
and U19040 (N_19040,N_18158,N_18592);
nand U19041 (N_19041,N_18216,N_18731);
nand U19042 (N_19042,N_18307,N_18277);
nor U19043 (N_19043,N_18542,N_18637);
xnor U19044 (N_19044,N_18404,N_18502);
or U19045 (N_19045,N_18469,N_18720);
nand U19046 (N_19046,N_18160,N_18455);
nor U19047 (N_19047,N_18619,N_18253);
nand U19048 (N_19048,N_18566,N_18705);
and U19049 (N_19049,N_18462,N_18665);
and U19050 (N_19050,N_18685,N_18400);
xnor U19051 (N_19051,N_18452,N_18576);
xnor U19052 (N_19052,N_18265,N_18655);
nand U19053 (N_19053,N_18210,N_18466);
or U19054 (N_19054,N_18687,N_18548);
xor U19055 (N_19055,N_18126,N_18445);
or U19056 (N_19056,N_18545,N_18675);
nor U19057 (N_19057,N_18737,N_18748);
xnor U19058 (N_19058,N_18550,N_18627);
or U19059 (N_19059,N_18306,N_18571);
nand U19060 (N_19060,N_18662,N_18171);
xor U19061 (N_19061,N_18442,N_18594);
nor U19062 (N_19062,N_18232,N_18341);
xnor U19063 (N_19063,N_18331,N_18436);
or U19064 (N_19064,N_18342,N_18314);
nand U19065 (N_19065,N_18727,N_18198);
and U19066 (N_19066,N_18248,N_18125);
or U19067 (N_19067,N_18410,N_18147);
nand U19068 (N_19068,N_18748,N_18511);
xnor U19069 (N_19069,N_18747,N_18140);
and U19070 (N_19070,N_18495,N_18230);
and U19071 (N_19071,N_18455,N_18310);
nand U19072 (N_19072,N_18457,N_18357);
nor U19073 (N_19073,N_18282,N_18431);
or U19074 (N_19074,N_18540,N_18654);
and U19075 (N_19075,N_18189,N_18279);
xnor U19076 (N_19076,N_18576,N_18262);
xor U19077 (N_19077,N_18652,N_18541);
xnor U19078 (N_19078,N_18728,N_18744);
xnor U19079 (N_19079,N_18701,N_18244);
xor U19080 (N_19080,N_18168,N_18716);
nor U19081 (N_19081,N_18133,N_18208);
or U19082 (N_19082,N_18318,N_18493);
nor U19083 (N_19083,N_18726,N_18223);
xnor U19084 (N_19084,N_18160,N_18641);
xnor U19085 (N_19085,N_18232,N_18632);
xor U19086 (N_19086,N_18312,N_18652);
nand U19087 (N_19087,N_18205,N_18353);
nor U19088 (N_19088,N_18173,N_18291);
nand U19089 (N_19089,N_18268,N_18343);
nand U19090 (N_19090,N_18421,N_18689);
nand U19091 (N_19091,N_18350,N_18684);
and U19092 (N_19092,N_18623,N_18223);
xor U19093 (N_19093,N_18528,N_18493);
and U19094 (N_19094,N_18156,N_18641);
nor U19095 (N_19095,N_18618,N_18393);
xnor U19096 (N_19096,N_18200,N_18290);
nand U19097 (N_19097,N_18536,N_18384);
xor U19098 (N_19098,N_18191,N_18536);
nor U19099 (N_19099,N_18597,N_18237);
nand U19100 (N_19100,N_18235,N_18268);
and U19101 (N_19101,N_18409,N_18237);
or U19102 (N_19102,N_18624,N_18378);
xnor U19103 (N_19103,N_18453,N_18175);
nor U19104 (N_19104,N_18703,N_18417);
nor U19105 (N_19105,N_18594,N_18260);
xor U19106 (N_19106,N_18474,N_18416);
or U19107 (N_19107,N_18461,N_18565);
and U19108 (N_19108,N_18135,N_18577);
nor U19109 (N_19109,N_18362,N_18464);
nand U19110 (N_19110,N_18384,N_18353);
and U19111 (N_19111,N_18584,N_18372);
or U19112 (N_19112,N_18230,N_18159);
xor U19113 (N_19113,N_18630,N_18349);
or U19114 (N_19114,N_18562,N_18271);
and U19115 (N_19115,N_18528,N_18357);
nor U19116 (N_19116,N_18326,N_18186);
nor U19117 (N_19117,N_18227,N_18419);
xor U19118 (N_19118,N_18685,N_18319);
xor U19119 (N_19119,N_18550,N_18581);
xnor U19120 (N_19120,N_18215,N_18499);
or U19121 (N_19121,N_18600,N_18280);
xor U19122 (N_19122,N_18522,N_18668);
nor U19123 (N_19123,N_18388,N_18742);
nor U19124 (N_19124,N_18199,N_18558);
and U19125 (N_19125,N_18196,N_18160);
nand U19126 (N_19126,N_18668,N_18439);
nand U19127 (N_19127,N_18645,N_18744);
nor U19128 (N_19128,N_18604,N_18343);
and U19129 (N_19129,N_18619,N_18417);
or U19130 (N_19130,N_18551,N_18141);
xor U19131 (N_19131,N_18222,N_18466);
nor U19132 (N_19132,N_18736,N_18435);
xor U19133 (N_19133,N_18396,N_18663);
nand U19134 (N_19134,N_18415,N_18304);
nor U19135 (N_19135,N_18183,N_18603);
and U19136 (N_19136,N_18429,N_18515);
nor U19137 (N_19137,N_18371,N_18748);
xor U19138 (N_19138,N_18553,N_18155);
nor U19139 (N_19139,N_18599,N_18442);
or U19140 (N_19140,N_18588,N_18210);
and U19141 (N_19141,N_18406,N_18372);
and U19142 (N_19142,N_18125,N_18620);
nand U19143 (N_19143,N_18511,N_18562);
nor U19144 (N_19144,N_18486,N_18479);
or U19145 (N_19145,N_18580,N_18663);
nor U19146 (N_19146,N_18315,N_18502);
or U19147 (N_19147,N_18430,N_18413);
and U19148 (N_19148,N_18368,N_18455);
xnor U19149 (N_19149,N_18433,N_18274);
and U19150 (N_19150,N_18496,N_18543);
nand U19151 (N_19151,N_18598,N_18399);
and U19152 (N_19152,N_18409,N_18660);
nand U19153 (N_19153,N_18644,N_18491);
nor U19154 (N_19154,N_18697,N_18563);
xnor U19155 (N_19155,N_18357,N_18596);
and U19156 (N_19156,N_18594,N_18600);
or U19157 (N_19157,N_18136,N_18159);
xnor U19158 (N_19158,N_18346,N_18392);
nand U19159 (N_19159,N_18561,N_18312);
nor U19160 (N_19160,N_18716,N_18159);
nor U19161 (N_19161,N_18261,N_18563);
xnor U19162 (N_19162,N_18164,N_18173);
or U19163 (N_19163,N_18569,N_18302);
xor U19164 (N_19164,N_18599,N_18460);
or U19165 (N_19165,N_18552,N_18394);
nor U19166 (N_19166,N_18416,N_18454);
or U19167 (N_19167,N_18741,N_18260);
or U19168 (N_19168,N_18370,N_18242);
nand U19169 (N_19169,N_18126,N_18635);
and U19170 (N_19170,N_18652,N_18448);
xor U19171 (N_19171,N_18215,N_18603);
and U19172 (N_19172,N_18193,N_18129);
and U19173 (N_19173,N_18719,N_18159);
nand U19174 (N_19174,N_18614,N_18152);
or U19175 (N_19175,N_18329,N_18552);
or U19176 (N_19176,N_18691,N_18322);
xor U19177 (N_19177,N_18207,N_18353);
xor U19178 (N_19178,N_18364,N_18663);
nand U19179 (N_19179,N_18184,N_18661);
and U19180 (N_19180,N_18614,N_18375);
or U19181 (N_19181,N_18208,N_18728);
nor U19182 (N_19182,N_18185,N_18271);
and U19183 (N_19183,N_18324,N_18690);
or U19184 (N_19184,N_18748,N_18237);
nand U19185 (N_19185,N_18206,N_18243);
nor U19186 (N_19186,N_18256,N_18315);
nand U19187 (N_19187,N_18162,N_18715);
or U19188 (N_19188,N_18567,N_18473);
or U19189 (N_19189,N_18264,N_18243);
and U19190 (N_19190,N_18393,N_18187);
xor U19191 (N_19191,N_18685,N_18706);
nand U19192 (N_19192,N_18314,N_18584);
and U19193 (N_19193,N_18224,N_18500);
and U19194 (N_19194,N_18237,N_18402);
xnor U19195 (N_19195,N_18146,N_18204);
nor U19196 (N_19196,N_18384,N_18245);
nor U19197 (N_19197,N_18244,N_18737);
xnor U19198 (N_19198,N_18175,N_18334);
and U19199 (N_19199,N_18242,N_18721);
and U19200 (N_19200,N_18194,N_18724);
nand U19201 (N_19201,N_18255,N_18219);
xnor U19202 (N_19202,N_18669,N_18618);
nand U19203 (N_19203,N_18530,N_18141);
or U19204 (N_19204,N_18562,N_18499);
nand U19205 (N_19205,N_18574,N_18348);
and U19206 (N_19206,N_18604,N_18611);
and U19207 (N_19207,N_18467,N_18697);
nand U19208 (N_19208,N_18705,N_18746);
and U19209 (N_19209,N_18695,N_18536);
and U19210 (N_19210,N_18695,N_18452);
nor U19211 (N_19211,N_18497,N_18733);
xor U19212 (N_19212,N_18291,N_18315);
nor U19213 (N_19213,N_18470,N_18282);
nor U19214 (N_19214,N_18237,N_18583);
or U19215 (N_19215,N_18659,N_18423);
and U19216 (N_19216,N_18377,N_18415);
nor U19217 (N_19217,N_18376,N_18195);
or U19218 (N_19218,N_18656,N_18286);
nand U19219 (N_19219,N_18522,N_18727);
nor U19220 (N_19220,N_18595,N_18539);
nor U19221 (N_19221,N_18591,N_18259);
nand U19222 (N_19222,N_18717,N_18656);
xor U19223 (N_19223,N_18238,N_18353);
or U19224 (N_19224,N_18181,N_18518);
nand U19225 (N_19225,N_18723,N_18512);
nor U19226 (N_19226,N_18139,N_18604);
or U19227 (N_19227,N_18588,N_18657);
nand U19228 (N_19228,N_18482,N_18287);
or U19229 (N_19229,N_18328,N_18130);
and U19230 (N_19230,N_18519,N_18320);
nand U19231 (N_19231,N_18134,N_18342);
or U19232 (N_19232,N_18423,N_18430);
or U19233 (N_19233,N_18264,N_18352);
nand U19234 (N_19234,N_18639,N_18676);
xnor U19235 (N_19235,N_18476,N_18278);
or U19236 (N_19236,N_18203,N_18477);
xnor U19237 (N_19237,N_18608,N_18661);
or U19238 (N_19238,N_18727,N_18355);
or U19239 (N_19239,N_18359,N_18538);
xnor U19240 (N_19240,N_18234,N_18164);
nand U19241 (N_19241,N_18452,N_18667);
and U19242 (N_19242,N_18647,N_18729);
xor U19243 (N_19243,N_18155,N_18562);
nor U19244 (N_19244,N_18515,N_18290);
nand U19245 (N_19245,N_18178,N_18583);
or U19246 (N_19246,N_18520,N_18427);
nor U19247 (N_19247,N_18328,N_18335);
and U19248 (N_19248,N_18736,N_18619);
and U19249 (N_19249,N_18283,N_18484);
nand U19250 (N_19250,N_18466,N_18430);
nand U19251 (N_19251,N_18393,N_18676);
nor U19252 (N_19252,N_18369,N_18634);
xor U19253 (N_19253,N_18669,N_18551);
or U19254 (N_19254,N_18576,N_18667);
or U19255 (N_19255,N_18537,N_18198);
nand U19256 (N_19256,N_18558,N_18661);
nand U19257 (N_19257,N_18709,N_18143);
xor U19258 (N_19258,N_18357,N_18666);
nor U19259 (N_19259,N_18545,N_18521);
and U19260 (N_19260,N_18540,N_18324);
or U19261 (N_19261,N_18389,N_18591);
or U19262 (N_19262,N_18578,N_18610);
and U19263 (N_19263,N_18591,N_18549);
nand U19264 (N_19264,N_18290,N_18535);
nand U19265 (N_19265,N_18481,N_18214);
and U19266 (N_19266,N_18144,N_18160);
or U19267 (N_19267,N_18568,N_18149);
nor U19268 (N_19268,N_18628,N_18557);
nand U19269 (N_19269,N_18585,N_18512);
xor U19270 (N_19270,N_18625,N_18659);
nand U19271 (N_19271,N_18598,N_18322);
and U19272 (N_19272,N_18243,N_18226);
xnor U19273 (N_19273,N_18316,N_18684);
nand U19274 (N_19274,N_18675,N_18597);
and U19275 (N_19275,N_18677,N_18642);
nor U19276 (N_19276,N_18559,N_18161);
and U19277 (N_19277,N_18432,N_18580);
nor U19278 (N_19278,N_18696,N_18178);
or U19279 (N_19279,N_18141,N_18242);
xnor U19280 (N_19280,N_18592,N_18629);
or U19281 (N_19281,N_18264,N_18513);
xnor U19282 (N_19282,N_18560,N_18572);
or U19283 (N_19283,N_18674,N_18678);
and U19284 (N_19284,N_18554,N_18548);
or U19285 (N_19285,N_18564,N_18127);
and U19286 (N_19286,N_18312,N_18581);
and U19287 (N_19287,N_18137,N_18606);
nor U19288 (N_19288,N_18498,N_18173);
and U19289 (N_19289,N_18718,N_18704);
or U19290 (N_19290,N_18294,N_18704);
or U19291 (N_19291,N_18312,N_18418);
and U19292 (N_19292,N_18221,N_18205);
nor U19293 (N_19293,N_18512,N_18185);
nand U19294 (N_19294,N_18446,N_18611);
and U19295 (N_19295,N_18444,N_18538);
or U19296 (N_19296,N_18410,N_18603);
or U19297 (N_19297,N_18650,N_18559);
and U19298 (N_19298,N_18664,N_18370);
nor U19299 (N_19299,N_18170,N_18436);
nor U19300 (N_19300,N_18410,N_18570);
and U19301 (N_19301,N_18184,N_18386);
nand U19302 (N_19302,N_18440,N_18297);
or U19303 (N_19303,N_18160,N_18740);
nor U19304 (N_19304,N_18142,N_18201);
and U19305 (N_19305,N_18174,N_18320);
xor U19306 (N_19306,N_18742,N_18412);
nor U19307 (N_19307,N_18306,N_18425);
xnor U19308 (N_19308,N_18410,N_18728);
and U19309 (N_19309,N_18129,N_18678);
or U19310 (N_19310,N_18438,N_18529);
and U19311 (N_19311,N_18653,N_18271);
and U19312 (N_19312,N_18684,N_18747);
nor U19313 (N_19313,N_18500,N_18164);
xnor U19314 (N_19314,N_18358,N_18177);
or U19315 (N_19315,N_18681,N_18283);
nand U19316 (N_19316,N_18747,N_18504);
nand U19317 (N_19317,N_18286,N_18746);
nand U19318 (N_19318,N_18613,N_18634);
or U19319 (N_19319,N_18572,N_18318);
nor U19320 (N_19320,N_18571,N_18661);
and U19321 (N_19321,N_18639,N_18439);
xnor U19322 (N_19322,N_18252,N_18452);
xnor U19323 (N_19323,N_18156,N_18150);
and U19324 (N_19324,N_18182,N_18714);
nand U19325 (N_19325,N_18508,N_18736);
and U19326 (N_19326,N_18624,N_18631);
nor U19327 (N_19327,N_18321,N_18425);
xor U19328 (N_19328,N_18545,N_18498);
xnor U19329 (N_19329,N_18432,N_18468);
and U19330 (N_19330,N_18722,N_18159);
xor U19331 (N_19331,N_18465,N_18497);
xor U19332 (N_19332,N_18533,N_18704);
nor U19333 (N_19333,N_18394,N_18196);
and U19334 (N_19334,N_18746,N_18637);
and U19335 (N_19335,N_18384,N_18210);
nor U19336 (N_19336,N_18525,N_18689);
xnor U19337 (N_19337,N_18483,N_18357);
xor U19338 (N_19338,N_18296,N_18403);
xor U19339 (N_19339,N_18520,N_18529);
and U19340 (N_19340,N_18151,N_18225);
nand U19341 (N_19341,N_18159,N_18205);
xnor U19342 (N_19342,N_18336,N_18334);
nor U19343 (N_19343,N_18310,N_18217);
xnor U19344 (N_19344,N_18399,N_18673);
nand U19345 (N_19345,N_18718,N_18603);
or U19346 (N_19346,N_18226,N_18157);
nand U19347 (N_19347,N_18137,N_18173);
nand U19348 (N_19348,N_18385,N_18239);
xor U19349 (N_19349,N_18525,N_18198);
nor U19350 (N_19350,N_18309,N_18674);
nor U19351 (N_19351,N_18737,N_18308);
and U19352 (N_19352,N_18665,N_18621);
and U19353 (N_19353,N_18682,N_18733);
nand U19354 (N_19354,N_18430,N_18545);
and U19355 (N_19355,N_18168,N_18379);
nor U19356 (N_19356,N_18652,N_18435);
xor U19357 (N_19357,N_18547,N_18515);
and U19358 (N_19358,N_18134,N_18222);
xor U19359 (N_19359,N_18379,N_18656);
nand U19360 (N_19360,N_18687,N_18633);
xor U19361 (N_19361,N_18563,N_18236);
or U19362 (N_19362,N_18564,N_18200);
and U19363 (N_19363,N_18419,N_18323);
xor U19364 (N_19364,N_18576,N_18509);
and U19365 (N_19365,N_18737,N_18624);
or U19366 (N_19366,N_18134,N_18635);
or U19367 (N_19367,N_18213,N_18553);
nor U19368 (N_19368,N_18191,N_18660);
xnor U19369 (N_19369,N_18610,N_18194);
or U19370 (N_19370,N_18133,N_18262);
nor U19371 (N_19371,N_18169,N_18463);
or U19372 (N_19372,N_18552,N_18430);
nand U19373 (N_19373,N_18236,N_18589);
nand U19374 (N_19374,N_18741,N_18444);
or U19375 (N_19375,N_18984,N_19317);
xor U19376 (N_19376,N_19308,N_19216);
nand U19377 (N_19377,N_18883,N_18890);
and U19378 (N_19378,N_19166,N_19069);
or U19379 (N_19379,N_19322,N_19088);
xnor U19380 (N_19380,N_19363,N_19296);
and U19381 (N_19381,N_19018,N_19295);
nor U19382 (N_19382,N_18829,N_18789);
nor U19383 (N_19383,N_19170,N_18995);
nor U19384 (N_19384,N_19168,N_19077);
nand U19385 (N_19385,N_19023,N_18940);
xor U19386 (N_19386,N_18976,N_19146);
or U19387 (N_19387,N_19114,N_19169);
nor U19388 (N_19388,N_18866,N_18760);
nor U19389 (N_19389,N_19218,N_18969);
or U19390 (N_19390,N_18844,N_19070);
nand U19391 (N_19391,N_19139,N_19068);
xor U19392 (N_19392,N_19151,N_19356);
nand U19393 (N_19393,N_19190,N_19150);
nor U19394 (N_19394,N_19210,N_19148);
nand U19395 (N_19395,N_18945,N_19051);
or U19396 (N_19396,N_19319,N_19050);
nor U19397 (N_19397,N_19145,N_18859);
xnor U19398 (N_19398,N_18788,N_18834);
and U19399 (N_19399,N_18861,N_18925);
nand U19400 (N_19400,N_18881,N_18944);
nand U19401 (N_19401,N_18784,N_19043);
xor U19402 (N_19402,N_18865,N_19113);
or U19403 (N_19403,N_19345,N_19231);
and U19404 (N_19404,N_18796,N_19233);
nor U19405 (N_19405,N_19312,N_18801);
or U19406 (N_19406,N_18943,N_19066);
xnor U19407 (N_19407,N_18767,N_19126);
and U19408 (N_19408,N_19336,N_18998);
nand U19409 (N_19409,N_18763,N_19161);
and U19410 (N_19410,N_19270,N_18899);
xnor U19411 (N_19411,N_18840,N_18850);
xor U19412 (N_19412,N_18773,N_18843);
nand U19413 (N_19413,N_18942,N_19264);
nor U19414 (N_19414,N_19232,N_19267);
nor U19415 (N_19415,N_18764,N_19222);
xnor U19416 (N_19416,N_19153,N_18957);
xnor U19417 (N_19417,N_18820,N_19331);
and U19418 (N_19418,N_18846,N_19368);
nor U19419 (N_19419,N_19341,N_19309);
or U19420 (N_19420,N_19040,N_19257);
nand U19421 (N_19421,N_18930,N_19038);
nand U19422 (N_19422,N_18931,N_18948);
xor U19423 (N_19423,N_18884,N_19326);
nand U19424 (N_19424,N_19243,N_19062);
and U19425 (N_19425,N_18937,N_19046);
or U19426 (N_19426,N_19122,N_18900);
and U19427 (N_19427,N_18830,N_19364);
xor U19428 (N_19428,N_19136,N_19199);
or U19429 (N_19429,N_19294,N_18776);
nand U19430 (N_19430,N_18867,N_18838);
nor U19431 (N_19431,N_18982,N_19022);
and U19432 (N_19432,N_19072,N_18818);
or U19433 (N_19433,N_18939,N_18911);
nor U19434 (N_19434,N_18888,N_19196);
xnor U19435 (N_19435,N_19286,N_19029);
and U19436 (N_19436,N_19047,N_19073);
nand U19437 (N_19437,N_18929,N_18825);
and U19438 (N_19438,N_18974,N_18821);
and U19439 (N_19439,N_18781,N_18882);
or U19440 (N_19440,N_19087,N_19223);
or U19441 (N_19441,N_19101,N_19017);
nand U19442 (N_19442,N_19310,N_19283);
xor U19443 (N_19443,N_19352,N_19133);
and U19444 (N_19444,N_19335,N_19256);
xor U19445 (N_19445,N_18753,N_18972);
or U19446 (N_19446,N_19240,N_19276);
xnor U19447 (N_19447,N_19093,N_18992);
nor U19448 (N_19448,N_18953,N_19221);
and U19449 (N_19449,N_18808,N_19273);
nand U19450 (N_19450,N_19001,N_18814);
or U19451 (N_19451,N_18980,N_18924);
and U19452 (N_19452,N_18828,N_18993);
or U19453 (N_19453,N_18868,N_18886);
or U19454 (N_19454,N_18895,N_18827);
or U19455 (N_19455,N_19275,N_18871);
xor U19456 (N_19456,N_19197,N_19289);
nand U19457 (N_19457,N_18935,N_18832);
nand U19458 (N_19458,N_19291,N_18938);
xor U19459 (N_19459,N_19086,N_18914);
nor U19460 (N_19460,N_19365,N_19002);
and U19461 (N_19461,N_19079,N_18877);
and U19462 (N_19462,N_18879,N_19155);
xor U19463 (N_19463,N_19127,N_19293);
or U19464 (N_19464,N_19280,N_18885);
xnor U19465 (N_19465,N_18936,N_19103);
xor U19466 (N_19466,N_18971,N_19315);
nand U19467 (N_19467,N_19193,N_19187);
or U19468 (N_19468,N_19229,N_19098);
or U19469 (N_19469,N_18810,N_18926);
xor U19470 (N_19470,N_19181,N_19048);
nor U19471 (N_19471,N_18787,N_19049);
or U19472 (N_19472,N_18874,N_19344);
or U19473 (N_19473,N_19281,N_18903);
nor U19474 (N_19474,N_18765,N_19074);
nand U19475 (N_19475,N_19194,N_18819);
or U19476 (N_19476,N_19369,N_18812);
and U19477 (N_19477,N_19235,N_18905);
xor U19478 (N_19478,N_19119,N_18824);
xnor U19479 (N_19479,N_19092,N_18927);
and U19480 (N_19480,N_19327,N_18896);
and U19481 (N_19481,N_19214,N_18994);
and U19482 (N_19482,N_18880,N_19238);
nor U19483 (N_19483,N_18949,N_18774);
or U19484 (N_19484,N_19207,N_19247);
nand U19485 (N_19485,N_19245,N_18851);
or U19486 (N_19486,N_18912,N_19096);
xnor U19487 (N_19487,N_18857,N_18910);
nand U19488 (N_19488,N_18970,N_18889);
or U19489 (N_19489,N_19024,N_19180);
nor U19490 (N_19490,N_18915,N_18964);
and U19491 (N_19491,N_19284,N_19012);
nor U19492 (N_19492,N_19129,N_19241);
or U19493 (N_19493,N_18941,N_18958);
xnor U19494 (N_19494,N_19158,N_18946);
nand U19495 (N_19495,N_19000,N_18775);
nor U19496 (N_19496,N_18755,N_19059);
nor U19497 (N_19497,N_18909,N_19274);
and U19498 (N_19498,N_19271,N_19003);
xnor U19499 (N_19499,N_18966,N_19147);
nand U19500 (N_19500,N_19120,N_19045);
nand U19501 (N_19501,N_19172,N_19300);
or U19502 (N_19502,N_19010,N_19228);
or U19503 (N_19503,N_19104,N_19340);
nor U19504 (N_19504,N_19361,N_18869);
nor U19505 (N_19505,N_19025,N_19277);
and U19506 (N_19506,N_19347,N_18963);
nor U19507 (N_19507,N_19099,N_19357);
or U19508 (N_19508,N_19107,N_19348);
or U19509 (N_19509,N_19313,N_19249);
and U19510 (N_19510,N_19329,N_18750);
or U19511 (N_19511,N_18959,N_18908);
nand U19512 (N_19512,N_19225,N_19167);
xnor U19513 (N_19513,N_19255,N_19203);
nor U19514 (N_19514,N_19005,N_19346);
nor U19515 (N_19515,N_19065,N_19115);
or U19516 (N_19516,N_19268,N_19324);
xor U19517 (N_19517,N_19008,N_19039);
and U19518 (N_19518,N_18987,N_18797);
xor U19519 (N_19519,N_19263,N_18862);
nand U19520 (N_19520,N_18907,N_19082);
or U19521 (N_19521,N_18779,N_19085);
nand U19522 (N_19522,N_19083,N_19164);
and U19523 (N_19523,N_18922,N_19041);
nor U19524 (N_19524,N_18758,N_18860);
nand U19525 (N_19525,N_18823,N_19063);
nor U19526 (N_19526,N_19032,N_18920);
or U19527 (N_19527,N_19011,N_19078);
and U19528 (N_19528,N_18836,N_18848);
xnor U19529 (N_19529,N_18921,N_18761);
and U19530 (N_19530,N_18816,N_18997);
nand U19531 (N_19531,N_18878,N_18780);
nand U19532 (N_19532,N_19185,N_18856);
nor U19533 (N_19533,N_19200,N_18973);
nor U19534 (N_19534,N_19044,N_19067);
nor U19535 (N_19535,N_18802,N_18975);
nor U19536 (N_19536,N_19258,N_19131);
nor U19537 (N_19537,N_19367,N_19355);
xnor U19538 (N_19538,N_19287,N_19060);
xnor U19539 (N_19539,N_19248,N_18923);
nand U19540 (N_19540,N_19090,N_18988);
and U19541 (N_19541,N_19349,N_19323);
xor U19542 (N_19542,N_19244,N_19316);
nor U19543 (N_19543,N_19236,N_19250);
xnor U19544 (N_19544,N_19163,N_18906);
nor U19545 (N_19545,N_18813,N_19124);
or U19546 (N_19546,N_18979,N_19261);
nor U19547 (N_19547,N_19128,N_18887);
xnor U19548 (N_19548,N_19290,N_19353);
nand U19549 (N_19549,N_19259,N_18845);
or U19550 (N_19550,N_18904,N_18955);
and U19551 (N_19551,N_19282,N_19108);
xor U19552 (N_19552,N_19125,N_18785);
xor U19553 (N_19553,N_18872,N_19301);
nand U19554 (N_19554,N_18918,N_19334);
or U19555 (N_19555,N_19303,N_18804);
nor U19556 (N_19556,N_19160,N_19373);
xor U19557 (N_19557,N_19095,N_19165);
and U19558 (N_19558,N_19156,N_19304);
and U19559 (N_19559,N_18817,N_19350);
nor U19560 (N_19560,N_19076,N_19297);
nand U19561 (N_19561,N_18919,N_19057);
nand U19562 (N_19562,N_19234,N_19354);
nand U19563 (N_19563,N_19054,N_18951);
xnor U19564 (N_19564,N_18902,N_19251);
xnor U19565 (N_19565,N_18960,N_18978);
nand U19566 (N_19566,N_18854,N_19298);
or U19567 (N_19567,N_18875,N_19112);
nand U19568 (N_19568,N_18913,N_19140);
xnor U19569 (N_19569,N_18800,N_19061);
and U19570 (N_19570,N_18989,N_19135);
xor U19571 (N_19571,N_18783,N_19053);
nor U19572 (N_19572,N_18996,N_19175);
nor U19573 (N_19573,N_19343,N_19342);
nor U19574 (N_19574,N_19253,N_18977);
xor U19575 (N_19575,N_19209,N_19184);
xnor U19576 (N_19576,N_18798,N_19182);
and U19577 (N_19577,N_19116,N_19254);
nand U19578 (N_19578,N_19097,N_19174);
or U19579 (N_19579,N_19089,N_19269);
xor U19580 (N_19580,N_19252,N_19036);
nor U19581 (N_19581,N_19366,N_19118);
or U19582 (N_19582,N_18756,N_18766);
xnor U19583 (N_19583,N_18847,N_18967);
nor U19584 (N_19584,N_19117,N_18901);
xor U19585 (N_19585,N_19035,N_19191);
xnor U19586 (N_19586,N_19004,N_19138);
and U19587 (N_19587,N_18870,N_19212);
nand U19588 (N_19588,N_18876,N_19007);
or U19589 (N_19589,N_19123,N_19102);
nor U19590 (N_19590,N_18757,N_19351);
nand U19591 (N_19591,N_18771,N_18954);
and U19592 (N_19592,N_19328,N_18891);
nor U19593 (N_19593,N_18752,N_19130);
and U19594 (N_19594,N_19056,N_19205);
xor U19595 (N_19595,N_18873,N_19279);
or U19596 (N_19596,N_19037,N_19265);
nand U19597 (N_19597,N_19305,N_18932);
nor U19598 (N_19598,N_19176,N_19262);
xor U19599 (N_19599,N_18839,N_19006);
xor U19600 (N_19600,N_19177,N_18950);
and U19601 (N_19601,N_19311,N_19278);
xnor U19602 (N_19602,N_18772,N_19217);
xnor U19603 (N_19603,N_18842,N_19084);
and U19604 (N_19604,N_19143,N_19110);
xor U19605 (N_19605,N_19159,N_19198);
nand U19606 (N_19606,N_18822,N_18807);
and U19607 (N_19607,N_18990,N_18999);
nor U19608 (N_19608,N_19173,N_19201);
nor U19609 (N_19609,N_19266,N_19224);
nor U19610 (N_19610,N_19299,N_19246);
nor U19611 (N_19611,N_18770,N_19220);
nand U19612 (N_19612,N_18986,N_18809);
and U19613 (N_19613,N_18898,N_19026);
xor U19614 (N_19614,N_19227,N_19171);
and U19615 (N_19615,N_19359,N_18790);
nor U19616 (N_19616,N_19080,N_19213);
and U19617 (N_19617,N_19332,N_18792);
and U19618 (N_19618,N_18852,N_19105);
or U19619 (N_19619,N_19318,N_19337);
and U19620 (N_19620,N_19015,N_18956);
nand U19621 (N_19621,N_19152,N_18928);
nand U19622 (N_19622,N_19307,N_19370);
xor U19623 (N_19623,N_19149,N_19042);
and U19624 (N_19624,N_18985,N_18892);
nor U19625 (N_19625,N_19157,N_18947);
nor U19626 (N_19626,N_18835,N_19142);
or U19627 (N_19627,N_18961,N_19333);
nor U19628 (N_19628,N_19064,N_19091);
or U19629 (N_19629,N_18983,N_19360);
xnor U19630 (N_19630,N_19215,N_18778);
and U19631 (N_19631,N_19206,N_18981);
or U19632 (N_19632,N_18768,N_19321);
or U19633 (N_19633,N_18962,N_19285);
nor U19634 (N_19634,N_18791,N_19211);
nand U19635 (N_19635,N_18786,N_19106);
xor U19636 (N_19636,N_18793,N_19195);
xor U19637 (N_19637,N_19179,N_18897);
nor U19638 (N_19638,N_18864,N_18799);
nor U19639 (N_19639,N_19027,N_19121);
and U19640 (N_19640,N_18769,N_18863);
xor U19641 (N_19641,N_19019,N_19202);
and U19642 (N_19642,N_19111,N_19141);
or U19643 (N_19643,N_18916,N_18853);
xnor U19644 (N_19644,N_19132,N_18805);
xnor U19645 (N_19645,N_18815,N_19100);
or U19646 (N_19646,N_18894,N_18893);
and U19647 (N_19647,N_19016,N_19109);
nand U19648 (N_19648,N_18794,N_19183);
nand U19649 (N_19649,N_18855,N_18841);
and U19650 (N_19650,N_19306,N_19137);
xnor U19651 (N_19651,N_19055,N_19239);
xor U19652 (N_19652,N_19320,N_19204);
and U19653 (N_19653,N_19028,N_18917);
nand U19654 (N_19654,N_18762,N_19081);
nor U19655 (N_19655,N_19020,N_19288);
nand U19656 (N_19656,N_19260,N_19154);
and U19657 (N_19657,N_18837,N_18806);
nand U19658 (N_19658,N_18831,N_19272);
or U19659 (N_19659,N_19330,N_18858);
nand U19660 (N_19660,N_19292,N_19325);
and U19661 (N_19661,N_19188,N_18968);
xor U19662 (N_19662,N_19021,N_19013);
nor U19663 (N_19663,N_19219,N_19237);
xor U19664 (N_19664,N_19362,N_19189);
and U19665 (N_19665,N_19058,N_19186);
and U19666 (N_19666,N_18965,N_19302);
and U19667 (N_19667,N_18991,N_19144);
nor U19668 (N_19668,N_19372,N_19208);
xnor U19669 (N_19669,N_18751,N_19371);
nand U19670 (N_19670,N_18803,N_18759);
nor U19671 (N_19671,N_18952,N_18933);
nand U19672 (N_19672,N_19009,N_19374);
nor U19673 (N_19673,N_18795,N_18782);
nand U19674 (N_19674,N_19242,N_19014);
nand U19675 (N_19675,N_18934,N_19358);
nand U19676 (N_19676,N_19339,N_19031);
xor U19677 (N_19677,N_18849,N_18833);
and U19678 (N_19678,N_19230,N_19134);
and U19679 (N_19679,N_19071,N_19338);
or U19680 (N_19680,N_18826,N_19162);
nand U19681 (N_19681,N_19030,N_19033);
or U19682 (N_19682,N_19178,N_18811);
nor U19683 (N_19683,N_19052,N_18777);
or U19684 (N_19684,N_19094,N_18754);
nor U19685 (N_19685,N_19075,N_19226);
nand U19686 (N_19686,N_19314,N_19192);
and U19687 (N_19687,N_19034,N_18848);
nand U19688 (N_19688,N_19288,N_18947);
xor U19689 (N_19689,N_18846,N_19067);
nor U19690 (N_19690,N_18810,N_18775);
xor U19691 (N_19691,N_19374,N_19027);
nand U19692 (N_19692,N_19050,N_19171);
nor U19693 (N_19693,N_18801,N_19044);
or U19694 (N_19694,N_19051,N_19166);
nor U19695 (N_19695,N_18961,N_19100);
and U19696 (N_19696,N_19151,N_18887);
nor U19697 (N_19697,N_18979,N_19216);
nor U19698 (N_19698,N_19005,N_18967);
or U19699 (N_19699,N_18930,N_19005);
xnor U19700 (N_19700,N_19334,N_19352);
or U19701 (N_19701,N_19183,N_19215);
and U19702 (N_19702,N_19345,N_19288);
and U19703 (N_19703,N_19220,N_19121);
xnor U19704 (N_19704,N_19114,N_19080);
nor U19705 (N_19705,N_19144,N_18877);
nand U19706 (N_19706,N_19107,N_18832);
xor U19707 (N_19707,N_18977,N_18863);
and U19708 (N_19708,N_19272,N_19158);
nand U19709 (N_19709,N_19344,N_18959);
or U19710 (N_19710,N_18955,N_19277);
or U19711 (N_19711,N_19359,N_19049);
nor U19712 (N_19712,N_18920,N_19354);
nand U19713 (N_19713,N_18900,N_19065);
and U19714 (N_19714,N_18909,N_19347);
and U19715 (N_19715,N_19110,N_19101);
nand U19716 (N_19716,N_19095,N_19371);
and U19717 (N_19717,N_19074,N_19283);
xor U19718 (N_19718,N_18750,N_19136);
xor U19719 (N_19719,N_18828,N_18781);
xor U19720 (N_19720,N_18949,N_19168);
xnor U19721 (N_19721,N_19313,N_19345);
nor U19722 (N_19722,N_19228,N_18846);
and U19723 (N_19723,N_19238,N_19122);
xor U19724 (N_19724,N_19197,N_19007);
nand U19725 (N_19725,N_18867,N_19361);
nand U19726 (N_19726,N_19292,N_18838);
or U19727 (N_19727,N_19242,N_19103);
nand U19728 (N_19728,N_19177,N_19220);
xnor U19729 (N_19729,N_18860,N_19032);
xor U19730 (N_19730,N_19283,N_18812);
and U19731 (N_19731,N_18902,N_19249);
xnor U19732 (N_19732,N_18756,N_19049);
xnor U19733 (N_19733,N_18832,N_19188);
or U19734 (N_19734,N_18996,N_19303);
or U19735 (N_19735,N_19299,N_19140);
or U19736 (N_19736,N_19286,N_19069);
or U19737 (N_19737,N_19186,N_19069);
or U19738 (N_19738,N_19270,N_18939);
and U19739 (N_19739,N_18913,N_18835);
or U19740 (N_19740,N_19234,N_19109);
and U19741 (N_19741,N_19156,N_19327);
or U19742 (N_19742,N_19156,N_18983);
xor U19743 (N_19743,N_19246,N_19065);
and U19744 (N_19744,N_18931,N_19118);
nand U19745 (N_19745,N_19108,N_19094);
xor U19746 (N_19746,N_18967,N_19321);
nand U19747 (N_19747,N_18912,N_19327);
xor U19748 (N_19748,N_19283,N_19357);
nand U19749 (N_19749,N_19198,N_18792);
nor U19750 (N_19750,N_19355,N_19066);
nand U19751 (N_19751,N_19272,N_18923);
or U19752 (N_19752,N_19315,N_18808);
nor U19753 (N_19753,N_18976,N_19110);
nor U19754 (N_19754,N_19224,N_19140);
and U19755 (N_19755,N_19153,N_19000);
xor U19756 (N_19756,N_18767,N_19134);
xnor U19757 (N_19757,N_18943,N_19177);
nor U19758 (N_19758,N_18997,N_19260);
xor U19759 (N_19759,N_19065,N_19001);
nand U19760 (N_19760,N_19195,N_19346);
and U19761 (N_19761,N_19356,N_19140);
nand U19762 (N_19762,N_19177,N_18751);
nor U19763 (N_19763,N_18908,N_18845);
and U19764 (N_19764,N_19141,N_18871);
and U19765 (N_19765,N_19013,N_18920);
or U19766 (N_19766,N_18940,N_18825);
or U19767 (N_19767,N_18994,N_18982);
nand U19768 (N_19768,N_19166,N_19221);
xor U19769 (N_19769,N_19001,N_19137);
xnor U19770 (N_19770,N_18994,N_19164);
or U19771 (N_19771,N_19247,N_19216);
and U19772 (N_19772,N_19160,N_18807);
xor U19773 (N_19773,N_19138,N_19356);
and U19774 (N_19774,N_18976,N_19322);
and U19775 (N_19775,N_18998,N_19330);
xor U19776 (N_19776,N_19297,N_19293);
nor U19777 (N_19777,N_19259,N_18943);
nand U19778 (N_19778,N_19047,N_19348);
or U19779 (N_19779,N_18788,N_19016);
nand U19780 (N_19780,N_19349,N_18794);
and U19781 (N_19781,N_19008,N_19064);
nor U19782 (N_19782,N_18881,N_19063);
or U19783 (N_19783,N_18770,N_18916);
and U19784 (N_19784,N_19255,N_19072);
and U19785 (N_19785,N_19003,N_19243);
and U19786 (N_19786,N_18964,N_18999);
and U19787 (N_19787,N_18815,N_19303);
and U19788 (N_19788,N_19012,N_19188);
and U19789 (N_19789,N_18915,N_19081);
nand U19790 (N_19790,N_19018,N_18888);
nor U19791 (N_19791,N_19251,N_18820);
or U19792 (N_19792,N_18802,N_19206);
nor U19793 (N_19793,N_19120,N_19082);
and U19794 (N_19794,N_19277,N_19062);
or U19795 (N_19795,N_19116,N_19042);
nand U19796 (N_19796,N_19162,N_18929);
xnor U19797 (N_19797,N_18987,N_19219);
and U19798 (N_19798,N_19234,N_19283);
and U19799 (N_19799,N_19350,N_18993);
xnor U19800 (N_19800,N_19254,N_19004);
nor U19801 (N_19801,N_19148,N_18887);
xnor U19802 (N_19802,N_18955,N_18818);
or U19803 (N_19803,N_19025,N_18991);
nand U19804 (N_19804,N_19062,N_19082);
and U19805 (N_19805,N_19176,N_18833);
nor U19806 (N_19806,N_18765,N_19179);
or U19807 (N_19807,N_18804,N_19075);
and U19808 (N_19808,N_19133,N_19069);
xnor U19809 (N_19809,N_19258,N_19105);
xor U19810 (N_19810,N_19079,N_19204);
xor U19811 (N_19811,N_19258,N_18841);
or U19812 (N_19812,N_18982,N_18873);
or U19813 (N_19813,N_18826,N_19372);
nor U19814 (N_19814,N_18885,N_19054);
nor U19815 (N_19815,N_18998,N_19143);
and U19816 (N_19816,N_19158,N_19089);
or U19817 (N_19817,N_19045,N_19131);
nor U19818 (N_19818,N_18826,N_18971);
xor U19819 (N_19819,N_18916,N_19166);
nand U19820 (N_19820,N_18996,N_19316);
nand U19821 (N_19821,N_19265,N_19014);
nand U19822 (N_19822,N_18817,N_19365);
xnor U19823 (N_19823,N_18970,N_18845);
nand U19824 (N_19824,N_19275,N_18977);
or U19825 (N_19825,N_18951,N_19276);
xor U19826 (N_19826,N_18948,N_18806);
nand U19827 (N_19827,N_18817,N_19221);
or U19828 (N_19828,N_18844,N_18788);
nand U19829 (N_19829,N_19199,N_19241);
nor U19830 (N_19830,N_18984,N_18845);
nor U19831 (N_19831,N_19145,N_19072);
nor U19832 (N_19832,N_18934,N_19331);
nor U19833 (N_19833,N_18917,N_19296);
and U19834 (N_19834,N_18843,N_19109);
nand U19835 (N_19835,N_19146,N_19124);
and U19836 (N_19836,N_18987,N_19347);
and U19837 (N_19837,N_18977,N_19266);
nand U19838 (N_19838,N_19371,N_18908);
and U19839 (N_19839,N_19118,N_18850);
or U19840 (N_19840,N_18982,N_19335);
or U19841 (N_19841,N_18838,N_18841);
and U19842 (N_19842,N_18820,N_19212);
and U19843 (N_19843,N_18757,N_18813);
xnor U19844 (N_19844,N_19191,N_19004);
or U19845 (N_19845,N_19313,N_19354);
xnor U19846 (N_19846,N_19236,N_18977);
and U19847 (N_19847,N_19123,N_18803);
nand U19848 (N_19848,N_18944,N_19057);
or U19849 (N_19849,N_18807,N_19247);
or U19850 (N_19850,N_18806,N_18899);
xnor U19851 (N_19851,N_18896,N_18814);
and U19852 (N_19852,N_19341,N_19314);
and U19853 (N_19853,N_18814,N_18772);
xor U19854 (N_19854,N_19032,N_19053);
nand U19855 (N_19855,N_19007,N_18933);
and U19856 (N_19856,N_19010,N_18756);
or U19857 (N_19857,N_18761,N_19264);
xor U19858 (N_19858,N_18883,N_19086);
nand U19859 (N_19859,N_19025,N_18822);
nand U19860 (N_19860,N_19347,N_18993);
and U19861 (N_19861,N_18864,N_18857);
or U19862 (N_19862,N_18958,N_19149);
xor U19863 (N_19863,N_18873,N_19363);
xnor U19864 (N_19864,N_19353,N_19356);
or U19865 (N_19865,N_19071,N_19348);
or U19866 (N_19866,N_18961,N_18807);
nand U19867 (N_19867,N_19072,N_18905);
nand U19868 (N_19868,N_18942,N_19211);
or U19869 (N_19869,N_18870,N_19218);
or U19870 (N_19870,N_19113,N_18879);
nor U19871 (N_19871,N_18931,N_19089);
xnor U19872 (N_19872,N_18889,N_19194);
nand U19873 (N_19873,N_19170,N_18863);
or U19874 (N_19874,N_19085,N_18951);
nand U19875 (N_19875,N_19344,N_19304);
or U19876 (N_19876,N_18869,N_19324);
or U19877 (N_19877,N_18831,N_18973);
or U19878 (N_19878,N_18954,N_19362);
nand U19879 (N_19879,N_19289,N_19057);
nand U19880 (N_19880,N_19019,N_18996);
nor U19881 (N_19881,N_19259,N_18803);
and U19882 (N_19882,N_18983,N_18786);
nor U19883 (N_19883,N_19141,N_18770);
nor U19884 (N_19884,N_18791,N_19319);
nand U19885 (N_19885,N_18957,N_19298);
and U19886 (N_19886,N_19033,N_18766);
nand U19887 (N_19887,N_19236,N_18875);
nand U19888 (N_19888,N_18750,N_18812);
nor U19889 (N_19889,N_19339,N_19071);
nand U19890 (N_19890,N_18850,N_19129);
nand U19891 (N_19891,N_18965,N_19020);
nor U19892 (N_19892,N_19145,N_18910);
nand U19893 (N_19893,N_19361,N_19329);
nor U19894 (N_19894,N_19276,N_18826);
nor U19895 (N_19895,N_19171,N_19239);
nand U19896 (N_19896,N_18783,N_18987);
nand U19897 (N_19897,N_19222,N_19162);
xor U19898 (N_19898,N_18898,N_19333);
or U19899 (N_19899,N_18998,N_19057);
and U19900 (N_19900,N_19134,N_19304);
and U19901 (N_19901,N_19019,N_19201);
xnor U19902 (N_19902,N_19230,N_18989);
and U19903 (N_19903,N_19109,N_18899);
and U19904 (N_19904,N_19073,N_19358);
or U19905 (N_19905,N_18913,N_19169);
and U19906 (N_19906,N_18984,N_18826);
nand U19907 (N_19907,N_19192,N_19364);
or U19908 (N_19908,N_19198,N_18932);
nand U19909 (N_19909,N_19231,N_18876);
or U19910 (N_19910,N_19100,N_18899);
and U19911 (N_19911,N_19054,N_19067);
nor U19912 (N_19912,N_18793,N_18804);
nor U19913 (N_19913,N_18938,N_19098);
nor U19914 (N_19914,N_19365,N_19162);
xnor U19915 (N_19915,N_19216,N_19081);
xnor U19916 (N_19916,N_18773,N_19116);
or U19917 (N_19917,N_19276,N_19175);
nor U19918 (N_19918,N_19312,N_19221);
nand U19919 (N_19919,N_19149,N_18948);
nor U19920 (N_19920,N_18912,N_18826);
xnor U19921 (N_19921,N_19228,N_18774);
xnor U19922 (N_19922,N_18971,N_19180);
and U19923 (N_19923,N_18890,N_19103);
nand U19924 (N_19924,N_19334,N_19002);
nor U19925 (N_19925,N_19308,N_18998);
nor U19926 (N_19926,N_18929,N_19355);
and U19927 (N_19927,N_18941,N_19284);
xnor U19928 (N_19928,N_18761,N_19291);
nand U19929 (N_19929,N_19347,N_18975);
nor U19930 (N_19930,N_18804,N_18971);
nand U19931 (N_19931,N_19127,N_19259);
nand U19932 (N_19932,N_19021,N_19357);
nand U19933 (N_19933,N_19263,N_19177);
or U19934 (N_19934,N_19104,N_19202);
and U19935 (N_19935,N_18936,N_19259);
and U19936 (N_19936,N_19081,N_19145);
xor U19937 (N_19937,N_19175,N_18906);
and U19938 (N_19938,N_19196,N_18852);
nand U19939 (N_19939,N_19078,N_18845);
and U19940 (N_19940,N_18862,N_19041);
nand U19941 (N_19941,N_18794,N_18782);
xor U19942 (N_19942,N_18851,N_19108);
nor U19943 (N_19943,N_18813,N_19103);
and U19944 (N_19944,N_19334,N_19133);
xor U19945 (N_19945,N_18763,N_19267);
nor U19946 (N_19946,N_19308,N_19179);
xor U19947 (N_19947,N_19214,N_18769);
and U19948 (N_19948,N_18832,N_19118);
xor U19949 (N_19949,N_18816,N_18956);
nand U19950 (N_19950,N_18841,N_19190);
nand U19951 (N_19951,N_18955,N_19176);
or U19952 (N_19952,N_19203,N_18807);
xor U19953 (N_19953,N_19169,N_18754);
nor U19954 (N_19954,N_18793,N_19068);
xor U19955 (N_19955,N_18931,N_19189);
or U19956 (N_19956,N_18959,N_19214);
or U19957 (N_19957,N_19063,N_18826);
or U19958 (N_19958,N_19013,N_18944);
nand U19959 (N_19959,N_19122,N_19131);
xor U19960 (N_19960,N_19133,N_19055);
and U19961 (N_19961,N_18912,N_19082);
nand U19962 (N_19962,N_18956,N_18838);
nor U19963 (N_19963,N_18930,N_18785);
nor U19964 (N_19964,N_18923,N_18934);
xor U19965 (N_19965,N_19372,N_18804);
and U19966 (N_19966,N_19219,N_19342);
nand U19967 (N_19967,N_18760,N_19167);
xnor U19968 (N_19968,N_18952,N_19200);
and U19969 (N_19969,N_18925,N_19103);
nor U19970 (N_19970,N_19048,N_19001);
nor U19971 (N_19971,N_18875,N_18971);
xnor U19972 (N_19972,N_19310,N_18783);
xnor U19973 (N_19973,N_19113,N_19263);
or U19974 (N_19974,N_18825,N_19104);
or U19975 (N_19975,N_19323,N_19135);
xnor U19976 (N_19976,N_19153,N_18886);
or U19977 (N_19977,N_19018,N_18763);
xnor U19978 (N_19978,N_18781,N_19126);
nand U19979 (N_19979,N_19316,N_19314);
or U19980 (N_19980,N_19350,N_19295);
or U19981 (N_19981,N_19044,N_18944);
or U19982 (N_19982,N_19263,N_19020);
xor U19983 (N_19983,N_19231,N_19173);
or U19984 (N_19984,N_18935,N_19200);
nand U19985 (N_19985,N_18757,N_18850);
and U19986 (N_19986,N_18977,N_19317);
and U19987 (N_19987,N_19167,N_18962);
or U19988 (N_19988,N_19070,N_18922);
or U19989 (N_19989,N_18962,N_19025);
or U19990 (N_19990,N_19324,N_19259);
nor U19991 (N_19991,N_19094,N_18993);
nor U19992 (N_19992,N_19007,N_18912);
or U19993 (N_19993,N_18958,N_19318);
nor U19994 (N_19994,N_19252,N_19128);
or U19995 (N_19995,N_19311,N_19226);
or U19996 (N_19996,N_19086,N_18829);
xnor U19997 (N_19997,N_18834,N_18796);
and U19998 (N_19998,N_19153,N_19048);
xnor U19999 (N_19999,N_19022,N_18797);
or U20000 (N_20000,N_19865,N_19923);
nor U20001 (N_20001,N_19728,N_19487);
or U20002 (N_20002,N_19604,N_19881);
nor U20003 (N_20003,N_19571,N_19933);
xor U20004 (N_20004,N_19917,N_19740);
nand U20005 (N_20005,N_19450,N_19593);
or U20006 (N_20006,N_19530,N_19555);
and U20007 (N_20007,N_19532,N_19935);
nand U20008 (N_20008,N_19391,N_19770);
nand U20009 (N_20009,N_19922,N_19485);
nor U20010 (N_20010,N_19803,N_19989);
xor U20011 (N_20011,N_19823,N_19381);
nor U20012 (N_20012,N_19410,N_19779);
nor U20013 (N_20013,N_19725,N_19375);
or U20014 (N_20014,N_19460,N_19417);
or U20015 (N_20015,N_19415,N_19925);
nor U20016 (N_20016,N_19936,N_19574);
nand U20017 (N_20017,N_19901,N_19378);
or U20018 (N_20018,N_19743,N_19746);
or U20019 (N_20019,N_19861,N_19760);
nand U20020 (N_20020,N_19491,N_19641);
nor U20021 (N_20021,N_19840,N_19634);
nor U20022 (N_20022,N_19851,N_19897);
nand U20023 (N_20023,N_19900,N_19787);
nand U20024 (N_20024,N_19958,N_19835);
xor U20025 (N_20025,N_19678,N_19553);
nor U20026 (N_20026,N_19658,N_19916);
nor U20027 (N_20027,N_19704,N_19686);
nor U20028 (N_20028,N_19612,N_19763);
xnor U20029 (N_20029,N_19581,N_19439);
and U20030 (N_20030,N_19878,N_19483);
or U20031 (N_20031,N_19996,N_19843);
nand U20032 (N_20032,N_19799,N_19719);
and U20033 (N_20033,N_19540,N_19440);
nand U20034 (N_20034,N_19846,N_19506);
nand U20035 (N_20035,N_19393,N_19499);
nor U20036 (N_20036,N_19937,N_19551);
xnor U20037 (N_20037,N_19462,N_19741);
and U20038 (N_20038,N_19665,N_19709);
nand U20039 (N_20039,N_19691,N_19722);
nand U20040 (N_20040,N_19498,N_19692);
nand U20041 (N_20041,N_19408,N_19489);
or U20042 (N_20042,N_19533,N_19784);
nand U20043 (N_20043,N_19972,N_19463);
xor U20044 (N_20044,N_19957,N_19667);
nand U20045 (N_20045,N_19880,N_19697);
xnor U20046 (N_20046,N_19405,N_19931);
or U20047 (N_20047,N_19761,N_19831);
xnor U20048 (N_20048,N_19479,N_19602);
xnor U20049 (N_20049,N_19973,N_19425);
nor U20050 (N_20050,N_19568,N_19449);
nor U20051 (N_20051,N_19857,N_19626);
nor U20052 (N_20052,N_19514,N_19982);
or U20053 (N_20053,N_19681,N_19815);
and U20054 (N_20054,N_19749,N_19587);
xor U20055 (N_20055,N_19909,N_19411);
nor U20056 (N_20056,N_19492,N_19519);
or U20057 (N_20057,N_19976,N_19652);
or U20058 (N_20058,N_19625,N_19580);
xor U20059 (N_20059,N_19536,N_19527);
and U20060 (N_20060,N_19594,N_19905);
or U20061 (N_20061,N_19511,N_19806);
nor U20062 (N_20062,N_19855,N_19507);
or U20063 (N_20063,N_19930,N_19643);
xor U20064 (N_20064,N_19856,N_19689);
or U20065 (N_20065,N_19377,N_19785);
xnor U20066 (N_20066,N_19836,N_19791);
xnor U20067 (N_20067,N_19899,N_19380);
nand U20068 (N_20068,N_19828,N_19622);
nand U20069 (N_20069,N_19804,N_19910);
or U20070 (N_20070,N_19517,N_19600);
nand U20071 (N_20071,N_19503,N_19703);
xnor U20072 (N_20072,N_19759,N_19550);
and U20073 (N_20073,N_19613,N_19558);
nor U20074 (N_20074,N_19453,N_19902);
and U20075 (N_20075,N_19452,N_19797);
and U20076 (N_20076,N_19591,N_19610);
nor U20077 (N_20077,N_19954,N_19750);
or U20078 (N_20078,N_19694,N_19446);
or U20079 (N_20079,N_19628,N_19995);
xor U20080 (N_20080,N_19466,N_19870);
xnor U20081 (N_20081,N_19685,N_19726);
nand U20082 (N_20082,N_19817,N_19968);
nand U20083 (N_20083,N_19911,N_19423);
nand U20084 (N_20084,N_19786,N_19397);
nand U20085 (N_20085,N_19898,N_19951);
xnor U20086 (N_20086,N_19734,N_19546);
or U20087 (N_20087,N_19673,N_19820);
nand U20088 (N_20088,N_19599,N_19642);
or U20089 (N_20089,N_19394,N_19971);
nand U20090 (N_20090,N_19758,N_19644);
or U20091 (N_20091,N_19890,N_19822);
xnor U20092 (N_20092,N_19829,N_19413);
xor U20093 (N_20093,N_19860,N_19541);
xor U20094 (N_20094,N_19648,N_19889);
nand U20095 (N_20095,N_19913,N_19619);
nand U20096 (N_20096,N_19987,N_19895);
or U20097 (N_20097,N_19941,N_19508);
and U20098 (N_20098,N_19493,N_19674);
nand U20099 (N_20099,N_19896,N_19950);
or U20100 (N_20100,N_19979,N_19780);
or U20101 (N_20101,N_19382,N_19608);
nor U20102 (N_20102,N_19929,N_19448);
xor U20103 (N_20103,N_19547,N_19427);
xor U20104 (N_20104,N_19486,N_19821);
and U20105 (N_20105,N_19653,N_19712);
and U20106 (N_20106,N_19967,N_19947);
or U20107 (N_20107,N_19502,N_19762);
xnor U20108 (N_20108,N_19592,N_19827);
and U20109 (N_20109,N_19755,N_19469);
and U20110 (N_20110,N_19969,N_19738);
nor U20111 (N_20111,N_19699,N_19818);
or U20112 (N_20112,N_19518,N_19504);
and U20113 (N_20113,N_19538,N_19980);
nand U20114 (N_20114,N_19419,N_19934);
nand U20115 (N_20115,N_19789,N_19396);
or U20116 (N_20116,N_19528,N_19904);
xor U20117 (N_20117,N_19430,N_19988);
nor U20118 (N_20118,N_19471,N_19490);
nand U20119 (N_20119,N_19675,N_19735);
or U20120 (N_20120,N_19757,N_19633);
or U20121 (N_20121,N_19565,N_19707);
nor U20122 (N_20122,N_19983,N_19556);
or U20123 (N_20123,N_19570,N_19970);
nor U20124 (N_20124,N_19867,N_19744);
nor U20125 (N_20125,N_19645,N_19801);
nor U20126 (N_20126,N_19386,N_19832);
nand U20127 (N_20127,N_19383,N_19621);
or U20128 (N_20128,N_19554,N_19876);
nor U20129 (N_20129,N_19721,N_19636);
nor U20130 (N_20130,N_19474,N_19447);
xnor U20131 (N_20131,N_19647,N_19847);
xor U20132 (N_20132,N_19616,N_19676);
nand U20133 (N_20133,N_19557,N_19908);
nand U20134 (N_20134,N_19809,N_19775);
or U20135 (N_20135,N_19814,N_19918);
nor U20136 (N_20136,N_19389,N_19960);
nand U20137 (N_20137,N_19919,N_19457);
xor U20138 (N_20138,N_19624,N_19404);
nor U20139 (N_20139,N_19614,N_19526);
xor U20140 (N_20140,N_19522,N_19588);
nor U20141 (N_20141,N_19742,N_19584);
or U20142 (N_20142,N_19903,N_19655);
and U20143 (N_20143,N_19595,N_19564);
nand U20144 (N_20144,N_19458,N_19777);
nor U20145 (N_20145,N_19577,N_19400);
nor U20146 (N_20146,N_19912,N_19959);
and U20147 (N_20147,N_19615,N_19724);
nand U20148 (N_20148,N_19467,N_19737);
xor U20149 (N_20149,N_19700,N_19552);
nor U20150 (N_20150,N_19566,N_19561);
or U20151 (N_20151,N_19945,N_19997);
xnor U20152 (N_20152,N_19690,N_19695);
nand U20153 (N_20153,N_19944,N_19589);
and U20154 (N_20154,N_19736,N_19906);
xnor U20155 (N_20155,N_19807,N_19590);
nand U20156 (N_20156,N_19718,N_19680);
nor U20157 (N_20157,N_19477,N_19651);
nand U20158 (N_20158,N_19974,N_19893);
xor U20159 (N_20159,N_19769,N_19716);
nand U20160 (N_20160,N_19495,N_19683);
nand U20161 (N_20161,N_19537,N_19949);
nor U20162 (N_20162,N_19454,N_19572);
xnor U20163 (N_20163,N_19781,N_19531);
nor U20164 (N_20164,N_19993,N_19871);
xnor U20165 (N_20165,N_19883,N_19384);
and U20166 (N_20166,N_19496,N_19834);
or U20167 (N_20167,N_19961,N_19659);
and U20168 (N_20168,N_19521,N_19459);
and U20169 (N_20169,N_19578,N_19745);
nor U20170 (N_20170,N_19729,N_19782);
or U20171 (N_20171,N_19481,N_19938);
and U20172 (N_20172,N_19875,N_19733);
xnor U20173 (N_20173,N_19392,N_19421);
nor U20174 (N_20174,N_19998,N_19409);
nand U20175 (N_20175,N_19940,N_19515);
xor U20176 (N_20176,N_19748,N_19582);
xnor U20177 (N_20177,N_19535,N_19765);
xnor U20178 (N_20178,N_19579,N_19387);
xor U20179 (N_20179,N_19739,N_19869);
xnor U20180 (N_20180,N_19990,N_19403);
xor U20181 (N_20181,N_19638,N_19630);
nor U20182 (N_20182,N_19402,N_19399);
xor U20183 (N_20183,N_19482,N_19907);
and U20184 (N_20184,N_19412,N_19476);
nand U20185 (N_20185,N_19464,N_19468);
nand U20186 (N_20186,N_19661,N_19854);
nor U20187 (N_20187,N_19756,N_19388);
or U20188 (N_20188,N_19629,N_19385);
nand U20189 (N_20189,N_19730,N_19776);
and U20190 (N_20190,N_19946,N_19723);
or U20191 (N_20191,N_19663,N_19442);
xnor U20192 (N_20192,N_19611,N_19698);
nor U20193 (N_20193,N_19977,N_19445);
nor U20194 (N_20194,N_19888,N_19943);
xor U20195 (N_20195,N_19708,N_19992);
nor U20196 (N_20196,N_19559,N_19682);
nor U20197 (N_20197,N_19792,N_19473);
or U20198 (N_20198,N_19434,N_19475);
or U20199 (N_20199,N_19747,N_19752);
or U20200 (N_20200,N_19632,N_19509);
and U20201 (N_20201,N_19705,N_19560);
and U20202 (N_20202,N_19848,N_19562);
and U20203 (N_20203,N_19573,N_19808);
nand U20204 (N_20204,N_19768,N_19882);
and U20205 (N_20205,N_19720,N_19955);
or U20206 (N_20206,N_19494,N_19926);
nor U20207 (N_20207,N_19414,N_19701);
and U20208 (N_20208,N_19839,N_19894);
nand U20209 (N_20209,N_19932,N_19985);
nor U20210 (N_20210,N_19606,N_19783);
and U20211 (N_20211,N_19966,N_19617);
xor U20212 (N_20212,N_19850,N_19841);
nand U20213 (N_20213,N_19852,N_19510);
xnor U20214 (N_20214,N_19607,N_19684);
or U20215 (N_20215,N_19443,N_19603);
or U20216 (N_20216,N_19920,N_19437);
xor U20217 (N_20217,N_19859,N_19623);
or U20218 (N_20218,N_19524,N_19948);
and U20219 (N_20219,N_19640,N_19986);
and U20220 (N_20220,N_19435,N_19398);
nand U20221 (N_20221,N_19395,N_19424);
nand U20222 (N_20222,N_19664,N_19879);
or U20223 (N_20223,N_19873,N_19764);
xnor U20224 (N_20224,N_19646,N_19795);
or U20225 (N_20225,N_19596,N_19732);
and U20226 (N_20226,N_19687,N_19953);
and U20227 (N_20227,N_19598,N_19862);
and U20228 (N_20228,N_19575,N_19431);
and U20229 (N_20229,N_19771,N_19984);
nor U20230 (N_20230,N_19505,N_19952);
nor U20231 (N_20231,N_19418,N_19497);
and U20232 (N_20232,N_19766,N_19872);
nand U20233 (N_20233,N_19849,N_19548);
or U20234 (N_20234,N_19833,N_19731);
nand U20235 (N_20235,N_19576,N_19545);
nand U20236 (N_20236,N_19438,N_19706);
nor U20237 (N_20237,N_19543,N_19451);
xor U20238 (N_20238,N_19877,N_19710);
nand U20239 (N_20239,N_19539,N_19868);
nor U20240 (N_20240,N_19627,N_19406);
nand U20241 (N_20241,N_19455,N_19767);
or U20242 (N_20242,N_19793,N_19714);
and U20243 (N_20243,N_19751,N_19853);
and U20244 (N_20244,N_19963,N_19677);
nand U20245 (N_20245,N_19939,N_19432);
xor U20246 (N_20246,N_19788,N_19654);
nor U20247 (N_20247,N_19800,N_19672);
and U20248 (N_20248,N_19884,N_19864);
and U20249 (N_20249,N_19461,N_19891);
nor U20250 (N_20250,N_19772,N_19656);
or U20251 (N_20251,N_19420,N_19816);
and U20252 (N_20252,N_19802,N_19962);
nor U20253 (N_20253,N_19794,N_19679);
nor U20254 (N_20254,N_19915,N_19994);
nand U20255 (N_20255,N_19422,N_19542);
and U20256 (N_20256,N_19688,N_19429);
or U20257 (N_20257,N_19597,N_19981);
nor U20258 (N_20258,N_19436,N_19858);
and U20259 (N_20259,N_19717,N_19826);
or U20260 (N_20260,N_19586,N_19639);
or U20261 (N_20261,N_19666,N_19842);
or U20262 (N_20262,N_19825,N_19928);
xor U20263 (N_20263,N_19631,N_19713);
xnor U20264 (N_20264,N_19914,N_19693);
and U20265 (N_20265,N_19774,N_19660);
nor U20266 (N_20266,N_19668,N_19866);
and U20267 (N_20267,N_19484,N_19441);
xnor U20268 (N_20268,N_19874,N_19812);
xor U20269 (N_20269,N_19978,N_19956);
and U20270 (N_20270,N_19379,N_19887);
nor U20271 (N_20271,N_19813,N_19671);
xnor U20272 (N_20272,N_19472,N_19609);
xor U20273 (N_20273,N_19796,N_19662);
nand U20274 (N_20274,N_19991,N_19727);
nand U20275 (N_20275,N_19601,N_19805);
and U20276 (N_20276,N_19401,N_19921);
or U20277 (N_20277,N_19567,N_19975);
nand U20278 (N_20278,N_19927,N_19620);
nor U20279 (N_20279,N_19965,N_19512);
nor U20280 (N_20280,N_19885,N_19456);
nor U20281 (N_20281,N_19516,N_19650);
nor U20282 (N_20282,N_19669,N_19863);
and U20283 (N_20283,N_19525,N_19790);
nor U20284 (N_20284,N_19618,N_19711);
nor U20285 (N_20285,N_19811,N_19773);
and U20286 (N_20286,N_19837,N_19715);
and U20287 (N_20287,N_19529,N_19838);
nand U20288 (N_20288,N_19844,N_19444);
or U20289 (N_20289,N_19778,N_19886);
xor U20290 (N_20290,N_19416,N_19754);
nor U20291 (N_20291,N_19488,N_19520);
and U20292 (N_20292,N_19470,N_19478);
nand U20293 (N_20293,N_19696,N_19798);
xor U20294 (N_20294,N_19390,N_19964);
xor U20295 (N_20295,N_19376,N_19657);
nand U20296 (N_20296,N_19605,N_19845);
and U20297 (N_20297,N_19563,N_19534);
xor U20298 (N_20298,N_19513,N_19500);
xor U20299 (N_20299,N_19702,N_19649);
and U20300 (N_20300,N_19942,N_19830);
nor U20301 (N_20301,N_19480,N_19637);
nand U20302 (N_20302,N_19824,N_19585);
nand U20303 (N_20303,N_19523,N_19426);
or U20304 (N_20304,N_19810,N_19999);
nor U20305 (N_20305,N_19433,N_19428);
nand U20306 (N_20306,N_19892,N_19924);
or U20307 (N_20307,N_19549,N_19753);
or U20308 (N_20308,N_19583,N_19670);
or U20309 (N_20309,N_19819,N_19465);
nor U20310 (N_20310,N_19635,N_19569);
nor U20311 (N_20311,N_19544,N_19501);
nor U20312 (N_20312,N_19407,N_19574);
xnor U20313 (N_20313,N_19587,N_19418);
nand U20314 (N_20314,N_19498,N_19606);
and U20315 (N_20315,N_19605,N_19579);
xor U20316 (N_20316,N_19968,N_19385);
and U20317 (N_20317,N_19949,N_19897);
or U20318 (N_20318,N_19385,N_19421);
and U20319 (N_20319,N_19643,N_19907);
nand U20320 (N_20320,N_19676,N_19651);
nor U20321 (N_20321,N_19682,N_19821);
xnor U20322 (N_20322,N_19473,N_19767);
or U20323 (N_20323,N_19957,N_19962);
or U20324 (N_20324,N_19756,N_19485);
and U20325 (N_20325,N_19405,N_19959);
nor U20326 (N_20326,N_19621,N_19842);
nand U20327 (N_20327,N_19383,N_19702);
or U20328 (N_20328,N_19414,N_19412);
nand U20329 (N_20329,N_19537,N_19518);
nor U20330 (N_20330,N_19682,N_19481);
nand U20331 (N_20331,N_19833,N_19865);
xnor U20332 (N_20332,N_19728,N_19430);
or U20333 (N_20333,N_19818,N_19843);
nor U20334 (N_20334,N_19679,N_19658);
or U20335 (N_20335,N_19487,N_19954);
and U20336 (N_20336,N_19620,N_19418);
and U20337 (N_20337,N_19630,N_19827);
nor U20338 (N_20338,N_19942,N_19606);
or U20339 (N_20339,N_19774,N_19598);
or U20340 (N_20340,N_19997,N_19600);
nor U20341 (N_20341,N_19581,N_19785);
and U20342 (N_20342,N_19883,N_19872);
xor U20343 (N_20343,N_19472,N_19792);
nand U20344 (N_20344,N_19659,N_19700);
or U20345 (N_20345,N_19509,N_19702);
and U20346 (N_20346,N_19659,N_19646);
or U20347 (N_20347,N_19682,N_19460);
nor U20348 (N_20348,N_19957,N_19619);
or U20349 (N_20349,N_19531,N_19740);
and U20350 (N_20350,N_19550,N_19596);
nor U20351 (N_20351,N_19975,N_19523);
xor U20352 (N_20352,N_19464,N_19771);
nor U20353 (N_20353,N_19886,N_19674);
and U20354 (N_20354,N_19949,N_19707);
xor U20355 (N_20355,N_19682,N_19602);
or U20356 (N_20356,N_19464,N_19952);
nor U20357 (N_20357,N_19679,N_19552);
nand U20358 (N_20358,N_19563,N_19633);
xnor U20359 (N_20359,N_19979,N_19576);
nand U20360 (N_20360,N_19725,N_19939);
or U20361 (N_20361,N_19477,N_19394);
nand U20362 (N_20362,N_19948,N_19778);
and U20363 (N_20363,N_19714,N_19927);
and U20364 (N_20364,N_19571,N_19656);
xnor U20365 (N_20365,N_19449,N_19768);
and U20366 (N_20366,N_19738,N_19412);
nor U20367 (N_20367,N_19496,N_19845);
xnor U20368 (N_20368,N_19673,N_19382);
and U20369 (N_20369,N_19401,N_19731);
nand U20370 (N_20370,N_19404,N_19397);
or U20371 (N_20371,N_19989,N_19762);
and U20372 (N_20372,N_19847,N_19505);
xor U20373 (N_20373,N_19718,N_19467);
nor U20374 (N_20374,N_19599,N_19726);
and U20375 (N_20375,N_19824,N_19445);
nand U20376 (N_20376,N_19579,N_19678);
nand U20377 (N_20377,N_19960,N_19516);
nand U20378 (N_20378,N_19928,N_19803);
nand U20379 (N_20379,N_19773,N_19446);
and U20380 (N_20380,N_19507,N_19812);
nand U20381 (N_20381,N_19379,N_19501);
and U20382 (N_20382,N_19607,N_19540);
and U20383 (N_20383,N_19395,N_19621);
nand U20384 (N_20384,N_19704,N_19392);
nand U20385 (N_20385,N_19848,N_19867);
nor U20386 (N_20386,N_19550,N_19488);
xor U20387 (N_20387,N_19570,N_19593);
and U20388 (N_20388,N_19507,N_19994);
or U20389 (N_20389,N_19389,N_19584);
xnor U20390 (N_20390,N_19967,N_19874);
nand U20391 (N_20391,N_19757,N_19452);
nor U20392 (N_20392,N_19556,N_19525);
xnor U20393 (N_20393,N_19636,N_19613);
xor U20394 (N_20394,N_19953,N_19474);
nand U20395 (N_20395,N_19766,N_19746);
nor U20396 (N_20396,N_19908,N_19762);
xnor U20397 (N_20397,N_19607,N_19829);
nor U20398 (N_20398,N_19671,N_19789);
nor U20399 (N_20399,N_19461,N_19900);
and U20400 (N_20400,N_19557,N_19715);
nor U20401 (N_20401,N_19389,N_19399);
nand U20402 (N_20402,N_19813,N_19495);
nor U20403 (N_20403,N_19536,N_19898);
and U20404 (N_20404,N_19907,N_19722);
and U20405 (N_20405,N_19683,N_19383);
nor U20406 (N_20406,N_19706,N_19537);
nor U20407 (N_20407,N_19972,N_19760);
nand U20408 (N_20408,N_19463,N_19799);
and U20409 (N_20409,N_19618,N_19480);
nand U20410 (N_20410,N_19723,N_19567);
or U20411 (N_20411,N_19810,N_19545);
or U20412 (N_20412,N_19634,N_19703);
nand U20413 (N_20413,N_19843,N_19663);
nand U20414 (N_20414,N_19445,N_19762);
nor U20415 (N_20415,N_19889,N_19717);
xor U20416 (N_20416,N_19408,N_19932);
or U20417 (N_20417,N_19497,N_19545);
and U20418 (N_20418,N_19998,N_19382);
nand U20419 (N_20419,N_19385,N_19460);
or U20420 (N_20420,N_19987,N_19616);
and U20421 (N_20421,N_19649,N_19404);
nor U20422 (N_20422,N_19434,N_19829);
nor U20423 (N_20423,N_19977,N_19739);
nand U20424 (N_20424,N_19654,N_19578);
and U20425 (N_20425,N_19626,N_19702);
xor U20426 (N_20426,N_19476,N_19497);
and U20427 (N_20427,N_19995,N_19713);
or U20428 (N_20428,N_19423,N_19998);
nor U20429 (N_20429,N_19432,N_19842);
xor U20430 (N_20430,N_19966,N_19465);
xnor U20431 (N_20431,N_19491,N_19772);
xnor U20432 (N_20432,N_19577,N_19730);
and U20433 (N_20433,N_19644,N_19857);
xnor U20434 (N_20434,N_19668,N_19422);
nor U20435 (N_20435,N_19897,N_19647);
and U20436 (N_20436,N_19899,N_19483);
and U20437 (N_20437,N_19694,N_19525);
xor U20438 (N_20438,N_19794,N_19709);
and U20439 (N_20439,N_19555,N_19559);
and U20440 (N_20440,N_19482,N_19952);
or U20441 (N_20441,N_19990,N_19722);
or U20442 (N_20442,N_19704,N_19986);
and U20443 (N_20443,N_19732,N_19696);
nand U20444 (N_20444,N_19380,N_19577);
nor U20445 (N_20445,N_19461,N_19465);
and U20446 (N_20446,N_19813,N_19959);
nor U20447 (N_20447,N_19583,N_19731);
and U20448 (N_20448,N_19539,N_19782);
nor U20449 (N_20449,N_19544,N_19478);
or U20450 (N_20450,N_19496,N_19732);
or U20451 (N_20451,N_19610,N_19957);
xor U20452 (N_20452,N_19864,N_19734);
or U20453 (N_20453,N_19492,N_19552);
xnor U20454 (N_20454,N_19583,N_19413);
xor U20455 (N_20455,N_19422,N_19855);
and U20456 (N_20456,N_19979,N_19792);
or U20457 (N_20457,N_19679,N_19772);
or U20458 (N_20458,N_19393,N_19643);
or U20459 (N_20459,N_19420,N_19528);
or U20460 (N_20460,N_19447,N_19566);
or U20461 (N_20461,N_19717,N_19734);
xnor U20462 (N_20462,N_19442,N_19383);
nand U20463 (N_20463,N_19533,N_19823);
nor U20464 (N_20464,N_19619,N_19821);
nor U20465 (N_20465,N_19601,N_19515);
nand U20466 (N_20466,N_19794,N_19941);
or U20467 (N_20467,N_19375,N_19911);
or U20468 (N_20468,N_19708,N_19721);
nor U20469 (N_20469,N_19955,N_19534);
xnor U20470 (N_20470,N_19720,N_19808);
xor U20471 (N_20471,N_19999,N_19484);
nor U20472 (N_20472,N_19981,N_19406);
nor U20473 (N_20473,N_19752,N_19980);
nand U20474 (N_20474,N_19647,N_19621);
xor U20475 (N_20475,N_19433,N_19634);
or U20476 (N_20476,N_19726,N_19523);
and U20477 (N_20477,N_19453,N_19722);
or U20478 (N_20478,N_19838,N_19479);
nand U20479 (N_20479,N_19926,N_19912);
or U20480 (N_20480,N_19757,N_19748);
and U20481 (N_20481,N_19982,N_19640);
nor U20482 (N_20482,N_19665,N_19997);
xnor U20483 (N_20483,N_19755,N_19567);
nand U20484 (N_20484,N_19730,N_19490);
or U20485 (N_20485,N_19494,N_19508);
and U20486 (N_20486,N_19862,N_19511);
or U20487 (N_20487,N_19659,N_19550);
xor U20488 (N_20488,N_19800,N_19461);
or U20489 (N_20489,N_19591,N_19747);
and U20490 (N_20490,N_19797,N_19660);
xnor U20491 (N_20491,N_19375,N_19776);
nand U20492 (N_20492,N_19841,N_19833);
nor U20493 (N_20493,N_19382,N_19981);
nor U20494 (N_20494,N_19679,N_19731);
and U20495 (N_20495,N_19836,N_19609);
and U20496 (N_20496,N_19947,N_19383);
nand U20497 (N_20497,N_19474,N_19763);
nand U20498 (N_20498,N_19771,N_19606);
or U20499 (N_20499,N_19807,N_19402);
xor U20500 (N_20500,N_19619,N_19782);
nor U20501 (N_20501,N_19996,N_19496);
nor U20502 (N_20502,N_19849,N_19816);
or U20503 (N_20503,N_19472,N_19478);
nand U20504 (N_20504,N_19655,N_19724);
nor U20505 (N_20505,N_19934,N_19724);
and U20506 (N_20506,N_19955,N_19566);
and U20507 (N_20507,N_19939,N_19743);
xnor U20508 (N_20508,N_19665,N_19504);
or U20509 (N_20509,N_19447,N_19472);
or U20510 (N_20510,N_19857,N_19696);
nor U20511 (N_20511,N_19531,N_19537);
nand U20512 (N_20512,N_19630,N_19383);
nor U20513 (N_20513,N_19833,N_19938);
nor U20514 (N_20514,N_19570,N_19590);
nand U20515 (N_20515,N_19998,N_19550);
nand U20516 (N_20516,N_19502,N_19623);
nor U20517 (N_20517,N_19594,N_19384);
nand U20518 (N_20518,N_19830,N_19715);
nor U20519 (N_20519,N_19671,N_19487);
or U20520 (N_20520,N_19694,N_19679);
nor U20521 (N_20521,N_19781,N_19900);
or U20522 (N_20522,N_19890,N_19899);
and U20523 (N_20523,N_19775,N_19463);
and U20524 (N_20524,N_19503,N_19971);
xor U20525 (N_20525,N_19847,N_19454);
nand U20526 (N_20526,N_19757,N_19604);
nor U20527 (N_20527,N_19970,N_19385);
or U20528 (N_20528,N_19502,N_19962);
nand U20529 (N_20529,N_19985,N_19466);
and U20530 (N_20530,N_19976,N_19640);
xor U20531 (N_20531,N_19492,N_19981);
xor U20532 (N_20532,N_19508,N_19884);
nand U20533 (N_20533,N_19731,N_19903);
or U20534 (N_20534,N_19739,N_19428);
nand U20535 (N_20535,N_19959,N_19459);
and U20536 (N_20536,N_19612,N_19421);
nor U20537 (N_20537,N_19460,N_19892);
and U20538 (N_20538,N_19599,N_19944);
or U20539 (N_20539,N_19681,N_19492);
nor U20540 (N_20540,N_19420,N_19697);
and U20541 (N_20541,N_19747,N_19845);
xnor U20542 (N_20542,N_19545,N_19559);
nor U20543 (N_20543,N_19758,N_19944);
and U20544 (N_20544,N_19660,N_19636);
or U20545 (N_20545,N_19608,N_19747);
xor U20546 (N_20546,N_19680,N_19811);
nand U20547 (N_20547,N_19659,N_19620);
and U20548 (N_20548,N_19621,N_19556);
nand U20549 (N_20549,N_19978,N_19778);
and U20550 (N_20550,N_19568,N_19937);
and U20551 (N_20551,N_19738,N_19927);
and U20552 (N_20552,N_19811,N_19474);
xnor U20553 (N_20553,N_19899,N_19922);
xnor U20554 (N_20554,N_19896,N_19525);
nor U20555 (N_20555,N_19523,N_19375);
or U20556 (N_20556,N_19855,N_19741);
nor U20557 (N_20557,N_19723,N_19593);
or U20558 (N_20558,N_19628,N_19625);
and U20559 (N_20559,N_19422,N_19948);
or U20560 (N_20560,N_19652,N_19568);
or U20561 (N_20561,N_19947,N_19746);
nor U20562 (N_20562,N_19859,N_19812);
nand U20563 (N_20563,N_19882,N_19783);
or U20564 (N_20564,N_19421,N_19922);
nor U20565 (N_20565,N_19677,N_19800);
nand U20566 (N_20566,N_19873,N_19742);
nor U20567 (N_20567,N_19769,N_19968);
nor U20568 (N_20568,N_19863,N_19883);
or U20569 (N_20569,N_19651,N_19476);
and U20570 (N_20570,N_19611,N_19865);
nand U20571 (N_20571,N_19953,N_19735);
nand U20572 (N_20572,N_19612,N_19628);
nor U20573 (N_20573,N_19563,N_19384);
or U20574 (N_20574,N_19505,N_19446);
nor U20575 (N_20575,N_19663,N_19385);
nor U20576 (N_20576,N_19783,N_19962);
and U20577 (N_20577,N_19875,N_19887);
or U20578 (N_20578,N_19910,N_19586);
or U20579 (N_20579,N_19931,N_19404);
nor U20580 (N_20580,N_19959,N_19656);
or U20581 (N_20581,N_19866,N_19630);
nor U20582 (N_20582,N_19733,N_19852);
and U20583 (N_20583,N_19939,N_19505);
or U20584 (N_20584,N_19633,N_19930);
nor U20585 (N_20585,N_19508,N_19511);
xnor U20586 (N_20586,N_19690,N_19903);
or U20587 (N_20587,N_19968,N_19900);
or U20588 (N_20588,N_19591,N_19393);
xor U20589 (N_20589,N_19942,N_19899);
and U20590 (N_20590,N_19693,N_19650);
nor U20591 (N_20591,N_19781,N_19867);
nor U20592 (N_20592,N_19842,N_19643);
nand U20593 (N_20593,N_19630,N_19903);
xor U20594 (N_20594,N_19608,N_19949);
and U20595 (N_20595,N_19820,N_19775);
or U20596 (N_20596,N_19589,N_19567);
xnor U20597 (N_20597,N_19694,N_19984);
or U20598 (N_20598,N_19702,N_19825);
nor U20599 (N_20599,N_19789,N_19662);
nand U20600 (N_20600,N_19479,N_19885);
nor U20601 (N_20601,N_19926,N_19454);
or U20602 (N_20602,N_19990,N_19655);
nand U20603 (N_20603,N_19580,N_19476);
nor U20604 (N_20604,N_19956,N_19684);
nor U20605 (N_20605,N_19802,N_19581);
and U20606 (N_20606,N_19944,N_19905);
and U20607 (N_20607,N_19911,N_19903);
nand U20608 (N_20608,N_19428,N_19414);
or U20609 (N_20609,N_19980,N_19459);
nor U20610 (N_20610,N_19575,N_19806);
nor U20611 (N_20611,N_19576,N_19510);
nand U20612 (N_20612,N_19747,N_19500);
and U20613 (N_20613,N_19417,N_19635);
xor U20614 (N_20614,N_19899,N_19674);
nand U20615 (N_20615,N_19572,N_19967);
and U20616 (N_20616,N_19478,N_19848);
nor U20617 (N_20617,N_19759,N_19544);
xnor U20618 (N_20618,N_19446,N_19898);
nand U20619 (N_20619,N_19876,N_19416);
or U20620 (N_20620,N_19458,N_19566);
nor U20621 (N_20621,N_19594,N_19861);
nand U20622 (N_20622,N_19618,N_19973);
nand U20623 (N_20623,N_19489,N_19568);
nand U20624 (N_20624,N_19587,N_19379);
nor U20625 (N_20625,N_20399,N_20514);
and U20626 (N_20626,N_20216,N_20576);
nand U20627 (N_20627,N_20362,N_20104);
and U20628 (N_20628,N_20616,N_20419);
nor U20629 (N_20629,N_20081,N_20134);
or U20630 (N_20630,N_20332,N_20085);
and U20631 (N_20631,N_20129,N_20249);
and U20632 (N_20632,N_20619,N_20184);
nor U20633 (N_20633,N_20586,N_20388);
nor U20634 (N_20634,N_20029,N_20326);
and U20635 (N_20635,N_20014,N_20527);
or U20636 (N_20636,N_20491,N_20082);
nor U20637 (N_20637,N_20079,N_20435);
nand U20638 (N_20638,N_20267,N_20522);
nor U20639 (N_20639,N_20109,N_20177);
and U20640 (N_20640,N_20568,N_20260);
xor U20641 (N_20641,N_20263,N_20063);
nand U20642 (N_20642,N_20212,N_20463);
or U20643 (N_20643,N_20307,N_20441);
nand U20644 (N_20644,N_20349,N_20154);
nor U20645 (N_20645,N_20116,N_20484);
nand U20646 (N_20646,N_20203,N_20471);
or U20647 (N_20647,N_20164,N_20380);
or U20648 (N_20648,N_20169,N_20246);
or U20649 (N_20649,N_20004,N_20548);
or U20650 (N_20650,N_20204,N_20453);
nand U20651 (N_20651,N_20052,N_20523);
nand U20652 (N_20652,N_20254,N_20364);
xor U20653 (N_20653,N_20108,N_20353);
or U20654 (N_20654,N_20042,N_20341);
nor U20655 (N_20655,N_20077,N_20464);
nand U20656 (N_20656,N_20274,N_20377);
and U20657 (N_20657,N_20327,N_20221);
xnor U20658 (N_20658,N_20596,N_20456);
and U20659 (N_20659,N_20028,N_20288);
xor U20660 (N_20660,N_20336,N_20444);
nor U20661 (N_20661,N_20386,N_20232);
and U20662 (N_20662,N_20525,N_20229);
nand U20663 (N_20663,N_20334,N_20322);
and U20664 (N_20664,N_20037,N_20241);
or U20665 (N_20665,N_20240,N_20546);
nor U20666 (N_20666,N_20436,N_20613);
or U20667 (N_20667,N_20478,N_20496);
and U20668 (N_20668,N_20461,N_20121);
or U20669 (N_20669,N_20114,N_20558);
xor U20670 (N_20670,N_20188,N_20163);
or U20671 (N_20671,N_20252,N_20292);
or U20672 (N_20672,N_20173,N_20495);
nor U20673 (N_20673,N_20166,N_20183);
nand U20674 (N_20674,N_20348,N_20107);
nor U20675 (N_20675,N_20617,N_20228);
or U20676 (N_20676,N_20595,N_20076);
xnor U20677 (N_20677,N_20505,N_20196);
xor U20678 (N_20678,N_20047,N_20370);
nor U20679 (N_20679,N_20090,N_20565);
nand U20680 (N_20680,N_20003,N_20499);
nor U20681 (N_20681,N_20128,N_20214);
xnor U20682 (N_20682,N_20224,N_20472);
xnor U20683 (N_20683,N_20497,N_20608);
nand U20684 (N_20684,N_20311,N_20536);
or U20685 (N_20685,N_20217,N_20567);
xnor U20686 (N_20686,N_20466,N_20160);
xnor U20687 (N_20687,N_20328,N_20507);
and U20688 (N_20688,N_20487,N_20226);
or U20689 (N_20689,N_20099,N_20598);
nand U20690 (N_20690,N_20285,N_20059);
nand U20691 (N_20691,N_20542,N_20331);
nand U20692 (N_20692,N_20513,N_20477);
or U20693 (N_20693,N_20137,N_20178);
or U20694 (N_20694,N_20279,N_20122);
or U20695 (N_20695,N_20033,N_20233);
xor U20696 (N_20696,N_20579,N_20300);
xor U20697 (N_20697,N_20385,N_20158);
xnor U20698 (N_20698,N_20281,N_20394);
xor U20699 (N_20699,N_20248,N_20208);
nand U20700 (N_20700,N_20105,N_20460);
and U20701 (N_20701,N_20492,N_20345);
nor U20702 (N_20702,N_20211,N_20430);
nor U20703 (N_20703,N_20193,N_20165);
nand U20704 (N_20704,N_20271,N_20272);
xnor U20705 (N_20705,N_20034,N_20594);
xor U20706 (N_20706,N_20395,N_20198);
and U20707 (N_20707,N_20044,N_20578);
or U20708 (N_20708,N_20131,N_20245);
and U20709 (N_20709,N_20575,N_20623);
nand U20710 (N_20710,N_20008,N_20438);
xor U20711 (N_20711,N_20482,N_20095);
nand U20712 (N_20712,N_20132,N_20220);
nor U20713 (N_20713,N_20058,N_20161);
xnor U20714 (N_20714,N_20309,N_20421);
or U20715 (N_20715,N_20148,N_20537);
or U20716 (N_20716,N_20553,N_20571);
nor U20717 (N_20717,N_20515,N_20045);
and U20718 (N_20718,N_20015,N_20084);
and U20719 (N_20719,N_20218,N_20144);
and U20720 (N_20720,N_20488,N_20053);
nand U20721 (N_20721,N_20367,N_20476);
nand U20722 (N_20722,N_20305,N_20019);
and U20723 (N_20723,N_20343,N_20383);
xnor U20724 (N_20724,N_20310,N_20175);
xor U20725 (N_20725,N_20040,N_20143);
and U20726 (N_20726,N_20428,N_20091);
nor U20727 (N_20727,N_20611,N_20573);
nor U20728 (N_20728,N_20206,N_20299);
xor U20729 (N_20729,N_20256,N_20602);
xnor U20730 (N_20730,N_20294,N_20470);
nor U20731 (N_20731,N_20335,N_20351);
xor U20732 (N_20732,N_20580,N_20247);
nand U20733 (N_20733,N_20168,N_20423);
and U20734 (N_20734,N_20321,N_20027);
nor U20735 (N_20735,N_20142,N_20100);
xnor U20736 (N_20736,N_20365,N_20133);
xor U20737 (N_20737,N_20315,N_20540);
xor U20738 (N_20738,N_20115,N_20006);
xor U20739 (N_20739,N_20469,N_20511);
nand U20740 (N_20740,N_20454,N_20250);
nor U20741 (N_20741,N_20396,N_20413);
nor U20742 (N_20742,N_20031,N_20219);
xnor U20743 (N_20743,N_20426,N_20170);
and U20744 (N_20744,N_20324,N_20518);
nand U20745 (N_20745,N_20439,N_20067);
or U20746 (N_20746,N_20140,N_20465);
or U20747 (N_20747,N_20519,N_20190);
xnor U20748 (N_20748,N_20582,N_20167);
nand U20749 (N_20749,N_20038,N_20237);
or U20750 (N_20750,N_20560,N_20201);
nor U20751 (N_20751,N_20360,N_20239);
nor U20752 (N_20752,N_20041,N_20411);
or U20753 (N_20753,N_20113,N_20024);
nor U20754 (N_20754,N_20480,N_20605);
or U20755 (N_20755,N_20127,N_20275);
nor U20756 (N_20756,N_20159,N_20251);
or U20757 (N_20757,N_20317,N_20117);
and U20758 (N_20758,N_20273,N_20624);
nor U20759 (N_20759,N_20500,N_20433);
and U20760 (N_20760,N_20032,N_20337);
nand U20761 (N_20761,N_20585,N_20384);
nor U20762 (N_20762,N_20185,N_20280);
and U20763 (N_20763,N_20347,N_20080);
nor U20764 (N_20764,N_20124,N_20389);
or U20765 (N_20765,N_20452,N_20025);
xnor U20766 (N_20766,N_20207,N_20431);
or U20767 (N_20767,N_20162,N_20012);
nor U20768 (N_20768,N_20236,N_20009);
or U20769 (N_20769,N_20179,N_20414);
and U20770 (N_20770,N_20528,N_20545);
or U20771 (N_20771,N_20401,N_20111);
nand U20772 (N_20772,N_20621,N_20570);
xnor U20773 (N_20773,N_20021,N_20533);
and U20774 (N_20774,N_20615,N_20535);
and U20775 (N_20775,N_20490,N_20330);
nor U20776 (N_20776,N_20287,N_20462);
nand U20777 (N_20777,N_20323,N_20001);
and U20778 (N_20778,N_20258,N_20412);
xor U20779 (N_20779,N_20342,N_20072);
nor U20780 (N_20780,N_20574,N_20308);
and U20781 (N_20781,N_20286,N_20510);
and U20782 (N_20782,N_20359,N_20096);
xnor U20783 (N_20783,N_20094,N_20151);
and U20784 (N_20784,N_20344,N_20136);
and U20785 (N_20785,N_20101,N_20358);
and U20786 (N_20786,N_20368,N_20126);
and U20787 (N_20787,N_20506,N_20340);
nand U20788 (N_20788,N_20225,N_20517);
nor U20789 (N_20789,N_20352,N_20564);
nor U20790 (N_20790,N_20410,N_20562);
xor U20791 (N_20791,N_20289,N_20603);
nor U20792 (N_20792,N_20516,N_20544);
xor U20793 (N_20793,N_20355,N_20123);
xnor U20794 (N_20794,N_20458,N_20120);
xor U20795 (N_20795,N_20375,N_20442);
nand U20796 (N_20796,N_20559,N_20422);
or U20797 (N_20797,N_20106,N_20152);
nor U20798 (N_20798,N_20155,N_20539);
nor U20799 (N_20799,N_20071,N_20093);
nor U20800 (N_20800,N_20209,N_20046);
or U20801 (N_20801,N_20291,N_20597);
and U20802 (N_20802,N_20073,N_20020);
nor U20803 (N_20803,N_20382,N_20538);
nor U20804 (N_20804,N_20083,N_20427);
nand U20805 (N_20805,N_20552,N_20607);
or U20806 (N_20806,N_20583,N_20023);
xnor U20807 (N_20807,N_20387,N_20504);
or U20808 (N_20808,N_20097,N_20405);
xnor U20809 (N_20809,N_20119,N_20103);
xnor U20810 (N_20810,N_20296,N_20282);
nor U20811 (N_20811,N_20056,N_20561);
nand U20812 (N_20812,N_20563,N_20443);
and U20813 (N_20813,N_20278,N_20325);
xnor U20814 (N_20814,N_20112,N_20489);
nand U20815 (N_20815,N_20264,N_20284);
and U20816 (N_20816,N_20534,N_20016);
xor U20817 (N_20817,N_20373,N_20622);
or U20818 (N_20818,N_20520,N_20261);
nor U20819 (N_20819,N_20593,N_20262);
nand U20820 (N_20820,N_20007,N_20521);
nand U20821 (N_20821,N_20210,N_20051);
nor U20822 (N_20822,N_20429,N_20147);
nor U20823 (N_20823,N_20529,N_20180);
xnor U20824 (N_20824,N_20145,N_20065);
nor U20825 (N_20825,N_20420,N_20393);
or U20826 (N_20826,N_20069,N_20609);
or U20827 (N_20827,N_20092,N_20205);
xor U20828 (N_20828,N_20054,N_20010);
xnor U20829 (N_20829,N_20587,N_20197);
xnor U20830 (N_20830,N_20588,N_20541);
and U20831 (N_20831,N_20242,N_20350);
nand U20832 (N_20832,N_20584,N_20473);
nand U20833 (N_20833,N_20153,N_20591);
or U20834 (N_20834,N_20366,N_20244);
nor U20835 (N_20835,N_20361,N_20475);
nor U20836 (N_20836,N_20234,N_20181);
nor U20837 (N_20837,N_20195,N_20074);
and U20838 (N_20838,N_20110,N_20118);
or U20839 (N_20839,N_20600,N_20599);
and U20840 (N_20840,N_20297,N_20416);
xor U20841 (N_20841,N_20610,N_20400);
or U20842 (N_20842,N_20057,N_20141);
xor U20843 (N_20843,N_20055,N_20374);
nand U20844 (N_20844,N_20277,N_20086);
and U20845 (N_20845,N_20526,N_20230);
xnor U20846 (N_20846,N_20138,N_20222);
nand U20847 (N_20847,N_20509,N_20298);
and U20848 (N_20848,N_20481,N_20479);
xnor U20849 (N_20849,N_20501,N_20030);
xnor U20850 (N_20850,N_20379,N_20089);
and U20851 (N_20851,N_20176,N_20356);
nor U20852 (N_20852,N_20457,N_20601);
or U20853 (N_20853,N_20449,N_20290);
and U20854 (N_20854,N_20171,N_20555);
nand U20855 (N_20855,N_20013,N_20199);
or U20856 (N_20856,N_20174,N_20146);
and U20857 (N_20857,N_20486,N_20318);
and U20858 (N_20858,N_20339,N_20455);
or U20859 (N_20859,N_20243,N_20532);
xor U20860 (N_20860,N_20397,N_20554);
and U20861 (N_20861,N_20022,N_20049);
and U20862 (N_20862,N_20172,N_20043);
nand U20863 (N_20863,N_20371,N_20149);
xnor U20864 (N_20864,N_20459,N_20446);
nand U20865 (N_20865,N_20606,N_20432);
xnor U20866 (N_20866,N_20451,N_20186);
nor U20867 (N_20867,N_20064,N_20139);
nor U20868 (N_20868,N_20550,N_20447);
and U20869 (N_20869,N_20313,N_20070);
nor U20870 (N_20870,N_20182,N_20235);
nand U20871 (N_20871,N_20039,N_20409);
or U20872 (N_20872,N_20036,N_20445);
nand U20873 (N_20873,N_20102,N_20440);
and U20874 (N_20874,N_20231,N_20075);
xor U20875 (N_20875,N_20376,N_20614);
nand U20876 (N_20876,N_20213,N_20403);
and U20877 (N_20877,N_20402,N_20130);
xnor U20878 (N_20878,N_20425,N_20238);
xnor U20879 (N_20879,N_20604,N_20581);
nand U20880 (N_20880,N_20406,N_20372);
nor U20881 (N_20881,N_20483,N_20088);
nand U20882 (N_20882,N_20391,N_20468);
or U20883 (N_20883,N_20276,N_20011);
and U20884 (N_20884,N_20078,N_20498);
xnor U20885 (N_20885,N_20590,N_20404);
or U20886 (N_20886,N_20061,N_20592);
and U20887 (N_20887,N_20191,N_20333);
nand U20888 (N_20888,N_20026,N_20531);
and U20889 (N_20889,N_20346,N_20398);
xnor U20890 (N_20890,N_20512,N_20194);
nor U20891 (N_20891,N_20485,N_20192);
xor U20892 (N_20892,N_20156,N_20316);
and U20893 (N_20893,N_20314,N_20612);
and U20894 (N_20894,N_20530,N_20303);
nor U20895 (N_20895,N_20467,N_20087);
or U20896 (N_20896,N_20474,N_20202);
and U20897 (N_20897,N_20551,N_20378);
nand U20898 (N_20898,N_20547,N_20189);
or U20899 (N_20899,N_20390,N_20524);
xor U20900 (N_20900,N_20255,N_20227);
or U20901 (N_20901,N_20266,N_20572);
and U20902 (N_20902,N_20259,N_20450);
nand U20903 (N_20903,N_20268,N_20618);
nor U20904 (N_20904,N_20257,N_20543);
and U20905 (N_20905,N_20508,N_20293);
xor U20906 (N_20906,N_20135,N_20295);
or U20907 (N_20907,N_20035,N_20493);
nor U20908 (N_20908,N_20503,N_20319);
xor U20909 (N_20909,N_20338,N_20329);
or U20910 (N_20910,N_20306,N_20018);
xnor U20911 (N_20911,N_20418,N_20304);
xor U20912 (N_20912,N_20270,N_20424);
or U20913 (N_20913,N_20566,N_20050);
nor U20914 (N_20914,N_20301,N_20620);
or U20915 (N_20915,N_20549,N_20068);
or U20916 (N_20916,N_20502,N_20150);
or U20917 (N_20917,N_20408,N_20000);
nor U20918 (N_20918,N_20312,N_20494);
nor U20919 (N_20919,N_20187,N_20569);
or U20920 (N_20920,N_20157,N_20269);
and U20921 (N_20921,N_20448,N_20556);
xor U20922 (N_20922,N_20415,N_20002);
nand U20923 (N_20923,N_20357,N_20283);
nand U20924 (N_20924,N_20060,N_20320);
nor U20925 (N_20925,N_20215,N_20066);
nor U20926 (N_20926,N_20005,N_20392);
nor U20927 (N_20927,N_20369,N_20048);
or U20928 (N_20928,N_20434,N_20200);
xnor U20929 (N_20929,N_20363,N_20577);
and U20930 (N_20930,N_20417,N_20098);
or U20931 (N_20931,N_20265,N_20125);
or U20932 (N_20932,N_20437,N_20589);
nand U20933 (N_20933,N_20407,N_20557);
xor U20934 (N_20934,N_20223,N_20062);
xnor U20935 (N_20935,N_20253,N_20381);
nor U20936 (N_20936,N_20354,N_20302);
xnor U20937 (N_20937,N_20017,N_20306);
nor U20938 (N_20938,N_20507,N_20607);
nand U20939 (N_20939,N_20149,N_20103);
nor U20940 (N_20940,N_20055,N_20150);
nand U20941 (N_20941,N_20291,N_20315);
nor U20942 (N_20942,N_20312,N_20541);
nand U20943 (N_20943,N_20016,N_20588);
nand U20944 (N_20944,N_20431,N_20376);
or U20945 (N_20945,N_20163,N_20514);
xor U20946 (N_20946,N_20197,N_20046);
and U20947 (N_20947,N_20497,N_20352);
or U20948 (N_20948,N_20620,N_20146);
nand U20949 (N_20949,N_20053,N_20031);
and U20950 (N_20950,N_20143,N_20162);
or U20951 (N_20951,N_20026,N_20392);
nor U20952 (N_20952,N_20382,N_20248);
xnor U20953 (N_20953,N_20229,N_20434);
and U20954 (N_20954,N_20342,N_20340);
and U20955 (N_20955,N_20275,N_20345);
and U20956 (N_20956,N_20522,N_20427);
nor U20957 (N_20957,N_20284,N_20127);
or U20958 (N_20958,N_20022,N_20324);
or U20959 (N_20959,N_20349,N_20550);
nand U20960 (N_20960,N_20601,N_20520);
or U20961 (N_20961,N_20165,N_20347);
or U20962 (N_20962,N_20067,N_20570);
nor U20963 (N_20963,N_20289,N_20562);
or U20964 (N_20964,N_20387,N_20109);
xor U20965 (N_20965,N_20569,N_20227);
or U20966 (N_20966,N_20014,N_20317);
nor U20967 (N_20967,N_20366,N_20415);
and U20968 (N_20968,N_20395,N_20041);
xnor U20969 (N_20969,N_20543,N_20368);
or U20970 (N_20970,N_20441,N_20480);
nor U20971 (N_20971,N_20488,N_20396);
or U20972 (N_20972,N_20040,N_20226);
nor U20973 (N_20973,N_20143,N_20303);
or U20974 (N_20974,N_20525,N_20024);
or U20975 (N_20975,N_20570,N_20252);
xnor U20976 (N_20976,N_20165,N_20091);
nor U20977 (N_20977,N_20191,N_20549);
nand U20978 (N_20978,N_20296,N_20410);
or U20979 (N_20979,N_20184,N_20530);
or U20980 (N_20980,N_20388,N_20095);
nand U20981 (N_20981,N_20214,N_20024);
or U20982 (N_20982,N_20175,N_20126);
xor U20983 (N_20983,N_20581,N_20423);
xor U20984 (N_20984,N_20561,N_20064);
and U20985 (N_20985,N_20173,N_20461);
xor U20986 (N_20986,N_20443,N_20336);
nor U20987 (N_20987,N_20428,N_20181);
or U20988 (N_20988,N_20085,N_20551);
and U20989 (N_20989,N_20142,N_20553);
or U20990 (N_20990,N_20139,N_20041);
and U20991 (N_20991,N_20336,N_20093);
or U20992 (N_20992,N_20258,N_20567);
nor U20993 (N_20993,N_20367,N_20168);
or U20994 (N_20994,N_20115,N_20082);
or U20995 (N_20995,N_20121,N_20213);
xnor U20996 (N_20996,N_20105,N_20322);
nand U20997 (N_20997,N_20275,N_20533);
or U20998 (N_20998,N_20046,N_20269);
and U20999 (N_20999,N_20441,N_20041);
and U21000 (N_21000,N_20413,N_20346);
or U21001 (N_21001,N_20185,N_20141);
or U21002 (N_21002,N_20171,N_20617);
or U21003 (N_21003,N_20162,N_20283);
or U21004 (N_21004,N_20436,N_20597);
nand U21005 (N_21005,N_20112,N_20465);
or U21006 (N_21006,N_20300,N_20513);
nand U21007 (N_21007,N_20601,N_20272);
xor U21008 (N_21008,N_20479,N_20399);
or U21009 (N_21009,N_20495,N_20179);
and U21010 (N_21010,N_20229,N_20198);
nand U21011 (N_21011,N_20203,N_20566);
nand U21012 (N_21012,N_20607,N_20223);
nand U21013 (N_21013,N_20266,N_20211);
xor U21014 (N_21014,N_20254,N_20466);
and U21015 (N_21015,N_20157,N_20422);
or U21016 (N_21016,N_20197,N_20474);
or U21017 (N_21017,N_20352,N_20436);
nor U21018 (N_21018,N_20498,N_20489);
xnor U21019 (N_21019,N_20134,N_20455);
or U21020 (N_21020,N_20624,N_20109);
xnor U21021 (N_21021,N_20176,N_20354);
xnor U21022 (N_21022,N_20238,N_20401);
or U21023 (N_21023,N_20454,N_20487);
or U21024 (N_21024,N_20058,N_20415);
nor U21025 (N_21025,N_20601,N_20247);
xnor U21026 (N_21026,N_20236,N_20375);
xnor U21027 (N_21027,N_20124,N_20291);
or U21028 (N_21028,N_20495,N_20169);
and U21029 (N_21029,N_20452,N_20559);
or U21030 (N_21030,N_20400,N_20282);
or U21031 (N_21031,N_20538,N_20394);
or U21032 (N_21032,N_20465,N_20081);
nand U21033 (N_21033,N_20063,N_20402);
or U21034 (N_21034,N_20411,N_20173);
or U21035 (N_21035,N_20362,N_20118);
xnor U21036 (N_21036,N_20598,N_20058);
nand U21037 (N_21037,N_20486,N_20599);
or U21038 (N_21038,N_20432,N_20482);
or U21039 (N_21039,N_20347,N_20425);
nand U21040 (N_21040,N_20119,N_20065);
or U21041 (N_21041,N_20109,N_20455);
xor U21042 (N_21042,N_20501,N_20359);
nor U21043 (N_21043,N_20253,N_20149);
or U21044 (N_21044,N_20124,N_20408);
nor U21045 (N_21045,N_20119,N_20507);
or U21046 (N_21046,N_20489,N_20356);
xnor U21047 (N_21047,N_20221,N_20116);
nand U21048 (N_21048,N_20439,N_20001);
xor U21049 (N_21049,N_20300,N_20420);
or U21050 (N_21050,N_20183,N_20575);
nor U21051 (N_21051,N_20468,N_20155);
xnor U21052 (N_21052,N_20551,N_20162);
nor U21053 (N_21053,N_20498,N_20210);
nor U21054 (N_21054,N_20368,N_20148);
and U21055 (N_21055,N_20159,N_20600);
nand U21056 (N_21056,N_20490,N_20578);
and U21057 (N_21057,N_20462,N_20337);
xor U21058 (N_21058,N_20125,N_20072);
or U21059 (N_21059,N_20131,N_20453);
xnor U21060 (N_21060,N_20374,N_20570);
and U21061 (N_21061,N_20496,N_20366);
nor U21062 (N_21062,N_20621,N_20003);
or U21063 (N_21063,N_20173,N_20474);
or U21064 (N_21064,N_20464,N_20241);
xor U21065 (N_21065,N_20176,N_20230);
and U21066 (N_21066,N_20084,N_20542);
xnor U21067 (N_21067,N_20189,N_20494);
or U21068 (N_21068,N_20601,N_20523);
xor U21069 (N_21069,N_20297,N_20601);
or U21070 (N_21070,N_20202,N_20127);
xor U21071 (N_21071,N_20042,N_20079);
xnor U21072 (N_21072,N_20622,N_20016);
xnor U21073 (N_21073,N_20498,N_20618);
nand U21074 (N_21074,N_20268,N_20613);
nor U21075 (N_21075,N_20301,N_20005);
or U21076 (N_21076,N_20464,N_20368);
and U21077 (N_21077,N_20047,N_20616);
and U21078 (N_21078,N_20515,N_20552);
nand U21079 (N_21079,N_20304,N_20354);
and U21080 (N_21080,N_20123,N_20541);
nor U21081 (N_21081,N_20395,N_20276);
and U21082 (N_21082,N_20512,N_20493);
nor U21083 (N_21083,N_20553,N_20580);
and U21084 (N_21084,N_20558,N_20176);
or U21085 (N_21085,N_20317,N_20174);
or U21086 (N_21086,N_20546,N_20439);
xor U21087 (N_21087,N_20552,N_20040);
nor U21088 (N_21088,N_20217,N_20152);
xnor U21089 (N_21089,N_20166,N_20357);
or U21090 (N_21090,N_20079,N_20205);
xnor U21091 (N_21091,N_20588,N_20139);
or U21092 (N_21092,N_20558,N_20404);
xor U21093 (N_21093,N_20357,N_20310);
xor U21094 (N_21094,N_20161,N_20501);
xor U21095 (N_21095,N_20601,N_20439);
nor U21096 (N_21096,N_20501,N_20022);
and U21097 (N_21097,N_20080,N_20079);
nand U21098 (N_21098,N_20617,N_20208);
or U21099 (N_21099,N_20229,N_20596);
or U21100 (N_21100,N_20589,N_20311);
nor U21101 (N_21101,N_20568,N_20054);
or U21102 (N_21102,N_20530,N_20572);
nor U21103 (N_21103,N_20612,N_20138);
and U21104 (N_21104,N_20566,N_20145);
xor U21105 (N_21105,N_20414,N_20305);
nand U21106 (N_21106,N_20480,N_20075);
nor U21107 (N_21107,N_20462,N_20174);
nand U21108 (N_21108,N_20103,N_20309);
and U21109 (N_21109,N_20479,N_20195);
xnor U21110 (N_21110,N_20168,N_20007);
or U21111 (N_21111,N_20512,N_20581);
or U21112 (N_21112,N_20399,N_20620);
nor U21113 (N_21113,N_20548,N_20361);
nand U21114 (N_21114,N_20482,N_20544);
xnor U21115 (N_21115,N_20307,N_20314);
xnor U21116 (N_21116,N_20543,N_20280);
nor U21117 (N_21117,N_20199,N_20196);
xnor U21118 (N_21118,N_20265,N_20024);
nor U21119 (N_21119,N_20166,N_20164);
nand U21120 (N_21120,N_20528,N_20360);
and U21121 (N_21121,N_20187,N_20394);
nor U21122 (N_21122,N_20274,N_20281);
and U21123 (N_21123,N_20262,N_20330);
and U21124 (N_21124,N_20294,N_20342);
nand U21125 (N_21125,N_20448,N_20046);
or U21126 (N_21126,N_20036,N_20111);
nor U21127 (N_21127,N_20117,N_20007);
nand U21128 (N_21128,N_20527,N_20299);
nor U21129 (N_21129,N_20591,N_20188);
and U21130 (N_21130,N_20170,N_20621);
or U21131 (N_21131,N_20209,N_20254);
and U21132 (N_21132,N_20276,N_20331);
and U21133 (N_21133,N_20246,N_20094);
nor U21134 (N_21134,N_20204,N_20197);
and U21135 (N_21135,N_20212,N_20603);
and U21136 (N_21136,N_20270,N_20136);
or U21137 (N_21137,N_20464,N_20578);
and U21138 (N_21138,N_20405,N_20610);
nand U21139 (N_21139,N_20128,N_20259);
or U21140 (N_21140,N_20529,N_20192);
or U21141 (N_21141,N_20087,N_20381);
or U21142 (N_21142,N_20375,N_20322);
xnor U21143 (N_21143,N_20242,N_20560);
and U21144 (N_21144,N_20597,N_20302);
nor U21145 (N_21145,N_20493,N_20562);
and U21146 (N_21146,N_20035,N_20516);
nand U21147 (N_21147,N_20132,N_20308);
and U21148 (N_21148,N_20551,N_20577);
or U21149 (N_21149,N_20130,N_20016);
nand U21150 (N_21150,N_20572,N_20316);
nand U21151 (N_21151,N_20167,N_20115);
and U21152 (N_21152,N_20026,N_20236);
or U21153 (N_21153,N_20379,N_20365);
or U21154 (N_21154,N_20497,N_20038);
or U21155 (N_21155,N_20347,N_20440);
or U21156 (N_21156,N_20486,N_20467);
or U21157 (N_21157,N_20575,N_20428);
nor U21158 (N_21158,N_20540,N_20616);
or U21159 (N_21159,N_20226,N_20001);
nand U21160 (N_21160,N_20042,N_20241);
and U21161 (N_21161,N_20140,N_20374);
xor U21162 (N_21162,N_20406,N_20148);
xor U21163 (N_21163,N_20170,N_20199);
nor U21164 (N_21164,N_20461,N_20499);
nand U21165 (N_21165,N_20558,N_20358);
nand U21166 (N_21166,N_20065,N_20011);
nand U21167 (N_21167,N_20446,N_20273);
and U21168 (N_21168,N_20485,N_20346);
and U21169 (N_21169,N_20044,N_20551);
xnor U21170 (N_21170,N_20219,N_20349);
or U21171 (N_21171,N_20617,N_20302);
and U21172 (N_21172,N_20618,N_20091);
nor U21173 (N_21173,N_20421,N_20059);
nand U21174 (N_21174,N_20343,N_20099);
and U21175 (N_21175,N_20548,N_20190);
xor U21176 (N_21176,N_20404,N_20327);
or U21177 (N_21177,N_20139,N_20563);
xor U21178 (N_21178,N_20542,N_20163);
nor U21179 (N_21179,N_20480,N_20001);
and U21180 (N_21180,N_20298,N_20495);
nor U21181 (N_21181,N_20413,N_20498);
nor U21182 (N_21182,N_20225,N_20426);
and U21183 (N_21183,N_20490,N_20123);
or U21184 (N_21184,N_20058,N_20404);
xnor U21185 (N_21185,N_20543,N_20495);
or U21186 (N_21186,N_20216,N_20042);
nor U21187 (N_21187,N_20578,N_20378);
xor U21188 (N_21188,N_20008,N_20442);
xor U21189 (N_21189,N_20201,N_20585);
or U21190 (N_21190,N_20525,N_20526);
and U21191 (N_21191,N_20414,N_20138);
nand U21192 (N_21192,N_20138,N_20584);
xnor U21193 (N_21193,N_20071,N_20300);
nand U21194 (N_21194,N_20458,N_20122);
xnor U21195 (N_21195,N_20208,N_20211);
xor U21196 (N_21196,N_20523,N_20155);
xnor U21197 (N_21197,N_20383,N_20288);
and U21198 (N_21198,N_20332,N_20178);
or U21199 (N_21199,N_20508,N_20519);
xnor U21200 (N_21200,N_20621,N_20252);
nor U21201 (N_21201,N_20541,N_20016);
and U21202 (N_21202,N_20093,N_20465);
nand U21203 (N_21203,N_20380,N_20247);
and U21204 (N_21204,N_20469,N_20039);
and U21205 (N_21205,N_20535,N_20207);
or U21206 (N_21206,N_20513,N_20227);
or U21207 (N_21207,N_20296,N_20606);
or U21208 (N_21208,N_20339,N_20130);
nor U21209 (N_21209,N_20058,N_20244);
nand U21210 (N_21210,N_20381,N_20175);
xnor U21211 (N_21211,N_20000,N_20282);
nand U21212 (N_21212,N_20416,N_20240);
or U21213 (N_21213,N_20607,N_20499);
nand U21214 (N_21214,N_20299,N_20597);
and U21215 (N_21215,N_20356,N_20129);
or U21216 (N_21216,N_20300,N_20329);
and U21217 (N_21217,N_20293,N_20128);
or U21218 (N_21218,N_20127,N_20196);
and U21219 (N_21219,N_20535,N_20146);
nor U21220 (N_21220,N_20330,N_20056);
nor U21221 (N_21221,N_20071,N_20055);
nand U21222 (N_21222,N_20205,N_20018);
or U21223 (N_21223,N_20590,N_20475);
nand U21224 (N_21224,N_20191,N_20398);
xor U21225 (N_21225,N_20238,N_20407);
and U21226 (N_21226,N_20541,N_20161);
xor U21227 (N_21227,N_20196,N_20177);
nor U21228 (N_21228,N_20180,N_20146);
nand U21229 (N_21229,N_20386,N_20230);
or U21230 (N_21230,N_20015,N_20524);
nor U21231 (N_21231,N_20473,N_20274);
nand U21232 (N_21232,N_20269,N_20000);
and U21233 (N_21233,N_20545,N_20591);
and U21234 (N_21234,N_20576,N_20149);
and U21235 (N_21235,N_20306,N_20097);
and U21236 (N_21236,N_20554,N_20279);
or U21237 (N_21237,N_20288,N_20036);
nand U21238 (N_21238,N_20568,N_20375);
and U21239 (N_21239,N_20587,N_20134);
nor U21240 (N_21240,N_20497,N_20506);
nand U21241 (N_21241,N_20516,N_20488);
xor U21242 (N_21242,N_20424,N_20399);
xor U21243 (N_21243,N_20512,N_20388);
xnor U21244 (N_21244,N_20031,N_20068);
xor U21245 (N_21245,N_20575,N_20071);
nand U21246 (N_21246,N_20107,N_20073);
and U21247 (N_21247,N_20461,N_20005);
or U21248 (N_21248,N_20264,N_20143);
nor U21249 (N_21249,N_20168,N_20299);
xnor U21250 (N_21250,N_21247,N_20954);
nand U21251 (N_21251,N_21156,N_20726);
nor U21252 (N_21252,N_21226,N_21071);
and U21253 (N_21253,N_21130,N_20710);
nand U21254 (N_21254,N_20955,N_20816);
nand U21255 (N_21255,N_20930,N_20885);
xnor U21256 (N_21256,N_21013,N_20774);
nor U21257 (N_21257,N_20731,N_20905);
and U21258 (N_21258,N_21181,N_20682);
and U21259 (N_21259,N_20755,N_20922);
nand U21260 (N_21260,N_20677,N_21033);
nand U21261 (N_21261,N_20762,N_21102);
xnor U21262 (N_21262,N_20758,N_20879);
xor U21263 (N_21263,N_21145,N_20988);
xor U21264 (N_21264,N_21056,N_20993);
or U21265 (N_21265,N_20749,N_20883);
or U21266 (N_21266,N_21179,N_20994);
and U21267 (N_21267,N_21195,N_20901);
and U21268 (N_21268,N_20788,N_20940);
nand U21269 (N_21269,N_20839,N_20824);
or U21270 (N_21270,N_21212,N_20983);
or U21271 (N_21271,N_20925,N_21141);
xor U21272 (N_21272,N_20972,N_21155);
nor U21273 (N_21273,N_21027,N_21018);
nand U21274 (N_21274,N_21135,N_20754);
and U21275 (N_21275,N_21140,N_20760);
and U21276 (N_21276,N_20927,N_20709);
nor U21277 (N_21277,N_20753,N_20951);
and U21278 (N_21278,N_20893,N_20923);
nand U21279 (N_21279,N_20696,N_20913);
nor U21280 (N_21280,N_21229,N_20832);
and U21281 (N_21281,N_21113,N_20803);
xor U21282 (N_21282,N_20685,N_21123);
or U21283 (N_21283,N_20843,N_20996);
nor U21284 (N_21284,N_20911,N_21088);
and U21285 (N_21285,N_21103,N_21132);
nor U21286 (N_21286,N_20667,N_21021);
or U21287 (N_21287,N_21170,N_21144);
or U21288 (N_21288,N_20875,N_20739);
xnor U21289 (N_21289,N_20786,N_20705);
or U21290 (N_21290,N_21243,N_20987);
nor U21291 (N_21291,N_20949,N_21126);
and U21292 (N_21292,N_20699,N_21238);
nand U21293 (N_21293,N_21178,N_20656);
nand U21294 (N_21294,N_20633,N_21177);
nand U21295 (N_21295,N_20694,N_21043);
nand U21296 (N_21296,N_21205,N_21202);
and U21297 (N_21297,N_21017,N_21114);
xor U21298 (N_21298,N_20907,N_21218);
xnor U21299 (N_21299,N_21194,N_20895);
xnor U21300 (N_21300,N_21072,N_20966);
nor U21301 (N_21301,N_20738,N_21068);
nand U21302 (N_21302,N_20891,N_21041);
xor U21303 (N_21303,N_21190,N_21036);
or U21304 (N_21304,N_21139,N_20759);
nor U21305 (N_21305,N_20757,N_20833);
nor U21306 (N_21306,N_21066,N_20952);
xor U21307 (N_21307,N_20890,N_20971);
nor U21308 (N_21308,N_21084,N_20747);
and U21309 (N_21309,N_20920,N_20926);
and U21310 (N_21310,N_20687,N_20770);
nor U21311 (N_21311,N_21022,N_21082);
xnor U21312 (N_21312,N_20767,N_20733);
nand U21313 (N_21313,N_20830,N_21023);
and U21314 (N_21314,N_21024,N_20887);
nand U21315 (N_21315,N_21115,N_21221);
and U21316 (N_21316,N_20918,N_21173);
or U21317 (N_21317,N_21049,N_21001);
and U21318 (N_21318,N_20724,N_20714);
xor U21319 (N_21319,N_21137,N_20836);
nand U21320 (N_21320,N_21215,N_20855);
or U21321 (N_21321,N_20676,N_21175);
nor U21322 (N_21322,N_20669,N_20625);
nand U21323 (N_21323,N_20878,N_21153);
or U21324 (N_21324,N_20799,N_21046);
xor U21325 (N_21325,N_21246,N_21163);
nor U21326 (N_21326,N_20736,N_20931);
and U21327 (N_21327,N_20730,N_21164);
nand U21328 (N_21328,N_21160,N_21138);
nand U21329 (N_21329,N_21191,N_21133);
nand U21330 (N_21330,N_21209,N_21165);
xnor U21331 (N_21331,N_20784,N_20691);
or U21332 (N_21332,N_20686,N_20640);
nand U21333 (N_21333,N_20795,N_21239);
and U21334 (N_21334,N_20702,N_21098);
nand U21335 (N_21335,N_20668,N_20792);
nand U21336 (N_21336,N_20825,N_21147);
or U21337 (N_21337,N_21070,N_20664);
and U21338 (N_21338,N_21000,N_20741);
or U21339 (N_21339,N_21249,N_21110);
or U21340 (N_21340,N_21047,N_20791);
and U21341 (N_21341,N_20756,N_20700);
or U21342 (N_21342,N_21231,N_20628);
nor U21343 (N_21343,N_20787,N_20977);
or U21344 (N_21344,N_20959,N_20750);
or U21345 (N_21345,N_21008,N_21146);
nand U21346 (N_21346,N_20894,N_20796);
or U21347 (N_21347,N_20998,N_20995);
and U21348 (N_21348,N_20812,N_20841);
nand U21349 (N_21349,N_20805,N_21025);
nor U21350 (N_21350,N_21196,N_20650);
nand U21351 (N_21351,N_21242,N_20642);
and U21352 (N_21352,N_21158,N_21223);
and U21353 (N_21353,N_21211,N_20829);
or U21354 (N_21354,N_20858,N_20910);
and U21355 (N_21355,N_20847,N_21093);
nor U21356 (N_21356,N_21125,N_21096);
nor U21357 (N_21357,N_21198,N_21105);
nand U21358 (N_21358,N_21055,N_21100);
xnor U21359 (N_21359,N_20933,N_20647);
and U21360 (N_21360,N_21121,N_21213);
nor U21361 (N_21361,N_21180,N_21142);
nand U21362 (N_21362,N_20678,N_20672);
or U21363 (N_21363,N_20725,N_21219);
nand U21364 (N_21364,N_20789,N_21091);
nor U21365 (N_21365,N_20990,N_20641);
xor U21366 (N_21366,N_21089,N_20899);
or U21367 (N_21367,N_20688,N_20826);
and U21368 (N_21368,N_21015,N_21062);
nand U21369 (N_21369,N_21232,N_21035);
nor U21370 (N_21370,N_21080,N_21048);
nor U21371 (N_21371,N_20752,N_20742);
and U21372 (N_21372,N_20908,N_20643);
and U21373 (N_21373,N_20635,N_20869);
xor U21374 (N_21374,N_20857,N_21065);
xnor U21375 (N_21375,N_20729,N_20882);
and U21376 (N_21376,N_20771,N_20960);
xor U21377 (N_21377,N_21006,N_20800);
nor U21378 (N_21378,N_20673,N_21183);
nand U21379 (N_21379,N_20946,N_20976);
nor U21380 (N_21380,N_20802,N_20835);
and U21381 (N_21381,N_21028,N_20906);
and U21382 (N_21382,N_21012,N_20680);
nand U21383 (N_21383,N_20775,N_20853);
nand U21384 (N_21384,N_20856,N_20982);
nor U21385 (N_21385,N_20860,N_20768);
and U21386 (N_21386,N_20881,N_21152);
xor U21387 (N_21387,N_20706,N_20684);
nor U21388 (N_21388,N_21003,N_20765);
xor U21389 (N_21389,N_21077,N_21154);
or U21390 (N_21390,N_20904,N_20840);
or U21391 (N_21391,N_20962,N_20711);
nand U21392 (N_21392,N_20675,N_20663);
xnor U21393 (N_21393,N_21007,N_20645);
xor U21394 (N_21394,N_20921,N_20766);
nand U21395 (N_21395,N_20790,N_21029);
nand U21396 (N_21396,N_20928,N_20867);
nor U21397 (N_21397,N_20704,N_21044);
xnor U21398 (N_21398,N_21095,N_20896);
and U21399 (N_21399,N_20818,N_20713);
nor U21400 (N_21400,N_20773,N_20877);
or U21401 (N_21401,N_21186,N_20892);
xnor U21402 (N_21402,N_20834,N_20880);
nand U21403 (N_21403,N_20813,N_21083);
xor U21404 (N_21404,N_20671,N_20652);
and U21405 (N_21405,N_20968,N_21149);
xnor U21406 (N_21406,N_20937,N_21002);
or U21407 (N_21407,N_21014,N_21225);
and U21408 (N_21408,N_21118,N_20900);
nor U21409 (N_21409,N_20958,N_21107);
and U21410 (N_21410,N_20953,N_20973);
or U21411 (N_21411,N_21074,N_20897);
or U21412 (N_21412,N_21159,N_20718);
xor U21413 (N_21413,N_20924,N_20939);
xor U21414 (N_21414,N_20785,N_21216);
nand U21415 (N_21415,N_21109,N_20817);
and U21416 (N_21416,N_20657,N_20779);
xnor U21417 (N_21417,N_20842,N_20655);
or U21418 (N_21418,N_20876,N_20707);
and U21419 (N_21419,N_21051,N_20720);
and U21420 (N_21420,N_21004,N_21050);
nand U21421 (N_21421,N_20764,N_20734);
xor U21422 (N_21422,N_20638,N_20965);
nor U21423 (N_21423,N_20991,N_21143);
or U21424 (N_21424,N_20852,N_20751);
or U21425 (N_21425,N_20941,N_21234);
xor U21426 (N_21426,N_21157,N_21206);
or U21427 (N_21427,N_20884,N_21201);
xor U21428 (N_21428,N_20659,N_20658);
or U21429 (N_21429,N_21053,N_21168);
and U21430 (N_21430,N_21244,N_20740);
xor U21431 (N_21431,N_21111,N_21167);
and U21432 (N_21432,N_21151,N_20814);
or U21433 (N_21433,N_20679,N_20654);
xor U21434 (N_21434,N_21199,N_21161);
nand U21435 (N_21435,N_20851,N_21052);
nor U21436 (N_21436,N_20936,N_21075);
nor U21437 (N_21437,N_20902,N_20723);
xnor U21438 (N_21438,N_20984,N_20938);
xor U21439 (N_21439,N_21009,N_21131);
and U21440 (N_21440,N_20828,N_21124);
nand U21441 (N_21441,N_21045,N_21136);
nor U21442 (N_21442,N_20948,N_20735);
nand U21443 (N_21443,N_20985,N_21188);
nand U21444 (N_21444,N_21092,N_20708);
nand U21445 (N_21445,N_20661,N_20957);
nand U21446 (N_21446,N_20997,N_20863);
and U21447 (N_21447,N_20660,N_20689);
nor U21448 (N_21448,N_20912,N_20989);
or U21449 (N_21449,N_20978,N_21122);
nor U21450 (N_21450,N_20945,N_21038);
xor U21451 (N_21451,N_20870,N_20916);
xnor U21452 (N_21452,N_21054,N_20632);
xnor U21453 (N_21453,N_20794,N_21117);
and U21454 (N_21454,N_21040,N_20859);
nor U21455 (N_21455,N_20961,N_20728);
xor U21456 (N_21456,N_20820,N_21034);
and U21457 (N_21457,N_21187,N_20837);
xor U21458 (N_21458,N_21245,N_20819);
nor U21459 (N_21459,N_21197,N_21097);
nand U21460 (N_21460,N_20862,N_20744);
or U21461 (N_21461,N_20992,N_21174);
nor U21462 (N_21462,N_21019,N_20967);
nor U21463 (N_21463,N_20888,N_20810);
or U21464 (N_21464,N_21189,N_20665);
and U21465 (N_21465,N_20737,N_20980);
nand U21466 (N_21466,N_20701,N_21090);
nor U21467 (N_21467,N_21063,N_21222);
nor U21468 (N_21468,N_21060,N_21057);
and U21469 (N_21469,N_20919,N_20864);
xnor U21470 (N_21470,N_20934,N_20849);
xnor U21471 (N_21471,N_21094,N_21228);
nor U21472 (N_21472,N_21087,N_20981);
and U21473 (N_21473,N_20693,N_20637);
or U21474 (N_21474,N_20801,N_20772);
or U21475 (N_21475,N_20964,N_21217);
and U21476 (N_21476,N_20850,N_20627);
and U21477 (N_21477,N_21058,N_21227);
nand U21478 (N_21478,N_21020,N_20646);
or U21479 (N_21479,N_21108,N_21112);
nand U21480 (N_21480,N_20662,N_20806);
nor U21481 (N_21481,N_21059,N_21042);
and U21482 (N_21482,N_20963,N_20846);
nor U21483 (N_21483,N_20644,N_20903);
xnor U21484 (N_21484,N_20909,N_20807);
xor U21485 (N_21485,N_21203,N_20782);
or U21486 (N_21486,N_20712,N_21171);
and U21487 (N_21487,N_21106,N_20808);
xnor U21488 (N_21488,N_20769,N_21240);
or U21489 (N_21489,N_21182,N_20732);
xnor U21490 (N_21490,N_21204,N_21011);
or U21491 (N_21491,N_20865,N_20692);
and U21492 (N_21492,N_20631,N_21236);
xor U21493 (N_21493,N_20653,N_20975);
and U21494 (N_21494,N_20698,N_20681);
or U21495 (N_21495,N_20827,N_20874);
or U21496 (N_21496,N_21210,N_20861);
or U21497 (N_21497,N_21005,N_20886);
nor U21498 (N_21498,N_21129,N_21193);
and U21499 (N_21499,N_20649,N_20697);
or U21500 (N_21500,N_21185,N_20917);
nor U21501 (N_21501,N_20703,N_20974);
or U21502 (N_21502,N_20871,N_21026);
or U21503 (N_21503,N_21184,N_21166);
nand U21504 (N_21504,N_21016,N_20778);
or U21505 (N_21505,N_21099,N_21208);
or U21506 (N_21506,N_21176,N_20722);
and U21507 (N_21507,N_21120,N_20873);
or U21508 (N_21508,N_21030,N_20748);
nand U21509 (N_21509,N_21241,N_21039);
and U21510 (N_21510,N_20690,N_20781);
xnor U21511 (N_21511,N_20715,N_20761);
xor U21512 (N_21512,N_20636,N_20845);
and U21513 (N_21513,N_21127,N_20815);
and U21514 (N_21514,N_21073,N_21031);
xor U21515 (N_21515,N_20629,N_21230);
or U21516 (N_21516,N_20763,N_21069);
nor U21517 (N_21517,N_20651,N_20695);
or U21518 (N_21518,N_21128,N_21086);
nand U21519 (N_21519,N_20979,N_20804);
or U21520 (N_21520,N_20719,N_20746);
xnor U21521 (N_21521,N_20745,N_20969);
nor U21522 (N_21522,N_20943,N_21104);
nor U21523 (N_21523,N_20783,N_21169);
nand U21524 (N_21524,N_21248,N_20780);
and U21525 (N_21525,N_21150,N_20872);
nand U21526 (N_21526,N_20683,N_21233);
nand U21527 (N_21527,N_21220,N_20942);
nand U21528 (N_21528,N_21061,N_20914);
nor U21529 (N_21529,N_20797,N_20743);
or U21530 (N_21530,N_20727,N_20999);
nor U21531 (N_21531,N_20777,N_20868);
nor U21532 (N_21532,N_20986,N_21085);
or U21533 (N_21533,N_20666,N_21162);
or U21534 (N_21534,N_21037,N_20630);
or U21535 (N_21535,N_20634,N_20970);
or U21536 (N_21536,N_20674,N_20944);
and U21537 (N_21537,N_21101,N_21192);
nand U21538 (N_21538,N_20889,N_20776);
nand U21539 (N_21539,N_21067,N_21079);
nor U21540 (N_21540,N_20947,N_20848);
xnor U21541 (N_21541,N_20932,N_20956);
or U21542 (N_21542,N_20935,N_20626);
xnor U21543 (N_21543,N_20809,N_21207);
or U21544 (N_21544,N_21116,N_21076);
or U21545 (N_21545,N_20844,N_20798);
nor U21546 (N_21546,N_21078,N_20822);
nand U21547 (N_21547,N_21237,N_21148);
or U21548 (N_21548,N_21119,N_20823);
and U21549 (N_21549,N_20811,N_21134);
and U21550 (N_21550,N_20821,N_20639);
or U21551 (N_21551,N_20950,N_20670);
or U21552 (N_21552,N_20831,N_20854);
and U21553 (N_21553,N_21214,N_20721);
nor U21554 (N_21554,N_20793,N_21172);
nor U21555 (N_21555,N_21224,N_21032);
nor U21556 (N_21556,N_21200,N_20866);
or U21557 (N_21557,N_21010,N_20838);
nand U21558 (N_21558,N_20929,N_21235);
and U21559 (N_21559,N_20898,N_20915);
nor U21560 (N_21560,N_21081,N_20716);
nor U21561 (N_21561,N_20648,N_21064);
nor U21562 (N_21562,N_20717,N_20755);
and U21563 (N_21563,N_21173,N_20676);
nand U21564 (N_21564,N_20886,N_21098);
nor U21565 (N_21565,N_20702,N_21014);
xnor U21566 (N_21566,N_20738,N_21190);
nand U21567 (N_21567,N_21108,N_21132);
nand U21568 (N_21568,N_20794,N_20811);
xnor U21569 (N_21569,N_20652,N_21186);
nand U21570 (N_21570,N_20872,N_20719);
and U21571 (N_21571,N_21021,N_21043);
nand U21572 (N_21572,N_20948,N_20718);
nand U21573 (N_21573,N_20750,N_20834);
nor U21574 (N_21574,N_20759,N_21181);
xnor U21575 (N_21575,N_20885,N_20977);
and U21576 (N_21576,N_20695,N_20784);
nand U21577 (N_21577,N_20878,N_21243);
nand U21578 (N_21578,N_21114,N_21122);
nor U21579 (N_21579,N_21185,N_21125);
nand U21580 (N_21580,N_20681,N_21025);
nor U21581 (N_21581,N_20826,N_21032);
and U21582 (N_21582,N_20820,N_20757);
xnor U21583 (N_21583,N_21131,N_21189);
xor U21584 (N_21584,N_20956,N_20920);
xnor U21585 (N_21585,N_20783,N_20678);
or U21586 (N_21586,N_21034,N_20770);
or U21587 (N_21587,N_20993,N_20677);
or U21588 (N_21588,N_21148,N_20819);
and U21589 (N_21589,N_21166,N_21165);
or U21590 (N_21590,N_21045,N_20691);
nor U21591 (N_21591,N_20676,N_20703);
xnor U21592 (N_21592,N_20717,N_21145);
or U21593 (N_21593,N_20754,N_20924);
and U21594 (N_21594,N_20941,N_20750);
or U21595 (N_21595,N_20804,N_20851);
xnor U21596 (N_21596,N_21157,N_20746);
or U21597 (N_21597,N_20750,N_20830);
xnor U21598 (N_21598,N_20693,N_21028);
nand U21599 (N_21599,N_21084,N_21086);
xor U21600 (N_21600,N_20997,N_20757);
and U21601 (N_21601,N_21166,N_21123);
nor U21602 (N_21602,N_21111,N_20920);
nand U21603 (N_21603,N_20756,N_21094);
and U21604 (N_21604,N_20837,N_20631);
xor U21605 (N_21605,N_21120,N_21005);
or U21606 (N_21606,N_20830,N_20798);
nand U21607 (N_21607,N_20679,N_20824);
and U21608 (N_21608,N_20680,N_20856);
xnor U21609 (N_21609,N_20646,N_20742);
xor U21610 (N_21610,N_20992,N_21192);
and U21611 (N_21611,N_20844,N_21212);
and U21612 (N_21612,N_20997,N_20989);
or U21613 (N_21613,N_20873,N_20992);
or U21614 (N_21614,N_20821,N_20905);
and U21615 (N_21615,N_20696,N_21099);
and U21616 (N_21616,N_21182,N_20841);
nor U21617 (N_21617,N_20995,N_20658);
and U21618 (N_21618,N_21200,N_20753);
nor U21619 (N_21619,N_21148,N_20889);
nand U21620 (N_21620,N_20805,N_21069);
xnor U21621 (N_21621,N_21161,N_21110);
xor U21622 (N_21622,N_20858,N_20917);
and U21623 (N_21623,N_20833,N_21139);
nor U21624 (N_21624,N_20770,N_21135);
xnor U21625 (N_21625,N_20870,N_21054);
and U21626 (N_21626,N_21114,N_21041);
xor U21627 (N_21627,N_20771,N_20811);
xnor U21628 (N_21628,N_21082,N_20670);
or U21629 (N_21629,N_21210,N_20700);
nor U21630 (N_21630,N_20876,N_20696);
nor U21631 (N_21631,N_21145,N_21211);
xor U21632 (N_21632,N_20980,N_20779);
and U21633 (N_21633,N_20807,N_20908);
and U21634 (N_21634,N_20658,N_20830);
nand U21635 (N_21635,N_20832,N_20842);
nor U21636 (N_21636,N_20947,N_21229);
and U21637 (N_21637,N_20949,N_20976);
xor U21638 (N_21638,N_21026,N_21162);
or U21639 (N_21639,N_21213,N_20890);
xor U21640 (N_21640,N_20991,N_21019);
or U21641 (N_21641,N_21088,N_20789);
or U21642 (N_21642,N_21031,N_20737);
nand U21643 (N_21643,N_20749,N_21050);
and U21644 (N_21644,N_21188,N_20857);
or U21645 (N_21645,N_20801,N_20859);
and U21646 (N_21646,N_21109,N_20865);
or U21647 (N_21647,N_20921,N_21219);
or U21648 (N_21648,N_20880,N_21064);
xor U21649 (N_21649,N_21038,N_21111);
nor U21650 (N_21650,N_20762,N_21007);
nand U21651 (N_21651,N_20993,N_21109);
and U21652 (N_21652,N_20875,N_21058);
nor U21653 (N_21653,N_21008,N_20955);
and U21654 (N_21654,N_20801,N_20918);
nand U21655 (N_21655,N_21079,N_20995);
nand U21656 (N_21656,N_21207,N_21138);
or U21657 (N_21657,N_20918,N_20932);
nor U21658 (N_21658,N_20782,N_20632);
xor U21659 (N_21659,N_21009,N_21038);
xnor U21660 (N_21660,N_21124,N_21032);
nand U21661 (N_21661,N_20883,N_20934);
or U21662 (N_21662,N_21144,N_21067);
nand U21663 (N_21663,N_20670,N_21140);
nor U21664 (N_21664,N_20991,N_20937);
xnor U21665 (N_21665,N_21019,N_21095);
nor U21666 (N_21666,N_20899,N_20873);
nor U21667 (N_21667,N_20862,N_21194);
or U21668 (N_21668,N_21178,N_20767);
or U21669 (N_21669,N_21247,N_20744);
xnor U21670 (N_21670,N_20866,N_20824);
or U21671 (N_21671,N_21004,N_21167);
xor U21672 (N_21672,N_20823,N_21102);
nand U21673 (N_21673,N_21113,N_21104);
xnor U21674 (N_21674,N_21087,N_21092);
xor U21675 (N_21675,N_20745,N_20840);
nor U21676 (N_21676,N_21170,N_20821);
or U21677 (N_21677,N_20919,N_21040);
xnor U21678 (N_21678,N_21178,N_20776);
and U21679 (N_21679,N_20697,N_21144);
nor U21680 (N_21680,N_21083,N_20736);
and U21681 (N_21681,N_20930,N_20689);
nand U21682 (N_21682,N_21126,N_21095);
xor U21683 (N_21683,N_20943,N_20660);
nor U21684 (N_21684,N_21221,N_21198);
nand U21685 (N_21685,N_20941,N_20865);
and U21686 (N_21686,N_21156,N_20869);
nor U21687 (N_21687,N_20826,N_20814);
nand U21688 (N_21688,N_20693,N_20957);
nor U21689 (N_21689,N_21213,N_21147);
and U21690 (N_21690,N_20858,N_20655);
or U21691 (N_21691,N_21180,N_21193);
and U21692 (N_21692,N_21199,N_21208);
nand U21693 (N_21693,N_20837,N_20890);
or U21694 (N_21694,N_20908,N_21037);
and U21695 (N_21695,N_20831,N_20948);
xnor U21696 (N_21696,N_20890,N_20811);
and U21697 (N_21697,N_20727,N_21242);
and U21698 (N_21698,N_20851,N_20713);
nor U21699 (N_21699,N_21051,N_21173);
or U21700 (N_21700,N_20994,N_20888);
nor U21701 (N_21701,N_20812,N_20800);
or U21702 (N_21702,N_20951,N_21196);
nand U21703 (N_21703,N_20821,N_20865);
nand U21704 (N_21704,N_20823,N_21183);
nor U21705 (N_21705,N_20844,N_20968);
and U21706 (N_21706,N_20883,N_20810);
xnor U21707 (N_21707,N_20844,N_21047);
nor U21708 (N_21708,N_20868,N_20867);
or U21709 (N_21709,N_20795,N_20852);
xor U21710 (N_21710,N_20815,N_21054);
and U21711 (N_21711,N_21145,N_20944);
nand U21712 (N_21712,N_21055,N_20967);
nor U21713 (N_21713,N_20795,N_20905);
nand U21714 (N_21714,N_21011,N_20693);
nand U21715 (N_21715,N_20978,N_20939);
nand U21716 (N_21716,N_21029,N_20644);
or U21717 (N_21717,N_20979,N_20848);
xnor U21718 (N_21718,N_20851,N_20834);
and U21719 (N_21719,N_20839,N_20681);
and U21720 (N_21720,N_20734,N_20730);
xnor U21721 (N_21721,N_20876,N_20736);
nand U21722 (N_21722,N_20719,N_21149);
xnor U21723 (N_21723,N_21042,N_21194);
nor U21724 (N_21724,N_20775,N_20774);
nor U21725 (N_21725,N_21073,N_21050);
or U21726 (N_21726,N_21240,N_21098);
and U21727 (N_21727,N_20825,N_21240);
or U21728 (N_21728,N_20699,N_20763);
nor U21729 (N_21729,N_20640,N_21109);
xnor U21730 (N_21730,N_20803,N_21028);
xor U21731 (N_21731,N_20635,N_20866);
xor U21732 (N_21732,N_20906,N_20774);
and U21733 (N_21733,N_20884,N_20712);
or U21734 (N_21734,N_20940,N_20667);
xnor U21735 (N_21735,N_21240,N_20995);
and U21736 (N_21736,N_20626,N_21131);
and U21737 (N_21737,N_20625,N_21171);
and U21738 (N_21738,N_21132,N_20916);
and U21739 (N_21739,N_21117,N_20891);
nor U21740 (N_21740,N_20858,N_20809);
and U21741 (N_21741,N_21054,N_20991);
xnor U21742 (N_21742,N_20935,N_21107);
xor U21743 (N_21743,N_21226,N_21096);
or U21744 (N_21744,N_20936,N_20822);
and U21745 (N_21745,N_20940,N_21101);
and U21746 (N_21746,N_20819,N_20724);
nand U21747 (N_21747,N_21147,N_21124);
nand U21748 (N_21748,N_20977,N_21168);
nor U21749 (N_21749,N_21177,N_21108);
or U21750 (N_21750,N_21121,N_21187);
xor U21751 (N_21751,N_21085,N_20936);
xnor U21752 (N_21752,N_20869,N_20803);
nor U21753 (N_21753,N_20933,N_20884);
or U21754 (N_21754,N_21097,N_21249);
nor U21755 (N_21755,N_20799,N_20809);
and U21756 (N_21756,N_20902,N_20919);
or U21757 (N_21757,N_20963,N_20852);
nor U21758 (N_21758,N_21155,N_21056);
and U21759 (N_21759,N_20674,N_20899);
and U21760 (N_21760,N_21050,N_20928);
nor U21761 (N_21761,N_20691,N_20834);
xnor U21762 (N_21762,N_20630,N_21021);
nor U21763 (N_21763,N_20634,N_20699);
nand U21764 (N_21764,N_20850,N_21113);
nor U21765 (N_21765,N_21229,N_21232);
nand U21766 (N_21766,N_20993,N_20806);
nand U21767 (N_21767,N_20870,N_20676);
or U21768 (N_21768,N_21149,N_20722);
nor U21769 (N_21769,N_20667,N_20911);
and U21770 (N_21770,N_20849,N_20630);
or U21771 (N_21771,N_21237,N_20940);
nor U21772 (N_21772,N_20685,N_20811);
or U21773 (N_21773,N_21211,N_20995);
nand U21774 (N_21774,N_20655,N_21249);
nand U21775 (N_21775,N_20964,N_21130);
nand U21776 (N_21776,N_21210,N_20934);
or U21777 (N_21777,N_21222,N_20710);
nand U21778 (N_21778,N_20735,N_20808);
and U21779 (N_21779,N_20656,N_20827);
nor U21780 (N_21780,N_20744,N_20718);
nand U21781 (N_21781,N_21221,N_21232);
xor U21782 (N_21782,N_21238,N_20954);
nor U21783 (N_21783,N_21229,N_21209);
nor U21784 (N_21784,N_21046,N_20692);
nor U21785 (N_21785,N_20886,N_21087);
or U21786 (N_21786,N_21131,N_20679);
xor U21787 (N_21787,N_21054,N_20742);
nand U21788 (N_21788,N_20934,N_20791);
xnor U21789 (N_21789,N_20744,N_20960);
and U21790 (N_21790,N_21216,N_21131);
xnor U21791 (N_21791,N_20802,N_20924);
and U21792 (N_21792,N_20746,N_21234);
and U21793 (N_21793,N_20731,N_20642);
and U21794 (N_21794,N_20634,N_21236);
or U21795 (N_21795,N_21059,N_21221);
and U21796 (N_21796,N_21067,N_20774);
or U21797 (N_21797,N_21230,N_20885);
xor U21798 (N_21798,N_20766,N_21189);
nand U21799 (N_21799,N_21246,N_20668);
or U21800 (N_21800,N_21103,N_20895);
nand U21801 (N_21801,N_21215,N_21140);
nor U21802 (N_21802,N_21209,N_20862);
nand U21803 (N_21803,N_20820,N_20681);
xor U21804 (N_21804,N_20723,N_20929);
or U21805 (N_21805,N_20896,N_20906);
nor U21806 (N_21806,N_20974,N_20724);
and U21807 (N_21807,N_21082,N_20757);
nand U21808 (N_21808,N_20739,N_21064);
xor U21809 (N_21809,N_21240,N_21074);
and U21810 (N_21810,N_20656,N_20855);
and U21811 (N_21811,N_20711,N_20931);
and U21812 (N_21812,N_21007,N_20913);
and U21813 (N_21813,N_20717,N_21115);
and U21814 (N_21814,N_20975,N_21202);
and U21815 (N_21815,N_21227,N_20889);
or U21816 (N_21816,N_20636,N_20638);
or U21817 (N_21817,N_21140,N_20761);
nand U21818 (N_21818,N_20965,N_20733);
and U21819 (N_21819,N_20763,N_20795);
and U21820 (N_21820,N_21156,N_20628);
or U21821 (N_21821,N_20744,N_21004);
or U21822 (N_21822,N_21045,N_20791);
nor U21823 (N_21823,N_20839,N_21205);
nor U21824 (N_21824,N_21230,N_21062);
xor U21825 (N_21825,N_21196,N_21141);
or U21826 (N_21826,N_20826,N_20843);
nor U21827 (N_21827,N_21238,N_21224);
xor U21828 (N_21828,N_20939,N_21181);
nand U21829 (N_21829,N_21048,N_20676);
or U21830 (N_21830,N_20802,N_20659);
or U21831 (N_21831,N_20892,N_20991);
nand U21832 (N_21832,N_21082,N_20811);
nor U21833 (N_21833,N_21132,N_21019);
xnor U21834 (N_21834,N_20893,N_21151);
nor U21835 (N_21835,N_21077,N_20943);
or U21836 (N_21836,N_20848,N_20712);
nor U21837 (N_21837,N_20916,N_20928);
nand U21838 (N_21838,N_20938,N_21184);
nor U21839 (N_21839,N_21136,N_21239);
and U21840 (N_21840,N_21226,N_21036);
nand U21841 (N_21841,N_20644,N_20783);
nor U21842 (N_21842,N_20753,N_20625);
nor U21843 (N_21843,N_20646,N_20908);
xnor U21844 (N_21844,N_20707,N_21127);
nor U21845 (N_21845,N_20830,N_21194);
nor U21846 (N_21846,N_21090,N_20838);
nand U21847 (N_21847,N_20789,N_20972);
nand U21848 (N_21848,N_20744,N_20763);
or U21849 (N_21849,N_20870,N_20959);
nand U21850 (N_21850,N_20686,N_20695);
nor U21851 (N_21851,N_20753,N_21078);
xnor U21852 (N_21852,N_21140,N_20852);
xnor U21853 (N_21853,N_21101,N_20867);
xor U21854 (N_21854,N_20803,N_20684);
and U21855 (N_21855,N_20875,N_20745);
or U21856 (N_21856,N_21016,N_20871);
nor U21857 (N_21857,N_20780,N_20682);
xnor U21858 (N_21858,N_20786,N_21030);
and U21859 (N_21859,N_21004,N_21178);
nor U21860 (N_21860,N_21248,N_20885);
nor U21861 (N_21861,N_20872,N_20959);
or U21862 (N_21862,N_21193,N_21133);
or U21863 (N_21863,N_21028,N_21151);
or U21864 (N_21864,N_21189,N_20647);
nand U21865 (N_21865,N_21059,N_20777);
or U21866 (N_21866,N_20666,N_20658);
nand U21867 (N_21867,N_20683,N_20817);
nor U21868 (N_21868,N_21242,N_20646);
nand U21869 (N_21869,N_20962,N_20922);
nor U21870 (N_21870,N_21056,N_20643);
xnor U21871 (N_21871,N_20631,N_20636);
nor U21872 (N_21872,N_20841,N_20840);
nand U21873 (N_21873,N_20780,N_21140);
nor U21874 (N_21874,N_20670,N_21072);
and U21875 (N_21875,N_21370,N_21250);
or U21876 (N_21876,N_21850,N_21281);
and U21877 (N_21877,N_21414,N_21856);
or U21878 (N_21878,N_21742,N_21279);
or U21879 (N_21879,N_21805,N_21393);
nor U21880 (N_21880,N_21710,N_21777);
nand U21881 (N_21881,N_21322,N_21613);
xnor U21882 (N_21882,N_21369,N_21470);
nor U21883 (N_21883,N_21706,N_21722);
or U21884 (N_21884,N_21530,N_21565);
xor U21885 (N_21885,N_21260,N_21251);
xor U21886 (N_21886,N_21581,N_21809);
and U21887 (N_21887,N_21665,N_21394);
and U21888 (N_21888,N_21511,N_21346);
or U21889 (N_21889,N_21738,N_21509);
and U21890 (N_21890,N_21574,N_21390);
xnor U21891 (N_21891,N_21841,N_21256);
nand U21892 (N_21892,N_21852,N_21277);
and U21893 (N_21893,N_21282,N_21596);
or U21894 (N_21894,N_21529,N_21763);
nor U21895 (N_21895,N_21448,N_21564);
xnor U21896 (N_21896,N_21378,N_21863);
nand U21897 (N_21897,N_21424,N_21327);
or U21898 (N_21898,N_21680,N_21491);
xnor U21899 (N_21899,N_21816,N_21363);
or U21900 (N_21900,N_21822,N_21569);
xnor U21901 (N_21901,N_21542,N_21261);
nand U21902 (N_21902,N_21811,N_21645);
nand U21903 (N_21903,N_21606,N_21373);
nor U21904 (N_21904,N_21496,N_21791);
xor U21905 (N_21905,N_21867,N_21612);
or U21906 (N_21906,N_21718,N_21588);
and U21907 (N_21907,N_21824,N_21702);
nand U21908 (N_21908,N_21679,N_21636);
xnor U21909 (N_21909,N_21506,N_21800);
nor U21910 (N_21910,N_21633,N_21745);
and U21911 (N_21911,N_21481,N_21550);
xor U21912 (N_21912,N_21731,N_21519);
and U21913 (N_21913,N_21659,N_21726);
xor U21914 (N_21914,N_21453,N_21799);
nor U21915 (N_21915,N_21642,N_21770);
xor U21916 (N_21916,N_21761,N_21562);
xor U21917 (N_21917,N_21720,N_21405);
or U21918 (N_21918,N_21591,N_21328);
and U21919 (N_21919,N_21338,N_21313);
xor U21920 (N_21920,N_21255,N_21868);
nor U21921 (N_21921,N_21634,N_21427);
xor U21922 (N_21922,N_21828,N_21662);
nand U21923 (N_21923,N_21418,N_21434);
and U21924 (N_21924,N_21455,N_21814);
xor U21925 (N_21925,N_21392,N_21570);
nand U21926 (N_21926,N_21437,N_21553);
or U21927 (N_21927,N_21810,N_21347);
or U21928 (N_21928,N_21334,N_21275);
xnor U21929 (N_21929,N_21433,N_21641);
nand U21930 (N_21930,N_21689,N_21525);
xnor U21931 (N_21931,N_21579,N_21778);
nor U21932 (N_21932,N_21836,N_21302);
or U21933 (N_21933,N_21727,N_21771);
nor U21934 (N_21934,N_21602,N_21871);
and U21935 (N_21935,N_21486,N_21395);
or U21936 (N_21936,N_21295,N_21305);
xor U21937 (N_21937,N_21270,N_21324);
xor U21938 (N_21938,N_21575,N_21499);
xor U21939 (N_21939,N_21479,N_21608);
nor U21940 (N_21940,N_21790,N_21497);
nor U21941 (N_21941,N_21618,N_21473);
and U21942 (N_21942,N_21838,N_21829);
xnor U21943 (N_21943,N_21339,N_21510);
or U21944 (N_21944,N_21257,N_21406);
nand U21945 (N_21945,N_21476,N_21292);
nand U21946 (N_21946,N_21254,N_21263);
and U21947 (N_21947,N_21644,N_21701);
nand U21948 (N_21948,N_21580,N_21619);
and U21949 (N_21949,N_21600,N_21735);
xor U21950 (N_21950,N_21541,N_21443);
nand U21951 (N_21951,N_21458,N_21681);
xnor U21952 (N_21952,N_21269,N_21274);
and U21953 (N_21953,N_21772,N_21375);
nand U21954 (N_21954,N_21306,N_21310);
nor U21955 (N_21955,N_21435,N_21801);
nand U21956 (N_21956,N_21563,N_21287);
xnor U21957 (N_21957,N_21278,N_21697);
xnor U21958 (N_21958,N_21625,N_21721);
nand U21959 (N_21959,N_21851,N_21766);
or U21960 (N_21960,N_21316,N_21262);
nor U21961 (N_21961,N_21603,N_21452);
and U21962 (N_21962,N_21594,N_21555);
nand U21963 (N_21963,N_21299,N_21289);
or U21964 (N_21964,N_21559,N_21482);
nor U21965 (N_21965,N_21821,N_21337);
xor U21966 (N_21966,N_21258,N_21410);
and U21967 (N_21967,N_21860,N_21391);
xor U21968 (N_21968,N_21558,N_21380);
xnor U21969 (N_21969,N_21853,N_21350);
nand U21970 (N_21970,N_21540,N_21691);
or U21971 (N_21971,N_21671,N_21818);
nand U21972 (N_21972,N_21782,N_21806);
xnor U21973 (N_21973,N_21366,N_21690);
nand U21974 (N_21974,N_21524,N_21477);
nand U21975 (N_21975,N_21503,N_21781);
or U21976 (N_21976,N_21705,N_21340);
xnor U21977 (N_21977,N_21667,N_21537);
xor U21978 (N_21978,N_21409,N_21398);
nand U21979 (N_21979,N_21445,N_21272);
and U21980 (N_21980,N_21514,N_21372);
and U21981 (N_21981,N_21283,N_21688);
nor U21982 (N_21982,N_21500,N_21732);
xor U21983 (N_21983,N_21360,N_21535);
xor U21984 (N_21984,N_21756,N_21533);
nor U21985 (N_21985,N_21297,N_21724);
xor U21986 (N_21986,N_21451,N_21787);
nand U21987 (N_21987,N_21684,N_21478);
and U21988 (N_21988,N_21592,N_21630);
or U21989 (N_21989,N_21517,N_21743);
nand U21990 (N_21990,N_21831,N_21751);
or U21991 (N_21991,N_21813,N_21512);
xnor U21992 (N_21992,N_21827,N_21741);
nor U21993 (N_21993,N_21872,N_21259);
xor U21994 (N_21994,N_21774,N_21627);
and U21995 (N_21995,N_21330,N_21361);
nand U21996 (N_21996,N_21861,N_21769);
and U21997 (N_21997,N_21859,N_21609);
and U21998 (N_21998,N_21488,N_21593);
and U21999 (N_21999,N_21447,N_21354);
and U22000 (N_22000,N_21615,N_21583);
and U22001 (N_22001,N_21472,N_21423);
nand U22002 (N_22002,N_21802,N_21561);
nand U22003 (N_22003,N_21397,N_21586);
or U22004 (N_22004,N_21400,N_21857);
or U22005 (N_22005,N_21573,N_21536);
xnor U22006 (N_22006,N_21749,N_21773);
and U22007 (N_22007,N_21661,N_21331);
xor U22008 (N_22008,N_21344,N_21484);
and U22009 (N_22009,N_21711,N_21543);
or U22010 (N_22010,N_21325,N_21385);
xor U22011 (N_22011,N_21620,N_21683);
or U22012 (N_22012,N_21696,N_21371);
nand U22013 (N_22013,N_21528,N_21265);
nand U22014 (N_22014,N_21675,N_21812);
nand U22015 (N_22015,N_21704,N_21566);
or U22016 (N_22016,N_21567,N_21759);
or U22017 (N_22017,N_21318,N_21288);
xor U22018 (N_22018,N_21725,N_21584);
xnor U22019 (N_22019,N_21660,N_21539);
nor U22020 (N_22020,N_21438,N_21786);
nor U22021 (N_22021,N_21797,N_21329);
xor U22022 (N_22022,N_21505,N_21436);
and U22023 (N_22023,N_21804,N_21678);
and U22024 (N_22024,N_21572,N_21650);
and U22025 (N_22025,N_21357,N_21485);
or U22026 (N_22026,N_21538,N_21674);
nor U22027 (N_22027,N_21723,N_21396);
xor U22028 (N_22028,N_21489,N_21601);
xnor U22029 (N_22029,N_21446,N_21707);
nor U22030 (N_22030,N_21686,N_21595);
or U22031 (N_22031,N_21532,N_21468);
nor U22032 (N_22032,N_21654,N_21590);
nor U22033 (N_22033,N_21404,N_21833);
and U22034 (N_22034,N_21652,N_21382);
and U22035 (N_22035,N_21623,N_21783);
or U22036 (N_22036,N_21425,N_21639);
or U22037 (N_22037,N_21317,N_21271);
or U22038 (N_22038,N_21646,N_21296);
xnor U22039 (N_22039,N_21546,N_21744);
nor U22040 (N_22040,N_21311,N_21483);
nand U22041 (N_22041,N_21268,N_21611);
and U22042 (N_22042,N_21577,N_21507);
or U22043 (N_22043,N_21647,N_21466);
xnor U22044 (N_22044,N_21359,N_21864);
nor U22045 (N_22045,N_21381,N_21557);
and U22046 (N_22046,N_21531,N_21544);
nor U22047 (N_22047,N_21374,N_21475);
and U22048 (N_22048,N_21501,N_21849);
or U22049 (N_22049,N_21534,N_21668);
nor U22050 (N_22050,N_21342,N_21432);
nor U22051 (N_22051,N_21714,N_21321);
and U22052 (N_22052,N_21740,N_21556);
or U22053 (N_22053,N_21267,N_21846);
nor U22054 (N_22054,N_21610,N_21670);
nor U22055 (N_22055,N_21355,N_21709);
or U22056 (N_22056,N_21307,N_21315);
or U22057 (N_22057,N_21440,N_21869);
or U22058 (N_22058,N_21789,N_21746);
nand U22059 (N_22059,N_21762,N_21461);
nand U22060 (N_22060,N_21874,N_21430);
xnor U22061 (N_22061,N_21284,N_21765);
nand U22062 (N_22062,N_21730,N_21421);
or U22063 (N_22063,N_21651,N_21356);
xnor U22064 (N_22064,N_21401,N_21293);
xor U22065 (N_22065,N_21492,N_21304);
nor U22066 (N_22066,N_21280,N_21419);
nand U22067 (N_22067,N_21784,N_21653);
and U22068 (N_22068,N_21819,N_21700);
and U22069 (N_22069,N_21621,N_21326);
or U22070 (N_22070,N_21605,N_21676);
or U22071 (N_22071,N_21286,N_21333);
xnor U22072 (N_22072,N_21444,N_21808);
and U22073 (N_22073,N_21467,N_21303);
xnor U22074 (N_22074,N_21693,N_21719);
or U22075 (N_22075,N_21367,N_21456);
xor U22076 (N_22076,N_21637,N_21495);
and U22077 (N_22077,N_21522,N_21403);
xor U22078 (N_22078,N_21264,N_21545);
xor U22079 (N_22079,N_21753,N_21527);
xnor U22080 (N_22080,N_21757,N_21521);
nor U22081 (N_22081,N_21792,N_21413);
nand U22082 (N_22082,N_21798,N_21717);
nor U22083 (N_22083,N_21854,N_21399);
or U22084 (N_22084,N_21632,N_21752);
nor U22085 (N_22085,N_21578,N_21649);
nand U22086 (N_22086,N_21471,N_21796);
nor U22087 (N_22087,N_21490,N_21739);
or U22088 (N_22088,N_21560,N_21803);
nand U22089 (N_22089,N_21388,N_21695);
nand U22090 (N_22090,N_21823,N_21494);
or U22091 (N_22091,N_21515,N_21729);
and U22092 (N_22092,N_21873,N_21622);
nor U22093 (N_22093,N_21733,N_21767);
and U22094 (N_22094,N_21628,N_21300);
xnor U22095 (N_22095,N_21498,N_21576);
nor U22096 (N_22096,N_21460,N_21638);
xor U22097 (N_22097,N_21459,N_21582);
and U22098 (N_22098,N_21826,N_21308);
nor U22099 (N_22099,N_21734,N_21516);
nor U22100 (N_22100,N_21407,N_21585);
nand U22101 (N_22101,N_21715,N_21520);
xnor U22102 (N_22102,N_21648,N_21411);
nor U22103 (N_22103,N_21698,N_21677);
xnor U22104 (N_22104,N_21664,N_21748);
nor U22105 (N_22105,N_21387,N_21865);
xnor U22106 (N_22106,N_21487,N_21549);
and U22107 (N_22107,N_21314,N_21480);
or U22108 (N_22108,N_21508,N_21844);
xnor U22109 (N_22109,N_21847,N_21760);
nand U22110 (N_22110,N_21755,N_21252);
nor U22111 (N_22111,N_21685,N_21384);
nand U22112 (N_22112,N_21794,N_21513);
xor U22113 (N_22113,N_21817,N_21416);
nor U22114 (N_22114,N_21820,N_21417);
xnor U22115 (N_22115,N_21353,N_21750);
and U22116 (N_22116,N_21319,N_21554);
xnor U22117 (N_22117,N_21383,N_21640);
or U22118 (N_22118,N_21377,N_21571);
or U22119 (N_22119,N_21764,N_21736);
nor U22120 (N_22120,N_21699,N_21568);
or U22121 (N_22121,N_21441,N_21362);
and U22122 (N_22122,N_21643,N_21673);
or U22123 (N_22123,N_21835,N_21551);
nor U22124 (N_22124,N_21703,N_21358);
and U22125 (N_22125,N_21815,N_21426);
and U22126 (N_22126,N_21523,N_21341);
or U22127 (N_22127,N_21309,N_21348);
xor U22128 (N_22128,N_21450,N_21708);
or U22129 (N_22129,N_21758,N_21276);
nand U22130 (N_22130,N_21807,N_21842);
or U22131 (N_22131,N_21830,N_21442);
or U22132 (N_22132,N_21768,N_21607);
or U22133 (N_22133,N_21352,N_21692);
xnor U22134 (N_22134,N_21598,N_21320);
nor U22135 (N_22135,N_21457,N_21291);
xnor U22136 (N_22136,N_21465,N_21716);
or U22137 (N_22137,N_21825,N_21449);
and U22138 (N_22138,N_21845,N_21469);
nand U22139 (N_22139,N_21290,N_21389);
and U22140 (N_22140,N_21843,N_21834);
nand U22141 (N_22141,N_21379,N_21518);
nand U22142 (N_22142,N_21712,N_21428);
and U22143 (N_22143,N_21332,N_21655);
xnor U22144 (N_22144,N_21657,N_21408);
or U22145 (N_22145,N_21463,N_21866);
and U22146 (N_22146,N_21616,N_21728);
xor U22147 (N_22147,N_21604,N_21349);
xor U22148 (N_22148,N_21775,N_21669);
and U22149 (N_22149,N_21858,N_21345);
xnor U22150 (N_22150,N_21713,N_21412);
nor U22151 (N_22151,N_21780,N_21658);
nand U22152 (N_22152,N_21754,N_21832);
nand U22153 (N_22153,N_21364,N_21386);
or U22154 (N_22154,N_21454,N_21694);
or U22155 (N_22155,N_21656,N_21464);
nor U22156 (N_22156,N_21666,N_21376);
nand U22157 (N_22157,N_21599,N_21848);
nand U22158 (N_22158,N_21439,N_21793);
nand U22159 (N_22159,N_21429,N_21431);
and U22160 (N_22160,N_21624,N_21548);
and U22161 (N_22161,N_21855,N_21266);
nor U22162 (N_22162,N_21462,N_21420);
or U22163 (N_22163,N_21587,N_21335);
and U22164 (N_22164,N_21870,N_21502);
xnor U22165 (N_22165,N_21672,N_21617);
xnor U22166 (N_22166,N_21839,N_21422);
and U22167 (N_22167,N_21526,N_21629);
and U22168 (N_22168,N_21402,N_21597);
nor U22169 (N_22169,N_21312,N_21323);
nand U22170 (N_22170,N_21365,N_21415);
nand U22171 (N_22171,N_21474,N_21368);
xnor U22172 (N_22172,N_21253,N_21493);
and U22173 (N_22173,N_21837,N_21285);
nor U22174 (N_22174,N_21682,N_21547);
nand U22175 (N_22175,N_21343,N_21776);
or U22176 (N_22176,N_21301,N_21840);
xnor U22177 (N_22177,N_21663,N_21785);
xor U22178 (N_22178,N_21687,N_21294);
xnor U22179 (N_22179,N_21552,N_21298);
xor U22180 (N_22180,N_21351,N_21631);
and U22181 (N_22181,N_21273,N_21626);
or U22182 (N_22182,N_21737,N_21589);
nand U22183 (N_22183,N_21635,N_21862);
or U22184 (N_22184,N_21336,N_21779);
nor U22185 (N_22185,N_21795,N_21747);
nand U22186 (N_22186,N_21788,N_21614);
nand U22187 (N_22187,N_21504,N_21850);
nor U22188 (N_22188,N_21435,N_21571);
nor U22189 (N_22189,N_21523,N_21829);
nor U22190 (N_22190,N_21513,N_21770);
xor U22191 (N_22191,N_21847,N_21786);
nor U22192 (N_22192,N_21418,N_21834);
nor U22193 (N_22193,N_21815,N_21305);
nand U22194 (N_22194,N_21630,N_21781);
nand U22195 (N_22195,N_21256,N_21636);
nand U22196 (N_22196,N_21409,N_21712);
and U22197 (N_22197,N_21769,N_21541);
or U22198 (N_22198,N_21642,N_21740);
and U22199 (N_22199,N_21527,N_21260);
nor U22200 (N_22200,N_21307,N_21545);
xor U22201 (N_22201,N_21336,N_21477);
and U22202 (N_22202,N_21496,N_21844);
and U22203 (N_22203,N_21253,N_21530);
and U22204 (N_22204,N_21746,N_21660);
xnor U22205 (N_22205,N_21354,N_21782);
or U22206 (N_22206,N_21814,N_21303);
nor U22207 (N_22207,N_21595,N_21354);
xnor U22208 (N_22208,N_21742,N_21778);
and U22209 (N_22209,N_21526,N_21814);
nand U22210 (N_22210,N_21481,N_21867);
nor U22211 (N_22211,N_21771,N_21394);
and U22212 (N_22212,N_21329,N_21653);
nor U22213 (N_22213,N_21440,N_21667);
nand U22214 (N_22214,N_21347,N_21868);
and U22215 (N_22215,N_21486,N_21763);
xor U22216 (N_22216,N_21597,N_21327);
nand U22217 (N_22217,N_21322,N_21773);
or U22218 (N_22218,N_21865,N_21722);
nor U22219 (N_22219,N_21790,N_21493);
xnor U22220 (N_22220,N_21790,N_21486);
and U22221 (N_22221,N_21788,N_21777);
nor U22222 (N_22222,N_21353,N_21846);
nor U22223 (N_22223,N_21589,N_21587);
or U22224 (N_22224,N_21557,N_21265);
nand U22225 (N_22225,N_21541,N_21551);
xnor U22226 (N_22226,N_21371,N_21590);
nor U22227 (N_22227,N_21343,N_21752);
nor U22228 (N_22228,N_21532,N_21381);
and U22229 (N_22229,N_21537,N_21318);
xnor U22230 (N_22230,N_21314,N_21270);
and U22231 (N_22231,N_21727,N_21804);
nor U22232 (N_22232,N_21325,N_21654);
nand U22233 (N_22233,N_21873,N_21541);
and U22234 (N_22234,N_21486,N_21605);
and U22235 (N_22235,N_21368,N_21250);
and U22236 (N_22236,N_21266,N_21451);
nor U22237 (N_22237,N_21793,N_21588);
or U22238 (N_22238,N_21507,N_21665);
nor U22239 (N_22239,N_21774,N_21753);
nand U22240 (N_22240,N_21731,N_21280);
nor U22241 (N_22241,N_21309,N_21743);
or U22242 (N_22242,N_21864,N_21844);
nor U22243 (N_22243,N_21594,N_21536);
nand U22244 (N_22244,N_21263,N_21703);
or U22245 (N_22245,N_21362,N_21437);
and U22246 (N_22246,N_21507,N_21336);
xor U22247 (N_22247,N_21790,N_21647);
or U22248 (N_22248,N_21750,N_21557);
nor U22249 (N_22249,N_21655,N_21321);
xnor U22250 (N_22250,N_21404,N_21665);
nand U22251 (N_22251,N_21624,N_21523);
or U22252 (N_22252,N_21451,N_21835);
xnor U22253 (N_22253,N_21426,N_21868);
nand U22254 (N_22254,N_21283,N_21479);
nand U22255 (N_22255,N_21623,N_21565);
or U22256 (N_22256,N_21730,N_21850);
nor U22257 (N_22257,N_21360,N_21659);
or U22258 (N_22258,N_21646,N_21391);
nor U22259 (N_22259,N_21574,N_21276);
or U22260 (N_22260,N_21310,N_21398);
xnor U22261 (N_22261,N_21755,N_21375);
and U22262 (N_22262,N_21722,N_21287);
or U22263 (N_22263,N_21806,N_21421);
nor U22264 (N_22264,N_21474,N_21779);
xor U22265 (N_22265,N_21365,N_21588);
and U22266 (N_22266,N_21518,N_21686);
nand U22267 (N_22267,N_21588,N_21314);
and U22268 (N_22268,N_21539,N_21394);
and U22269 (N_22269,N_21507,N_21312);
xor U22270 (N_22270,N_21829,N_21340);
nand U22271 (N_22271,N_21260,N_21662);
xnor U22272 (N_22272,N_21618,N_21320);
nand U22273 (N_22273,N_21351,N_21839);
and U22274 (N_22274,N_21415,N_21622);
or U22275 (N_22275,N_21518,N_21418);
and U22276 (N_22276,N_21266,N_21453);
nand U22277 (N_22277,N_21852,N_21671);
nor U22278 (N_22278,N_21765,N_21366);
xnor U22279 (N_22279,N_21366,N_21650);
xnor U22280 (N_22280,N_21848,N_21590);
nand U22281 (N_22281,N_21444,N_21686);
or U22282 (N_22282,N_21676,N_21407);
nor U22283 (N_22283,N_21301,N_21859);
nand U22284 (N_22284,N_21633,N_21429);
nand U22285 (N_22285,N_21713,N_21744);
or U22286 (N_22286,N_21372,N_21473);
or U22287 (N_22287,N_21672,N_21527);
and U22288 (N_22288,N_21631,N_21654);
and U22289 (N_22289,N_21291,N_21777);
or U22290 (N_22290,N_21571,N_21448);
or U22291 (N_22291,N_21591,N_21741);
and U22292 (N_22292,N_21424,N_21838);
nor U22293 (N_22293,N_21496,N_21869);
and U22294 (N_22294,N_21582,N_21299);
xnor U22295 (N_22295,N_21776,N_21642);
xnor U22296 (N_22296,N_21839,N_21535);
nor U22297 (N_22297,N_21669,N_21370);
xor U22298 (N_22298,N_21546,N_21463);
and U22299 (N_22299,N_21797,N_21792);
or U22300 (N_22300,N_21811,N_21747);
nor U22301 (N_22301,N_21506,N_21736);
nand U22302 (N_22302,N_21293,N_21642);
and U22303 (N_22303,N_21623,N_21779);
and U22304 (N_22304,N_21550,N_21463);
or U22305 (N_22305,N_21463,N_21632);
xor U22306 (N_22306,N_21681,N_21723);
nor U22307 (N_22307,N_21542,N_21434);
nand U22308 (N_22308,N_21785,N_21399);
or U22309 (N_22309,N_21503,N_21838);
xnor U22310 (N_22310,N_21484,N_21797);
xnor U22311 (N_22311,N_21456,N_21348);
xor U22312 (N_22312,N_21761,N_21665);
and U22313 (N_22313,N_21825,N_21672);
and U22314 (N_22314,N_21758,N_21639);
or U22315 (N_22315,N_21828,N_21707);
nor U22316 (N_22316,N_21671,N_21706);
or U22317 (N_22317,N_21796,N_21287);
nand U22318 (N_22318,N_21375,N_21823);
and U22319 (N_22319,N_21688,N_21620);
or U22320 (N_22320,N_21251,N_21751);
or U22321 (N_22321,N_21573,N_21257);
xor U22322 (N_22322,N_21792,N_21845);
xor U22323 (N_22323,N_21589,N_21486);
nor U22324 (N_22324,N_21606,N_21280);
or U22325 (N_22325,N_21724,N_21417);
and U22326 (N_22326,N_21647,N_21343);
xor U22327 (N_22327,N_21541,N_21398);
or U22328 (N_22328,N_21605,N_21737);
nand U22329 (N_22329,N_21333,N_21812);
and U22330 (N_22330,N_21868,N_21525);
xnor U22331 (N_22331,N_21268,N_21683);
or U22332 (N_22332,N_21735,N_21704);
nor U22333 (N_22333,N_21703,N_21825);
nor U22334 (N_22334,N_21604,N_21471);
nand U22335 (N_22335,N_21632,N_21261);
or U22336 (N_22336,N_21509,N_21442);
nor U22337 (N_22337,N_21495,N_21822);
xor U22338 (N_22338,N_21405,N_21672);
xor U22339 (N_22339,N_21833,N_21499);
or U22340 (N_22340,N_21621,N_21568);
xor U22341 (N_22341,N_21737,N_21590);
xor U22342 (N_22342,N_21270,N_21415);
nor U22343 (N_22343,N_21251,N_21450);
nor U22344 (N_22344,N_21400,N_21703);
xor U22345 (N_22345,N_21369,N_21726);
or U22346 (N_22346,N_21257,N_21502);
or U22347 (N_22347,N_21470,N_21393);
nand U22348 (N_22348,N_21672,N_21492);
nor U22349 (N_22349,N_21624,N_21440);
nand U22350 (N_22350,N_21855,N_21600);
and U22351 (N_22351,N_21359,N_21552);
xnor U22352 (N_22352,N_21663,N_21866);
nand U22353 (N_22353,N_21858,N_21660);
nor U22354 (N_22354,N_21389,N_21713);
xnor U22355 (N_22355,N_21254,N_21859);
and U22356 (N_22356,N_21700,N_21657);
nor U22357 (N_22357,N_21274,N_21735);
nand U22358 (N_22358,N_21773,N_21380);
and U22359 (N_22359,N_21526,N_21264);
xnor U22360 (N_22360,N_21582,N_21291);
nor U22361 (N_22361,N_21813,N_21778);
nor U22362 (N_22362,N_21841,N_21815);
xor U22363 (N_22363,N_21286,N_21785);
and U22364 (N_22364,N_21424,N_21730);
or U22365 (N_22365,N_21538,N_21629);
nand U22366 (N_22366,N_21426,N_21712);
or U22367 (N_22367,N_21643,N_21813);
nor U22368 (N_22368,N_21555,N_21279);
nor U22369 (N_22369,N_21536,N_21292);
xnor U22370 (N_22370,N_21754,N_21409);
and U22371 (N_22371,N_21870,N_21858);
nor U22372 (N_22372,N_21743,N_21820);
or U22373 (N_22373,N_21611,N_21729);
nand U22374 (N_22374,N_21501,N_21300);
xnor U22375 (N_22375,N_21867,N_21694);
nor U22376 (N_22376,N_21488,N_21604);
or U22377 (N_22377,N_21568,N_21516);
xor U22378 (N_22378,N_21354,N_21312);
or U22379 (N_22379,N_21856,N_21618);
and U22380 (N_22380,N_21465,N_21680);
nor U22381 (N_22381,N_21805,N_21614);
xnor U22382 (N_22382,N_21801,N_21353);
nand U22383 (N_22383,N_21736,N_21781);
and U22384 (N_22384,N_21865,N_21797);
and U22385 (N_22385,N_21516,N_21253);
and U22386 (N_22386,N_21749,N_21780);
and U22387 (N_22387,N_21623,N_21616);
nand U22388 (N_22388,N_21302,N_21324);
or U22389 (N_22389,N_21363,N_21859);
nand U22390 (N_22390,N_21356,N_21565);
nor U22391 (N_22391,N_21490,N_21492);
nor U22392 (N_22392,N_21524,N_21323);
xor U22393 (N_22393,N_21631,N_21713);
or U22394 (N_22394,N_21388,N_21591);
nor U22395 (N_22395,N_21440,N_21832);
nand U22396 (N_22396,N_21833,N_21800);
xor U22397 (N_22397,N_21287,N_21828);
or U22398 (N_22398,N_21348,N_21630);
xor U22399 (N_22399,N_21489,N_21323);
nand U22400 (N_22400,N_21835,N_21250);
nand U22401 (N_22401,N_21812,N_21606);
and U22402 (N_22402,N_21397,N_21796);
nor U22403 (N_22403,N_21543,N_21847);
and U22404 (N_22404,N_21607,N_21433);
or U22405 (N_22405,N_21871,N_21646);
or U22406 (N_22406,N_21863,N_21812);
nand U22407 (N_22407,N_21658,N_21624);
nor U22408 (N_22408,N_21344,N_21654);
xnor U22409 (N_22409,N_21705,N_21509);
nor U22410 (N_22410,N_21356,N_21566);
or U22411 (N_22411,N_21754,N_21672);
and U22412 (N_22412,N_21333,N_21577);
nand U22413 (N_22413,N_21370,N_21597);
nand U22414 (N_22414,N_21266,N_21571);
nor U22415 (N_22415,N_21465,N_21617);
xnor U22416 (N_22416,N_21726,N_21622);
or U22417 (N_22417,N_21668,N_21360);
or U22418 (N_22418,N_21855,N_21486);
or U22419 (N_22419,N_21509,N_21359);
nand U22420 (N_22420,N_21673,N_21623);
or U22421 (N_22421,N_21434,N_21255);
and U22422 (N_22422,N_21678,N_21542);
nor U22423 (N_22423,N_21250,N_21673);
xnor U22424 (N_22424,N_21291,N_21528);
and U22425 (N_22425,N_21258,N_21484);
and U22426 (N_22426,N_21560,N_21323);
and U22427 (N_22427,N_21258,N_21308);
and U22428 (N_22428,N_21340,N_21383);
xor U22429 (N_22429,N_21739,N_21640);
and U22430 (N_22430,N_21409,N_21617);
and U22431 (N_22431,N_21661,N_21690);
or U22432 (N_22432,N_21740,N_21870);
and U22433 (N_22433,N_21439,N_21473);
nor U22434 (N_22434,N_21513,N_21674);
and U22435 (N_22435,N_21412,N_21646);
nor U22436 (N_22436,N_21868,N_21745);
xor U22437 (N_22437,N_21535,N_21388);
xor U22438 (N_22438,N_21759,N_21766);
nor U22439 (N_22439,N_21468,N_21418);
nand U22440 (N_22440,N_21440,N_21332);
xnor U22441 (N_22441,N_21472,N_21536);
nand U22442 (N_22442,N_21766,N_21349);
xor U22443 (N_22443,N_21381,N_21771);
or U22444 (N_22444,N_21316,N_21655);
xor U22445 (N_22445,N_21407,N_21251);
nand U22446 (N_22446,N_21263,N_21710);
and U22447 (N_22447,N_21447,N_21802);
xnor U22448 (N_22448,N_21614,N_21505);
nor U22449 (N_22449,N_21695,N_21283);
xor U22450 (N_22450,N_21832,N_21554);
xnor U22451 (N_22451,N_21480,N_21798);
nand U22452 (N_22452,N_21360,N_21635);
or U22453 (N_22453,N_21577,N_21511);
nand U22454 (N_22454,N_21807,N_21821);
or U22455 (N_22455,N_21650,N_21740);
or U22456 (N_22456,N_21499,N_21517);
nand U22457 (N_22457,N_21615,N_21430);
nand U22458 (N_22458,N_21744,N_21561);
and U22459 (N_22459,N_21525,N_21497);
or U22460 (N_22460,N_21561,N_21752);
xnor U22461 (N_22461,N_21258,N_21294);
or U22462 (N_22462,N_21740,N_21281);
and U22463 (N_22463,N_21404,N_21666);
nor U22464 (N_22464,N_21707,N_21520);
nand U22465 (N_22465,N_21288,N_21442);
and U22466 (N_22466,N_21757,N_21544);
nand U22467 (N_22467,N_21501,N_21523);
nand U22468 (N_22468,N_21693,N_21520);
or U22469 (N_22469,N_21866,N_21459);
xnor U22470 (N_22470,N_21491,N_21422);
and U22471 (N_22471,N_21812,N_21345);
nor U22472 (N_22472,N_21552,N_21806);
nor U22473 (N_22473,N_21526,N_21622);
and U22474 (N_22474,N_21420,N_21623);
nand U22475 (N_22475,N_21368,N_21812);
or U22476 (N_22476,N_21772,N_21782);
nand U22477 (N_22477,N_21686,N_21616);
xnor U22478 (N_22478,N_21596,N_21313);
xnor U22479 (N_22479,N_21676,N_21626);
or U22480 (N_22480,N_21558,N_21306);
nand U22481 (N_22481,N_21710,N_21332);
nor U22482 (N_22482,N_21398,N_21278);
nand U22483 (N_22483,N_21282,N_21663);
or U22484 (N_22484,N_21289,N_21652);
nand U22485 (N_22485,N_21282,N_21723);
nor U22486 (N_22486,N_21706,N_21589);
xnor U22487 (N_22487,N_21548,N_21347);
or U22488 (N_22488,N_21661,N_21515);
or U22489 (N_22489,N_21685,N_21533);
and U22490 (N_22490,N_21786,N_21465);
nand U22491 (N_22491,N_21530,N_21729);
nand U22492 (N_22492,N_21864,N_21603);
and U22493 (N_22493,N_21640,N_21699);
and U22494 (N_22494,N_21458,N_21300);
or U22495 (N_22495,N_21866,N_21597);
nand U22496 (N_22496,N_21658,N_21832);
nor U22497 (N_22497,N_21299,N_21710);
and U22498 (N_22498,N_21583,N_21619);
and U22499 (N_22499,N_21648,N_21563);
xnor U22500 (N_22500,N_22384,N_22075);
xnor U22501 (N_22501,N_21964,N_22452);
or U22502 (N_22502,N_22252,N_22122);
nor U22503 (N_22503,N_22158,N_22131);
nand U22504 (N_22504,N_22145,N_22410);
or U22505 (N_22505,N_21917,N_22454);
nor U22506 (N_22506,N_22062,N_21912);
and U22507 (N_22507,N_21987,N_22343);
nor U22508 (N_22508,N_22306,N_21908);
nor U22509 (N_22509,N_22060,N_22048);
nand U22510 (N_22510,N_22399,N_21875);
xor U22511 (N_22511,N_22245,N_22271);
or U22512 (N_22512,N_21993,N_22157);
or U22513 (N_22513,N_22416,N_21907);
xor U22514 (N_22514,N_21977,N_21920);
nand U22515 (N_22515,N_22007,N_22202);
or U22516 (N_22516,N_22216,N_22173);
and U22517 (N_22517,N_22152,N_22228);
and U22518 (N_22518,N_22290,N_21927);
nand U22519 (N_22519,N_21923,N_22334);
and U22520 (N_22520,N_22016,N_22379);
and U22521 (N_22521,N_22256,N_22344);
xor U22522 (N_22522,N_22451,N_21929);
or U22523 (N_22523,N_22365,N_21959);
xnor U22524 (N_22524,N_22025,N_22052);
nand U22525 (N_22525,N_21913,N_22413);
xor U22526 (N_22526,N_22423,N_22296);
nand U22527 (N_22527,N_22026,N_22420);
nor U22528 (N_22528,N_21968,N_21883);
or U22529 (N_22529,N_22066,N_22303);
nor U22530 (N_22530,N_21992,N_22023);
nand U22531 (N_22531,N_22323,N_22310);
nor U22532 (N_22532,N_22392,N_22337);
and U22533 (N_22533,N_22087,N_22236);
xnor U22534 (N_22534,N_22000,N_22434);
nand U22535 (N_22535,N_22233,N_22091);
or U22536 (N_22536,N_22426,N_22286);
xnor U22537 (N_22537,N_22431,N_22329);
xnor U22538 (N_22538,N_21990,N_22141);
or U22539 (N_22539,N_22218,N_22128);
and U22540 (N_22540,N_22328,N_22136);
nand U22541 (N_22541,N_21909,N_22312);
xor U22542 (N_22542,N_22439,N_22429);
and U22543 (N_22543,N_22243,N_22054);
or U22544 (N_22544,N_22241,N_22248);
or U22545 (N_22545,N_21889,N_22130);
or U22546 (N_22546,N_22073,N_21954);
and U22547 (N_22547,N_22222,N_22186);
or U22548 (N_22548,N_22436,N_22076);
or U22549 (N_22549,N_22321,N_22240);
nor U22550 (N_22550,N_22193,N_22474);
and U22551 (N_22551,N_22069,N_21884);
and U22552 (N_22552,N_21942,N_22398);
nor U22553 (N_22553,N_22095,N_22368);
nor U22554 (N_22554,N_22466,N_22383);
nor U22555 (N_22555,N_22288,N_22083);
nor U22556 (N_22556,N_21994,N_22209);
nand U22557 (N_22557,N_22235,N_22278);
and U22558 (N_22558,N_22031,N_22144);
or U22559 (N_22559,N_22302,N_22096);
and U22560 (N_22560,N_22184,N_22100);
nor U22561 (N_22561,N_22492,N_22146);
xnor U22562 (N_22562,N_22124,N_22332);
xor U22563 (N_22563,N_21886,N_22497);
or U22564 (N_22564,N_22089,N_22009);
and U22565 (N_22565,N_22159,N_22020);
and U22566 (N_22566,N_22353,N_22113);
or U22567 (N_22567,N_21926,N_22160);
and U22568 (N_22568,N_22041,N_21985);
and U22569 (N_22569,N_22307,N_21998);
xnor U22570 (N_22570,N_22059,N_22443);
xnor U22571 (N_22571,N_21940,N_22195);
nand U22572 (N_22572,N_22148,N_21970);
and U22573 (N_22573,N_22281,N_22320);
nand U22574 (N_22574,N_22473,N_22494);
and U22575 (N_22575,N_22199,N_22357);
xor U22576 (N_22576,N_22211,N_22396);
nand U22577 (N_22577,N_22116,N_22154);
or U22578 (N_22578,N_22422,N_22464);
nand U22579 (N_22579,N_22458,N_22393);
nand U22580 (N_22580,N_22004,N_21988);
and U22581 (N_22581,N_21910,N_22168);
nor U22582 (N_22582,N_22018,N_22080);
xor U22583 (N_22583,N_21951,N_22200);
and U22584 (N_22584,N_22305,N_22250);
nand U22585 (N_22585,N_22378,N_22441);
nand U22586 (N_22586,N_22292,N_22298);
nor U22587 (N_22587,N_21948,N_21921);
nor U22588 (N_22588,N_22289,N_22155);
nand U22589 (N_22589,N_22061,N_21960);
xor U22590 (N_22590,N_22486,N_21891);
xor U22591 (N_22591,N_22215,N_22489);
nor U22592 (N_22592,N_22177,N_22462);
nand U22593 (N_22593,N_22265,N_22283);
xor U22594 (N_22594,N_22401,N_22263);
nor U22595 (N_22595,N_22125,N_22478);
or U22596 (N_22596,N_22389,N_22325);
nor U22597 (N_22597,N_22139,N_22395);
nand U22598 (N_22598,N_22427,N_22455);
or U22599 (N_22599,N_22121,N_22417);
nand U22600 (N_22600,N_22185,N_22264);
xor U22601 (N_22601,N_21966,N_22435);
nor U22602 (N_22602,N_21949,N_22493);
xor U22603 (N_22603,N_22287,N_22418);
nor U22604 (N_22604,N_22212,N_22063);
or U22605 (N_22605,N_22270,N_21906);
nand U22606 (N_22606,N_22050,N_22453);
nand U22607 (N_22607,N_21955,N_22359);
xnor U22608 (N_22608,N_22170,N_21878);
xnor U22609 (N_22609,N_21934,N_22447);
nor U22610 (N_22610,N_22174,N_22491);
or U22611 (N_22611,N_22346,N_22279);
and U22612 (N_22612,N_22088,N_22472);
and U22613 (N_22613,N_22364,N_21935);
or U22614 (N_22614,N_22126,N_22267);
nor U22615 (N_22615,N_21946,N_22386);
or U22616 (N_22616,N_22496,N_22324);
and U22617 (N_22617,N_21885,N_22268);
nor U22618 (N_22618,N_22077,N_22065);
and U22619 (N_22619,N_21894,N_22183);
and U22620 (N_22620,N_22207,N_21996);
xor U22621 (N_22621,N_22499,N_22227);
or U22622 (N_22622,N_22104,N_22381);
xnor U22623 (N_22623,N_22445,N_22475);
nand U22624 (N_22624,N_22327,N_22099);
and U22625 (N_22625,N_22414,N_21974);
nand U22626 (N_22626,N_22049,N_22345);
nand U22627 (N_22627,N_22118,N_21905);
nand U22628 (N_22628,N_22360,N_22382);
nor U22629 (N_22629,N_22165,N_22463);
xor U22630 (N_22630,N_22341,N_22335);
and U22631 (N_22631,N_22338,N_22068);
and U22632 (N_22632,N_22484,N_21941);
or U22633 (N_22633,N_22354,N_22074);
and U22634 (N_22634,N_21932,N_22457);
nor U22635 (N_22635,N_21947,N_22319);
nand U22636 (N_22636,N_22244,N_22203);
or U22637 (N_22637,N_22400,N_22367);
and U22638 (N_22638,N_22098,N_22019);
and U22639 (N_22639,N_22112,N_22032);
xnor U22640 (N_22640,N_21911,N_22220);
xnor U22641 (N_22641,N_22421,N_22348);
nand U22642 (N_22642,N_22142,N_22385);
or U22643 (N_22643,N_22316,N_22039);
nand U22644 (N_22644,N_22111,N_22079);
or U22645 (N_22645,N_22394,N_22487);
nor U22646 (N_22646,N_22008,N_22027);
and U22647 (N_22647,N_22123,N_22110);
or U22648 (N_22648,N_21965,N_21978);
nand U22649 (N_22649,N_22390,N_22311);
nand U22650 (N_22650,N_21887,N_22356);
nand U22651 (N_22651,N_22053,N_22376);
nor U22652 (N_22652,N_21931,N_21928);
or U22653 (N_22653,N_21899,N_22115);
nand U22654 (N_22654,N_21957,N_22430);
nor U22655 (N_22655,N_22133,N_21997);
and U22656 (N_22656,N_22415,N_22055);
and U22657 (N_22657,N_22047,N_22072);
and U22658 (N_22658,N_21890,N_22260);
xor U22659 (N_22659,N_21981,N_22274);
nor U22660 (N_22660,N_21904,N_21995);
nand U22661 (N_22661,N_22214,N_21963);
nand U22662 (N_22662,N_22397,N_22238);
nand U22663 (N_22663,N_22370,N_22369);
nand U22664 (N_22664,N_22219,N_22239);
xnor U22665 (N_22665,N_22064,N_21914);
or U22666 (N_22666,N_21922,N_22084);
nand U22667 (N_22667,N_22372,N_21973);
and U22668 (N_22668,N_22037,N_22082);
nand U22669 (N_22669,N_22167,N_22189);
and U22670 (N_22670,N_22010,N_22432);
and U22671 (N_22671,N_22045,N_22304);
nor U22672 (N_22672,N_22469,N_21980);
and U22673 (N_22673,N_21930,N_22442);
nand U22674 (N_22674,N_22085,N_22021);
nor U22675 (N_22675,N_22269,N_21976);
and U22676 (N_22676,N_22034,N_22366);
or U22677 (N_22677,N_22355,N_22003);
and U22678 (N_22678,N_22446,N_22038);
xnor U22679 (N_22679,N_21945,N_22150);
xnor U22680 (N_22680,N_22205,N_22282);
and U22681 (N_22681,N_22424,N_22229);
nor U22682 (N_22682,N_21936,N_21983);
nand U22683 (N_22683,N_22483,N_22127);
nor U22684 (N_22684,N_22058,N_22028);
and U22685 (N_22685,N_22153,N_22460);
nand U22686 (N_22686,N_21969,N_22490);
nand U22687 (N_22687,N_21989,N_21991);
and U22688 (N_22688,N_21882,N_22291);
xnor U22689 (N_22689,N_22450,N_22164);
nand U22690 (N_22690,N_22375,N_21897);
nor U22691 (N_22691,N_22103,N_22140);
or U22692 (N_22692,N_21918,N_22237);
and U22693 (N_22693,N_21915,N_22407);
xnor U22694 (N_22694,N_22336,N_22317);
nand U22695 (N_22695,N_22371,N_22197);
and U22696 (N_22696,N_22119,N_22191);
nand U22697 (N_22697,N_22482,N_22419);
and U22698 (N_22698,N_21919,N_22409);
or U22699 (N_22699,N_22230,N_22221);
nor U22700 (N_22700,N_22261,N_22071);
or U22701 (N_22701,N_22471,N_22280);
nor U22702 (N_22702,N_21961,N_22358);
nand U22703 (N_22703,N_21898,N_22408);
and U22704 (N_22704,N_22156,N_21933);
xnor U22705 (N_22705,N_21888,N_22258);
or U22706 (N_22706,N_22456,N_22070);
and U22707 (N_22707,N_22011,N_22086);
and U22708 (N_22708,N_22459,N_22030);
or U22709 (N_22709,N_21902,N_21986);
or U22710 (N_22710,N_22097,N_22495);
xnor U22711 (N_22711,N_22318,N_22347);
nor U22712 (N_22712,N_21895,N_22067);
xor U22713 (N_22713,N_22051,N_21893);
nand U22714 (N_22714,N_22388,N_22107);
nor U22715 (N_22715,N_22406,N_22242);
or U22716 (N_22716,N_22300,N_22294);
and U22717 (N_22717,N_22137,N_22313);
xor U22718 (N_22718,N_22194,N_22106);
or U22719 (N_22719,N_22391,N_22470);
or U22720 (N_22720,N_21938,N_22437);
nand U22721 (N_22721,N_22326,N_21880);
xor U22722 (N_22722,N_21962,N_22108);
or U22723 (N_22723,N_22012,N_22340);
nand U22724 (N_22724,N_22182,N_22259);
or U22725 (N_22725,N_22330,N_21953);
or U22726 (N_22726,N_22322,N_22465);
nand U22727 (N_22727,N_22301,N_21900);
xor U22728 (N_22728,N_21971,N_22204);
xnor U22729 (N_22729,N_22090,N_21943);
and U22730 (N_22730,N_22135,N_22006);
xnor U22731 (N_22731,N_22249,N_22129);
nor U22732 (N_22732,N_22210,N_21979);
nor U22733 (N_22733,N_22093,N_22213);
and U22734 (N_22734,N_22187,N_22105);
or U22735 (N_22735,N_22299,N_22295);
xor U22736 (N_22736,N_22308,N_21999);
nor U22737 (N_22737,N_22377,N_22277);
nor U22738 (N_22738,N_22285,N_22251);
or U22739 (N_22739,N_22351,N_21958);
and U22740 (N_22740,N_22246,N_21967);
and U22741 (N_22741,N_22223,N_21950);
or U22742 (N_22742,N_22425,N_22151);
or U22743 (N_22743,N_22339,N_22479);
xnor U22744 (N_22744,N_22373,N_21892);
and U22745 (N_22745,N_21903,N_22014);
xor U22746 (N_22746,N_22109,N_21877);
and U22747 (N_22747,N_22476,N_22024);
or U22748 (N_22748,N_22266,N_22498);
nor U22749 (N_22749,N_22078,N_21975);
nor U22750 (N_22750,N_21901,N_22402);
or U22751 (N_22751,N_22192,N_21924);
nor U22752 (N_22752,N_22043,N_22081);
or U22753 (N_22753,N_22225,N_22275);
and U22754 (N_22754,N_22331,N_22057);
and U22755 (N_22755,N_22309,N_22440);
or U22756 (N_22756,N_22273,N_22387);
xnor U22757 (N_22757,N_22171,N_22175);
nor U22758 (N_22758,N_22485,N_22232);
nor U22759 (N_22759,N_21881,N_22002);
nand U22760 (N_22760,N_22480,N_22179);
nor U22761 (N_22761,N_21896,N_22257);
nor U22762 (N_22762,N_22433,N_22132);
nor U22763 (N_22763,N_21952,N_22297);
nor U22764 (N_22764,N_22488,N_22315);
nand U22765 (N_22765,N_22362,N_22224);
nor U22766 (N_22766,N_22017,N_21944);
and U22767 (N_22767,N_22461,N_22046);
xor U22768 (N_22768,N_22293,N_22134);
nand U22769 (N_22769,N_22138,N_22481);
or U22770 (N_22770,N_22253,N_22044);
or U22771 (N_22771,N_22349,N_22056);
or U22772 (N_22772,N_22042,N_22217);
nand U22773 (N_22773,N_22196,N_22147);
nand U22774 (N_22774,N_22477,N_22262);
nor U22775 (N_22775,N_22314,N_21939);
nor U22776 (N_22776,N_22380,N_22255);
and U22777 (N_22777,N_22206,N_22117);
nand U22778 (N_22778,N_22208,N_22102);
and U22779 (N_22779,N_22352,N_22094);
xnor U22780 (N_22780,N_22226,N_21879);
or U22781 (N_22781,N_22143,N_22163);
and U22782 (N_22782,N_22405,N_22231);
or U22783 (N_22783,N_22350,N_22188);
or U22784 (N_22784,N_22438,N_22467);
or U22785 (N_22785,N_22404,N_22449);
nor U22786 (N_22786,N_22444,N_22172);
and U22787 (N_22787,N_22178,N_22176);
or U22788 (N_22788,N_21916,N_22374);
nand U22789 (N_22789,N_22180,N_22190);
nor U22790 (N_22790,N_22169,N_22201);
and U22791 (N_22791,N_22114,N_21937);
nor U22792 (N_22792,N_22342,N_22333);
and U22793 (N_22793,N_21876,N_22101);
or U22794 (N_22794,N_22361,N_22015);
xor U22795 (N_22795,N_22254,N_22276);
xnor U22796 (N_22796,N_22412,N_22149);
nor U22797 (N_22797,N_21956,N_22198);
and U22798 (N_22798,N_22162,N_22181);
and U22799 (N_22799,N_22161,N_21925);
nor U22800 (N_22800,N_22022,N_22029);
or U22801 (N_22801,N_21984,N_21972);
xnor U22802 (N_22802,N_21982,N_22363);
and U22803 (N_22803,N_22428,N_22120);
and U22804 (N_22804,N_22403,N_22272);
nor U22805 (N_22805,N_22033,N_22035);
xor U22806 (N_22806,N_22092,N_22013);
and U22807 (N_22807,N_22247,N_22448);
xor U22808 (N_22808,N_22001,N_22036);
nor U22809 (N_22809,N_22284,N_22005);
nor U22810 (N_22810,N_22468,N_22234);
nor U22811 (N_22811,N_22040,N_22166);
xor U22812 (N_22812,N_22411,N_22272);
nor U22813 (N_22813,N_22124,N_22257);
or U22814 (N_22814,N_22103,N_21914);
nand U22815 (N_22815,N_22260,N_21931);
xnor U22816 (N_22816,N_22166,N_22407);
nand U22817 (N_22817,N_21920,N_22030);
and U22818 (N_22818,N_22424,N_22118);
xnor U22819 (N_22819,N_22113,N_22230);
nor U22820 (N_22820,N_22129,N_21946);
nand U22821 (N_22821,N_22017,N_22389);
xor U22822 (N_22822,N_22348,N_21905);
xor U22823 (N_22823,N_21937,N_21996);
xor U22824 (N_22824,N_22385,N_22465);
or U22825 (N_22825,N_22412,N_21926);
or U22826 (N_22826,N_22276,N_22293);
and U22827 (N_22827,N_22382,N_22078);
nor U22828 (N_22828,N_21997,N_22099);
or U22829 (N_22829,N_21924,N_21886);
nor U22830 (N_22830,N_22303,N_22005);
or U22831 (N_22831,N_21899,N_22462);
xnor U22832 (N_22832,N_22315,N_22325);
nor U22833 (N_22833,N_22158,N_22428);
or U22834 (N_22834,N_22020,N_22176);
and U22835 (N_22835,N_21926,N_22161);
nand U22836 (N_22836,N_22346,N_22430);
and U22837 (N_22837,N_22293,N_21992);
nor U22838 (N_22838,N_21990,N_22405);
and U22839 (N_22839,N_22033,N_22411);
or U22840 (N_22840,N_22064,N_22223);
nor U22841 (N_22841,N_22396,N_22174);
xnor U22842 (N_22842,N_21968,N_22282);
xnor U22843 (N_22843,N_21928,N_22001);
xnor U22844 (N_22844,N_21921,N_22222);
nand U22845 (N_22845,N_21965,N_21887);
or U22846 (N_22846,N_22073,N_22146);
xnor U22847 (N_22847,N_21948,N_22211);
nand U22848 (N_22848,N_22060,N_22077);
nor U22849 (N_22849,N_22436,N_22374);
and U22850 (N_22850,N_22110,N_21982);
nand U22851 (N_22851,N_22087,N_22484);
or U22852 (N_22852,N_21894,N_22306);
and U22853 (N_22853,N_21942,N_22107);
nor U22854 (N_22854,N_21897,N_22192);
nand U22855 (N_22855,N_22437,N_22029);
nand U22856 (N_22856,N_22130,N_21929);
nor U22857 (N_22857,N_22265,N_22028);
or U22858 (N_22858,N_22267,N_22094);
or U22859 (N_22859,N_22309,N_21981);
xor U22860 (N_22860,N_22459,N_22224);
or U22861 (N_22861,N_21891,N_22009);
nand U22862 (N_22862,N_22000,N_22181);
or U22863 (N_22863,N_21925,N_22436);
nor U22864 (N_22864,N_22359,N_21926);
nand U22865 (N_22865,N_22364,N_21943);
xnor U22866 (N_22866,N_21885,N_22203);
xor U22867 (N_22867,N_21958,N_21993);
and U22868 (N_22868,N_22215,N_22323);
or U22869 (N_22869,N_22431,N_21895);
and U22870 (N_22870,N_22160,N_22161);
xor U22871 (N_22871,N_22054,N_22205);
xor U22872 (N_22872,N_22052,N_22369);
and U22873 (N_22873,N_22273,N_22421);
nor U22874 (N_22874,N_22310,N_21952);
or U22875 (N_22875,N_22422,N_22498);
or U22876 (N_22876,N_22202,N_21970);
nor U22877 (N_22877,N_21984,N_22194);
xnor U22878 (N_22878,N_22028,N_22071);
nor U22879 (N_22879,N_21934,N_22120);
xnor U22880 (N_22880,N_22292,N_22301);
xnor U22881 (N_22881,N_22246,N_22291);
or U22882 (N_22882,N_22021,N_22456);
xor U22883 (N_22883,N_22325,N_22364);
or U22884 (N_22884,N_22410,N_22398);
nor U22885 (N_22885,N_21995,N_22459);
nor U22886 (N_22886,N_22231,N_21941);
nor U22887 (N_22887,N_22357,N_22452);
or U22888 (N_22888,N_22364,N_22343);
and U22889 (N_22889,N_22205,N_22002);
nor U22890 (N_22890,N_22225,N_21895);
nor U22891 (N_22891,N_22152,N_21919);
and U22892 (N_22892,N_22098,N_22028);
or U22893 (N_22893,N_21947,N_22476);
nand U22894 (N_22894,N_22455,N_21933);
xor U22895 (N_22895,N_22187,N_22075);
nand U22896 (N_22896,N_21972,N_22071);
xnor U22897 (N_22897,N_21947,N_22341);
and U22898 (N_22898,N_22478,N_21918);
nor U22899 (N_22899,N_21882,N_22406);
xnor U22900 (N_22900,N_22130,N_21959);
or U22901 (N_22901,N_22397,N_22285);
nand U22902 (N_22902,N_22274,N_22195);
and U22903 (N_22903,N_22417,N_21884);
or U22904 (N_22904,N_22146,N_22179);
and U22905 (N_22905,N_22246,N_22089);
xnor U22906 (N_22906,N_21934,N_22497);
nand U22907 (N_22907,N_22042,N_22194);
and U22908 (N_22908,N_22042,N_22295);
nand U22909 (N_22909,N_22425,N_22398);
nor U22910 (N_22910,N_21901,N_22230);
xnor U22911 (N_22911,N_22260,N_22123);
nor U22912 (N_22912,N_21986,N_21886);
and U22913 (N_22913,N_22380,N_22030);
nor U22914 (N_22914,N_22252,N_22322);
and U22915 (N_22915,N_21935,N_21976);
xor U22916 (N_22916,N_21875,N_22169);
or U22917 (N_22917,N_22287,N_22387);
nor U22918 (N_22918,N_22467,N_21881);
nor U22919 (N_22919,N_22395,N_22155);
and U22920 (N_22920,N_22475,N_22419);
xnor U22921 (N_22921,N_22215,N_22191);
or U22922 (N_22922,N_22363,N_22017);
or U22923 (N_22923,N_22329,N_22158);
or U22924 (N_22924,N_22004,N_21982);
nand U22925 (N_22925,N_22454,N_22245);
xor U22926 (N_22926,N_22355,N_22474);
xnor U22927 (N_22927,N_22123,N_22120);
xnor U22928 (N_22928,N_22055,N_22440);
nand U22929 (N_22929,N_22345,N_22385);
nor U22930 (N_22930,N_22457,N_22147);
xor U22931 (N_22931,N_21929,N_22039);
nor U22932 (N_22932,N_22161,N_22375);
nor U22933 (N_22933,N_22216,N_21978);
xnor U22934 (N_22934,N_22381,N_22126);
nand U22935 (N_22935,N_22272,N_21997);
nand U22936 (N_22936,N_22316,N_22393);
nor U22937 (N_22937,N_22348,N_22297);
nand U22938 (N_22938,N_21940,N_22460);
xnor U22939 (N_22939,N_22048,N_22104);
or U22940 (N_22940,N_22173,N_22145);
or U22941 (N_22941,N_22251,N_22244);
nand U22942 (N_22942,N_22094,N_22315);
nor U22943 (N_22943,N_22379,N_22473);
nand U22944 (N_22944,N_21879,N_22476);
xnor U22945 (N_22945,N_22219,N_22491);
nor U22946 (N_22946,N_22063,N_22035);
nor U22947 (N_22947,N_22273,N_22308);
nand U22948 (N_22948,N_22286,N_22131);
nand U22949 (N_22949,N_22473,N_22257);
nor U22950 (N_22950,N_22270,N_22035);
or U22951 (N_22951,N_22088,N_22327);
nor U22952 (N_22952,N_21880,N_21909);
nand U22953 (N_22953,N_22451,N_21908);
xor U22954 (N_22954,N_22161,N_22439);
or U22955 (N_22955,N_21884,N_22309);
and U22956 (N_22956,N_22263,N_22360);
or U22957 (N_22957,N_22313,N_21890);
xor U22958 (N_22958,N_22114,N_22172);
or U22959 (N_22959,N_21957,N_22136);
nor U22960 (N_22960,N_22128,N_22311);
nand U22961 (N_22961,N_22398,N_22464);
nor U22962 (N_22962,N_22479,N_22188);
xor U22963 (N_22963,N_22324,N_22056);
nor U22964 (N_22964,N_22363,N_22106);
nand U22965 (N_22965,N_22234,N_22136);
nor U22966 (N_22966,N_22417,N_22230);
nand U22967 (N_22967,N_22283,N_22154);
nor U22968 (N_22968,N_22272,N_22275);
xor U22969 (N_22969,N_22484,N_22388);
xor U22970 (N_22970,N_22298,N_22169);
or U22971 (N_22971,N_22290,N_22193);
or U22972 (N_22972,N_22274,N_22016);
nand U22973 (N_22973,N_22075,N_22304);
nand U22974 (N_22974,N_22065,N_22449);
nand U22975 (N_22975,N_22443,N_22041);
xnor U22976 (N_22976,N_22471,N_22326);
or U22977 (N_22977,N_21927,N_22304);
xnor U22978 (N_22978,N_21899,N_22358);
or U22979 (N_22979,N_22262,N_22467);
and U22980 (N_22980,N_22261,N_21896);
xor U22981 (N_22981,N_22315,N_22365);
nor U22982 (N_22982,N_22220,N_22063);
or U22983 (N_22983,N_22489,N_22323);
or U22984 (N_22984,N_22282,N_22459);
nor U22985 (N_22985,N_21919,N_22344);
or U22986 (N_22986,N_22160,N_21982);
xor U22987 (N_22987,N_22155,N_21968);
nand U22988 (N_22988,N_22485,N_22002);
nand U22989 (N_22989,N_22176,N_22048);
nor U22990 (N_22990,N_22151,N_22069);
or U22991 (N_22991,N_21878,N_21934);
nand U22992 (N_22992,N_22352,N_21917);
nor U22993 (N_22993,N_22450,N_21984);
nand U22994 (N_22994,N_22216,N_22003);
xnor U22995 (N_22995,N_21935,N_22053);
or U22996 (N_22996,N_22066,N_22174);
nand U22997 (N_22997,N_21889,N_22068);
xor U22998 (N_22998,N_21930,N_22453);
and U22999 (N_22999,N_22442,N_21933);
xnor U23000 (N_23000,N_22202,N_22156);
and U23001 (N_23001,N_22249,N_22234);
nand U23002 (N_23002,N_22022,N_22374);
or U23003 (N_23003,N_22073,N_21966);
xnor U23004 (N_23004,N_22218,N_22419);
and U23005 (N_23005,N_22375,N_21876);
or U23006 (N_23006,N_22276,N_22114);
nor U23007 (N_23007,N_22072,N_22133);
or U23008 (N_23008,N_21933,N_22248);
or U23009 (N_23009,N_21997,N_22485);
xor U23010 (N_23010,N_22057,N_22047);
nor U23011 (N_23011,N_22248,N_22287);
nand U23012 (N_23012,N_21971,N_22289);
nand U23013 (N_23013,N_21908,N_22080);
xnor U23014 (N_23014,N_22148,N_22060);
nor U23015 (N_23015,N_22178,N_22395);
xnor U23016 (N_23016,N_22199,N_22303);
xor U23017 (N_23017,N_22064,N_22000);
and U23018 (N_23018,N_21968,N_22273);
nor U23019 (N_23019,N_22407,N_22275);
nand U23020 (N_23020,N_22401,N_22472);
nand U23021 (N_23021,N_22182,N_21976);
xor U23022 (N_23022,N_21940,N_21882);
and U23023 (N_23023,N_22456,N_22402);
or U23024 (N_23024,N_22436,N_21918);
or U23025 (N_23025,N_22320,N_22330);
or U23026 (N_23026,N_22080,N_22127);
nand U23027 (N_23027,N_22464,N_21926);
nand U23028 (N_23028,N_22410,N_21916);
xnor U23029 (N_23029,N_22100,N_22324);
nor U23030 (N_23030,N_22051,N_22123);
nor U23031 (N_23031,N_22150,N_22040);
or U23032 (N_23032,N_22183,N_22171);
or U23033 (N_23033,N_21895,N_22289);
nor U23034 (N_23034,N_22485,N_22467);
nor U23035 (N_23035,N_22069,N_21905);
nor U23036 (N_23036,N_22155,N_22329);
nand U23037 (N_23037,N_22075,N_22329);
and U23038 (N_23038,N_22065,N_22321);
nand U23039 (N_23039,N_22086,N_22046);
or U23040 (N_23040,N_21883,N_22020);
nand U23041 (N_23041,N_21898,N_22478);
nand U23042 (N_23042,N_22469,N_22321);
nand U23043 (N_23043,N_22327,N_21884);
and U23044 (N_23044,N_21885,N_22458);
and U23045 (N_23045,N_22121,N_22423);
nor U23046 (N_23046,N_22206,N_22327);
xnor U23047 (N_23047,N_21931,N_22344);
xor U23048 (N_23048,N_22062,N_22253);
nand U23049 (N_23049,N_21996,N_22094);
xnor U23050 (N_23050,N_22156,N_22295);
nand U23051 (N_23051,N_22252,N_22349);
and U23052 (N_23052,N_21912,N_22031);
nor U23053 (N_23053,N_22042,N_22424);
xor U23054 (N_23054,N_22377,N_22362);
xor U23055 (N_23055,N_22236,N_22064);
and U23056 (N_23056,N_22351,N_22342);
nor U23057 (N_23057,N_22284,N_22412);
nand U23058 (N_23058,N_22180,N_22476);
or U23059 (N_23059,N_22202,N_22164);
or U23060 (N_23060,N_21906,N_22020);
nand U23061 (N_23061,N_22424,N_21914);
xnor U23062 (N_23062,N_21876,N_22393);
nand U23063 (N_23063,N_22285,N_21949);
nor U23064 (N_23064,N_22177,N_22402);
nand U23065 (N_23065,N_22251,N_22468);
nand U23066 (N_23066,N_22090,N_22079);
and U23067 (N_23067,N_21987,N_21917);
nand U23068 (N_23068,N_22314,N_21875);
and U23069 (N_23069,N_22490,N_22467);
nand U23070 (N_23070,N_22282,N_22045);
xnor U23071 (N_23071,N_22466,N_22145);
xor U23072 (N_23072,N_22038,N_22228);
nor U23073 (N_23073,N_22069,N_22084);
or U23074 (N_23074,N_22353,N_22158);
nor U23075 (N_23075,N_22393,N_22397);
xnor U23076 (N_23076,N_22307,N_22488);
nor U23077 (N_23077,N_21960,N_22153);
nand U23078 (N_23078,N_22154,N_22461);
nand U23079 (N_23079,N_22250,N_22064);
xnor U23080 (N_23080,N_22221,N_22050);
and U23081 (N_23081,N_22059,N_22024);
nor U23082 (N_23082,N_22496,N_22131);
and U23083 (N_23083,N_22277,N_22376);
nor U23084 (N_23084,N_22081,N_22098);
nand U23085 (N_23085,N_22410,N_21980);
and U23086 (N_23086,N_22016,N_22300);
xnor U23087 (N_23087,N_22495,N_22151);
or U23088 (N_23088,N_22097,N_22203);
and U23089 (N_23089,N_22433,N_22251);
or U23090 (N_23090,N_21948,N_22210);
or U23091 (N_23091,N_22402,N_21890);
nand U23092 (N_23092,N_22221,N_22247);
and U23093 (N_23093,N_22095,N_22013);
or U23094 (N_23094,N_22191,N_22409);
nor U23095 (N_23095,N_22299,N_22112);
xnor U23096 (N_23096,N_22461,N_21995);
or U23097 (N_23097,N_22328,N_21943);
nand U23098 (N_23098,N_22402,N_22054);
nand U23099 (N_23099,N_22063,N_21968);
xor U23100 (N_23100,N_22489,N_22151);
xnor U23101 (N_23101,N_22245,N_22498);
and U23102 (N_23102,N_22317,N_22258);
nor U23103 (N_23103,N_22388,N_22211);
xnor U23104 (N_23104,N_22136,N_21908);
nand U23105 (N_23105,N_22392,N_22464);
and U23106 (N_23106,N_21931,N_22119);
or U23107 (N_23107,N_22051,N_22249);
and U23108 (N_23108,N_22050,N_22199);
nor U23109 (N_23109,N_22239,N_21977);
nand U23110 (N_23110,N_22300,N_22095);
xnor U23111 (N_23111,N_21883,N_22472);
or U23112 (N_23112,N_22274,N_22300);
nor U23113 (N_23113,N_22154,N_22125);
and U23114 (N_23114,N_22028,N_22453);
nor U23115 (N_23115,N_22232,N_22236);
and U23116 (N_23116,N_22463,N_22199);
and U23117 (N_23117,N_22167,N_21900);
nand U23118 (N_23118,N_22067,N_22212);
or U23119 (N_23119,N_22098,N_22477);
nor U23120 (N_23120,N_22002,N_22186);
nand U23121 (N_23121,N_22315,N_22090);
nor U23122 (N_23122,N_22431,N_22231);
xnor U23123 (N_23123,N_21952,N_22205);
nor U23124 (N_23124,N_21973,N_22061);
xor U23125 (N_23125,N_22782,N_22674);
nand U23126 (N_23126,N_22758,N_22853);
or U23127 (N_23127,N_22553,N_22742);
nor U23128 (N_23128,N_22880,N_22883);
nor U23129 (N_23129,N_22551,N_22893);
xor U23130 (N_23130,N_22860,N_22799);
and U23131 (N_23131,N_22868,N_22672);
nand U23132 (N_23132,N_23087,N_22554);
and U23133 (N_23133,N_22818,N_22733);
nand U23134 (N_23134,N_23081,N_22980);
and U23135 (N_23135,N_23031,N_22641);
nor U23136 (N_23136,N_23078,N_22747);
nand U23137 (N_23137,N_23082,N_22690);
xnor U23138 (N_23138,N_23062,N_23022);
nand U23139 (N_23139,N_22710,N_22970);
and U23140 (N_23140,N_22723,N_22768);
nor U23141 (N_23141,N_22812,N_23013);
nand U23142 (N_23142,N_22685,N_22502);
nor U23143 (N_23143,N_22523,N_22531);
nor U23144 (N_23144,N_22509,N_22585);
nand U23145 (N_23145,N_22850,N_22726);
or U23146 (N_23146,N_22587,N_22591);
or U23147 (N_23147,N_22953,N_22656);
and U23148 (N_23148,N_22937,N_23079);
and U23149 (N_23149,N_22678,N_22862);
xor U23150 (N_23150,N_22790,N_22892);
or U23151 (N_23151,N_22962,N_22612);
and U23152 (N_23152,N_22786,N_22569);
nor U23153 (N_23153,N_22722,N_22595);
nand U23154 (N_23154,N_22965,N_22615);
or U23155 (N_23155,N_23097,N_23024);
xor U23156 (N_23156,N_22944,N_22545);
xnor U23157 (N_23157,N_22929,N_23027);
nor U23158 (N_23158,N_22597,N_22703);
nand U23159 (N_23159,N_22817,N_22847);
and U23160 (N_23160,N_23019,N_23110);
and U23161 (N_23161,N_23069,N_23007);
nor U23162 (N_23162,N_22671,N_22842);
nand U23163 (N_23163,N_22661,N_22804);
nor U23164 (N_23164,N_22986,N_22665);
nor U23165 (N_23165,N_23074,N_22631);
nand U23166 (N_23166,N_22992,N_23002);
nand U23167 (N_23167,N_23039,N_22561);
nor U23168 (N_23168,N_22739,N_22990);
and U23169 (N_23169,N_22697,N_22568);
xnor U23170 (N_23170,N_22634,N_23124);
xnor U23171 (N_23171,N_22759,N_23016);
xnor U23172 (N_23172,N_22978,N_22844);
or U23173 (N_23173,N_22838,N_22789);
or U23174 (N_23174,N_22760,N_22874);
nor U23175 (N_23175,N_22548,N_22550);
nor U23176 (N_23176,N_22943,N_23015);
nor U23177 (N_23177,N_23086,N_22624);
and U23178 (N_23178,N_22754,N_22834);
or U23179 (N_23179,N_23080,N_22610);
nor U23180 (N_23180,N_22598,N_22859);
and U23181 (N_23181,N_22903,N_22899);
nor U23182 (N_23182,N_22865,N_22887);
nor U23183 (N_23183,N_22907,N_22520);
or U23184 (N_23184,N_22813,N_22642);
and U23185 (N_23185,N_23041,N_22904);
or U23186 (N_23186,N_22711,N_22777);
and U23187 (N_23187,N_23059,N_23049);
or U23188 (N_23188,N_22967,N_22979);
xnor U23189 (N_23189,N_22781,N_22919);
and U23190 (N_23190,N_22830,N_22625);
xor U23191 (N_23191,N_22575,N_22906);
or U23192 (N_23192,N_22651,N_22670);
nand U23193 (N_23193,N_22994,N_22989);
xor U23194 (N_23194,N_22511,N_22749);
xor U23195 (N_23195,N_22572,N_22856);
or U23196 (N_23196,N_22900,N_23088);
and U23197 (N_23197,N_22521,N_22636);
or U23198 (N_23198,N_22748,N_22622);
or U23199 (N_23199,N_22829,N_22995);
nor U23200 (N_23200,N_22955,N_22730);
or U23201 (N_23201,N_22767,N_22629);
nor U23202 (N_23202,N_22846,N_22526);
nand U23203 (N_23203,N_22596,N_22996);
and U23204 (N_23204,N_23004,N_22626);
and U23205 (N_23205,N_22650,N_23073);
or U23206 (N_23206,N_22512,N_22924);
and U23207 (N_23207,N_22773,N_22620);
or U23208 (N_23208,N_22774,N_22869);
or U23209 (N_23209,N_22934,N_22873);
or U23210 (N_23210,N_23030,N_23018);
nor U23211 (N_23211,N_22713,N_23098);
nand U23212 (N_23212,N_22762,N_22606);
nand U23213 (N_23213,N_22617,N_22926);
nand U23214 (N_23214,N_22673,N_23050);
or U23215 (N_23215,N_22562,N_22699);
nor U23216 (N_23216,N_22503,N_22588);
xor U23217 (N_23217,N_23120,N_22770);
nand U23218 (N_23218,N_22935,N_23076);
or U23219 (N_23219,N_23113,N_22542);
or U23220 (N_23220,N_22825,N_22788);
and U23221 (N_23221,N_22821,N_22922);
nor U23222 (N_23222,N_22677,N_23033);
nand U23223 (N_23223,N_22779,N_22913);
or U23224 (N_23224,N_22780,N_22957);
nor U23225 (N_23225,N_23001,N_22513);
or U23226 (N_23226,N_23063,N_22536);
or U23227 (N_23227,N_22753,N_22810);
nand U23228 (N_23228,N_22566,N_22921);
and U23229 (N_23229,N_23005,N_22993);
nor U23230 (N_23230,N_23053,N_22556);
nand U23231 (N_23231,N_22910,N_22525);
or U23232 (N_23232,N_22707,N_22614);
xor U23233 (N_23233,N_22586,N_23023);
or U23234 (N_23234,N_22991,N_22682);
nand U23235 (N_23235,N_22949,N_22756);
and U23236 (N_23236,N_22816,N_22579);
nor U23237 (N_23237,N_22982,N_22832);
nand U23238 (N_23238,N_22942,N_22558);
nand U23239 (N_23239,N_22669,N_22696);
or U23240 (N_23240,N_22911,N_22960);
or U23241 (N_23241,N_22776,N_23020);
and U23242 (N_23242,N_22968,N_22538);
and U23243 (N_23243,N_22839,N_22959);
nor U23244 (N_23244,N_22765,N_22801);
or U23245 (N_23245,N_22950,N_22695);
or U23246 (N_23246,N_22952,N_22643);
xor U23247 (N_23247,N_22743,N_22735);
xor U23248 (N_23248,N_22870,N_22852);
nor U23249 (N_23249,N_22964,N_22826);
nor U23250 (N_23250,N_23094,N_23077);
xnor U23251 (N_23251,N_22909,N_22985);
nand U23252 (N_23252,N_22981,N_22527);
or U23253 (N_23253,N_23012,N_22941);
nor U23254 (N_23254,N_22824,N_22709);
nand U23255 (N_23255,N_23032,N_22951);
and U23256 (N_23256,N_22702,N_22731);
nand U23257 (N_23257,N_22803,N_23105);
nor U23258 (N_23258,N_23096,N_22795);
nand U23259 (N_23259,N_22515,N_22637);
nand U23260 (N_23260,N_22822,N_22508);
xor U23261 (N_23261,N_22772,N_23090);
xnor U23262 (N_23262,N_23047,N_22918);
nand U23263 (N_23263,N_22505,N_23009);
xor U23264 (N_23264,N_22717,N_23035);
and U23265 (N_23265,N_23104,N_22895);
nor U23266 (N_23266,N_22741,N_22891);
or U23267 (N_23267,N_22655,N_22882);
nand U23268 (N_23268,N_22798,N_23021);
xnor U23269 (N_23269,N_22657,N_22744);
nor U23270 (N_23270,N_22963,N_22507);
xor U23271 (N_23271,N_22712,N_22524);
or U23272 (N_23272,N_22522,N_22623);
and U23273 (N_23273,N_22608,N_22987);
nor U23274 (N_23274,N_22835,N_22914);
or U23275 (N_23275,N_22532,N_22787);
nor U23276 (N_23276,N_22607,N_22500);
or U23277 (N_23277,N_22886,N_22871);
nand U23278 (N_23278,N_22947,N_22530);
xnor U23279 (N_23279,N_22881,N_22589);
xnor U23280 (N_23280,N_22808,N_22931);
or U23281 (N_23281,N_22783,N_22755);
or U23282 (N_23282,N_22890,N_22724);
nand U23283 (N_23283,N_22611,N_23109);
xnor U23284 (N_23284,N_23122,N_22750);
nand U23285 (N_23285,N_22577,N_22796);
nor U23286 (N_23286,N_22855,N_22811);
and U23287 (N_23287,N_22872,N_22815);
nand U23288 (N_23288,N_22592,N_22889);
xnor U23289 (N_23289,N_22543,N_22720);
nand U23290 (N_23290,N_22590,N_23048);
nand U23291 (N_23291,N_22653,N_23101);
and U23292 (N_23292,N_22603,N_22570);
nand U23293 (N_23293,N_22529,N_22763);
and U23294 (N_23294,N_22633,N_22836);
or U23295 (N_23295,N_22605,N_22833);
and U23296 (N_23296,N_22721,N_23107);
and U23297 (N_23297,N_22948,N_23034);
or U23298 (N_23298,N_22632,N_22698);
or U23299 (N_23299,N_22557,N_22706);
and U23300 (N_23300,N_22769,N_23055);
or U23301 (N_23301,N_22567,N_22714);
and U23302 (N_23302,N_23091,N_22635);
or U23303 (N_23303,N_22686,N_23085);
or U23304 (N_23304,N_22564,N_23067);
and U23305 (N_23305,N_22814,N_22761);
and U23306 (N_23306,N_22679,N_23075);
and U23307 (N_23307,N_22877,N_22849);
nor U23308 (N_23308,N_22647,N_23036);
xor U23309 (N_23309,N_23052,N_22501);
nor U23310 (N_23310,N_22648,N_22676);
nand U23311 (N_23311,N_23008,N_22885);
nand U23312 (N_23312,N_22738,N_23037);
nor U23313 (N_23313,N_22716,N_22820);
and U23314 (N_23314,N_22983,N_22658);
xnor U23315 (N_23315,N_22583,N_22694);
or U23316 (N_23316,N_22547,N_22976);
xor U23317 (N_23317,N_22519,N_22728);
nand U23318 (N_23318,N_22969,N_22928);
nor U23319 (N_23319,N_22565,N_22664);
nor U23320 (N_23320,N_22863,N_23111);
or U23321 (N_23321,N_23014,N_22546);
xnor U23322 (N_23322,N_22932,N_22923);
xor U23323 (N_23323,N_22560,N_22571);
and U23324 (N_23324,N_22630,N_23003);
nor U23325 (N_23325,N_23084,N_22876);
nor U23326 (N_23326,N_22725,N_22604);
nor U23327 (N_23327,N_22708,N_23100);
nand U23328 (N_23328,N_22660,N_22884);
and U23329 (N_23329,N_22974,N_22927);
and U23330 (N_23330,N_22640,N_23000);
and U23331 (N_23331,N_23102,N_23011);
nand U23332 (N_23332,N_22866,N_22574);
nor U23333 (N_23333,N_23114,N_22602);
nand U23334 (N_23334,N_22514,N_22966);
or U23335 (N_23335,N_22535,N_23006);
nor U23336 (N_23336,N_22652,N_23061);
nor U23337 (N_23337,N_22766,N_22794);
nand U23338 (N_23338,N_22687,N_22659);
and U23339 (N_23339,N_22867,N_22563);
xnor U23340 (N_23340,N_22619,N_22840);
xor U23341 (N_23341,N_22704,N_22896);
nor U23342 (N_23342,N_22800,N_22613);
xor U23343 (N_23343,N_22516,N_22930);
xnor U23344 (N_23344,N_22646,N_22997);
and U23345 (N_23345,N_22792,N_22578);
or U23346 (N_23346,N_23068,N_22977);
nand U23347 (N_23347,N_22912,N_22793);
or U23348 (N_23348,N_22719,N_23043);
and U23349 (N_23349,N_22837,N_22946);
nor U23350 (N_23350,N_22540,N_22681);
nor U23351 (N_23351,N_23115,N_22878);
nand U23352 (N_23352,N_23064,N_22544);
or U23353 (N_23353,N_23093,N_22954);
xor U23354 (N_23354,N_22864,N_23108);
nand U23355 (N_23355,N_22601,N_22654);
and U23356 (N_23356,N_22745,N_22666);
and U23357 (N_23357,N_23025,N_22639);
xor U23358 (N_23358,N_22933,N_22580);
nand U23359 (N_23359,N_22584,N_23042);
nor U23360 (N_23360,N_22541,N_22823);
nor U23361 (N_23361,N_22689,N_23071);
or U23362 (N_23362,N_23095,N_23044);
xnor U23363 (N_23363,N_22938,N_23103);
and U23364 (N_23364,N_22549,N_22667);
xor U23365 (N_23365,N_22688,N_22925);
or U23366 (N_23366,N_22843,N_23058);
nand U23367 (N_23367,N_22668,N_23051);
xor U23368 (N_23368,N_22751,N_22700);
nand U23369 (N_23369,N_22827,N_22573);
or U23370 (N_23370,N_22675,N_22627);
and U23371 (N_23371,N_23038,N_23028);
or U23372 (N_23372,N_22740,N_22854);
nor U23373 (N_23373,N_22785,N_22888);
or U23374 (N_23374,N_22845,N_22936);
and U23375 (N_23375,N_22851,N_22701);
or U23376 (N_23376,N_22594,N_22528);
and U23377 (N_23377,N_22534,N_23045);
nor U23378 (N_23378,N_23070,N_23119);
and U23379 (N_23379,N_22680,N_22757);
or U23380 (N_23380,N_23057,N_22807);
and U23381 (N_23381,N_22752,N_22533);
nor U23382 (N_23382,N_22539,N_22555);
nand U23383 (N_23383,N_22537,N_22736);
or U23384 (N_23384,N_23099,N_22894);
or U23385 (N_23385,N_22645,N_22662);
or U23386 (N_23386,N_22729,N_22940);
nor U23387 (N_23387,N_22841,N_23066);
xor U23388 (N_23388,N_23060,N_23121);
nand U23389 (N_23389,N_23117,N_23083);
nor U23390 (N_23390,N_22809,N_22999);
nor U23391 (N_23391,N_22879,N_23072);
or U23392 (N_23392,N_22691,N_22504);
and U23393 (N_23393,N_23118,N_22599);
and U23394 (N_23394,N_22732,N_23092);
nand U23395 (N_23395,N_22971,N_22975);
nand U23396 (N_23396,N_22734,N_23046);
and U23397 (N_23397,N_22908,N_23010);
nor U23398 (N_23398,N_22897,N_23017);
nor U23399 (N_23399,N_22791,N_22684);
nor U23400 (N_23400,N_23040,N_22618);
xor U23401 (N_23401,N_22875,N_22663);
or U23402 (N_23402,N_22559,N_23112);
and U23403 (N_23403,N_22784,N_22915);
or U23404 (N_23404,N_22984,N_22857);
or U23405 (N_23405,N_22902,N_22806);
or U23406 (N_23406,N_22693,N_22861);
xor U23407 (N_23407,N_22746,N_22621);
nor U23408 (N_23408,N_22972,N_23029);
and U23409 (N_23409,N_22958,N_22998);
or U23410 (N_23410,N_23089,N_22988);
nand U23411 (N_23411,N_22973,N_23026);
xor U23412 (N_23412,N_22778,N_22775);
and U23413 (N_23413,N_23054,N_22805);
xor U23414 (N_23414,N_22901,N_22715);
nand U23415 (N_23415,N_22848,N_22920);
nand U23416 (N_23416,N_22916,N_23056);
and U23417 (N_23417,N_22518,N_22939);
xor U23418 (N_23418,N_22510,N_22797);
nor U23419 (N_23419,N_23123,N_22517);
nand U23420 (N_23420,N_22616,N_22905);
and U23421 (N_23421,N_22718,N_22764);
xnor U23422 (N_23422,N_22945,N_23065);
and U23423 (N_23423,N_22858,N_22581);
nand U23424 (N_23424,N_22506,N_22600);
and U23425 (N_23425,N_22831,N_22705);
nand U23426 (N_23426,N_22582,N_22638);
and U23427 (N_23427,N_22737,N_22609);
or U23428 (N_23428,N_22683,N_22644);
xnor U23429 (N_23429,N_22961,N_22898);
xnor U23430 (N_23430,N_22649,N_22828);
and U23431 (N_23431,N_22956,N_22771);
and U23432 (N_23432,N_22692,N_23116);
and U23433 (N_23433,N_22628,N_22802);
xor U23434 (N_23434,N_23106,N_22917);
nand U23435 (N_23435,N_22819,N_22593);
xor U23436 (N_23436,N_22727,N_22552);
nand U23437 (N_23437,N_22576,N_22650);
nor U23438 (N_23438,N_22751,N_22832);
and U23439 (N_23439,N_22549,N_22899);
and U23440 (N_23440,N_22799,N_22701);
nand U23441 (N_23441,N_22544,N_23069);
and U23442 (N_23442,N_22572,N_22865);
or U23443 (N_23443,N_22714,N_22894);
or U23444 (N_23444,N_22780,N_22774);
xnor U23445 (N_23445,N_22863,N_23106);
nand U23446 (N_23446,N_22900,N_22865);
or U23447 (N_23447,N_22739,N_22750);
and U23448 (N_23448,N_23028,N_23037);
nor U23449 (N_23449,N_22597,N_22958);
and U23450 (N_23450,N_22626,N_22738);
nand U23451 (N_23451,N_22502,N_23036);
nand U23452 (N_23452,N_22938,N_22577);
xor U23453 (N_23453,N_23081,N_23049);
or U23454 (N_23454,N_22872,N_22520);
nor U23455 (N_23455,N_22642,N_23062);
and U23456 (N_23456,N_22698,N_23065);
nor U23457 (N_23457,N_22693,N_22617);
xnor U23458 (N_23458,N_22865,N_22531);
and U23459 (N_23459,N_22992,N_22870);
nor U23460 (N_23460,N_23088,N_22575);
and U23461 (N_23461,N_22566,N_23036);
nand U23462 (N_23462,N_23115,N_22911);
and U23463 (N_23463,N_22863,N_22884);
or U23464 (N_23464,N_23093,N_22837);
nand U23465 (N_23465,N_22901,N_22742);
nor U23466 (N_23466,N_22509,N_22919);
xor U23467 (N_23467,N_23117,N_22934);
or U23468 (N_23468,N_22943,N_22664);
xor U23469 (N_23469,N_22846,N_22593);
or U23470 (N_23470,N_22707,N_23018);
nand U23471 (N_23471,N_22582,N_22831);
or U23472 (N_23472,N_22669,N_22975);
nor U23473 (N_23473,N_22800,N_22815);
or U23474 (N_23474,N_23039,N_22674);
or U23475 (N_23475,N_23016,N_22987);
nor U23476 (N_23476,N_22699,N_22829);
and U23477 (N_23477,N_22634,N_22564);
nand U23478 (N_23478,N_22829,N_23044);
nor U23479 (N_23479,N_23079,N_22729);
xor U23480 (N_23480,N_22760,N_22960);
xor U23481 (N_23481,N_22538,N_22858);
or U23482 (N_23482,N_22616,N_22797);
nand U23483 (N_23483,N_23123,N_23078);
nor U23484 (N_23484,N_23060,N_23095);
xnor U23485 (N_23485,N_22968,N_22713);
nor U23486 (N_23486,N_22684,N_23019);
xnor U23487 (N_23487,N_22759,N_22800);
nand U23488 (N_23488,N_22702,N_23101);
and U23489 (N_23489,N_22780,N_22631);
or U23490 (N_23490,N_22987,N_22857);
nor U23491 (N_23491,N_22500,N_22546);
xor U23492 (N_23492,N_23001,N_22875);
xor U23493 (N_23493,N_23078,N_22658);
nand U23494 (N_23494,N_23053,N_23122);
or U23495 (N_23495,N_22606,N_22723);
or U23496 (N_23496,N_23019,N_23068);
nor U23497 (N_23497,N_22830,N_23066);
xnor U23498 (N_23498,N_22808,N_23106);
or U23499 (N_23499,N_22594,N_22598);
nor U23500 (N_23500,N_23019,N_22763);
or U23501 (N_23501,N_23034,N_22533);
or U23502 (N_23502,N_22688,N_22733);
nor U23503 (N_23503,N_23013,N_22622);
and U23504 (N_23504,N_22898,N_22956);
nor U23505 (N_23505,N_22745,N_23026);
nand U23506 (N_23506,N_23039,N_23052);
nand U23507 (N_23507,N_22553,N_23058);
and U23508 (N_23508,N_22848,N_23075);
nand U23509 (N_23509,N_22918,N_22788);
nand U23510 (N_23510,N_22649,N_22553);
xnor U23511 (N_23511,N_23089,N_23037);
or U23512 (N_23512,N_22931,N_22723);
and U23513 (N_23513,N_22986,N_22594);
or U23514 (N_23514,N_22596,N_23117);
or U23515 (N_23515,N_22617,N_22508);
nor U23516 (N_23516,N_22859,N_22534);
and U23517 (N_23517,N_22862,N_22505);
or U23518 (N_23518,N_22663,N_22603);
or U23519 (N_23519,N_22830,N_22941);
and U23520 (N_23520,N_22703,N_22975);
nor U23521 (N_23521,N_22738,N_22682);
and U23522 (N_23522,N_22759,N_22732);
xnor U23523 (N_23523,N_22579,N_22695);
and U23524 (N_23524,N_22842,N_22567);
nor U23525 (N_23525,N_22572,N_23050);
nand U23526 (N_23526,N_23092,N_22677);
nand U23527 (N_23527,N_22911,N_22808);
or U23528 (N_23528,N_22624,N_22972);
nand U23529 (N_23529,N_23002,N_22900);
nand U23530 (N_23530,N_22562,N_22852);
xor U23531 (N_23531,N_22568,N_23050);
and U23532 (N_23532,N_22823,N_23014);
or U23533 (N_23533,N_22788,N_22999);
nand U23534 (N_23534,N_22589,N_22588);
xor U23535 (N_23535,N_22979,N_22781);
xor U23536 (N_23536,N_22581,N_22698);
or U23537 (N_23537,N_22685,N_22872);
nor U23538 (N_23538,N_23026,N_23045);
and U23539 (N_23539,N_23046,N_23074);
nor U23540 (N_23540,N_22625,N_22991);
nand U23541 (N_23541,N_22678,N_22713);
nand U23542 (N_23542,N_22636,N_22870);
nand U23543 (N_23543,N_22803,N_22521);
nor U23544 (N_23544,N_22731,N_22938);
or U23545 (N_23545,N_22684,N_23029);
xnor U23546 (N_23546,N_23104,N_22786);
xnor U23547 (N_23547,N_22695,N_22525);
xor U23548 (N_23548,N_22589,N_22750);
nor U23549 (N_23549,N_22849,N_22822);
nand U23550 (N_23550,N_22530,N_22698);
nand U23551 (N_23551,N_22759,N_22880);
or U23552 (N_23552,N_22515,N_23071);
and U23553 (N_23553,N_22902,N_22613);
nand U23554 (N_23554,N_22561,N_22918);
nor U23555 (N_23555,N_23064,N_22513);
nand U23556 (N_23556,N_22943,N_22749);
and U23557 (N_23557,N_22542,N_22835);
or U23558 (N_23558,N_22938,N_22969);
xor U23559 (N_23559,N_22802,N_22850);
nand U23560 (N_23560,N_23080,N_22786);
xor U23561 (N_23561,N_22538,N_23025);
nor U23562 (N_23562,N_23119,N_23012);
or U23563 (N_23563,N_22980,N_22808);
and U23564 (N_23564,N_22578,N_22591);
or U23565 (N_23565,N_22636,N_22538);
xnor U23566 (N_23566,N_23054,N_22595);
nand U23567 (N_23567,N_22818,N_22675);
nor U23568 (N_23568,N_22526,N_22902);
and U23569 (N_23569,N_22956,N_23076);
xnor U23570 (N_23570,N_22916,N_23010);
xnor U23571 (N_23571,N_22966,N_22624);
or U23572 (N_23572,N_22659,N_22542);
nor U23573 (N_23573,N_22568,N_22879);
or U23574 (N_23574,N_23077,N_22770);
or U23575 (N_23575,N_22654,N_22671);
nor U23576 (N_23576,N_23110,N_22614);
nor U23577 (N_23577,N_23036,N_22974);
nor U23578 (N_23578,N_22727,N_22864);
nor U23579 (N_23579,N_22673,N_22768);
xnor U23580 (N_23580,N_22700,N_22950);
xor U23581 (N_23581,N_22710,N_22707);
nand U23582 (N_23582,N_22588,N_22662);
nand U23583 (N_23583,N_22647,N_22619);
and U23584 (N_23584,N_22868,N_23093);
xor U23585 (N_23585,N_23066,N_22757);
nand U23586 (N_23586,N_22934,N_22635);
xnor U23587 (N_23587,N_22554,N_22661);
or U23588 (N_23588,N_22659,N_22890);
and U23589 (N_23589,N_22598,N_22960);
and U23590 (N_23590,N_22675,N_22768);
and U23591 (N_23591,N_22786,N_22789);
or U23592 (N_23592,N_22918,N_22995);
nand U23593 (N_23593,N_22789,N_22839);
nor U23594 (N_23594,N_22724,N_22990);
nand U23595 (N_23595,N_23052,N_22799);
xnor U23596 (N_23596,N_22917,N_22642);
xnor U23597 (N_23597,N_23115,N_22985);
and U23598 (N_23598,N_22760,N_22504);
and U23599 (N_23599,N_22622,N_22886);
or U23600 (N_23600,N_23003,N_22948);
xor U23601 (N_23601,N_22548,N_22845);
nor U23602 (N_23602,N_22730,N_22907);
or U23603 (N_23603,N_22635,N_22748);
or U23604 (N_23604,N_22924,N_22691);
nor U23605 (N_23605,N_22916,N_22798);
and U23606 (N_23606,N_22727,N_23050);
and U23607 (N_23607,N_22857,N_23009);
or U23608 (N_23608,N_22790,N_22842);
or U23609 (N_23609,N_22985,N_23004);
nor U23610 (N_23610,N_22962,N_22633);
or U23611 (N_23611,N_22982,N_23024);
nor U23612 (N_23612,N_22875,N_22675);
nor U23613 (N_23613,N_22862,N_22811);
nor U23614 (N_23614,N_23035,N_22839);
nor U23615 (N_23615,N_22537,N_23094);
or U23616 (N_23616,N_23073,N_23007);
nand U23617 (N_23617,N_22653,N_22748);
xor U23618 (N_23618,N_22717,N_22800);
xnor U23619 (N_23619,N_22671,N_23084);
nor U23620 (N_23620,N_22730,N_22593);
nor U23621 (N_23621,N_23058,N_22780);
and U23622 (N_23622,N_22964,N_22635);
nand U23623 (N_23623,N_22798,N_23084);
xnor U23624 (N_23624,N_22755,N_22753);
nand U23625 (N_23625,N_23045,N_22989);
nor U23626 (N_23626,N_22606,N_23095);
and U23627 (N_23627,N_22558,N_22964);
and U23628 (N_23628,N_22970,N_22954);
and U23629 (N_23629,N_22883,N_23088);
nand U23630 (N_23630,N_23037,N_22677);
or U23631 (N_23631,N_22552,N_22691);
nor U23632 (N_23632,N_22536,N_22510);
or U23633 (N_23633,N_22573,N_22628);
nand U23634 (N_23634,N_22629,N_22916);
xnor U23635 (N_23635,N_23051,N_22808);
nand U23636 (N_23636,N_22508,N_23080);
and U23637 (N_23637,N_22537,N_22898);
or U23638 (N_23638,N_22885,N_22537);
and U23639 (N_23639,N_22752,N_23016);
xor U23640 (N_23640,N_22563,N_22568);
and U23641 (N_23641,N_23049,N_22518);
nand U23642 (N_23642,N_22972,N_22930);
xor U23643 (N_23643,N_22995,N_22901);
or U23644 (N_23644,N_23087,N_22810);
xor U23645 (N_23645,N_22574,N_22816);
and U23646 (N_23646,N_22729,N_22616);
xor U23647 (N_23647,N_22924,N_22693);
xnor U23648 (N_23648,N_22553,N_22699);
or U23649 (N_23649,N_22822,N_23102);
and U23650 (N_23650,N_23110,N_22794);
and U23651 (N_23651,N_23083,N_22526);
or U23652 (N_23652,N_22756,N_22988);
nor U23653 (N_23653,N_22825,N_22567);
nor U23654 (N_23654,N_23099,N_22659);
nor U23655 (N_23655,N_22545,N_22522);
and U23656 (N_23656,N_22889,N_22751);
nor U23657 (N_23657,N_22987,N_22559);
nand U23658 (N_23658,N_22915,N_22877);
or U23659 (N_23659,N_22530,N_22710);
nand U23660 (N_23660,N_23051,N_22818);
or U23661 (N_23661,N_22590,N_23031);
and U23662 (N_23662,N_22803,N_22990);
nor U23663 (N_23663,N_22894,N_22994);
nand U23664 (N_23664,N_22871,N_22831);
or U23665 (N_23665,N_22618,N_22764);
xnor U23666 (N_23666,N_22797,N_22985);
nand U23667 (N_23667,N_22795,N_22606);
nor U23668 (N_23668,N_22566,N_22890);
or U23669 (N_23669,N_22660,N_22978);
xor U23670 (N_23670,N_22669,N_22980);
nor U23671 (N_23671,N_22895,N_22804);
and U23672 (N_23672,N_22723,N_22534);
and U23673 (N_23673,N_22860,N_22859);
nand U23674 (N_23674,N_22797,N_23011);
xor U23675 (N_23675,N_22651,N_22977);
and U23676 (N_23676,N_22827,N_22758);
xnor U23677 (N_23677,N_22561,N_22653);
nor U23678 (N_23678,N_22848,N_22678);
nand U23679 (N_23679,N_22869,N_22648);
xnor U23680 (N_23680,N_23105,N_22741);
nor U23681 (N_23681,N_22574,N_23035);
nand U23682 (N_23682,N_22868,N_22691);
or U23683 (N_23683,N_22540,N_22653);
and U23684 (N_23684,N_22871,N_22954);
nor U23685 (N_23685,N_22530,N_22909);
nor U23686 (N_23686,N_22851,N_22672);
nand U23687 (N_23687,N_22578,N_22728);
nor U23688 (N_23688,N_22531,N_23080);
or U23689 (N_23689,N_22743,N_23120);
and U23690 (N_23690,N_22630,N_22869);
or U23691 (N_23691,N_22573,N_22760);
or U23692 (N_23692,N_22939,N_22896);
and U23693 (N_23693,N_22597,N_23040);
or U23694 (N_23694,N_22760,N_22863);
xnor U23695 (N_23695,N_22850,N_22848);
nor U23696 (N_23696,N_22928,N_22735);
nand U23697 (N_23697,N_22516,N_23080);
and U23698 (N_23698,N_22928,N_22846);
nand U23699 (N_23699,N_22901,N_22892);
or U23700 (N_23700,N_23038,N_22835);
and U23701 (N_23701,N_22598,N_22503);
and U23702 (N_23702,N_22698,N_22659);
nor U23703 (N_23703,N_22575,N_23083);
or U23704 (N_23704,N_22885,N_22674);
nand U23705 (N_23705,N_22684,N_22790);
and U23706 (N_23706,N_22536,N_22563);
and U23707 (N_23707,N_22689,N_22690);
or U23708 (N_23708,N_22595,N_22979);
and U23709 (N_23709,N_22567,N_22605);
or U23710 (N_23710,N_22923,N_23073);
or U23711 (N_23711,N_22747,N_22968);
and U23712 (N_23712,N_23106,N_23064);
or U23713 (N_23713,N_22948,N_22958);
xnor U23714 (N_23714,N_23006,N_23055);
and U23715 (N_23715,N_23069,N_22662);
or U23716 (N_23716,N_22659,N_22896);
nor U23717 (N_23717,N_23083,N_22696);
and U23718 (N_23718,N_22719,N_22893);
and U23719 (N_23719,N_22586,N_23119);
and U23720 (N_23720,N_22624,N_22823);
or U23721 (N_23721,N_22967,N_22560);
and U23722 (N_23722,N_22994,N_22647);
nand U23723 (N_23723,N_22503,N_22744);
and U23724 (N_23724,N_23098,N_22911);
or U23725 (N_23725,N_22759,N_23032);
nor U23726 (N_23726,N_22725,N_23056);
and U23727 (N_23727,N_22946,N_22684);
and U23728 (N_23728,N_23105,N_22784);
xnor U23729 (N_23729,N_22968,N_22564);
nand U23730 (N_23730,N_22668,N_22644);
nor U23731 (N_23731,N_23051,N_22964);
and U23732 (N_23732,N_22815,N_22509);
or U23733 (N_23733,N_22547,N_22772);
and U23734 (N_23734,N_23088,N_22521);
nand U23735 (N_23735,N_23061,N_22696);
xor U23736 (N_23736,N_23070,N_23080);
or U23737 (N_23737,N_22511,N_22935);
nor U23738 (N_23738,N_22659,N_23049);
nand U23739 (N_23739,N_22882,N_23121);
nor U23740 (N_23740,N_22738,N_23053);
or U23741 (N_23741,N_22842,N_22779);
nor U23742 (N_23742,N_22615,N_22980);
xnor U23743 (N_23743,N_22944,N_22769);
and U23744 (N_23744,N_22808,N_23105);
nor U23745 (N_23745,N_23014,N_22611);
xnor U23746 (N_23746,N_22793,N_22500);
or U23747 (N_23747,N_22520,N_22678);
or U23748 (N_23748,N_22679,N_22795);
or U23749 (N_23749,N_22589,N_22808);
nor U23750 (N_23750,N_23647,N_23172);
or U23751 (N_23751,N_23686,N_23415);
nand U23752 (N_23752,N_23641,N_23526);
nor U23753 (N_23753,N_23562,N_23365);
or U23754 (N_23754,N_23490,N_23561);
xor U23755 (N_23755,N_23195,N_23136);
xnor U23756 (N_23756,N_23705,N_23229);
nor U23757 (N_23757,N_23653,N_23461);
nand U23758 (N_23758,N_23338,N_23693);
and U23759 (N_23759,N_23629,N_23446);
and U23760 (N_23760,N_23720,N_23486);
and U23761 (N_23761,N_23580,N_23379);
nand U23762 (N_23762,N_23314,N_23531);
xor U23763 (N_23763,N_23740,N_23383);
nor U23764 (N_23764,N_23303,N_23423);
nand U23765 (N_23765,N_23492,N_23339);
or U23766 (N_23766,N_23679,N_23322);
or U23767 (N_23767,N_23616,N_23215);
and U23768 (N_23768,N_23578,N_23293);
or U23769 (N_23769,N_23373,N_23261);
or U23770 (N_23770,N_23455,N_23198);
or U23771 (N_23771,N_23161,N_23541);
and U23772 (N_23772,N_23714,N_23358);
and U23773 (N_23773,N_23405,N_23552);
and U23774 (N_23774,N_23672,N_23197);
and U23775 (N_23775,N_23267,N_23235);
nor U23776 (N_23776,N_23301,N_23256);
and U23777 (N_23777,N_23420,N_23570);
and U23778 (N_23778,N_23707,N_23619);
and U23779 (N_23779,N_23481,N_23724);
and U23780 (N_23780,N_23634,N_23620);
or U23781 (N_23781,N_23363,N_23436);
nand U23782 (N_23782,N_23696,N_23700);
and U23783 (N_23783,N_23290,N_23219);
xor U23784 (N_23784,N_23665,N_23512);
or U23785 (N_23785,N_23231,N_23376);
nor U23786 (N_23786,N_23668,N_23288);
or U23787 (N_23787,N_23252,N_23159);
nand U23788 (N_23788,N_23599,N_23522);
nor U23789 (N_23789,N_23637,N_23190);
xnor U23790 (N_23790,N_23142,N_23579);
nand U23791 (N_23791,N_23721,N_23263);
or U23792 (N_23792,N_23702,N_23581);
and U23793 (N_23793,N_23621,N_23277);
xor U23794 (N_23794,N_23281,N_23410);
and U23795 (N_23795,N_23251,N_23183);
or U23796 (N_23796,N_23408,N_23186);
nor U23797 (N_23797,N_23398,N_23594);
nor U23798 (N_23798,N_23321,N_23725);
and U23799 (N_23799,N_23704,N_23337);
or U23800 (N_23800,N_23294,N_23126);
and U23801 (N_23801,N_23335,N_23207);
nor U23802 (N_23802,N_23135,N_23203);
nor U23803 (N_23803,N_23155,N_23457);
nor U23804 (N_23804,N_23598,N_23151);
nand U23805 (N_23805,N_23140,N_23743);
nand U23806 (N_23806,N_23268,N_23600);
xor U23807 (N_23807,N_23566,N_23317);
nor U23808 (N_23808,N_23516,N_23176);
xor U23809 (N_23809,N_23305,N_23460);
xnor U23810 (N_23810,N_23242,N_23501);
and U23811 (N_23811,N_23445,N_23595);
and U23812 (N_23812,N_23432,N_23661);
nand U23813 (N_23813,N_23572,N_23617);
nand U23814 (N_23814,N_23153,N_23631);
xor U23815 (N_23815,N_23318,N_23507);
and U23816 (N_23816,N_23625,N_23417);
or U23817 (N_23817,N_23636,N_23593);
nand U23818 (N_23818,N_23144,N_23329);
nand U23819 (N_23819,N_23453,N_23476);
nor U23820 (N_23820,N_23264,N_23749);
nand U23821 (N_23821,N_23659,N_23208);
nor U23822 (N_23822,N_23241,N_23166);
xor U23823 (N_23823,N_23421,N_23418);
xnor U23824 (N_23824,N_23540,N_23657);
nor U23825 (N_23825,N_23138,N_23664);
nor U23826 (N_23826,N_23509,N_23643);
or U23827 (N_23827,N_23746,N_23291);
nor U23828 (N_23828,N_23255,N_23532);
nand U23829 (N_23829,N_23296,N_23736);
and U23830 (N_23830,N_23528,N_23710);
nor U23831 (N_23831,N_23385,N_23478);
nor U23832 (N_23832,N_23613,N_23554);
nand U23833 (N_23833,N_23442,N_23278);
or U23834 (N_23834,N_23504,N_23237);
nor U23835 (N_23835,N_23349,N_23244);
or U23836 (N_23836,N_23609,N_23745);
nand U23837 (N_23837,N_23544,N_23299);
xor U23838 (N_23838,N_23644,N_23205);
nand U23839 (N_23839,N_23431,N_23717);
nand U23840 (N_23840,N_23688,N_23530);
xnor U23841 (N_23841,N_23134,N_23345);
and U23842 (N_23842,N_23353,N_23539);
and U23843 (N_23843,N_23143,N_23196);
or U23844 (N_23844,N_23269,N_23677);
xnor U23845 (N_23845,N_23171,N_23556);
nand U23846 (N_23846,N_23611,N_23650);
nor U23847 (N_23847,N_23663,N_23535);
or U23848 (N_23848,N_23744,N_23259);
and U23849 (N_23849,N_23178,N_23475);
or U23850 (N_23850,N_23605,N_23226);
and U23851 (N_23851,N_23217,N_23536);
nand U23852 (N_23852,N_23282,N_23260);
xor U23853 (N_23853,N_23715,N_23179);
nand U23854 (N_23854,N_23346,N_23239);
nor U23855 (N_23855,N_23312,N_23316);
nand U23856 (N_23856,N_23549,N_23187);
and U23857 (N_23857,N_23440,N_23716);
xor U23858 (N_23858,N_23515,N_23382);
nand U23859 (N_23859,N_23697,N_23466);
and U23860 (N_23860,N_23300,N_23655);
nor U23861 (N_23861,N_23538,N_23499);
nor U23862 (N_23862,N_23563,N_23163);
nor U23863 (N_23863,N_23494,N_23271);
nand U23864 (N_23864,N_23343,N_23675);
nor U23865 (N_23865,N_23395,N_23451);
or U23866 (N_23866,N_23170,N_23520);
nor U23867 (N_23867,N_23748,N_23156);
and U23868 (N_23868,N_23206,N_23292);
nor U23869 (N_23869,N_23713,N_23742);
and U23870 (N_23870,N_23250,N_23689);
or U23871 (N_23871,N_23364,N_23220);
or U23872 (N_23872,N_23551,N_23510);
or U23873 (N_23873,N_23518,N_23607);
nand U23874 (N_23874,N_23564,N_23498);
xnor U23875 (N_23875,N_23414,N_23646);
xor U23876 (N_23876,N_23500,N_23154);
xor U23877 (N_23877,N_23633,N_23212);
xor U23878 (N_23878,N_23439,N_23334);
or U23879 (N_23879,N_23435,N_23351);
or U23880 (N_23880,N_23222,N_23680);
nand U23881 (N_23881,N_23149,N_23354);
or U23882 (N_23882,N_23331,N_23368);
xor U23883 (N_23883,N_23571,N_23690);
or U23884 (N_23884,N_23380,N_23673);
or U23885 (N_23885,N_23645,N_23200);
xor U23886 (N_23886,N_23181,N_23639);
nor U23887 (N_23887,N_23589,N_23437);
or U23888 (N_23888,N_23369,N_23622);
and U23889 (N_23889,N_23150,N_23430);
xnor U23890 (N_23890,N_23602,N_23488);
or U23891 (N_23891,N_23576,N_23547);
and U23892 (N_23892,N_23524,N_23590);
and U23893 (N_23893,N_23262,N_23586);
nor U23894 (N_23894,N_23464,N_23582);
nor U23895 (N_23895,N_23584,N_23550);
or U23896 (N_23896,N_23184,N_23158);
and U23897 (N_23897,N_23228,N_23670);
xnor U23898 (N_23898,N_23685,N_23273);
nand U23899 (N_23899,N_23517,N_23201);
xnor U23900 (N_23900,N_23592,N_23729);
or U23901 (N_23901,N_23402,N_23730);
or U23902 (N_23902,N_23708,N_23361);
nand U23903 (N_23903,N_23258,N_23392);
xor U23904 (N_23904,N_23422,N_23573);
nor U23905 (N_23905,N_23221,N_23627);
nor U23906 (N_23906,N_23546,N_23396);
and U23907 (N_23907,N_23375,N_23315);
and U23908 (N_23908,N_23447,N_23493);
xnor U23909 (N_23909,N_23505,N_23468);
or U23910 (N_23910,N_23474,N_23387);
or U23911 (N_23911,N_23608,N_23127);
and U23912 (N_23912,N_23238,N_23678);
xnor U23913 (N_23913,N_23378,N_23428);
nor U23914 (N_23914,N_23545,N_23254);
nor U23915 (N_23915,N_23284,N_23157);
and U23916 (N_23916,N_23132,N_23519);
or U23917 (N_23917,N_23674,N_23306);
nor U23918 (N_23918,N_23667,N_23719);
nand U23919 (N_23919,N_23372,N_23359);
and U23920 (N_23920,N_23413,N_23640);
xor U23921 (N_23921,N_23604,N_23472);
nor U23922 (N_23922,N_23406,N_23287);
nand U23923 (N_23923,N_23129,N_23601);
or U23924 (N_23924,N_23128,N_23747);
and U23925 (N_23925,N_23313,N_23443);
and U23926 (N_23926,N_23403,N_23211);
xor U23927 (N_23927,N_23167,N_23189);
and U23928 (N_23928,N_23374,N_23390);
or U23929 (N_23929,N_23448,N_23272);
and U23930 (N_23930,N_23147,N_23204);
nand U23931 (N_23931,N_23394,N_23233);
nand U23932 (N_23932,N_23703,N_23735);
and U23933 (N_23933,N_23706,N_23433);
and U23934 (N_23934,N_23738,N_23371);
or U23935 (N_23935,N_23558,N_23712);
nor U23936 (N_23936,N_23630,N_23388);
nor U23937 (N_23937,N_23304,N_23467);
nand U23938 (N_23938,N_23626,N_23444);
or U23939 (N_23939,N_23389,N_23537);
nand U23940 (N_23940,N_23514,N_23297);
xnor U23941 (N_23941,N_23656,N_23502);
or U23942 (N_23942,N_23691,N_23542);
nand U23943 (N_23943,N_23606,N_23367);
xnor U23944 (N_23944,N_23612,N_23245);
xnor U23945 (N_23945,N_23699,N_23357);
nor U23946 (N_23946,N_23458,N_23434);
nand U23947 (N_23947,N_23356,N_23569);
and U23948 (N_23948,N_23722,N_23618);
or U23949 (N_23949,N_23711,N_23588);
or U23950 (N_23950,N_23404,N_23401);
or U23951 (N_23951,N_23575,N_23477);
nand U23952 (N_23952,N_23734,N_23130);
and U23953 (N_23953,N_23479,N_23463);
and U23954 (N_23954,N_23429,N_23283);
or U23955 (N_23955,N_23249,N_23295);
nand U23956 (N_23956,N_23534,N_23642);
xor U23957 (N_23957,N_23279,N_23651);
nand U23958 (N_23958,N_23209,N_23587);
xnor U23959 (N_23959,N_23683,N_23169);
or U23960 (N_23960,N_23180,N_23511);
nor U23961 (N_23961,N_23459,N_23192);
xnor U23962 (N_23962,N_23286,N_23173);
or U23963 (N_23963,N_23559,N_23662);
nand U23964 (N_23964,N_23328,N_23366);
or U23965 (N_23965,N_23565,N_23230);
nor U23966 (N_23966,N_23324,N_23308);
or U23967 (N_23967,N_23302,N_23560);
xnor U23968 (N_23968,N_23342,N_23285);
nand U23969 (N_23969,N_23658,N_23289);
or U23970 (N_23970,N_23497,N_23182);
xor U23971 (N_23971,N_23265,N_23638);
nor U23972 (N_23972,N_23483,N_23596);
nand U23973 (N_23973,N_23568,N_23399);
nand U23974 (N_23974,N_23424,N_23553);
nand U23975 (N_23975,N_23449,N_23583);
nor U23976 (N_23976,N_23174,N_23320);
xor U23977 (N_23977,N_23216,N_23723);
nand U23978 (N_23978,N_23311,N_23350);
nor U23979 (N_23979,N_23164,N_23480);
nand U23980 (N_23980,N_23384,N_23411);
or U23981 (N_23981,N_23362,N_23125);
nand U23982 (N_23982,N_23452,N_23175);
or U23983 (N_23983,N_23393,N_23603);
nand U23984 (N_23984,N_23506,N_23733);
or U23985 (N_23985,N_23145,N_23543);
and U23986 (N_23986,N_23741,N_23257);
xor U23987 (N_23987,N_23628,N_23694);
or U23988 (N_23988,N_23332,N_23591);
xor U23989 (N_23989,N_23557,N_23682);
or U23990 (N_23990,N_23513,N_23521);
xor U23991 (N_23991,N_23266,N_23185);
xnor U23992 (N_23992,N_23165,N_23623);
nand U23993 (N_23993,N_23523,N_23326);
or U23994 (N_23994,N_23527,N_23577);
nor U23995 (N_23995,N_23236,N_23327);
xnor U23996 (N_23996,N_23397,N_23218);
and U23997 (N_23997,N_23309,N_23276);
or U23998 (N_23998,N_23223,N_23487);
and U23999 (N_23999,N_23333,N_23232);
nor U24000 (N_24000,N_23597,N_23652);
nor U24001 (N_24001,N_23137,N_23469);
nand U24002 (N_24002,N_23400,N_23495);
or U24003 (N_24003,N_23471,N_23344);
nor U24004 (N_24004,N_23274,N_23687);
or U24005 (N_24005,N_23348,N_23425);
nor U24006 (N_24006,N_23482,N_23162);
and U24007 (N_24007,N_23234,N_23146);
nor U24008 (N_24008,N_23191,N_23496);
nor U24009 (N_24009,N_23412,N_23298);
or U24010 (N_24010,N_23695,N_23484);
xnor U24011 (N_24011,N_23726,N_23352);
or U24012 (N_24012,N_23210,N_23407);
nand U24013 (N_24013,N_23709,N_23177);
nor U24014 (N_24014,N_23632,N_23671);
nor U24015 (N_24015,N_23489,N_23727);
or U24016 (N_24016,N_23275,N_23202);
xnor U24017 (N_24017,N_23227,N_23548);
and U24018 (N_24018,N_23585,N_23438);
or U24019 (N_24019,N_23319,N_23567);
xor U24020 (N_24020,N_23427,N_23491);
nor U24021 (N_24021,N_23199,N_23139);
xor U24022 (N_24022,N_23529,N_23193);
and U24023 (N_24023,N_23731,N_23648);
and U24024 (N_24024,N_23377,N_23336);
or U24025 (N_24025,N_23660,N_23610);
nor U24026 (N_24026,N_23214,N_23701);
and U24027 (N_24027,N_23409,N_23462);
nor U24028 (N_24028,N_23441,N_23370);
xnor U24029 (N_24029,N_23684,N_23450);
nor U24030 (N_24030,N_23225,N_23168);
nand U24031 (N_24031,N_23419,N_23485);
xor U24032 (N_24032,N_23624,N_23473);
and U24033 (N_24033,N_23681,N_23470);
nand U24034 (N_24034,N_23635,N_23307);
nor U24035 (N_24035,N_23692,N_23160);
nand U24036 (N_24036,N_23360,N_23728);
or U24037 (N_24037,N_23240,N_23654);
nand U24038 (N_24038,N_23533,N_23732);
xnor U24039 (N_24039,N_23247,N_23280);
nor U24040 (N_24040,N_23243,N_23391);
or U24041 (N_24041,N_23246,N_23426);
or U24042 (N_24042,N_23465,N_23270);
nor U24043 (N_24043,N_23340,N_23347);
or U24044 (N_24044,N_23386,N_23148);
or U24045 (N_24045,N_23341,N_23456);
and U24046 (N_24046,N_23381,N_23508);
and U24047 (N_24047,N_23614,N_23615);
nor U24048 (N_24048,N_23194,N_23739);
and U24049 (N_24049,N_23555,N_23355);
xnor U24050 (N_24050,N_23454,N_23669);
nor U24051 (N_24051,N_23310,N_23330);
and U24052 (N_24052,N_23248,N_23224);
or U24053 (N_24053,N_23503,N_23323);
nand U24054 (N_24054,N_23737,N_23676);
xnor U24055 (N_24055,N_23213,N_23525);
xor U24056 (N_24056,N_23325,N_23133);
nand U24057 (N_24057,N_23666,N_23416);
nor U24058 (N_24058,N_23152,N_23131);
nor U24059 (N_24059,N_23141,N_23698);
or U24060 (N_24060,N_23574,N_23718);
nor U24061 (N_24061,N_23649,N_23188);
xnor U24062 (N_24062,N_23253,N_23563);
nor U24063 (N_24063,N_23554,N_23249);
xnor U24064 (N_24064,N_23379,N_23361);
xor U24065 (N_24065,N_23347,N_23260);
nor U24066 (N_24066,N_23708,N_23384);
or U24067 (N_24067,N_23264,N_23340);
nor U24068 (N_24068,N_23676,N_23305);
nand U24069 (N_24069,N_23291,N_23487);
nor U24070 (N_24070,N_23182,N_23183);
and U24071 (N_24071,N_23210,N_23284);
and U24072 (N_24072,N_23205,N_23517);
or U24073 (N_24073,N_23678,N_23585);
nand U24074 (N_24074,N_23610,N_23574);
nor U24075 (N_24075,N_23469,N_23708);
xor U24076 (N_24076,N_23567,N_23219);
xnor U24077 (N_24077,N_23667,N_23704);
and U24078 (N_24078,N_23362,N_23622);
nor U24079 (N_24079,N_23490,N_23597);
nand U24080 (N_24080,N_23456,N_23403);
and U24081 (N_24081,N_23299,N_23619);
or U24082 (N_24082,N_23307,N_23455);
or U24083 (N_24083,N_23262,N_23588);
and U24084 (N_24084,N_23320,N_23688);
or U24085 (N_24085,N_23473,N_23617);
or U24086 (N_24086,N_23691,N_23686);
xor U24087 (N_24087,N_23281,N_23227);
nor U24088 (N_24088,N_23659,N_23289);
or U24089 (N_24089,N_23310,N_23237);
and U24090 (N_24090,N_23453,N_23734);
nor U24091 (N_24091,N_23392,N_23157);
xnor U24092 (N_24092,N_23327,N_23749);
xnor U24093 (N_24093,N_23167,N_23635);
and U24094 (N_24094,N_23540,N_23550);
nand U24095 (N_24095,N_23426,N_23305);
and U24096 (N_24096,N_23748,N_23633);
and U24097 (N_24097,N_23595,N_23709);
xor U24098 (N_24098,N_23506,N_23558);
xnor U24099 (N_24099,N_23425,N_23686);
or U24100 (N_24100,N_23568,N_23558);
xnor U24101 (N_24101,N_23614,N_23230);
and U24102 (N_24102,N_23727,N_23284);
and U24103 (N_24103,N_23489,N_23411);
nor U24104 (N_24104,N_23445,N_23398);
and U24105 (N_24105,N_23741,N_23408);
nor U24106 (N_24106,N_23483,N_23204);
or U24107 (N_24107,N_23723,N_23139);
nand U24108 (N_24108,N_23562,N_23578);
xnor U24109 (N_24109,N_23651,N_23440);
or U24110 (N_24110,N_23344,N_23542);
nor U24111 (N_24111,N_23404,N_23319);
and U24112 (N_24112,N_23428,N_23646);
xnor U24113 (N_24113,N_23329,N_23673);
and U24114 (N_24114,N_23720,N_23230);
nand U24115 (N_24115,N_23492,N_23572);
nor U24116 (N_24116,N_23680,N_23648);
xnor U24117 (N_24117,N_23314,N_23436);
or U24118 (N_24118,N_23696,N_23620);
nor U24119 (N_24119,N_23525,N_23528);
nor U24120 (N_24120,N_23225,N_23311);
or U24121 (N_24121,N_23477,N_23281);
xor U24122 (N_24122,N_23164,N_23394);
nand U24123 (N_24123,N_23642,N_23540);
and U24124 (N_24124,N_23502,N_23478);
or U24125 (N_24125,N_23234,N_23646);
or U24126 (N_24126,N_23178,N_23727);
xnor U24127 (N_24127,N_23334,N_23248);
xor U24128 (N_24128,N_23636,N_23434);
nor U24129 (N_24129,N_23457,N_23382);
nor U24130 (N_24130,N_23459,N_23159);
and U24131 (N_24131,N_23641,N_23134);
nor U24132 (N_24132,N_23276,N_23216);
nand U24133 (N_24133,N_23158,N_23355);
and U24134 (N_24134,N_23277,N_23465);
and U24135 (N_24135,N_23628,N_23370);
or U24136 (N_24136,N_23162,N_23487);
xnor U24137 (N_24137,N_23722,N_23685);
xor U24138 (N_24138,N_23435,N_23577);
and U24139 (N_24139,N_23565,N_23737);
or U24140 (N_24140,N_23192,N_23196);
or U24141 (N_24141,N_23387,N_23614);
or U24142 (N_24142,N_23222,N_23733);
or U24143 (N_24143,N_23133,N_23506);
or U24144 (N_24144,N_23262,N_23238);
nor U24145 (N_24145,N_23173,N_23394);
and U24146 (N_24146,N_23475,N_23163);
nand U24147 (N_24147,N_23443,N_23450);
xnor U24148 (N_24148,N_23665,N_23443);
or U24149 (N_24149,N_23429,N_23225);
nor U24150 (N_24150,N_23644,N_23343);
and U24151 (N_24151,N_23437,N_23701);
xor U24152 (N_24152,N_23608,N_23376);
and U24153 (N_24153,N_23218,N_23181);
nor U24154 (N_24154,N_23496,N_23611);
nor U24155 (N_24155,N_23595,N_23379);
nand U24156 (N_24156,N_23394,N_23613);
or U24157 (N_24157,N_23724,N_23406);
and U24158 (N_24158,N_23130,N_23412);
or U24159 (N_24159,N_23507,N_23727);
nor U24160 (N_24160,N_23439,N_23742);
or U24161 (N_24161,N_23160,N_23441);
nor U24162 (N_24162,N_23178,N_23585);
nand U24163 (N_24163,N_23648,N_23478);
nand U24164 (N_24164,N_23166,N_23571);
xor U24165 (N_24165,N_23446,N_23172);
xor U24166 (N_24166,N_23455,N_23746);
or U24167 (N_24167,N_23422,N_23146);
and U24168 (N_24168,N_23304,N_23318);
or U24169 (N_24169,N_23663,N_23361);
or U24170 (N_24170,N_23393,N_23143);
nand U24171 (N_24171,N_23299,N_23559);
and U24172 (N_24172,N_23468,N_23663);
or U24173 (N_24173,N_23142,N_23648);
xnor U24174 (N_24174,N_23266,N_23662);
or U24175 (N_24175,N_23597,N_23409);
and U24176 (N_24176,N_23494,N_23136);
xnor U24177 (N_24177,N_23464,N_23730);
or U24178 (N_24178,N_23333,N_23362);
and U24179 (N_24179,N_23455,N_23142);
and U24180 (N_24180,N_23511,N_23616);
xnor U24181 (N_24181,N_23327,N_23571);
xnor U24182 (N_24182,N_23525,N_23392);
nor U24183 (N_24183,N_23291,N_23234);
or U24184 (N_24184,N_23165,N_23257);
xor U24185 (N_24185,N_23134,N_23250);
and U24186 (N_24186,N_23645,N_23175);
nor U24187 (N_24187,N_23600,N_23504);
xnor U24188 (N_24188,N_23315,N_23552);
xor U24189 (N_24189,N_23169,N_23220);
nor U24190 (N_24190,N_23682,N_23651);
and U24191 (N_24191,N_23384,N_23265);
and U24192 (N_24192,N_23268,N_23239);
nor U24193 (N_24193,N_23716,N_23242);
xnor U24194 (N_24194,N_23489,N_23507);
xor U24195 (N_24195,N_23346,N_23402);
xnor U24196 (N_24196,N_23543,N_23572);
nand U24197 (N_24197,N_23557,N_23419);
or U24198 (N_24198,N_23593,N_23655);
or U24199 (N_24199,N_23335,N_23156);
xnor U24200 (N_24200,N_23354,N_23231);
or U24201 (N_24201,N_23262,N_23737);
or U24202 (N_24202,N_23313,N_23647);
nor U24203 (N_24203,N_23242,N_23502);
nor U24204 (N_24204,N_23485,N_23660);
nor U24205 (N_24205,N_23236,N_23160);
or U24206 (N_24206,N_23565,N_23744);
and U24207 (N_24207,N_23688,N_23494);
nor U24208 (N_24208,N_23431,N_23176);
and U24209 (N_24209,N_23624,N_23358);
nand U24210 (N_24210,N_23264,N_23514);
or U24211 (N_24211,N_23410,N_23674);
or U24212 (N_24212,N_23684,N_23447);
or U24213 (N_24213,N_23567,N_23198);
and U24214 (N_24214,N_23136,N_23478);
nand U24215 (N_24215,N_23455,N_23469);
nor U24216 (N_24216,N_23137,N_23564);
xor U24217 (N_24217,N_23561,N_23585);
xnor U24218 (N_24218,N_23632,N_23144);
xnor U24219 (N_24219,N_23214,N_23306);
nand U24220 (N_24220,N_23213,N_23542);
nand U24221 (N_24221,N_23692,N_23717);
nand U24222 (N_24222,N_23357,N_23136);
xor U24223 (N_24223,N_23445,N_23482);
xnor U24224 (N_24224,N_23523,N_23217);
nand U24225 (N_24225,N_23152,N_23199);
nand U24226 (N_24226,N_23535,N_23706);
xor U24227 (N_24227,N_23156,N_23696);
or U24228 (N_24228,N_23661,N_23181);
nor U24229 (N_24229,N_23661,N_23255);
or U24230 (N_24230,N_23169,N_23268);
nor U24231 (N_24231,N_23513,N_23680);
and U24232 (N_24232,N_23137,N_23607);
xnor U24233 (N_24233,N_23210,N_23358);
nor U24234 (N_24234,N_23481,N_23148);
nor U24235 (N_24235,N_23215,N_23163);
nor U24236 (N_24236,N_23665,N_23208);
and U24237 (N_24237,N_23190,N_23154);
nand U24238 (N_24238,N_23736,N_23272);
xor U24239 (N_24239,N_23310,N_23295);
or U24240 (N_24240,N_23518,N_23723);
or U24241 (N_24241,N_23392,N_23343);
and U24242 (N_24242,N_23707,N_23221);
nor U24243 (N_24243,N_23182,N_23266);
xnor U24244 (N_24244,N_23279,N_23557);
xor U24245 (N_24245,N_23745,N_23410);
nand U24246 (N_24246,N_23663,N_23526);
or U24247 (N_24247,N_23333,N_23159);
nand U24248 (N_24248,N_23559,N_23212);
nand U24249 (N_24249,N_23433,N_23587);
or U24250 (N_24250,N_23240,N_23685);
nor U24251 (N_24251,N_23632,N_23173);
nor U24252 (N_24252,N_23382,N_23623);
and U24253 (N_24253,N_23601,N_23525);
or U24254 (N_24254,N_23738,N_23209);
and U24255 (N_24255,N_23568,N_23220);
xnor U24256 (N_24256,N_23451,N_23704);
xnor U24257 (N_24257,N_23200,N_23705);
nand U24258 (N_24258,N_23194,N_23492);
nand U24259 (N_24259,N_23287,N_23701);
nor U24260 (N_24260,N_23566,N_23293);
xnor U24261 (N_24261,N_23179,N_23523);
xnor U24262 (N_24262,N_23595,N_23186);
xor U24263 (N_24263,N_23552,N_23157);
xor U24264 (N_24264,N_23317,N_23707);
xor U24265 (N_24265,N_23202,N_23152);
or U24266 (N_24266,N_23307,N_23294);
nand U24267 (N_24267,N_23147,N_23555);
nand U24268 (N_24268,N_23709,N_23454);
or U24269 (N_24269,N_23685,N_23547);
nor U24270 (N_24270,N_23147,N_23492);
xor U24271 (N_24271,N_23211,N_23729);
or U24272 (N_24272,N_23514,N_23459);
or U24273 (N_24273,N_23649,N_23701);
nand U24274 (N_24274,N_23148,N_23172);
nor U24275 (N_24275,N_23287,N_23266);
nor U24276 (N_24276,N_23154,N_23558);
and U24277 (N_24277,N_23653,N_23503);
nand U24278 (N_24278,N_23263,N_23661);
and U24279 (N_24279,N_23614,N_23723);
nor U24280 (N_24280,N_23442,N_23308);
xnor U24281 (N_24281,N_23724,N_23264);
nand U24282 (N_24282,N_23571,N_23184);
nand U24283 (N_24283,N_23690,N_23487);
and U24284 (N_24284,N_23221,N_23403);
nand U24285 (N_24285,N_23274,N_23513);
or U24286 (N_24286,N_23363,N_23642);
and U24287 (N_24287,N_23285,N_23593);
or U24288 (N_24288,N_23477,N_23232);
nor U24289 (N_24289,N_23604,N_23293);
xor U24290 (N_24290,N_23350,N_23405);
nor U24291 (N_24291,N_23719,N_23505);
and U24292 (N_24292,N_23550,N_23374);
nand U24293 (N_24293,N_23638,N_23465);
and U24294 (N_24294,N_23665,N_23555);
and U24295 (N_24295,N_23735,N_23188);
nor U24296 (N_24296,N_23592,N_23323);
and U24297 (N_24297,N_23224,N_23367);
nand U24298 (N_24298,N_23305,N_23386);
nand U24299 (N_24299,N_23665,N_23294);
nor U24300 (N_24300,N_23328,N_23636);
xor U24301 (N_24301,N_23529,N_23504);
and U24302 (N_24302,N_23177,N_23349);
nor U24303 (N_24303,N_23575,N_23218);
or U24304 (N_24304,N_23459,N_23156);
nor U24305 (N_24305,N_23242,N_23361);
xor U24306 (N_24306,N_23302,N_23265);
xor U24307 (N_24307,N_23538,N_23510);
and U24308 (N_24308,N_23413,N_23155);
and U24309 (N_24309,N_23708,N_23156);
nor U24310 (N_24310,N_23553,N_23475);
xnor U24311 (N_24311,N_23138,N_23349);
or U24312 (N_24312,N_23615,N_23486);
nand U24313 (N_24313,N_23389,N_23168);
nand U24314 (N_24314,N_23189,N_23130);
or U24315 (N_24315,N_23678,N_23414);
nand U24316 (N_24316,N_23384,N_23749);
nor U24317 (N_24317,N_23642,N_23445);
nor U24318 (N_24318,N_23162,N_23313);
nand U24319 (N_24319,N_23408,N_23516);
or U24320 (N_24320,N_23398,N_23726);
or U24321 (N_24321,N_23688,N_23336);
and U24322 (N_24322,N_23384,N_23608);
and U24323 (N_24323,N_23131,N_23243);
nor U24324 (N_24324,N_23689,N_23261);
xnor U24325 (N_24325,N_23234,N_23664);
nand U24326 (N_24326,N_23468,N_23521);
nand U24327 (N_24327,N_23392,N_23247);
and U24328 (N_24328,N_23230,N_23746);
xnor U24329 (N_24329,N_23415,N_23253);
and U24330 (N_24330,N_23633,N_23458);
xnor U24331 (N_24331,N_23311,N_23599);
and U24332 (N_24332,N_23446,N_23609);
xor U24333 (N_24333,N_23212,N_23734);
nor U24334 (N_24334,N_23127,N_23168);
xor U24335 (N_24335,N_23268,N_23458);
or U24336 (N_24336,N_23177,N_23389);
xor U24337 (N_24337,N_23687,N_23507);
nor U24338 (N_24338,N_23386,N_23447);
or U24339 (N_24339,N_23487,N_23692);
and U24340 (N_24340,N_23654,N_23360);
or U24341 (N_24341,N_23331,N_23624);
nor U24342 (N_24342,N_23444,N_23174);
nand U24343 (N_24343,N_23293,N_23345);
and U24344 (N_24344,N_23647,N_23250);
nand U24345 (N_24345,N_23399,N_23498);
nor U24346 (N_24346,N_23260,N_23187);
xnor U24347 (N_24347,N_23310,N_23338);
nand U24348 (N_24348,N_23230,N_23434);
or U24349 (N_24349,N_23268,N_23412);
nor U24350 (N_24350,N_23652,N_23224);
or U24351 (N_24351,N_23468,N_23605);
nand U24352 (N_24352,N_23744,N_23334);
nor U24353 (N_24353,N_23293,N_23384);
nor U24354 (N_24354,N_23685,N_23283);
nand U24355 (N_24355,N_23616,N_23561);
xor U24356 (N_24356,N_23459,N_23401);
or U24357 (N_24357,N_23464,N_23338);
nand U24358 (N_24358,N_23353,N_23330);
and U24359 (N_24359,N_23408,N_23503);
nor U24360 (N_24360,N_23263,N_23424);
or U24361 (N_24361,N_23600,N_23585);
nand U24362 (N_24362,N_23251,N_23695);
nand U24363 (N_24363,N_23326,N_23312);
and U24364 (N_24364,N_23609,N_23393);
xnor U24365 (N_24365,N_23233,N_23189);
and U24366 (N_24366,N_23471,N_23549);
nor U24367 (N_24367,N_23218,N_23382);
and U24368 (N_24368,N_23430,N_23319);
nor U24369 (N_24369,N_23390,N_23519);
xor U24370 (N_24370,N_23303,N_23377);
and U24371 (N_24371,N_23343,N_23664);
xnor U24372 (N_24372,N_23229,N_23402);
nor U24373 (N_24373,N_23380,N_23695);
and U24374 (N_24374,N_23298,N_23503);
or U24375 (N_24375,N_23877,N_24315);
or U24376 (N_24376,N_24141,N_24271);
and U24377 (N_24377,N_23769,N_24331);
or U24378 (N_24378,N_24082,N_24263);
nand U24379 (N_24379,N_23751,N_23894);
nand U24380 (N_24380,N_23750,N_24325);
or U24381 (N_24381,N_24114,N_23910);
nor U24382 (N_24382,N_24200,N_23757);
xnor U24383 (N_24383,N_23808,N_23830);
and U24384 (N_24384,N_23921,N_24094);
and U24385 (N_24385,N_24179,N_23856);
or U24386 (N_24386,N_24195,N_24298);
nand U24387 (N_24387,N_24065,N_23837);
nor U24388 (N_24388,N_24233,N_24256);
and U24389 (N_24389,N_24085,N_24228);
xnor U24390 (N_24390,N_23949,N_24300);
nor U24391 (N_24391,N_23860,N_24064);
or U24392 (N_24392,N_24088,N_24342);
nand U24393 (N_24393,N_23807,N_24178);
nand U24394 (N_24394,N_24235,N_23780);
nand U24395 (N_24395,N_24329,N_23899);
or U24396 (N_24396,N_24108,N_24214);
nand U24397 (N_24397,N_23785,N_24186);
xor U24398 (N_24398,N_23835,N_24283);
nor U24399 (N_24399,N_23886,N_23915);
nand U24400 (N_24400,N_23933,N_24265);
nand U24401 (N_24401,N_24270,N_24297);
or U24402 (N_24402,N_24275,N_23789);
nand U24403 (N_24403,N_23799,N_23811);
and U24404 (N_24404,N_24241,N_24160);
or U24405 (N_24405,N_23754,N_24115);
or U24406 (N_24406,N_23779,N_23756);
nand U24407 (N_24407,N_23936,N_24007);
xnor U24408 (N_24408,N_24351,N_23991);
and U24409 (N_24409,N_23794,N_24251);
nor U24410 (N_24410,N_23996,N_24166);
and U24411 (N_24411,N_23889,N_24272);
nand U24412 (N_24412,N_23904,N_24148);
nand U24413 (N_24413,N_23952,N_24238);
nor U24414 (N_24414,N_24062,N_24180);
or U24415 (N_24415,N_23842,N_24185);
xor U24416 (N_24416,N_24015,N_23943);
nand U24417 (N_24417,N_24360,N_23917);
nand U24418 (N_24418,N_24028,N_23988);
nor U24419 (N_24419,N_24110,N_24106);
nor U24420 (N_24420,N_24116,N_23844);
xnor U24421 (N_24421,N_24054,N_23839);
nand U24422 (N_24422,N_24107,N_24137);
or U24423 (N_24423,N_24039,N_24059);
nand U24424 (N_24424,N_24125,N_23876);
nand U24425 (N_24425,N_23895,N_24244);
and U24426 (N_24426,N_24104,N_24146);
and U24427 (N_24427,N_24018,N_23793);
and U24428 (N_24428,N_24058,N_24132);
or U24429 (N_24429,N_23864,N_24305);
or U24430 (N_24430,N_24339,N_24068);
nand U24431 (N_24431,N_24227,N_23992);
and U24432 (N_24432,N_23822,N_24196);
xnor U24433 (N_24433,N_23908,N_23901);
xnor U24434 (N_24434,N_24136,N_24012);
nor U24435 (N_24435,N_24348,N_24359);
xnor U24436 (N_24436,N_23800,N_24143);
nand U24437 (N_24437,N_24316,N_23932);
xor U24438 (N_24438,N_24176,N_24181);
xor U24439 (N_24439,N_23871,N_23848);
or U24440 (N_24440,N_23846,N_24129);
and U24441 (N_24441,N_23783,N_24296);
or U24442 (N_24442,N_24057,N_24282);
nor U24443 (N_24443,N_24310,N_24205);
nor U24444 (N_24444,N_23859,N_24017);
xor U24445 (N_24445,N_23953,N_24060);
xnor U24446 (N_24446,N_24211,N_23858);
nor U24447 (N_24447,N_24063,N_24051);
xor U24448 (N_24448,N_24152,N_24303);
and U24449 (N_24449,N_24119,N_23818);
or U24450 (N_24450,N_24313,N_23984);
nand U24451 (N_24451,N_24358,N_24027);
nand U24452 (N_24452,N_24309,N_24191);
or U24453 (N_24453,N_23972,N_24301);
nor U24454 (N_24454,N_24144,N_24229);
nand U24455 (N_24455,N_23878,N_23752);
xor U24456 (N_24456,N_24264,N_23964);
and U24457 (N_24457,N_24187,N_23965);
nand U24458 (N_24458,N_23887,N_24083);
nor U24459 (N_24459,N_23993,N_24019);
xnor U24460 (N_24460,N_24239,N_24101);
nor U24461 (N_24461,N_23814,N_24081);
or U24462 (N_24462,N_24162,N_23890);
nand U24463 (N_24463,N_24212,N_23888);
xor U24464 (N_24464,N_24291,N_23817);
and U24465 (N_24465,N_24193,N_24292);
nor U24466 (N_24466,N_24145,N_24092);
nand U24467 (N_24467,N_24373,N_24131);
nor U24468 (N_24468,N_23884,N_24221);
xor U24469 (N_24469,N_23841,N_24338);
or U24470 (N_24470,N_23960,N_23782);
nand U24471 (N_24471,N_24231,N_24258);
and U24472 (N_24472,N_24167,N_24075);
or U24473 (N_24473,N_24128,N_24078);
or U24474 (N_24474,N_24069,N_24124);
or U24475 (N_24475,N_23771,N_23914);
xnor U24476 (N_24476,N_23853,N_23806);
nand U24477 (N_24477,N_24267,N_24295);
or U24478 (N_24478,N_24154,N_24142);
and U24479 (N_24479,N_23998,N_24366);
or U24480 (N_24480,N_23913,N_23903);
and U24481 (N_24481,N_23919,N_24175);
xor U24482 (N_24482,N_23755,N_24053);
nand U24483 (N_24483,N_24090,N_24159);
or U24484 (N_24484,N_24209,N_23843);
nor U24485 (N_24485,N_24259,N_24333);
nor U24486 (N_24486,N_24335,N_23893);
and U24487 (N_24487,N_23790,N_24287);
nand U24488 (N_24488,N_23766,N_24035);
xor U24489 (N_24489,N_24367,N_24198);
and U24490 (N_24490,N_24025,N_24147);
and U24491 (N_24491,N_23954,N_24080);
nor U24492 (N_24492,N_24197,N_24319);
and U24493 (N_24493,N_23999,N_23906);
xnor U24494 (N_24494,N_24207,N_24153);
or U24495 (N_24495,N_23924,N_24280);
nor U24496 (N_24496,N_24356,N_23868);
and U24497 (N_24497,N_23824,N_24236);
xor U24498 (N_24498,N_24232,N_23941);
or U24499 (N_24499,N_24248,N_23963);
nand U24500 (N_24500,N_24243,N_23946);
and U24501 (N_24501,N_24347,N_24361);
xnor U24502 (N_24502,N_23770,N_23945);
nand U24503 (N_24503,N_23840,N_24311);
xor U24504 (N_24504,N_24150,N_23944);
nor U24505 (N_24505,N_24262,N_24001);
or U24506 (N_24506,N_23865,N_24317);
xor U24507 (N_24507,N_24074,N_23762);
nor U24508 (N_24508,N_24014,N_23997);
nor U24509 (N_24509,N_23761,N_23776);
xor U24510 (N_24510,N_23951,N_23786);
nor U24511 (N_24511,N_24169,N_23845);
nand U24512 (N_24512,N_24052,N_24293);
nor U24513 (N_24513,N_24066,N_24004);
and U24514 (N_24514,N_24322,N_24032);
xnor U24515 (N_24515,N_24071,N_24257);
xor U24516 (N_24516,N_24318,N_24255);
xor U24517 (N_24517,N_23855,N_24173);
and U24518 (N_24518,N_23760,N_24284);
nand U24519 (N_24519,N_23816,N_24008);
xnor U24520 (N_24520,N_23851,N_23950);
and U24521 (N_24521,N_24299,N_24246);
nor U24522 (N_24522,N_24113,N_24208);
and U24523 (N_24523,N_24218,N_23819);
nand U24524 (N_24524,N_24345,N_23956);
nand U24525 (N_24525,N_24023,N_24149);
xnor U24526 (N_24526,N_23881,N_23891);
xor U24527 (N_24527,N_23986,N_24364);
nor U24528 (N_24528,N_24033,N_23938);
nand U24529 (N_24529,N_24121,N_23882);
and U24530 (N_24530,N_24135,N_23907);
xor U24531 (N_24531,N_23923,N_24273);
nor U24532 (N_24532,N_24072,N_23929);
and U24533 (N_24533,N_24006,N_24168);
nor U24534 (N_24534,N_23897,N_24111);
nor U24535 (N_24535,N_24031,N_23764);
and U24536 (N_24536,N_23788,N_24084);
or U24537 (N_24537,N_23866,N_24230);
and U24538 (N_24538,N_24163,N_24034);
xor U24539 (N_24539,N_24127,N_24079);
or U24540 (N_24540,N_23940,N_23832);
nor U24541 (N_24541,N_24130,N_24048);
xor U24542 (N_24542,N_24278,N_24118);
and U24543 (N_24543,N_24013,N_24038);
nand U24544 (N_24544,N_23812,N_24030);
or U24545 (N_24545,N_23980,N_24242);
nand U24546 (N_24546,N_23815,N_23928);
or U24547 (N_24547,N_24206,N_24139);
nand U24548 (N_24548,N_24247,N_24174);
nand U24549 (N_24549,N_24155,N_24097);
nand U24550 (N_24550,N_23968,N_24047);
or U24551 (N_24551,N_23753,N_23784);
xnor U24552 (N_24552,N_24372,N_23867);
and U24553 (N_24553,N_24215,N_24281);
nand U24554 (N_24554,N_24192,N_23834);
xor U24555 (N_24555,N_24040,N_24126);
nand U24556 (N_24556,N_23765,N_23905);
xor U24557 (N_24557,N_24353,N_24341);
and U24558 (N_24558,N_24334,N_24354);
and U24559 (N_24559,N_24164,N_24240);
nand U24560 (N_24560,N_24357,N_23979);
or U24561 (N_24561,N_24049,N_23879);
and U24562 (N_24562,N_23970,N_24201);
and U24563 (N_24563,N_24067,N_24182);
xor U24564 (N_24564,N_24224,N_24105);
nor U24565 (N_24565,N_23983,N_23971);
nor U24566 (N_24566,N_23768,N_24276);
xor U24567 (N_24567,N_23778,N_24061);
nor U24568 (N_24568,N_23829,N_23920);
nor U24569 (N_24569,N_23838,N_24171);
or U24570 (N_24570,N_24268,N_24157);
nand U24571 (N_24571,N_24330,N_24210);
or U24572 (N_24572,N_23777,N_23759);
xor U24573 (N_24573,N_24252,N_24253);
nand U24574 (N_24574,N_24024,N_24009);
nand U24575 (N_24575,N_24266,N_24103);
xor U24576 (N_24576,N_24044,N_23987);
nand U24577 (N_24577,N_23826,N_23792);
xnor U24578 (N_24578,N_23820,N_23927);
xnor U24579 (N_24579,N_23930,N_24374);
nand U24580 (N_24580,N_24288,N_24093);
or U24581 (N_24581,N_24037,N_24188);
xor U24582 (N_24582,N_24323,N_23973);
or U24583 (N_24583,N_24056,N_24355);
xnor U24584 (N_24584,N_23763,N_24086);
xnor U24585 (N_24585,N_24324,N_23836);
nand U24586 (N_24586,N_24223,N_24099);
or U24587 (N_24587,N_23828,N_24260);
or U24588 (N_24588,N_23801,N_24026);
nor U24589 (N_24589,N_23821,N_24011);
and U24590 (N_24590,N_24219,N_24226);
nor U24591 (N_24591,N_23911,N_24087);
and U24592 (N_24592,N_24327,N_24100);
or U24593 (N_24593,N_23798,N_23898);
or U24594 (N_24594,N_23847,N_23863);
nand U24595 (N_24595,N_24350,N_24172);
or U24596 (N_24596,N_24320,N_24363);
nor U24597 (N_24597,N_23797,N_24368);
nand U24598 (N_24598,N_24213,N_23978);
or U24599 (N_24599,N_24203,N_24000);
xor U24600 (N_24600,N_23925,N_23900);
or U24601 (N_24601,N_24204,N_24123);
nand U24602 (N_24602,N_24274,N_24286);
and U24603 (N_24603,N_23931,N_23975);
or U24604 (N_24604,N_23995,N_23775);
nand U24605 (N_24605,N_23880,N_23869);
nand U24606 (N_24606,N_23922,N_23795);
nor U24607 (N_24607,N_24234,N_24189);
nor U24608 (N_24608,N_23981,N_24220);
xnor U24609 (N_24609,N_24005,N_24073);
nand U24610 (N_24610,N_23861,N_23967);
and U24611 (N_24611,N_23976,N_24183);
and U24612 (N_24612,N_23854,N_23787);
and U24613 (N_24613,N_24290,N_24308);
nand U24614 (N_24614,N_23883,N_24098);
nand U24615 (N_24615,N_24370,N_23977);
and U24616 (N_24616,N_23962,N_24254);
nor U24617 (N_24617,N_24307,N_24042);
nor U24618 (N_24618,N_24285,N_24328);
xnor U24619 (N_24619,N_23809,N_24041);
nor U24620 (N_24620,N_23875,N_23773);
and U24621 (N_24621,N_23994,N_24277);
nand U24622 (N_24622,N_23805,N_24091);
or U24623 (N_24623,N_23813,N_23985);
or U24624 (N_24624,N_24020,N_23850);
and U24625 (N_24625,N_24055,N_24250);
and U24626 (N_24626,N_23781,N_23912);
nand U24627 (N_24627,N_24177,N_24036);
nand U24628 (N_24628,N_24002,N_24352);
and U24629 (N_24629,N_23833,N_24337);
and U24630 (N_24630,N_23937,N_23852);
xnor U24631 (N_24631,N_24120,N_23947);
xor U24632 (N_24632,N_24237,N_24222);
nor U24633 (N_24633,N_24109,N_23955);
or U24634 (N_24634,N_23827,N_23873);
nand U24635 (N_24635,N_23892,N_24321);
nand U24636 (N_24636,N_23935,N_24261);
nand U24637 (N_24637,N_24158,N_24371);
or U24638 (N_24638,N_24362,N_23948);
xor U24639 (N_24639,N_23942,N_23823);
or U24640 (N_24640,N_24096,N_23989);
or U24641 (N_24641,N_23831,N_24312);
nor U24642 (N_24642,N_24134,N_23969);
nand U24643 (N_24643,N_24249,N_24245);
or U24644 (N_24644,N_24202,N_24022);
or U24645 (N_24645,N_24184,N_24343);
and U24646 (N_24646,N_24340,N_24151);
and U24647 (N_24647,N_24046,N_24170);
or U24648 (N_24648,N_23909,N_24190);
nand U24649 (N_24649,N_23803,N_24076);
nor U24650 (N_24650,N_23885,N_23774);
nor U24651 (N_24651,N_24365,N_23966);
xor U24652 (N_24652,N_24156,N_24095);
nor U24653 (N_24653,N_23961,N_24029);
or U24654 (N_24654,N_24043,N_23974);
xnor U24655 (N_24655,N_24138,N_24336);
nor U24656 (N_24656,N_24216,N_24344);
xor U24657 (N_24657,N_24117,N_24349);
nor U24658 (N_24658,N_24122,N_23804);
nand U24659 (N_24659,N_23870,N_24102);
xor U24660 (N_24660,N_24050,N_23791);
nand U24661 (N_24661,N_23902,N_24199);
nand U24662 (N_24662,N_24294,N_24021);
nor U24663 (N_24663,N_24326,N_24225);
and U24664 (N_24664,N_24217,N_24112);
and U24665 (N_24665,N_24161,N_24314);
and U24666 (N_24666,N_23959,N_23862);
nor U24667 (N_24667,N_24194,N_24165);
or U24668 (N_24668,N_24045,N_23918);
or U24669 (N_24669,N_23758,N_24070);
xor U24670 (N_24670,N_23958,N_24306);
and U24671 (N_24671,N_24003,N_23796);
and U24672 (N_24672,N_24279,N_24077);
nor U24673 (N_24673,N_24016,N_23849);
nand U24674 (N_24674,N_24289,N_24133);
nand U24675 (N_24675,N_23926,N_23939);
or U24676 (N_24676,N_23772,N_24332);
nand U24677 (N_24677,N_23767,N_24346);
and U24678 (N_24678,N_24369,N_24089);
nand U24679 (N_24679,N_24304,N_24140);
nor U24680 (N_24680,N_23916,N_23957);
or U24681 (N_24681,N_23872,N_23810);
and U24682 (N_24682,N_23874,N_24010);
and U24683 (N_24683,N_23990,N_23896);
nor U24684 (N_24684,N_23802,N_24269);
xnor U24685 (N_24685,N_23825,N_23857);
xnor U24686 (N_24686,N_24302,N_23982);
or U24687 (N_24687,N_23934,N_24260);
nor U24688 (N_24688,N_24179,N_24260);
nor U24689 (N_24689,N_23878,N_24077);
and U24690 (N_24690,N_24224,N_23890);
and U24691 (N_24691,N_24285,N_23969);
xnor U24692 (N_24692,N_24098,N_24267);
and U24693 (N_24693,N_23840,N_24244);
or U24694 (N_24694,N_23984,N_23816);
xnor U24695 (N_24695,N_24332,N_24019);
nor U24696 (N_24696,N_24080,N_24064);
nor U24697 (N_24697,N_23891,N_23985);
and U24698 (N_24698,N_24150,N_24266);
nor U24699 (N_24699,N_24340,N_24363);
nand U24700 (N_24700,N_24185,N_23859);
xor U24701 (N_24701,N_24012,N_24275);
xor U24702 (N_24702,N_24030,N_24087);
nor U24703 (N_24703,N_24195,N_24309);
xor U24704 (N_24704,N_24309,N_24156);
xor U24705 (N_24705,N_24284,N_24232);
nor U24706 (N_24706,N_23789,N_23890);
xnor U24707 (N_24707,N_24017,N_24362);
or U24708 (N_24708,N_24052,N_24120);
or U24709 (N_24709,N_24182,N_23834);
xnor U24710 (N_24710,N_24361,N_24024);
and U24711 (N_24711,N_24300,N_24051);
nand U24712 (N_24712,N_24032,N_23766);
xor U24713 (N_24713,N_24278,N_24286);
or U24714 (N_24714,N_24285,N_23985);
and U24715 (N_24715,N_24100,N_24079);
nand U24716 (N_24716,N_23906,N_23775);
and U24717 (N_24717,N_23774,N_24350);
xnor U24718 (N_24718,N_24234,N_24176);
xor U24719 (N_24719,N_23858,N_24128);
xor U24720 (N_24720,N_24069,N_24208);
nor U24721 (N_24721,N_24258,N_24143);
and U24722 (N_24722,N_24277,N_24289);
nand U24723 (N_24723,N_24114,N_23909);
and U24724 (N_24724,N_24079,N_23889);
and U24725 (N_24725,N_24367,N_23804);
nand U24726 (N_24726,N_24090,N_24197);
nor U24727 (N_24727,N_24367,N_24195);
nand U24728 (N_24728,N_23960,N_23990);
or U24729 (N_24729,N_24144,N_23807);
and U24730 (N_24730,N_23913,N_23884);
and U24731 (N_24731,N_24055,N_24057);
nor U24732 (N_24732,N_23827,N_24286);
nor U24733 (N_24733,N_23932,N_23905);
nand U24734 (N_24734,N_24158,N_24330);
xor U24735 (N_24735,N_23877,N_23848);
or U24736 (N_24736,N_23811,N_23885);
xor U24737 (N_24737,N_24324,N_24019);
and U24738 (N_24738,N_23856,N_24056);
nor U24739 (N_24739,N_23974,N_23948);
or U24740 (N_24740,N_23777,N_23980);
nand U24741 (N_24741,N_24109,N_24234);
nor U24742 (N_24742,N_24121,N_23835);
and U24743 (N_24743,N_24368,N_24136);
or U24744 (N_24744,N_24260,N_24314);
nand U24745 (N_24745,N_24335,N_24189);
nor U24746 (N_24746,N_24318,N_24193);
nor U24747 (N_24747,N_23857,N_23986);
nor U24748 (N_24748,N_23872,N_24068);
nor U24749 (N_24749,N_24316,N_24003);
or U24750 (N_24750,N_24080,N_24286);
and U24751 (N_24751,N_24022,N_24339);
xnor U24752 (N_24752,N_23766,N_23987);
and U24753 (N_24753,N_23999,N_24268);
or U24754 (N_24754,N_24226,N_23795);
nand U24755 (N_24755,N_23905,N_24131);
nand U24756 (N_24756,N_23907,N_23892);
nand U24757 (N_24757,N_23854,N_24302);
and U24758 (N_24758,N_24147,N_24201);
or U24759 (N_24759,N_24096,N_24275);
xnor U24760 (N_24760,N_24262,N_24048);
or U24761 (N_24761,N_24336,N_24244);
nand U24762 (N_24762,N_23964,N_24101);
xnor U24763 (N_24763,N_24316,N_24353);
or U24764 (N_24764,N_24262,N_24339);
nor U24765 (N_24765,N_24245,N_23767);
or U24766 (N_24766,N_23953,N_24337);
nand U24767 (N_24767,N_24102,N_24319);
nand U24768 (N_24768,N_24115,N_23890);
nor U24769 (N_24769,N_23948,N_24091);
xnor U24770 (N_24770,N_24215,N_24268);
nor U24771 (N_24771,N_23895,N_24270);
nor U24772 (N_24772,N_24059,N_24170);
nand U24773 (N_24773,N_23756,N_24215);
or U24774 (N_24774,N_23849,N_23966);
nor U24775 (N_24775,N_23868,N_24106);
and U24776 (N_24776,N_24058,N_24248);
and U24777 (N_24777,N_24355,N_23935);
and U24778 (N_24778,N_24053,N_24093);
or U24779 (N_24779,N_23757,N_24236);
and U24780 (N_24780,N_24103,N_24172);
or U24781 (N_24781,N_23978,N_23752);
nand U24782 (N_24782,N_24225,N_23910);
and U24783 (N_24783,N_23826,N_23986);
and U24784 (N_24784,N_24055,N_23946);
nor U24785 (N_24785,N_23788,N_23972);
and U24786 (N_24786,N_23956,N_23919);
and U24787 (N_24787,N_23836,N_23939);
xor U24788 (N_24788,N_24232,N_24129);
nand U24789 (N_24789,N_24122,N_24062);
or U24790 (N_24790,N_24234,N_23907);
or U24791 (N_24791,N_23961,N_24277);
nor U24792 (N_24792,N_23866,N_24247);
nor U24793 (N_24793,N_23821,N_24053);
nor U24794 (N_24794,N_24085,N_24101);
nand U24795 (N_24795,N_24153,N_24129);
nor U24796 (N_24796,N_23960,N_24064);
or U24797 (N_24797,N_24251,N_24319);
or U24798 (N_24798,N_23786,N_24271);
nand U24799 (N_24799,N_23808,N_24178);
xor U24800 (N_24800,N_23997,N_24282);
nor U24801 (N_24801,N_23928,N_24024);
nor U24802 (N_24802,N_23826,N_24331);
nor U24803 (N_24803,N_23880,N_24010);
nand U24804 (N_24804,N_23936,N_24233);
nand U24805 (N_24805,N_23952,N_23782);
and U24806 (N_24806,N_23885,N_23909);
and U24807 (N_24807,N_23813,N_23949);
nand U24808 (N_24808,N_23768,N_24154);
and U24809 (N_24809,N_24053,N_24008);
or U24810 (N_24810,N_24314,N_23955);
nor U24811 (N_24811,N_24348,N_23939);
nand U24812 (N_24812,N_23923,N_24088);
nand U24813 (N_24813,N_23843,N_24347);
nand U24814 (N_24814,N_24251,N_24187);
nor U24815 (N_24815,N_24044,N_23821);
nor U24816 (N_24816,N_24024,N_23937);
nand U24817 (N_24817,N_24203,N_24219);
nand U24818 (N_24818,N_24197,N_24011);
and U24819 (N_24819,N_24087,N_24110);
or U24820 (N_24820,N_24003,N_24246);
xor U24821 (N_24821,N_24041,N_24210);
xnor U24822 (N_24822,N_24322,N_24209);
or U24823 (N_24823,N_23883,N_24088);
or U24824 (N_24824,N_24313,N_24233);
nor U24825 (N_24825,N_24065,N_24269);
nand U24826 (N_24826,N_24215,N_24343);
xor U24827 (N_24827,N_23875,N_24332);
and U24828 (N_24828,N_23829,N_23785);
nand U24829 (N_24829,N_24293,N_23764);
xor U24830 (N_24830,N_23813,N_23939);
nand U24831 (N_24831,N_24342,N_24017);
nor U24832 (N_24832,N_24187,N_24269);
or U24833 (N_24833,N_24249,N_23984);
nand U24834 (N_24834,N_24290,N_24317);
and U24835 (N_24835,N_23858,N_24025);
nor U24836 (N_24836,N_24192,N_24042);
nand U24837 (N_24837,N_23761,N_24284);
nor U24838 (N_24838,N_24228,N_23891);
xnor U24839 (N_24839,N_24294,N_24244);
nand U24840 (N_24840,N_24349,N_23838);
or U24841 (N_24841,N_23956,N_24083);
and U24842 (N_24842,N_23952,N_23786);
xnor U24843 (N_24843,N_24323,N_24237);
or U24844 (N_24844,N_24338,N_24268);
and U24845 (N_24845,N_24006,N_24159);
or U24846 (N_24846,N_23843,N_23796);
and U24847 (N_24847,N_24248,N_24220);
and U24848 (N_24848,N_23781,N_23878);
or U24849 (N_24849,N_23994,N_24136);
nand U24850 (N_24850,N_24087,N_24262);
nor U24851 (N_24851,N_23777,N_24360);
nand U24852 (N_24852,N_23884,N_24345);
xor U24853 (N_24853,N_24237,N_24342);
xnor U24854 (N_24854,N_24371,N_23970);
xor U24855 (N_24855,N_24148,N_23811);
or U24856 (N_24856,N_24063,N_24118);
and U24857 (N_24857,N_24013,N_24225);
nor U24858 (N_24858,N_23829,N_24369);
nand U24859 (N_24859,N_23986,N_23888);
xnor U24860 (N_24860,N_23806,N_23946);
nor U24861 (N_24861,N_23815,N_24207);
and U24862 (N_24862,N_23822,N_24371);
and U24863 (N_24863,N_24049,N_24035);
or U24864 (N_24864,N_24343,N_24327);
nand U24865 (N_24865,N_24339,N_24319);
nor U24866 (N_24866,N_24017,N_23887);
nor U24867 (N_24867,N_23906,N_23833);
nor U24868 (N_24868,N_24188,N_24329);
nand U24869 (N_24869,N_23777,N_24348);
and U24870 (N_24870,N_23776,N_24022);
nand U24871 (N_24871,N_24317,N_24009);
or U24872 (N_24872,N_23785,N_24247);
nor U24873 (N_24873,N_23940,N_24327);
xor U24874 (N_24874,N_23965,N_24244);
nor U24875 (N_24875,N_23793,N_24292);
xnor U24876 (N_24876,N_23923,N_24238);
and U24877 (N_24877,N_24343,N_23777);
nand U24878 (N_24878,N_24171,N_23955);
or U24879 (N_24879,N_24183,N_23812);
nand U24880 (N_24880,N_23960,N_23766);
or U24881 (N_24881,N_23751,N_24256);
and U24882 (N_24882,N_23974,N_23935);
or U24883 (N_24883,N_24255,N_23927);
xor U24884 (N_24884,N_23800,N_23977);
xor U24885 (N_24885,N_23857,N_24028);
and U24886 (N_24886,N_24230,N_23901);
xnor U24887 (N_24887,N_24264,N_24265);
nand U24888 (N_24888,N_23790,N_24061);
xnor U24889 (N_24889,N_24255,N_24048);
nor U24890 (N_24890,N_24340,N_24371);
nand U24891 (N_24891,N_23834,N_24063);
nand U24892 (N_24892,N_23874,N_24038);
nor U24893 (N_24893,N_23909,N_23817);
nand U24894 (N_24894,N_24184,N_23972);
and U24895 (N_24895,N_24328,N_24255);
nand U24896 (N_24896,N_24246,N_23933);
or U24897 (N_24897,N_23883,N_23948);
nand U24898 (N_24898,N_24224,N_23907);
and U24899 (N_24899,N_23782,N_24226);
nand U24900 (N_24900,N_24271,N_24200);
or U24901 (N_24901,N_23766,N_24073);
and U24902 (N_24902,N_24286,N_23983);
xor U24903 (N_24903,N_24196,N_24161);
xnor U24904 (N_24904,N_24207,N_24362);
xor U24905 (N_24905,N_24357,N_24216);
xnor U24906 (N_24906,N_23903,N_24129);
nor U24907 (N_24907,N_24359,N_24169);
and U24908 (N_24908,N_24231,N_23953);
or U24909 (N_24909,N_23904,N_24103);
nand U24910 (N_24910,N_23814,N_23974);
or U24911 (N_24911,N_24009,N_23952);
xor U24912 (N_24912,N_24243,N_24212);
and U24913 (N_24913,N_23977,N_24356);
and U24914 (N_24914,N_24044,N_23799);
nor U24915 (N_24915,N_24293,N_24227);
xor U24916 (N_24916,N_23948,N_24030);
nand U24917 (N_24917,N_23772,N_24069);
nor U24918 (N_24918,N_24030,N_23982);
nor U24919 (N_24919,N_24279,N_24075);
xor U24920 (N_24920,N_24201,N_23915);
or U24921 (N_24921,N_23957,N_24231);
and U24922 (N_24922,N_23922,N_23855);
xor U24923 (N_24923,N_24161,N_23860);
nand U24924 (N_24924,N_23999,N_23762);
nor U24925 (N_24925,N_24159,N_24180);
nor U24926 (N_24926,N_23928,N_23821);
nand U24927 (N_24927,N_24321,N_24167);
nor U24928 (N_24928,N_24063,N_23961);
nor U24929 (N_24929,N_23868,N_23756);
nand U24930 (N_24930,N_24227,N_23884);
nand U24931 (N_24931,N_24008,N_24107);
or U24932 (N_24932,N_23798,N_23843);
and U24933 (N_24933,N_23816,N_23827);
and U24934 (N_24934,N_24313,N_24055);
xor U24935 (N_24935,N_24352,N_24068);
xnor U24936 (N_24936,N_23906,N_24111);
nor U24937 (N_24937,N_24096,N_24221);
nand U24938 (N_24938,N_24365,N_23888);
nor U24939 (N_24939,N_24220,N_23923);
nor U24940 (N_24940,N_24191,N_24335);
nor U24941 (N_24941,N_23863,N_24003);
nand U24942 (N_24942,N_23799,N_24273);
nor U24943 (N_24943,N_24137,N_23787);
and U24944 (N_24944,N_24184,N_24324);
nor U24945 (N_24945,N_23969,N_24080);
or U24946 (N_24946,N_24099,N_24302);
nor U24947 (N_24947,N_23885,N_23959);
nor U24948 (N_24948,N_24118,N_24358);
nand U24949 (N_24949,N_23862,N_24153);
and U24950 (N_24950,N_23981,N_24319);
nand U24951 (N_24951,N_24180,N_24261);
or U24952 (N_24952,N_24159,N_24338);
nor U24953 (N_24953,N_23982,N_24121);
xnor U24954 (N_24954,N_24211,N_24195);
nor U24955 (N_24955,N_24262,N_23769);
nor U24956 (N_24956,N_24220,N_23907);
nand U24957 (N_24957,N_23794,N_24198);
xor U24958 (N_24958,N_24198,N_23874);
xor U24959 (N_24959,N_24176,N_24012);
xor U24960 (N_24960,N_24194,N_23756);
and U24961 (N_24961,N_24057,N_24222);
xnor U24962 (N_24962,N_23947,N_23874);
xnor U24963 (N_24963,N_23764,N_24163);
and U24964 (N_24964,N_23861,N_24104);
and U24965 (N_24965,N_24340,N_24026);
or U24966 (N_24966,N_24213,N_23863);
and U24967 (N_24967,N_24343,N_24096);
or U24968 (N_24968,N_24361,N_24275);
and U24969 (N_24969,N_23777,N_23994);
nor U24970 (N_24970,N_23931,N_23861);
xnor U24971 (N_24971,N_24299,N_23858);
nor U24972 (N_24972,N_23855,N_24225);
and U24973 (N_24973,N_24158,N_23978);
nand U24974 (N_24974,N_24032,N_24206);
xnor U24975 (N_24975,N_23761,N_24324);
nand U24976 (N_24976,N_23752,N_24004);
and U24977 (N_24977,N_23954,N_24249);
nand U24978 (N_24978,N_23968,N_24198);
or U24979 (N_24979,N_23753,N_23757);
xor U24980 (N_24980,N_23950,N_23998);
and U24981 (N_24981,N_24193,N_24209);
xnor U24982 (N_24982,N_24074,N_23772);
nand U24983 (N_24983,N_23975,N_23901);
xnor U24984 (N_24984,N_23900,N_24072);
xnor U24985 (N_24985,N_23977,N_23933);
nand U24986 (N_24986,N_23921,N_23755);
or U24987 (N_24987,N_23967,N_23757);
xnor U24988 (N_24988,N_23966,N_24175);
nor U24989 (N_24989,N_24213,N_23912);
nand U24990 (N_24990,N_23977,N_23755);
and U24991 (N_24991,N_24064,N_24084);
nor U24992 (N_24992,N_23804,N_23922);
and U24993 (N_24993,N_24300,N_24027);
xor U24994 (N_24994,N_24289,N_23823);
and U24995 (N_24995,N_24012,N_23918);
nor U24996 (N_24996,N_24225,N_24334);
or U24997 (N_24997,N_23831,N_24193);
and U24998 (N_24998,N_23941,N_24031);
xnor U24999 (N_24999,N_23929,N_23835);
and UO_0 (O_0,N_24872,N_24828);
xor UO_1 (O_1,N_24810,N_24502);
or UO_2 (O_2,N_24498,N_24980);
nand UO_3 (O_3,N_24838,N_24598);
or UO_4 (O_4,N_24744,N_24734);
and UO_5 (O_5,N_24645,N_24543);
xor UO_6 (O_6,N_24903,N_24932);
and UO_7 (O_7,N_24576,N_24457);
nor UO_8 (O_8,N_24473,N_24622);
or UO_9 (O_9,N_24845,N_24822);
nand UO_10 (O_10,N_24833,N_24879);
nor UO_11 (O_11,N_24672,N_24963);
nor UO_12 (O_12,N_24491,N_24794);
or UO_13 (O_13,N_24504,N_24820);
nor UO_14 (O_14,N_24816,N_24894);
nor UO_15 (O_15,N_24818,N_24505);
nor UO_16 (O_16,N_24771,N_24391);
xor UO_17 (O_17,N_24933,N_24913);
or UO_18 (O_18,N_24501,N_24817);
or UO_19 (O_19,N_24411,N_24472);
nor UO_20 (O_20,N_24451,N_24722);
and UO_21 (O_21,N_24625,N_24954);
nor UO_22 (O_22,N_24615,N_24521);
or UO_23 (O_23,N_24563,N_24799);
xor UO_24 (O_24,N_24808,N_24789);
nand UO_25 (O_25,N_24958,N_24815);
and UO_26 (O_26,N_24507,N_24747);
and UO_27 (O_27,N_24623,N_24648);
or UO_28 (O_28,N_24780,N_24924);
xor UO_29 (O_29,N_24436,N_24417);
nor UO_30 (O_30,N_24635,N_24555);
xor UO_31 (O_31,N_24401,N_24392);
or UO_32 (O_32,N_24773,N_24668);
nor UO_33 (O_33,N_24616,N_24809);
xor UO_34 (O_34,N_24936,N_24530);
and UO_35 (O_35,N_24721,N_24937);
xor UO_36 (O_36,N_24792,N_24618);
or UO_37 (O_37,N_24603,N_24770);
nand UO_38 (O_38,N_24713,N_24741);
xnor UO_39 (O_39,N_24998,N_24513);
xnor UO_40 (O_40,N_24431,N_24655);
nand UO_41 (O_41,N_24915,N_24891);
xor UO_42 (O_42,N_24724,N_24581);
nor UO_43 (O_43,N_24824,N_24865);
xor UO_44 (O_44,N_24536,N_24985);
xor UO_45 (O_45,N_24531,N_24447);
nor UO_46 (O_46,N_24596,N_24953);
xor UO_47 (O_47,N_24571,N_24979);
nand UO_48 (O_48,N_24628,N_24404);
or UO_49 (O_49,N_24664,N_24493);
nand UO_50 (O_50,N_24446,N_24853);
and UO_51 (O_51,N_24701,N_24437);
or UO_52 (O_52,N_24720,N_24606);
or UO_53 (O_53,N_24978,N_24757);
nor UO_54 (O_54,N_24477,N_24442);
or UO_55 (O_55,N_24718,N_24674);
nand UO_56 (O_56,N_24604,N_24786);
or UO_57 (O_57,N_24777,N_24611);
nand UO_58 (O_58,N_24752,N_24990);
nand UO_59 (O_59,N_24454,N_24423);
or UO_60 (O_60,N_24515,N_24609);
nand UO_61 (O_61,N_24970,N_24884);
nand UO_62 (O_62,N_24443,N_24561);
xnor UO_63 (O_63,N_24841,N_24753);
or UO_64 (O_64,N_24659,N_24748);
or UO_65 (O_65,N_24935,N_24601);
and UO_66 (O_66,N_24863,N_24983);
nor UO_67 (O_67,N_24756,N_24389);
and UO_68 (O_68,N_24877,N_24661);
xnor UO_69 (O_69,N_24699,N_24846);
and UO_70 (O_70,N_24396,N_24790);
nor UO_71 (O_71,N_24567,N_24545);
nand UO_72 (O_72,N_24572,N_24565);
xnor UO_73 (O_73,N_24727,N_24984);
xor UO_74 (O_74,N_24564,N_24868);
xor UO_75 (O_75,N_24407,N_24675);
nand UO_76 (O_76,N_24842,N_24586);
xnor UO_77 (O_77,N_24728,N_24951);
nor UO_78 (O_78,N_24918,N_24669);
nor UO_79 (O_79,N_24427,N_24408);
or UO_80 (O_80,N_24546,N_24731);
nor UO_81 (O_81,N_24957,N_24766);
xor UO_82 (O_82,N_24969,N_24484);
xnor UO_83 (O_83,N_24959,N_24854);
nand UO_84 (O_84,N_24716,N_24459);
nand UO_85 (O_85,N_24919,N_24509);
xnor UO_86 (O_86,N_24730,N_24435);
and UO_87 (O_87,N_24923,N_24767);
nor UO_88 (O_88,N_24776,N_24573);
nor UO_89 (O_89,N_24551,N_24445);
nor UO_90 (O_90,N_24859,N_24589);
nand UO_91 (O_91,N_24517,N_24631);
nand UO_92 (O_92,N_24848,N_24483);
nand UO_93 (O_93,N_24626,N_24761);
nor UO_94 (O_94,N_24488,N_24580);
and UO_95 (O_95,N_24544,N_24649);
nand UO_96 (O_96,N_24482,N_24821);
nand UO_97 (O_97,N_24795,N_24432);
nor UO_98 (O_98,N_24585,N_24926);
and UO_99 (O_99,N_24746,N_24945);
xor UO_100 (O_100,N_24568,N_24535);
or UO_101 (O_101,N_24996,N_24578);
nor UO_102 (O_102,N_24697,N_24575);
xor UO_103 (O_103,N_24434,N_24928);
nor UO_104 (O_104,N_24931,N_24930);
nand UO_105 (O_105,N_24634,N_24642);
nor UO_106 (O_106,N_24395,N_24869);
and UO_107 (O_107,N_24896,N_24736);
or UO_108 (O_108,N_24384,N_24494);
xnor UO_109 (O_109,N_24774,N_24554);
xor UO_110 (O_110,N_24480,N_24782);
or UO_111 (O_111,N_24379,N_24876);
nand UO_112 (O_112,N_24624,N_24909);
or UO_113 (O_113,N_24765,N_24485);
nor UO_114 (O_114,N_24512,N_24698);
xor UO_115 (O_115,N_24523,N_24988);
or UO_116 (O_116,N_24764,N_24883);
nand UO_117 (O_117,N_24667,N_24652);
or UO_118 (O_118,N_24421,N_24579);
nor UO_119 (O_119,N_24745,N_24556);
nand UO_120 (O_120,N_24995,N_24525);
and UO_121 (O_121,N_24663,N_24438);
nor UO_122 (O_122,N_24662,N_24458);
and UO_123 (O_123,N_24908,N_24592);
or UO_124 (O_124,N_24973,N_24644);
or UO_125 (O_125,N_24733,N_24600);
nor UO_126 (O_126,N_24981,N_24653);
or UO_127 (O_127,N_24882,N_24855);
nor UO_128 (O_128,N_24916,N_24922);
or UO_129 (O_129,N_24834,N_24450);
and UO_130 (O_130,N_24813,N_24583);
or UO_131 (O_131,N_24430,N_24617);
and UO_132 (O_132,N_24852,N_24656);
xor UO_133 (O_133,N_24867,N_24938);
nor UO_134 (O_134,N_24866,N_24738);
xnor UO_135 (O_135,N_24829,N_24641);
or UO_136 (O_136,N_24380,N_24499);
or UO_137 (O_137,N_24775,N_24461);
xnor UO_138 (O_138,N_24428,N_24468);
and UO_139 (O_139,N_24467,N_24570);
or UO_140 (O_140,N_24832,N_24489);
xor UO_141 (O_141,N_24900,N_24386);
nand UO_142 (O_142,N_24519,N_24574);
or UO_143 (O_143,N_24940,N_24463);
nand UO_144 (O_144,N_24510,N_24768);
xor UO_145 (O_145,N_24708,N_24495);
nor UO_146 (O_146,N_24976,N_24385);
nor UO_147 (O_147,N_24582,N_24986);
nand UO_148 (O_148,N_24650,N_24388);
xor UO_149 (O_149,N_24381,N_24812);
nor UO_150 (O_150,N_24857,N_24696);
nand UO_151 (O_151,N_24426,N_24899);
and UO_152 (O_152,N_24383,N_24398);
nor UO_153 (O_153,N_24952,N_24681);
nand UO_154 (O_154,N_24717,N_24693);
xor UO_155 (O_155,N_24605,N_24471);
and UO_156 (O_156,N_24397,N_24703);
nand UO_157 (O_157,N_24440,N_24711);
or UO_158 (O_158,N_24943,N_24419);
or UO_159 (O_159,N_24588,N_24885);
xor UO_160 (O_160,N_24704,N_24971);
and UO_161 (O_161,N_24939,N_24898);
nor UO_162 (O_162,N_24783,N_24814);
or UO_163 (O_163,N_24539,N_24695);
or UO_164 (O_164,N_24679,N_24686);
nor UO_165 (O_165,N_24878,N_24566);
or UO_166 (O_166,N_24921,N_24715);
or UO_167 (O_167,N_24627,N_24590);
nor UO_168 (O_168,N_24464,N_24726);
and UO_169 (O_169,N_24929,N_24439);
or UO_170 (O_170,N_24714,N_24997);
or UO_171 (O_171,N_24897,N_24914);
and UO_172 (O_172,N_24678,N_24851);
xor UO_173 (O_173,N_24961,N_24562);
and UO_174 (O_174,N_24524,N_24462);
xor UO_175 (O_175,N_24880,N_24413);
or UO_176 (O_176,N_24839,N_24974);
and UO_177 (O_177,N_24784,N_24497);
nand UO_178 (O_178,N_24415,N_24861);
xor UO_179 (O_179,N_24665,N_24874);
or UO_180 (O_180,N_24862,N_24781);
xnor UO_181 (O_181,N_24827,N_24390);
nand UO_182 (O_182,N_24557,N_24797);
and UO_183 (O_183,N_24378,N_24599);
nor UO_184 (O_184,N_24890,N_24393);
and UO_185 (O_185,N_24503,N_24705);
or UO_186 (O_186,N_24420,N_24685);
nor UO_187 (O_187,N_24910,N_24907);
or UO_188 (O_188,N_24492,N_24860);
and UO_189 (O_189,N_24700,N_24691);
nand UO_190 (O_190,N_24772,N_24858);
or UO_191 (O_191,N_24620,N_24487);
nor UO_192 (O_192,N_24619,N_24706);
nand UO_193 (O_193,N_24873,N_24640);
nor UO_194 (O_194,N_24399,N_24762);
xor UO_195 (O_195,N_24486,N_24466);
or UO_196 (O_196,N_24830,N_24893);
xor UO_197 (O_197,N_24688,N_24725);
nor UO_198 (O_198,N_24680,N_24966);
nand UO_199 (O_199,N_24840,N_24707);
nor UO_200 (O_200,N_24751,N_24904);
nor UO_201 (O_201,N_24825,N_24710);
nand UO_202 (O_202,N_24514,N_24887);
or UO_203 (O_203,N_24750,N_24496);
nor UO_204 (O_204,N_24759,N_24989);
or UO_205 (O_205,N_24632,N_24831);
nand UO_206 (O_206,N_24844,N_24796);
nand UO_207 (O_207,N_24376,N_24591);
nand UO_208 (O_208,N_24490,N_24638);
or UO_209 (O_209,N_24944,N_24740);
xnor UO_210 (O_210,N_24526,N_24889);
nand UO_211 (O_211,N_24453,N_24422);
nor UO_212 (O_212,N_24639,N_24947);
or UO_213 (O_213,N_24418,N_24843);
and UO_214 (O_214,N_24850,N_24875);
and UO_215 (O_215,N_24394,N_24478);
nor UO_216 (O_216,N_24684,N_24597);
nor UO_217 (O_217,N_24529,N_24595);
or UO_218 (O_218,N_24927,N_24637);
and UO_219 (O_219,N_24456,N_24612);
and UO_220 (O_220,N_24798,N_24587);
and UO_221 (O_221,N_24677,N_24712);
xor UO_222 (O_222,N_24569,N_24801);
nor UO_223 (O_223,N_24965,N_24630);
nand UO_224 (O_224,N_24802,N_24651);
nor UO_225 (O_225,N_24755,N_24476);
nor UO_226 (O_226,N_24892,N_24694);
nor UO_227 (O_227,N_24646,N_24778);
xor UO_228 (O_228,N_24607,N_24425);
xor UO_229 (O_229,N_24534,N_24673);
nor UO_230 (O_230,N_24823,N_24657);
or UO_231 (O_231,N_24807,N_24584);
or UO_232 (O_232,N_24416,N_24743);
or UO_233 (O_233,N_24593,N_24560);
and UO_234 (O_234,N_24402,N_24660);
xnor UO_235 (O_235,N_24956,N_24542);
nand UO_236 (O_236,N_24621,N_24702);
nand UO_237 (O_237,N_24779,N_24805);
xnor UO_238 (O_238,N_24739,N_24479);
nand UO_239 (O_239,N_24690,N_24683);
xor UO_240 (O_240,N_24760,N_24475);
or UO_241 (O_241,N_24934,N_24559);
nand UO_242 (O_242,N_24785,N_24469);
and UO_243 (O_243,N_24671,N_24452);
nand UO_244 (O_244,N_24888,N_24835);
nand UO_245 (O_245,N_24803,N_24837);
and UO_246 (O_246,N_24474,N_24553);
and UO_247 (O_247,N_24993,N_24964);
nand UO_248 (O_248,N_24847,N_24955);
xnor UO_249 (O_249,N_24800,N_24414);
nor UO_250 (O_250,N_24975,N_24441);
nor UO_251 (O_251,N_24972,N_24682);
nand UO_252 (O_252,N_24749,N_24901);
and UO_253 (O_253,N_24946,N_24527);
and UO_254 (O_254,N_24577,N_24613);
or UO_255 (O_255,N_24532,N_24806);
and UO_256 (O_256,N_24382,N_24870);
nand UO_257 (O_257,N_24948,N_24643);
and UO_258 (O_258,N_24737,N_24917);
nand UO_259 (O_259,N_24925,N_24787);
or UO_260 (O_260,N_24856,N_24732);
nor UO_261 (O_261,N_24670,N_24886);
xor UO_262 (O_262,N_24864,N_24788);
and UO_263 (O_263,N_24522,N_24742);
xnor UO_264 (O_264,N_24518,N_24541);
xor UO_265 (O_265,N_24511,N_24412);
and UO_266 (O_266,N_24528,N_24836);
or UO_267 (O_267,N_24791,N_24537);
nand UO_268 (O_268,N_24455,N_24602);
nand UO_269 (O_269,N_24424,N_24444);
xor UO_270 (O_270,N_24552,N_24547);
and UO_271 (O_271,N_24448,N_24538);
nand UO_272 (O_272,N_24811,N_24968);
or UO_273 (O_273,N_24949,N_24709);
xor UO_274 (O_274,N_24941,N_24647);
and UO_275 (O_275,N_24375,N_24719);
nand UO_276 (O_276,N_24689,N_24905);
or UO_277 (O_277,N_24594,N_24520);
nor UO_278 (O_278,N_24912,N_24902);
or UO_279 (O_279,N_24377,N_24793);
nor UO_280 (O_280,N_24999,N_24735);
or UO_281 (O_281,N_24881,N_24449);
xnor UO_282 (O_282,N_24403,N_24994);
or UO_283 (O_283,N_24769,N_24687);
and UO_284 (O_284,N_24723,N_24614);
or UO_285 (O_285,N_24506,N_24992);
and UO_286 (O_286,N_24508,N_24540);
and UO_287 (O_287,N_24991,N_24465);
and UO_288 (O_288,N_24558,N_24654);
nor UO_289 (O_289,N_24516,N_24533);
xnor UO_290 (O_290,N_24460,N_24610);
nand UO_291 (O_291,N_24920,N_24549);
xor UO_292 (O_292,N_24942,N_24633);
xnor UO_293 (O_293,N_24550,N_24895);
nand UO_294 (O_294,N_24826,N_24763);
or UO_295 (O_295,N_24729,N_24950);
xnor UO_296 (O_296,N_24977,N_24849);
and UO_297 (O_297,N_24758,N_24692);
nand UO_298 (O_298,N_24982,N_24629);
xor UO_299 (O_299,N_24967,N_24410);
nor UO_300 (O_300,N_24911,N_24500);
or UO_301 (O_301,N_24429,N_24676);
nand UO_302 (O_302,N_24409,N_24960);
and UO_303 (O_303,N_24405,N_24658);
nor UO_304 (O_304,N_24433,N_24636);
and UO_305 (O_305,N_24470,N_24548);
nand UO_306 (O_306,N_24481,N_24871);
and UO_307 (O_307,N_24400,N_24819);
nand UO_308 (O_308,N_24987,N_24754);
and UO_309 (O_309,N_24906,N_24608);
nor UO_310 (O_310,N_24804,N_24962);
xnor UO_311 (O_311,N_24666,N_24406);
xnor UO_312 (O_312,N_24387,N_24698);
nand UO_313 (O_313,N_24781,N_24530);
xnor UO_314 (O_314,N_24481,N_24692);
or UO_315 (O_315,N_24977,N_24682);
or UO_316 (O_316,N_24974,N_24967);
nor UO_317 (O_317,N_24571,N_24696);
nor UO_318 (O_318,N_24473,N_24436);
nor UO_319 (O_319,N_24690,N_24611);
nand UO_320 (O_320,N_24432,N_24592);
or UO_321 (O_321,N_24675,N_24866);
nor UO_322 (O_322,N_24850,N_24589);
nor UO_323 (O_323,N_24717,N_24896);
nor UO_324 (O_324,N_24700,N_24513);
nand UO_325 (O_325,N_24752,N_24767);
nor UO_326 (O_326,N_24797,N_24878);
or UO_327 (O_327,N_24693,N_24808);
nor UO_328 (O_328,N_24764,N_24808);
nand UO_329 (O_329,N_24448,N_24804);
and UO_330 (O_330,N_24568,N_24845);
xor UO_331 (O_331,N_24969,N_24791);
xnor UO_332 (O_332,N_24796,N_24996);
nand UO_333 (O_333,N_24946,N_24976);
and UO_334 (O_334,N_24740,N_24828);
xnor UO_335 (O_335,N_24830,N_24636);
nand UO_336 (O_336,N_24952,N_24671);
or UO_337 (O_337,N_24710,N_24635);
xor UO_338 (O_338,N_24448,N_24990);
xor UO_339 (O_339,N_24634,N_24911);
nor UO_340 (O_340,N_24933,N_24600);
and UO_341 (O_341,N_24909,N_24876);
nand UO_342 (O_342,N_24883,N_24745);
and UO_343 (O_343,N_24728,N_24775);
xnor UO_344 (O_344,N_24453,N_24791);
and UO_345 (O_345,N_24849,N_24426);
or UO_346 (O_346,N_24840,N_24714);
xnor UO_347 (O_347,N_24539,N_24900);
and UO_348 (O_348,N_24702,N_24889);
nand UO_349 (O_349,N_24659,N_24873);
xor UO_350 (O_350,N_24704,N_24891);
or UO_351 (O_351,N_24684,N_24654);
and UO_352 (O_352,N_24668,N_24932);
and UO_353 (O_353,N_24391,N_24524);
or UO_354 (O_354,N_24923,N_24660);
and UO_355 (O_355,N_24494,N_24538);
and UO_356 (O_356,N_24592,N_24574);
xnor UO_357 (O_357,N_24881,N_24628);
and UO_358 (O_358,N_24993,N_24635);
nor UO_359 (O_359,N_24717,N_24850);
nand UO_360 (O_360,N_24938,N_24575);
or UO_361 (O_361,N_24910,N_24521);
xnor UO_362 (O_362,N_24758,N_24960);
nor UO_363 (O_363,N_24722,N_24432);
xnor UO_364 (O_364,N_24487,N_24667);
xnor UO_365 (O_365,N_24483,N_24669);
or UO_366 (O_366,N_24677,N_24460);
nand UO_367 (O_367,N_24780,N_24447);
or UO_368 (O_368,N_24587,N_24616);
nand UO_369 (O_369,N_24964,N_24517);
nand UO_370 (O_370,N_24427,N_24450);
nor UO_371 (O_371,N_24690,N_24448);
and UO_372 (O_372,N_24866,N_24895);
nand UO_373 (O_373,N_24601,N_24749);
nand UO_374 (O_374,N_24859,N_24502);
nor UO_375 (O_375,N_24963,N_24695);
nor UO_376 (O_376,N_24770,N_24427);
and UO_377 (O_377,N_24807,N_24758);
xor UO_378 (O_378,N_24616,N_24406);
nor UO_379 (O_379,N_24939,N_24812);
and UO_380 (O_380,N_24932,N_24443);
nor UO_381 (O_381,N_24452,N_24517);
nor UO_382 (O_382,N_24780,N_24422);
xor UO_383 (O_383,N_24784,N_24783);
nor UO_384 (O_384,N_24554,N_24693);
nand UO_385 (O_385,N_24428,N_24761);
nor UO_386 (O_386,N_24772,N_24514);
nand UO_387 (O_387,N_24509,N_24910);
and UO_388 (O_388,N_24848,N_24473);
xnor UO_389 (O_389,N_24669,N_24566);
or UO_390 (O_390,N_24475,N_24743);
nor UO_391 (O_391,N_24958,N_24694);
nand UO_392 (O_392,N_24853,N_24814);
nand UO_393 (O_393,N_24484,N_24712);
or UO_394 (O_394,N_24700,N_24672);
nor UO_395 (O_395,N_24436,N_24985);
nor UO_396 (O_396,N_24976,N_24416);
and UO_397 (O_397,N_24667,N_24502);
xor UO_398 (O_398,N_24450,N_24522);
or UO_399 (O_399,N_24887,N_24664);
xor UO_400 (O_400,N_24625,N_24914);
nor UO_401 (O_401,N_24574,N_24704);
nor UO_402 (O_402,N_24434,N_24979);
and UO_403 (O_403,N_24789,N_24822);
or UO_404 (O_404,N_24977,N_24662);
nor UO_405 (O_405,N_24481,N_24552);
xnor UO_406 (O_406,N_24481,N_24550);
or UO_407 (O_407,N_24890,N_24641);
xnor UO_408 (O_408,N_24798,N_24939);
or UO_409 (O_409,N_24500,N_24733);
or UO_410 (O_410,N_24799,N_24725);
xor UO_411 (O_411,N_24905,N_24421);
nor UO_412 (O_412,N_24562,N_24537);
nor UO_413 (O_413,N_24666,N_24434);
or UO_414 (O_414,N_24445,N_24626);
or UO_415 (O_415,N_24975,N_24529);
or UO_416 (O_416,N_24667,N_24513);
xor UO_417 (O_417,N_24936,N_24606);
nor UO_418 (O_418,N_24603,N_24393);
or UO_419 (O_419,N_24632,N_24942);
and UO_420 (O_420,N_24941,N_24397);
and UO_421 (O_421,N_24436,N_24841);
xor UO_422 (O_422,N_24546,N_24895);
xnor UO_423 (O_423,N_24827,N_24525);
and UO_424 (O_424,N_24919,N_24528);
or UO_425 (O_425,N_24580,N_24712);
nand UO_426 (O_426,N_24964,N_24767);
xor UO_427 (O_427,N_24571,N_24601);
xor UO_428 (O_428,N_24644,N_24826);
nor UO_429 (O_429,N_24435,N_24776);
nor UO_430 (O_430,N_24867,N_24837);
xnor UO_431 (O_431,N_24482,N_24816);
nand UO_432 (O_432,N_24760,N_24672);
nor UO_433 (O_433,N_24572,N_24508);
or UO_434 (O_434,N_24419,N_24841);
nand UO_435 (O_435,N_24540,N_24671);
and UO_436 (O_436,N_24936,N_24552);
nor UO_437 (O_437,N_24926,N_24399);
nand UO_438 (O_438,N_24390,N_24889);
nand UO_439 (O_439,N_24439,N_24939);
nand UO_440 (O_440,N_24687,N_24429);
nand UO_441 (O_441,N_24875,N_24673);
and UO_442 (O_442,N_24862,N_24637);
or UO_443 (O_443,N_24515,N_24773);
nand UO_444 (O_444,N_24913,N_24729);
or UO_445 (O_445,N_24801,N_24405);
nand UO_446 (O_446,N_24476,N_24824);
xor UO_447 (O_447,N_24575,N_24846);
or UO_448 (O_448,N_24384,N_24441);
xor UO_449 (O_449,N_24677,N_24412);
nor UO_450 (O_450,N_24851,N_24933);
or UO_451 (O_451,N_24385,N_24397);
nor UO_452 (O_452,N_24713,N_24628);
and UO_453 (O_453,N_24574,N_24671);
and UO_454 (O_454,N_24876,N_24777);
nand UO_455 (O_455,N_24396,N_24432);
or UO_456 (O_456,N_24912,N_24473);
and UO_457 (O_457,N_24521,N_24883);
or UO_458 (O_458,N_24577,N_24579);
and UO_459 (O_459,N_24976,N_24458);
nor UO_460 (O_460,N_24981,N_24760);
nor UO_461 (O_461,N_24466,N_24424);
nand UO_462 (O_462,N_24983,N_24911);
nor UO_463 (O_463,N_24797,N_24396);
or UO_464 (O_464,N_24848,N_24570);
xnor UO_465 (O_465,N_24774,N_24967);
or UO_466 (O_466,N_24483,N_24892);
xnor UO_467 (O_467,N_24741,N_24458);
nor UO_468 (O_468,N_24668,N_24712);
and UO_469 (O_469,N_24647,N_24987);
and UO_470 (O_470,N_24503,N_24479);
nor UO_471 (O_471,N_24970,N_24994);
xnor UO_472 (O_472,N_24827,N_24970);
xor UO_473 (O_473,N_24981,N_24561);
or UO_474 (O_474,N_24671,N_24430);
or UO_475 (O_475,N_24544,N_24652);
nand UO_476 (O_476,N_24622,N_24750);
nand UO_477 (O_477,N_24789,N_24818);
nand UO_478 (O_478,N_24979,N_24452);
and UO_479 (O_479,N_24814,N_24392);
nor UO_480 (O_480,N_24950,N_24975);
and UO_481 (O_481,N_24852,N_24989);
nand UO_482 (O_482,N_24802,N_24467);
nand UO_483 (O_483,N_24586,N_24489);
xor UO_484 (O_484,N_24952,N_24429);
xnor UO_485 (O_485,N_24625,N_24903);
nand UO_486 (O_486,N_24486,N_24477);
and UO_487 (O_487,N_24899,N_24496);
nor UO_488 (O_488,N_24963,N_24798);
and UO_489 (O_489,N_24782,N_24597);
or UO_490 (O_490,N_24660,N_24962);
or UO_491 (O_491,N_24910,N_24593);
and UO_492 (O_492,N_24993,N_24807);
or UO_493 (O_493,N_24851,N_24534);
or UO_494 (O_494,N_24663,N_24783);
or UO_495 (O_495,N_24760,N_24611);
nor UO_496 (O_496,N_24546,N_24754);
nor UO_497 (O_497,N_24805,N_24520);
xor UO_498 (O_498,N_24998,N_24578);
and UO_499 (O_499,N_24807,N_24638);
nor UO_500 (O_500,N_24460,N_24734);
nor UO_501 (O_501,N_24627,N_24753);
nor UO_502 (O_502,N_24805,N_24725);
nor UO_503 (O_503,N_24862,N_24676);
and UO_504 (O_504,N_24920,N_24580);
nand UO_505 (O_505,N_24745,N_24442);
and UO_506 (O_506,N_24995,N_24427);
nor UO_507 (O_507,N_24663,N_24981);
xnor UO_508 (O_508,N_24828,N_24963);
nor UO_509 (O_509,N_24866,N_24710);
or UO_510 (O_510,N_24459,N_24697);
nand UO_511 (O_511,N_24905,N_24539);
and UO_512 (O_512,N_24829,N_24830);
and UO_513 (O_513,N_24957,N_24921);
nor UO_514 (O_514,N_24990,N_24405);
and UO_515 (O_515,N_24448,N_24431);
xnor UO_516 (O_516,N_24439,N_24954);
xor UO_517 (O_517,N_24920,N_24595);
nand UO_518 (O_518,N_24408,N_24384);
nor UO_519 (O_519,N_24674,N_24739);
xor UO_520 (O_520,N_24896,N_24613);
xnor UO_521 (O_521,N_24443,N_24787);
or UO_522 (O_522,N_24811,N_24742);
nand UO_523 (O_523,N_24419,N_24932);
or UO_524 (O_524,N_24906,N_24668);
nand UO_525 (O_525,N_24535,N_24798);
xnor UO_526 (O_526,N_24634,N_24761);
nor UO_527 (O_527,N_24381,N_24614);
and UO_528 (O_528,N_24938,N_24445);
nand UO_529 (O_529,N_24936,N_24545);
or UO_530 (O_530,N_24451,N_24860);
xnor UO_531 (O_531,N_24615,N_24881);
nand UO_532 (O_532,N_24946,N_24780);
nand UO_533 (O_533,N_24552,N_24646);
or UO_534 (O_534,N_24777,N_24680);
xor UO_535 (O_535,N_24444,N_24954);
nor UO_536 (O_536,N_24460,N_24556);
and UO_537 (O_537,N_24838,N_24526);
xor UO_538 (O_538,N_24846,N_24869);
or UO_539 (O_539,N_24696,N_24626);
xor UO_540 (O_540,N_24765,N_24834);
nor UO_541 (O_541,N_24618,N_24722);
or UO_542 (O_542,N_24852,N_24433);
nand UO_543 (O_543,N_24762,N_24999);
nand UO_544 (O_544,N_24605,N_24889);
nor UO_545 (O_545,N_24888,N_24549);
xor UO_546 (O_546,N_24422,N_24507);
or UO_547 (O_547,N_24569,N_24921);
or UO_548 (O_548,N_24916,N_24989);
and UO_549 (O_549,N_24470,N_24809);
nand UO_550 (O_550,N_24432,N_24960);
xor UO_551 (O_551,N_24792,N_24730);
nor UO_552 (O_552,N_24408,N_24964);
and UO_553 (O_553,N_24784,N_24814);
nor UO_554 (O_554,N_24792,N_24994);
or UO_555 (O_555,N_24837,N_24480);
or UO_556 (O_556,N_24937,N_24740);
and UO_557 (O_557,N_24704,N_24629);
xor UO_558 (O_558,N_24948,N_24583);
nand UO_559 (O_559,N_24767,N_24466);
nand UO_560 (O_560,N_24394,N_24415);
and UO_561 (O_561,N_24999,N_24675);
nor UO_562 (O_562,N_24488,N_24968);
and UO_563 (O_563,N_24929,N_24375);
xor UO_564 (O_564,N_24624,N_24782);
or UO_565 (O_565,N_24873,N_24568);
or UO_566 (O_566,N_24465,N_24381);
xnor UO_567 (O_567,N_24960,N_24713);
and UO_568 (O_568,N_24390,N_24554);
nand UO_569 (O_569,N_24762,N_24884);
nand UO_570 (O_570,N_24830,N_24532);
nand UO_571 (O_571,N_24381,N_24705);
nor UO_572 (O_572,N_24943,N_24579);
or UO_573 (O_573,N_24827,N_24715);
or UO_574 (O_574,N_24771,N_24825);
or UO_575 (O_575,N_24725,N_24573);
or UO_576 (O_576,N_24877,N_24712);
or UO_577 (O_577,N_24701,N_24832);
nor UO_578 (O_578,N_24423,N_24988);
or UO_579 (O_579,N_24872,N_24581);
nor UO_580 (O_580,N_24663,N_24964);
nand UO_581 (O_581,N_24540,N_24969);
nor UO_582 (O_582,N_24746,N_24758);
nor UO_583 (O_583,N_24635,N_24770);
and UO_584 (O_584,N_24810,N_24890);
xor UO_585 (O_585,N_24992,N_24559);
xnor UO_586 (O_586,N_24940,N_24971);
xor UO_587 (O_587,N_24847,N_24651);
nor UO_588 (O_588,N_24863,N_24469);
xor UO_589 (O_589,N_24427,N_24625);
nand UO_590 (O_590,N_24817,N_24441);
nand UO_591 (O_591,N_24609,N_24455);
nand UO_592 (O_592,N_24965,N_24949);
xor UO_593 (O_593,N_24908,N_24793);
nor UO_594 (O_594,N_24565,N_24698);
nand UO_595 (O_595,N_24787,N_24894);
nand UO_596 (O_596,N_24712,N_24632);
xnor UO_597 (O_597,N_24528,N_24616);
xor UO_598 (O_598,N_24878,N_24477);
nor UO_599 (O_599,N_24960,N_24729);
and UO_600 (O_600,N_24527,N_24660);
nand UO_601 (O_601,N_24617,N_24381);
nor UO_602 (O_602,N_24485,N_24961);
or UO_603 (O_603,N_24677,N_24989);
nor UO_604 (O_604,N_24733,N_24565);
and UO_605 (O_605,N_24604,N_24929);
nand UO_606 (O_606,N_24815,N_24428);
xnor UO_607 (O_607,N_24809,N_24736);
and UO_608 (O_608,N_24988,N_24974);
nor UO_609 (O_609,N_24605,N_24478);
nor UO_610 (O_610,N_24698,N_24935);
xor UO_611 (O_611,N_24965,N_24534);
nand UO_612 (O_612,N_24795,N_24609);
nor UO_613 (O_613,N_24937,N_24855);
and UO_614 (O_614,N_24822,N_24775);
nand UO_615 (O_615,N_24634,N_24742);
nor UO_616 (O_616,N_24576,N_24820);
xor UO_617 (O_617,N_24443,N_24467);
xnor UO_618 (O_618,N_24886,N_24538);
nand UO_619 (O_619,N_24941,N_24775);
or UO_620 (O_620,N_24951,N_24973);
nand UO_621 (O_621,N_24979,N_24428);
and UO_622 (O_622,N_24715,N_24468);
and UO_623 (O_623,N_24656,N_24649);
or UO_624 (O_624,N_24734,N_24526);
and UO_625 (O_625,N_24913,N_24739);
nor UO_626 (O_626,N_24620,N_24748);
xor UO_627 (O_627,N_24677,N_24859);
and UO_628 (O_628,N_24925,N_24736);
or UO_629 (O_629,N_24947,N_24995);
and UO_630 (O_630,N_24410,N_24925);
nor UO_631 (O_631,N_24967,N_24935);
and UO_632 (O_632,N_24658,N_24735);
and UO_633 (O_633,N_24546,N_24925);
nor UO_634 (O_634,N_24740,N_24395);
nand UO_635 (O_635,N_24667,N_24680);
nor UO_636 (O_636,N_24855,N_24580);
or UO_637 (O_637,N_24631,N_24692);
nand UO_638 (O_638,N_24700,N_24632);
nand UO_639 (O_639,N_24763,N_24598);
nand UO_640 (O_640,N_24682,N_24737);
or UO_641 (O_641,N_24480,N_24712);
or UO_642 (O_642,N_24512,N_24557);
nor UO_643 (O_643,N_24552,N_24735);
xor UO_644 (O_644,N_24669,N_24692);
or UO_645 (O_645,N_24417,N_24652);
xnor UO_646 (O_646,N_24413,N_24931);
xor UO_647 (O_647,N_24812,N_24679);
nand UO_648 (O_648,N_24543,N_24727);
nand UO_649 (O_649,N_24847,N_24815);
and UO_650 (O_650,N_24492,N_24993);
xnor UO_651 (O_651,N_24974,N_24671);
and UO_652 (O_652,N_24851,N_24890);
nor UO_653 (O_653,N_24990,N_24835);
xor UO_654 (O_654,N_24776,N_24827);
xnor UO_655 (O_655,N_24478,N_24422);
nor UO_656 (O_656,N_24886,N_24922);
xor UO_657 (O_657,N_24962,N_24728);
nor UO_658 (O_658,N_24697,N_24658);
or UO_659 (O_659,N_24970,N_24419);
or UO_660 (O_660,N_24510,N_24408);
xnor UO_661 (O_661,N_24721,N_24772);
and UO_662 (O_662,N_24970,N_24394);
nand UO_663 (O_663,N_24521,N_24451);
xor UO_664 (O_664,N_24762,N_24714);
and UO_665 (O_665,N_24481,N_24598);
xnor UO_666 (O_666,N_24529,N_24646);
nand UO_667 (O_667,N_24654,N_24850);
nor UO_668 (O_668,N_24951,N_24739);
or UO_669 (O_669,N_24512,N_24973);
nor UO_670 (O_670,N_24584,N_24814);
and UO_671 (O_671,N_24386,N_24777);
or UO_672 (O_672,N_24385,N_24971);
or UO_673 (O_673,N_24432,N_24939);
xnor UO_674 (O_674,N_24917,N_24517);
or UO_675 (O_675,N_24614,N_24455);
nand UO_676 (O_676,N_24941,N_24544);
nor UO_677 (O_677,N_24781,N_24966);
and UO_678 (O_678,N_24987,N_24567);
and UO_679 (O_679,N_24989,N_24808);
and UO_680 (O_680,N_24387,N_24986);
or UO_681 (O_681,N_24966,N_24949);
or UO_682 (O_682,N_24494,N_24402);
nand UO_683 (O_683,N_24852,N_24465);
xor UO_684 (O_684,N_24602,N_24580);
and UO_685 (O_685,N_24693,N_24815);
and UO_686 (O_686,N_24805,N_24584);
nand UO_687 (O_687,N_24918,N_24817);
or UO_688 (O_688,N_24853,N_24722);
xor UO_689 (O_689,N_24585,N_24659);
nor UO_690 (O_690,N_24912,N_24538);
nor UO_691 (O_691,N_24658,N_24745);
or UO_692 (O_692,N_24427,N_24472);
nor UO_693 (O_693,N_24924,N_24903);
nor UO_694 (O_694,N_24977,N_24997);
xor UO_695 (O_695,N_24510,N_24749);
nor UO_696 (O_696,N_24412,N_24484);
and UO_697 (O_697,N_24511,N_24720);
xnor UO_698 (O_698,N_24826,N_24577);
xor UO_699 (O_699,N_24858,N_24468);
nand UO_700 (O_700,N_24632,N_24913);
and UO_701 (O_701,N_24418,N_24588);
nor UO_702 (O_702,N_24443,N_24733);
nand UO_703 (O_703,N_24380,N_24940);
nand UO_704 (O_704,N_24915,N_24563);
nor UO_705 (O_705,N_24694,N_24637);
or UO_706 (O_706,N_24984,N_24455);
nand UO_707 (O_707,N_24452,N_24588);
and UO_708 (O_708,N_24684,N_24416);
xor UO_709 (O_709,N_24525,N_24773);
nand UO_710 (O_710,N_24567,N_24752);
and UO_711 (O_711,N_24632,N_24588);
and UO_712 (O_712,N_24863,N_24472);
xnor UO_713 (O_713,N_24719,N_24811);
nand UO_714 (O_714,N_24392,N_24868);
and UO_715 (O_715,N_24804,N_24820);
nand UO_716 (O_716,N_24498,N_24934);
nand UO_717 (O_717,N_24418,N_24758);
xor UO_718 (O_718,N_24889,N_24584);
nor UO_719 (O_719,N_24550,N_24576);
xor UO_720 (O_720,N_24970,N_24917);
and UO_721 (O_721,N_24449,N_24791);
and UO_722 (O_722,N_24695,N_24919);
nand UO_723 (O_723,N_24822,N_24782);
nor UO_724 (O_724,N_24651,N_24998);
xnor UO_725 (O_725,N_24703,N_24704);
and UO_726 (O_726,N_24696,N_24450);
or UO_727 (O_727,N_24609,N_24413);
and UO_728 (O_728,N_24482,N_24573);
xor UO_729 (O_729,N_24562,N_24441);
nand UO_730 (O_730,N_24764,N_24590);
and UO_731 (O_731,N_24851,N_24645);
or UO_732 (O_732,N_24748,N_24649);
xnor UO_733 (O_733,N_24475,N_24890);
nand UO_734 (O_734,N_24544,N_24934);
and UO_735 (O_735,N_24503,N_24793);
or UO_736 (O_736,N_24416,N_24697);
or UO_737 (O_737,N_24823,N_24777);
and UO_738 (O_738,N_24943,N_24808);
nor UO_739 (O_739,N_24415,N_24590);
and UO_740 (O_740,N_24464,N_24840);
nor UO_741 (O_741,N_24588,N_24430);
or UO_742 (O_742,N_24406,N_24933);
xnor UO_743 (O_743,N_24594,N_24558);
or UO_744 (O_744,N_24971,N_24709);
nand UO_745 (O_745,N_24661,N_24595);
nor UO_746 (O_746,N_24498,N_24985);
nor UO_747 (O_747,N_24424,N_24948);
and UO_748 (O_748,N_24883,N_24580);
nand UO_749 (O_749,N_24428,N_24461);
nand UO_750 (O_750,N_24610,N_24981);
nor UO_751 (O_751,N_24773,N_24434);
nand UO_752 (O_752,N_24584,N_24843);
nor UO_753 (O_753,N_24957,N_24768);
nand UO_754 (O_754,N_24412,N_24699);
xnor UO_755 (O_755,N_24618,N_24668);
or UO_756 (O_756,N_24926,N_24455);
nor UO_757 (O_757,N_24550,N_24411);
and UO_758 (O_758,N_24383,N_24574);
and UO_759 (O_759,N_24481,N_24663);
xnor UO_760 (O_760,N_24442,N_24866);
nor UO_761 (O_761,N_24831,N_24518);
or UO_762 (O_762,N_24769,N_24625);
and UO_763 (O_763,N_24951,N_24418);
and UO_764 (O_764,N_24985,N_24796);
nor UO_765 (O_765,N_24903,N_24600);
nor UO_766 (O_766,N_24490,N_24551);
xnor UO_767 (O_767,N_24685,N_24564);
xnor UO_768 (O_768,N_24588,N_24898);
nor UO_769 (O_769,N_24881,N_24710);
nand UO_770 (O_770,N_24518,N_24822);
nand UO_771 (O_771,N_24474,N_24567);
nor UO_772 (O_772,N_24621,N_24875);
nand UO_773 (O_773,N_24646,N_24875);
nand UO_774 (O_774,N_24459,N_24968);
or UO_775 (O_775,N_24631,N_24916);
or UO_776 (O_776,N_24658,N_24571);
or UO_777 (O_777,N_24666,N_24687);
or UO_778 (O_778,N_24796,N_24739);
or UO_779 (O_779,N_24753,N_24732);
nand UO_780 (O_780,N_24771,N_24767);
xnor UO_781 (O_781,N_24672,N_24923);
and UO_782 (O_782,N_24536,N_24980);
or UO_783 (O_783,N_24476,N_24861);
and UO_784 (O_784,N_24918,N_24501);
nor UO_785 (O_785,N_24782,N_24518);
or UO_786 (O_786,N_24851,N_24538);
nor UO_787 (O_787,N_24746,N_24774);
nand UO_788 (O_788,N_24917,N_24492);
and UO_789 (O_789,N_24973,N_24926);
and UO_790 (O_790,N_24817,N_24708);
nor UO_791 (O_791,N_24517,N_24455);
nand UO_792 (O_792,N_24999,N_24955);
or UO_793 (O_793,N_24966,N_24422);
nand UO_794 (O_794,N_24378,N_24563);
or UO_795 (O_795,N_24877,N_24799);
or UO_796 (O_796,N_24719,N_24445);
nand UO_797 (O_797,N_24833,N_24508);
or UO_798 (O_798,N_24783,N_24605);
and UO_799 (O_799,N_24385,N_24871);
nand UO_800 (O_800,N_24999,N_24779);
xnor UO_801 (O_801,N_24656,N_24757);
and UO_802 (O_802,N_24715,N_24960);
nand UO_803 (O_803,N_24390,N_24912);
nor UO_804 (O_804,N_24402,N_24834);
nand UO_805 (O_805,N_24972,N_24770);
or UO_806 (O_806,N_24985,N_24409);
or UO_807 (O_807,N_24840,N_24825);
or UO_808 (O_808,N_24401,N_24798);
xor UO_809 (O_809,N_24896,N_24927);
nand UO_810 (O_810,N_24624,N_24573);
and UO_811 (O_811,N_24467,N_24515);
and UO_812 (O_812,N_24714,N_24435);
xor UO_813 (O_813,N_24885,N_24919);
xor UO_814 (O_814,N_24823,N_24888);
and UO_815 (O_815,N_24768,N_24692);
nand UO_816 (O_816,N_24657,N_24803);
nor UO_817 (O_817,N_24923,N_24894);
nand UO_818 (O_818,N_24723,N_24620);
and UO_819 (O_819,N_24936,N_24493);
xor UO_820 (O_820,N_24858,N_24960);
nand UO_821 (O_821,N_24859,N_24877);
nor UO_822 (O_822,N_24712,N_24399);
or UO_823 (O_823,N_24487,N_24507);
xor UO_824 (O_824,N_24407,N_24765);
and UO_825 (O_825,N_24418,N_24832);
or UO_826 (O_826,N_24837,N_24714);
or UO_827 (O_827,N_24827,N_24538);
or UO_828 (O_828,N_24896,N_24678);
and UO_829 (O_829,N_24686,N_24856);
xor UO_830 (O_830,N_24565,N_24928);
or UO_831 (O_831,N_24375,N_24612);
or UO_832 (O_832,N_24725,N_24403);
nor UO_833 (O_833,N_24432,N_24620);
nor UO_834 (O_834,N_24560,N_24588);
nand UO_835 (O_835,N_24883,N_24613);
or UO_836 (O_836,N_24705,N_24939);
or UO_837 (O_837,N_24782,N_24576);
nand UO_838 (O_838,N_24869,N_24939);
or UO_839 (O_839,N_24383,N_24942);
nor UO_840 (O_840,N_24770,N_24450);
nand UO_841 (O_841,N_24573,N_24603);
nor UO_842 (O_842,N_24943,N_24428);
xnor UO_843 (O_843,N_24543,N_24689);
xnor UO_844 (O_844,N_24693,N_24625);
nor UO_845 (O_845,N_24788,N_24789);
xnor UO_846 (O_846,N_24452,N_24600);
nand UO_847 (O_847,N_24580,N_24549);
nand UO_848 (O_848,N_24577,N_24700);
and UO_849 (O_849,N_24565,N_24482);
and UO_850 (O_850,N_24569,N_24476);
and UO_851 (O_851,N_24447,N_24918);
and UO_852 (O_852,N_24898,N_24862);
xnor UO_853 (O_853,N_24552,N_24791);
and UO_854 (O_854,N_24664,N_24974);
xor UO_855 (O_855,N_24806,N_24458);
or UO_856 (O_856,N_24995,N_24826);
nor UO_857 (O_857,N_24527,N_24891);
nor UO_858 (O_858,N_24697,N_24681);
and UO_859 (O_859,N_24984,N_24616);
xor UO_860 (O_860,N_24431,N_24685);
nor UO_861 (O_861,N_24441,N_24552);
nor UO_862 (O_862,N_24531,N_24906);
xnor UO_863 (O_863,N_24746,N_24760);
and UO_864 (O_864,N_24579,N_24489);
or UO_865 (O_865,N_24595,N_24727);
or UO_866 (O_866,N_24418,N_24585);
xnor UO_867 (O_867,N_24870,N_24804);
and UO_868 (O_868,N_24922,N_24847);
nand UO_869 (O_869,N_24403,N_24689);
xor UO_870 (O_870,N_24588,N_24837);
or UO_871 (O_871,N_24380,N_24388);
nand UO_872 (O_872,N_24511,N_24855);
nor UO_873 (O_873,N_24786,N_24609);
or UO_874 (O_874,N_24857,N_24709);
or UO_875 (O_875,N_24392,N_24702);
or UO_876 (O_876,N_24758,N_24414);
xnor UO_877 (O_877,N_24776,N_24814);
or UO_878 (O_878,N_24732,N_24525);
nand UO_879 (O_879,N_24885,N_24415);
xnor UO_880 (O_880,N_24476,N_24585);
or UO_881 (O_881,N_24557,N_24440);
or UO_882 (O_882,N_24386,N_24948);
or UO_883 (O_883,N_24627,N_24723);
and UO_884 (O_884,N_24751,N_24994);
or UO_885 (O_885,N_24810,N_24635);
nor UO_886 (O_886,N_24748,N_24723);
nand UO_887 (O_887,N_24654,N_24872);
xnor UO_888 (O_888,N_24454,N_24576);
xor UO_889 (O_889,N_24387,N_24471);
nand UO_890 (O_890,N_24408,N_24732);
or UO_891 (O_891,N_24416,N_24973);
nand UO_892 (O_892,N_24867,N_24438);
nor UO_893 (O_893,N_24584,N_24777);
or UO_894 (O_894,N_24495,N_24758);
nor UO_895 (O_895,N_24393,N_24476);
and UO_896 (O_896,N_24893,N_24920);
and UO_897 (O_897,N_24712,N_24469);
nor UO_898 (O_898,N_24846,N_24873);
nor UO_899 (O_899,N_24540,N_24935);
and UO_900 (O_900,N_24799,N_24871);
nand UO_901 (O_901,N_24872,N_24917);
nor UO_902 (O_902,N_24489,N_24768);
or UO_903 (O_903,N_24604,N_24674);
xnor UO_904 (O_904,N_24732,N_24701);
and UO_905 (O_905,N_24575,N_24393);
or UO_906 (O_906,N_24483,N_24969);
nor UO_907 (O_907,N_24719,N_24898);
xor UO_908 (O_908,N_24640,N_24932);
nand UO_909 (O_909,N_24853,N_24549);
nand UO_910 (O_910,N_24710,N_24474);
or UO_911 (O_911,N_24763,N_24540);
xor UO_912 (O_912,N_24477,N_24434);
nor UO_913 (O_913,N_24890,N_24880);
or UO_914 (O_914,N_24499,N_24853);
nor UO_915 (O_915,N_24553,N_24987);
xor UO_916 (O_916,N_24482,N_24657);
nand UO_917 (O_917,N_24899,N_24523);
and UO_918 (O_918,N_24767,N_24517);
and UO_919 (O_919,N_24457,N_24431);
and UO_920 (O_920,N_24391,N_24789);
or UO_921 (O_921,N_24476,N_24454);
nor UO_922 (O_922,N_24654,N_24661);
nor UO_923 (O_923,N_24776,N_24647);
xnor UO_924 (O_924,N_24681,N_24411);
nand UO_925 (O_925,N_24446,N_24759);
nor UO_926 (O_926,N_24459,N_24681);
and UO_927 (O_927,N_24714,N_24697);
or UO_928 (O_928,N_24902,N_24980);
or UO_929 (O_929,N_24878,N_24896);
and UO_930 (O_930,N_24809,N_24455);
and UO_931 (O_931,N_24926,N_24433);
or UO_932 (O_932,N_24949,N_24744);
xnor UO_933 (O_933,N_24730,N_24877);
xnor UO_934 (O_934,N_24521,N_24945);
xor UO_935 (O_935,N_24376,N_24847);
or UO_936 (O_936,N_24540,N_24502);
nand UO_937 (O_937,N_24709,N_24831);
or UO_938 (O_938,N_24401,N_24514);
and UO_939 (O_939,N_24518,N_24638);
nor UO_940 (O_940,N_24393,N_24566);
or UO_941 (O_941,N_24616,N_24678);
or UO_942 (O_942,N_24522,N_24931);
xor UO_943 (O_943,N_24863,N_24710);
and UO_944 (O_944,N_24801,N_24541);
or UO_945 (O_945,N_24954,N_24806);
nand UO_946 (O_946,N_24836,N_24738);
xor UO_947 (O_947,N_24501,N_24766);
nand UO_948 (O_948,N_24442,N_24883);
or UO_949 (O_949,N_24921,N_24688);
nand UO_950 (O_950,N_24566,N_24916);
nand UO_951 (O_951,N_24985,N_24494);
nor UO_952 (O_952,N_24835,N_24377);
and UO_953 (O_953,N_24436,N_24693);
nand UO_954 (O_954,N_24920,N_24695);
xor UO_955 (O_955,N_24913,N_24404);
nand UO_956 (O_956,N_24481,N_24754);
nor UO_957 (O_957,N_24964,N_24888);
and UO_958 (O_958,N_24864,N_24650);
or UO_959 (O_959,N_24715,N_24881);
nor UO_960 (O_960,N_24788,N_24753);
and UO_961 (O_961,N_24986,N_24398);
and UO_962 (O_962,N_24692,N_24503);
nor UO_963 (O_963,N_24854,N_24791);
or UO_964 (O_964,N_24643,N_24605);
xnor UO_965 (O_965,N_24913,N_24388);
nor UO_966 (O_966,N_24391,N_24770);
xnor UO_967 (O_967,N_24632,N_24648);
or UO_968 (O_968,N_24694,N_24761);
xnor UO_969 (O_969,N_24766,N_24911);
xnor UO_970 (O_970,N_24805,N_24585);
nor UO_971 (O_971,N_24640,N_24692);
nor UO_972 (O_972,N_24764,N_24401);
nand UO_973 (O_973,N_24878,N_24463);
nor UO_974 (O_974,N_24835,N_24507);
nand UO_975 (O_975,N_24452,N_24952);
and UO_976 (O_976,N_24946,N_24730);
nor UO_977 (O_977,N_24743,N_24648);
and UO_978 (O_978,N_24519,N_24937);
nor UO_979 (O_979,N_24439,N_24627);
xnor UO_980 (O_980,N_24995,N_24402);
xnor UO_981 (O_981,N_24547,N_24577);
nand UO_982 (O_982,N_24805,N_24763);
and UO_983 (O_983,N_24428,N_24909);
xor UO_984 (O_984,N_24656,N_24402);
xnor UO_985 (O_985,N_24420,N_24629);
or UO_986 (O_986,N_24451,N_24547);
xnor UO_987 (O_987,N_24604,N_24854);
nand UO_988 (O_988,N_24462,N_24887);
xnor UO_989 (O_989,N_24473,N_24773);
nand UO_990 (O_990,N_24885,N_24391);
and UO_991 (O_991,N_24491,N_24681);
nor UO_992 (O_992,N_24933,N_24705);
xor UO_993 (O_993,N_24904,N_24555);
and UO_994 (O_994,N_24699,N_24437);
xnor UO_995 (O_995,N_24879,N_24412);
and UO_996 (O_996,N_24899,N_24902);
and UO_997 (O_997,N_24882,N_24560);
xnor UO_998 (O_998,N_24901,N_24801);
and UO_999 (O_999,N_24519,N_24643);
and UO_1000 (O_1000,N_24541,N_24537);
nand UO_1001 (O_1001,N_24728,N_24380);
or UO_1002 (O_1002,N_24933,N_24601);
nor UO_1003 (O_1003,N_24438,N_24714);
nand UO_1004 (O_1004,N_24687,N_24888);
nand UO_1005 (O_1005,N_24501,N_24588);
xor UO_1006 (O_1006,N_24753,N_24915);
or UO_1007 (O_1007,N_24858,N_24709);
or UO_1008 (O_1008,N_24879,N_24975);
nand UO_1009 (O_1009,N_24694,N_24801);
xnor UO_1010 (O_1010,N_24586,N_24456);
nand UO_1011 (O_1011,N_24534,N_24893);
nand UO_1012 (O_1012,N_24380,N_24977);
or UO_1013 (O_1013,N_24888,N_24392);
xor UO_1014 (O_1014,N_24640,N_24955);
nand UO_1015 (O_1015,N_24398,N_24758);
or UO_1016 (O_1016,N_24811,N_24558);
nand UO_1017 (O_1017,N_24760,N_24968);
nand UO_1018 (O_1018,N_24616,N_24525);
nor UO_1019 (O_1019,N_24410,N_24381);
xor UO_1020 (O_1020,N_24447,N_24916);
xor UO_1021 (O_1021,N_24564,N_24643);
and UO_1022 (O_1022,N_24991,N_24749);
nor UO_1023 (O_1023,N_24495,N_24668);
nor UO_1024 (O_1024,N_24557,N_24938);
or UO_1025 (O_1025,N_24556,N_24870);
or UO_1026 (O_1026,N_24879,N_24820);
nor UO_1027 (O_1027,N_24952,N_24718);
nor UO_1028 (O_1028,N_24869,N_24849);
nor UO_1029 (O_1029,N_24648,N_24380);
nand UO_1030 (O_1030,N_24575,N_24970);
nand UO_1031 (O_1031,N_24507,N_24421);
nand UO_1032 (O_1032,N_24697,N_24712);
xor UO_1033 (O_1033,N_24790,N_24792);
nand UO_1034 (O_1034,N_24973,N_24989);
and UO_1035 (O_1035,N_24859,N_24573);
nor UO_1036 (O_1036,N_24536,N_24480);
nand UO_1037 (O_1037,N_24830,N_24706);
nand UO_1038 (O_1038,N_24943,N_24873);
xor UO_1039 (O_1039,N_24938,N_24667);
or UO_1040 (O_1040,N_24538,N_24965);
or UO_1041 (O_1041,N_24874,N_24508);
or UO_1042 (O_1042,N_24966,N_24790);
xor UO_1043 (O_1043,N_24986,N_24759);
and UO_1044 (O_1044,N_24810,N_24723);
or UO_1045 (O_1045,N_24399,N_24867);
nor UO_1046 (O_1046,N_24595,N_24479);
or UO_1047 (O_1047,N_24786,N_24952);
nor UO_1048 (O_1048,N_24737,N_24816);
or UO_1049 (O_1049,N_24996,N_24448);
nor UO_1050 (O_1050,N_24827,N_24869);
nand UO_1051 (O_1051,N_24908,N_24870);
nand UO_1052 (O_1052,N_24848,N_24833);
nor UO_1053 (O_1053,N_24926,N_24965);
and UO_1054 (O_1054,N_24844,N_24842);
nand UO_1055 (O_1055,N_24850,N_24684);
nor UO_1056 (O_1056,N_24418,N_24408);
or UO_1057 (O_1057,N_24793,N_24711);
nand UO_1058 (O_1058,N_24852,N_24958);
and UO_1059 (O_1059,N_24588,N_24855);
nand UO_1060 (O_1060,N_24943,N_24831);
xnor UO_1061 (O_1061,N_24802,N_24481);
nand UO_1062 (O_1062,N_24624,N_24452);
nor UO_1063 (O_1063,N_24620,N_24608);
nand UO_1064 (O_1064,N_24596,N_24910);
xnor UO_1065 (O_1065,N_24702,N_24655);
nor UO_1066 (O_1066,N_24657,N_24739);
and UO_1067 (O_1067,N_24996,N_24821);
nor UO_1068 (O_1068,N_24772,N_24575);
and UO_1069 (O_1069,N_24440,N_24798);
or UO_1070 (O_1070,N_24864,N_24713);
nand UO_1071 (O_1071,N_24401,N_24810);
and UO_1072 (O_1072,N_24760,N_24390);
and UO_1073 (O_1073,N_24986,N_24623);
or UO_1074 (O_1074,N_24705,N_24753);
or UO_1075 (O_1075,N_24821,N_24978);
nand UO_1076 (O_1076,N_24914,N_24931);
and UO_1077 (O_1077,N_24937,N_24810);
nor UO_1078 (O_1078,N_24491,N_24553);
nor UO_1079 (O_1079,N_24926,N_24617);
and UO_1080 (O_1080,N_24815,N_24925);
nand UO_1081 (O_1081,N_24391,N_24584);
or UO_1082 (O_1082,N_24491,N_24625);
nand UO_1083 (O_1083,N_24668,N_24628);
or UO_1084 (O_1084,N_24393,N_24752);
and UO_1085 (O_1085,N_24743,N_24752);
and UO_1086 (O_1086,N_24943,N_24989);
or UO_1087 (O_1087,N_24650,N_24904);
xor UO_1088 (O_1088,N_24908,N_24889);
nor UO_1089 (O_1089,N_24465,N_24676);
nand UO_1090 (O_1090,N_24533,N_24597);
nor UO_1091 (O_1091,N_24822,N_24823);
or UO_1092 (O_1092,N_24795,N_24542);
xor UO_1093 (O_1093,N_24716,N_24534);
or UO_1094 (O_1094,N_24917,N_24503);
nor UO_1095 (O_1095,N_24644,N_24518);
and UO_1096 (O_1096,N_24401,N_24751);
nor UO_1097 (O_1097,N_24602,N_24512);
xnor UO_1098 (O_1098,N_24629,N_24886);
nand UO_1099 (O_1099,N_24585,N_24738);
and UO_1100 (O_1100,N_24619,N_24866);
nand UO_1101 (O_1101,N_24840,N_24627);
or UO_1102 (O_1102,N_24805,N_24604);
nand UO_1103 (O_1103,N_24585,N_24458);
xnor UO_1104 (O_1104,N_24467,N_24958);
or UO_1105 (O_1105,N_24596,N_24744);
and UO_1106 (O_1106,N_24679,N_24956);
xor UO_1107 (O_1107,N_24938,N_24758);
xnor UO_1108 (O_1108,N_24572,N_24859);
xor UO_1109 (O_1109,N_24710,N_24573);
nand UO_1110 (O_1110,N_24670,N_24919);
nor UO_1111 (O_1111,N_24667,N_24424);
nor UO_1112 (O_1112,N_24768,N_24797);
nor UO_1113 (O_1113,N_24910,N_24375);
or UO_1114 (O_1114,N_24848,N_24503);
nand UO_1115 (O_1115,N_24852,N_24741);
xor UO_1116 (O_1116,N_24662,N_24403);
and UO_1117 (O_1117,N_24996,N_24889);
nor UO_1118 (O_1118,N_24512,N_24491);
xnor UO_1119 (O_1119,N_24696,N_24828);
nand UO_1120 (O_1120,N_24640,N_24695);
nand UO_1121 (O_1121,N_24553,N_24530);
and UO_1122 (O_1122,N_24379,N_24858);
nor UO_1123 (O_1123,N_24903,N_24841);
nand UO_1124 (O_1124,N_24397,N_24903);
and UO_1125 (O_1125,N_24386,N_24435);
and UO_1126 (O_1126,N_24733,N_24482);
nor UO_1127 (O_1127,N_24878,N_24594);
nor UO_1128 (O_1128,N_24953,N_24824);
or UO_1129 (O_1129,N_24725,N_24638);
xnor UO_1130 (O_1130,N_24594,N_24940);
and UO_1131 (O_1131,N_24498,N_24732);
nor UO_1132 (O_1132,N_24435,N_24391);
and UO_1133 (O_1133,N_24436,N_24659);
nand UO_1134 (O_1134,N_24445,N_24848);
nor UO_1135 (O_1135,N_24991,N_24953);
xor UO_1136 (O_1136,N_24949,N_24684);
and UO_1137 (O_1137,N_24764,N_24643);
xnor UO_1138 (O_1138,N_24993,N_24449);
and UO_1139 (O_1139,N_24799,N_24598);
or UO_1140 (O_1140,N_24664,N_24655);
or UO_1141 (O_1141,N_24514,N_24457);
or UO_1142 (O_1142,N_24696,N_24765);
nand UO_1143 (O_1143,N_24656,N_24899);
nand UO_1144 (O_1144,N_24537,N_24674);
nor UO_1145 (O_1145,N_24552,N_24966);
or UO_1146 (O_1146,N_24955,N_24705);
nor UO_1147 (O_1147,N_24605,N_24496);
xnor UO_1148 (O_1148,N_24887,N_24963);
nand UO_1149 (O_1149,N_24813,N_24787);
xor UO_1150 (O_1150,N_24644,N_24592);
or UO_1151 (O_1151,N_24538,N_24704);
nand UO_1152 (O_1152,N_24801,N_24476);
and UO_1153 (O_1153,N_24652,N_24701);
xnor UO_1154 (O_1154,N_24436,N_24823);
nor UO_1155 (O_1155,N_24727,N_24925);
nor UO_1156 (O_1156,N_24662,N_24465);
xor UO_1157 (O_1157,N_24884,N_24540);
nor UO_1158 (O_1158,N_24417,N_24879);
xor UO_1159 (O_1159,N_24787,N_24425);
nor UO_1160 (O_1160,N_24697,N_24867);
or UO_1161 (O_1161,N_24851,N_24522);
nor UO_1162 (O_1162,N_24938,N_24809);
and UO_1163 (O_1163,N_24639,N_24750);
nand UO_1164 (O_1164,N_24805,N_24525);
or UO_1165 (O_1165,N_24932,N_24697);
xor UO_1166 (O_1166,N_24689,N_24889);
and UO_1167 (O_1167,N_24596,N_24521);
or UO_1168 (O_1168,N_24835,N_24869);
nand UO_1169 (O_1169,N_24684,N_24400);
or UO_1170 (O_1170,N_24392,N_24889);
nand UO_1171 (O_1171,N_24641,N_24709);
nand UO_1172 (O_1172,N_24487,N_24691);
xor UO_1173 (O_1173,N_24930,N_24413);
nor UO_1174 (O_1174,N_24709,N_24672);
and UO_1175 (O_1175,N_24588,N_24803);
xor UO_1176 (O_1176,N_24806,N_24570);
xor UO_1177 (O_1177,N_24698,N_24498);
xor UO_1178 (O_1178,N_24869,N_24588);
nand UO_1179 (O_1179,N_24419,N_24499);
nand UO_1180 (O_1180,N_24668,N_24517);
and UO_1181 (O_1181,N_24862,N_24804);
nand UO_1182 (O_1182,N_24914,N_24564);
xor UO_1183 (O_1183,N_24930,N_24792);
nor UO_1184 (O_1184,N_24727,N_24622);
xnor UO_1185 (O_1185,N_24982,N_24920);
or UO_1186 (O_1186,N_24620,N_24703);
and UO_1187 (O_1187,N_24629,N_24808);
xor UO_1188 (O_1188,N_24868,N_24632);
or UO_1189 (O_1189,N_24833,N_24554);
and UO_1190 (O_1190,N_24884,N_24924);
nor UO_1191 (O_1191,N_24572,N_24914);
and UO_1192 (O_1192,N_24851,N_24769);
or UO_1193 (O_1193,N_24395,N_24787);
nor UO_1194 (O_1194,N_24792,N_24668);
nand UO_1195 (O_1195,N_24917,N_24548);
nand UO_1196 (O_1196,N_24759,N_24632);
or UO_1197 (O_1197,N_24482,N_24823);
and UO_1198 (O_1198,N_24989,N_24669);
xor UO_1199 (O_1199,N_24820,N_24625);
nor UO_1200 (O_1200,N_24932,N_24405);
nand UO_1201 (O_1201,N_24413,N_24404);
and UO_1202 (O_1202,N_24808,N_24883);
nand UO_1203 (O_1203,N_24428,N_24779);
and UO_1204 (O_1204,N_24419,N_24665);
or UO_1205 (O_1205,N_24945,N_24996);
nand UO_1206 (O_1206,N_24598,N_24490);
and UO_1207 (O_1207,N_24384,N_24892);
xor UO_1208 (O_1208,N_24927,N_24747);
and UO_1209 (O_1209,N_24554,N_24701);
nor UO_1210 (O_1210,N_24836,N_24764);
xnor UO_1211 (O_1211,N_24665,N_24994);
or UO_1212 (O_1212,N_24698,N_24758);
nand UO_1213 (O_1213,N_24422,N_24624);
or UO_1214 (O_1214,N_24577,N_24667);
nor UO_1215 (O_1215,N_24789,N_24948);
and UO_1216 (O_1216,N_24978,N_24993);
xnor UO_1217 (O_1217,N_24927,N_24645);
and UO_1218 (O_1218,N_24708,N_24499);
nand UO_1219 (O_1219,N_24762,N_24727);
nand UO_1220 (O_1220,N_24518,N_24740);
nor UO_1221 (O_1221,N_24445,N_24552);
or UO_1222 (O_1222,N_24528,N_24830);
xor UO_1223 (O_1223,N_24521,N_24637);
or UO_1224 (O_1224,N_24493,N_24615);
nor UO_1225 (O_1225,N_24910,N_24377);
nand UO_1226 (O_1226,N_24385,N_24746);
and UO_1227 (O_1227,N_24575,N_24548);
xor UO_1228 (O_1228,N_24996,N_24872);
or UO_1229 (O_1229,N_24888,N_24777);
or UO_1230 (O_1230,N_24545,N_24645);
or UO_1231 (O_1231,N_24907,N_24534);
nand UO_1232 (O_1232,N_24618,N_24503);
nor UO_1233 (O_1233,N_24995,N_24550);
xnor UO_1234 (O_1234,N_24863,N_24955);
nor UO_1235 (O_1235,N_24806,N_24602);
nand UO_1236 (O_1236,N_24775,N_24764);
nand UO_1237 (O_1237,N_24870,N_24895);
nand UO_1238 (O_1238,N_24828,N_24733);
and UO_1239 (O_1239,N_24643,N_24840);
or UO_1240 (O_1240,N_24761,N_24393);
xnor UO_1241 (O_1241,N_24662,N_24996);
nor UO_1242 (O_1242,N_24409,N_24766);
nor UO_1243 (O_1243,N_24542,N_24946);
xor UO_1244 (O_1244,N_24951,N_24814);
xnor UO_1245 (O_1245,N_24604,N_24672);
xor UO_1246 (O_1246,N_24793,N_24847);
nor UO_1247 (O_1247,N_24980,N_24882);
nor UO_1248 (O_1248,N_24750,N_24936);
nor UO_1249 (O_1249,N_24739,N_24998);
and UO_1250 (O_1250,N_24995,N_24895);
xor UO_1251 (O_1251,N_24873,N_24435);
nand UO_1252 (O_1252,N_24592,N_24469);
xnor UO_1253 (O_1253,N_24587,N_24773);
nand UO_1254 (O_1254,N_24992,N_24920);
nand UO_1255 (O_1255,N_24579,N_24412);
or UO_1256 (O_1256,N_24726,N_24704);
and UO_1257 (O_1257,N_24849,N_24445);
xnor UO_1258 (O_1258,N_24706,N_24943);
xor UO_1259 (O_1259,N_24587,N_24696);
xnor UO_1260 (O_1260,N_24725,N_24921);
nor UO_1261 (O_1261,N_24749,N_24864);
xor UO_1262 (O_1262,N_24396,N_24810);
nand UO_1263 (O_1263,N_24442,N_24817);
or UO_1264 (O_1264,N_24385,N_24690);
nand UO_1265 (O_1265,N_24559,N_24743);
xor UO_1266 (O_1266,N_24906,N_24389);
or UO_1267 (O_1267,N_24565,N_24398);
nor UO_1268 (O_1268,N_24812,N_24913);
or UO_1269 (O_1269,N_24567,N_24530);
or UO_1270 (O_1270,N_24528,N_24922);
xor UO_1271 (O_1271,N_24963,N_24551);
and UO_1272 (O_1272,N_24714,N_24719);
and UO_1273 (O_1273,N_24970,N_24588);
xor UO_1274 (O_1274,N_24483,N_24461);
nor UO_1275 (O_1275,N_24886,N_24934);
or UO_1276 (O_1276,N_24525,N_24383);
or UO_1277 (O_1277,N_24877,N_24910);
and UO_1278 (O_1278,N_24505,N_24602);
xor UO_1279 (O_1279,N_24488,N_24869);
nor UO_1280 (O_1280,N_24420,N_24925);
nor UO_1281 (O_1281,N_24874,N_24634);
and UO_1282 (O_1282,N_24468,N_24937);
nand UO_1283 (O_1283,N_24566,N_24922);
and UO_1284 (O_1284,N_24777,N_24612);
and UO_1285 (O_1285,N_24398,N_24785);
nor UO_1286 (O_1286,N_24644,N_24885);
or UO_1287 (O_1287,N_24632,N_24524);
xnor UO_1288 (O_1288,N_24546,N_24511);
nand UO_1289 (O_1289,N_24999,N_24962);
nor UO_1290 (O_1290,N_24429,N_24889);
nand UO_1291 (O_1291,N_24926,N_24441);
nand UO_1292 (O_1292,N_24814,N_24870);
nand UO_1293 (O_1293,N_24979,N_24476);
nor UO_1294 (O_1294,N_24929,N_24870);
or UO_1295 (O_1295,N_24837,N_24555);
nand UO_1296 (O_1296,N_24756,N_24409);
and UO_1297 (O_1297,N_24901,N_24935);
xor UO_1298 (O_1298,N_24981,N_24688);
or UO_1299 (O_1299,N_24807,N_24489);
nand UO_1300 (O_1300,N_24583,N_24701);
xnor UO_1301 (O_1301,N_24565,N_24709);
and UO_1302 (O_1302,N_24457,N_24966);
or UO_1303 (O_1303,N_24492,N_24598);
nor UO_1304 (O_1304,N_24939,N_24632);
nor UO_1305 (O_1305,N_24838,N_24527);
nand UO_1306 (O_1306,N_24722,N_24946);
and UO_1307 (O_1307,N_24499,N_24563);
nor UO_1308 (O_1308,N_24917,N_24499);
and UO_1309 (O_1309,N_24606,N_24768);
or UO_1310 (O_1310,N_24418,N_24676);
and UO_1311 (O_1311,N_24490,N_24901);
xnor UO_1312 (O_1312,N_24858,N_24844);
and UO_1313 (O_1313,N_24498,N_24780);
and UO_1314 (O_1314,N_24705,N_24954);
nand UO_1315 (O_1315,N_24572,N_24604);
nand UO_1316 (O_1316,N_24542,N_24409);
and UO_1317 (O_1317,N_24708,N_24745);
nand UO_1318 (O_1318,N_24804,N_24661);
nor UO_1319 (O_1319,N_24573,N_24516);
nor UO_1320 (O_1320,N_24638,N_24522);
xor UO_1321 (O_1321,N_24741,N_24511);
or UO_1322 (O_1322,N_24508,N_24553);
nand UO_1323 (O_1323,N_24827,N_24711);
or UO_1324 (O_1324,N_24609,N_24546);
nand UO_1325 (O_1325,N_24858,N_24542);
nand UO_1326 (O_1326,N_24816,N_24868);
and UO_1327 (O_1327,N_24521,N_24460);
xor UO_1328 (O_1328,N_24960,N_24730);
nand UO_1329 (O_1329,N_24430,N_24636);
nor UO_1330 (O_1330,N_24425,N_24441);
and UO_1331 (O_1331,N_24987,N_24457);
or UO_1332 (O_1332,N_24647,N_24885);
or UO_1333 (O_1333,N_24544,N_24451);
xor UO_1334 (O_1334,N_24735,N_24567);
xnor UO_1335 (O_1335,N_24929,N_24595);
and UO_1336 (O_1336,N_24851,N_24659);
xnor UO_1337 (O_1337,N_24613,N_24819);
nor UO_1338 (O_1338,N_24678,N_24465);
nand UO_1339 (O_1339,N_24905,N_24400);
nand UO_1340 (O_1340,N_24734,N_24920);
xor UO_1341 (O_1341,N_24701,N_24388);
and UO_1342 (O_1342,N_24439,N_24673);
or UO_1343 (O_1343,N_24626,N_24897);
xnor UO_1344 (O_1344,N_24856,N_24644);
or UO_1345 (O_1345,N_24978,N_24624);
and UO_1346 (O_1346,N_24794,N_24666);
or UO_1347 (O_1347,N_24820,N_24945);
or UO_1348 (O_1348,N_24966,N_24993);
nand UO_1349 (O_1349,N_24984,N_24475);
nand UO_1350 (O_1350,N_24874,N_24621);
or UO_1351 (O_1351,N_24518,N_24497);
xor UO_1352 (O_1352,N_24431,N_24497);
xnor UO_1353 (O_1353,N_24679,N_24440);
and UO_1354 (O_1354,N_24411,N_24908);
nor UO_1355 (O_1355,N_24991,N_24426);
and UO_1356 (O_1356,N_24425,N_24628);
and UO_1357 (O_1357,N_24732,N_24727);
xor UO_1358 (O_1358,N_24549,N_24439);
or UO_1359 (O_1359,N_24794,N_24919);
and UO_1360 (O_1360,N_24391,N_24417);
xnor UO_1361 (O_1361,N_24398,N_24674);
nand UO_1362 (O_1362,N_24464,N_24717);
nand UO_1363 (O_1363,N_24918,N_24798);
nor UO_1364 (O_1364,N_24627,N_24722);
xor UO_1365 (O_1365,N_24569,N_24702);
nand UO_1366 (O_1366,N_24792,N_24863);
and UO_1367 (O_1367,N_24816,N_24418);
nor UO_1368 (O_1368,N_24492,N_24892);
nand UO_1369 (O_1369,N_24464,N_24489);
and UO_1370 (O_1370,N_24631,N_24516);
xor UO_1371 (O_1371,N_24390,N_24717);
nand UO_1372 (O_1372,N_24743,N_24698);
nor UO_1373 (O_1373,N_24546,N_24709);
or UO_1374 (O_1374,N_24452,N_24817);
nand UO_1375 (O_1375,N_24839,N_24657);
or UO_1376 (O_1376,N_24655,N_24813);
and UO_1377 (O_1377,N_24665,N_24885);
nand UO_1378 (O_1378,N_24800,N_24462);
and UO_1379 (O_1379,N_24554,N_24715);
or UO_1380 (O_1380,N_24657,N_24515);
xor UO_1381 (O_1381,N_24810,N_24925);
xnor UO_1382 (O_1382,N_24899,N_24597);
and UO_1383 (O_1383,N_24635,N_24604);
or UO_1384 (O_1384,N_24429,N_24920);
nor UO_1385 (O_1385,N_24384,N_24673);
nor UO_1386 (O_1386,N_24398,N_24883);
and UO_1387 (O_1387,N_24385,N_24698);
or UO_1388 (O_1388,N_24969,N_24870);
nor UO_1389 (O_1389,N_24651,N_24654);
or UO_1390 (O_1390,N_24540,N_24633);
xnor UO_1391 (O_1391,N_24759,N_24659);
nand UO_1392 (O_1392,N_24763,N_24967);
and UO_1393 (O_1393,N_24722,N_24498);
nand UO_1394 (O_1394,N_24545,N_24637);
xnor UO_1395 (O_1395,N_24758,N_24627);
and UO_1396 (O_1396,N_24645,N_24447);
and UO_1397 (O_1397,N_24656,N_24933);
nor UO_1398 (O_1398,N_24577,N_24959);
xor UO_1399 (O_1399,N_24952,N_24734);
nand UO_1400 (O_1400,N_24731,N_24862);
xor UO_1401 (O_1401,N_24493,N_24487);
or UO_1402 (O_1402,N_24496,N_24728);
or UO_1403 (O_1403,N_24962,N_24425);
and UO_1404 (O_1404,N_24954,N_24769);
and UO_1405 (O_1405,N_24999,N_24436);
and UO_1406 (O_1406,N_24378,N_24935);
or UO_1407 (O_1407,N_24413,N_24941);
nand UO_1408 (O_1408,N_24376,N_24392);
or UO_1409 (O_1409,N_24955,N_24477);
nand UO_1410 (O_1410,N_24920,N_24619);
nor UO_1411 (O_1411,N_24931,N_24809);
xor UO_1412 (O_1412,N_24756,N_24867);
nand UO_1413 (O_1413,N_24429,N_24385);
and UO_1414 (O_1414,N_24802,N_24907);
and UO_1415 (O_1415,N_24579,N_24965);
or UO_1416 (O_1416,N_24485,N_24457);
or UO_1417 (O_1417,N_24402,N_24622);
xnor UO_1418 (O_1418,N_24507,N_24916);
or UO_1419 (O_1419,N_24579,N_24465);
nand UO_1420 (O_1420,N_24430,N_24772);
xnor UO_1421 (O_1421,N_24535,N_24789);
xor UO_1422 (O_1422,N_24726,N_24378);
nand UO_1423 (O_1423,N_24850,N_24948);
xnor UO_1424 (O_1424,N_24527,N_24980);
or UO_1425 (O_1425,N_24757,N_24440);
xnor UO_1426 (O_1426,N_24423,N_24785);
xor UO_1427 (O_1427,N_24899,N_24618);
nand UO_1428 (O_1428,N_24648,N_24975);
nand UO_1429 (O_1429,N_24908,N_24819);
nand UO_1430 (O_1430,N_24527,N_24803);
and UO_1431 (O_1431,N_24822,N_24893);
nor UO_1432 (O_1432,N_24664,N_24414);
xor UO_1433 (O_1433,N_24703,N_24451);
nand UO_1434 (O_1434,N_24704,N_24723);
xnor UO_1435 (O_1435,N_24990,N_24470);
xnor UO_1436 (O_1436,N_24894,N_24560);
or UO_1437 (O_1437,N_24441,N_24979);
nand UO_1438 (O_1438,N_24461,N_24462);
nor UO_1439 (O_1439,N_24931,N_24545);
nand UO_1440 (O_1440,N_24675,N_24872);
xor UO_1441 (O_1441,N_24491,N_24470);
nor UO_1442 (O_1442,N_24924,N_24404);
nand UO_1443 (O_1443,N_24938,N_24534);
nor UO_1444 (O_1444,N_24762,N_24390);
xnor UO_1445 (O_1445,N_24720,N_24880);
xnor UO_1446 (O_1446,N_24945,N_24997);
or UO_1447 (O_1447,N_24427,N_24954);
or UO_1448 (O_1448,N_24766,N_24999);
and UO_1449 (O_1449,N_24411,N_24670);
xnor UO_1450 (O_1450,N_24636,N_24390);
and UO_1451 (O_1451,N_24507,N_24508);
nand UO_1452 (O_1452,N_24692,N_24845);
nor UO_1453 (O_1453,N_24597,N_24908);
nand UO_1454 (O_1454,N_24759,N_24509);
or UO_1455 (O_1455,N_24669,N_24753);
or UO_1456 (O_1456,N_24539,N_24793);
nor UO_1457 (O_1457,N_24865,N_24952);
nor UO_1458 (O_1458,N_24698,N_24428);
nand UO_1459 (O_1459,N_24848,N_24633);
nand UO_1460 (O_1460,N_24460,N_24537);
nor UO_1461 (O_1461,N_24630,N_24496);
nor UO_1462 (O_1462,N_24829,N_24523);
xor UO_1463 (O_1463,N_24494,N_24408);
or UO_1464 (O_1464,N_24628,N_24823);
xnor UO_1465 (O_1465,N_24731,N_24891);
or UO_1466 (O_1466,N_24800,N_24968);
nand UO_1467 (O_1467,N_24535,N_24807);
and UO_1468 (O_1468,N_24521,N_24533);
xnor UO_1469 (O_1469,N_24965,N_24998);
nor UO_1470 (O_1470,N_24511,N_24950);
nor UO_1471 (O_1471,N_24822,N_24992);
and UO_1472 (O_1472,N_24895,N_24794);
or UO_1473 (O_1473,N_24402,N_24836);
or UO_1474 (O_1474,N_24637,N_24671);
and UO_1475 (O_1475,N_24989,N_24945);
and UO_1476 (O_1476,N_24436,N_24583);
and UO_1477 (O_1477,N_24743,N_24650);
or UO_1478 (O_1478,N_24675,N_24894);
nand UO_1479 (O_1479,N_24925,N_24563);
nand UO_1480 (O_1480,N_24403,N_24749);
or UO_1481 (O_1481,N_24677,N_24399);
xor UO_1482 (O_1482,N_24851,N_24824);
nand UO_1483 (O_1483,N_24827,N_24712);
nor UO_1484 (O_1484,N_24827,N_24746);
xnor UO_1485 (O_1485,N_24809,N_24399);
xor UO_1486 (O_1486,N_24901,N_24496);
nand UO_1487 (O_1487,N_24792,N_24617);
nor UO_1488 (O_1488,N_24997,N_24516);
nor UO_1489 (O_1489,N_24448,N_24604);
xor UO_1490 (O_1490,N_24697,N_24595);
and UO_1491 (O_1491,N_24425,N_24517);
and UO_1492 (O_1492,N_24724,N_24777);
and UO_1493 (O_1493,N_24427,N_24911);
nand UO_1494 (O_1494,N_24456,N_24868);
xnor UO_1495 (O_1495,N_24964,N_24979);
xor UO_1496 (O_1496,N_24615,N_24668);
or UO_1497 (O_1497,N_24712,N_24576);
xnor UO_1498 (O_1498,N_24846,N_24757);
or UO_1499 (O_1499,N_24730,N_24667);
xnor UO_1500 (O_1500,N_24888,N_24779);
or UO_1501 (O_1501,N_24478,N_24572);
or UO_1502 (O_1502,N_24976,N_24788);
xor UO_1503 (O_1503,N_24917,N_24669);
xnor UO_1504 (O_1504,N_24461,N_24908);
and UO_1505 (O_1505,N_24780,N_24628);
or UO_1506 (O_1506,N_24428,N_24824);
or UO_1507 (O_1507,N_24713,N_24647);
nor UO_1508 (O_1508,N_24675,N_24902);
or UO_1509 (O_1509,N_24549,N_24592);
or UO_1510 (O_1510,N_24572,N_24846);
nor UO_1511 (O_1511,N_24741,N_24603);
nor UO_1512 (O_1512,N_24474,N_24753);
and UO_1513 (O_1513,N_24553,N_24880);
nor UO_1514 (O_1514,N_24693,N_24498);
nor UO_1515 (O_1515,N_24855,N_24709);
or UO_1516 (O_1516,N_24824,N_24461);
nor UO_1517 (O_1517,N_24654,N_24735);
xor UO_1518 (O_1518,N_24954,N_24787);
nand UO_1519 (O_1519,N_24509,N_24502);
nand UO_1520 (O_1520,N_24814,N_24377);
nand UO_1521 (O_1521,N_24972,N_24747);
nor UO_1522 (O_1522,N_24594,N_24850);
nor UO_1523 (O_1523,N_24681,N_24532);
or UO_1524 (O_1524,N_24609,N_24384);
or UO_1525 (O_1525,N_24973,N_24675);
nand UO_1526 (O_1526,N_24776,N_24773);
and UO_1527 (O_1527,N_24706,N_24565);
and UO_1528 (O_1528,N_24865,N_24825);
xnor UO_1529 (O_1529,N_24464,N_24995);
nor UO_1530 (O_1530,N_24588,N_24571);
nor UO_1531 (O_1531,N_24959,N_24843);
or UO_1532 (O_1532,N_24510,N_24950);
nand UO_1533 (O_1533,N_24748,N_24772);
nor UO_1534 (O_1534,N_24506,N_24573);
and UO_1535 (O_1535,N_24599,N_24645);
xnor UO_1536 (O_1536,N_24868,N_24984);
nor UO_1537 (O_1537,N_24868,N_24901);
and UO_1538 (O_1538,N_24717,N_24900);
xor UO_1539 (O_1539,N_24459,N_24597);
nand UO_1540 (O_1540,N_24845,N_24783);
or UO_1541 (O_1541,N_24874,N_24405);
and UO_1542 (O_1542,N_24665,N_24945);
xnor UO_1543 (O_1543,N_24861,N_24422);
xor UO_1544 (O_1544,N_24915,N_24665);
and UO_1545 (O_1545,N_24903,N_24988);
and UO_1546 (O_1546,N_24518,N_24879);
or UO_1547 (O_1547,N_24802,N_24598);
xnor UO_1548 (O_1548,N_24700,N_24457);
and UO_1549 (O_1549,N_24817,N_24548);
xor UO_1550 (O_1550,N_24876,N_24756);
or UO_1551 (O_1551,N_24562,N_24669);
nor UO_1552 (O_1552,N_24948,N_24904);
nand UO_1553 (O_1553,N_24418,N_24670);
nand UO_1554 (O_1554,N_24922,N_24780);
nor UO_1555 (O_1555,N_24399,N_24476);
xnor UO_1556 (O_1556,N_24591,N_24501);
nand UO_1557 (O_1557,N_24777,N_24867);
and UO_1558 (O_1558,N_24583,N_24798);
or UO_1559 (O_1559,N_24711,N_24407);
nand UO_1560 (O_1560,N_24804,N_24998);
xnor UO_1561 (O_1561,N_24876,N_24652);
and UO_1562 (O_1562,N_24658,N_24456);
nand UO_1563 (O_1563,N_24873,N_24633);
nor UO_1564 (O_1564,N_24593,N_24666);
or UO_1565 (O_1565,N_24933,N_24899);
and UO_1566 (O_1566,N_24603,N_24777);
xnor UO_1567 (O_1567,N_24380,N_24976);
nand UO_1568 (O_1568,N_24639,N_24974);
xor UO_1569 (O_1569,N_24399,N_24831);
and UO_1570 (O_1570,N_24885,N_24658);
nor UO_1571 (O_1571,N_24746,N_24612);
nand UO_1572 (O_1572,N_24877,N_24971);
or UO_1573 (O_1573,N_24388,N_24759);
nand UO_1574 (O_1574,N_24552,N_24956);
xnor UO_1575 (O_1575,N_24543,N_24568);
and UO_1576 (O_1576,N_24962,N_24857);
xnor UO_1577 (O_1577,N_24399,N_24675);
nand UO_1578 (O_1578,N_24428,N_24404);
xor UO_1579 (O_1579,N_24762,N_24610);
nor UO_1580 (O_1580,N_24674,N_24382);
xnor UO_1581 (O_1581,N_24883,N_24751);
nand UO_1582 (O_1582,N_24745,N_24642);
and UO_1583 (O_1583,N_24779,N_24568);
xor UO_1584 (O_1584,N_24678,N_24994);
or UO_1585 (O_1585,N_24476,N_24812);
nor UO_1586 (O_1586,N_24708,N_24540);
nand UO_1587 (O_1587,N_24496,N_24986);
and UO_1588 (O_1588,N_24673,N_24611);
or UO_1589 (O_1589,N_24759,N_24383);
and UO_1590 (O_1590,N_24414,N_24599);
nand UO_1591 (O_1591,N_24441,N_24429);
or UO_1592 (O_1592,N_24799,N_24883);
nor UO_1593 (O_1593,N_24740,N_24640);
nor UO_1594 (O_1594,N_24748,N_24918);
or UO_1595 (O_1595,N_24706,N_24947);
nor UO_1596 (O_1596,N_24387,N_24791);
nor UO_1597 (O_1597,N_24524,N_24912);
and UO_1598 (O_1598,N_24479,N_24835);
and UO_1599 (O_1599,N_24769,N_24814);
and UO_1600 (O_1600,N_24399,N_24626);
nand UO_1601 (O_1601,N_24388,N_24637);
and UO_1602 (O_1602,N_24827,N_24822);
or UO_1603 (O_1603,N_24643,N_24972);
and UO_1604 (O_1604,N_24929,N_24866);
xnor UO_1605 (O_1605,N_24732,N_24848);
nand UO_1606 (O_1606,N_24984,N_24601);
nand UO_1607 (O_1607,N_24415,N_24606);
xnor UO_1608 (O_1608,N_24584,N_24460);
xor UO_1609 (O_1609,N_24702,N_24698);
nor UO_1610 (O_1610,N_24467,N_24985);
nor UO_1611 (O_1611,N_24715,N_24848);
or UO_1612 (O_1612,N_24812,N_24907);
xor UO_1613 (O_1613,N_24937,N_24508);
and UO_1614 (O_1614,N_24486,N_24411);
nor UO_1615 (O_1615,N_24848,N_24494);
and UO_1616 (O_1616,N_24534,N_24636);
nand UO_1617 (O_1617,N_24561,N_24548);
or UO_1618 (O_1618,N_24769,N_24394);
xor UO_1619 (O_1619,N_24658,N_24453);
nand UO_1620 (O_1620,N_24807,N_24851);
nand UO_1621 (O_1621,N_24388,N_24898);
and UO_1622 (O_1622,N_24886,N_24988);
nand UO_1623 (O_1623,N_24873,N_24459);
xor UO_1624 (O_1624,N_24979,N_24704);
xor UO_1625 (O_1625,N_24667,N_24635);
or UO_1626 (O_1626,N_24709,N_24733);
xor UO_1627 (O_1627,N_24516,N_24653);
nand UO_1628 (O_1628,N_24764,N_24811);
and UO_1629 (O_1629,N_24661,N_24945);
or UO_1630 (O_1630,N_24462,N_24584);
and UO_1631 (O_1631,N_24573,N_24680);
nor UO_1632 (O_1632,N_24978,N_24525);
nor UO_1633 (O_1633,N_24836,N_24459);
or UO_1634 (O_1634,N_24865,N_24608);
xor UO_1635 (O_1635,N_24547,N_24469);
nor UO_1636 (O_1636,N_24655,N_24394);
or UO_1637 (O_1637,N_24387,N_24806);
or UO_1638 (O_1638,N_24620,N_24663);
nand UO_1639 (O_1639,N_24710,N_24816);
xor UO_1640 (O_1640,N_24786,N_24474);
and UO_1641 (O_1641,N_24625,N_24600);
nand UO_1642 (O_1642,N_24998,N_24812);
nor UO_1643 (O_1643,N_24850,N_24480);
nor UO_1644 (O_1644,N_24614,N_24747);
nand UO_1645 (O_1645,N_24550,N_24716);
or UO_1646 (O_1646,N_24393,N_24420);
xnor UO_1647 (O_1647,N_24858,N_24982);
xnor UO_1648 (O_1648,N_24814,N_24715);
nor UO_1649 (O_1649,N_24375,N_24804);
nor UO_1650 (O_1650,N_24704,N_24552);
nor UO_1651 (O_1651,N_24379,N_24774);
nor UO_1652 (O_1652,N_24630,N_24607);
nor UO_1653 (O_1653,N_24618,N_24990);
xnor UO_1654 (O_1654,N_24842,N_24980);
nor UO_1655 (O_1655,N_24554,N_24863);
and UO_1656 (O_1656,N_24856,N_24617);
or UO_1657 (O_1657,N_24637,N_24872);
or UO_1658 (O_1658,N_24610,N_24983);
xor UO_1659 (O_1659,N_24860,N_24651);
and UO_1660 (O_1660,N_24715,N_24569);
xor UO_1661 (O_1661,N_24393,N_24824);
nor UO_1662 (O_1662,N_24401,N_24852);
and UO_1663 (O_1663,N_24598,N_24911);
and UO_1664 (O_1664,N_24513,N_24863);
nand UO_1665 (O_1665,N_24764,N_24639);
nand UO_1666 (O_1666,N_24458,N_24688);
nand UO_1667 (O_1667,N_24995,N_24534);
nor UO_1668 (O_1668,N_24423,N_24481);
or UO_1669 (O_1669,N_24704,N_24611);
xor UO_1670 (O_1670,N_24552,N_24442);
nand UO_1671 (O_1671,N_24645,N_24974);
nor UO_1672 (O_1672,N_24405,N_24665);
xor UO_1673 (O_1673,N_24537,N_24602);
nand UO_1674 (O_1674,N_24866,N_24450);
nor UO_1675 (O_1675,N_24874,N_24871);
xnor UO_1676 (O_1676,N_24969,N_24930);
and UO_1677 (O_1677,N_24839,N_24566);
nand UO_1678 (O_1678,N_24416,N_24770);
nand UO_1679 (O_1679,N_24891,N_24400);
nor UO_1680 (O_1680,N_24720,N_24701);
or UO_1681 (O_1681,N_24912,N_24443);
nand UO_1682 (O_1682,N_24606,N_24470);
and UO_1683 (O_1683,N_24768,N_24973);
xor UO_1684 (O_1684,N_24517,N_24512);
nand UO_1685 (O_1685,N_24449,N_24751);
or UO_1686 (O_1686,N_24981,N_24460);
xor UO_1687 (O_1687,N_24976,N_24783);
and UO_1688 (O_1688,N_24494,N_24862);
and UO_1689 (O_1689,N_24630,N_24793);
xnor UO_1690 (O_1690,N_24951,N_24636);
nor UO_1691 (O_1691,N_24409,N_24836);
and UO_1692 (O_1692,N_24992,N_24634);
xnor UO_1693 (O_1693,N_24581,N_24897);
nand UO_1694 (O_1694,N_24416,N_24936);
nor UO_1695 (O_1695,N_24444,N_24951);
nor UO_1696 (O_1696,N_24645,N_24899);
nand UO_1697 (O_1697,N_24798,N_24571);
xnor UO_1698 (O_1698,N_24886,N_24533);
nand UO_1699 (O_1699,N_24642,N_24619);
nor UO_1700 (O_1700,N_24642,N_24418);
and UO_1701 (O_1701,N_24928,N_24397);
nand UO_1702 (O_1702,N_24407,N_24569);
or UO_1703 (O_1703,N_24548,N_24823);
nand UO_1704 (O_1704,N_24651,N_24596);
xnor UO_1705 (O_1705,N_24839,N_24773);
and UO_1706 (O_1706,N_24695,N_24618);
or UO_1707 (O_1707,N_24850,N_24499);
nand UO_1708 (O_1708,N_24417,N_24797);
xor UO_1709 (O_1709,N_24875,N_24555);
xnor UO_1710 (O_1710,N_24989,N_24860);
and UO_1711 (O_1711,N_24410,N_24421);
xor UO_1712 (O_1712,N_24773,N_24451);
nand UO_1713 (O_1713,N_24619,N_24707);
and UO_1714 (O_1714,N_24779,N_24885);
and UO_1715 (O_1715,N_24468,N_24426);
nand UO_1716 (O_1716,N_24813,N_24667);
nor UO_1717 (O_1717,N_24667,N_24520);
or UO_1718 (O_1718,N_24938,N_24831);
and UO_1719 (O_1719,N_24536,N_24615);
xor UO_1720 (O_1720,N_24880,N_24565);
or UO_1721 (O_1721,N_24666,N_24441);
or UO_1722 (O_1722,N_24811,N_24591);
nor UO_1723 (O_1723,N_24646,N_24517);
or UO_1724 (O_1724,N_24561,N_24544);
nand UO_1725 (O_1725,N_24794,N_24495);
xor UO_1726 (O_1726,N_24679,N_24420);
or UO_1727 (O_1727,N_24449,N_24490);
xor UO_1728 (O_1728,N_24536,N_24795);
or UO_1729 (O_1729,N_24398,N_24946);
xor UO_1730 (O_1730,N_24920,N_24764);
xnor UO_1731 (O_1731,N_24871,N_24779);
or UO_1732 (O_1732,N_24850,N_24636);
xnor UO_1733 (O_1733,N_24795,N_24631);
nand UO_1734 (O_1734,N_24622,N_24480);
nand UO_1735 (O_1735,N_24585,N_24718);
xor UO_1736 (O_1736,N_24755,N_24847);
nand UO_1737 (O_1737,N_24510,N_24733);
and UO_1738 (O_1738,N_24618,N_24656);
and UO_1739 (O_1739,N_24438,N_24907);
nand UO_1740 (O_1740,N_24386,N_24525);
nor UO_1741 (O_1741,N_24554,N_24672);
nor UO_1742 (O_1742,N_24706,N_24702);
nand UO_1743 (O_1743,N_24619,N_24946);
nand UO_1744 (O_1744,N_24543,N_24718);
and UO_1745 (O_1745,N_24846,N_24966);
nand UO_1746 (O_1746,N_24725,N_24997);
xor UO_1747 (O_1747,N_24942,N_24915);
nor UO_1748 (O_1748,N_24465,N_24740);
or UO_1749 (O_1749,N_24545,N_24978);
and UO_1750 (O_1750,N_24508,N_24645);
nor UO_1751 (O_1751,N_24996,N_24473);
xnor UO_1752 (O_1752,N_24788,N_24687);
nand UO_1753 (O_1753,N_24878,N_24875);
xnor UO_1754 (O_1754,N_24811,N_24938);
and UO_1755 (O_1755,N_24829,N_24660);
and UO_1756 (O_1756,N_24884,N_24942);
and UO_1757 (O_1757,N_24462,N_24958);
nand UO_1758 (O_1758,N_24835,N_24776);
nor UO_1759 (O_1759,N_24833,N_24825);
nand UO_1760 (O_1760,N_24691,N_24853);
and UO_1761 (O_1761,N_24900,N_24391);
and UO_1762 (O_1762,N_24980,N_24611);
nand UO_1763 (O_1763,N_24902,N_24698);
nand UO_1764 (O_1764,N_24635,N_24490);
and UO_1765 (O_1765,N_24446,N_24881);
nor UO_1766 (O_1766,N_24902,N_24621);
or UO_1767 (O_1767,N_24982,N_24671);
and UO_1768 (O_1768,N_24599,N_24381);
nand UO_1769 (O_1769,N_24538,N_24385);
and UO_1770 (O_1770,N_24458,N_24661);
xor UO_1771 (O_1771,N_24428,N_24691);
or UO_1772 (O_1772,N_24883,N_24487);
and UO_1773 (O_1773,N_24534,N_24747);
and UO_1774 (O_1774,N_24615,N_24616);
and UO_1775 (O_1775,N_24799,N_24738);
nand UO_1776 (O_1776,N_24959,N_24602);
or UO_1777 (O_1777,N_24387,N_24554);
and UO_1778 (O_1778,N_24564,N_24483);
or UO_1779 (O_1779,N_24465,N_24801);
nand UO_1780 (O_1780,N_24629,N_24946);
nand UO_1781 (O_1781,N_24525,N_24456);
nand UO_1782 (O_1782,N_24495,N_24968);
xnor UO_1783 (O_1783,N_24842,N_24944);
nor UO_1784 (O_1784,N_24745,N_24586);
or UO_1785 (O_1785,N_24894,N_24401);
or UO_1786 (O_1786,N_24939,N_24906);
nor UO_1787 (O_1787,N_24494,N_24780);
xor UO_1788 (O_1788,N_24615,N_24612);
nand UO_1789 (O_1789,N_24731,N_24527);
xnor UO_1790 (O_1790,N_24857,N_24683);
nor UO_1791 (O_1791,N_24467,N_24776);
or UO_1792 (O_1792,N_24738,N_24721);
or UO_1793 (O_1793,N_24656,N_24590);
nand UO_1794 (O_1794,N_24731,N_24953);
and UO_1795 (O_1795,N_24682,N_24541);
nand UO_1796 (O_1796,N_24424,N_24438);
nor UO_1797 (O_1797,N_24400,N_24878);
and UO_1798 (O_1798,N_24394,N_24382);
and UO_1799 (O_1799,N_24403,N_24675);
or UO_1800 (O_1800,N_24983,N_24467);
or UO_1801 (O_1801,N_24574,N_24612);
or UO_1802 (O_1802,N_24523,N_24606);
nand UO_1803 (O_1803,N_24703,N_24597);
and UO_1804 (O_1804,N_24456,N_24534);
or UO_1805 (O_1805,N_24967,N_24960);
or UO_1806 (O_1806,N_24564,N_24796);
or UO_1807 (O_1807,N_24768,N_24426);
nand UO_1808 (O_1808,N_24582,N_24511);
nor UO_1809 (O_1809,N_24542,N_24787);
nand UO_1810 (O_1810,N_24401,N_24794);
xnor UO_1811 (O_1811,N_24791,N_24663);
nand UO_1812 (O_1812,N_24599,N_24697);
or UO_1813 (O_1813,N_24533,N_24900);
and UO_1814 (O_1814,N_24622,N_24618);
nand UO_1815 (O_1815,N_24877,N_24713);
and UO_1816 (O_1816,N_24964,N_24896);
and UO_1817 (O_1817,N_24767,N_24962);
nor UO_1818 (O_1818,N_24710,N_24432);
nand UO_1819 (O_1819,N_24686,N_24687);
nor UO_1820 (O_1820,N_24646,N_24758);
or UO_1821 (O_1821,N_24787,N_24974);
xor UO_1822 (O_1822,N_24833,N_24566);
nor UO_1823 (O_1823,N_24748,N_24379);
nor UO_1824 (O_1824,N_24969,N_24853);
nor UO_1825 (O_1825,N_24534,N_24547);
xnor UO_1826 (O_1826,N_24774,N_24878);
nor UO_1827 (O_1827,N_24988,N_24504);
xor UO_1828 (O_1828,N_24422,N_24857);
nor UO_1829 (O_1829,N_24823,N_24974);
or UO_1830 (O_1830,N_24966,N_24536);
nor UO_1831 (O_1831,N_24585,N_24658);
or UO_1832 (O_1832,N_24924,N_24394);
nor UO_1833 (O_1833,N_24903,N_24627);
nor UO_1834 (O_1834,N_24847,N_24585);
nor UO_1835 (O_1835,N_24703,N_24536);
nand UO_1836 (O_1836,N_24999,N_24433);
nor UO_1837 (O_1837,N_24761,N_24435);
nand UO_1838 (O_1838,N_24830,N_24907);
nor UO_1839 (O_1839,N_24691,N_24833);
xnor UO_1840 (O_1840,N_24612,N_24984);
nor UO_1841 (O_1841,N_24954,N_24579);
xor UO_1842 (O_1842,N_24866,N_24521);
nand UO_1843 (O_1843,N_24910,N_24740);
and UO_1844 (O_1844,N_24507,N_24635);
and UO_1845 (O_1845,N_24533,N_24570);
or UO_1846 (O_1846,N_24499,N_24533);
and UO_1847 (O_1847,N_24915,N_24379);
nor UO_1848 (O_1848,N_24703,N_24710);
xnor UO_1849 (O_1849,N_24872,N_24790);
nand UO_1850 (O_1850,N_24623,N_24746);
and UO_1851 (O_1851,N_24963,N_24424);
or UO_1852 (O_1852,N_24884,N_24843);
nand UO_1853 (O_1853,N_24593,N_24978);
nand UO_1854 (O_1854,N_24592,N_24595);
xor UO_1855 (O_1855,N_24454,N_24780);
and UO_1856 (O_1856,N_24511,N_24656);
and UO_1857 (O_1857,N_24547,N_24504);
xor UO_1858 (O_1858,N_24444,N_24656);
or UO_1859 (O_1859,N_24525,N_24481);
and UO_1860 (O_1860,N_24758,N_24820);
xor UO_1861 (O_1861,N_24501,N_24571);
xor UO_1862 (O_1862,N_24756,N_24714);
nor UO_1863 (O_1863,N_24516,N_24913);
nand UO_1864 (O_1864,N_24944,N_24408);
and UO_1865 (O_1865,N_24746,N_24771);
or UO_1866 (O_1866,N_24792,N_24893);
and UO_1867 (O_1867,N_24730,N_24407);
and UO_1868 (O_1868,N_24963,N_24419);
xnor UO_1869 (O_1869,N_24834,N_24883);
xor UO_1870 (O_1870,N_24743,N_24958);
or UO_1871 (O_1871,N_24779,N_24980);
nand UO_1872 (O_1872,N_24843,N_24853);
and UO_1873 (O_1873,N_24628,N_24971);
or UO_1874 (O_1874,N_24601,N_24489);
and UO_1875 (O_1875,N_24779,N_24804);
xor UO_1876 (O_1876,N_24621,N_24392);
or UO_1877 (O_1877,N_24518,N_24685);
and UO_1878 (O_1878,N_24580,N_24626);
nor UO_1879 (O_1879,N_24925,N_24408);
nor UO_1880 (O_1880,N_24894,N_24561);
and UO_1881 (O_1881,N_24892,N_24514);
or UO_1882 (O_1882,N_24435,N_24476);
nor UO_1883 (O_1883,N_24579,N_24708);
xor UO_1884 (O_1884,N_24887,N_24428);
and UO_1885 (O_1885,N_24938,N_24964);
nor UO_1886 (O_1886,N_24585,N_24529);
or UO_1887 (O_1887,N_24606,N_24424);
or UO_1888 (O_1888,N_24867,N_24653);
nand UO_1889 (O_1889,N_24414,N_24868);
nand UO_1890 (O_1890,N_24625,N_24382);
and UO_1891 (O_1891,N_24701,N_24479);
or UO_1892 (O_1892,N_24724,N_24504);
and UO_1893 (O_1893,N_24940,N_24967);
xnor UO_1894 (O_1894,N_24932,N_24418);
or UO_1895 (O_1895,N_24414,N_24493);
xor UO_1896 (O_1896,N_24438,N_24390);
xnor UO_1897 (O_1897,N_24759,N_24998);
nor UO_1898 (O_1898,N_24621,N_24769);
nor UO_1899 (O_1899,N_24607,N_24965);
and UO_1900 (O_1900,N_24683,N_24773);
nand UO_1901 (O_1901,N_24703,N_24787);
or UO_1902 (O_1902,N_24546,N_24811);
and UO_1903 (O_1903,N_24572,N_24927);
nand UO_1904 (O_1904,N_24796,N_24610);
xor UO_1905 (O_1905,N_24639,N_24530);
nor UO_1906 (O_1906,N_24379,N_24664);
nand UO_1907 (O_1907,N_24758,N_24653);
xnor UO_1908 (O_1908,N_24854,N_24896);
or UO_1909 (O_1909,N_24950,N_24668);
nand UO_1910 (O_1910,N_24868,N_24439);
nand UO_1911 (O_1911,N_24837,N_24520);
nand UO_1912 (O_1912,N_24751,N_24874);
nand UO_1913 (O_1913,N_24862,N_24950);
nand UO_1914 (O_1914,N_24500,N_24507);
nand UO_1915 (O_1915,N_24755,N_24720);
or UO_1916 (O_1916,N_24695,N_24460);
nor UO_1917 (O_1917,N_24485,N_24701);
nand UO_1918 (O_1918,N_24833,N_24690);
nand UO_1919 (O_1919,N_24489,N_24914);
xor UO_1920 (O_1920,N_24396,N_24705);
or UO_1921 (O_1921,N_24955,N_24834);
or UO_1922 (O_1922,N_24905,N_24644);
nor UO_1923 (O_1923,N_24468,N_24615);
or UO_1924 (O_1924,N_24604,N_24729);
or UO_1925 (O_1925,N_24521,N_24737);
nor UO_1926 (O_1926,N_24431,N_24990);
nor UO_1927 (O_1927,N_24477,N_24765);
xnor UO_1928 (O_1928,N_24874,N_24846);
and UO_1929 (O_1929,N_24430,N_24610);
nor UO_1930 (O_1930,N_24649,N_24456);
or UO_1931 (O_1931,N_24831,N_24467);
xnor UO_1932 (O_1932,N_24821,N_24440);
or UO_1933 (O_1933,N_24617,N_24601);
or UO_1934 (O_1934,N_24806,N_24609);
or UO_1935 (O_1935,N_24424,N_24867);
or UO_1936 (O_1936,N_24699,N_24852);
or UO_1937 (O_1937,N_24736,N_24826);
xor UO_1938 (O_1938,N_24973,N_24773);
nand UO_1939 (O_1939,N_24766,N_24989);
or UO_1940 (O_1940,N_24951,N_24666);
and UO_1941 (O_1941,N_24729,N_24631);
xnor UO_1942 (O_1942,N_24566,N_24485);
xor UO_1943 (O_1943,N_24636,N_24432);
nand UO_1944 (O_1944,N_24620,N_24762);
or UO_1945 (O_1945,N_24901,N_24684);
nor UO_1946 (O_1946,N_24766,N_24567);
and UO_1947 (O_1947,N_24646,N_24766);
or UO_1948 (O_1948,N_24402,N_24791);
xnor UO_1949 (O_1949,N_24883,N_24441);
or UO_1950 (O_1950,N_24800,N_24878);
nand UO_1951 (O_1951,N_24909,N_24882);
nor UO_1952 (O_1952,N_24597,N_24639);
nor UO_1953 (O_1953,N_24938,N_24698);
and UO_1954 (O_1954,N_24746,N_24848);
nand UO_1955 (O_1955,N_24905,N_24814);
nand UO_1956 (O_1956,N_24595,N_24533);
nor UO_1957 (O_1957,N_24623,N_24945);
xor UO_1958 (O_1958,N_24872,N_24689);
and UO_1959 (O_1959,N_24809,N_24414);
nor UO_1960 (O_1960,N_24421,N_24649);
nor UO_1961 (O_1961,N_24845,N_24724);
or UO_1962 (O_1962,N_24392,N_24553);
or UO_1963 (O_1963,N_24819,N_24741);
or UO_1964 (O_1964,N_24595,N_24419);
nor UO_1965 (O_1965,N_24800,N_24393);
xor UO_1966 (O_1966,N_24681,N_24754);
nand UO_1967 (O_1967,N_24432,N_24402);
nand UO_1968 (O_1968,N_24793,N_24832);
nor UO_1969 (O_1969,N_24978,N_24764);
or UO_1970 (O_1970,N_24544,N_24465);
xor UO_1971 (O_1971,N_24613,N_24935);
nand UO_1972 (O_1972,N_24399,N_24765);
or UO_1973 (O_1973,N_24689,N_24627);
nor UO_1974 (O_1974,N_24992,N_24623);
nand UO_1975 (O_1975,N_24982,N_24686);
xor UO_1976 (O_1976,N_24693,N_24547);
nand UO_1977 (O_1977,N_24744,N_24674);
nor UO_1978 (O_1978,N_24650,N_24535);
nor UO_1979 (O_1979,N_24834,N_24909);
and UO_1980 (O_1980,N_24713,N_24403);
and UO_1981 (O_1981,N_24607,N_24435);
xor UO_1982 (O_1982,N_24989,N_24551);
xor UO_1983 (O_1983,N_24783,N_24850);
or UO_1984 (O_1984,N_24648,N_24942);
nand UO_1985 (O_1985,N_24402,N_24820);
nand UO_1986 (O_1986,N_24989,N_24500);
xor UO_1987 (O_1987,N_24759,N_24738);
xor UO_1988 (O_1988,N_24543,N_24842);
xnor UO_1989 (O_1989,N_24439,N_24757);
and UO_1990 (O_1990,N_24686,N_24477);
xnor UO_1991 (O_1991,N_24402,N_24668);
nor UO_1992 (O_1992,N_24894,N_24867);
nor UO_1993 (O_1993,N_24696,N_24874);
xor UO_1994 (O_1994,N_24853,N_24517);
and UO_1995 (O_1995,N_24769,N_24381);
xnor UO_1996 (O_1996,N_24881,N_24482);
nand UO_1997 (O_1997,N_24406,N_24554);
or UO_1998 (O_1998,N_24549,N_24466);
nor UO_1999 (O_1999,N_24422,N_24432);
and UO_2000 (O_2000,N_24493,N_24580);
or UO_2001 (O_2001,N_24569,N_24789);
or UO_2002 (O_2002,N_24833,N_24523);
nor UO_2003 (O_2003,N_24947,N_24722);
or UO_2004 (O_2004,N_24698,N_24579);
xor UO_2005 (O_2005,N_24917,N_24939);
nor UO_2006 (O_2006,N_24758,N_24761);
and UO_2007 (O_2007,N_24635,N_24567);
nor UO_2008 (O_2008,N_24583,N_24714);
nand UO_2009 (O_2009,N_24777,N_24774);
or UO_2010 (O_2010,N_24479,N_24870);
or UO_2011 (O_2011,N_24945,N_24906);
nor UO_2012 (O_2012,N_24760,N_24508);
and UO_2013 (O_2013,N_24844,N_24483);
nor UO_2014 (O_2014,N_24844,N_24900);
or UO_2015 (O_2015,N_24889,N_24684);
nor UO_2016 (O_2016,N_24467,N_24959);
or UO_2017 (O_2017,N_24492,N_24406);
or UO_2018 (O_2018,N_24794,N_24922);
or UO_2019 (O_2019,N_24515,N_24982);
or UO_2020 (O_2020,N_24527,N_24428);
or UO_2021 (O_2021,N_24516,N_24959);
or UO_2022 (O_2022,N_24390,N_24998);
nor UO_2023 (O_2023,N_24934,N_24382);
nand UO_2024 (O_2024,N_24667,N_24634);
nor UO_2025 (O_2025,N_24507,N_24881);
nor UO_2026 (O_2026,N_24588,N_24851);
xor UO_2027 (O_2027,N_24469,N_24868);
or UO_2028 (O_2028,N_24611,N_24613);
nand UO_2029 (O_2029,N_24821,N_24909);
or UO_2030 (O_2030,N_24972,N_24780);
or UO_2031 (O_2031,N_24658,N_24421);
xnor UO_2032 (O_2032,N_24476,N_24712);
and UO_2033 (O_2033,N_24603,N_24836);
and UO_2034 (O_2034,N_24676,N_24985);
nand UO_2035 (O_2035,N_24586,N_24507);
nand UO_2036 (O_2036,N_24685,N_24951);
nand UO_2037 (O_2037,N_24645,N_24997);
and UO_2038 (O_2038,N_24802,N_24610);
nand UO_2039 (O_2039,N_24660,N_24403);
or UO_2040 (O_2040,N_24562,N_24426);
nand UO_2041 (O_2041,N_24991,N_24551);
nor UO_2042 (O_2042,N_24531,N_24811);
xnor UO_2043 (O_2043,N_24809,N_24678);
nor UO_2044 (O_2044,N_24987,N_24852);
xor UO_2045 (O_2045,N_24631,N_24574);
and UO_2046 (O_2046,N_24511,N_24571);
and UO_2047 (O_2047,N_24438,N_24881);
nand UO_2048 (O_2048,N_24953,N_24402);
xnor UO_2049 (O_2049,N_24895,N_24857);
or UO_2050 (O_2050,N_24674,N_24644);
nand UO_2051 (O_2051,N_24767,N_24490);
or UO_2052 (O_2052,N_24943,N_24519);
and UO_2053 (O_2053,N_24858,N_24697);
nand UO_2054 (O_2054,N_24434,N_24492);
nor UO_2055 (O_2055,N_24642,N_24524);
and UO_2056 (O_2056,N_24416,N_24810);
xnor UO_2057 (O_2057,N_24600,N_24458);
nor UO_2058 (O_2058,N_24581,N_24456);
xnor UO_2059 (O_2059,N_24409,N_24551);
or UO_2060 (O_2060,N_24774,N_24738);
xnor UO_2061 (O_2061,N_24649,N_24996);
and UO_2062 (O_2062,N_24681,N_24858);
and UO_2063 (O_2063,N_24904,N_24916);
xnor UO_2064 (O_2064,N_24420,N_24515);
nand UO_2065 (O_2065,N_24749,N_24759);
xor UO_2066 (O_2066,N_24566,N_24723);
nor UO_2067 (O_2067,N_24403,N_24659);
nand UO_2068 (O_2068,N_24945,N_24587);
xor UO_2069 (O_2069,N_24431,N_24907);
nor UO_2070 (O_2070,N_24824,N_24708);
or UO_2071 (O_2071,N_24410,N_24937);
xor UO_2072 (O_2072,N_24379,N_24626);
nand UO_2073 (O_2073,N_24924,N_24654);
nand UO_2074 (O_2074,N_24983,N_24702);
nor UO_2075 (O_2075,N_24689,N_24615);
nor UO_2076 (O_2076,N_24963,N_24612);
nor UO_2077 (O_2077,N_24920,N_24966);
or UO_2078 (O_2078,N_24423,N_24432);
nor UO_2079 (O_2079,N_24673,N_24561);
nand UO_2080 (O_2080,N_24482,N_24558);
nand UO_2081 (O_2081,N_24644,N_24907);
nor UO_2082 (O_2082,N_24614,N_24375);
and UO_2083 (O_2083,N_24388,N_24415);
and UO_2084 (O_2084,N_24739,N_24468);
nor UO_2085 (O_2085,N_24520,N_24880);
nor UO_2086 (O_2086,N_24536,N_24759);
or UO_2087 (O_2087,N_24859,N_24907);
xor UO_2088 (O_2088,N_24915,N_24671);
and UO_2089 (O_2089,N_24676,N_24675);
and UO_2090 (O_2090,N_24566,N_24747);
xor UO_2091 (O_2091,N_24766,N_24820);
nor UO_2092 (O_2092,N_24839,N_24757);
nand UO_2093 (O_2093,N_24620,N_24635);
or UO_2094 (O_2094,N_24666,N_24795);
nor UO_2095 (O_2095,N_24649,N_24755);
nor UO_2096 (O_2096,N_24994,N_24974);
and UO_2097 (O_2097,N_24997,N_24526);
xnor UO_2098 (O_2098,N_24530,N_24798);
or UO_2099 (O_2099,N_24452,N_24446);
and UO_2100 (O_2100,N_24431,N_24562);
or UO_2101 (O_2101,N_24460,N_24396);
or UO_2102 (O_2102,N_24787,N_24495);
and UO_2103 (O_2103,N_24860,N_24634);
and UO_2104 (O_2104,N_24789,N_24723);
nand UO_2105 (O_2105,N_24515,N_24523);
nand UO_2106 (O_2106,N_24963,N_24592);
and UO_2107 (O_2107,N_24928,N_24782);
nor UO_2108 (O_2108,N_24850,N_24675);
and UO_2109 (O_2109,N_24682,N_24428);
nor UO_2110 (O_2110,N_24743,N_24941);
and UO_2111 (O_2111,N_24654,N_24591);
xnor UO_2112 (O_2112,N_24810,N_24713);
nand UO_2113 (O_2113,N_24652,N_24670);
nor UO_2114 (O_2114,N_24669,N_24767);
nor UO_2115 (O_2115,N_24688,N_24499);
or UO_2116 (O_2116,N_24599,N_24776);
nor UO_2117 (O_2117,N_24826,N_24404);
xor UO_2118 (O_2118,N_24379,N_24860);
nand UO_2119 (O_2119,N_24388,N_24901);
nand UO_2120 (O_2120,N_24697,N_24774);
xor UO_2121 (O_2121,N_24662,N_24867);
and UO_2122 (O_2122,N_24582,N_24743);
or UO_2123 (O_2123,N_24740,N_24834);
or UO_2124 (O_2124,N_24879,N_24795);
and UO_2125 (O_2125,N_24706,N_24644);
nand UO_2126 (O_2126,N_24492,N_24696);
nand UO_2127 (O_2127,N_24608,N_24883);
xnor UO_2128 (O_2128,N_24678,N_24970);
or UO_2129 (O_2129,N_24836,N_24602);
nand UO_2130 (O_2130,N_24957,N_24538);
and UO_2131 (O_2131,N_24938,N_24808);
nand UO_2132 (O_2132,N_24862,N_24932);
and UO_2133 (O_2133,N_24930,N_24922);
nor UO_2134 (O_2134,N_24432,N_24689);
nor UO_2135 (O_2135,N_24765,N_24476);
nand UO_2136 (O_2136,N_24706,N_24787);
or UO_2137 (O_2137,N_24984,N_24704);
or UO_2138 (O_2138,N_24413,N_24859);
xor UO_2139 (O_2139,N_24993,N_24636);
nor UO_2140 (O_2140,N_24916,N_24720);
nand UO_2141 (O_2141,N_24860,N_24446);
nor UO_2142 (O_2142,N_24715,N_24404);
xor UO_2143 (O_2143,N_24947,N_24905);
nor UO_2144 (O_2144,N_24386,N_24873);
nor UO_2145 (O_2145,N_24731,N_24410);
or UO_2146 (O_2146,N_24624,N_24614);
nor UO_2147 (O_2147,N_24642,N_24507);
nand UO_2148 (O_2148,N_24840,N_24668);
or UO_2149 (O_2149,N_24767,N_24453);
nor UO_2150 (O_2150,N_24516,N_24513);
and UO_2151 (O_2151,N_24475,N_24384);
nor UO_2152 (O_2152,N_24693,N_24679);
xnor UO_2153 (O_2153,N_24565,N_24666);
xor UO_2154 (O_2154,N_24975,N_24420);
or UO_2155 (O_2155,N_24660,N_24543);
and UO_2156 (O_2156,N_24461,N_24987);
or UO_2157 (O_2157,N_24647,N_24862);
nand UO_2158 (O_2158,N_24843,N_24715);
or UO_2159 (O_2159,N_24643,N_24572);
xor UO_2160 (O_2160,N_24516,N_24859);
nor UO_2161 (O_2161,N_24557,N_24529);
or UO_2162 (O_2162,N_24742,N_24611);
nor UO_2163 (O_2163,N_24473,N_24613);
xnor UO_2164 (O_2164,N_24466,N_24607);
or UO_2165 (O_2165,N_24851,N_24414);
and UO_2166 (O_2166,N_24808,N_24906);
nor UO_2167 (O_2167,N_24879,N_24872);
and UO_2168 (O_2168,N_24685,N_24964);
and UO_2169 (O_2169,N_24546,N_24876);
and UO_2170 (O_2170,N_24453,N_24946);
nor UO_2171 (O_2171,N_24930,N_24403);
nor UO_2172 (O_2172,N_24499,N_24653);
and UO_2173 (O_2173,N_24936,N_24894);
xnor UO_2174 (O_2174,N_24406,N_24919);
nand UO_2175 (O_2175,N_24780,N_24745);
or UO_2176 (O_2176,N_24480,N_24943);
or UO_2177 (O_2177,N_24682,N_24445);
nor UO_2178 (O_2178,N_24556,N_24861);
xnor UO_2179 (O_2179,N_24692,N_24514);
nor UO_2180 (O_2180,N_24878,N_24684);
nor UO_2181 (O_2181,N_24461,N_24411);
or UO_2182 (O_2182,N_24637,N_24432);
and UO_2183 (O_2183,N_24897,N_24697);
xor UO_2184 (O_2184,N_24663,N_24516);
nor UO_2185 (O_2185,N_24564,N_24944);
nand UO_2186 (O_2186,N_24894,N_24613);
and UO_2187 (O_2187,N_24762,N_24619);
and UO_2188 (O_2188,N_24647,N_24908);
xor UO_2189 (O_2189,N_24741,N_24733);
xor UO_2190 (O_2190,N_24923,N_24548);
or UO_2191 (O_2191,N_24724,N_24607);
xnor UO_2192 (O_2192,N_24555,N_24567);
nor UO_2193 (O_2193,N_24897,N_24979);
or UO_2194 (O_2194,N_24461,N_24811);
nor UO_2195 (O_2195,N_24805,N_24755);
xor UO_2196 (O_2196,N_24547,N_24572);
and UO_2197 (O_2197,N_24601,N_24862);
nand UO_2198 (O_2198,N_24862,N_24836);
nor UO_2199 (O_2199,N_24659,N_24409);
nor UO_2200 (O_2200,N_24845,N_24422);
and UO_2201 (O_2201,N_24676,N_24997);
xor UO_2202 (O_2202,N_24457,N_24742);
nor UO_2203 (O_2203,N_24522,N_24810);
and UO_2204 (O_2204,N_24601,N_24434);
and UO_2205 (O_2205,N_24568,N_24634);
nand UO_2206 (O_2206,N_24714,N_24941);
nor UO_2207 (O_2207,N_24889,N_24703);
and UO_2208 (O_2208,N_24658,N_24740);
and UO_2209 (O_2209,N_24569,N_24500);
xor UO_2210 (O_2210,N_24837,N_24598);
nor UO_2211 (O_2211,N_24862,N_24552);
nor UO_2212 (O_2212,N_24816,N_24963);
and UO_2213 (O_2213,N_24750,N_24632);
nor UO_2214 (O_2214,N_24494,N_24980);
nand UO_2215 (O_2215,N_24646,N_24520);
nand UO_2216 (O_2216,N_24592,N_24807);
nand UO_2217 (O_2217,N_24468,N_24392);
xor UO_2218 (O_2218,N_24616,N_24641);
xor UO_2219 (O_2219,N_24773,N_24964);
and UO_2220 (O_2220,N_24685,N_24843);
and UO_2221 (O_2221,N_24497,N_24629);
xor UO_2222 (O_2222,N_24690,N_24528);
xor UO_2223 (O_2223,N_24850,N_24393);
nor UO_2224 (O_2224,N_24984,N_24710);
nor UO_2225 (O_2225,N_24883,N_24940);
and UO_2226 (O_2226,N_24950,N_24563);
nor UO_2227 (O_2227,N_24416,N_24754);
or UO_2228 (O_2228,N_24658,N_24702);
nor UO_2229 (O_2229,N_24525,N_24501);
nor UO_2230 (O_2230,N_24877,N_24418);
xnor UO_2231 (O_2231,N_24405,N_24849);
nor UO_2232 (O_2232,N_24398,N_24964);
and UO_2233 (O_2233,N_24762,N_24990);
or UO_2234 (O_2234,N_24765,N_24899);
xor UO_2235 (O_2235,N_24415,N_24598);
nand UO_2236 (O_2236,N_24426,N_24404);
nor UO_2237 (O_2237,N_24581,N_24919);
and UO_2238 (O_2238,N_24826,N_24997);
and UO_2239 (O_2239,N_24427,N_24619);
xor UO_2240 (O_2240,N_24432,N_24508);
nand UO_2241 (O_2241,N_24923,N_24873);
and UO_2242 (O_2242,N_24448,N_24437);
nand UO_2243 (O_2243,N_24549,N_24665);
xor UO_2244 (O_2244,N_24565,N_24460);
nand UO_2245 (O_2245,N_24945,N_24657);
or UO_2246 (O_2246,N_24541,N_24659);
nor UO_2247 (O_2247,N_24910,N_24912);
nor UO_2248 (O_2248,N_24910,N_24409);
or UO_2249 (O_2249,N_24763,N_24407);
nand UO_2250 (O_2250,N_24857,N_24837);
nor UO_2251 (O_2251,N_24578,N_24991);
and UO_2252 (O_2252,N_24629,N_24669);
nor UO_2253 (O_2253,N_24459,N_24779);
and UO_2254 (O_2254,N_24907,N_24464);
xor UO_2255 (O_2255,N_24589,N_24743);
and UO_2256 (O_2256,N_24692,N_24455);
or UO_2257 (O_2257,N_24965,N_24799);
or UO_2258 (O_2258,N_24901,N_24662);
xnor UO_2259 (O_2259,N_24504,N_24923);
or UO_2260 (O_2260,N_24470,N_24561);
nor UO_2261 (O_2261,N_24730,N_24530);
and UO_2262 (O_2262,N_24760,N_24573);
nor UO_2263 (O_2263,N_24488,N_24931);
and UO_2264 (O_2264,N_24932,N_24492);
and UO_2265 (O_2265,N_24520,N_24508);
xor UO_2266 (O_2266,N_24687,N_24730);
nand UO_2267 (O_2267,N_24406,N_24804);
or UO_2268 (O_2268,N_24582,N_24837);
and UO_2269 (O_2269,N_24414,N_24637);
nor UO_2270 (O_2270,N_24426,N_24989);
and UO_2271 (O_2271,N_24484,N_24927);
xor UO_2272 (O_2272,N_24504,N_24711);
nand UO_2273 (O_2273,N_24560,N_24790);
nor UO_2274 (O_2274,N_24578,N_24698);
or UO_2275 (O_2275,N_24539,N_24591);
and UO_2276 (O_2276,N_24493,N_24471);
and UO_2277 (O_2277,N_24746,N_24661);
nand UO_2278 (O_2278,N_24566,N_24801);
nand UO_2279 (O_2279,N_24827,N_24958);
nor UO_2280 (O_2280,N_24412,N_24858);
nand UO_2281 (O_2281,N_24745,N_24835);
nand UO_2282 (O_2282,N_24480,N_24757);
or UO_2283 (O_2283,N_24805,N_24761);
xnor UO_2284 (O_2284,N_24773,N_24553);
nand UO_2285 (O_2285,N_24906,N_24565);
xor UO_2286 (O_2286,N_24952,N_24922);
or UO_2287 (O_2287,N_24636,N_24451);
and UO_2288 (O_2288,N_24756,N_24619);
nand UO_2289 (O_2289,N_24422,N_24948);
xnor UO_2290 (O_2290,N_24443,N_24417);
nor UO_2291 (O_2291,N_24382,N_24563);
and UO_2292 (O_2292,N_24736,N_24935);
and UO_2293 (O_2293,N_24497,N_24650);
or UO_2294 (O_2294,N_24393,N_24829);
nand UO_2295 (O_2295,N_24739,N_24733);
nand UO_2296 (O_2296,N_24783,N_24563);
or UO_2297 (O_2297,N_24424,N_24771);
and UO_2298 (O_2298,N_24533,N_24795);
nand UO_2299 (O_2299,N_24716,N_24652);
xnor UO_2300 (O_2300,N_24608,N_24735);
nor UO_2301 (O_2301,N_24852,N_24908);
or UO_2302 (O_2302,N_24746,N_24766);
xnor UO_2303 (O_2303,N_24395,N_24724);
nand UO_2304 (O_2304,N_24471,N_24753);
and UO_2305 (O_2305,N_24742,N_24755);
or UO_2306 (O_2306,N_24547,N_24812);
xnor UO_2307 (O_2307,N_24640,N_24845);
nand UO_2308 (O_2308,N_24411,N_24930);
and UO_2309 (O_2309,N_24613,N_24791);
nor UO_2310 (O_2310,N_24485,N_24487);
nand UO_2311 (O_2311,N_24642,N_24949);
and UO_2312 (O_2312,N_24846,N_24381);
and UO_2313 (O_2313,N_24626,N_24724);
and UO_2314 (O_2314,N_24452,N_24812);
or UO_2315 (O_2315,N_24838,N_24468);
or UO_2316 (O_2316,N_24737,N_24881);
and UO_2317 (O_2317,N_24959,N_24763);
xnor UO_2318 (O_2318,N_24619,N_24509);
and UO_2319 (O_2319,N_24665,N_24776);
and UO_2320 (O_2320,N_24723,N_24388);
nor UO_2321 (O_2321,N_24701,N_24601);
nor UO_2322 (O_2322,N_24651,N_24638);
nand UO_2323 (O_2323,N_24937,N_24603);
xor UO_2324 (O_2324,N_24728,N_24878);
xnor UO_2325 (O_2325,N_24975,N_24397);
xnor UO_2326 (O_2326,N_24644,N_24408);
xnor UO_2327 (O_2327,N_24669,N_24652);
xor UO_2328 (O_2328,N_24562,N_24781);
nor UO_2329 (O_2329,N_24574,N_24453);
nor UO_2330 (O_2330,N_24384,N_24615);
nor UO_2331 (O_2331,N_24409,N_24816);
and UO_2332 (O_2332,N_24545,N_24434);
or UO_2333 (O_2333,N_24703,N_24667);
nor UO_2334 (O_2334,N_24872,N_24869);
nor UO_2335 (O_2335,N_24687,N_24918);
nand UO_2336 (O_2336,N_24938,N_24425);
xor UO_2337 (O_2337,N_24662,N_24785);
nand UO_2338 (O_2338,N_24677,N_24977);
nor UO_2339 (O_2339,N_24725,N_24755);
xor UO_2340 (O_2340,N_24919,N_24419);
and UO_2341 (O_2341,N_24885,N_24449);
xor UO_2342 (O_2342,N_24647,N_24978);
and UO_2343 (O_2343,N_24504,N_24524);
nor UO_2344 (O_2344,N_24897,N_24536);
xor UO_2345 (O_2345,N_24542,N_24576);
or UO_2346 (O_2346,N_24442,N_24877);
nor UO_2347 (O_2347,N_24640,N_24669);
xnor UO_2348 (O_2348,N_24641,N_24435);
nor UO_2349 (O_2349,N_24390,N_24870);
and UO_2350 (O_2350,N_24646,N_24528);
nand UO_2351 (O_2351,N_24409,N_24751);
and UO_2352 (O_2352,N_24810,N_24806);
xor UO_2353 (O_2353,N_24457,N_24547);
or UO_2354 (O_2354,N_24468,N_24751);
xnor UO_2355 (O_2355,N_24994,N_24428);
or UO_2356 (O_2356,N_24731,N_24594);
and UO_2357 (O_2357,N_24972,N_24844);
or UO_2358 (O_2358,N_24611,N_24756);
xnor UO_2359 (O_2359,N_24640,N_24902);
nor UO_2360 (O_2360,N_24728,N_24784);
xnor UO_2361 (O_2361,N_24904,N_24730);
and UO_2362 (O_2362,N_24986,N_24972);
xnor UO_2363 (O_2363,N_24681,N_24930);
and UO_2364 (O_2364,N_24666,N_24954);
and UO_2365 (O_2365,N_24688,N_24788);
or UO_2366 (O_2366,N_24622,N_24900);
nand UO_2367 (O_2367,N_24936,N_24763);
xor UO_2368 (O_2368,N_24442,N_24536);
nand UO_2369 (O_2369,N_24873,N_24975);
or UO_2370 (O_2370,N_24978,N_24429);
xnor UO_2371 (O_2371,N_24853,N_24613);
and UO_2372 (O_2372,N_24722,N_24797);
xnor UO_2373 (O_2373,N_24638,N_24769);
and UO_2374 (O_2374,N_24745,N_24761);
nand UO_2375 (O_2375,N_24748,N_24510);
and UO_2376 (O_2376,N_24543,N_24708);
nor UO_2377 (O_2377,N_24910,N_24605);
and UO_2378 (O_2378,N_24732,N_24639);
nor UO_2379 (O_2379,N_24416,N_24932);
or UO_2380 (O_2380,N_24735,N_24912);
and UO_2381 (O_2381,N_24941,N_24914);
nor UO_2382 (O_2382,N_24837,N_24630);
or UO_2383 (O_2383,N_24539,N_24992);
and UO_2384 (O_2384,N_24920,N_24692);
xor UO_2385 (O_2385,N_24643,N_24701);
or UO_2386 (O_2386,N_24753,N_24928);
and UO_2387 (O_2387,N_24921,N_24464);
and UO_2388 (O_2388,N_24429,N_24979);
or UO_2389 (O_2389,N_24792,N_24891);
xor UO_2390 (O_2390,N_24826,N_24779);
nand UO_2391 (O_2391,N_24903,N_24384);
or UO_2392 (O_2392,N_24433,N_24879);
nor UO_2393 (O_2393,N_24714,N_24523);
nand UO_2394 (O_2394,N_24558,N_24546);
or UO_2395 (O_2395,N_24914,N_24482);
or UO_2396 (O_2396,N_24572,N_24427);
nor UO_2397 (O_2397,N_24584,N_24859);
nand UO_2398 (O_2398,N_24613,N_24860);
or UO_2399 (O_2399,N_24472,N_24446);
nor UO_2400 (O_2400,N_24965,N_24959);
xnor UO_2401 (O_2401,N_24864,N_24431);
xnor UO_2402 (O_2402,N_24742,N_24843);
xnor UO_2403 (O_2403,N_24874,N_24883);
nor UO_2404 (O_2404,N_24768,N_24950);
nand UO_2405 (O_2405,N_24455,N_24435);
nor UO_2406 (O_2406,N_24677,N_24467);
nand UO_2407 (O_2407,N_24887,N_24893);
and UO_2408 (O_2408,N_24590,N_24867);
nand UO_2409 (O_2409,N_24722,N_24839);
xnor UO_2410 (O_2410,N_24760,N_24815);
xor UO_2411 (O_2411,N_24392,N_24552);
nand UO_2412 (O_2412,N_24969,N_24954);
nor UO_2413 (O_2413,N_24961,N_24680);
xor UO_2414 (O_2414,N_24763,N_24572);
nand UO_2415 (O_2415,N_24740,N_24671);
nor UO_2416 (O_2416,N_24434,N_24793);
nand UO_2417 (O_2417,N_24590,N_24979);
xnor UO_2418 (O_2418,N_24678,N_24946);
and UO_2419 (O_2419,N_24815,N_24385);
nor UO_2420 (O_2420,N_24756,N_24543);
xor UO_2421 (O_2421,N_24781,N_24509);
and UO_2422 (O_2422,N_24511,N_24393);
xor UO_2423 (O_2423,N_24392,N_24622);
nor UO_2424 (O_2424,N_24394,N_24543);
and UO_2425 (O_2425,N_24833,N_24412);
nor UO_2426 (O_2426,N_24786,N_24550);
and UO_2427 (O_2427,N_24611,N_24897);
or UO_2428 (O_2428,N_24958,N_24546);
or UO_2429 (O_2429,N_24724,N_24852);
or UO_2430 (O_2430,N_24889,N_24733);
nor UO_2431 (O_2431,N_24416,N_24432);
nand UO_2432 (O_2432,N_24723,N_24510);
nor UO_2433 (O_2433,N_24994,N_24703);
nand UO_2434 (O_2434,N_24776,N_24755);
and UO_2435 (O_2435,N_24926,N_24854);
xor UO_2436 (O_2436,N_24435,N_24859);
nor UO_2437 (O_2437,N_24441,N_24972);
nand UO_2438 (O_2438,N_24960,N_24975);
nand UO_2439 (O_2439,N_24563,N_24586);
and UO_2440 (O_2440,N_24447,N_24912);
or UO_2441 (O_2441,N_24426,N_24971);
nand UO_2442 (O_2442,N_24859,N_24715);
xor UO_2443 (O_2443,N_24544,N_24836);
and UO_2444 (O_2444,N_24819,N_24388);
xnor UO_2445 (O_2445,N_24599,N_24609);
and UO_2446 (O_2446,N_24591,N_24675);
or UO_2447 (O_2447,N_24974,N_24425);
nand UO_2448 (O_2448,N_24584,N_24553);
nor UO_2449 (O_2449,N_24665,N_24582);
nor UO_2450 (O_2450,N_24796,N_24382);
or UO_2451 (O_2451,N_24619,N_24684);
and UO_2452 (O_2452,N_24535,N_24888);
nor UO_2453 (O_2453,N_24952,N_24701);
nor UO_2454 (O_2454,N_24774,N_24468);
or UO_2455 (O_2455,N_24625,N_24596);
nand UO_2456 (O_2456,N_24790,N_24893);
xnor UO_2457 (O_2457,N_24410,N_24466);
nand UO_2458 (O_2458,N_24953,N_24845);
xnor UO_2459 (O_2459,N_24599,N_24614);
nand UO_2460 (O_2460,N_24702,N_24975);
xor UO_2461 (O_2461,N_24403,N_24702);
and UO_2462 (O_2462,N_24509,N_24426);
xor UO_2463 (O_2463,N_24641,N_24477);
nand UO_2464 (O_2464,N_24644,N_24467);
xor UO_2465 (O_2465,N_24919,N_24950);
nand UO_2466 (O_2466,N_24740,N_24796);
or UO_2467 (O_2467,N_24430,N_24861);
and UO_2468 (O_2468,N_24538,N_24780);
or UO_2469 (O_2469,N_24900,N_24867);
or UO_2470 (O_2470,N_24588,N_24921);
nand UO_2471 (O_2471,N_24572,N_24935);
nor UO_2472 (O_2472,N_24690,N_24375);
xnor UO_2473 (O_2473,N_24844,N_24518);
or UO_2474 (O_2474,N_24614,N_24632);
nand UO_2475 (O_2475,N_24807,N_24745);
and UO_2476 (O_2476,N_24684,N_24859);
nand UO_2477 (O_2477,N_24836,N_24700);
or UO_2478 (O_2478,N_24951,N_24450);
and UO_2479 (O_2479,N_24523,N_24478);
xnor UO_2480 (O_2480,N_24405,N_24603);
nand UO_2481 (O_2481,N_24403,N_24481);
and UO_2482 (O_2482,N_24715,N_24764);
nand UO_2483 (O_2483,N_24606,N_24750);
nor UO_2484 (O_2484,N_24629,N_24745);
xor UO_2485 (O_2485,N_24875,N_24441);
or UO_2486 (O_2486,N_24621,N_24900);
or UO_2487 (O_2487,N_24443,N_24505);
nand UO_2488 (O_2488,N_24517,N_24872);
nor UO_2489 (O_2489,N_24848,N_24835);
nand UO_2490 (O_2490,N_24945,N_24691);
xor UO_2491 (O_2491,N_24490,N_24517);
nand UO_2492 (O_2492,N_24652,N_24815);
nand UO_2493 (O_2493,N_24438,N_24675);
nor UO_2494 (O_2494,N_24946,N_24798);
nand UO_2495 (O_2495,N_24753,N_24592);
nand UO_2496 (O_2496,N_24795,N_24641);
xor UO_2497 (O_2497,N_24452,N_24798);
nor UO_2498 (O_2498,N_24477,N_24880);
nand UO_2499 (O_2499,N_24427,N_24639);
xnor UO_2500 (O_2500,N_24491,N_24960);
nand UO_2501 (O_2501,N_24538,N_24550);
nor UO_2502 (O_2502,N_24682,N_24731);
nor UO_2503 (O_2503,N_24884,N_24434);
nor UO_2504 (O_2504,N_24920,N_24987);
or UO_2505 (O_2505,N_24861,N_24810);
and UO_2506 (O_2506,N_24867,N_24729);
xnor UO_2507 (O_2507,N_24833,N_24899);
or UO_2508 (O_2508,N_24924,N_24972);
xnor UO_2509 (O_2509,N_24930,N_24625);
nor UO_2510 (O_2510,N_24552,N_24951);
xor UO_2511 (O_2511,N_24579,N_24772);
nand UO_2512 (O_2512,N_24534,N_24813);
nor UO_2513 (O_2513,N_24646,N_24471);
and UO_2514 (O_2514,N_24715,N_24749);
nor UO_2515 (O_2515,N_24888,N_24801);
xnor UO_2516 (O_2516,N_24789,N_24835);
nor UO_2517 (O_2517,N_24409,N_24922);
and UO_2518 (O_2518,N_24478,N_24720);
nor UO_2519 (O_2519,N_24931,N_24769);
and UO_2520 (O_2520,N_24755,N_24985);
nand UO_2521 (O_2521,N_24757,N_24648);
or UO_2522 (O_2522,N_24472,N_24937);
nand UO_2523 (O_2523,N_24879,N_24654);
nor UO_2524 (O_2524,N_24644,N_24801);
xor UO_2525 (O_2525,N_24962,N_24942);
nand UO_2526 (O_2526,N_24969,N_24507);
or UO_2527 (O_2527,N_24499,N_24682);
xnor UO_2528 (O_2528,N_24630,N_24827);
xor UO_2529 (O_2529,N_24952,N_24390);
nand UO_2530 (O_2530,N_24495,N_24484);
or UO_2531 (O_2531,N_24647,N_24612);
and UO_2532 (O_2532,N_24757,N_24826);
nand UO_2533 (O_2533,N_24937,N_24494);
xor UO_2534 (O_2534,N_24923,N_24752);
xor UO_2535 (O_2535,N_24577,N_24759);
and UO_2536 (O_2536,N_24541,N_24977);
or UO_2537 (O_2537,N_24768,N_24735);
and UO_2538 (O_2538,N_24692,N_24991);
nand UO_2539 (O_2539,N_24823,N_24843);
nor UO_2540 (O_2540,N_24881,N_24861);
nand UO_2541 (O_2541,N_24657,N_24513);
xor UO_2542 (O_2542,N_24547,N_24982);
xor UO_2543 (O_2543,N_24858,N_24656);
or UO_2544 (O_2544,N_24436,N_24604);
and UO_2545 (O_2545,N_24883,N_24806);
or UO_2546 (O_2546,N_24639,N_24963);
nand UO_2547 (O_2547,N_24866,N_24603);
or UO_2548 (O_2548,N_24935,N_24997);
nand UO_2549 (O_2549,N_24805,N_24549);
nor UO_2550 (O_2550,N_24433,N_24634);
nand UO_2551 (O_2551,N_24757,N_24694);
nor UO_2552 (O_2552,N_24617,N_24785);
nand UO_2553 (O_2553,N_24549,N_24425);
nor UO_2554 (O_2554,N_24559,N_24902);
and UO_2555 (O_2555,N_24476,N_24957);
and UO_2556 (O_2556,N_24787,N_24921);
and UO_2557 (O_2557,N_24681,N_24644);
and UO_2558 (O_2558,N_24566,N_24670);
nor UO_2559 (O_2559,N_24487,N_24697);
nor UO_2560 (O_2560,N_24756,N_24942);
xnor UO_2561 (O_2561,N_24604,N_24446);
and UO_2562 (O_2562,N_24593,N_24589);
nand UO_2563 (O_2563,N_24768,N_24895);
nor UO_2564 (O_2564,N_24668,N_24528);
nor UO_2565 (O_2565,N_24541,N_24655);
nor UO_2566 (O_2566,N_24916,N_24730);
and UO_2567 (O_2567,N_24958,N_24954);
xor UO_2568 (O_2568,N_24877,N_24469);
xor UO_2569 (O_2569,N_24944,N_24781);
xor UO_2570 (O_2570,N_24739,N_24815);
and UO_2571 (O_2571,N_24620,N_24476);
and UO_2572 (O_2572,N_24653,N_24417);
and UO_2573 (O_2573,N_24469,N_24431);
xor UO_2574 (O_2574,N_24616,N_24892);
nor UO_2575 (O_2575,N_24485,N_24590);
nor UO_2576 (O_2576,N_24852,N_24630);
or UO_2577 (O_2577,N_24878,N_24659);
or UO_2578 (O_2578,N_24872,N_24784);
xnor UO_2579 (O_2579,N_24702,N_24507);
and UO_2580 (O_2580,N_24805,N_24412);
nand UO_2581 (O_2581,N_24649,N_24843);
nand UO_2582 (O_2582,N_24516,N_24610);
xor UO_2583 (O_2583,N_24692,N_24964);
xor UO_2584 (O_2584,N_24619,N_24594);
or UO_2585 (O_2585,N_24852,N_24664);
and UO_2586 (O_2586,N_24377,N_24475);
nor UO_2587 (O_2587,N_24838,N_24952);
or UO_2588 (O_2588,N_24931,N_24492);
nor UO_2589 (O_2589,N_24937,N_24906);
nor UO_2590 (O_2590,N_24862,N_24590);
and UO_2591 (O_2591,N_24613,N_24438);
nor UO_2592 (O_2592,N_24589,N_24715);
nor UO_2593 (O_2593,N_24872,N_24788);
nor UO_2594 (O_2594,N_24834,N_24567);
or UO_2595 (O_2595,N_24841,N_24593);
and UO_2596 (O_2596,N_24586,N_24533);
and UO_2597 (O_2597,N_24939,N_24584);
xor UO_2598 (O_2598,N_24615,N_24735);
or UO_2599 (O_2599,N_24516,N_24425);
nand UO_2600 (O_2600,N_24514,N_24377);
or UO_2601 (O_2601,N_24518,N_24602);
and UO_2602 (O_2602,N_24400,N_24937);
nand UO_2603 (O_2603,N_24822,N_24484);
xnor UO_2604 (O_2604,N_24487,N_24745);
and UO_2605 (O_2605,N_24728,N_24754);
xor UO_2606 (O_2606,N_24875,N_24386);
or UO_2607 (O_2607,N_24438,N_24491);
or UO_2608 (O_2608,N_24680,N_24636);
and UO_2609 (O_2609,N_24419,N_24818);
nor UO_2610 (O_2610,N_24630,N_24834);
xor UO_2611 (O_2611,N_24654,N_24391);
xor UO_2612 (O_2612,N_24723,N_24897);
and UO_2613 (O_2613,N_24855,N_24496);
nand UO_2614 (O_2614,N_24933,N_24414);
and UO_2615 (O_2615,N_24711,N_24526);
nand UO_2616 (O_2616,N_24385,N_24508);
nand UO_2617 (O_2617,N_24581,N_24964);
and UO_2618 (O_2618,N_24590,N_24436);
and UO_2619 (O_2619,N_24750,N_24401);
xnor UO_2620 (O_2620,N_24786,N_24836);
xor UO_2621 (O_2621,N_24775,N_24916);
or UO_2622 (O_2622,N_24800,N_24519);
nor UO_2623 (O_2623,N_24629,N_24710);
xor UO_2624 (O_2624,N_24512,N_24612);
nand UO_2625 (O_2625,N_24811,N_24574);
or UO_2626 (O_2626,N_24480,N_24497);
or UO_2627 (O_2627,N_24814,N_24638);
nor UO_2628 (O_2628,N_24539,N_24694);
xnor UO_2629 (O_2629,N_24899,N_24878);
or UO_2630 (O_2630,N_24912,N_24626);
and UO_2631 (O_2631,N_24389,N_24610);
xor UO_2632 (O_2632,N_24880,N_24932);
xnor UO_2633 (O_2633,N_24612,N_24961);
nor UO_2634 (O_2634,N_24620,N_24806);
nor UO_2635 (O_2635,N_24966,N_24592);
and UO_2636 (O_2636,N_24787,N_24593);
nand UO_2637 (O_2637,N_24737,N_24460);
xnor UO_2638 (O_2638,N_24670,N_24414);
nor UO_2639 (O_2639,N_24780,N_24404);
or UO_2640 (O_2640,N_24797,N_24581);
xor UO_2641 (O_2641,N_24407,N_24840);
or UO_2642 (O_2642,N_24770,N_24961);
nand UO_2643 (O_2643,N_24838,N_24780);
nor UO_2644 (O_2644,N_24401,N_24923);
nor UO_2645 (O_2645,N_24795,N_24732);
nand UO_2646 (O_2646,N_24489,N_24749);
xnor UO_2647 (O_2647,N_24867,N_24481);
or UO_2648 (O_2648,N_24535,N_24903);
xnor UO_2649 (O_2649,N_24424,N_24757);
or UO_2650 (O_2650,N_24972,N_24388);
xnor UO_2651 (O_2651,N_24656,N_24700);
nor UO_2652 (O_2652,N_24481,N_24499);
nor UO_2653 (O_2653,N_24839,N_24772);
and UO_2654 (O_2654,N_24904,N_24561);
or UO_2655 (O_2655,N_24917,N_24741);
nor UO_2656 (O_2656,N_24857,N_24462);
nor UO_2657 (O_2657,N_24466,N_24800);
or UO_2658 (O_2658,N_24716,N_24504);
xor UO_2659 (O_2659,N_24781,N_24660);
xnor UO_2660 (O_2660,N_24659,N_24893);
nor UO_2661 (O_2661,N_24503,N_24895);
nor UO_2662 (O_2662,N_24409,N_24747);
nand UO_2663 (O_2663,N_24606,N_24616);
or UO_2664 (O_2664,N_24571,N_24633);
and UO_2665 (O_2665,N_24740,N_24599);
xor UO_2666 (O_2666,N_24512,N_24384);
nand UO_2667 (O_2667,N_24678,N_24695);
xnor UO_2668 (O_2668,N_24424,N_24449);
nor UO_2669 (O_2669,N_24989,N_24589);
and UO_2670 (O_2670,N_24798,N_24869);
xor UO_2671 (O_2671,N_24816,N_24516);
nand UO_2672 (O_2672,N_24423,N_24799);
or UO_2673 (O_2673,N_24967,N_24524);
and UO_2674 (O_2674,N_24412,N_24715);
or UO_2675 (O_2675,N_24656,N_24688);
and UO_2676 (O_2676,N_24568,N_24862);
or UO_2677 (O_2677,N_24930,N_24604);
nor UO_2678 (O_2678,N_24810,N_24936);
nand UO_2679 (O_2679,N_24859,N_24917);
xnor UO_2680 (O_2680,N_24440,N_24635);
nor UO_2681 (O_2681,N_24560,N_24891);
xor UO_2682 (O_2682,N_24734,N_24820);
and UO_2683 (O_2683,N_24591,N_24387);
and UO_2684 (O_2684,N_24712,N_24824);
or UO_2685 (O_2685,N_24641,N_24860);
nand UO_2686 (O_2686,N_24821,N_24670);
xnor UO_2687 (O_2687,N_24503,N_24822);
and UO_2688 (O_2688,N_24701,N_24977);
nand UO_2689 (O_2689,N_24517,N_24601);
nand UO_2690 (O_2690,N_24523,N_24928);
nand UO_2691 (O_2691,N_24717,N_24511);
nand UO_2692 (O_2692,N_24551,N_24448);
nand UO_2693 (O_2693,N_24963,N_24767);
and UO_2694 (O_2694,N_24957,N_24678);
xnor UO_2695 (O_2695,N_24980,N_24817);
nand UO_2696 (O_2696,N_24532,N_24674);
or UO_2697 (O_2697,N_24449,N_24928);
or UO_2698 (O_2698,N_24584,N_24722);
nor UO_2699 (O_2699,N_24787,N_24415);
nand UO_2700 (O_2700,N_24772,N_24656);
nor UO_2701 (O_2701,N_24389,N_24776);
xnor UO_2702 (O_2702,N_24799,N_24596);
nand UO_2703 (O_2703,N_24426,N_24572);
xor UO_2704 (O_2704,N_24844,N_24730);
nor UO_2705 (O_2705,N_24585,N_24433);
and UO_2706 (O_2706,N_24793,N_24874);
nor UO_2707 (O_2707,N_24772,N_24687);
xnor UO_2708 (O_2708,N_24394,N_24399);
nor UO_2709 (O_2709,N_24834,N_24859);
nor UO_2710 (O_2710,N_24808,N_24603);
or UO_2711 (O_2711,N_24467,N_24551);
nor UO_2712 (O_2712,N_24865,N_24440);
nand UO_2713 (O_2713,N_24817,N_24710);
xnor UO_2714 (O_2714,N_24970,N_24596);
nand UO_2715 (O_2715,N_24592,N_24780);
nor UO_2716 (O_2716,N_24459,N_24825);
nor UO_2717 (O_2717,N_24439,N_24538);
nand UO_2718 (O_2718,N_24867,N_24647);
or UO_2719 (O_2719,N_24713,N_24615);
or UO_2720 (O_2720,N_24415,N_24978);
nand UO_2721 (O_2721,N_24945,N_24488);
nor UO_2722 (O_2722,N_24607,N_24456);
and UO_2723 (O_2723,N_24670,N_24948);
and UO_2724 (O_2724,N_24906,N_24416);
and UO_2725 (O_2725,N_24383,N_24958);
nand UO_2726 (O_2726,N_24637,N_24574);
or UO_2727 (O_2727,N_24393,N_24700);
nand UO_2728 (O_2728,N_24919,N_24506);
nor UO_2729 (O_2729,N_24461,N_24944);
nor UO_2730 (O_2730,N_24646,N_24501);
nand UO_2731 (O_2731,N_24960,N_24408);
xnor UO_2732 (O_2732,N_24715,N_24530);
or UO_2733 (O_2733,N_24590,N_24377);
nor UO_2734 (O_2734,N_24934,N_24852);
xor UO_2735 (O_2735,N_24382,N_24451);
and UO_2736 (O_2736,N_24684,N_24745);
nand UO_2737 (O_2737,N_24576,N_24916);
nand UO_2738 (O_2738,N_24873,N_24856);
or UO_2739 (O_2739,N_24731,N_24897);
and UO_2740 (O_2740,N_24479,N_24400);
or UO_2741 (O_2741,N_24963,N_24594);
xnor UO_2742 (O_2742,N_24664,N_24405);
or UO_2743 (O_2743,N_24414,N_24576);
and UO_2744 (O_2744,N_24682,N_24695);
xnor UO_2745 (O_2745,N_24826,N_24426);
nor UO_2746 (O_2746,N_24445,N_24456);
nor UO_2747 (O_2747,N_24558,N_24895);
nor UO_2748 (O_2748,N_24791,N_24506);
xor UO_2749 (O_2749,N_24561,N_24553);
nor UO_2750 (O_2750,N_24522,N_24541);
nor UO_2751 (O_2751,N_24688,N_24924);
nand UO_2752 (O_2752,N_24825,N_24411);
nand UO_2753 (O_2753,N_24427,N_24788);
nor UO_2754 (O_2754,N_24867,N_24799);
and UO_2755 (O_2755,N_24501,N_24445);
xnor UO_2756 (O_2756,N_24808,N_24594);
nand UO_2757 (O_2757,N_24493,N_24563);
nor UO_2758 (O_2758,N_24534,N_24623);
nand UO_2759 (O_2759,N_24719,N_24859);
or UO_2760 (O_2760,N_24497,N_24820);
nand UO_2761 (O_2761,N_24999,N_24420);
nor UO_2762 (O_2762,N_24861,N_24524);
or UO_2763 (O_2763,N_24689,N_24748);
or UO_2764 (O_2764,N_24465,N_24945);
xnor UO_2765 (O_2765,N_24398,N_24991);
xor UO_2766 (O_2766,N_24434,N_24823);
or UO_2767 (O_2767,N_24544,N_24669);
or UO_2768 (O_2768,N_24552,N_24537);
or UO_2769 (O_2769,N_24916,N_24899);
or UO_2770 (O_2770,N_24881,N_24423);
nor UO_2771 (O_2771,N_24618,N_24626);
xnor UO_2772 (O_2772,N_24821,N_24572);
nand UO_2773 (O_2773,N_24763,N_24579);
xor UO_2774 (O_2774,N_24451,N_24680);
nand UO_2775 (O_2775,N_24734,N_24782);
and UO_2776 (O_2776,N_24775,N_24542);
nor UO_2777 (O_2777,N_24531,N_24974);
xor UO_2778 (O_2778,N_24845,N_24495);
nor UO_2779 (O_2779,N_24402,N_24473);
xnor UO_2780 (O_2780,N_24942,N_24488);
nor UO_2781 (O_2781,N_24745,N_24558);
and UO_2782 (O_2782,N_24663,N_24751);
or UO_2783 (O_2783,N_24739,N_24500);
nand UO_2784 (O_2784,N_24595,N_24692);
xor UO_2785 (O_2785,N_24828,N_24466);
or UO_2786 (O_2786,N_24496,N_24447);
and UO_2787 (O_2787,N_24897,N_24654);
xnor UO_2788 (O_2788,N_24506,N_24881);
or UO_2789 (O_2789,N_24794,N_24492);
or UO_2790 (O_2790,N_24618,N_24615);
or UO_2791 (O_2791,N_24967,N_24633);
or UO_2792 (O_2792,N_24543,N_24414);
and UO_2793 (O_2793,N_24642,N_24517);
nor UO_2794 (O_2794,N_24758,N_24947);
or UO_2795 (O_2795,N_24406,N_24854);
xnor UO_2796 (O_2796,N_24990,N_24442);
xor UO_2797 (O_2797,N_24925,N_24963);
nand UO_2798 (O_2798,N_24529,N_24629);
nand UO_2799 (O_2799,N_24970,N_24976);
or UO_2800 (O_2800,N_24657,N_24896);
and UO_2801 (O_2801,N_24731,N_24969);
nor UO_2802 (O_2802,N_24825,N_24721);
xnor UO_2803 (O_2803,N_24491,N_24901);
nor UO_2804 (O_2804,N_24447,N_24653);
xnor UO_2805 (O_2805,N_24500,N_24762);
or UO_2806 (O_2806,N_24502,N_24914);
or UO_2807 (O_2807,N_24949,N_24538);
or UO_2808 (O_2808,N_24421,N_24561);
xor UO_2809 (O_2809,N_24566,N_24734);
nand UO_2810 (O_2810,N_24712,N_24717);
or UO_2811 (O_2811,N_24526,N_24857);
nor UO_2812 (O_2812,N_24957,N_24471);
and UO_2813 (O_2813,N_24447,N_24776);
or UO_2814 (O_2814,N_24908,N_24941);
xor UO_2815 (O_2815,N_24894,N_24944);
nand UO_2816 (O_2816,N_24400,N_24798);
or UO_2817 (O_2817,N_24721,N_24943);
nand UO_2818 (O_2818,N_24668,N_24855);
or UO_2819 (O_2819,N_24681,N_24538);
xor UO_2820 (O_2820,N_24688,N_24501);
nor UO_2821 (O_2821,N_24620,N_24983);
nor UO_2822 (O_2822,N_24725,N_24969);
xor UO_2823 (O_2823,N_24784,N_24503);
nor UO_2824 (O_2824,N_24594,N_24793);
nand UO_2825 (O_2825,N_24709,N_24595);
nor UO_2826 (O_2826,N_24882,N_24750);
or UO_2827 (O_2827,N_24753,N_24799);
nand UO_2828 (O_2828,N_24823,N_24796);
nor UO_2829 (O_2829,N_24925,N_24771);
or UO_2830 (O_2830,N_24995,N_24951);
nand UO_2831 (O_2831,N_24826,N_24486);
and UO_2832 (O_2832,N_24502,N_24724);
nor UO_2833 (O_2833,N_24424,N_24752);
or UO_2834 (O_2834,N_24627,N_24619);
and UO_2835 (O_2835,N_24812,N_24716);
nand UO_2836 (O_2836,N_24689,N_24883);
or UO_2837 (O_2837,N_24645,N_24889);
or UO_2838 (O_2838,N_24411,N_24941);
xnor UO_2839 (O_2839,N_24428,N_24471);
xor UO_2840 (O_2840,N_24638,N_24434);
nand UO_2841 (O_2841,N_24870,N_24453);
and UO_2842 (O_2842,N_24404,N_24770);
xor UO_2843 (O_2843,N_24800,N_24931);
nand UO_2844 (O_2844,N_24789,N_24927);
nor UO_2845 (O_2845,N_24883,N_24850);
and UO_2846 (O_2846,N_24534,N_24868);
and UO_2847 (O_2847,N_24518,N_24972);
and UO_2848 (O_2848,N_24559,N_24542);
xnor UO_2849 (O_2849,N_24422,N_24441);
nor UO_2850 (O_2850,N_24917,N_24442);
xor UO_2851 (O_2851,N_24698,N_24850);
and UO_2852 (O_2852,N_24632,N_24843);
xor UO_2853 (O_2853,N_24937,N_24626);
xnor UO_2854 (O_2854,N_24995,N_24639);
nand UO_2855 (O_2855,N_24671,N_24859);
and UO_2856 (O_2856,N_24375,N_24634);
and UO_2857 (O_2857,N_24874,N_24384);
nor UO_2858 (O_2858,N_24583,N_24860);
nand UO_2859 (O_2859,N_24699,N_24461);
nand UO_2860 (O_2860,N_24971,N_24435);
nand UO_2861 (O_2861,N_24785,N_24774);
or UO_2862 (O_2862,N_24840,N_24920);
and UO_2863 (O_2863,N_24798,N_24924);
nand UO_2864 (O_2864,N_24751,N_24917);
or UO_2865 (O_2865,N_24476,N_24735);
and UO_2866 (O_2866,N_24627,N_24552);
nand UO_2867 (O_2867,N_24467,N_24726);
or UO_2868 (O_2868,N_24794,N_24448);
nand UO_2869 (O_2869,N_24861,N_24926);
nor UO_2870 (O_2870,N_24595,N_24637);
nand UO_2871 (O_2871,N_24890,N_24885);
and UO_2872 (O_2872,N_24739,N_24833);
nor UO_2873 (O_2873,N_24887,N_24749);
and UO_2874 (O_2874,N_24855,N_24618);
or UO_2875 (O_2875,N_24420,N_24606);
or UO_2876 (O_2876,N_24450,N_24400);
nor UO_2877 (O_2877,N_24678,N_24783);
xnor UO_2878 (O_2878,N_24642,N_24734);
nor UO_2879 (O_2879,N_24451,N_24942);
and UO_2880 (O_2880,N_24605,N_24982);
or UO_2881 (O_2881,N_24418,N_24603);
and UO_2882 (O_2882,N_24941,N_24964);
and UO_2883 (O_2883,N_24395,N_24733);
nor UO_2884 (O_2884,N_24678,N_24922);
or UO_2885 (O_2885,N_24375,N_24684);
and UO_2886 (O_2886,N_24436,N_24576);
xor UO_2887 (O_2887,N_24813,N_24605);
nor UO_2888 (O_2888,N_24855,N_24569);
and UO_2889 (O_2889,N_24668,N_24927);
nor UO_2890 (O_2890,N_24999,N_24456);
xnor UO_2891 (O_2891,N_24880,N_24554);
or UO_2892 (O_2892,N_24575,N_24819);
or UO_2893 (O_2893,N_24519,N_24683);
and UO_2894 (O_2894,N_24933,N_24881);
or UO_2895 (O_2895,N_24447,N_24672);
nand UO_2896 (O_2896,N_24460,N_24466);
and UO_2897 (O_2897,N_24804,N_24801);
nand UO_2898 (O_2898,N_24656,N_24377);
or UO_2899 (O_2899,N_24607,N_24921);
nand UO_2900 (O_2900,N_24741,N_24891);
nor UO_2901 (O_2901,N_24721,N_24790);
and UO_2902 (O_2902,N_24736,N_24388);
xnor UO_2903 (O_2903,N_24435,N_24498);
and UO_2904 (O_2904,N_24949,N_24911);
nor UO_2905 (O_2905,N_24436,N_24386);
or UO_2906 (O_2906,N_24599,N_24874);
xnor UO_2907 (O_2907,N_24813,N_24870);
and UO_2908 (O_2908,N_24381,N_24712);
xnor UO_2909 (O_2909,N_24673,N_24388);
xor UO_2910 (O_2910,N_24870,N_24715);
nand UO_2911 (O_2911,N_24887,N_24707);
xor UO_2912 (O_2912,N_24924,N_24708);
nor UO_2913 (O_2913,N_24551,N_24958);
nor UO_2914 (O_2914,N_24981,N_24770);
nand UO_2915 (O_2915,N_24394,N_24659);
xor UO_2916 (O_2916,N_24760,N_24715);
nand UO_2917 (O_2917,N_24677,N_24861);
and UO_2918 (O_2918,N_24638,N_24711);
xor UO_2919 (O_2919,N_24388,N_24408);
or UO_2920 (O_2920,N_24408,N_24867);
nor UO_2921 (O_2921,N_24849,N_24408);
and UO_2922 (O_2922,N_24505,N_24824);
nand UO_2923 (O_2923,N_24519,N_24817);
nor UO_2924 (O_2924,N_24863,N_24818);
and UO_2925 (O_2925,N_24691,N_24786);
xor UO_2926 (O_2926,N_24989,N_24913);
and UO_2927 (O_2927,N_24638,N_24695);
nor UO_2928 (O_2928,N_24599,N_24581);
nor UO_2929 (O_2929,N_24754,N_24922);
and UO_2930 (O_2930,N_24978,N_24971);
and UO_2931 (O_2931,N_24799,N_24636);
or UO_2932 (O_2932,N_24743,N_24629);
and UO_2933 (O_2933,N_24957,N_24413);
and UO_2934 (O_2934,N_24674,N_24467);
xnor UO_2935 (O_2935,N_24531,N_24451);
xor UO_2936 (O_2936,N_24758,N_24694);
nor UO_2937 (O_2937,N_24566,N_24789);
xnor UO_2938 (O_2938,N_24569,N_24657);
nor UO_2939 (O_2939,N_24899,N_24946);
nand UO_2940 (O_2940,N_24619,N_24408);
nor UO_2941 (O_2941,N_24959,N_24589);
nor UO_2942 (O_2942,N_24377,N_24605);
nand UO_2943 (O_2943,N_24795,N_24464);
xnor UO_2944 (O_2944,N_24996,N_24535);
or UO_2945 (O_2945,N_24806,N_24761);
and UO_2946 (O_2946,N_24722,N_24856);
and UO_2947 (O_2947,N_24821,N_24679);
and UO_2948 (O_2948,N_24809,N_24829);
nor UO_2949 (O_2949,N_24920,N_24565);
and UO_2950 (O_2950,N_24646,N_24635);
nand UO_2951 (O_2951,N_24617,N_24555);
and UO_2952 (O_2952,N_24409,N_24801);
xnor UO_2953 (O_2953,N_24423,N_24865);
xor UO_2954 (O_2954,N_24565,N_24719);
or UO_2955 (O_2955,N_24429,N_24448);
nor UO_2956 (O_2956,N_24966,N_24962);
xnor UO_2957 (O_2957,N_24795,N_24481);
xnor UO_2958 (O_2958,N_24983,N_24493);
or UO_2959 (O_2959,N_24408,N_24539);
xor UO_2960 (O_2960,N_24540,N_24627);
nand UO_2961 (O_2961,N_24597,N_24562);
nor UO_2962 (O_2962,N_24646,N_24982);
nand UO_2963 (O_2963,N_24740,N_24621);
nor UO_2964 (O_2964,N_24726,N_24644);
nor UO_2965 (O_2965,N_24620,N_24780);
and UO_2966 (O_2966,N_24422,N_24865);
xor UO_2967 (O_2967,N_24678,N_24663);
nand UO_2968 (O_2968,N_24961,N_24767);
nand UO_2969 (O_2969,N_24836,N_24984);
nor UO_2970 (O_2970,N_24762,N_24528);
nor UO_2971 (O_2971,N_24730,N_24637);
xor UO_2972 (O_2972,N_24996,N_24406);
and UO_2973 (O_2973,N_24866,N_24498);
nand UO_2974 (O_2974,N_24467,N_24488);
nor UO_2975 (O_2975,N_24400,N_24889);
nor UO_2976 (O_2976,N_24816,N_24933);
xor UO_2977 (O_2977,N_24740,N_24679);
and UO_2978 (O_2978,N_24514,N_24543);
nor UO_2979 (O_2979,N_24904,N_24457);
or UO_2980 (O_2980,N_24380,N_24946);
nand UO_2981 (O_2981,N_24456,N_24570);
xnor UO_2982 (O_2982,N_24559,N_24985);
nand UO_2983 (O_2983,N_24642,N_24708);
or UO_2984 (O_2984,N_24995,N_24978);
nand UO_2985 (O_2985,N_24982,N_24631);
nand UO_2986 (O_2986,N_24685,N_24517);
or UO_2987 (O_2987,N_24657,N_24959);
nand UO_2988 (O_2988,N_24381,N_24603);
and UO_2989 (O_2989,N_24706,N_24892);
and UO_2990 (O_2990,N_24962,N_24598);
nor UO_2991 (O_2991,N_24950,N_24767);
xnor UO_2992 (O_2992,N_24631,N_24408);
or UO_2993 (O_2993,N_24471,N_24814);
xor UO_2994 (O_2994,N_24618,N_24827);
xor UO_2995 (O_2995,N_24967,N_24942);
and UO_2996 (O_2996,N_24601,N_24936);
or UO_2997 (O_2997,N_24838,N_24622);
xnor UO_2998 (O_2998,N_24833,N_24982);
nand UO_2999 (O_2999,N_24443,N_24688);
endmodule