module basic_750_5000_1000_2_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2512,N_2516,N_2517,N_2518,N_2519,N_2520,N_2522,N_2523,N_2525,N_2526,N_2527,N_2528,N_2530,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2540,N_2541,N_2542,N_2543,N_2544,N_2546,N_2547,N_2549,N_2550,N_2551,N_2554,N_2555,N_2556,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2567,N_2568,N_2570,N_2571,N_2573,N_2575,N_2576,N_2577,N_2578,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2596,N_2597,N_2598,N_2599,N_2601,N_2603,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2617,N_2618,N_2620,N_2621,N_2622,N_2625,N_2627,N_2628,N_2629,N_2630,N_2632,N_2633,N_2634,N_2636,N_2638,N_2640,N_2642,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2661,N_2662,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2712,N_2713,N_2714,N_2715,N_2717,N_2718,N_2719,N_2720,N_2724,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2753,N_2756,N_2757,N_2759,N_2760,N_2761,N_2763,N_2764,N_2766,N_2768,N_2769,N_2770,N_2771,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2793,N_2794,N_2795,N_2796,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2816,N_2817,N_2818,N_2819,N_2822,N_2823,N_2824,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2836,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2845,N_2846,N_2848,N_2849,N_2850,N_2851,N_2852,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2873,N_2874,N_2875,N_2877,N_2878,N_2879,N_2880,N_2881,N_2883,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2896,N_2897,N_2898,N_2900,N_2901,N_2902,N_2903,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2922,N_2923,N_2924,N_2926,N_2928,N_2929,N_2930,N_2931,N_2932,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2942,N_2944,N_2945,N_2946,N_2947,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2962,N_2963,N_2964,N_2965,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2975,N_2976,N_2978,N_2980,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_3000,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3016,N_3017,N_3019,N_3020,N_3021,N_3022,N_3025,N_3026,N_3028,N_3030,N_3031,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3052,N_3053,N_3054,N_3055,N_3056,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3067,N_3068,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3087,N_3089,N_3090,N_3091,N_3093,N_3094,N_3095,N_3096,N_3098,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3116,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3138,N_3139,N_3140,N_3142,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3195,N_3196,N_3197,N_3199,N_3200,N_3203,N_3204,N_3207,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3230,N_3231,N_3232,N_3234,N_3236,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3269,N_3270,N_3272,N_3273,N_3275,N_3276,N_3277,N_3278,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3294,N_3295,N_3297,N_3298,N_3300,N_3301,N_3302,N_3303,N_3305,N_3308,N_3309,N_3310,N_3312,N_3314,N_3315,N_3316,N_3317,N_3318,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3329,N_3331,N_3332,N_3334,N_3335,N_3336,N_3338,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3356,N_3357,N_3359,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3369,N_3370,N_3372,N_3373,N_3374,N_3375,N_3376,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3404,N_3407,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3416,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3448,N_3450,N_3451,N_3454,N_3456,N_3457,N_3459,N_3460,N_3462,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3472,N_3473,N_3475,N_3477,N_3478,N_3480,N_3481,N_3482,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3511,N_3512,N_3513,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3525,N_3526,N_3527,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3537,N_3538,N_3540,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3556,N_3558,N_3559,N_3560,N_3561,N_3562,N_3564,N_3565,N_3567,N_3568,N_3569,N_3570,N_3572,N_3574,N_3575,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3587,N_3588,N_3592,N_3593,N_3594,N_3596,N_3598,N_3599,N_3600,N_3601,N_3602,N_3605,N_3606,N_3607,N_3609,N_3610,N_3612,N_3613,N_3614,N_3616,N_3617,N_3618,N_3619,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3640,N_3641,N_3643,N_3644,N_3645,N_3646,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3657,N_3658,N_3659,N_3660,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3674,N_3675,N_3676,N_3678,N_3679,N_3680,N_3682,N_3683,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3707,N_3708,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3728,N_3729,N_3730,N_3731,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3745,N_3746,N_3747,N_3748,N_3749,N_3752,N_3753,N_3755,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3788,N_3789,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3814,N_3815,N_3816,N_3818,N_3819,N_3820,N_3821,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3840,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3861,N_3862,N_3864,N_3865,N_3866,N_3868,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3879,N_3882,N_3883,N_3886,N_3887,N_3888,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3900,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3909,N_3910,N_3911,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3920,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3943,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3971,N_3973,N_3975,N_3976,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3993,N_3994,N_3998,N_3999,N_4000,N_4001,N_4003,N_4004,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4021,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4034,N_4035,N_4036,N_4039,N_4040,N_4041,N_4042,N_4043,N_4045,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4065,N_4066,N_4067,N_4069,N_4070,N_4072,N_4073,N_4074,N_4075,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4086,N_4087,N_4088,N_4089,N_4090,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4104,N_4105,N_4106,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4120,N_4121,N_4122,N_4123,N_4124,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4136,N_4137,N_4138,N_4140,N_4141,N_4142,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4153,N_4155,N_4156,N_4157,N_4158,N_4160,N_4161,N_4162,N_4163,N_4164,N_4166,N_4167,N_4168,N_4169,N_4171,N_4172,N_4173,N_4174,N_4176,N_4177,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4189,N_4190,N_4191,N_4192,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4202,N_4203,N_4204,N_4205,N_4207,N_4208,N_4209,N_4210,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4227,N_4228,N_4230,N_4231,N_4233,N_4234,N_4235,N_4236,N_4237,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4254,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4286,N_4287,N_4288,N_4290,N_4291,N_4292,N_4293,N_4294,N_4296,N_4297,N_4298,N_4300,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4315,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4339,N_4340,N_4341,N_4342,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4382,N_4383,N_4384,N_4385,N_4387,N_4388,N_4389,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4399,N_4400,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4440,N_4443,N_4444,N_4445,N_4446,N_4448,N_4449,N_4450,N_4451,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4472,N_4473,N_4474,N_4477,N_4478,N_4481,N_4482,N_4483,N_4484,N_4486,N_4487,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4496,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4515,N_4517,N_4518,N_4519,N_4520,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4529,N_4530,N_4531,N_4532,N_4533,N_4535,N_4537,N_4538,N_4539,N_4540,N_4542,N_4545,N_4546,N_4547,N_4548,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4568,N_4573,N_4575,N_4576,N_4577,N_4578,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4601,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4612,N_4613,N_4614,N_4616,N_4617,N_4620,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4631,N_4632,N_4633,N_4634,N_4635,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4654,N_4655,N_4656,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4668,N_4669,N_4671,N_4672,N_4673,N_4674,N_4677,N_4678,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4707,N_4708,N_4709,N_4710,N_4712,N_4713,N_4716,N_4717,N_4718,N_4720,N_4721,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4730,N_4731,N_4734,N_4735,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4748,N_4749,N_4750,N_4753,N_4755,N_4756,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4765,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4778,N_4780,N_4781,N_4782,N_4784,N_4785,N_4786,N_4787,N_4789,N_4790,N_4791,N_4792,N_4796,N_4797,N_4800,N_4801,N_4805,N_4807,N_4808,N_4809,N_4811,N_4812,N_4814,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4826,N_4827,N_4828,N_4829,N_4830,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4839,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4855,N_4856,N_4857,N_4858,N_4859,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4874,N_4875,N_4876,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4894,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4905,N_4906,N_4907,N_4908,N_4910,N_4911,N_4912,N_4913,N_4914,N_4916,N_4918,N_4919,N_4920,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4948,N_4949,N_4950,N_4951,N_4953,N_4956,N_4957,N_4958,N_4959,N_4962,N_4965,N_4966,N_4967,N_4968,N_4970,N_4971,N_4972,N_4973,N_4975,N_4977,N_4978,N_4980,N_4981,N_4982,N_4985,N_4988,N_4989,N_4991,N_4992,N_4994,N_4995,N_4997,N_4998,N_4999;
nor U0 (N_0,In_317,In_229);
nand U1 (N_1,In_202,In_621);
or U2 (N_2,In_501,In_97);
nand U3 (N_3,In_337,In_710);
nand U4 (N_4,In_51,In_165);
and U5 (N_5,In_577,In_392);
nor U6 (N_6,In_103,In_705);
nor U7 (N_7,In_595,In_480);
nand U8 (N_8,In_167,In_45);
nand U9 (N_9,In_401,In_358);
and U10 (N_10,In_459,In_110);
or U11 (N_11,In_38,In_302);
or U12 (N_12,In_84,In_277);
or U13 (N_13,In_406,In_518);
nor U14 (N_14,In_515,In_101);
or U15 (N_15,In_367,In_386);
or U16 (N_16,In_136,In_275);
nand U17 (N_17,In_464,In_677);
or U18 (N_18,In_570,In_409);
or U19 (N_19,In_19,In_525);
and U20 (N_20,In_373,In_379);
or U21 (N_21,In_81,In_419);
and U22 (N_22,In_179,In_296);
or U23 (N_23,In_531,In_697);
nand U24 (N_24,In_173,In_711);
nand U25 (N_25,In_55,In_224);
nor U26 (N_26,In_481,In_635);
and U27 (N_27,In_550,In_478);
nand U28 (N_28,In_345,In_408);
or U29 (N_29,In_495,In_100);
or U30 (N_30,In_633,In_16);
or U31 (N_31,In_238,In_685);
or U32 (N_32,In_605,In_511);
nand U33 (N_33,In_598,In_215);
or U34 (N_34,In_643,In_145);
and U35 (N_35,In_143,In_484);
or U36 (N_36,In_382,In_311);
and U37 (N_37,In_542,In_32);
nand U38 (N_38,In_407,In_79);
nand U39 (N_39,In_551,In_727);
and U40 (N_40,In_673,In_395);
nand U41 (N_41,In_323,In_613);
nor U42 (N_42,In_660,In_470);
xnor U43 (N_43,In_329,In_606);
or U44 (N_44,In_290,In_712);
or U45 (N_45,In_394,In_76);
and U46 (N_46,In_522,In_371);
or U47 (N_47,In_69,In_618);
or U48 (N_48,In_144,In_342);
nor U49 (N_49,In_225,In_61);
nand U50 (N_50,In_429,In_295);
and U51 (N_51,In_370,In_365);
nor U52 (N_52,In_562,In_509);
and U53 (N_53,In_161,In_403);
nand U54 (N_54,In_194,In_380);
nor U55 (N_55,In_502,In_310);
xnor U56 (N_56,In_280,In_252);
or U57 (N_57,In_230,In_472);
or U58 (N_58,In_738,In_182);
nand U59 (N_59,In_266,In_695);
and U60 (N_60,In_183,In_322);
nor U61 (N_61,In_546,In_418);
nor U62 (N_62,In_92,In_284);
nand U63 (N_63,In_324,In_232);
or U64 (N_64,In_421,In_314);
nor U65 (N_65,In_514,In_628);
and U66 (N_66,In_734,In_554);
nand U67 (N_67,In_244,In_0);
nor U68 (N_68,In_544,In_684);
and U69 (N_69,In_30,In_29);
nor U70 (N_70,In_652,In_216);
or U71 (N_71,In_288,In_616);
and U72 (N_72,In_474,In_354);
nand U73 (N_73,In_485,In_294);
nor U74 (N_74,In_552,In_350);
nand U75 (N_75,In_453,In_339);
nor U76 (N_76,In_490,In_548);
nand U77 (N_77,In_125,In_438);
nor U78 (N_78,In_188,In_178);
nor U79 (N_79,In_739,In_447);
nor U80 (N_80,In_220,In_368);
and U81 (N_81,In_217,In_483);
nand U82 (N_82,In_22,In_261);
nor U83 (N_83,In_579,In_471);
nor U84 (N_84,In_547,In_247);
and U85 (N_85,In_720,In_571);
nand U86 (N_86,In_190,In_78);
nand U87 (N_87,In_309,In_576);
or U88 (N_88,In_132,In_398);
nor U89 (N_89,In_469,In_431);
nor U90 (N_90,In_328,In_640);
and U91 (N_91,In_538,In_71);
nand U92 (N_92,In_59,In_332);
nor U93 (N_93,In_463,In_87);
nor U94 (N_94,In_535,In_653);
and U95 (N_95,In_199,In_413);
nand U96 (N_96,In_213,In_638);
nor U97 (N_97,In_6,In_718);
nor U98 (N_98,In_211,In_164);
nand U99 (N_99,In_286,In_208);
nor U100 (N_100,In_135,In_526);
nor U101 (N_101,In_214,In_253);
nand U102 (N_102,In_42,In_320);
nor U103 (N_103,In_661,In_270);
nand U104 (N_104,In_376,In_316);
nand U105 (N_105,In_9,In_257);
or U106 (N_106,In_675,In_326);
nor U107 (N_107,In_96,In_475);
nand U108 (N_108,In_708,In_505);
and U109 (N_109,In_404,In_93);
nor U110 (N_110,In_37,In_555);
and U111 (N_111,In_40,In_352);
nand U112 (N_112,In_581,In_111);
nand U113 (N_113,In_427,In_636);
and U114 (N_114,In_107,In_556);
or U115 (N_115,In_2,In_619);
or U116 (N_116,In_597,In_749);
and U117 (N_117,In_665,In_489);
or U118 (N_118,In_428,In_558);
nor U119 (N_119,In_434,In_693);
nand U120 (N_120,In_351,In_1);
and U121 (N_121,In_48,In_251);
or U122 (N_122,In_246,In_264);
nand U123 (N_123,In_433,In_703);
or U124 (N_124,In_692,In_493);
nand U125 (N_125,In_702,In_44);
or U126 (N_126,In_644,In_707);
and U127 (N_127,In_35,In_155);
or U128 (N_128,In_271,In_362);
or U129 (N_129,In_701,In_601);
nor U130 (N_130,In_612,In_249);
and U131 (N_131,In_713,In_443);
nor U132 (N_132,In_455,In_654);
or U133 (N_133,In_139,In_435);
or U134 (N_134,In_282,In_686);
nand U135 (N_135,In_527,In_304);
nand U136 (N_136,In_212,In_565);
xnor U137 (N_137,In_70,In_627);
nand U138 (N_138,In_651,In_742);
nor U139 (N_139,In_709,In_449);
or U140 (N_140,In_385,In_85);
and U141 (N_141,In_735,In_670);
and U142 (N_142,In_451,In_11);
or U143 (N_143,In_440,In_344);
or U144 (N_144,In_250,In_115);
nand U145 (N_145,In_159,In_667);
or U146 (N_146,In_426,In_436);
or U147 (N_147,In_587,In_584);
nor U148 (N_148,In_624,In_72);
nand U149 (N_149,In_133,In_620);
and U150 (N_150,In_27,In_729);
nor U151 (N_151,In_89,In_414);
and U152 (N_152,In_355,In_726);
nor U153 (N_153,In_321,In_245);
or U154 (N_154,In_561,In_530);
nand U155 (N_155,In_402,In_108);
or U156 (N_156,In_637,In_596);
or U157 (N_157,In_346,In_461);
and U158 (N_158,In_679,In_491);
or U159 (N_159,In_719,In_539);
nor U160 (N_160,In_218,In_26);
and U161 (N_161,In_348,In_457);
nand U162 (N_162,In_534,In_98);
and U163 (N_163,In_174,In_241);
and U164 (N_164,In_13,In_333);
and U165 (N_165,In_566,In_417);
and U166 (N_166,In_121,In_671);
or U167 (N_167,In_338,In_390);
nand U168 (N_168,In_528,In_73);
nand U169 (N_169,In_240,In_682);
nor U170 (N_170,In_383,In_147);
nand U171 (N_171,In_88,In_31);
nor U172 (N_172,In_313,In_99);
nor U173 (N_173,In_192,In_722);
and U174 (N_174,In_140,In_169);
nand U175 (N_175,In_142,In_510);
and U176 (N_176,In_617,In_196);
nand U177 (N_177,In_114,In_151);
and U178 (N_178,In_152,In_715);
nand U179 (N_179,In_123,In_185);
or U180 (N_180,In_500,In_156);
or U181 (N_181,In_248,In_122);
or U182 (N_182,In_649,In_582);
or U183 (N_183,In_118,In_378);
nand U184 (N_184,In_126,In_425);
and U185 (N_185,In_209,In_423);
nor U186 (N_186,In_590,In_393);
nand U187 (N_187,In_743,In_634);
nand U188 (N_188,In_14,In_442);
and U189 (N_189,In_728,In_458);
nor U190 (N_190,In_293,In_492);
or U191 (N_191,In_256,In_517);
nand U192 (N_192,In_267,In_460);
nand U193 (N_193,In_327,In_521);
nor U194 (N_194,In_23,In_691);
and U195 (N_195,In_177,In_242);
xor U196 (N_196,In_53,In_353);
xor U197 (N_197,In_391,In_319);
or U198 (N_198,In_243,In_39);
nand U199 (N_199,In_529,In_357);
and U200 (N_200,In_662,In_171);
nand U201 (N_201,In_137,In_415);
nand U202 (N_202,In_630,In_564);
or U203 (N_203,In_255,In_462);
and U204 (N_204,In_396,In_519);
nor U205 (N_205,In_669,In_34);
and U206 (N_206,In_681,In_54);
nor U207 (N_207,In_659,In_52);
nor U208 (N_208,In_674,In_235);
nor U209 (N_209,In_600,In_77);
and U210 (N_210,In_520,In_102);
nor U211 (N_211,In_149,In_721);
and U212 (N_212,In_334,In_153);
nand U213 (N_213,In_283,In_74);
nand U214 (N_214,In_113,In_359);
nor U215 (N_215,In_746,In_732);
nand U216 (N_216,In_306,In_441);
or U217 (N_217,In_331,In_83);
and U218 (N_218,In_205,In_377);
and U219 (N_219,In_58,In_273);
and U220 (N_220,In_172,In_268);
nand U221 (N_221,In_274,In_698);
and U222 (N_222,In_642,In_7);
nor U223 (N_223,In_128,In_399);
nor U224 (N_224,In_374,In_731);
and U225 (N_225,In_592,In_303);
nand U226 (N_226,In_523,In_237);
or U227 (N_227,In_347,In_615);
and U228 (N_228,In_513,In_154);
nand U229 (N_229,In_593,In_387);
nor U230 (N_230,In_18,In_725);
and U231 (N_231,In_170,In_315);
nor U232 (N_232,In_747,In_678);
and U233 (N_233,In_536,In_664);
nor U234 (N_234,In_305,In_599);
and U235 (N_235,In_210,In_646);
xor U236 (N_236,In_278,In_714);
or U237 (N_237,In_532,In_400);
and U238 (N_238,In_405,In_25);
nand U239 (N_239,In_625,In_160);
nor U240 (N_240,In_696,In_559);
nor U241 (N_241,In_437,In_176);
or U242 (N_242,In_200,In_384);
or U243 (N_243,In_325,In_467);
nand U244 (N_244,In_704,In_560);
and U245 (N_245,In_219,In_254);
and U246 (N_246,In_341,In_263);
and U247 (N_247,In_363,In_629);
and U248 (N_248,In_609,In_279);
xor U249 (N_249,In_668,In_446);
or U250 (N_250,In_297,In_448);
nand U251 (N_251,In_90,In_388);
xnor U252 (N_252,In_411,In_737);
nand U253 (N_253,In_572,In_687);
nor U254 (N_254,In_195,In_496);
and U255 (N_255,In_226,In_588);
nand U256 (N_256,In_468,In_507);
nor U257 (N_257,In_187,In_138);
nor U258 (N_258,In_336,In_207);
and U259 (N_259,In_260,In_360);
or U260 (N_260,In_62,In_723);
and U261 (N_261,In_583,In_580);
nand U262 (N_262,In_308,In_745);
and U263 (N_263,In_477,In_676);
and U264 (N_264,In_228,In_589);
or U265 (N_265,In_197,In_281);
nor U266 (N_266,In_206,In_222);
nand U267 (N_267,In_389,In_80);
or U268 (N_268,In_504,In_129);
nor U269 (N_269,In_64,In_569);
and U270 (N_270,In_15,In_330);
nor U271 (N_271,In_553,In_131);
and U272 (N_272,In_4,In_416);
or U273 (N_273,In_680,In_689);
nor U274 (N_274,In_444,In_198);
nand U275 (N_275,In_239,In_41);
or U276 (N_276,In_163,In_366);
or U277 (N_277,In_650,In_65);
or U278 (N_278,In_227,In_432);
nand U279 (N_279,In_75,In_655);
nand U280 (N_280,In_20,In_412);
or U281 (N_281,In_186,In_318);
and U282 (N_282,In_748,In_473);
nand U283 (N_283,In_307,In_568);
nor U284 (N_284,In_86,In_632);
or U285 (N_285,In_47,In_201);
and U286 (N_286,In_381,In_603);
nand U287 (N_287,In_109,In_586);
nor U288 (N_288,In_94,In_666);
xnor U289 (N_289,In_10,In_486);
nand U290 (N_290,In_508,In_68);
and U291 (N_291,In_312,In_361);
xor U292 (N_292,In_12,In_291);
or U293 (N_293,In_567,In_541);
nor U294 (N_294,In_607,In_614);
nor U295 (N_295,In_104,In_700);
nand U296 (N_296,In_631,In_193);
or U297 (N_297,In_744,In_503);
xnor U298 (N_298,In_690,In_298);
or U299 (N_299,In_540,In_641);
nand U300 (N_300,In_5,In_658);
or U301 (N_301,In_730,In_130);
and U302 (N_302,In_49,In_424);
nor U303 (N_303,In_46,In_33);
or U304 (N_304,In_119,In_694);
nor U305 (N_305,In_549,In_465);
and U306 (N_306,In_66,In_120);
nor U307 (N_307,In_112,In_258);
or U308 (N_308,In_231,In_639);
nor U309 (N_309,In_91,In_56);
or U310 (N_310,In_466,In_439);
and U311 (N_311,In_657,In_494);
nor U312 (N_312,In_106,In_223);
nand U313 (N_313,In_604,In_236);
or U314 (N_314,In_364,In_397);
nand U315 (N_315,In_656,In_299);
nor U316 (N_316,In_533,In_146);
nor U317 (N_317,In_168,In_623);
nor U318 (N_318,In_375,In_602);
nand U319 (N_319,In_28,In_272);
or U320 (N_320,In_116,In_482);
nor U321 (N_321,In_82,In_63);
or U322 (N_322,In_573,In_292);
or U323 (N_323,In_716,In_706);
or U324 (N_324,In_516,In_134);
or U325 (N_325,In_608,In_105);
or U326 (N_326,In_578,In_343);
nand U327 (N_327,In_626,In_150);
nand U328 (N_328,In_148,In_349);
and U329 (N_329,In_512,In_124);
nor U330 (N_330,In_157,In_454);
nand U331 (N_331,In_594,In_672);
xnor U332 (N_332,In_203,In_479);
and U333 (N_333,In_610,In_184);
nand U334 (N_334,In_233,In_741);
nor U335 (N_335,In_189,In_234);
nand U336 (N_336,In_557,In_175);
nor U337 (N_337,In_162,In_356);
nor U338 (N_338,In_24,In_127);
and U339 (N_339,In_497,In_21);
nor U340 (N_340,In_488,In_17);
and U341 (N_341,In_545,In_648);
and U342 (N_342,In_499,In_166);
nor U343 (N_343,In_3,In_300);
and U344 (N_344,In_287,In_585);
or U345 (N_345,In_269,In_699);
xnor U346 (N_346,In_733,In_335);
xor U347 (N_347,In_141,In_591);
and U348 (N_348,In_180,In_191);
or U349 (N_349,In_340,In_717);
nand U350 (N_350,In_420,In_611);
nand U351 (N_351,In_683,In_204);
and U352 (N_352,In_221,In_8);
and U353 (N_353,In_476,In_259);
xnor U354 (N_354,In_524,In_563);
and U355 (N_355,In_487,In_181);
nand U356 (N_356,In_301,In_740);
and U357 (N_357,In_647,In_422);
and U358 (N_358,In_67,In_450);
nand U359 (N_359,In_724,In_117);
nand U360 (N_360,In_57,In_645);
nor U361 (N_361,In_95,In_574);
or U362 (N_362,In_430,In_537);
and U363 (N_363,In_43,In_285);
nor U364 (N_364,In_736,In_410);
nor U365 (N_365,In_452,In_663);
nand U366 (N_366,In_622,In_575);
and U367 (N_367,In_506,In_688);
and U368 (N_368,In_445,In_50);
and U369 (N_369,In_369,In_158);
or U370 (N_370,In_276,In_36);
nand U371 (N_371,In_372,In_265);
or U372 (N_372,In_456,In_498);
nand U373 (N_373,In_60,In_289);
nor U374 (N_374,In_543,In_262);
or U375 (N_375,In_116,In_642);
nand U376 (N_376,In_685,In_157);
nand U377 (N_377,In_54,In_627);
and U378 (N_378,In_741,In_277);
and U379 (N_379,In_116,In_581);
or U380 (N_380,In_383,In_126);
and U381 (N_381,In_212,In_552);
nand U382 (N_382,In_496,In_420);
and U383 (N_383,In_475,In_452);
nand U384 (N_384,In_601,In_625);
nor U385 (N_385,In_635,In_198);
nor U386 (N_386,In_690,In_646);
and U387 (N_387,In_448,In_377);
nand U388 (N_388,In_539,In_199);
nand U389 (N_389,In_560,In_143);
and U390 (N_390,In_369,In_135);
or U391 (N_391,In_484,In_718);
nor U392 (N_392,In_211,In_368);
or U393 (N_393,In_134,In_665);
or U394 (N_394,In_635,In_347);
and U395 (N_395,In_189,In_548);
nand U396 (N_396,In_98,In_689);
nor U397 (N_397,In_472,In_4);
nand U398 (N_398,In_350,In_533);
or U399 (N_399,In_631,In_387);
and U400 (N_400,In_469,In_201);
nor U401 (N_401,In_259,In_451);
and U402 (N_402,In_267,In_129);
or U403 (N_403,In_622,In_2);
or U404 (N_404,In_706,In_111);
nand U405 (N_405,In_266,In_637);
nand U406 (N_406,In_532,In_570);
or U407 (N_407,In_100,In_622);
or U408 (N_408,In_98,In_499);
or U409 (N_409,In_608,In_683);
nor U410 (N_410,In_262,In_604);
nand U411 (N_411,In_529,In_123);
nor U412 (N_412,In_386,In_606);
nor U413 (N_413,In_268,In_417);
nand U414 (N_414,In_733,In_299);
nor U415 (N_415,In_748,In_654);
and U416 (N_416,In_336,In_31);
nand U417 (N_417,In_722,In_316);
or U418 (N_418,In_173,In_497);
and U419 (N_419,In_559,In_256);
or U420 (N_420,In_432,In_558);
and U421 (N_421,In_661,In_74);
or U422 (N_422,In_470,In_201);
xnor U423 (N_423,In_505,In_613);
nor U424 (N_424,In_569,In_93);
nand U425 (N_425,In_345,In_556);
nand U426 (N_426,In_649,In_396);
or U427 (N_427,In_140,In_48);
nor U428 (N_428,In_344,In_135);
nand U429 (N_429,In_331,In_245);
nand U430 (N_430,In_8,In_182);
and U431 (N_431,In_562,In_143);
or U432 (N_432,In_135,In_472);
nor U433 (N_433,In_556,In_427);
or U434 (N_434,In_474,In_255);
nor U435 (N_435,In_572,In_160);
nor U436 (N_436,In_352,In_299);
and U437 (N_437,In_676,In_479);
and U438 (N_438,In_578,In_225);
nor U439 (N_439,In_27,In_491);
or U440 (N_440,In_633,In_331);
nor U441 (N_441,In_495,In_373);
or U442 (N_442,In_644,In_651);
or U443 (N_443,In_478,In_42);
nor U444 (N_444,In_318,In_308);
nand U445 (N_445,In_615,In_296);
or U446 (N_446,In_702,In_488);
or U447 (N_447,In_117,In_326);
and U448 (N_448,In_649,In_62);
xnor U449 (N_449,In_579,In_83);
nor U450 (N_450,In_159,In_315);
nor U451 (N_451,In_199,In_20);
nor U452 (N_452,In_348,In_571);
nand U453 (N_453,In_134,In_540);
nand U454 (N_454,In_702,In_400);
or U455 (N_455,In_672,In_597);
and U456 (N_456,In_256,In_246);
or U457 (N_457,In_326,In_515);
and U458 (N_458,In_402,In_210);
or U459 (N_459,In_390,In_172);
nor U460 (N_460,In_566,In_257);
or U461 (N_461,In_43,In_588);
nand U462 (N_462,In_583,In_637);
and U463 (N_463,In_505,In_378);
nand U464 (N_464,In_123,In_358);
nand U465 (N_465,In_369,In_527);
nand U466 (N_466,In_113,In_265);
nand U467 (N_467,In_527,In_655);
and U468 (N_468,In_138,In_213);
nand U469 (N_469,In_294,In_626);
and U470 (N_470,In_34,In_82);
nor U471 (N_471,In_544,In_745);
or U472 (N_472,In_652,In_298);
and U473 (N_473,In_655,In_672);
nand U474 (N_474,In_218,In_437);
and U475 (N_475,In_220,In_696);
and U476 (N_476,In_336,In_551);
or U477 (N_477,In_404,In_205);
nand U478 (N_478,In_586,In_77);
nor U479 (N_479,In_285,In_356);
nand U480 (N_480,In_266,In_700);
nand U481 (N_481,In_386,In_372);
nand U482 (N_482,In_231,In_223);
nor U483 (N_483,In_3,In_677);
and U484 (N_484,In_612,In_686);
and U485 (N_485,In_254,In_661);
nor U486 (N_486,In_287,In_269);
nor U487 (N_487,In_251,In_576);
nor U488 (N_488,In_711,In_29);
and U489 (N_489,In_716,In_51);
nand U490 (N_490,In_654,In_575);
and U491 (N_491,In_624,In_5);
and U492 (N_492,In_724,In_586);
nand U493 (N_493,In_706,In_83);
nand U494 (N_494,In_247,In_402);
nand U495 (N_495,In_536,In_74);
and U496 (N_496,In_163,In_619);
xnor U497 (N_497,In_234,In_145);
or U498 (N_498,In_92,In_611);
and U499 (N_499,In_111,In_568);
and U500 (N_500,In_306,In_310);
nand U501 (N_501,In_399,In_123);
and U502 (N_502,In_351,In_532);
and U503 (N_503,In_150,In_714);
nand U504 (N_504,In_605,In_444);
and U505 (N_505,In_413,In_308);
nand U506 (N_506,In_313,In_435);
xor U507 (N_507,In_651,In_355);
xnor U508 (N_508,In_293,In_60);
nand U509 (N_509,In_49,In_494);
and U510 (N_510,In_321,In_575);
or U511 (N_511,In_227,In_632);
and U512 (N_512,In_624,In_558);
nand U513 (N_513,In_508,In_253);
nand U514 (N_514,In_75,In_366);
and U515 (N_515,In_82,In_443);
nor U516 (N_516,In_124,In_350);
nor U517 (N_517,In_469,In_400);
nor U518 (N_518,In_312,In_317);
and U519 (N_519,In_729,In_644);
and U520 (N_520,In_127,In_208);
or U521 (N_521,In_28,In_652);
nor U522 (N_522,In_100,In_414);
or U523 (N_523,In_677,In_137);
or U524 (N_524,In_459,In_44);
nand U525 (N_525,In_460,In_512);
or U526 (N_526,In_343,In_202);
and U527 (N_527,In_375,In_257);
and U528 (N_528,In_355,In_433);
and U529 (N_529,In_46,In_254);
and U530 (N_530,In_503,In_413);
nor U531 (N_531,In_243,In_171);
or U532 (N_532,In_537,In_85);
nor U533 (N_533,In_554,In_647);
and U534 (N_534,In_154,In_437);
and U535 (N_535,In_260,In_492);
nor U536 (N_536,In_566,In_166);
nand U537 (N_537,In_44,In_531);
nor U538 (N_538,In_320,In_449);
nor U539 (N_539,In_350,In_413);
and U540 (N_540,In_2,In_504);
and U541 (N_541,In_390,In_375);
nand U542 (N_542,In_641,In_345);
or U543 (N_543,In_415,In_595);
xnor U544 (N_544,In_418,In_662);
nand U545 (N_545,In_291,In_583);
and U546 (N_546,In_229,In_724);
and U547 (N_547,In_637,In_593);
or U548 (N_548,In_169,In_172);
nand U549 (N_549,In_458,In_344);
and U550 (N_550,In_200,In_302);
nand U551 (N_551,In_382,In_399);
or U552 (N_552,In_146,In_251);
or U553 (N_553,In_350,In_106);
and U554 (N_554,In_520,In_505);
nor U555 (N_555,In_548,In_266);
and U556 (N_556,In_250,In_524);
and U557 (N_557,In_672,In_443);
nor U558 (N_558,In_175,In_330);
xor U559 (N_559,In_621,In_580);
nor U560 (N_560,In_379,In_96);
or U561 (N_561,In_713,In_414);
and U562 (N_562,In_2,In_446);
and U563 (N_563,In_721,In_454);
xor U564 (N_564,In_683,In_481);
nand U565 (N_565,In_367,In_394);
nand U566 (N_566,In_221,In_341);
nand U567 (N_567,In_270,In_169);
nand U568 (N_568,In_264,In_499);
nand U569 (N_569,In_193,In_441);
and U570 (N_570,In_470,In_613);
or U571 (N_571,In_625,In_390);
nand U572 (N_572,In_394,In_669);
or U573 (N_573,In_168,In_17);
or U574 (N_574,In_562,In_335);
nor U575 (N_575,In_688,In_603);
or U576 (N_576,In_736,In_229);
and U577 (N_577,In_582,In_526);
and U578 (N_578,In_674,In_288);
nor U579 (N_579,In_496,In_648);
nand U580 (N_580,In_585,In_607);
nand U581 (N_581,In_599,In_315);
and U582 (N_582,In_284,In_115);
or U583 (N_583,In_12,In_20);
nand U584 (N_584,In_75,In_257);
nor U585 (N_585,In_650,In_340);
nand U586 (N_586,In_178,In_27);
and U587 (N_587,In_518,In_265);
and U588 (N_588,In_4,In_443);
nor U589 (N_589,In_509,In_453);
or U590 (N_590,In_577,In_248);
xor U591 (N_591,In_133,In_86);
nor U592 (N_592,In_229,In_671);
or U593 (N_593,In_672,In_289);
nand U594 (N_594,In_291,In_99);
nand U595 (N_595,In_240,In_441);
or U596 (N_596,In_175,In_423);
nor U597 (N_597,In_377,In_36);
or U598 (N_598,In_342,In_126);
nor U599 (N_599,In_725,In_108);
and U600 (N_600,In_537,In_619);
xnor U601 (N_601,In_318,In_702);
nor U602 (N_602,In_631,In_474);
nand U603 (N_603,In_471,In_372);
nand U604 (N_604,In_299,In_407);
and U605 (N_605,In_693,In_510);
or U606 (N_606,In_465,In_433);
nand U607 (N_607,In_398,In_427);
or U608 (N_608,In_265,In_129);
nor U609 (N_609,In_481,In_2);
and U610 (N_610,In_453,In_689);
nand U611 (N_611,In_81,In_139);
nor U612 (N_612,In_532,In_438);
or U613 (N_613,In_156,In_287);
nand U614 (N_614,In_354,In_356);
nor U615 (N_615,In_550,In_25);
nand U616 (N_616,In_747,In_397);
nand U617 (N_617,In_332,In_221);
nor U618 (N_618,In_539,In_80);
or U619 (N_619,In_488,In_575);
nor U620 (N_620,In_683,In_20);
nand U621 (N_621,In_372,In_563);
or U622 (N_622,In_652,In_293);
nand U623 (N_623,In_39,In_748);
or U624 (N_624,In_230,In_108);
or U625 (N_625,In_530,In_8);
or U626 (N_626,In_283,In_718);
and U627 (N_627,In_41,In_410);
and U628 (N_628,In_129,In_577);
and U629 (N_629,In_448,In_260);
or U630 (N_630,In_108,In_62);
or U631 (N_631,In_99,In_565);
nor U632 (N_632,In_519,In_419);
and U633 (N_633,In_508,In_428);
and U634 (N_634,In_43,In_203);
or U635 (N_635,In_546,In_306);
and U636 (N_636,In_467,In_276);
and U637 (N_637,In_692,In_684);
nand U638 (N_638,In_105,In_74);
and U639 (N_639,In_704,In_312);
or U640 (N_640,In_403,In_356);
nor U641 (N_641,In_581,In_613);
or U642 (N_642,In_348,In_73);
nor U643 (N_643,In_592,In_272);
nand U644 (N_644,In_724,In_507);
or U645 (N_645,In_89,In_307);
nand U646 (N_646,In_185,In_706);
or U647 (N_647,In_280,In_489);
nor U648 (N_648,In_276,In_536);
and U649 (N_649,In_559,In_592);
xnor U650 (N_650,In_367,In_359);
and U651 (N_651,In_171,In_349);
and U652 (N_652,In_745,In_445);
or U653 (N_653,In_333,In_209);
nand U654 (N_654,In_545,In_184);
nand U655 (N_655,In_467,In_105);
nand U656 (N_656,In_309,In_333);
and U657 (N_657,In_609,In_425);
and U658 (N_658,In_292,In_451);
nand U659 (N_659,In_295,In_371);
and U660 (N_660,In_583,In_345);
or U661 (N_661,In_501,In_564);
nand U662 (N_662,In_581,In_690);
or U663 (N_663,In_717,In_377);
nand U664 (N_664,In_196,In_8);
nand U665 (N_665,In_308,In_133);
nand U666 (N_666,In_430,In_61);
nand U667 (N_667,In_161,In_686);
nand U668 (N_668,In_260,In_418);
or U669 (N_669,In_728,In_509);
and U670 (N_670,In_609,In_674);
nand U671 (N_671,In_341,In_637);
and U672 (N_672,In_131,In_402);
and U673 (N_673,In_161,In_215);
or U674 (N_674,In_12,In_538);
and U675 (N_675,In_246,In_253);
nand U676 (N_676,In_431,In_561);
or U677 (N_677,In_76,In_96);
nor U678 (N_678,In_635,In_181);
and U679 (N_679,In_589,In_314);
and U680 (N_680,In_7,In_102);
and U681 (N_681,In_85,In_515);
nand U682 (N_682,In_209,In_231);
nor U683 (N_683,In_633,In_78);
nand U684 (N_684,In_372,In_641);
nor U685 (N_685,In_374,In_491);
and U686 (N_686,In_113,In_246);
and U687 (N_687,In_75,In_86);
and U688 (N_688,In_33,In_394);
or U689 (N_689,In_618,In_341);
and U690 (N_690,In_187,In_133);
nand U691 (N_691,In_722,In_616);
nand U692 (N_692,In_129,In_164);
or U693 (N_693,In_287,In_548);
nor U694 (N_694,In_486,In_467);
nand U695 (N_695,In_181,In_540);
nand U696 (N_696,In_232,In_523);
nor U697 (N_697,In_563,In_628);
nor U698 (N_698,In_166,In_367);
or U699 (N_699,In_650,In_592);
and U700 (N_700,In_219,In_678);
nor U701 (N_701,In_10,In_407);
nand U702 (N_702,In_643,In_345);
nor U703 (N_703,In_184,In_467);
nand U704 (N_704,In_214,In_411);
or U705 (N_705,In_52,In_182);
nor U706 (N_706,In_408,In_503);
and U707 (N_707,In_58,In_140);
and U708 (N_708,In_558,In_505);
nor U709 (N_709,In_261,In_601);
nand U710 (N_710,In_633,In_530);
nor U711 (N_711,In_107,In_217);
and U712 (N_712,In_515,In_627);
nor U713 (N_713,In_690,In_476);
nand U714 (N_714,In_82,In_105);
nor U715 (N_715,In_549,In_512);
or U716 (N_716,In_721,In_258);
xor U717 (N_717,In_602,In_569);
nor U718 (N_718,In_724,In_159);
or U719 (N_719,In_721,In_140);
or U720 (N_720,In_360,In_313);
and U721 (N_721,In_344,In_383);
and U722 (N_722,In_273,In_628);
nor U723 (N_723,In_493,In_536);
nand U724 (N_724,In_40,In_557);
and U725 (N_725,In_103,In_639);
nor U726 (N_726,In_746,In_191);
nor U727 (N_727,In_220,In_319);
nor U728 (N_728,In_680,In_2);
nand U729 (N_729,In_484,In_2);
and U730 (N_730,In_86,In_464);
nand U731 (N_731,In_484,In_235);
nor U732 (N_732,In_75,In_378);
nor U733 (N_733,In_523,In_604);
and U734 (N_734,In_157,In_325);
nor U735 (N_735,In_650,In_140);
or U736 (N_736,In_269,In_104);
or U737 (N_737,In_537,In_110);
and U738 (N_738,In_145,In_660);
nor U739 (N_739,In_379,In_135);
nor U740 (N_740,In_483,In_230);
xnor U741 (N_741,In_735,In_537);
nand U742 (N_742,In_285,In_637);
or U743 (N_743,In_481,In_656);
nand U744 (N_744,In_164,In_286);
or U745 (N_745,In_598,In_373);
nor U746 (N_746,In_159,In_624);
or U747 (N_747,In_379,In_239);
xor U748 (N_748,In_273,In_572);
nand U749 (N_749,In_213,In_497);
or U750 (N_750,In_512,In_613);
or U751 (N_751,In_404,In_723);
and U752 (N_752,In_179,In_102);
nand U753 (N_753,In_207,In_257);
and U754 (N_754,In_419,In_714);
and U755 (N_755,In_325,In_545);
or U756 (N_756,In_344,In_599);
and U757 (N_757,In_144,In_579);
and U758 (N_758,In_688,In_282);
or U759 (N_759,In_423,In_58);
nand U760 (N_760,In_453,In_222);
nand U761 (N_761,In_128,In_479);
or U762 (N_762,In_146,In_294);
nand U763 (N_763,In_468,In_585);
and U764 (N_764,In_602,In_663);
nand U765 (N_765,In_460,In_222);
nor U766 (N_766,In_244,In_453);
and U767 (N_767,In_369,In_47);
nor U768 (N_768,In_322,In_626);
or U769 (N_769,In_420,In_648);
nor U770 (N_770,In_300,In_65);
and U771 (N_771,In_631,In_209);
and U772 (N_772,In_593,In_429);
or U773 (N_773,In_131,In_55);
or U774 (N_774,In_268,In_60);
nor U775 (N_775,In_81,In_392);
nor U776 (N_776,In_56,In_124);
nor U777 (N_777,In_330,In_526);
nor U778 (N_778,In_565,In_625);
nor U779 (N_779,In_232,In_564);
nand U780 (N_780,In_480,In_441);
nand U781 (N_781,In_244,In_399);
nor U782 (N_782,In_90,In_315);
nand U783 (N_783,In_152,In_367);
nor U784 (N_784,In_688,In_281);
or U785 (N_785,In_588,In_675);
and U786 (N_786,In_131,In_679);
nand U787 (N_787,In_348,In_443);
nand U788 (N_788,In_452,In_493);
or U789 (N_789,In_648,In_233);
nor U790 (N_790,In_80,In_50);
nand U791 (N_791,In_676,In_128);
and U792 (N_792,In_163,In_321);
and U793 (N_793,In_371,In_57);
nand U794 (N_794,In_511,In_134);
nor U795 (N_795,In_676,In_470);
and U796 (N_796,In_549,In_183);
nor U797 (N_797,In_298,In_421);
or U798 (N_798,In_336,In_238);
nor U799 (N_799,In_489,In_536);
or U800 (N_800,In_97,In_707);
nand U801 (N_801,In_665,In_446);
nor U802 (N_802,In_653,In_663);
nor U803 (N_803,In_189,In_112);
nor U804 (N_804,In_105,In_487);
or U805 (N_805,In_447,In_702);
or U806 (N_806,In_169,In_162);
nor U807 (N_807,In_692,In_351);
or U808 (N_808,In_473,In_93);
nor U809 (N_809,In_736,In_264);
nor U810 (N_810,In_213,In_46);
nand U811 (N_811,In_470,In_644);
or U812 (N_812,In_164,In_75);
nor U813 (N_813,In_306,In_504);
and U814 (N_814,In_69,In_558);
or U815 (N_815,In_728,In_576);
or U816 (N_816,In_236,In_91);
nor U817 (N_817,In_566,In_366);
nand U818 (N_818,In_350,In_539);
and U819 (N_819,In_527,In_348);
and U820 (N_820,In_502,In_603);
xnor U821 (N_821,In_223,In_260);
or U822 (N_822,In_266,In_366);
or U823 (N_823,In_626,In_257);
or U824 (N_824,In_249,In_358);
and U825 (N_825,In_689,In_522);
nor U826 (N_826,In_279,In_523);
nand U827 (N_827,In_534,In_71);
nor U828 (N_828,In_469,In_335);
nand U829 (N_829,In_377,In_111);
nor U830 (N_830,In_209,In_308);
or U831 (N_831,In_73,In_378);
or U832 (N_832,In_743,In_748);
or U833 (N_833,In_215,In_614);
nand U834 (N_834,In_569,In_483);
nor U835 (N_835,In_64,In_290);
nand U836 (N_836,In_254,In_165);
and U837 (N_837,In_456,In_273);
or U838 (N_838,In_736,In_349);
nor U839 (N_839,In_678,In_9);
or U840 (N_840,In_162,In_727);
and U841 (N_841,In_513,In_239);
nand U842 (N_842,In_537,In_348);
or U843 (N_843,In_442,In_406);
nor U844 (N_844,In_87,In_556);
nand U845 (N_845,In_458,In_62);
and U846 (N_846,In_612,In_351);
nand U847 (N_847,In_325,In_254);
and U848 (N_848,In_129,In_418);
or U849 (N_849,In_193,In_108);
and U850 (N_850,In_490,In_355);
nand U851 (N_851,In_662,In_163);
or U852 (N_852,In_259,In_678);
or U853 (N_853,In_607,In_135);
and U854 (N_854,In_620,In_610);
and U855 (N_855,In_246,In_616);
nand U856 (N_856,In_119,In_142);
nor U857 (N_857,In_96,In_632);
nor U858 (N_858,In_59,In_570);
or U859 (N_859,In_341,In_332);
and U860 (N_860,In_429,In_156);
nand U861 (N_861,In_722,In_12);
or U862 (N_862,In_257,In_654);
nor U863 (N_863,In_1,In_517);
and U864 (N_864,In_118,In_736);
nor U865 (N_865,In_508,In_204);
and U866 (N_866,In_424,In_433);
nor U867 (N_867,In_725,In_562);
nand U868 (N_868,In_417,In_212);
and U869 (N_869,In_252,In_493);
or U870 (N_870,In_586,In_0);
or U871 (N_871,In_371,In_230);
nor U872 (N_872,In_270,In_721);
or U873 (N_873,In_459,In_495);
nor U874 (N_874,In_365,In_571);
or U875 (N_875,In_344,In_111);
nor U876 (N_876,In_306,In_242);
nand U877 (N_877,In_704,In_56);
and U878 (N_878,In_188,In_360);
nor U879 (N_879,In_215,In_296);
and U880 (N_880,In_88,In_712);
and U881 (N_881,In_77,In_93);
and U882 (N_882,In_276,In_229);
nand U883 (N_883,In_629,In_9);
nand U884 (N_884,In_80,In_232);
or U885 (N_885,In_578,In_395);
and U886 (N_886,In_507,In_463);
and U887 (N_887,In_13,In_5);
nand U888 (N_888,In_335,In_129);
nand U889 (N_889,In_731,In_713);
or U890 (N_890,In_653,In_659);
nor U891 (N_891,In_304,In_182);
and U892 (N_892,In_92,In_653);
or U893 (N_893,In_689,In_234);
or U894 (N_894,In_252,In_154);
nor U895 (N_895,In_211,In_502);
nand U896 (N_896,In_717,In_645);
nor U897 (N_897,In_467,In_111);
nor U898 (N_898,In_122,In_44);
nor U899 (N_899,In_427,In_159);
nor U900 (N_900,In_503,In_8);
nand U901 (N_901,In_216,In_508);
and U902 (N_902,In_615,In_543);
nor U903 (N_903,In_115,In_544);
or U904 (N_904,In_271,In_618);
and U905 (N_905,In_649,In_536);
or U906 (N_906,In_108,In_579);
nor U907 (N_907,In_474,In_622);
nand U908 (N_908,In_401,In_238);
or U909 (N_909,In_272,In_411);
nor U910 (N_910,In_475,In_309);
or U911 (N_911,In_466,In_370);
nand U912 (N_912,In_275,In_402);
or U913 (N_913,In_747,In_583);
or U914 (N_914,In_469,In_553);
or U915 (N_915,In_11,In_499);
and U916 (N_916,In_165,In_559);
or U917 (N_917,In_301,In_79);
nor U918 (N_918,In_646,In_514);
and U919 (N_919,In_449,In_70);
and U920 (N_920,In_463,In_289);
nor U921 (N_921,In_656,In_729);
nor U922 (N_922,In_166,In_160);
and U923 (N_923,In_588,In_567);
nand U924 (N_924,In_411,In_228);
nand U925 (N_925,In_455,In_170);
nor U926 (N_926,In_614,In_740);
and U927 (N_927,In_527,In_532);
nand U928 (N_928,In_413,In_291);
or U929 (N_929,In_290,In_321);
nor U930 (N_930,In_190,In_73);
or U931 (N_931,In_575,In_602);
nand U932 (N_932,In_439,In_572);
and U933 (N_933,In_504,In_51);
nor U934 (N_934,In_543,In_645);
or U935 (N_935,In_29,In_109);
and U936 (N_936,In_374,In_248);
and U937 (N_937,In_127,In_82);
xor U938 (N_938,In_387,In_336);
and U939 (N_939,In_749,In_507);
or U940 (N_940,In_104,In_102);
nor U941 (N_941,In_458,In_448);
nor U942 (N_942,In_422,In_494);
nand U943 (N_943,In_187,In_289);
nand U944 (N_944,In_480,In_368);
and U945 (N_945,In_554,In_728);
and U946 (N_946,In_214,In_364);
nor U947 (N_947,In_621,In_128);
and U948 (N_948,In_503,In_352);
nor U949 (N_949,In_597,In_588);
nand U950 (N_950,In_295,In_694);
nor U951 (N_951,In_106,In_635);
and U952 (N_952,In_119,In_253);
nand U953 (N_953,In_541,In_508);
and U954 (N_954,In_430,In_227);
nor U955 (N_955,In_101,In_531);
or U956 (N_956,In_257,In_167);
and U957 (N_957,In_179,In_468);
or U958 (N_958,In_458,In_139);
and U959 (N_959,In_103,In_676);
and U960 (N_960,In_653,In_726);
nand U961 (N_961,In_510,In_672);
nor U962 (N_962,In_272,In_86);
or U963 (N_963,In_654,In_446);
or U964 (N_964,In_589,In_9);
or U965 (N_965,In_642,In_303);
nor U966 (N_966,In_285,In_661);
xnor U967 (N_967,In_706,In_355);
nand U968 (N_968,In_348,In_642);
and U969 (N_969,In_620,In_74);
or U970 (N_970,In_345,In_684);
nand U971 (N_971,In_369,In_240);
nand U972 (N_972,In_472,In_125);
nor U973 (N_973,In_61,In_127);
nand U974 (N_974,In_44,In_295);
and U975 (N_975,In_716,In_577);
or U976 (N_976,In_76,In_332);
and U977 (N_977,In_451,In_353);
and U978 (N_978,In_431,In_605);
nor U979 (N_979,In_50,In_201);
nor U980 (N_980,In_240,In_85);
nand U981 (N_981,In_582,In_97);
and U982 (N_982,In_130,In_749);
nand U983 (N_983,In_216,In_684);
nand U984 (N_984,In_389,In_495);
nand U985 (N_985,In_330,In_177);
or U986 (N_986,In_195,In_744);
and U987 (N_987,In_322,In_703);
nor U988 (N_988,In_696,In_83);
or U989 (N_989,In_712,In_119);
nand U990 (N_990,In_75,In_180);
and U991 (N_991,In_600,In_375);
or U992 (N_992,In_588,In_72);
nor U993 (N_993,In_118,In_491);
nand U994 (N_994,In_40,In_294);
or U995 (N_995,In_588,In_17);
or U996 (N_996,In_38,In_45);
and U997 (N_997,In_158,In_60);
and U998 (N_998,In_160,In_339);
nor U999 (N_999,In_483,In_363);
or U1000 (N_1000,In_528,In_537);
xor U1001 (N_1001,In_405,In_589);
nor U1002 (N_1002,In_252,In_401);
nand U1003 (N_1003,In_416,In_677);
nor U1004 (N_1004,In_386,In_26);
or U1005 (N_1005,In_1,In_97);
or U1006 (N_1006,In_167,In_441);
nand U1007 (N_1007,In_101,In_697);
nor U1008 (N_1008,In_647,In_614);
nor U1009 (N_1009,In_337,In_192);
nor U1010 (N_1010,In_448,In_386);
nor U1011 (N_1011,In_482,In_347);
and U1012 (N_1012,In_614,In_638);
and U1013 (N_1013,In_588,In_256);
nand U1014 (N_1014,In_523,In_569);
nor U1015 (N_1015,In_340,In_470);
nand U1016 (N_1016,In_271,In_346);
nand U1017 (N_1017,In_439,In_564);
and U1018 (N_1018,In_235,In_357);
or U1019 (N_1019,In_356,In_640);
or U1020 (N_1020,In_141,In_405);
or U1021 (N_1021,In_560,In_145);
and U1022 (N_1022,In_212,In_484);
nand U1023 (N_1023,In_463,In_231);
nor U1024 (N_1024,In_538,In_390);
nor U1025 (N_1025,In_151,In_161);
nor U1026 (N_1026,In_385,In_195);
nand U1027 (N_1027,In_744,In_477);
or U1028 (N_1028,In_623,In_408);
and U1029 (N_1029,In_455,In_157);
nand U1030 (N_1030,In_497,In_283);
nor U1031 (N_1031,In_161,In_204);
or U1032 (N_1032,In_481,In_18);
or U1033 (N_1033,In_14,In_736);
nor U1034 (N_1034,In_725,In_221);
nor U1035 (N_1035,In_79,In_472);
and U1036 (N_1036,In_502,In_611);
nor U1037 (N_1037,In_743,In_360);
or U1038 (N_1038,In_499,In_475);
or U1039 (N_1039,In_104,In_175);
nor U1040 (N_1040,In_14,In_634);
nand U1041 (N_1041,In_744,In_80);
or U1042 (N_1042,In_587,In_391);
or U1043 (N_1043,In_583,In_200);
or U1044 (N_1044,In_238,In_624);
or U1045 (N_1045,In_550,In_270);
and U1046 (N_1046,In_420,In_562);
and U1047 (N_1047,In_591,In_728);
nor U1048 (N_1048,In_689,In_88);
nor U1049 (N_1049,In_747,In_194);
and U1050 (N_1050,In_387,In_425);
and U1051 (N_1051,In_119,In_244);
or U1052 (N_1052,In_127,In_167);
nor U1053 (N_1053,In_513,In_78);
nand U1054 (N_1054,In_715,In_403);
or U1055 (N_1055,In_353,In_488);
or U1056 (N_1056,In_596,In_364);
nand U1057 (N_1057,In_156,In_710);
nor U1058 (N_1058,In_500,In_351);
nor U1059 (N_1059,In_101,In_112);
or U1060 (N_1060,In_369,In_140);
nor U1061 (N_1061,In_380,In_172);
nand U1062 (N_1062,In_16,In_536);
and U1063 (N_1063,In_505,In_26);
and U1064 (N_1064,In_91,In_413);
nor U1065 (N_1065,In_159,In_27);
and U1066 (N_1066,In_424,In_612);
and U1067 (N_1067,In_25,In_630);
nor U1068 (N_1068,In_189,In_107);
nor U1069 (N_1069,In_636,In_371);
nor U1070 (N_1070,In_601,In_106);
and U1071 (N_1071,In_739,In_410);
nor U1072 (N_1072,In_573,In_101);
xnor U1073 (N_1073,In_371,In_134);
nand U1074 (N_1074,In_124,In_625);
nand U1075 (N_1075,In_107,In_315);
and U1076 (N_1076,In_579,In_521);
nor U1077 (N_1077,In_92,In_570);
nand U1078 (N_1078,In_47,In_33);
and U1079 (N_1079,In_168,In_373);
and U1080 (N_1080,In_34,In_575);
or U1081 (N_1081,In_62,In_725);
and U1082 (N_1082,In_679,In_652);
nor U1083 (N_1083,In_688,In_187);
and U1084 (N_1084,In_745,In_190);
and U1085 (N_1085,In_537,In_637);
nand U1086 (N_1086,In_378,In_291);
and U1087 (N_1087,In_162,In_649);
nor U1088 (N_1088,In_101,In_729);
nand U1089 (N_1089,In_266,In_379);
or U1090 (N_1090,In_338,In_144);
nor U1091 (N_1091,In_75,In_357);
and U1092 (N_1092,In_82,In_406);
or U1093 (N_1093,In_102,In_408);
or U1094 (N_1094,In_213,In_399);
and U1095 (N_1095,In_177,In_670);
and U1096 (N_1096,In_556,In_579);
or U1097 (N_1097,In_314,In_137);
and U1098 (N_1098,In_31,In_89);
and U1099 (N_1099,In_263,In_479);
and U1100 (N_1100,In_383,In_299);
or U1101 (N_1101,In_601,In_398);
or U1102 (N_1102,In_545,In_560);
or U1103 (N_1103,In_82,In_222);
nor U1104 (N_1104,In_393,In_622);
and U1105 (N_1105,In_368,In_63);
or U1106 (N_1106,In_409,In_528);
or U1107 (N_1107,In_43,In_174);
or U1108 (N_1108,In_378,In_611);
nor U1109 (N_1109,In_180,In_557);
nor U1110 (N_1110,In_664,In_321);
nor U1111 (N_1111,In_364,In_507);
or U1112 (N_1112,In_418,In_248);
nor U1113 (N_1113,In_706,In_567);
or U1114 (N_1114,In_92,In_507);
nor U1115 (N_1115,In_605,In_24);
and U1116 (N_1116,In_257,In_602);
or U1117 (N_1117,In_108,In_647);
nand U1118 (N_1118,In_689,In_414);
nand U1119 (N_1119,In_153,In_481);
nand U1120 (N_1120,In_458,In_613);
nand U1121 (N_1121,In_727,In_660);
and U1122 (N_1122,In_142,In_54);
nand U1123 (N_1123,In_502,In_646);
or U1124 (N_1124,In_219,In_286);
nor U1125 (N_1125,In_294,In_201);
nor U1126 (N_1126,In_47,In_464);
nor U1127 (N_1127,In_265,In_235);
or U1128 (N_1128,In_155,In_491);
or U1129 (N_1129,In_7,In_368);
or U1130 (N_1130,In_154,In_2);
and U1131 (N_1131,In_162,In_655);
nor U1132 (N_1132,In_308,In_369);
nand U1133 (N_1133,In_711,In_49);
or U1134 (N_1134,In_529,In_326);
nand U1135 (N_1135,In_426,In_494);
nor U1136 (N_1136,In_462,In_222);
nand U1137 (N_1137,In_654,In_228);
and U1138 (N_1138,In_462,In_99);
and U1139 (N_1139,In_293,In_106);
nor U1140 (N_1140,In_636,In_329);
and U1141 (N_1141,In_748,In_144);
and U1142 (N_1142,In_240,In_308);
or U1143 (N_1143,In_239,In_740);
nand U1144 (N_1144,In_386,In_385);
nand U1145 (N_1145,In_209,In_105);
or U1146 (N_1146,In_710,In_373);
and U1147 (N_1147,In_346,In_729);
nor U1148 (N_1148,In_280,In_350);
nor U1149 (N_1149,In_282,In_67);
or U1150 (N_1150,In_181,In_157);
and U1151 (N_1151,In_202,In_443);
nand U1152 (N_1152,In_561,In_134);
nor U1153 (N_1153,In_537,In_576);
or U1154 (N_1154,In_214,In_19);
nor U1155 (N_1155,In_17,In_143);
and U1156 (N_1156,In_581,In_641);
and U1157 (N_1157,In_20,In_187);
nand U1158 (N_1158,In_286,In_213);
nand U1159 (N_1159,In_414,In_315);
nand U1160 (N_1160,In_457,In_104);
or U1161 (N_1161,In_335,In_559);
or U1162 (N_1162,In_512,In_1);
nand U1163 (N_1163,In_455,In_307);
and U1164 (N_1164,In_724,In_190);
nor U1165 (N_1165,In_337,In_449);
nand U1166 (N_1166,In_188,In_679);
nor U1167 (N_1167,In_679,In_633);
nand U1168 (N_1168,In_441,In_643);
or U1169 (N_1169,In_555,In_30);
nand U1170 (N_1170,In_357,In_573);
nor U1171 (N_1171,In_686,In_411);
nor U1172 (N_1172,In_540,In_479);
and U1173 (N_1173,In_302,In_576);
nand U1174 (N_1174,In_310,In_169);
nand U1175 (N_1175,In_677,In_272);
nand U1176 (N_1176,In_704,In_162);
and U1177 (N_1177,In_211,In_347);
or U1178 (N_1178,In_386,In_156);
nor U1179 (N_1179,In_0,In_293);
nand U1180 (N_1180,In_225,In_234);
or U1181 (N_1181,In_219,In_104);
nor U1182 (N_1182,In_5,In_301);
and U1183 (N_1183,In_560,In_271);
nand U1184 (N_1184,In_633,In_322);
or U1185 (N_1185,In_544,In_537);
and U1186 (N_1186,In_324,In_400);
nand U1187 (N_1187,In_165,In_497);
and U1188 (N_1188,In_54,In_626);
and U1189 (N_1189,In_580,In_161);
and U1190 (N_1190,In_586,In_646);
nand U1191 (N_1191,In_552,In_460);
and U1192 (N_1192,In_360,In_383);
or U1193 (N_1193,In_536,In_76);
nor U1194 (N_1194,In_548,In_308);
nor U1195 (N_1195,In_117,In_536);
nor U1196 (N_1196,In_276,In_75);
nand U1197 (N_1197,In_376,In_522);
and U1198 (N_1198,In_203,In_622);
and U1199 (N_1199,In_455,In_87);
nor U1200 (N_1200,In_159,In_145);
nand U1201 (N_1201,In_226,In_22);
or U1202 (N_1202,In_406,In_38);
nor U1203 (N_1203,In_733,In_624);
and U1204 (N_1204,In_342,In_36);
or U1205 (N_1205,In_373,In_207);
and U1206 (N_1206,In_102,In_472);
and U1207 (N_1207,In_671,In_250);
nand U1208 (N_1208,In_601,In_181);
or U1209 (N_1209,In_536,In_113);
or U1210 (N_1210,In_304,In_15);
or U1211 (N_1211,In_497,In_685);
and U1212 (N_1212,In_129,In_373);
or U1213 (N_1213,In_460,In_396);
and U1214 (N_1214,In_97,In_248);
nand U1215 (N_1215,In_318,In_113);
or U1216 (N_1216,In_636,In_23);
nand U1217 (N_1217,In_577,In_368);
xor U1218 (N_1218,In_505,In_224);
nor U1219 (N_1219,In_608,In_601);
nand U1220 (N_1220,In_184,In_358);
and U1221 (N_1221,In_111,In_628);
nand U1222 (N_1222,In_255,In_448);
nor U1223 (N_1223,In_452,In_155);
or U1224 (N_1224,In_375,In_160);
or U1225 (N_1225,In_234,In_319);
or U1226 (N_1226,In_695,In_132);
nor U1227 (N_1227,In_57,In_39);
and U1228 (N_1228,In_722,In_232);
or U1229 (N_1229,In_397,In_306);
or U1230 (N_1230,In_15,In_275);
nand U1231 (N_1231,In_66,In_599);
nand U1232 (N_1232,In_189,In_141);
or U1233 (N_1233,In_88,In_606);
or U1234 (N_1234,In_45,In_632);
and U1235 (N_1235,In_274,In_518);
nor U1236 (N_1236,In_143,In_392);
nand U1237 (N_1237,In_711,In_404);
or U1238 (N_1238,In_558,In_193);
nor U1239 (N_1239,In_604,In_133);
nand U1240 (N_1240,In_708,In_441);
xor U1241 (N_1241,In_326,In_715);
nor U1242 (N_1242,In_159,In_496);
nor U1243 (N_1243,In_564,In_82);
and U1244 (N_1244,In_37,In_613);
or U1245 (N_1245,In_321,In_460);
nor U1246 (N_1246,In_434,In_33);
and U1247 (N_1247,In_702,In_230);
xor U1248 (N_1248,In_716,In_319);
and U1249 (N_1249,In_245,In_633);
nand U1250 (N_1250,In_111,In_196);
or U1251 (N_1251,In_276,In_13);
and U1252 (N_1252,In_702,In_449);
and U1253 (N_1253,In_596,In_524);
nand U1254 (N_1254,In_243,In_303);
and U1255 (N_1255,In_277,In_666);
nand U1256 (N_1256,In_209,In_12);
nor U1257 (N_1257,In_660,In_135);
nor U1258 (N_1258,In_401,In_91);
and U1259 (N_1259,In_116,In_566);
nor U1260 (N_1260,In_404,In_375);
and U1261 (N_1261,In_166,In_711);
nand U1262 (N_1262,In_342,In_658);
or U1263 (N_1263,In_123,In_654);
nor U1264 (N_1264,In_454,In_350);
nand U1265 (N_1265,In_147,In_543);
nand U1266 (N_1266,In_300,In_321);
or U1267 (N_1267,In_156,In_451);
nor U1268 (N_1268,In_380,In_528);
nor U1269 (N_1269,In_646,In_14);
xor U1270 (N_1270,In_503,In_125);
nand U1271 (N_1271,In_230,In_240);
or U1272 (N_1272,In_227,In_608);
or U1273 (N_1273,In_472,In_283);
nor U1274 (N_1274,In_688,In_466);
nor U1275 (N_1275,In_586,In_110);
nor U1276 (N_1276,In_171,In_271);
nor U1277 (N_1277,In_703,In_474);
or U1278 (N_1278,In_141,In_284);
nand U1279 (N_1279,In_276,In_292);
and U1280 (N_1280,In_562,In_641);
nand U1281 (N_1281,In_55,In_143);
nand U1282 (N_1282,In_194,In_227);
and U1283 (N_1283,In_330,In_78);
or U1284 (N_1284,In_530,In_232);
nor U1285 (N_1285,In_664,In_655);
or U1286 (N_1286,In_414,In_552);
or U1287 (N_1287,In_629,In_82);
nand U1288 (N_1288,In_202,In_719);
nand U1289 (N_1289,In_416,In_661);
or U1290 (N_1290,In_499,In_333);
nor U1291 (N_1291,In_126,In_45);
or U1292 (N_1292,In_453,In_447);
nand U1293 (N_1293,In_19,In_293);
and U1294 (N_1294,In_461,In_230);
or U1295 (N_1295,In_198,In_274);
nor U1296 (N_1296,In_199,In_477);
or U1297 (N_1297,In_147,In_87);
or U1298 (N_1298,In_481,In_495);
or U1299 (N_1299,In_69,In_230);
or U1300 (N_1300,In_89,In_21);
or U1301 (N_1301,In_441,In_78);
or U1302 (N_1302,In_625,In_325);
nor U1303 (N_1303,In_627,In_591);
and U1304 (N_1304,In_203,In_141);
nor U1305 (N_1305,In_294,In_444);
or U1306 (N_1306,In_123,In_248);
nand U1307 (N_1307,In_110,In_453);
nand U1308 (N_1308,In_317,In_288);
nor U1309 (N_1309,In_152,In_202);
nand U1310 (N_1310,In_411,In_230);
nor U1311 (N_1311,In_183,In_716);
or U1312 (N_1312,In_169,In_322);
or U1313 (N_1313,In_445,In_347);
or U1314 (N_1314,In_297,In_413);
or U1315 (N_1315,In_607,In_163);
nand U1316 (N_1316,In_411,In_372);
nor U1317 (N_1317,In_334,In_575);
nand U1318 (N_1318,In_560,In_746);
nand U1319 (N_1319,In_419,In_399);
nand U1320 (N_1320,In_317,In_306);
nand U1321 (N_1321,In_268,In_647);
and U1322 (N_1322,In_148,In_697);
nor U1323 (N_1323,In_583,In_183);
and U1324 (N_1324,In_213,In_724);
and U1325 (N_1325,In_527,In_1);
nand U1326 (N_1326,In_697,In_542);
nand U1327 (N_1327,In_27,In_202);
nand U1328 (N_1328,In_728,In_363);
xnor U1329 (N_1329,In_512,In_594);
or U1330 (N_1330,In_80,In_278);
nand U1331 (N_1331,In_734,In_422);
and U1332 (N_1332,In_189,In_428);
nor U1333 (N_1333,In_660,In_156);
nand U1334 (N_1334,In_744,In_578);
nor U1335 (N_1335,In_75,In_285);
or U1336 (N_1336,In_226,In_31);
nor U1337 (N_1337,In_671,In_201);
or U1338 (N_1338,In_194,In_419);
and U1339 (N_1339,In_210,In_22);
and U1340 (N_1340,In_596,In_335);
nand U1341 (N_1341,In_269,In_554);
nor U1342 (N_1342,In_480,In_470);
and U1343 (N_1343,In_380,In_68);
or U1344 (N_1344,In_338,In_406);
nor U1345 (N_1345,In_513,In_19);
nor U1346 (N_1346,In_36,In_641);
or U1347 (N_1347,In_569,In_263);
nand U1348 (N_1348,In_92,In_4);
or U1349 (N_1349,In_400,In_570);
and U1350 (N_1350,In_73,In_159);
and U1351 (N_1351,In_316,In_175);
nor U1352 (N_1352,In_647,In_608);
nand U1353 (N_1353,In_91,In_192);
or U1354 (N_1354,In_45,In_397);
nand U1355 (N_1355,In_517,In_90);
and U1356 (N_1356,In_460,In_500);
xor U1357 (N_1357,In_127,In_427);
or U1358 (N_1358,In_54,In_699);
nand U1359 (N_1359,In_462,In_502);
nand U1360 (N_1360,In_594,In_566);
nor U1361 (N_1361,In_196,In_734);
or U1362 (N_1362,In_733,In_304);
or U1363 (N_1363,In_191,In_527);
and U1364 (N_1364,In_557,In_72);
nand U1365 (N_1365,In_271,In_371);
nand U1366 (N_1366,In_137,In_683);
or U1367 (N_1367,In_41,In_201);
nand U1368 (N_1368,In_672,In_686);
nand U1369 (N_1369,In_530,In_668);
or U1370 (N_1370,In_370,In_586);
or U1371 (N_1371,In_319,In_104);
nor U1372 (N_1372,In_80,In_297);
or U1373 (N_1373,In_412,In_615);
or U1374 (N_1374,In_346,In_204);
nor U1375 (N_1375,In_426,In_329);
and U1376 (N_1376,In_654,In_241);
nor U1377 (N_1377,In_401,In_735);
or U1378 (N_1378,In_602,In_61);
nand U1379 (N_1379,In_704,In_259);
or U1380 (N_1380,In_486,In_337);
xnor U1381 (N_1381,In_747,In_396);
nand U1382 (N_1382,In_559,In_591);
nand U1383 (N_1383,In_205,In_316);
and U1384 (N_1384,In_50,In_19);
nand U1385 (N_1385,In_639,In_52);
and U1386 (N_1386,In_656,In_355);
or U1387 (N_1387,In_621,In_88);
nand U1388 (N_1388,In_394,In_183);
and U1389 (N_1389,In_422,In_343);
nand U1390 (N_1390,In_497,In_80);
nand U1391 (N_1391,In_234,In_743);
and U1392 (N_1392,In_414,In_135);
and U1393 (N_1393,In_188,In_212);
and U1394 (N_1394,In_340,In_369);
nor U1395 (N_1395,In_335,In_550);
or U1396 (N_1396,In_379,In_298);
nand U1397 (N_1397,In_88,In_708);
nand U1398 (N_1398,In_357,In_739);
nand U1399 (N_1399,In_705,In_735);
or U1400 (N_1400,In_39,In_24);
or U1401 (N_1401,In_200,In_61);
nand U1402 (N_1402,In_730,In_312);
or U1403 (N_1403,In_708,In_96);
and U1404 (N_1404,In_651,In_632);
or U1405 (N_1405,In_382,In_611);
and U1406 (N_1406,In_138,In_231);
nor U1407 (N_1407,In_749,In_519);
and U1408 (N_1408,In_690,In_97);
and U1409 (N_1409,In_429,In_530);
or U1410 (N_1410,In_622,In_667);
or U1411 (N_1411,In_71,In_715);
nand U1412 (N_1412,In_460,In_296);
nor U1413 (N_1413,In_631,In_691);
nand U1414 (N_1414,In_126,In_124);
nor U1415 (N_1415,In_199,In_707);
or U1416 (N_1416,In_372,In_230);
nand U1417 (N_1417,In_551,In_501);
or U1418 (N_1418,In_100,In_547);
and U1419 (N_1419,In_565,In_473);
nand U1420 (N_1420,In_197,In_426);
or U1421 (N_1421,In_196,In_310);
nand U1422 (N_1422,In_642,In_664);
or U1423 (N_1423,In_101,In_111);
nand U1424 (N_1424,In_87,In_16);
or U1425 (N_1425,In_498,In_378);
nand U1426 (N_1426,In_405,In_104);
xnor U1427 (N_1427,In_728,In_346);
nand U1428 (N_1428,In_299,In_25);
nor U1429 (N_1429,In_710,In_590);
or U1430 (N_1430,In_534,In_35);
and U1431 (N_1431,In_732,In_54);
nand U1432 (N_1432,In_524,In_552);
or U1433 (N_1433,In_356,In_416);
nor U1434 (N_1434,In_257,In_443);
nand U1435 (N_1435,In_684,In_636);
nand U1436 (N_1436,In_209,In_339);
or U1437 (N_1437,In_464,In_717);
and U1438 (N_1438,In_491,In_715);
nand U1439 (N_1439,In_225,In_63);
and U1440 (N_1440,In_249,In_185);
xor U1441 (N_1441,In_642,In_93);
nand U1442 (N_1442,In_121,In_461);
nor U1443 (N_1443,In_430,In_27);
nand U1444 (N_1444,In_457,In_380);
nor U1445 (N_1445,In_279,In_405);
and U1446 (N_1446,In_581,In_654);
or U1447 (N_1447,In_673,In_508);
nor U1448 (N_1448,In_126,In_492);
and U1449 (N_1449,In_417,In_529);
or U1450 (N_1450,In_91,In_158);
nand U1451 (N_1451,In_105,In_95);
nor U1452 (N_1452,In_103,In_508);
and U1453 (N_1453,In_288,In_239);
nand U1454 (N_1454,In_329,In_343);
nor U1455 (N_1455,In_283,In_178);
nand U1456 (N_1456,In_657,In_59);
or U1457 (N_1457,In_352,In_118);
nand U1458 (N_1458,In_99,In_514);
nand U1459 (N_1459,In_228,In_127);
and U1460 (N_1460,In_384,In_360);
xnor U1461 (N_1461,In_489,In_84);
and U1462 (N_1462,In_349,In_518);
xnor U1463 (N_1463,In_595,In_357);
and U1464 (N_1464,In_479,In_329);
nand U1465 (N_1465,In_567,In_527);
nor U1466 (N_1466,In_120,In_422);
nand U1467 (N_1467,In_239,In_132);
and U1468 (N_1468,In_112,In_670);
nor U1469 (N_1469,In_692,In_10);
and U1470 (N_1470,In_370,In_712);
nor U1471 (N_1471,In_583,In_545);
nor U1472 (N_1472,In_315,In_394);
and U1473 (N_1473,In_339,In_606);
or U1474 (N_1474,In_248,In_537);
or U1475 (N_1475,In_446,In_54);
nor U1476 (N_1476,In_404,In_368);
and U1477 (N_1477,In_283,In_591);
nand U1478 (N_1478,In_135,In_208);
nor U1479 (N_1479,In_171,In_245);
and U1480 (N_1480,In_743,In_526);
and U1481 (N_1481,In_585,In_367);
or U1482 (N_1482,In_448,In_682);
and U1483 (N_1483,In_253,In_469);
nand U1484 (N_1484,In_740,In_256);
and U1485 (N_1485,In_735,In_395);
nand U1486 (N_1486,In_379,In_32);
nor U1487 (N_1487,In_542,In_222);
nand U1488 (N_1488,In_42,In_126);
nor U1489 (N_1489,In_18,In_650);
nand U1490 (N_1490,In_308,In_646);
and U1491 (N_1491,In_273,In_617);
nor U1492 (N_1492,In_27,In_466);
or U1493 (N_1493,In_67,In_524);
and U1494 (N_1494,In_565,In_172);
and U1495 (N_1495,In_73,In_226);
nor U1496 (N_1496,In_38,In_181);
nor U1497 (N_1497,In_647,In_159);
and U1498 (N_1498,In_493,In_736);
nand U1499 (N_1499,In_522,In_331);
nor U1500 (N_1500,In_52,In_422);
nand U1501 (N_1501,In_685,In_202);
and U1502 (N_1502,In_676,In_341);
nand U1503 (N_1503,In_18,In_240);
or U1504 (N_1504,In_712,In_217);
or U1505 (N_1505,In_55,In_100);
nor U1506 (N_1506,In_264,In_198);
nand U1507 (N_1507,In_548,In_292);
and U1508 (N_1508,In_469,In_622);
and U1509 (N_1509,In_727,In_699);
nor U1510 (N_1510,In_342,In_161);
and U1511 (N_1511,In_308,In_482);
and U1512 (N_1512,In_538,In_189);
nand U1513 (N_1513,In_28,In_230);
or U1514 (N_1514,In_515,In_262);
and U1515 (N_1515,In_272,In_311);
or U1516 (N_1516,In_687,In_6);
nand U1517 (N_1517,In_456,In_651);
and U1518 (N_1518,In_447,In_115);
nor U1519 (N_1519,In_363,In_134);
nor U1520 (N_1520,In_389,In_190);
and U1521 (N_1521,In_245,In_575);
and U1522 (N_1522,In_185,In_214);
nor U1523 (N_1523,In_39,In_485);
nand U1524 (N_1524,In_251,In_312);
or U1525 (N_1525,In_438,In_231);
nor U1526 (N_1526,In_518,In_50);
or U1527 (N_1527,In_461,In_539);
or U1528 (N_1528,In_538,In_724);
or U1529 (N_1529,In_180,In_566);
or U1530 (N_1530,In_583,In_409);
nor U1531 (N_1531,In_419,In_628);
and U1532 (N_1532,In_7,In_172);
nand U1533 (N_1533,In_31,In_52);
nand U1534 (N_1534,In_634,In_38);
and U1535 (N_1535,In_294,In_28);
or U1536 (N_1536,In_666,In_715);
nand U1537 (N_1537,In_464,In_152);
nand U1538 (N_1538,In_584,In_732);
nor U1539 (N_1539,In_88,In_628);
and U1540 (N_1540,In_707,In_675);
xor U1541 (N_1541,In_121,In_59);
and U1542 (N_1542,In_218,In_467);
or U1543 (N_1543,In_1,In_566);
nand U1544 (N_1544,In_600,In_455);
and U1545 (N_1545,In_618,In_167);
or U1546 (N_1546,In_26,In_221);
nor U1547 (N_1547,In_709,In_460);
and U1548 (N_1548,In_364,In_653);
nor U1549 (N_1549,In_653,In_300);
and U1550 (N_1550,In_521,In_425);
and U1551 (N_1551,In_377,In_384);
nand U1552 (N_1552,In_403,In_290);
nand U1553 (N_1553,In_556,In_198);
or U1554 (N_1554,In_29,In_418);
or U1555 (N_1555,In_300,In_9);
and U1556 (N_1556,In_298,In_638);
nor U1557 (N_1557,In_127,In_714);
or U1558 (N_1558,In_492,In_481);
and U1559 (N_1559,In_642,In_561);
nand U1560 (N_1560,In_16,In_665);
nor U1561 (N_1561,In_65,In_560);
nor U1562 (N_1562,In_456,In_414);
nor U1563 (N_1563,In_719,In_433);
and U1564 (N_1564,In_172,In_629);
nor U1565 (N_1565,In_530,In_159);
xor U1566 (N_1566,In_262,In_233);
nand U1567 (N_1567,In_155,In_582);
or U1568 (N_1568,In_280,In_329);
nand U1569 (N_1569,In_356,In_512);
and U1570 (N_1570,In_357,In_719);
nor U1571 (N_1571,In_350,In_347);
and U1572 (N_1572,In_304,In_738);
nand U1573 (N_1573,In_324,In_14);
nor U1574 (N_1574,In_341,In_706);
nand U1575 (N_1575,In_317,In_282);
xnor U1576 (N_1576,In_412,In_492);
nor U1577 (N_1577,In_741,In_215);
nand U1578 (N_1578,In_451,In_409);
nand U1579 (N_1579,In_545,In_260);
and U1580 (N_1580,In_463,In_100);
or U1581 (N_1581,In_728,In_658);
nor U1582 (N_1582,In_326,In_418);
nand U1583 (N_1583,In_240,In_362);
and U1584 (N_1584,In_132,In_166);
nor U1585 (N_1585,In_349,In_494);
and U1586 (N_1586,In_567,In_171);
nor U1587 (N_1587,In_700,In_747);
nor U1588 (N_1588,In_620,In_183);
or U1589 (N_1589,In_339,In_276);
and U1590 (N_1590,In_218,In_549);
or U1591 (N_1591,In_67,In_61);
and U1592 (N_1592,In_490,In_504);
or U1593 (N_1593,In_61,In_91);
xor U1594 (N_1594,In_567,In_545);
nand U1595 (N_1595,In_190,In_155);
nor U1596 (N_1596,In_741,In_168);
nor U1597 (N_1597,In_475,In_213);
and U1598 (N_1598,In_30,In_537);
nand U1599 (N_1599,In_395,In_425);
or U1600 (N_1600,In_634,In_2);
nor U1601 (N_1601,In_5,In_77);
xor U1602 (N_1602,In_228,In_198);
and U1603 (N_1603,In_354,In_596);
nor U1604 (N_1604,In_364,In_565);
nor U1605 (N_1605,In_400,In_662);
nand U1606 (N_1606,In_418,In_291);
xor U1607 (N_1607,In_621,In_497);
or U1608 (N_1608,In_305,In_646);
nor U1609 (N_1609,In_381,In_322);
or U1610 (N_1610,In_708,In_115);
and U1611 (N_1611,In_716,In_707);
and U1612 (N_1612,In_86,In_110);
or U1613 (N_1613,In_431,In_182);
and U1614 (N_1614,In_650,In_692);
nand U1615 (N_1615,In_405,In_749);
or U1616 (N_1616,In_249,In_645);
nand U1617 (N_1617,In_460,In_189);
nand U1618 (N_1618,In_265,In_645);
xnor U1619 (N_1619,In_26,In_281);
nor U1620 (N_1620,In_568,In_725);
or U1621 (N_1621,In_618,In_162);
or U1622 (N_1622,In_676,In_710);
nand U1623 (N_1623,In_255,In_653);
nand U1624 (N_1624,In_654,In_131);
or U1625 (N_1625,In_60,In_625);
or U1626 (N_1626,In_308,In_713);
nor U1627 (N_1627,In_572,In_391);
and U1628 (N_1628,In_700,In_491);
or U1629 (N_1629,In_704,In_673);
and U1630 (N_1630,In_522,In_23);
and U1631 (N_1631,In_344,In_568);
nand U1632 (N_1632,In_370,In_255);
nand U1633 (N_1633,In_277,In_380);
or U1634 (N_1634,In_557,In_326);
nand U1635 (N_1635,In_244,In_61);
or U1636 (N_1636,In_41,In_310);
nand U1637 (N_1637,In_675,In_536);
and U1638 (N_1638,In_22,In_83);
or U1639 (N_1639,In_154,In_457);
and U1640 (N_1640,In_306,In_236);
xnor U1641 (N_1641,In_107,In_745);
nand U1642 (N_1642,In_144,In_528);
nor U1643 (N_1643,In_573,In_597);
and U1644 (N_1644,In_504,In_577);
nand U1645 (N_1645,In_568,In_528);
nor U1646 (N_1646,In_195,In_651);
or U1647 (N_1647,In_345,In_550);
and U1648 (N_1648,In_561,In_344);
nor U1649 (N_1649,In_73,In_425);
or U1650 (N_1650,In_188,In_309);
nor U1651 (N_1651,In_214,In_525);
or U1652 (N_1652,In_0,In_119);
and U1653 (N_1653,In_107,In_178);
or U1654 (N_1654,In_326,In_347);
or U1655 (N_1655,In_610,In_397);
or U1656 (N_1656,In_111,In_383);
nor U1657 (N_1657,In_410,In_4);
and U1658 (N_1658,In_388,In_579);
and U1659 (N_1659,In_221,In_404);
nor U1660 (N_1660,In_175,In_656);
and U1661 (N_1661,In_197,In_63);
or U1662 (N_1662,In_178,In_292);
nand U1663 (N_1663,In_413,In_22);
and U1664 (N_1664,In_306,In_41);
nand U1665 (N_1665,In_681,In_460);
or U1666 (N_1666,In_46,In_222);
nor U1667 (N_1667,In_364,In_738);
nand U1668 (N_1668,In_403,In_409);
or U1669 (N_1669,In_58,In_478);
nor U1670 (N_1670,In_589,In_221);
nor U1671 (N_1671,In_655,In_11);
or U1672 (N_1672,In_186,In_467);
xor U1673 (N_1673,In_352,In_170);
nand U1674 (N_1674,In_303,In_716);
nor U1675 (N_1675,In_220,In_495);
nand U1676 (N_1676,In_377,In_25);
and U1677 (N_1677,In_667,In_534);
and U1678 (N_1678,In_153,In_485);
and U1679 (N_1679,In_210,In_163);
or U1680 (N_1680,In_393,In_566);
and U1681 (N_1681,In_697,In_86);
nor U1682 (N_1682,In_149,In_407);
and U1683 (N_1683,In_609,In_462);
or U1684 (N_1684,In_369,In_631);
or U1685 (N_1685,In_78,In_426);
and U1686 (N_1686,In_607,In_137);
nand U1687 (N_1687,In_218,In_692);
and U1688 (N_1688,In_395,In_640);
nand U1689 (N_1689,In_59,In_139);
and U1690 (N_1690,In_615,In_606);
and U1691 (N_1691,In_114,In_190);
nor U1692 (N_1692,In_329,In_319);
or U1693 (N_1693,In_368,In_623);
nor U1694 (N_1694,In_489,In_263);
nor U1695 (N_1695,In_415,In_387);
nand U1696 (N_1696,In_470,In_678);
nor U1697 (N_1697,In_152,In_18);
nor U1698 (N_1698,In_140,In_22);
nor U1699 (N_1699,In_124,In_180);
and U1700 (N_1700,In_266,In_336);
nand U1701 (N_1701,In_276,In_576);
nand U1702 (N_1702,In_322,In_682);
nand U1703 (N_1703,In_326,In_502);
and U1704 (N_1704,In_263,In_300);
or U1705 (N_1705,In_648,In_323);
nor U1706 (N_1706,In_255,In_550);
nand U1707 (N_1707,In_726,In_578);
or U1708 (N_1708,In_573,In_340);
nor U1709 (N_1709,In_174,In_183);
nand U1710 (N_1710,In_520,In_278);
nor U1711 (N_1711,In_466,In_673);
or U1712 (N_1712,In_99,In_72);
nor U1713 (N_1713,In_600,In_404);
or U1714 (N_1714,In_168,In_526);
or U1715 (N_1715,In_352,In_537);
or U1716 (N_1716,In_200,In_406);
nor U1717 (N_1717,In_494,In_383);
and U1718 (N_1718,In_707,In_744);
nor U1719 (N_1719,In_555,In_685);
xor U1720 (N_1720,In_130,In_671);
xor U1721 (N_1721,In_670,In_373);
nand U1722 (N_1722,In_112,In_476);
or U1723 (N_1723,In_269,In_578);
nand U1724 (N_1724,In_302,In_607);
or U1725 (N_1725,In_363,In_654);
or U1726 (N_1726,In_432,In_667);
nor U1727 (N_1727,In_333,In_161);
nor U1728 (N_1728,In_700,In_560);
nor U1729 (N_1729,In_663,In_39);
nor U1730 (N_1730,In_426,In_195);
and U1731 (N_1731,In_688,In_146);
or U1732 (N_1732,In_358,In_200);
nand U1733 (N_1733,In_538,In_46);
or U1734 (N_1734,In_417,In_626);
xor U1735 (N_1735,In_612,In_256);
nand U1736 (N_1736,In_324,In_4);
nand U1737 (N_1737,In_89,In_1);
nand U1738 (N_1738,In_118,In_223);
or U1739 (N_1739,In_323,In_189);
nor U1740 (N_1740,In_191,In_194);
nor U1741 (N_1741,In_534,In_745);
nand U1742 (N_1742,In_521,In_624);
or U1743 (N_1743,In_585,In_474);
nor U1744 (N_1744,In_637,In_657);
xor U1745 (N_1745,In_518,In_738);
nor U1746 (N_1746,In_643,In_115);
nor U1747 (N_1747,In_60,In_362);
nor U1748 (N_1748,In_41,In_735);
nor U1749 (N_1749,In_168,In_227);
and U1750 (N_1750,In_377,In_536);
or U1751 (N_1751,In_488,In_103);
or U1752 (N_1752,In_60,In_736);
nand U1753 (N_1753,In_431,In_477);
nand U1754 (N_1754,In_583,In_31);
and U1755 (N_1755,In_613,In_644);
nand U1756 (N_1756,In_38,In_4);
and U1757 (N_1757,In_93,In_351);
nor U1758 (N_1758,In_706,In_365);
or U1759 (N_1759,In_106,In_423);
nand U1760 (N_1760,In_264,In_444);
or U1761 (N_1761,In_111,In_619);
or U1762 (N_1762,In_487,In_628);
nor U1763 (N_1763,In_662,In_477);
nor U1764 (N_1764,In_298,In_531);
or U1765 (N_1765,In_472,In_588);
or U1766 (N_1766,In_675,In_503);
nor U1767 (N_1767,In_408,In_641);
or U1768 (N_1768,In_594,In_323);
xor U1769 (N_1769,In_381,In_633);
and U1770 (N_1770,In_563,In_138);
and U1771 (N_1771,In_283,In_33);
nor U1772 (N_1772,In_468,In_12);
or U1773 (N_1773,In_313,In_271);
and U1774 (N_1774,In_640,In_39);
and U1775 (N_1775,In_157,In_27);
nand U1776 (N_1776,In_594,In_448);
nand U1777 (N_1777,In_327,In_58);
nor U1778 (N_1778,In_706,In_629);
or U1779 (N_1779,In_679,In_338);
nand U1780 (N_1780,In_13,In_71);
nor U1781 (N_1781,In_408,In_130);
or U1782 (N_1782,In_32,In_725);
nand U1783 (N_1783,In_39,In_106);
or U1784 (N_1784,In_633,In_275);
nor U1785 (N_1785,In_742,In_288);
and U1786 (N_1786,In_659,In_622);
nand U1787 (N_1787,In_621,In_558);
nor U1788 (N_1788,In_390,In_73);
or U1789 (N_1789,In_687,In_163);
nand U1790 (N_1790,In_350,In_284);
nand U1791 (N_1791,In_7,In_142);
nor U1792 (N_1792,In_678,In_392);
nor U1793 (N_1793,In_194,In_399);
nor U1794 (N_1794,In_585,In_710);
and U1795 (N_1795,In_335,In_222);
and U1796 (N_1796,In_133,In_637);
nand U1797 (N_1797,In_540,In_47);
nor U1798 (N_1798,In_231,In_104);
nor U1799 (N_1799,In_601,In_193);
nand U1800 (N_1800,In_425,In_600);
or U1801 (N_1801,In_316,In_231);
xor U1802 (N_1802,In_302,In_145);
or U1803 (N_1803,In_592,In_316);
and U1804 (N_1804,In_459,In_639);
and U1805 (N_1805,In_531,In_411);
nor U1806 (N_1806,In_159,In_67);
and U1807 (N_1807,In_152,In_253);
or U1808 (N_1808,In_589,In_539);
nand U1809 (N_1809,In_220,In_492);
or U1810 (N_1810,In_584,In_467);
or U1811 (N_1811,In_555,In_90);
and U1812 (N_1812,In_104,In_96);
or U1813 (N_1813,In_547,In_314);
nor U1814 (N_1814,In_271,In_27);
nand U1815 (N_1815,In_742,In_167);
nand U1816 (N_1816,In_330,In_531);
nor U1817 (N_1817,In_425,In_292);
or U1818 (N_1818,In_466,In_453);
nor U1819 (N_1819,In_30,In_371);
or U1820 (N_1820,In_562,In_251);
nand U1821 (N_1821,In_612,In_2);
nand U1822 (N_1822,In_454,In_328);
nand U1823 (N_1823,In_739,In_434);
nand U1824 (N_1824,In_525,In_391);
nand U1825 (N_1825,In_529,In_125);
or U1826 (N_1826,In_110,In_344);
nor U1827 (N_1827,In_426,In_13);
and U1828 (N_1828,In_15,In_181);
and U1829 (N_1829,In_589,In_676);
or U1830 (N_1830,In_711,In_77);
nand U1831 (N_1831,In_222,In_95);
nand U1832 (N_1832,In_209,In_420);
nand U1833 (N_1833,In_626,In_612);
or U1834 (N_1834,In_254,In_530);
nand U1835 (N_1835,In_222,In_635);
or U1836 (N_1836,In_288,In_177);
or U1837 (N_1837,In_357,In_188);
and U1838 (N_1838,In_162,In_342);
or U1839 (N_1839,In_253,In_296);
and U1840 (N_1840,In_736,In_89);
nor U1841 (N_1841,In_226,In_131);
and U1842 (N_1842,In_53,In_169);
nand U1843 (N_1843,In_332,In_150);
or U1844 (N_1844,In_278,In_64);
nor U1845 (N_1845,In_215,In_86);
and U1846 (N_1846,In_587,In_732);
nand U1847 (N_1847,In_440,In_262);
nor U1848 (N_1848,In_417,In_150);
or U1849 (N_1849,In_167,In_747);
nor U1850 (N_1850,In_250,In_586);
and U1851 (N_1851,In_720,In_476);
nand U1852 (N_1852,In_262,In_279);
nand U1853 (N_1853,In_749,In_354);
xnor U1854 (N_1854,In_597,In_530);
nor U1855 (N_1855,In_283,In_628);
nand U1856 (N_1856,In_4,In_203);
nand U1857 (N_1857,In_368,In_435);
and U1858 (N_1858,In_483,In_154);
nand U1859 (N_1859,In_744,In_496);
nor U1860 (N_1860,In_688,In_210);
or U1861 (N_1861,In_517,In_717);
nor U1862 (N_1862,In_305,In_738);
nor U1863 (N_1863,In_1,In_575);
and U1864 (N_1864,In_178,In_488);
nand U1865 (N_1865,In_718,In_613);
nand U1866 (N_1866,In_569,In_346);
or U1867 (N_1867,In_210,In_426);
and U1868 (N_1868,In_434,In_100);
nor U1869 (N_1869,In_552,In_713);
or U1870 (N_1870,In_693,In_203);
nor U1871 (N_1871,In_155,In_676);
and U1872 (N_1872,In_730,In_406);
or U1873 (N_1873,In_222,In_576);
nand U1874 (N_1874,In_264,In_250);
or U1875 (N_1875,In_265,In_629);
and U1876 (N_1876,In_533,In_306);
and U1877 (N_1877,In_387,In_7);
nor U1878 (N_1878,In_460,In_297);
nor U1879 (N_1879,In_178,In_310);
nand U1880 (N_1880,In_255,In_623);
and U1881 (N_1881,In_665,In_730);
nand U1882 (N_1882,In_545,In_182);
and U1883 (N_1883,In_10,In_490);
or U1884 (N_1884,In_697,In_550);
and U1885 (N_1885,In_737,In_254);
nand U1886 (N_1886,In_79,In_421);
nor U1887 (N_1887,In_42,In_672);
or U1888 (N_1888,In_131,In_722);
or U1889 (N_1889,In_589,In_12);
and U1890 (N_1890,In_138,In_698);
or U1891 (N_1891,In_205,In_400);
nand U1892 (N_1892,In_485,In_269);
or U1893 (N_1893,In_680,In_490);
or U1894 (N_1894,In_96,In_106);
or U1895 (N_1895,In_328,In_457);
nor U1896 (N_1896,In_326,In_503);
and U1897 (N_1897,In_747,In_339);
nand U1898 (N_1898,In_45,In_376);
and U1899 (N_1899,In_201,In_278);
nor U1900 (N_1900,In_418,In_568);
and U1901 (N_1901,In_358,In_352);
nand U1902 (N_1902,In_20,In_189);
or U1903 (N_1903,In_717,In_527);
and U1904 (N_1904,In_300,In_435);
or U1905 (N_1905,In_532,In_604);
or U1906 (N_1906,In_710,In_569);
nand U1907 (N_1907,In_481,In_257);
and U1908 (N_1908,In_405,In_285);
or U1909 (N_1909,In_366,In_478);
nor U1910 (N_1910,In_288,In_552);
nand U1911 (N_1911,In_358,In_744);
or U1912 (N_1912,In_388,In_266);
nor U1913 (N_1913,In_130,In_198);
and U1914 (N_1914,In_468,In_640);
and U1915 (N_1915,In_497,In_147);
and U1916 (N_1916,In_667,In_520);
nor U1917 (N_1917,In_502,In_552);
or U1918 (N_1918,In_506,In_679);
or U1919 (N_1919,In_461,In_502);
or U1920 (N_1920,In_168,In_258);
or U1921 (N_1921,In_98,In_341);
nand U1922 (N_1922,In_728,In_492);
or U1923 (N_1923,In_707,In_492);
and U1924 (N_1924,In_35,In_728);
and U1925 (N_1925,In_75,In_130);
nor U1926 (N_1926,In_664,In_110);
nor U1927 (N_1927,In_227,In_553);
or U1928 (N_1928,In_354,In_694);
or U1929 (N_1929,In_163,In_711);
and U1930 (N_1930,In_348,In_218);
nand U1931 (N_1931,In_521,In_546);
nand U1932 (N_1932,In_419,In_232);
or U1933 (N_1933,In_703,In_227);
nand U1934 (N_1934,In_30,In_126);
or U1935 (N_1935,In_180,In_171);
or U1936 (N_1936,In_223,In_619);
or U1937 (N_1937,In_492,In_159);
and U1938 (N_1938,In_733,In_1);
nor U1939 (N_1939,In_490,In_377);
or U1940 (N_1940,In_463,In_53);
nor U1941 (N_1941,In_350,In_532);
or U1942 (N_1942,In_509,In_722);
nand U1943 (N_1943,In_585,In_283);
nor U1944 (N_1944,In_364,In_505);
or U1945 (N_1945,In_178,In_26);
and U1946 (N_1946,In_280,In_335);
nand U1947 (N_1947,In_126,In_235);
nor U1948 (N_1948,In_600,In_158);
and U1949 (N_1949,In_345,In_262);
or U1950 (N_1950,In_426,In_622);
and U1951 (N_1951,In_84,In_582);
nand U1952 (N_1952,In_55,In_401);
and U1953 (N_1953,In_58,In_553);
and U1954 (N_1954,In_34,In_400);
nand U1955 (N_1955,In_280,In_716);
nand U1956 (N_1956,In_278,In_664);
xor U1957 (N_1957,In_332,In_676);
and U1958 (N_1958,In_552,In_344);
and U1959 (N_1959,In_629,In_371);
nor U1960 (N_1960,In_184,In_351);
nand U1961 (N_1961,In_626,In_517);
and U1962 (N_1962,In_473,In_0);
or U1963 (N_1963,In_25,In_67);
nand U1964 (N_1964,In_276,In_644);
or U1965 (N_1965,In_117,In_567);
or U1966 (N_1966,In_665,In_603);
or U1967 (N_1967,In_337,In_521);
and U1968 (N_1968,In_211,In_741);
nand U1969 (N_1969,In_449,In_142);
nand U1970 (N_1970,In_243,In_227);
nor U1971 (N_1971,In_509,In_711);
nand U1972 (N_1972,In_273,In_422);
nand U1973 (N_1973,In_470,In_738);
nand U1974 (N_1974,In_283,In_736);
and U1975 (N_1975,In_611,In_540);
or U1976 (N_1976,In_216,In_336);
and U1977 (N_1977,In_576,In_565);
or U1978 (N_1978,In_730,In_538);
nor U1979 (N_1979,In_39,In_123);
nor U1980 (N_1980,In_77,In_289);
nor U1981 (N_1981,In_577,In_328);
nand U1982 (N_1982,In_145,In_308);
nor U1983 (N_1983,In_301,In_138);
nand U1984 (N_1984,In_440,In_631);
nor U1985 (N_1985,In_161,In_387);
nor U1986 (N_1986,In_571,In_526);
or U1987 (N_1987,In_181,In_652);
and U1988 (N_1988,In_60,In_449);
nor U1989 (N_1989,In_465,In_569);
and U1990 (N_1990,In_560,In_749);
and U1991 (N_1991,In_217,In_302);
or U1992 (N_1992,In_120,In_703);
and U1993 (N_1993,In_409,In_587);
nand U1994 (N_1994,In_150,In_0);
or U1995 (N_1995,In_498,In_627);
nor U1996 (N_1996,In_575,In_735);
nor U1997 (N_1997,In_729,In_748);
nand U1998 (N_1998,In_228,In_107);
and U1999 (N_1999,In_91,In_20);
or U2000 (N_2000,In_503,In_148);
nand U2001 (N_2001,In_710,In_129);
nor U2002 (N_2002,In_148,In_207);
nor U2003 (N_2003,In_134,In_218);
nand U2004 (N_2004,In_489,In_456);
nor U2005 (N_2005,In_282,In_469);
xnor U2006 (N_2006,In_272,In_588);
nor U2007 (N_2007,In_478,In_658);
and U2008 (N_2008,In_280,In_714);
and U2009 (N_2009,In_565,In_501);
or U2010 (N_2010,In_501,In_625);
nand U2011 (N_2011,In_346,In_619);
and U2012 (N_2012,In_636,In_82);
or U2013 (N_2013,In_1,In_369);
or U2014 (N_2014,In_90,In_22);
nand U2015 (N_2015,In_294,In_195);
nor U2016 (N_2016,In_122,In_481);
and U2017 (N_2017,In_156,In_458);
nor U2018 (N_2018,In_463,In_396);
nand U2019 (N_2019,In_350,In_636);
nor U2020 (N_2020,In_620,In_310);
nor U2021 (N_2021,In_565,In_267);
or U2022 (N_2022,In_671,In_343);
nor U2023 (N_2023,In_371,In_742);
xnor U2024 (N_2024,In_449,In_74);
nand U2025 (N_2025,In_350,In_406);
and U2026 (N_2026,In_556,In_696);
and U2027 (N_2027,In_353,In_408);
nand U2028 (N_2028,In_92,In_666);
and U2029 (N_2029,In_158,In_547);
xor U2030 (N_2030,In_441,In_283);
nor U2031 (N_2031,In_556,In_131);
nor U2032 (N_2032,In_566,In_71);
nand U2033 (N_2033,In_18,In_541);
nand U2034 (N_2034,In_63,In_373);
nor U2035 (N_2035,In_493,In_63);
or U2036 (N_2036,In_188,In_560);
nand U2037 (N_2037,In_137,In_544);
nand U2038 (N_2038,In_594,In_445);
nand U2039 (N_2039,In_313,In_507);
and U2040 (N_2040,In_259,In_427);
nor U2041 (N_2041,In_643,In_322);
nand U2042 (N_2042,In_396,In_254);
nor U2043 (N_2043,In_277,In_251);
nor U2044 (N_2044,In_440,In_26);
and U2045 (N_2045,In_379,In_735);
or U2046 (N_2046,In_629,In_551);
or U2047 (N_2047,In_291,In_217);
nor U2048 (N_2048,In_179,In_53);
nor U2049 (N_2049,In_527,In_128);
and U2050 (N_2050,In_374,In_257);
and U2051 (N_2051,In_267,In_362);
nand U2052 (N_2052,In_248,In_435);
nand U2053 (N_2053,In_137,In_288);
and U2054 (N_2054,In_413,In_365);
nor U2055 (N_2055,In_454,In_440);
or U2056 (N_2056,In_657,In_555);
nor U2057 (N_2057,In_516,In_24);
and U2058 (N_2058,In_303,In_170);
or U2059 (N_2059,In_229,In_603);
nand U2060 (N_2060,In_480,In_505);
nor U2061 (N_2061,In_602,In_606);
or U2062 (N_2062,In_637,In_678);
and U2063 (N_2063,In_392,In_670);
and U2064 (N_2064,In_685,In_251);
or U2065 (N_2065,In_80,In_45);
or U2066 (N_2066,In_34,In_603);
nand U2067 (N_2067,In_622,In_191);
or U2068 (N_2068,In_429,In_615);
nor U2069 (N_2069,In_273,In_229);
or U2070 (N_2070,In_230,In_367);
nor U2071 (N_2071,In_454,In_67);
and U2072 (N_2072,In_10,In_473);
nand U2073 (N_2073,In_385,In_543);
nor U2074 (N_2074,In_359,In_118);
nor U2075 (N_2075,In_512,In_580);
xor U2076 (N_2076,In_466,In_232);
nor U2077 (N_2077,In_641,In_690);
nand U2078 (N_2078,In_616,In_330);
nand U2079 (N_2079,In_546,In_0);
or U2080 (N_2080,In_652,In_117);
nor U2081 (N_2081,In_368,In_70);
nor U2082 (N_2082,In_201,In_330);
nand U2083 (N_2083,In_551,In_33);
or U2084 (N_2084,In_744,In_687);
nor U2085 (N_2085,In_67,In_126);
nor U2086 (N_2086,In_711,In_589);
nand U2087 (N_2087,In_141,In_124);
and U2088 (N_2088,In_219,In_694);
and U2089 (N_2089,In_683,In_458);
and U2090 (N_2090,In_462,In_132);
and U2091 (N_2091,In_95,In_639);
or U2092 (N_2092,In_359,In_503);
nor U2093 (N_2093,In_163,In_749);
xnor U2094 (N_2094,In_284,In_485);
or U2095 (N_2095,In_58,In_601);
nor U2096 (N_2096,In_236,In_713);
and U2097 (N_2097,In_54,In_202);
nor U2098 (N_2098,In_496,In_209);
nand U2099 (N_2099,In_85,In_318);
and U2100 (N_2100,In_311,In_132);
nand U2101 (N_2101,In_591,In_194);
xor U2102 (N_2102,In_394,In_578);
or U2103 (N_2103,In_479,In_33);
and U2104 (N_2104,In_133,In_4);
or U2105 (N_2105,In_308,In_16);
nand U2106 (N_2106,In_323,In_333);
xor U2107 (N_2107,In_45,In_636);
nand U2108 (N_2108,In_310,In_344);
or U2109 (N_2109,In_567,In_188);
or U2110 (N_2110,In_290,In_26);
nand U2111 (N_2111,In_210,In_439);
and U2112 (N_2112,In_110,In_602);
or U2113 (N_2113,In_613,In_112);
nand U2114 (N_2114,In_2,In_308);
or U2115 (N_2115,In_408,In_575);
nor U2116 (N_2116,In_527,In_193);
or U2117 (N_2117,In_343,In_567);
nor U2118 (N_2118,In_202,In_230);
or U2119 (N_2119,In_512,In_34);
and U2120 (N_2120,In_749,In_283);
and U2121 (N_2121,In_33,In_31);
nand U2122 (N_2122,In_313,In_81);
nor U2123 (N_2123,In_446,In_157);
nand U2124 (N_2124,In_702,In_102);
nor U2125 (N_2125,In_59,In_303);
and U2126 (N_2126,In_592,In_80);
nand U2127 (N_2127,In_318,In_104);
xnor U2128 (N_2128,In_417,In_333);
nand U2129 (N_2129,In_101,In_624);
or U2130 (N_2130,In_64,In_235);
and U2131 (N_2131,In_161,In_94);
nand U2132 (N_2132,In_122,In_624);
nor U2133 (N_2133,In_627,In_480);
nand U2134 (N_2134,In_427,In_472);
or U2135 (N_2135,In_319,In_342);
and U2136 (N_2136,In_346,In_555);
nand U2137 (N_2137,In_522,In_509);
nand U2138 (N_2138,In_612,In_286);
and U2139 (N_2139,In_229,In_557);
nand U2140 (N_2140,In_55,In_733);
or U2141 (N_2141,In_122,In_424);
or U2142 (N_2142,In_516,In_632);
or U2143 (N_2143,In_284,In_160);
or U2144 (N_2144,In_48,In_660);
xor U2145 (N_2145,In_599,In_92);
and U2146 (N_2146,In_692,In_363);
nand U2147 (N_2147,In_26,In_97);
or U2148 (N_2148,In_637,In_335);
nand U2149 (N_2149,In_589,In_96);
or U2150 (N_2150,In_446,In_148);
nand U2151 (N_2151,In_24,In_723);
nand U2152 (N_2152,In_637,In_30);
nand U2153 (N_2153,In_730,In_116);
nand U2154 (N_2154,In_193,In_328);
and U2155 (N_2155,In_255,In_701);
and U2156 (N_2156,In_600,In_506);
or U2157 (N_2157,In_105,In_373);
nand U2158 (N_2158,In_691,In_662);
nor U2159 (N_2159,In_584,In_666);
nor U2160 (N_2160,In_308,In_81);
nor U2161 (N_2161,In_224,In_685);
or U2162 (N_2162,In_457,In_163);
xnor U2163 (N_2163,In_700,In_78);
nor U2164 (N_2164,In_390,In_173);
nand U2165 (N_2165,In_606,In_118);
xnor U2166 (N_2166,In_558,In_94);
nand U2167 (N_2167,In_107,In_184);
and U2168 (N_2168,In_531,In_642);
nor U2169 (N_2169,In_448,In_661);
and U2170 (N_2170,In_49,In_712);
nand U2171 (N_2171,In_241,In_477);
and U2172 (N_2172,In_283,In_490);
or U2173 (N_2173,In_521,In_60);
or U2174 (N_2174,In_92,In_354);
and U2175 (N_2175,In_248,In_156);
xnor U2176 (N_2176,In_417,In_299);
nand U2177 (N_2177,In_530,In_234);
nor U2178 (N_2178,In_322,In_203);
nor U2179 (N_2179,In_475,In_327);
and U2180 (N_2180,In_493,In_277);
nor U2181 (N_2181,In_231,In_484);
nand U2182 (N_2182,In_730,In_17);
nand U2183 (N_2183,In_247,In_613);
or U2184 (N_2184,In_145,In_427);
nor U2185 (N_2185,In_154,In_277);
xnor U2186 (N_2186,In_637,In_265);
or U2187 (N_2187,In_539,In_131);
nor U2188 (N_2188,In_41,In_440);
nand U2189 (N_2189,In_523,In_641);
or U2190 (N_2190,In_186,In_174);
or U2191 (N_2191,In_116,In_571);
or U2192 (N_2192,In_172,In_121);
or U2193 (N_2193,In_617,In_492);
nor U2194 (N_2194,In_178,In_644);
and U2195 (N_2195,In_552,In_387);
nor U2196 (N_2196,In_298,In_146);
nand U2197 (N_2197,In_709,In_213);
nand U2198 (N_2198,In_19,In_541);
or U2199 (N_2199,In_264,In_746);
or U2200 (N_2200,In_221,In_497);
or U2201 (N_2201,In_454,In_645);
nor U2202 (N_2202,In_388,In_437);
or U2203 (N_2203,In_59,In_626);
and U2204 (N_2204,In_178,In_305);
nand U2205 (N_2205,In_700,In_733);
xor U2206 (N_2206,In_87,In_361);
and U2207 (N_2207,In_93,In_585);
and U2208 (N_2208,In_130,In_239);
nand U2209 (N_2209,In_378,In_237);
nand U2210 (N_2210,In_536,In_562);
and U2211 (N_2211,In_551,In_412);
or U2212 (N_2212,In_515,In_222);
nand U2213 (N_2213,In_495,In_697);
xor U2214 (N_2214,In_121,In_383);
and U2215 (N_2215,In_4,In_519);
nand U2216 (N_2216,In_237,In_48);
nand U2217 (N_2217,In_633,In_300);
or U2218 (N_2218,In_129,In_549);
nand U2219 (N_2219,In_637,In_131);
nand U2220 (N_2220,In_268,In_86);
or U2221 (N_2221,In_550,In_689);
or U2222 (N_2222,In_731,In_627);
or U2223 (N_2223,In_680,In_43);
and U2224 (N_2224,In_181,In_42);
or U2225 (N_2225,In_566,In_207);
nor U2226 (N_2226,In_75,In_532);
nand U2227 (N_2227,In_611,In_296);
and U2228 (N_2228,In_619,In_326);
nor U2229 (N_2229,In_4,In_531);
and U2230 (N_2230,In_694,In_171);
nand U2231 (N_2231,In_647,In_507);
nor U2232 (N_2232,In_91,In_40);
and U2233 (N_2233,In_167,In_229);
nand U2234 (N_2234,In_736,In_670);
and U2235 (N_2235,In_235,In_617);
nor U2236 (N_2236,In_187,In_585);
nand U2237 (N_2237,In_413,In_146);
nand U2238 (N_2238,In_134,In_329);
nand U2239 (N_2239,In_8,In_536);
or U2240 (N_2240,In_530,In_529);
or U2241 (N_2241,In_564,In_200);
and U2242 (N_2242,In_712,In_177);
nor U2243 (N_2243,In_744,In_81);
nor U2244 (N_2244,In_478,In_328);
or U2245 (N_2245,In_623,In_478);
or U2246 (N_2246,In_17,In_704);
xor U2247 (N_2247,In_359,In_342);
or U2248 (N_2248,In_720,In_592);
or U2249 (N_2249,In_206,In_468);
nand U2250 (N_2250,In_183,In_70);
or U2251 (N_2251,In_695,In_579);
nor U2252 (N_2252,In_64,In_622);
nand U2253 (N_2253,In_232,In_30);
nor U2254 (N_2254,In_280,In_261);
and U2255 (N_2255,In_163,In_328);
or U2256 (N_2256,In_14,In_173);
and U2257 (N_2257,In_170,In_423);
and U2258 (N_2258,In_545,In_8);
or U2259 (N_2259,In_121,In_576);
nand U2260 (N_2260,In_60,In_90);
and U2261 (N_2261,In_735,In_307);
and U2262 (N_2262,In_164,In_87);
or U2263 (N_2263,In_318,In_330);
nand U2264 (N_2264,In_648,In_255);
and U2265 (N_2265,In_314,In_337);
and U2266 (N_2266,In_477,In_603);
or U2267 (N_2267,In_639,In_676);
and U2268 (N_2268,In_364,In_101);
nand U2269 (N_2269,In_600,In_337);
and U2270 (N_2270,In_174,In_4);
nor U2271 (N_2271,In_227,In_745);
or U2272 (N_2272,In_364,In_263);
and U2273 (N_2273,In_325,In_515);
xnor U2274 (N_2274,In_418,In_449);
xnor U2275 (N_2275,In_311,In_733);
nor U2276 (N_2276,In_424,In_390);
nor U2277 (N_2277,In_440,In_702);
or U2278 (N_2278,In_135,In_91);
xor U2279 (N_2279,In_493,In_315);
nor U2280 (N_2280,In_149,In_336);
nand U2281 (N_2281,In_311,In_267);
nor U2282 (N_2282,In_629,In_341);
and U2283 (N_2283,In_496,In_743);
and U2284 (N_2284,In_276,In_582);
and U2285 (N_2285,In_474,In_273);
nor U2286 (N_2286,In_427,In_511);
and U2287 (N_2287,In_636,In_600);
and U2288 (N_2288,In_11,In_231);
or U2289 (N_2289,In_70,In_587);
and U2290 (N_2290,In_658,In_726);
and U2291 (N_2291,In_145,In_386);
and U2292 (N_2292,In_518,In_253);
and U2293 (N_2293,In_729,In_155);
nand U2294 (N_2294,In_533,In_422);
nand U2295 (N_2295,In_737,In_8);
and U2296 (N_2296,In_369,In_407);
nand U2297 (N_2297,In_482,In_576);
or U2298 (N_2298,In_186,In_158);
nand U2299 (N_2299,In_308,In_399);
nand U2300 (N_2300,In_287,In_188);
nor U2301 (N_2301,In_309,In_325);
or U2302 (N_2302,In_492,In_693);
nor U2303 (N_2303,In_272,In_565);
and U2304 (N_2304,In_647,In_182);
nand U2305 (N_2305,In_235,In_226);
or U2306 (N_2306,In_398,In_88);
nor U2307 (N_2307,In_37,In_732);
nor U2308 (N_2308,In_634,In_517);
nand U2309 (N_2309,In_581,In_458);
and U2310 (N_2310,In_281,In_87);
nor U2311 (N_2311,In_22,In_291);
nand U2312 (N_2312,In_400,In_123);
and U2313 (N_2313,In_60,In_577);
and U2314 (N_2314,In_175,In_285);
and U2315 (N_2315,In_553,In_11);
nor U2316 (N_2316,In_368,In_351);
and U2317 (N_2317,In_712,In_645);
or U2318 (N_2318,In_407,In_636);
nor U2319 (N_2319,In_519,In_469);
nor U2320 (N_2320,In_102,In_704);
and U2321 (N_2321,In_691,In_417);
or U2322 (N_2322,In_284,In_652);
nand U2323 (N_2323,In_342,In_537);
nand U2324 (N_2324,In_160,In_632);
and U2325 (N_2325,In_371,In_613);
xor U2326 (N_2326,In_730,In_637);
xor U2327 (N_2327,In_682,In_237);
or U2328 (N_2328,In_455,In_346);
nor U2329 (N_2329,In_359,In_427);
nand U2330 (N_2330,In_131,In_344);
or U2331 (N_2331,In_707,In_559);
nand U2332 (N_2332,In_148,In_482);
and U2333 (N_2333,In_731,In_677);
nor U2334 (N_2334,In_474,In_694);
nand U2335 (N_2335,In_355,In_605);
and U2336 (N_2336,In_733,In_434);
nand U2337 (N_2337,In_385,In_285);
or U2338 (N_2338,In_307,In_667);
nand U2339 (N_2339,In_185,In_86);
and U2340 (N_2340,In_221,In_413);
nor U2341 (N_2341,In_49,In_117);
nor U2342 (N_2342,In_480,In_72);
or U2343 (N_2343,In_530,In_491);
nor U2344 (N_2344,In_285,In_150);
or U2345 (N_2345,In_158,In_135);
nor U2346 (N_2346,In_667,In_181);
and U2347 (N_2347,In_54,In_311);
or U2348 (N_2348,In_208,In_635);
nand U2349 (N_2349,In_236,In_179);
or U2350 (N_2350,In_476,In_678);
or U2351 (N_2351,In_405,In_346);
and U2352 (N_2352,In_586,In_61);
or U2353 (N_2353,In_197,In_199);
nand U2354 (N_2354,In_140,In_581);
and U2355 (N_2355,In_335,In_711);
nand U2356 (N_2356,In_388,In_159);
nor U2357 (N_2357,In_201,In_218);
nor U2358 (N_2358,In_407,In_223);
nand U2359 (N_2359,In_434,In_382);
xor U2360 (N_2360,In_681,In_332);
and U2361 (N_2361,In_595,In_7);
or U2362 (N_2362,In_418,In_319);
or U2363 (N_2363,In_673,In_417);
nand U2364 (N_2364,In_192,In_334);
nand U2365 (N_2365,In_495,In_624);
xnor U2366 (N_2366,In_112,In_519);
and U2367 (N_2367,In_650,In_621);
nand U2368 (N_2368,In_146,In_549);
nand U2369 (N_2369,In_143,In_252);
xor U2370 (N_2370,In_178,In_373);
nand U2371 (N_2371,In_596,In_696);
and U2372 (N_2372,In_29,In_748);
or U2373 (N_2373,In_391,In_322);
nor U2374 (N_2374,In_724,In_618);
or U2375 (N_2375,In_55,In_70);
nor U2376 (N_2376,In_213,In_433);
nor U2377 (N_2377,In_404,In_506);
nor U2378 (N_2378,In_745,In_586);
and U2379 (N_2379,In_572,In_305);
nor U2380 (N_2380,In_96,In_186);
or U2381 (N_2381,In_603,In_711);
nand U2382 (N_2382,In_596,In_463);
or U2383 (N_2383,In_637,In_119);
or U2384 (N_2384,In_691,In_502);
or U2385 (N_2385,In_313,In_308);
nor U2386 (N_2386,In_103,In_476);
or U2387 (N_2387,In_381,In_314);
nor U2388 (N_2388,In_589,In_164);
or U2389 (N_2389,In_687,In_67);
and U2390 (N_2390,In_310,In_145);
nand U2391 (N_2391,In_487,In_402);
nor U2392 (N_2392,In_414,In_225);
nand U2393 (N_2393,In_276,In_605);
nor U2394 (N_2394,In_460,In_351);
nand U2395 (N_2395,In_157,In_671);
nor U2396 (N_2396,In_692,In_689);
or U2397 (N_2397,In_690,In_605);
nor U2398 (N_2398,In_555,In_56);
nor U2399 (N_2399,In_344,In_452);
nand U2400 (N_2400,In_190,In_372);
or U2401 (N_2401,In_387,In_541);
or U2402 (N_2402,In_0,In_156);
and U2403 (N_2403,In_151,In_564);
nor U2404 (N_2404,In_538,In_330);
nand U2405 (N_2405,In_165,In_506);
or U2406 (N_2406,In_398,In_173);
and U2407 (N_2407,In_431,In_254);
nor U2408 (N_2408,In_172,In_503);
nor U2409 (N_2409,In_99,In_464);
nand U2410 (N_2410,In_489,In_212);
and U2411 (N_2411,In_320,In_598);
nor U2412 (N_2412,In_369,In_70);
nand U2413 (N_2413,In_380,In_595);
xnor U2414 (N_2414,In_518,In_668);
nor U2415 (N_2415,In_369,In_104);
nor U2416 (N_2416,In_317,In_342);
nand U2417 (N_2417,In_112,In_168);
and U2418 (N_2418,In_369,In_601);
and U2419 (N_2419,In_272,In_268);
or U2420 (N_2420,In_423,In_404);
nand U2421 (N_2421,In_516,In_227);
nor U2422 (N_2422,In_336,In_55);
xnor U2423 (N_2423,In_146,In_302);
nand U2424 (N_2424,In_411,In_482);
nor U2425 (N_2425,In_224,In_515);
nand U2426 (N_2426,In_519,In_64);
nand U2427 (N_2427,In_181,In_142);
and U2428 (N_2428,In_442,In_451);
and U2429 (N_2429,In_348,In_88);
nand U2430 (N_2430,In_679,In_34);
nor U2431 (N_2431,In_615,In_329);
nor U2432 (N_2432,In_573,In_389);
nor U2433 (N_2433,In_472,In_60);
or U2434 (N_2434,In_51,In_341);
or U2435 (N_2435,In_724,In_508);
xor U2436 (N_2436,In_327,In_281);
nor U2437 (N_2437,In_259,In_404);
and U2438 (N_2438,In_106,In_459);
nand U2439 (N_2439,In_87,In_647);
and U2440 (N_2440,In_544,In_576);
and U2441 (N_2441,In_532,In_542);
or U2442 (N_2442,In_118,In_236);
nor U2443 (N_2443,In_563,In_294);
nor U2444 (N_2444,In_390,In_218);
nor U2445 (N_2445,In_371,In_647);
and U2446 (N_2446,In_102,In_431);
and U2447 (N_2447,In_283,In_378);
nor U2448 (N_2448,In_27,In_703);
nand U2449 (N_2449,In_351,In_520);
nor U2450 (N_2450,In_336,In_47);
or U2451 (N_2451,In_544,In_305);
nand U2452 (N_2452,In_106,In_622);
or U2453 (N_2453,In_557,In_192);
and U2454 (N_2454,In_735,In_736);
nor U2455 (N_2455,In_639,In_741);
nand U2456 (N_2456,In_437,In_512);
nor U2457 (N_2457,In_210,In_86);
or U2458 (N_2458,In_512,In_162);
nand U2459 (N_2459,In_532,In_424);
and U2460 (N_2460,In_563,In_541);
nand U2461 (N_2461,In_538,In_480);
nand U2462 (N_2462,In_709,In_94);
nand U2463 (N_2463,In_447,In_728);
or U2464 (N_2464,In_181,In_308);
nand U2465 (N_2465,In_118,In_595);
and U2466 (N_2466,In_79,In_143);
nand U2467 (N_2467,In_140,In_275);
nor U2468 (N_2468,In_164,In_193);
nor U2469 (N_2469,In_586,In_351);
and U2470 (N_2470,In_729,In_642);
nand U2471 (N_2471,In_152,In_121);
nor U2472 (N_2472,In_532,In_659);
nor U2473 (N_2473,In_514,In_186);
or U2474 (N_2474,In_578,In_471);
nor U2475 (N_2475,In_694,In_112);
and U2476 (N_2476,In_595,In_730);
or U2477 (N_2477,In_475,In_640);
nor U2478 (N_2478,In_542,In_442);
or U2479 (N_2479,In_286,In_152);
or U2480 (N_2480,In_400,In_218);
or U2481 (N_2481,In_676,In_130);
nor U2482 (N_2482,In_634,In_54);
nand U2483 (N_2483,In_671,In_76);
and U2484 (N_2484,In_320,In_208);
nand U2485 (N_2485,In_309,In_4);
and U2486 (N_2486,In_636,In_410);
nor U2487 (N_2487,In_489,In_114);
or U2488 (N_2488,In_195,In_543);
and U2489 (N_2489,In_152,In_353);
or U2490 (N_2490,In_251,In_81);
xnor U2491 (N_2491,In_646,In_5);
nand U2492 (N_2492,In_378,In_297);
nand U2493 (N_2493,In_19,In_153);
nor U2494 (N_2494,In_186,In_375);
nand U2495 (N_2495,In_366,In_228);
and U2496 (N_2496,In_43,In_657);
nand U2497 (N_2497,In_697,In_129);
or U2498 (N_2498,In_742,In_22);
nand U2499 (N_2499,In_122,In_423);
or U2500 (N_2500,N_2088,N_2337);
nand U2501 (N_2501,N_1877,N_968);
or U2502 (N_2502,N_290,N_84);
and U2503 (N_2503,N_986,N_2129);
and U2504 (N_2504,N_698,N_625);
or U2505 (N_2505,N_1982,N_2352);
or U2506 (N_2506,N_1572,N_568);
nor U2507 (N_2507,N_1955,N_1782);
and U2508 (N_2508,N_2307,N_1013);
xnor U2509 (N_2509,N_509,N_2189);
nor U2510 (N_2510,N_268,N_734);
or U2511 (N_2511,N_862,N_1454);
nor U2512 (N_2512,N_1661,N_1904);
and U2513 (N_2513,N_471,N_832);
and U2514 (N_2514,N_876,N_532);
nor U2515 (N_2515,N_487,N_1155);
or U2516 (N_2516,N_1591,N_1914);
nand U2517 (N_2517,N_2494,N_1519);
and U2518 (N_2518,N_1028,N_2117);
nand U2519 (N_2519,N_114,N_230);
nor U2520 (N_2520,N_1565,N_1074);
nor U2521 (N_2521,N_2095,N_712);
or U2522 (N_2522,N_1638,N_1487);
nand U2523 (N_2523,N_443,N_737);
and U2524 (N_2524,N_482,N_933);
nand U2525 (N_2525,N_1405,N_2047);
or U2526 (N_2526,N_234,N_939);
or U2527 (N_2527,N_785,N_1919);
or U2528 (N_2528,N_1809,N_1459);
or U2529 (N_2529,N_305,N_152);
nand U2530 (N_2530,N_2140,N_559);
nor U2531 (N_2531,N_970,N_502);
nor U2532 (N_2532,N_1320,N_1732);
and U2533 (N_2533,N_2378,N_1184);
and U2534 (N_2534,N_2439,N_2179);
nor U2535 (N_2535,N_446,N_1107);
xor U2536 (N_2536,N_78,N_895);
nor U2537 (N_2537,N_1431,N_1747);
nor U2538 (N_2538,N_924,N_815);
and U2539 (N_2539,N_730,N_1892);
nor U2540 (N_2540,N_1868,N_1059);
nand U2541 (N_2541,N_30,N_1971);
and U2542 (N_2542,N_1635,N_1962);
or U2543 (N_2543,N_14,N_1414);
nor U2544 (N_2544,N_936,N_1835);
nor U2545 (N_2545,N_1704,N_600);
and U2546 (N_2546,N_1945,N_2050);
nand U2547 (N_2547,N_907,N_1277);
nor U2548 (N_2548,N_2321,N_2397);
nor U2549 (N_2549,N_1413,N_1273);
nor U2550 (N_2550,N_1756,N_2027);
or U2551 (N_2551,N_1621,N_2485);
and U2552 (N_2552,N_636,N_1167);
and U2553 (N_2553,N_997,N_1967);
nor U2554 (N_2554,N_2417,N_1777);
and U2555 (N_2555,N_2253,N_1372);
and U2556 (N_2556,N_1946,N_1048);
nor U2557 (N_2557,N_1585,N_547);
or U2558 (N_2558,N_1518,N_535);
nor U2559 (N_2559,N_165,N_791);
nor U2560 (N_2560,N_1345,N_1037);
nand U2561 (N_2561,N_29,N_411);
or U2562 (N_2562,N_2454,N_1287);
nand U2563 (N_2563,N_1787,N_941);
nor U2564 (N_2564,N_2142,N_2053);
or U2565 (N_2565,N_937,N_1568);
nor U2566 (N_2566,N_1795,N_453);
and U2567 (N_2567,N_407,N_1103);
or U2568 (N_2568,N_2110,N_2167);
nand U2569 (N_2569,N_250,N_858);
nand U2570 (N_2570,N_1639,N_197);
and U2571 (N_2571,N_2232,N_423);
nand U2572 (N_2572,N_386,N_1783);
and U2573 (N_2573,N_1199,N_464);
and U2574 (N_2574,N_665,N_1631);
or U2575 (N_2575,N_1110,N_893);
or U2576 (N_2576,N_1402,N_2305);
and U2577 (N_2577,N_308,N_479);
nand U2578 (N_2578,N_1820,N_2162);
nand U2579 (N_2579,N_156,N_1853);
and U2580 (N_2580,N_384,N_1563);
nand U2581 (N_2581,N_1357,N_208);
nor U2582 (N_2582,N_1736,N_905);
and U2583 (N_2583,N_455,N_387);
nor U2584 (N_2584,N_1776,N_2296);
and U2585 (N_2585,N_321,N_2301);
and U2586 (N_2586,N_1988,N_1913);
xor U2587 (N_2587,N_1089,N_596);
nor U2588 (N_2588,N_1505,N_1856);
and U2589 (N_2589,N_1440,N_531);
and U2590 (N_2590,N_1527,N_2463);
nand U2591 (N_2591,N_2197,N_2492);
or U2592 (N_2592,N_518,N_1650);
or U2593 (N_2593,N_1220,N_2458);
and U2594 (N_2594,N_1181,N_796);
or U2595 (N_2595,N_2278,N_454);
nand U2596 (N_2596,N_2353,N_2498);
and U2597 (N_2597,N_703,N_2123);
or U2598 (N_2598,N_1701,N_2244);
nand U2599 (N_2599,N_633,N_2163);
and U2600 (N_2600,N_161,N_2132);
nand U2601 (N_2601,N_1232,N_1275);
nor U2602 (N_2602,N_1739,N_1011);
and U2603 (N_2603,N_1611,N_452);
or U2604 (N_2604,N_719,N_1290);
or U2605 (N_2605,N_2032,N_1619);
and U2606 (N_2606,N_2291,N_817);
and U2607 (N_2607,N_2039,N_1685);
nor U2608 (N_2608,N_163,N_2255);
nand U2609 (N_2609,N_1449,N_2090);
and U2610 (N_2610,N_526,N_344);
or U2611 (N_2611,N_133,N_853);
nand U2612 (N_2612,N_34,N_909);
and U2613 (N_2613,N_1969,N_356);
nor U2614 (N_2614,N_866,N_147);
nand U2615 (N_2615,N_99,N_558);
nor U2616 (N_2616,N_1396,N_1420);
and U2617 (N_2617,N_1212,N_1806);
nand U2618 (N_2618,N_974,N_1972);
nand U2619 (N_2619,N_1911,N_2387);
nand U2620 (N_2620,N_548,N_1418);
nand U2621 (N_2621,N_2225,N_1271);
and U2622 (N_2622,N_962,N_638);
or U2623 (N_2623,N_604,N_555);
nor U2624 (N_2624,N_1857,N_1131);
and U2625 (N_2625,N_821,N_2106);
nand U2626 (N_2626,N_887,N_1860);
and U2627 (N_2627,N_1258,N_1239);
and U2628 (N_2628,N_337,N_2407);
and U2629 (N_2629,N_1375,N_1775);
and U2630 (N_2630,N_2011,N_2356);
nand U2631 (N_2631,N_1965,N_1778);
nand U2632 (N_2632,N_1752,N_1749);
nor U2633 (N_2633,N_2341,N_1762);
and U2634 (N_2634,N_1342,N_2384);
nor U2635 (N_2635,N_507,N_819);
nand U2636 (N_2636,N_162,N_196);
nand U2637 (N_2637,N_2234,N_2351);
or U2638 (N_2638,N_794,N_262);
nor U2639 (N_2639,N_1368,N_173);
nor U2640 (N_2640,N_1690,N_808);
nand U2641 (N_2641,N_1132,N_1818);
and U2642 (N_2642,N_1244,N_1664);
or U2643 (N_2643,N_708,N_1143);
and U2644 (N_2644,N_2187,N_2456);
or U2645 (N_2645,N_105,N_1090);
or U2646 (N_2646,N_1634,N_103);
nor U2647 (N_2647,N_2005,N_1076);
nor U2648 (N_2648,N_1334,N_505);
nand U2649 (N_2649,N_1769,N_247);
and U2650 (N_2650,N_2248,N_1313);
and U2651 (N_2651,N_1931,N_630);
nand U2652 (N_2652,N_1697,N_884);
nand U2653 (N_2653,N_1360,N_1146);
or U2654 (N_2654,N_679,N_1502);
or U2655 (N_2655,N_657,N_1168);
nor U2656 (N_2656,N_2450,N_1054);
nor U2657 (N_2657,N_1427,N_488);
nor U2658 (N_2658,N_850,N_1937);
nor U2659 (N_2659,N_2486,N_1622);
nor U2660 (N_2660,N_1719,N_1952);
and U2661 (N_2661,N_799,N_1178);
and U2662 (N_2662,N_1772,N_1468);
nor U2663 (N_2663,N_1633,N_233);
and U2664 (N_2664,N_1022,N_367);
nor U2665 (N_2665,N_919,N_9);
nand U2666 (N_2666,N_1763,N_626);
or U2667 (N_2667,N_2262,N_2211);
nor U2668 (N_2668,N_2017,N_2335);
nor U2669 (N_2669,N_1123,N_2467);
and U2670 (N_2670,N_1890,N_1388);
nor U2671 (N_2671,N_1524,N_1326);
nand U2672 (N_2672,N_2431,N_1190);
nand U2673 (N_2673,N_959,N_877);
or U2674 (N_2674,N_61,N_503);
and U2675 (N_2675,N_1259,N_134);
or U2676 (N_2676,N_1014,N_1461);
and U2677 (N_2677,N_217,N_978);
nand U2678 (N_2678,N_956,N_1490);
nand U2679 (N_2679,N_2202,N_660);
nand U2680 (N_2680,N_754,N_1613);
nand U2681 (N_2681,N_1497,N_1246);
or U2682 (N_2682,N_2459,N_1799);
nand U2683 (N_2683,N_1715,N_1285);
nand U2684 (N_2684,N_2041,N_2394);
nor U2685 (N_2685,N_529,N_709);
xnor U2686 (N_2686,N_1233,N_259);
and U2687 (N_2687,N_766,N_969);
and U2688 (N_2688,N_1910,N_1863);
and U2689 (N_2689,N_1636,N_135);
and U2690 (N_2690,N_894,N_91);
and U2691 (N_2691,N_699,N_1520);
nand U2692 (N_2692,N_1078,N_1506);
or U2693 (N_2693,N_1223,N_35);
or U2694 (N_2694,N_1925,N_1198);
and U2695 (N_2695,N_226,N_494);
and U2696 (N_2696,N_2020,N_1305);
nand U2697 (N_2697,N_788,N_1169);
xnor U2698 (N_2698,N_85,N_2084);
nand U2699 (N_2699,N_1175,N_774);
and U2700 (N_2700,N_1987,N_1475);
and U2701 (N_2701,N_767,N_2121);
or U2702 (N_2702,N_1121,N_89);
nor U2703 (N_2703,N_1786,N_2379);
nand U2704 (N_2704,N_87,N_2361);
or U2705 (N_2705,N_1219,N_174);
or U2706 (N_2706,N_1193,N_2007);
or U2707 (N_2707,N_622,N_982);
nor U2708 (N_2708,N_2477,N_2266);
nand U2709 (N_2709,N_44,N_566);
and U2710 (N_2710,N_2240,N_1446);
and U2711 (N_2711,N_1927,N_587);
nor U2712 (N_2712,N_92,N_1185);
nor U2713 (N_2713,N_1555,N_257);
nand U2714 (N_2714,N_1416,N_2480);
or U2715 (N_2715,N_1679,N_1836);
nor U2716 (N_2716,N_1928,N_1828);
nor U2717 (N_2717,N_425,N_1854);
nand U2718 (N_2718,N_616,N_2009);
nand U2719 (N_2719,N_2437,N_610);
nor U2720 (N_2720,N_789,N_760);
and U2721 (N_2721,N_1130,N_691);
or U2722 (N_2722,N_1789,N_70);
nand U2723 (N_2723,N_750,N_183);
nand U2724 (N_2724,N_2228,N_1392);
nand U2725 (N_2725,N_1730,N_1589);
and U2726 (N_2726,N_1323,N_2408);
nor U2727 (N_2727,N_641,N_1324);
nor U2728 (N_2728,N_1383,N_1709);
and U2729 (N_2729,N_1660,N_1231);
and U2730 (N_2730,N_2029,N_601);
nand U2731 (N_2731,N_846,N_2306);
nand U2732 (N_2732,N_1872,N_830);
nor U2733 (N_2733,N_926,N_560);
and U2734 (N_2734,N_1105,N_649);
and U2735 (N_2735,N_802,N_2194);
and U2736 (N_2736,N_820,N_2182);
nor U2737 (N_2737,N_1848,N_1455);
or U2738 (N_2738,N_1738,N_2038);
or U2739 (N_2739,N_1288,N_705);
nand U2740 (N_2740,N_2369,N_2413);
nor U2741 (N_2741,N_977,N_2183);
and U2742 (N_2742,N_1302,N_2471);
or U2743 (N_2743,N_1441,N_1678);
and U2744 (N_2744,N_1163,N_2006);
and U2745 (N_2745,N_449,N_110);
or U2746 (N_2746,N_1917,N_2282);
and U2747 (N_2747,N_1476,N_198);
or U2748 (N_2748,N_722,N_2375);
and U2749 (N_2749,N_261,N_2340);
nor U2750 (N_2750,N_1055,N_1614);
and U2751 (N_2751,N_2294,N_757);
or U2752 (N_2752,N_2316,N_2448);
nor U2753 (N_2753,N_1746,N_1080);
nor U2754 (N_2754,N_2287,N_2256);
or U2755 (N_2755,N_205,N_711);
nor U2756 (N_2756,N_281,N_1874);
or U2757 (N_2757,N_1210,N_1997);
xnor U2758 (N_2758,N_1717,N_2388);
nand U2759 (N_2759,N_2461,N_2160);
nand U2760 (N_2760,N_779,N_724);
or U2761 (N_2761,N_1807,N_836);
and U2762 (N_2762,N_1049,N_1844);
or U2763 (N_2763,N_1469,N_1587);
and U2764 (N_2764,N_1453,N_1092);
nor U2765 (N_2765,N_1692,N_1617);
nor U2766 (N_2766,N_1842,N_2409);
nor U2767 (N_2767,N_2138,N_1279);
nand U2768 (N_2768,N_2345,N_120);
nand U2769 (N_2769,N_1194,N_1124);
and U2770 (N_2770,N_1995,N_872);
or U2771 (N_2771,N_42,N_748);
nand U2772 (N_2772,N_2373,N_1716);
or U2773 (N_2773,N_1008,N_662);
or U2774 (N_2774,N_975,N_984);
or U2775 (N_2775,N_2231,N_733);
nand U2776 (N_2776,N_949,N_2243);
or U2777 (N_2777,N_390,N_1827);
xor U2778 (N_2778,N_2175,N_1042);
nor U2779 (N_2779,N_311,N_139);
and U2780 (N_2780,N_2393,N_383);
and U2781 (N_2781,N_1733,N_914);
and U2782 (N_2782,N_1098,N_1333);
nor U2783 (N_2783,N_825,N_979);
nor U2784 (N_2784,N_1542,N_59);
and U2785 (N_2785,N_618,N_1083);
and U2786 (N_2786,N_228,N_1269);
and U2787 (N_2787,N_379,N_170);
and U2788 (N_2788,N_1794,N_973);
or U2789 (N_2789,N_2030,N_1801);
and U2790 (N_2790,N_410,N_857);
nor U2791 (N_2791,N_611,N_2031);
nand U2792 (N_2792,N_2441,N_382);
nand U2793 (N_2793,N_1349,N_689);
nand U2794 (N_2794,N_1951,N_1415);
nor U2795 (N_2795,N_852,N_781);
nand U2796 (N_2796,N_1980,N_1020);
nand U2797 (N_2797,N_950,N_348);
or U2798 (N_2798,N_277,N_1241);
nor U2799 (N_2799,N_73,N_2045);
and U2800 (N_2800,N_2258,N_2060);
or U2801 (N_2801,N_421,N_1695);
and U2802 (N_2802,N_1039,N_1669);
nand U2803 (N_2803,N_1126,N_1532);
and U2804 (N_2804,N_182,N_2216);
and U2805 (N_2805,N_336,N_359);
nor U2806 (N_2806,N_1430,N_2099);
and U2807 (N_2807,N_1566,N_1332);
nand U2808 (N_2808,N_2024,N_1979);
and U2809 (N_2809,N_1940,N_1850);
nand U2810 (N_2810,N_694,N_1843);
and U2811 (N_2811,N_1050,N_851);
or U2812 (N_2812,N_1816,N_957);
or U2813 (N_2813,N_2018,N_2086);
or U2814 (N_2814,N_1165,N_1869);
or U2815 (N_2815,N_1765,N_1580);
nor U2816 (N_2816,N_0,N_178);
nand U2817 (N_2817,N_1521,N_1706);
and U2818 (N_2818,N_184,N_238);
nor U2819 (N_2819,N_631,N_2418);
or U2820 (N_2820,N_2276,N_1329);
and U2821 (N_2821,N_2205,N_546);
nor U2822 (N_2822,N_1941,N_1379);
nand U2823 (N_2823,N_1289,N_829);
and U2824 (N_2824,N_1522,N_1113);
and U2825 (N_2825,N_755,N_2396);
or U2826 (N_2826,N_1016,N_2360);
or U2827 (N_2827,N_1391,N_827);
or U2828 (N_2828,N_2219,N_373);
nor U2829 (N_2829,N_1834,N_1768);
nand U2830 (N_2830,N_1883,N_1017);
xor U2831 (N_2831,N_445,N_1295);
nand U2832 (N_2832,N_1545,N_1590);
and U2833 (N_2833,N_1494,N_1671);
or U2834 (N_2834,N_1096,N_805);
or U2835 (N_2835,N_2136,N_1511);
nor U2836 (N_2836,N_874,N_412);
nor U2837 (N_2837,N_1084,N_242);
nor U2838 (N_2838,N_116,N_504);
nor U2839 (N_2839,N_1403,N_897);
and U2840 (N_2840,N_1463,N_1560);
nor U2841 (N_2841,N_1479,N_1918);
and U2842 (N_2842,N_22,N_1297);
or U2843 (N_2843,N_391,N_80);
or U2844 (N_2844,N_1546,N_1451);
or U2845 (N_2845,N_2073,N_1822);
nand U2846 (N_2846,N_300,N_345);
or U2847 (N_2847,N_1993,N_2333);
and U2848 (N_2848,N_839,N_1564);
nor U2849 (N_2849,N_2453,N_438);
or U2850 (N_2850,N_1376,N_540);
nor U2851 (N_2851,N_868,N_1426);
nor U2852 (N_2852,N_1529,N_227);
nand U2853 (N_2853,N_1906,N_324);
or U2854 (N_2854,N_25,N_1482);
and U2855 (N_2855,N_1102,N_1129);
and U2856 (N_2856,N_1120,N_1133);
nor U2857 (N_2857,N_1743,N_119);
nor U2858 (N_2858,N_2004,N_2066);
or U2859 (N_2859,N_1314,N_1003);
nor U2860 (N_2860,N_1724,N_717);
nor U2861 (N_2861,N_1935,N_1653);
nand U2862 (N_2862,N_557,N_253);
and U2863 (N_2863,N_1895,N_63);
or U2864 (N_2864,N_2166,N_988);
nor U2865 (N_2865,N_1294,N_1203);
nand U2866 (N_2866,N_1432,N_573);
or U2867 (N_2867,N_1009,N_1139);
nand U2868 (N_2868,N_339,N_1659);
nand U2869 (N_2869,N_1336,N_692);
or U2870 (N_2870,N_1171,N_1977);
nand U2871 (N_2871,N_1921,N_741);
nor U2872 (N_2872,N_1007,N_813);
nand U2873 (N_2873,N_2368,N_2227);
nor U2874 (N_2874,N_1112,N_759);
nand U2875 (N_2875,N_681,N_2101);
nand U2876 (N_2876,N_1371,N_1046);
nand U2877 (N_2877,N_1643,N_1579);
and U2878 (N_2878,N_710,N_2043);
nand U2879 (N_2879,N_2061,N_2082);
nor U2880 (N_2880,N_112,N_1051);
and U2881 (N_2881,N_1923,N_646);
nand U2882 (N_2882,N_2199,N_1151);
nand U2883 (N_2883,N_2108,N_896);
or U2884 (N_2884,N_1849,N_1672);
nor U2885 (N_2885,N_420,N_334);
xor U2886 (N_2886,N_1681,N_1975);
nor U2887 (N_2887,N_1605,N_744);
nand U2888 (N_2888,N_659,N_2493);
nor U2889 (N_2889,N_960,N_1788);
or U2890 (N_2890,N_1157,N_484);
and U2891 (N_2891,N_623,N_1994);
and U2892 (N_2892,N_2295,N_1040);
nand U2893 (N_2893,N_7,N_1693);
nor U2894 (N_2894,N_1839,N_8);
and U2895 (N_2895,N_58,N_2057);
or U2896 (N_2896,N_1548,N_512);
and U2897 (N_2897,N_39,N_280);
nand U2898 (N_2898,N_1832,N_2481);
nand U2899 (N_2899,N_1798,N_921);
nor U2900 (N_2900,N_81,N_388);
or U2901 (N_2901,N_2089,N_911);
and U2902 (N_2902,N_1553,N_2042);
or U2903 (N_2903,N_1478,N_1531);
and U2904 (N_2904,N_2303,N_1864);
nand U2905 (N_2905,N_1991,N_1640);
nor U2906 (N_2906,N_1144,N_1929);
nor U2907 (N_2907,N_1260,N_1227);
or U2908 (N_2908,N_291,N_922);
and U2909 (N_2909,N_447,N_577);
xnor U2910 (N_2910,N_628,N_1894);
and U2911 (N_2911,N_1445,N_270);
and U2912 (N_2912,N_1472,N_295);
and U2913 (N_2913,N_1840,N_435);
or U2914 (N_2914,N_2400,N_111);
nor U2915 (N_2915,N_1412,N_2170);
and U2916 (N_2916,N_1351,N_2188);
and U2917 (N_2917,N_1108,N_2449);
nor U2918 (N_2918,N_350,N_1343);
nand U2919 (N_2919,N_1740,N_2280);
nor U2920 (N_2920,N_1556,N_1754);
nand U2921 (N_2921,N_2403,N_450);
or U2922 (N_2922,N_1593,N_963);
nor U2923 (N_2923,N_1547,N_1069);
or U2924 (N_2924,N_849,N_1915);
nand U2925 (N_2925,N_2433,N_1065);
and U2926 (N_2926,N_782,N_1907);
or U2927 (N_2927,N_713,N_287);
and U2928 (N_2928,N_1025,N_609);
nor U2929 (N_2929,N_1214,N_758);
nor U2930 (N_2930,N_2048,N_1606);
or U2931 (N_2931,N_140,N_1408);
nand U2932 (N_2932,N_1073,N_181);
and U2933 (N_2933,N_1201,N_780);
nor U2934 (N_2934,N_1251,N_1213);
nor U2935 (N_2935,N_1905,N_1041);
or U2936 (N_2936,N_2016,N_1189);
nand U2937 (N_2937,N_322,N_840);
and U2938 (N_2938,N_1488,N_523);
and U2939 (N_2939,N_1082,N_508);
or U2940 (N_2940,N_1934,N_915);
nor U2941 (N_2941,N_1027,N_2425);
xnor U2942 (N_2942,N_2195,N_580);
nand U2943 (N_2943,N_2468,N_2128);
nand U2944 (N_2944,N_2065,N_885);
xnor U2945 (N_2945,N_327,N_860);
and U2946 (N_2946,N_82,N_1081);
nor U2947 (N_2947,N_776,N_591);
and U2948 (N_2948,N_833,N_2440);
or U2949 (N_2949,N_160,N_961);
and U2950 (N_2950,N_214,N_946);
and U2951 (N_2951,N_229,N_899);
nor U2952 (N_2952,N_795,N_64);
nand U2953 (N_2953,N_166,N_1192);
nand U2954 (N_2954,N_2134,N_1578);
nand U2955 (N_2955,N_1068,N_1793);
and U2956 (N_2956,N_522,N_125);
or U2957 (N_2957,N_2247,N_1604);
and U2958 (N_2958,N_1549,N_2028);
and U2959 (N_2959,N_2092,N_481);
nor U2960 (N_2960,N_627,N_1757);
or U2961 (N_2961,N_1533,N_1099);
and U2962 (N_2962,N_2318,N_570);
nor U2963 (N_2963,N_714,N_2081);
or U2964 (N_2964,N_151,N_1085);
nand U2965 (N_2965,N_2357,N_1974);
or U2966 (N_2966,N_999,N_2242);
and U2967 (N_2967,N_702,N_1615);
nand U2968 (N_2968,N_1276,N_1428);
and U2969 (N_2969,N_1452,N_1183);
and U2970 (N_2970,N_1610,N_727);
nor U2971 (N_2971,N_4,N_2422);
or U2972 (N_2972,N_10,N_521);
nor U2973 (N_2973,N_1903,N_480);
nor U2974 (N_2974,N_158,N_1395);
and U2975 (N_2975,N_1154,N_989);
nor U2976 (N_2976,N_442,N_686);
or U2977 (N_2977,N_1460,N_927);
and U2978 (N_2978,N_971,N_2259);
and U2979 (N_2979,N_1922,N_1912);
and U2980 (N_2980,N_2217,N_1176);
nor U2981 (N_2981,N_2328,N_221);
and U2982 (N_2982,N_1662,N_1398);
and U2983 (N_2983,N_695,N_923);
nor U2984 (N_2984,N_415,N_1422);
or U2985 (N_2985,N_424,N_108);
and U2986 (N_2986,N_444,N_2118);
nand U2987 (N_2987,N_2405,N_154);
nand U2988 (N_2988,N_2487,N_1557);
or U2989 (N_2989,N_793,N_1741);
and U2990 (N_2990,N_643,N_500);
nor U2991 (N_2991,N_2213,N_574);
nand U2992 (N_2992,N_2473,N_2430);
or U2993 (N_2993,N_426,N_680);
nand U2994 (N_2994,N_211,N_739);
nand U2995 (N_2995,N_1325,N_1767);
or U2996 (N_2996,N_2046,N_2212);
and U2997 (N_2997,N_1963,N_1675);
nor U2998 (N_2998,N_770,N_2358);
and U2999 (N_2999,N_1071,N_298);
or U3000 (N_3000,N_806,N_1734);
or U3001 (N_3001,N_475,N_2392);
or U3002 (N_3002,N_368,N_2386);
and U3003 (N_3003,N_525,N_683);
and U3004 (N_3004,N_272,N_1286);
and U3005 (N_3005,N_1718,N_1471);
nor U3006 (N_3006,N_474,N_1808);
and U3007 (N_3007,N_1278,N_17);
nor U3008 (N_3008,N_380,N_477);
nand U3009 (N_3009,N_392,N_980);
and U3010 (N_3010,N_394,N_457);
xnor U3011 (N_3011,N_2338,N_1386);
nand U3012 (N_3012,N_289,N_1909);
or U3013 (N_3013,N_1920,N_100);
nor U3014 (N_3014,N_787,N_1682);
or U3015 (N_3015,N_1599,N_2355);
nand U3016 (N_3016,N_1135,N_847);
and U3017 (N_3017,N_1688,N_844);
nor U3018 (N_3018,N_2033,N_1932);
nor U3019 (N_3019,N_293,N_1562);
nor U3020 (N_3020,N_2210,N_1939);
nand U3021 (N_3021,N_2435,N_878);
nor U3022 (N_3022,N_1796,N_1380);
and U3023 (N_3023,N_1270,N_2349);
or U3024 (N_3024,N_1296,N_146);
or U3025 (N_3025,N_908,N_1683);
or U3026 (N_3026,N_2474,N_2124);
or U3027 (N_3027,N_1652,N_718);
and U3028 (N_3028,N_2096,N_1871);
and U3029 (N_3029,N_2331,N_1526);
nor U3030 (N_3030,N_448,N_288);
and U3031 (N_3031,N_1225,N_854);
xor U3032 (N_3032,N_55,N_565);
and U3033 (N_3033,N_2343,N_60);
xor U3034 (N_3034,N_1882,N_72);
and U3035 (N_3035,N_223,N_1036);
nand U3036 (N_3036,N_1484,N_121);
or U3037 (N_3037,N_731,N_2462);
nand U3038 (N_3038,N_1696,N_2315);
nand U3039 (N_3039,N_1291,N_1421);
nor U3040 (N_3040,N_1846,N_2236);
or U3041 (N_3041,N_2401,N_912);
or U3042 (N_3042,N_1293,N_2252);
nand U3043 (N_3043,N_1541,N_1249);
or U3044 (N_3044,N_725,N_200);
or U3045 (N_3045,N_841,N_1031);
nand U3046 (N_3046,N_1893,N_1318);
nand U3047 (N_3047,N_243,N_735);
nand U3048 (N_3048,N_318,N_2308);
and U3049 (N_3049,N_224,N_1819);
xnor U3050 (N_3050,N_2036,N_1677);
and U3051 (N_3051,N_966,N_1356);
or U3052 (N_3052,N_1128,N_1142);
xnor U3053 (N_3053,N_1348,N_690);
nor U3054 (N_3054,N_1115,N_1021);
or U3055 (N_3055,N_1052,N_564);
nor U3056 (N_3056,N_69,N_256);
nor U3057 (N_3057,N_2472,N_1355);
and U3058 (N_3058,N_2279,N_1180);
xnor U3059 (N_3059,N_1339,N_1773);
nand U3060 (N_3060,N_549,N_47);
and U3061 (N_3061,N_539,N_2344);
and U3062 (N_3062,N_1150,N_1668);
nand U3063 (N_3063,N_2436,N_1004);
or U3064 (N_3064,N_1425,N_2067);
or U3065 (N_3065,N_1221,N_413);
xnor U3066 (N_3066,N_2114,N_1957);
or U3067 (N_3067,N_417,N_436);
and U3068 (N_3068,N_143,N_2071);
and U3069 (N_3069,N_427,N_1012);
and U3070 (N_3070,N_511,N_1581);
and U3071 (N_3071,N_206,N_1409);
nor U3072 (N_3072,N_1322,N_67);
nor U3073 (N_3073,N_1570,N_632);
and U3074 (N_3074,N_1953,N_2374);
or U3075 (N_3075,N_1207,N_2191);
nand U3076 (N_3076,N_513,N_2113);
xnor U3077 (N_3077,N_273,N_1236);
or U3078 (N_3078,N_1256,N_1361);
and U3079 (N_3079,N_2257,N_1802);
and U3080 (N_3080,N_1010,N_620);
or U3081 (N_3081,N_985,N_1725);
nand U3082 (N_3082,N_1389,N_998);
nand U3083 (N_3083,N_131,N_1464);
nand U3084 (N_3084,N_1623,N_1626);
or U3085 (N_3085,N_684,N_2319);
nor U3086 (N_3086,N_1845,N_786);
nor U3087 (N_3087,N_902,N_1034);
and U3088 (N_3088,N_2275,N_231);
and U3089 (N_3089,N_2021,N_2058);
and U3090 (N_3090,N_361,N_1174);
nor U3091 (N_3091,N_251,N_650);
nand U3092 (N_3092,N_742,N_2415);
nand U3093 (N_3093,N_306,N_2285);
nand U3094 (N_3094,N_74,N_1859);
xor U3095 (N_3095,N_1908,N_880);
and U3096 (N_3096,N_1779,N_2497);
nor U3097 (N_3097,N_910,N_478);
or U3098 (N_3098,N_654,N_335);
nand U3099 (N_3099,N_1624,N_629);
nand U3100 (N_3100,N_2270,N_2063);
nor U3101 (N_3101,N_195,N_590);
nor U3102 (N_3102,N_606,N_1986);
and U3103 (N_3103,N_1238,N_2054);
nor U3104 (N_3104,N_865,N_2158);
nand U3105 (N_3105,N_409,N_2271);
or U3106 (N_3106,N_818,N_374);
nor U3107 (N_3107,N_1535,N_1340);
or U3108 (N_3108,N_883,N_1858);
or U3109 (N_3109,N_276,N_249);
and U3110 (N_3110,N_768,N_1516);
or U3111 (N_3111,N_869,N_1751);
nand U3112 (N_3112,N_1829,N_2366);
nand U3113 (N_3113,N_258,N_873);
or U3114 (N_3114,N_1438,N_589);
or U3115 (N_3115,N_2325,N_1208);
nand U3116 (N_3116,N_1205,N_1517);
xor U3117 (N_3117,N_1899,N_728);
or U3118 (N_3118,N_2171,N_283);
nand U3119 (N_3119,N_863,N_1364);
nand U3120 (N_3120,N_2336,N_1493);
nand U3121 (N_3121,N_738,N_1222);
and U3122 (N_3122,N_102,N_207);
and U3123 (N_3123,N_77,N_1554);
nand U3124 (N_3124,N_2475,N_1592);
and U3125 (N_3125,N_1486,N_1862);
xnor U3126 (N_3126,N_1536,N_1385);
nor U3127 (N_3127,N_2250,N_550);
and U3128 (N_3128,N_506,N_595);
or U3129 (N_3129,N_1457,N_682);
nand U3130 (N_3130,N_2302,N_1594);
nand U3131 (N_3131,N_1436,N_106);
nand U3132 (N_3132,N_2311,N_1655);
nor U3133 (N_3133,N_1444,N_519);
nor U3134 (N_3134,N_366,N_332);
and U3135 (N_3135,N_1873,N_2483);
and U3136 (N_3136,N_677,N_1195);
and U3137 (N_3137,N_2034,N_2359);
and U3138 (N_3138,N_1166,N_1359);
nand U3139 (N_3139,N_472,N_1363);
nor U3140 (N_3140,N_210,N_2268);
nor U3141 (N_3141,N_434,N_3);
nor U3142 (N_3142,N_816,N_2141);
and U3143 (N_3143,N_736,N_581);
and U3144 (N_3144,N_1825,N_1647);
nand U3145 (N_3145,N_2001,N_365);
and U3146 (N_3146,N_826,N_153);
and U3147 (N_3147,N_408,N_1401);
nor U3148 (N_3148,N_2223,N_1933);
xor U3149 (N_3149,N_301,N_1938);
nor U3150 (N_3150,N_814,N_2348);
nor U3151 (N_3151,N_1960,N_1137);
or U3152 (N_3152,N_1710,N_252);
and U3153 (N_3153,N_1792,N_1111);
and U3154 (N_3154,N_354,N_1503);
or U3155 (N_3155,N_2445,N_1608);
nand U3156 (N_3156,N_2432,N_2416);
and U3157 (N_3157,N_900,N_1983);
nor U3158 (N_3158,N_2363,N_740);
and U3159 (N_3159,N_1540,N_124);
nor U3160 (N_3160,N_1916,N_54);
nor U3161 (N_3161,N_1387,N_351);
or U3162 (N_3162,N_938,N_658);
and U3163 (N_3163,N_667,N_2093);
nand U3164 (N_3164,N_562,N_569);
and U3165 (N_3165,N_215,N_219);
or U3166 (N_3166,N_2466,N_2426);
nand U3167 (N_3167,N_2290,N_2169);
nor U3168 (N_3168,N_342,N_778);
nand U3169 (N_3169,N_1720,N_489);
and U3170 (N_3170,N_634,N_804);
nor U3171 (N_3171,N_20,N_1310);
nand U3172 (N_3172,N_1803,N_232);
and U3173 (N_3173,N_598,N_1537);
nand U3174 (N_3174,N_1030,N_2420);
nand U3175 (N_3175,N_2220,N_12);
or U3176 (N_3176,N_483,N_1211);
nand U3177 (N_3177,N_118,N_1884);
or U3178 (N_3178,N_1712,N_1458);
or U3179 (N_3179,N_810,N_2476);
nand U3180 (N_3180,N_430,N_349);
nor U3181 (N_3181,N_216,N_843);
and U3182 (N_3182,N_1880,N_2273);
and U3183 (N_3183,N_1805,N_2406);
nor U3184 (N_3184,N_732,N_254);
nor U3185 (N_3185,N_552,N_1429);
and U3186 (N_3186,N_282,N_2284);
and U3187 (N_3187,N_278,N_1229);
or U3188 (N_3188,N_1841,N_1254);
nor U3189 (N_3189,N_2402,N_2224);
xor U3190 (N_3190,N_19,N_485);
or U3191 (N_3191,N_1309,N_612);
nor U3192 (N_3192,N_2245,N_1824);
and U3193 (N_3193,N_991,N_1179);
nand U3194 (N_3194,N_624,N_2320);
nand U3195 (N_3195,N_2354,N_369);
nor U3196 (N_3196,N_1936,N_2389);
xnor U3197 (N_3197,N_371,N_1216);
nand U3198 (N_3198,N_1240,N_2087);
nor U3199 (N_3199,N_362,N_2151);
and U3200 (N_3200,N_675,N_904);
and U3201 (N_3201,N_1663,N_2068);
and U3202 (N_3202,N_541,N_1966);
or U3203 (N_3203,N_1708,N_2078);
and U3204 (N_3204,N_501,N_397);
nand U3205 (N_3205,N_1627,N_1152);
and U3206 (N_3206,N_1657,N_2145);
nor U3207 (N_3207,N_1628,N_2125);
xor U3208 (N_3208,N_1950,N_1000);
nand U3209 (N_3209,N_18,N_1694);
nand U3210 (N_3210,N_1875,N_2329);
nor U3211 (N_3211,N_1196,N_2310);
nand U3212 (N_3212,N_666,N_378);
or U3213 (N_3213,N_2109,N_615);
and U3214 (N_3214,N_2111,N_1182);
nor U3215 (N_3215,N_777,N_101);
or U3216 (N_3216,N_1838,N_189);
or U3217 (N_3217,N_2370,N_180);
and U3218 (N_3218,N_2246,N_976);
or U3219 (N_3219,N_1419,N_142);
nand U3220 (N_3220,N_617,N_130);
or U3221 (N_3221,N_1066,N_2442);
nor U3222 (N_3222,N_992,N_190);
nor U3223 (N_3223,N_2317,N_2342);
nand U3224 (N_3224,N_1237,N_138);
xor U3225 (N_3225,N_1637,N_1433);
nand U3226 (N_3226,N_642,N_2404);
nand U3227 (N_3227,N_1393,N_1056);
nor U3228 (N_3228,N_2350,N_1400);
nor U3229 (N_3229,N_309,N_1268);
or U3230 (N_3230,N_191,N_593);
or U3231 (N_3231,N_1900,N_432);
nor U3232 (N_3232,N_1583,N_2180);
or U3233 (N_3233,N_71,N_172);
and U3234 (N_3234,N_1970,N_6);
or U3235 (N_3235,N_1327,N_1140);
and U3236 (N_3236,N_891,N_1390);
nor U3237 (N_3237,N_1218,N_1507);
nand U3238 (N_3238,N_930,N_468);
nand U3239 (N_3239,N_104,N_2470);
and U3240 (N_3240,N_86,N_43);
nand U3241 (N_3241,N_2176,N_1867);
or U3242 (N_3242,N_2249,N_2237);
nand U3243 (N_3243,N_377,N_2447);
or U3244 (N_3244,N_1691,N_326);
and U3245 (N_3245,N_700,N_1753);
and U3246 (N_3246,N_1879,N_1341);
nand U3247 (N_3247,N_1149,N_137);
nor U3248 (N_3248,N_1070,N_1337);
nand U3249 (N_3249,N_715,N_496);
nand U3250 (N_3250,N_1317,N_1813);
nor U3251 (N_3251,N_11,N_2174);
or U3252 (N_3252,N_2206,N_265);
nand U3253 (N_3253,N_1255,N_1217);
xor U3254 (N_3254,N_1063,N_1093);
nor U3255 (N_3255,N_310,N_1281);
nand U3256 (N_3256,N_2488,N_245);
nor U3257 (N_3257,N_1713,N_2383);
or U3258 (N_3258,N_1978,N_451);
and U3259 (N_3259,N_578,N_685);
xor U3260 (N_3260,N_983,N_1353);
xor U3261 (N_3261,N_1886,N_1600);
nand U3262 (N_3262,N_772,N_1780);
and U3263 (N_3263,N_2277,N_40);
nor U3264 (N_3264,N_459,N_1072);
or U3265 (N_3265,N_194,N_2104);
nand U3266 (N_3266,N_1292,N_202);
nand U3267 (N_3267,N_95,N_931);
nand U3268 (N_3268,N_1439,N_2127);
or U3269 (N_3269,N_2122,N_1996);
and U3270 (N_3270,N_1499,N_1423);
or U3271 (N_3271,N_823,N_2421);
nor U3272 (N_3272,N_136,N_2465);
nand U3273 (N_3273,N_648,N_784);
nor U3274 (N_3274,N_2309,N_404);
nand U3275 (N_3275,N_925,N_1498);
or U3276 (N_3276,N_62,N_1676);
and U3277 (N_3277,N_1758,N_1406);
or U3278 (N_3278,N_460,N_1550);
or U3279 (N_3279,N_2299,N_1670);
or U3280 (N_3280,N_316,N_1735);
or U3281 (N_3281,N_1766,N_2126);
or U3282 (N_3282,N_285,N_995);
and U3283 (N_3283,N_1033,N_749);
nand U3284 (N_3284,N_1607,N_1926);
or U3285 (N_3285,N_2064,N_385);
nor U3286 (N_3286,N_673,N_26);
and U3287 (N_3287,N_2326,N_406);
or U3288 (N_3288,N_955,N_932);
or U3289 (N_3289,N_2080,N_2209);
nand U3290 (N_3290,N_746,N_514);
nor U3291 (N_3291,N_1215,N_1759);
nor U3292 (N_3292,N_1771,N_996);
or U3293 (N_3293,N_967,N_790);
and U3294 (N_3294,N_331,N_1723);
or U3295 (N_3295,N_644,N_31);
nor U3296 (N_3296,N_495,N_945);
and U3297 (N_3297,N_721,N_701);
or U3298 (N_3298,N_176,N_704);
nor U3299 (N_3299,N_2261,N_313);
nand U3300 (N_3300,N_621,N_1596);
or U3301 (N_3301,N_1861,N_1437);
or U3302 (N_3302,N_2131,N_2015);
nor U3303 (N_3303,N_1667,N_1119);
nand U3304 (N_3304,N_1703,N_1629);
or U3305 (N_3305,N_1417,N_493);
or U3306 (N_3306,N_1384,N_2491);
nor U3307 (N_3307,N_2003,N_1117);
or U3308 (N_3308,N_236,N_661);
and U3309 (N_3309,N_2490,N_275);
nand U3310 (N_3310,N_1514,N_2489);
nand U3311 (N_3311,N_203,N_2372);
nand U3312 (N_3312,N_1958,N_1870);
nor U3313 (N_3313,N_1206,N_1721);
nand U3314 (N_3314,N_2214,N_2238);
and U3315 (N_3315,N_1397,N_889);
nor U3316 (N_3316,N_1847,N_994);
nor U3317 (N_3317,N_1673,N_1878);
nand U3318 (N_3318,N_1272,N_663);
nor U3319 (N_3319,N_2446,N_113);
and U3320 (N_3320,N_1298,N_571);
nor U3321 (N_3321,N_670,N_346);
and U3322 (N_3322,N_1588,N_1350);
nand U3323 (N_3323,N_1821,N_319);
nor U3324 (N_3324,N_109,N_1365);
nand U3325 (N_3325,N_1815,N_2443);
nand U3326 (N_3326,N_773,N_2172);
nor U3327 (N_3327,N_1887,N_347);
nand U3328 (N_3328,N_588,N_355);
or U3329 (N_3329,N_1257,N_314);
nand U3330 (N_3330,N_720,N_2239);
nor U3331 (N_3331,N_1601,N_1496);
nor U3332 (N_3332,N_422,N_651);
xnor U3333 (N_3333,N_204,N_149);
or U3334 (N_3334,N_429,N_1586);
nand U3335 (N_3335,N_890,N_2139);
nand U3336 (N_3336,N_2499,N_2293);
or U3337 (N_3337,N_1299,N_1574);
or U3338 (N_3338,N_993,N_400);
nor U3339 (N_3339,N_1015,N_1087);
nand U3340 (N_3340,N_90,N_2012);
nor U3341 (N_3341,N_1265,N_1959);
nor U3342 (N_3342,N_837,N_652);
and U3343 (N_3343,N_1755,N_2460);
and U3344 (N_3344,N_241,N_613);
nor U3345 (N_3345,N_551,N_1346);
nor U3346 (N_3346,N_1094,N_1158);
nor U3347 (N_3347,N_1477,N_440);
nand U3348 (N_3348,N_542,N_418);
nand U3349 (N_3349,N_2207,N_745);
nand U3350 (N_3350,N_2165,N_1095);
nand U3351 (N_3351,N_187,N_2037);
nand U3352 (N_3352,N_403,N_2203);
or U3353 (N_3353,N_2390,N_1525);
or U3354 (N_3354,N_1086,N_490);
nand U3355 (N_3355,N_402,N_2192);
or U3356 (N_3356,N_942,N_544);
or U3357 (N_3357,N_2263,N_831);
or U3358 (N_3358,N_2391,N_2161);
nand U3359 (N_3359,N_2074,N_1618);
or U3360 (N_3360,N_416,N_2283);
or U3361 (N_3361,N_1358,N_1450);
or U3362 (N_3362,N_2190,N_1247);
or U3363 (N_3363,N_1998,N_1261);
nand U3364 (N_3364,N_317,N_2144);
nor U3365 (N_3365,N_2323,N_330);
nor U3366 (N_3366,N_1316,N_45);
nand U3367 (N_3367,N_2035,N_697);
or U3368 (N_3368,N_2102,N_553);
or U3369 (N_3369,N_1250,N_315);
or U3370 (N_3370,N_753,N_1252);
nor U3371 (N_3371,N_2479,N_803);
nor U3372 (N_3372,N_1489,N_1930);
nor U3373 (N_3373,N_2495,N_297);
and U3374 (N_3374,N_263,N_1684);
and U3375 (N_3375,N_1748,N_98);
nand U3376 (N_3376,N_461,N_1761);
nand U3377 (N_3377,N_128,N_1362);
nor U3378 (N_3378,N_127,N_1984);
and U3379 (N_3379,N_465,N_370);
and U3380 (N_3380,N_145,N_56);
nor U3381 (N_3381,N_1253,N_267);
and U3382 (N_3382,N_307,N_1301);
nand U3383 (N_3383,N_88,N_2147);
nand U3384 (N_3384,N_463,N_2347);
or U3385 (N_3385,N_1035,N_2008);
nor U3386 (N_3386,N_1897,N_2382);
nor U3387 (N_3387,N_798,N_2105);
nand U3388 (N_3388,N_1136,N_1501);
or U3389 (N_3389,N_2385,N_352);
nand U3390 (N_3390,N_13,N_1731);
nand U3391 (N_3391,N_2164,N_2133);
nor U3392 (N_3392,N_1114,N_2428);
xnor U3393 (N_3393,N_1774,N_954);
nor U3394 (N_3394,N_414,N_1367);
or U3395 (N_3395,N_2419,N_2380);
nand U3396 (N_3396,N_1539,N_1370);
nor U3397 (N_3397,N_1138,N_1976);
nor U3398 (N_3398,N_1528,N_1029);
and U3399 (N_3399,N_747,N_2457);
and U3400 (N_3400,N_168,N_1315);
nor U3401 (N_3401,N_1961,N_2269);
nand U3402 (N_3402,N_375,N_597);
or U3403 (N_3403,N_2056,N_296);
or U3404 (N_3404,N_1344,N_1658);
nor U3405 (N_3405,N_668,N_567);
and U3406 (N_3406,N_2322,N_235);
xor U3407 (N_3407,N_1410,N_1188);
nor U3408 (N_3408,N_1164,N_175);
and U3409 (N_3409,N_1597,N_1785);
nand U3410 (N_3410,N_2451,N_2484);
nor U3411 (N_3411,N_2168,N_1473);
xnor U3412 (N_3412,N_2365,N_586);
nor U3413 (N_3413,N_75,N_1106);
nand U3414 (N_3414,N_1577,N_486);
nor U3415 (N_3415,N_901,N_376);
and U3416 (N_3416,N_1837,N_1656);
nor U3417 (N_3417,N_2288,N_1038);
and U3418 (N_3418,N_2156,N_756);
and U3419 (N_3419,N_1264,N_1665);
nand U3420 (N_3420,N_1335,N_906);
nor U3421 (N_3421,N_1148,N_2265);
or U3422 (N_3422,N_1234,N_157);
nand U3423 (N_3423,N_50,N_97);
or U3424 (N_3424,N_1830,N_1582);
nand U3425 (N_3425,N_23,N_437);
nor U3426 (N_3426,N_2215,N_534);
and U3427 (N_3427,N_1989,N_2272);
nor U3428 (N_3428,N_199,N_943);
nor U3429 (N_3429,N_2204,N_1330);
nand U3430 (N_3430,N_1544,N_575);
nor U3431 (N_3431,N_903,N_1162);
and U3432 (N_3432,N_57,N_917);
nor U3433 (N_3433,N_2229,N_1209);
and U3434 (N_3434,N_1510,N_1191);
nand U3435 (N_3435,N_599,N_473);
nor U3436 (N_3436,N_1134,N_1352);
and U3437 (N_3437,N_209,N_561);
and U3438 (N_3438,N_1248,N_491);
nor U3439 (N_3439,N_1999,N_159);
xor U3440 (N_3440,N_537,N_2281);
nand U3441 (N_3441,N_396,N_1153);
and U3442 (N_3442,N_186,N_1512);
or U3443 (N_3443,N_879,N_1263);
or U3444 (N_3444,N_855,N_2181);
and U3445 (N_3445,N_706,N_1504);
nand U3446 (N_3446,N_886,N_1064);
nor U3447 (N_3447,N_2072,N_2201);
nand U3448 (N_3448,N_533,N_5);
or U3449 (N_3449,N_1811,N_115);
nor U3450 (N_3450,N_647,N_192);
nor U3451 (N_3451,N_1032,N_1674);
nand U3452 (N_3452,N_1077,N_929);
or U3453 (N_3453,N_1101,N_838);
or U3454 (N_3454,N_2381,N_2137);
xnor U3455 (N_3455,N_401,N_1262);
xnor U3456 (N_3456,N_2075,N_1968);
xnor U3457 (N_3457,N_1399,N_1187);
or U3458 (N_3458,N_2044,N_835);
nand U3459 (N_3459,N_834,N_1047);
and U3460 (N_3460,N_1561,N_2019);
or U3461 (N_3461,N_1947,N_1833);
and U3462 (N_3462,N_1267,N_1062);
nor U3463 (N_3463,N_2185,N_1680);
or U3464 (N_3464,N_1442,N_1160);
nand U3465 (N_3465,N_940,N_576);
nor U3466 (N_3466,N_2346,N_645);
and U3467 (N_3467,N_167,N_2010);
or U3468 (N_3468,N_2221,N_1943);
nor U3469 (N_3469,N_1790,N_2115);
nor U3470 (N_3470,N_2097,N_2159);
nand U3471 (N_3471,N_323,N_1283);
and U3472 (N_3472,N_1866,N_678);
and U3473 (N_3473,N_1045,N_255);
nand U3474 (N_3474,N_2119,N_510);
nand U3475 (N_3475,N_2052,N_1053);
nor U3476 (N_3476,N_2173,N_981);
xor U3477 (N_3477,N_1855,N_935);
nand U3478 (N_3478,N_2222,N_1235);
and U3479 (N_3479,N_1284,N_2330);
nand U3480 (N_3480,N_2286,N_947);
or U3481 (N_3481,N_2304,N_2062);
and U3482 (N_3482,N_2274,N_1944);
or U3483 (N_3483,N_225,N_329);
nor U3484 (N_3484,N_1889,N_2143);
or U3485 (N_3485,N_1538,N_294);
and U3486 (N_3486,N_2154,N_2339);
or U3487 (N_3487,N_1876,N_1630);
nor U3488 (N_3488,N_2178,N_2423);
or U3489 (N_3489,N_1300,N_1170);
nand U3490 (N_3490,N_2376,N_762);
nand U3491 (N_3491,N_185,N_266);
nor U3492 (N_3492,N_605,N_1443);
nor U3493 (N_3493,N_150,N_1973);
nand U3494 (N_3494,N_304,N_1800);
nor U3495 (N_3495,N_845,N_171);
and U3496 (N_3496,N_1483,N_1104);
and U3497 (N_3497,N_274,N_1625);
and U3498 (N_3498,N_1303,N_1924);
and U3499 (N_3499,N_572,N_68);
xor U3500 (N_3500,N_696,N_1609);
nor U3501 (N_3501,N_286,N_248);
or U3502 (N_3502,N_1891,N_2177);
nor U3503 (N_3503,N_144,N_24);
nor U3504 (N_3504,N_2241,N_2002);
or U3505 (N_3505,N_888,N_1186);
nand U3506 (N_3506,N_619,N_1534);
and U3507 (N_3507,N_2208,N_357);
or U3508 (N_3508,N_1814,N_987);
nor U3509 (N_3509,N_856,N_1100);
or U3510 (N_3510,N_462,N_1651);
nor U3511 (N_3511,N_1781,N_1026);
nand U3512 (N_3512,N_284,N_1981);
nand U3513 (N_3513,N_246,N_1411);
nor U3514 (N_3514,N_1687,N_515);
xnor U3515 (N_3515,N_2371,N_179);
and U3516 (N_3516,N_2297,N_2414);
nor U3517 (N_3517,N_2332,N_1728);
nand U3518 (N_3518,N_828,N_169);
or U3519 (N_3519,N_1902,N_360);
nand U3520 (N_3520,N_439,N_1616);
nor U3521 (N_3521,N_1147,N_320);
or U3522 (N_3522,N_2076,N_870);
nand U3523 (N_3523,N_358,N_764);
nand U3524 (N_3524,N_279,N_1177);
and U3525 (N_3525,N_859,N_340);
nand U3526 (N_3526,N_1700,N_1760);
or U3527 (N_3527,N_2200,N_2);
nor U3528 (N_3528,N_499,N_220);
nor U3529 (N_3529,N_21,N_65);
or U3530 (N_3530,N_1491,N_2077);
nand U3531 (N_3531,N_1727,N_1689);
nor U3532 (N_3532,N_1159,N_1942);
nor U3533 (N_3533,N_1826,N_664);
nand U3534 (N_3534,N_15,N_188);
nor U3535 (N_3535,N_1804,N_2395);
nor U3536 (N_3536,N_655,N_240);
nor U3537 (N_3537,N_1075,N_129);
nand U3538 (N_3538,N_1424,N_965);
and U3539 (N_3539,N_1881,N_458);
nor U3540 (N_3540,N_1646,N_27);
and U3541 (N_3541,N_2334,N_2478);
or U3542 (N_3542,N_898,N_79);
and U3543 (N_3543,N_2452,N_341);
nor U3544 (N_3544,N_1024,N_972);
nor U3545 (N_3545,N_2362,N_671);
nand U3546 (N_3546,N_16,N_498);
nor U3547 (N_3547,N_1373,N_726);
or U3548 (N_3548,N_2148,N_1744);
nor U3549 (N_3549,N_1434,N_1448);
or U3550 (N_3550,N_1764,N_1992);
or U3551 (N_3551,N_1058,N_545);
xnor U3552 (N_3552,N_2112,N_2411);
and U3553 (N_3553,N_1515,N_1831);
nand U3554 (N_3554,N_693,N_1127);
or U3555 (N_3555,N_2424,N_2059);
and U3556 (N_3556,N_2150,N_1649);
nand U3557 (N_3557,N_1242,N_637);
or U3558 (N_3558,N_1745,N_2193);
or U3559 (N_3559,N_2410,N_83);
and U3560 (N_3560,N_676,N_1797);
nor U3561 (N_3561,N_1851,N_1369);
nor U3562 (N_3562,N_325,N_2412);
and U3563 (N_3563,N_1645,N_807);
and U3564 (N_3564,N_2399,N_76);
or U3565 (N_3565,N_338,N_2079);
nand U3566 (N_3566,N_497,N_2146);
nand U3567 (N_3567,N_264,N_892);
and U3568 (N_3568,N_1328,N_871);
nand U3569 (N_3569,N_1374,N_2100);
and U3570 (N_3570,N_126,N_848);
or U3571 (N_3571,N_96,N_2434);
nand U3572 (N_3572,N_953,N_1714);
and U3573 (N_3573,N_2000,N_769);
or U3574 (N_3574,N_1852,N_1571);
nor U3575 (N_3575,N_952,N_1784);
nand U3576 (N_3576,N_303,N_492);
nand U3577 (N_3577,N_751,N_842);
xor U3578 (N_3578,N_1686,N_723);
or U3579 (N_3579,N_2298,N_951);
nor U3580 (N_3580,N_1523,N_1509);
and U3581 (N_3581,N_1091,N_1109);
and U3582 (N_3582,N_93,N_237);
nand U3583 (N_3583,N_372,N_1559);
and U3584 (N_3584,N_1500,N_1002);
nand U3585 (N_3585,N_2218,N_1474);
or U3586 (N_3586,N_1061,N_2364);
and U3587 (N_3587,N_1641,N_809);
and U3588 (N_3588,N_2289,N_1274);
and U3589 (N_3589,N_428,N_395);
nor U3590 (N_3590,N_2313,N_213);
xnor U3591 (N_3591,N_2130,N_1282);
nor U3592 (N_3592,N_1366,N_1005);
nor U3593 (N_3593,N_405,N_1122);
or U3594 (N_3594,N_2264,N_2196);
nand U3595 (N_3595,N_1060,N_1595);
and U3596 (N_3596,N_861,N_1575);
or U3597 (N_3597,N_53,N_1204);
and U3598 (N_3598,N_1948,N_1567);
nor U3599 (N_3599,N_913,N_528);
nand U3600 (N_3600,N_1266,N_2083);
or U3601 (N_3601,N_583,N_867);
and U3602 (N_3602,N_1569,N_1067);
nor U3603 (N_3603,N_1173,N_132);
nor U3604 (N_3604,N_2051,N_1823);
or U3605 (N_3605,N_881,N_674);
nand U3606 (N_3606,N_1481,N_556);
nand U3607 (N_3607,N_2157,N_882);
or U3608 (N_3608,N_1492,N_2429);
and U3609 (N_3609,N_1485,N_269);
and U3610 (N_3610,N_792,N_328);
or U3611 (N_3611,N_2198,N_1722);
and U3612 (N_3612,N_212,N_1810);
and U3613 (N_3613,N_1228,N_1057);
nor U3614 (N_3614,N_2184,N_1705);
nor U3615 (N_3615,N_603,N_1304);
nor U3616 (N_3616,N_771,N_775);
and U3617 (N_3617,N_672,N_1001);
nand U3618 (N_3618,N_1311,N_1307);
or U3619 (N_3619,N_1018,N_38);
or U3620 (N_3620,N_1707,N_1230);
xnor U3621 (N_3621,N_653,N_1382);
and U3622 (N_3622,N_1985,N_1200);
or U3623 (N_3623,N_222,N_1791);
nor U3624 (N_3624,N_687,N_164);
and U3625 (N_3625,N_1602,N_812);
nand U3626 (N_3626,N_585,N_958);
nor U3627 (N_3627,N_530,N_1698);
and U3628 (N_3628,N_1381,N_1812);
or U3629 (N_3629,N_1817,N_752);
and U3630 (N_3630,N_399,N_343);
nor U3631 (N_3631,N_2026,N_1949);
nand U3632 (N_3632,N_1394,N_536);
and U3633 (N_3633,N_2152,N_543);
nand U3634 (N_3634,N_2254,N_2482);
xor U3635 (N_3635,N_1990,N_2292);
and U3636 (N_3636,N_1642,N_1954);
or U3637 (N_3637,N_456,N_669);
and U3638 (N_3638,N_1770,N_1023);
nand U3639 (N_3639,N_1197,N_466);
and U3640 (N_3640,N_1726,N_353);
or U3641 (N_3641,N_1598,N_239);
nand U3642 (N_3642,N_1116,N_563);
and U3643 (N_3643,N_2377,N_1508);
and U3644 (N_3644,N_2070,N_1558);
and U3645 (N_3645,N_2300,N_1456);
or U3646 (N_3646,N_602,N_141);
or U3647 (N_3647,N_1172,N_1145);
and U3648 (N_3648,N_2438,N_864);
nor U3649 (N_3649,N_1,N_419);
nor U3650 (N_3650,N_1648,N_1006);
and U3651 (N_3651,N_2098,N_1612);
nand U3652 (N_3652,N_2120,N_2013);
or U3653 (N_3653,N_1467,N_1584);
nand U3654 (N_3654,N_2233,N_1125);
or U3655 (N_3655,N_765,N_2085);
or U3656 (N_3656,N_783,N_2055);
nor U3657 (N_3657,N_1202,N_1699);
nand U3658 (N_3658,N_364,N_1321);
or U3659 (N_3659,N_1495,N_656);
and U3660 (N_3660,N_48,N_431);
or U3661 (N_3661,N_33,N_524);
nand U3662 (N_3662,N_1543,N_1319);
or U3663 (N_3663,N_640,N_32);
and U3664 (N_3664,N_1603,N_635);
or U3665 (N_3665,N_1513,N_707);
and U3666 (N_3666,N_1576,N_1378);
and U3667 (N_3667,N_470,N_1750);
nor U3668 (N_3668,N_1573,N_389);
nor U3669 (N_3669,N_1964,N_1308);
and U3670 (N_3670,N_1632,N_990);
or U3671 (N_3671,N_292,N_582);
or U3672 (N_3672,N_218,N_822);
nor U3673 (N_3673,N_2235,N_2069);
or U3674 (N_3674,N_155,N_1280);
and U3675 (N_3675,N_2469,N_2444);
nor U3676 (N_3676,N_1666,N_1462);
nand U3677 (N_3677,N_2314,N_1480);
and U3678 (N_3678,N_2091,N_1097);
and U3679 (N_3679,N_1702,N_2023);
nor U3680 (N_3680,N_516,N_1865);
or U3681 (N_3681,N_193,N_2153);
nor U3682 (N_3682,N_2022,N_333);
nor U3683 (N_3683,N_467,N_1156);
nand U3684 (N_3684,N_1079,N_1088);
nand U3685 (N_3685,N_1141,N_2149);
and U3686 (N_3686,N_614,N_2367);
and U3687 (N_3687,N_1407,N_1306);
nor U3688 (N_3688,N_476,N_2230);
nor U3689 (N_3689,N_441,N_28);
nand U3690 (N_3690,N_2226,N_639);
nand U3691 (N_3691,N_763,N_2260);
or U3692 (N_3692,N_1551,N_538);
and U3693 (N_3693,N_177,N_1898);
nor U3694 (N_3694,N_554,N_2116);
or U3695 (N_3695,N_1377,N_594);
or U3696 (N_3696,N_2251,N_1224);
and U3697 (N_3697,N_824,N_934);
and U3698 (N_3698,N_928,N_761);
xor U3699 (N_3699,N_1956,N_1552);
or U3700 (N_3700,N_811,N_1888);
or U3701 (N_3701,N_1354,N_94);
or U3702 (N_3702,N_1742,N_41);
or U3703 (N_3703,N_2025,N_2324);
nand U3704 (N_3704,N_1245,N_579);
nor U3705 (N_3705,N_1019,N_1331);
and U3706 (N_3706,N_1447,N_117);
and U3707 (N_3707,N_37,N_743);
nor U3708 (N_3708,N_2135,N_948);
or U3709 (N_3709,N_517,N_260);
nor U3710 (N_3710,N_312,N_918);
or U3711 (N_3711,N_1161,N_2107);
nand U3712 (N_3712,N_1312,N_1711);
and U3713 (N_3713,N_716,N_2155);
or U3714 (N_3714,N_2455,N_398);
nand U3715 (N_3715,N_299,N_1044);
nand U3716 (N_3716,N_1530,N_381);
and U3717 (N_3717,N_433,N_2094);
and U3718 (N_3718,N_1729,N_608);
and U3719 (N_3719,N_1465,N_1901);
and U3720 (N_3720,N_271,N_1243);
nor U3721 (N_3721,N_520,N_244);
nor U3722 (N_3722,N_2186,N_1338);
nor U3723 (N_3723,N_797,N_49);
nand U3724 (N_3724,N_2014,N_1347);
and U3725 (N_3725,N_2103,N_107);
nand U3726 (N_3726,N_46,N_688);
or U3727 (N_3727,N_607,N_2398);
nor U3728 (N_3728,N_66,N_393);
nand U3729 (N_3729,N_1404,N_729);
or U3730 (N_3730,N_36,N_800);
nor U3731 (N_3731,N_584,N_1226);
nor U3732 (N_3732,N_2464,N_363);
nor U3733 (N_3733,N_964,N_801);
or U3734 (N_3734,N_1654,N_2427);
and U3735 (N_3735,N_2496,N_1644);
nand U3736 (N_3736,N_592,N_2049);
nand U3737 (N_3737,N_2327,N_527);
or U3738 (N_3738,N_1737,N_1896);
and U3739 (N_3739,N_148,N_51);
nor U3740 (N_3740,N_944,N_875);
and U3741 (N_3741,N_2267,N_1470);
and U3742 (N_3742,N_52,N_916);
nor U3743 (N_3743,N_123,N_1043);
or U3744 (N_3744,N_1435,N_1885);
or U3745 (N_3745,N_1620,N_302);
or U3746 (N_3746,N_2040,N_1118);
nand U3747 (N_3747,N_2312,N_201);
nand U3748 (N_3748,N_122,N_469);
and U3749 (N_3749,N_920,N_1466);
nor U3750 (N_3750,N_2003,N_433);
and U3751 (N_3751,N_776,N_1548);
and U3752 (N_3752,N_1691,N_2465);
nand U3753 (N_3753,N_2129,N_1759);
and U3754 (N_3754,N_685,N_841);
nor U3755 (N_3755,N_1848,N_1486);
nand U3756 (N_3756,N_2386,N_1481);
and U3757 (N_3757,N_1715,N_828);
and U3758 (N_3758,N_1149,N_2352);
nand U3759 (N_3759,N_2099,N_2367);
and U3760 (N_3760,N_1463,N_843);
or U3761 (N_3761,N_1568,N_1005);
and U3762 (N_3762,N_2313,N_2109);
or U3763 (N_3763,N_474,N_2209);
nand U3764 (N_3764,N_2416,N_1853);
nor U3765 (N_3765,N_1780,N_920);
nand U3766 (N_3766,N_1281,N_1659);
or U3767 (N_3767,N_862,N_705);
and U3768 (N_3768,N_346,N_1321);
nand U3769 (N_3769,N_909,N_1966);
nor U3770 (N_3770,N_1148,N_1934);
nor U3771 (N_3771,N_1778,N_165);
or U3772 (N_3772,N_1157,N_178);
or U3773 (N_3773,N_796,N_1857);
and U3774 (N_3774,N_2384,N_1938);
and U3775 (N_3775,N_438,N_2250);
nor U3776 (N_3776,N_1712,N_330);
nor U3777 (N_3777,N_316,N_801);
nor U3778 (N_3778,N_758,N_1335);
nand U3779 (N_3779,N_499,N_2200);
and U3780 (N_3780,N_641,N_2264);
nor U3781 (N_3781,N_2431,N_674);
or U3782 (N_3782,N_1789,N_290);
and U3783 (N_3783,N_1317,N_1309);
and U3784 (N_3784,N_1188,N_214);
and U3785 (N_3785,N_1202,N_487);
xor U3786 (N_3786,N_2184,N_919);
or U3787 (N_3787,N_864,N_1324);
or U3788 (N_3788,N_781,N_624);
and U3789 (N_3789,N_2310,N_507);
nor U3790 (N_3790,N_400,N_1858);
and U3791 (N_3791,N_1539,N_1610);
nor U3792 (N_3792,N_331,N_432);
nor U3793 (N_3793,N_627,N_83);
and U3794 (N_3794,N_2491,N_2475);
or U3795 (N_3795,N_585,N_1657);
nand U3796 (N_3796,N_2413,N_1620);
or U3797 (N_3797,N_1344,N_1191);
or U3798 (N_3798,N_2404,N_1649);
and U3799 (N_3799,N_1686,N_1701);
or U3800 (N_3800,N_171,N_16);
nor U3801 (N_3801,N_339,N_1631);
and U3802 (N_3802,N_365,N_1730);
nand U3803 (N_3803,N_1845,N_507);
nand U3804 (N_3804,N_1679,N_1219);
and U3805 (N_3805,N_619,N_360);
and U3806 (N_3806,N_1847,N_698);
nor U3807 (N_3807,N_1196,N_2365);
or U3808 (N_3808,N_1120,N_1356);
nor U3809 (N_3809,N_751,N_862);
and U3810 (N_3810,N_1824,N_59);
or U3811 (N_3811,N_358,N_570);
or U3812 (N_3812,N_303,N_315);
xnor U3813 (N_3813,N_1661,N_2267);
and U3814 (N_3814,N_2294,N_47);
nor U3815 (N_3815,N_1001,N_1551);
nor U3816 (N_3816,N_1132,N_2228);
and U3817 (N_3817,N_2089,N_2371);
or U3818 (N_3818,N_528,N_927);
nor U3819 (N_3819,N_1775,N_367);
nor U3820 (N_3820,N_1918,N_88);
nand U3821 (N_3821,N_1211,N_1452);
nor U3822 (N_3822,N_1509,N_1093);
nand U3823 (N_3823,N_1688,N_768);
nor U3824 (N_3824,N_497,N_1974);
nor U3825 (N_3825,N_1856,N_1814);
nand U3826 (N_3826,N_2486,N_1387);
nor U3827 (N_3827,N_1969,N_1729);
nand U3828 (N_3828,N_1076,N_2196);
and U3829 (N_3829,N_447,N_247);
nand U3830 (N_3830,N_2452,N_2214);
and U3831 (N_3831,N_1485,N_1607);
or U3832 (N_3832,N_2456,N_1254);
or U3833 (N_3833,N_2059,N_179);
or U3834 (N_3834,N_1392,N_293);
nor U3835 (N_3835,N_568,N_1151);
or U3836 (N_3836,N_1585,N_119);
nor U3837 (N_3837,N_704,N_253);
and U3838 (N_3838,N_1477,N_1436);
nand U3839 (N_3839,N_1883,N_881);
nand U3840 (N_3840,N_1977,N_176);
and U3841 (N_3841,N_946,N_1687);
or U3842 (N_3842,N_1791,N_1691);
and U3843 (N_3843,N_1357,N_872);
nand U3844 (N_3844,N_2275,N_989);
or U3845 (N_3845,N_1371,N_1383);
and U3846 (N_3846,N_1206,N_1456);
nand U3847 (N_3847,N_508,N_1015);
nand U3848 (N_3848,N_1729,N_1242);
nor U3849 (N_3849,N_2483,N_1329);
or U3850 (N_3850,N_499,N_1392);
and U3851 (N_3851,N_1445,N_2389);
nand U3852 (N_3852,N_379,N_2233);
nor U3853 (N_3853,N_1487,N_1557);
nor U3854 (N_3854,N_230,N_1873);
xor U3855 (N_3855,N_323,N_45);
or U3856 (N_3856,N_692,N_1481);
or U3857 (N_3857,N_1053,N_2216);
or U3858 (N_3858,N_1975,N_1810);
nand U3859 (N_3859,N_1356,N_1324);
nand U3860 (N_3860,N_1093,N_1297);
nand U3861 (N_3861,N_208,N_1549);
nand U3862 (N_3862,N_256,N_74);
or U3863 (N_3863,N_850,N_984);
and U3864 (N_3864,N_2031,N_96);
or U3865 (N_3865,N_241,N_2279);
and U3866 (N_3866,N_2271,N_144);
or U3867 (N_3867,N_1358,N_853);
and U3868 (N_3868,N_1724,N_1602);
nor U3869 (N_3869,N_2284,N_348);
nand U3870 (N_3870,N_1784,N_2433);
nor U3871 (N_3871,N_2474,N_2064);
nand U3872 (N_3872,N_998,N_1745);
nand U3873 (N_3873,N_1869,N_789);
or U3874 (N_3874,N_1518,N_342);
or U3875 (N_3875,N_1494,N_1674);
or U3876 (N_3876,N_819,N_49);
nor U3877 (N_3877,N_445,N_738);
and U3878 (N_3878,N_742,N_1346);
and U3879 (N_3879,N_2349,N_1688);
and U3880 (N_3880,N_1503,N_2304);
nor U3881 (N_3881,N_356,N_1490);
or U3882 (N_3882,N_507,N_2419);
or U3883 (N_3883,N_2046,N_2377);
nor U3884 (N_3884,N_2444,N_2331);
or U3885 (N_3885,N_954,N_634);
nor U3886 (N_3886,N_302,N_1238);
nor U3887 (N_3887,N_1023,N_1697);
or U3888 (N_3888,N_733,N_1406);
nand U3889 (N_3889,N_2224,N_1776);
and U3890 (N_3890,N_2226,N_698);
nand U3891 (N_3891,N_1370,N_1500);
xnor U3892 (N_3892,N_2105,N_1000);
or U3893 (N_3893,N_2486,N_127);
and U3894 (N_3894,N_643,N_2197);
and U3895 (N_3895,N_313,N_1234);
nand U3896 (N_3896,N_2446,N_574);
and U3897 (N_3897,N_1008,N_359);
and U3898 (N_3898,N_2351,N_2083);
nor U3899 (N_3899,N_1455,N_1465);
nor U3900 (N_3900,N_2485,N_1119);
or U3901 (N_3901,N_986,N_245);
nand U3902 (N_3902,N_791,N_1271);
nor U3903 (N_3903,N_1614,N_582);
nor U3904 (N_3904,N_2027,N_448);
nand U3905 (N_3905,N_1227,N_2093);
and U3906 (N_3906,N_1825,N_2046);
xnor U3907 (N_3907,N_2104,N_110);
or U3908 (N_3908,N_153,N_2049);
and U3909 (N_3909,N_1322,N_109);
and U3910 (N_3910,N_318,N_1278);
nand U3911 (N_3911,N_1342,N_249);
and U3912 (N_3912,N_572,N_2181);
nand U3913 (N_3913,N_860,N_1062);
and U3914 (N_3914,N_2008,N_741);
nand U3915 (N_3915,N_730,N_120);
or U3916 (N_3916,N_2159,N_2064);
nor U3917 (N_3917,N_2146,N_1846);
and U3918 (N_3918,N_2206,N_2226);
nand U3919 (N_3919,N_417,N_2316);
nand U3920 (N_3920,N_1083,N_2);
nor U3921 (N_3921,N_1391,N_912);
nor U3922 (N_3922,N_72,N_482);
or U3923 (N_3923,N_721,N_1961);
and U3924 (N_3924,N_1610,N_2181);
or U3925 (N_3925,N_1922,N_1483);
nand U3926 (N_3926,N_71,N_1942);
xnor U3927 (N_3927,N_1825,N_2424);
and U3928 (N_3928,N_1387,N_2017);
or U3929 (N_3929,N_1861,N_107);
nand U3930 (N_3930,N_687,N_1598);
or U3931 (N_3931,N_1414,N_1293);
or U3932 (N_3932,N_1202,N_199);
and U3933 (N_3933,N_1645,N_2330);
nor U3934 (N_3934,N_581,N_1764);
and U3935 (N_3935,N_933,N_201);
and U3936 (N_3936,N_633,N_546);
nand U3937 (N_3937,N_762,N_211);
nand U3938 (N_3938,N_950,N_1097);
or U3939 (N_3939,N_1683,N_2130);
and U3940 (N_3940,N_1138,N_987);
nand U3941 (N_3941,N_1752,N_2407);
and U3942 (N_3942,N_1126,N_83);
or U3943 (N_3943,N_1084,N_1887);
nand U3944 (N_3944,N_1126,N_2021);
nand U3945 (N_3945,N_1646,N_1358);
nand U3946 (N_3946,N_2042,N_37);
nand U3947 (N_3947,N_95,N_2070);
nor U3948 (N_3948,N_1325,N_846);
or U3949 (N_3949,N_2359,N_2157);
and U3950 (N_3950,N_1841,N_844);
nand U3951 (N_3951,N_9,N_2061);
or U3952 (N_3952,N_557,N_2178);
nor U3953 (N_3953,N_421,N_2187);
or U3954 (N_3954,N_100,N_690);
and U3955 (N_3955,N_119,N_797);
nor U3956 (N_3956,N_1279,N_69);
nor U3957 (N_3957,N_1311,N_1874);
nor U3958 (N_3958,N_655,N_271);
nand U3959 (N_3959,N_372,N_1499);
nand U3960 (N_3960,N_1848,N_2057);
nand U3961 (N_3961,N_416,N_291);
and U3962 (N_3962,N_718,N_1898);
nand U3963 (N_3963,N_2181,N_1739);
and U3964 (N_3964,N_2054,N_767);
or U3965 (N_3965,N_303,N_1273);
nand U3966 (N_3966,N_2068,N_2348);
and U3967 (N_3967,N_854,N_1060);
nand U3968 (N_3968,N_1938,N_2364);
or U3969 (N_3969,N_613,N_2497);
and U3970 (N_3970,N_78,N_869);
nand U3971 (N_3971,N_971,N_2098);
and U3972 (N_3972,N_1651,N_1509);
nand U3973 (N_3973,N_1616,N_1562);
nand U3974 (N_3974,N_522,N_2158);
nand U3975 (N_3975,N_300,N_2235);
nand U3976 (N_3976,N_2155,N_141);
and U3977 (N_3977,N_2132,N_872);
nor U3978 (N_3978,N_2255,N_1797);
nor U3979 (N_3979,N_398,N_1411);
or U3980 (N_3980,N_2372,N_2101);
or U3981 (N_3981,N_691,N_903);
and U3982 (N_3982,N_1654,N_468);
or U3983 (N_3983,N_1005,N_320);
or U3984 (N_3984,N_888,N_850);
nor U3985 (N_3985,N_2458,N_1262);
nand U3986 (N_3986,N_32,N_746);
or U3987 (N_3987,N_867,N_2345);
or U3988 (N_3988,N_1526,N_944);
nand U3989 (N_3989,N_1359,N_2268);
nor U3990 (N_3990,N_165,N_2085);
and U3991 (N_3991,N_542,N_2492);
nor U3992 (N_3992,N_334,N_261);
or U3993 (N_3993,N_2453,N_805);
nand U3994 (N_3994,N_2379,N_2203);
nor U3995 (N_3995,N_1374,N_424);
nand U3996 (N_3996,N_2396,N_806);
nor U3997 (N_3997,N_471,N_211);
or U3998 (N_3998,N_1946,N_2431);
nand U3999 (N_3999,N_535,N_1381);
or U4000 (N_4000,N_1922,N_725);
or U4001 (N_4001,N_1196,N_1862);
nand U4002 (N_4002,N_1757,N_1476);
nand U4003 (N_4003,N_1816,N_850);
nand U4004 (N_4004,N_2091,N_677);
and U4005 (N_4005,N_2282,N_1865);
nor U4006 (N_4006,N_391,N_2062);
nand U4007 (N_4007,N_1761,N_1572);
or U4008 (N_4008,N_217,N_2123);
nand U4009 (N_4009,N_758,N_328);
nor U4010 (N_4010,N_2113,N_2311);
or U4011 (N_4011,N_908,N_2006);
nor U4012 (N_4012,N_444,N_818);
nor U4013 (N_4013,N_415,N_1402);
or U4014 (N_4014,N_642,N_2173);
nor U4015 (N_4015,N_812,N_9);
and U4016 (N_4016,N_948,N_319);
nand U4017 (N_4017,N_2396,N_658);
nor U4018 (N_4018,N_643,N_364);
nor U4019 (N_4019,N_709,N_678);
or U4020 (N_4020,N_2184,N_1965);
and U4021 (N_4021,N_90,N_1276);
or U4022 (N_4022,N_1442,N_591);
nor U4023 (N_4023,N_393,N_676);
and U4024 (N_4024,N_944,N_1157);
and U4025 (N_4025,N_1706,N_554);
nor U4026 (N_4026,N_837,N_1897);
nor U4027 (N_4027,N_773,N_391);
and U4028 (N_4028,N_1968,N_295);
or U4029 (N_4029,N_887,N_317);
and U4030 (N_4030,N_139,N_702);
or U4031 (N_4031,N_1352,N_2413);
and U4032 (N_4032,N_3,N_725);
nor U4033 (N_4033,N_2403,N_953);
nor U4034 (N_4034,N_748,N_1032);
xnor U4035 (N_4035,N_53,N_1470);
nand U4036 (N_4036,N_1010,N_1135);
nor U4037 (N_4037,N_1061,N_2214);
or U4038 (N_4038,N_1604,N_225);
nor U4039 (N_4039,N_2424,N_1387);
and U4040 (N_4040,N_1796,N_1026);
nor U4041 (N_4041,N_300,N_1312);
or U4042 (N_4042,N_229,N_46);
and U4043 (N_4043,N_2047,N_1547);
nand U4044 (N_4044,N_2065,N_558);
and U4045 (N_4045,N_2196,N_1849);
nor U4046 (N_4046,N_791,N_2331);
and U4047 (N_4047,N_1848,N_996);
or U4048 (N_4048,N_1352,N_1372);
nand U4049 (N_4049,N_589,N_867);
and U4050 (N_4050,N_1284,N_235);
or U4051 (N_4051,N_39,N_199);
or U4052 (N_4052,N_982,N_1968);
or U4053 (N_4053,N_2155,N_2012);
nor U4054 (N_4054,N_1381,N_2305);
nand U4055 (N_4055,N_1030,N_2240);
nor U4056 (N_4056,N_1891,N_1852);
or U4057 (N_4057,N_711,N_1265);
nand U4058 (N_4058,N_1914,N_1989);
nor U4059 (N_4059,N_1464,N_1344);
and U4060 (N_4060,N_251,N_532);
nand U4061 (N_4061,N_616,N_1741);
or U4062 (N_4062,N_1838,N_903);
or U4063 (N_4063,N_110,N_127);
or U4064 (N_4064,N_794,N_284);
and U4065 (N_4065,N_1322,N_909);
nand U4066 (N_4066,N_358,N_643);
xnor U4067 (N_4067,N_68,N_904);
and U4068 (N_4068,N_1627,N_933);
and U4069 (N_4069,N_281,N_661);
and U4070 (N_4070,N_1564,N_2268);
or U4071 (N_4071,N_1684,N_503);
and U4072 (N_4072,N_1771,N_216);
nor U4073 (N_4073,N_808,N_2464);
xor U4074 (N_4074,N_1378,N_160);
and U4075 (N_4075,N_1440,N_2410);
nor U4076 (N_4076,N_1140,N_867);
and U4077 (N_4077,N_195,N_885);
or U4078 (N_4078,N_1170,N_874);
xnor U4079 (N_4079,N_985,N_770);
nor U4080 (N_4080,N_1015,N_1985);
nand U4081 (N_4081,N_2238,N_848);
nand U4082 (N_4082,N_1714,N_1118);
and U4083 (N_4083,N_1877,N_2123);
nor U4084 (N_4084,N_1442,N_416);
nand U4085 (N_4085,N_1747,N_1646);
nor U4086 (N_4086,N_1706,N_1695);
nor U4087 (N_4087,N_2353,N_2259);
nand U4088 (N_4088,N_720,N_2171);
and U4089 (N_4089,N_987,N_1939);
and U4090 (N_4090,N_819,N_1130);
xor U4091 (N_4091,N_1297,N_1539);
nor U4092 (N_4092,N_1381,N_1077);
and U4093 (N_4093,N_647,N_2294);
nand U4094 (N_4094,N_1754,N_677);
and U4095 (N_4095,N_1462,N_147);
nor U4096 (N_4096,N_184,N_963);
or U4097 (N_4097,N_1214,N_840);
nor U4098 (N_4098,N_2203,N_2316);
and U4099 (N_4099,N_1527,N_1197);
and U4100 (N_4100,N_535,N_751);
and U4101 (N_4101,N_1065,N_75);
and U4102 (N_4102,N_2175,N_553);
or U4103 (N_4103,N_1568,N_1908);
nor U4104 (N_4104,N_528,N_1338);
and U4105 (N_4105,N_216,N_1145);
nor U4106 (N_4106,N_1179,N_2462);
or U4107 (N_4107,N_1856,N_2265);
or U4108 (N_4108,N_1630,N_1540);
or U4109 (N_4109,N_770,N_1630);
nand U4110 (N_4110,N_1055,N_882);
and U4111 (N_4111,N_8,N_1382);
and U4112 (N_4112,N_86,N_2036);
or U4113 (N_4113,N_1432,N_1821);
nand U4114 (N_4114,N_2150,N_145);
or U4115 (N_4115,N_1533,N_1126);
nand U4116 (N_4116,N_2404,N_1560);
xnor U4117 (N_4117,N_2086,N_1315);
nor U4118 (N_4118,N_331,N_554);
nand U4119 (N_4119,N_2024,N_165);
and U4120 (N_4120,N_113,N_1361);
and U4121 (N_4121,N_1717,N_674);
or U4122 (N_4122,N_1135,N_1613);
or U4123 (N_4123,N_430,N_114);
or U4124 (N_4124,N_865,N_2020);
xor U4125 (N_4125,N_119,N_2126);
and U4126 (N_4126,N_777,N_776);
nor U4127 (N_4127,N_883,N_74);
nor U4128 (N_4128,N_2483,N_1278);
and U4129 (N_4129,N_2468,N_2249);
nand U4130 (N_4130,N_1345,N_493);
nor U4131 (N_4131,N_664,N_1134);
nor U4132 (N_4132,N_1010,N_2430);
nand U4133 (N_4133,N_2301,N_1650);
and U4134 (N_4134,N_31,N_988);
nor U4135 (N_4135,N_847,N_321);
nor U4136 (N_4136,N_357,N_2391);
nand U4137 (N_4137,N_2044,N_605);
or U4138 (N_4138,N_2407,N_1321);
or U4139 (N_4139,N_1004,N_897);
and U4140 (N_4140,N_187,N_2272);
or U4141 (N_4141,N_591,N_2089);
or U4142 (N_4142,N_1090,N_1485);
or U4143 (N_4143,N_528,N_2036);
or U4144 (N_4144,N_1399,N_1653);
or U4145 (N_4145,N_1105,N_983);
and U4146 (N_4146,N_659,N_1092);
nor U4147 (N_4147,N_689,N_946);
nand U4148 (N_4148,N_2408,N_1806);
or U4149 (N_4149,N_639,N_620);
or U4150 (N_4150,N_1559,N_1475);
nor U4151 (N_4151,N_1207,N_1898);
or U4152 (N_4152,N_1062,N_1557);
and U4153 (N_4153,N_2389,N_1269);
and U4154 (N_4154,N_25,N_1901);
or U4155 (N_4155,N_53,N_228);
nor U4156 (N_4156,N_443,N_237);
and U4157 (N_4157,N_1502,N_649);
and U4158 (N_4158,N_1597,N_322);
nor U4159 (N_4159,N_1371,N_346);
xor U4160 (N_4160,N_1046,N_830);
nand U4161 (N_4161,N_1632,N_671);
and U4162 (N_4162,N_86,N_2412);
xnor U4163 (N_4163,N_1654,N_573);
nor U4164 (N_4164,N_1646,N_2058);
nand U4165 (N_4165,N_468,N_406);
or U4166 (N_4166,N_90,N_1116);
and U4167 (N_4167,N_797,N_1526);
nand U4168 (N_4168,N_900,N_2077);
nand U4169 (N_4169,N_1064,N_1502);
or U4170 (N_4170,N_267,N_381);
nor U4171 (N_4171,N_1368,N_2237);
nor U4172 (N_4172,N_1619,N_1555);
or U4173 (N_4173,N_1162,N_2219);
xor U4174 (N_4174,N_350,N_1432);
nor U4175 (N_4175,N_986,N_1750);
nand U4176 (N_4176,N_1967,N_285);
and U4177 (N_4177,N_736,N_738);
nor U4178 (N_4178,N_2108,N_2043);
and U4179 (N_4179,N_2437,N_1347);
or U4180 (N_4180,N_2464,N_1427);
nor U4181 (N_4181,N_2427,N_395);
nor U4182 (N_4182,N_56,N_241);
or U4183 (N_4183,N_815,N_259);
nand U4184 (N_4184,N_1716,N_441);
or U4185 (N_4185,N_2224,N_2498);
and U4186 (N_4186,N_1356,N_2070);
nor U4187 (N_4187,N_1620,N_2383);
nand U4188 (N_4188,N_2388,N_1883);
nand U4189 (N_4189,N_67,N_48);
nand U4190 (N_4190,N_1304,N_2243);
and U4191 (N_4191,N_136,N_1368);
nand U4192 (N_4192,N_2302,N_1974);
and U4193 (N_4193,N_2236,N_384);
and U4194 (N_4194,N_1707,N_849);
nor U4195 (N_4195,N_1029,N_1504);
nor U4196 (N_4196,N_1654,N_772);
nor U4197 (N_4197,N_710,N_448);
or U4198 (N_4198,N_2001,N_741);
and U4199 (N_4199,N_1297,N_866);
or U4200 (N_4200,N_2364,N_1182);
nor U4201 (N_4201,N_355,N_1563);
or U4202 (N_4202,N_1453,N_2327);
and U4203 (N_4203,N_76,N_1090);
xnor U4204 (N_4204,N_1047,N_1261);
xnor U4205 (N_4205,N_1074,N_260);
nand U4206 (N_4206,N_999,N_179);
and U4207 (N_4207,N_668,N_1069);
or U4208 (N_4208,N_166,N_1426);
nor U4209 (N_4209,N_15,N_1704);
nor U4210 (N_4210,N_72,N_2266);
nand U4211 (N_4211,N_1536,N_729);
nand U4212 (N_4212,N_21,N_953);
nand U4213 (N_4213,N_1354,N_1455);
nand U4214 (N_4214,N_345,N_1939);
and U4215 (N_4215,N_290,N_114);
nor U4216 (N_4216,N_1538,N_346);
or U4217 (N_4217,N_1848,N_512);
nor U4218 (N_4218,N_1917,N_1304);
or U4219 (N_4219,N_516,N_2257);
nor U4220 (N_4220,N_872,N_1637);
nand U4221 (N_4221,N_389,N_2205);
and U4222 (N_4222,N_1279,N_1951);
or U4223 (N_4223,N_836,N_1270);
nor U4224 (N_4224,N_1756,N_2265);
nor U4225 (N_4225,N_2166,N_1168);
and U4226 (N_4226,N_512,N_992);
nand U4227 (N_4227,N_2297,N_1776);
or U4228 (N_4228,N_1908,N_1818);
and U4229 (N_4229,N_1583,N_2095);
nand U4230 (N_4230,N_523,N_2026);
nand U4231 (N_4231,N_883,N_301);
nor U4232 (N_4232,N_1494,N_678);
or U4233 (N_4233,N_116,N_2286);
or U4234 (N_4234,N_1047,N_648);
or U4235 (N_4235,N_2262,N_851);
and U4236 (N_4236,N_2102,N_775);
xnor U4237 (N_4237,N_2439,N_2328);
or U4238 (N_4238,N_2442,N_835);
nand U4239 (N_4239,N_2250,N_1028);
nand U4240 (N_4240,N_128,N_14);
nor U4241 (N_4241,N_1746,N_377);
nor U4242 (N_4242,N_2487,N_611);
xnor U4243 (N_4243,N_1484,N_1233);
nand U4244 (N_4244,N_720,N_972);
and U4245 (N_4245,N_1420,N_901);
or U4246 (N_4246,N_1566,N_362);
nor U4247 (N_4247,N_1065,N_232);
or U4248 (N_4248,N_434,N_1728);
xor U4249 (N_4249,N_321,N_1429);
nor U4250 (N_4250,N_1253,N_1577);
nand U4251 (N_4251,N_2038,N_1260);
and U4252 (N_4252,N_2462,N_1619);
or U4253 (N_4253,N_787,N_910);
and U4254 (N_4254,N_1347,N_2060);
or U4255 (N_4255,N_1294,N_728);
nand U4256 (N_4256,N_1085,N_890);
nor U4257 (N_4257,N_1704,N_1093);
or U4258 (N_4258,N_1436,N_527);
nor U4259 (N_4259,N_25,N_816);
nor U4260 (N_4260,N_1612,N_1280);
and U4261 (N_4261,N_582,N_1833);
nand U4262 (N_4262,N_572,N_1423);
nor U4263 (N_4263,N_1042,N_1069);
nor U4264 (N_4264,N_1962,N_758);
nor U4265 (N_4265,N_528,N_2219);
nand U4266 (N_4266,N_1119,N_244);
nor U4267 (N_4267,N_26,N_903);
nor U4268 (N_4268,N_1261,N_1689);
or U4269 (N_4269,N_399,N_1570);
nor U4270 (N_4270,N_1089,N_1792);
or U4271 (N_4271,N_804,N_797);
nand U4272 (N_4272,N_1297,N_99);
and U4273 (N_4273,N_2022,N_1615);
or U4274 (N_4274,N_438,N_1262);
nor U4275 (N_4275,N_536,N_1668);
and U4276 (N_4276,N_1748,N_1791);
and U4277 (N_4277,N_981,N_375);
nand U4278 (N_4278,N_682,N_1099);
and U4279 (N_4279,N_1780,N_165);
xnor U4280 (N_4280,N_1078,N_620);
or U4281 (N_4281,N_1235,N_675);
and U4282 (N_4282,N_2246,N_1373);
and U4283 (N_4283,N_2406,N_144);
or U4284 (N_4284,N_506,N_423);
and U4285 (N_4285,N_323,N_101);
nor U4286 (N_4286,N_1566,N_1393);
and U4287 (N_4287,N_1744,N_499);
nor U4288 (N_4288,N_2230,N_4);
and U4289 (N_4289,N_1173,N_2434);
nor U4290 (N_4290,N_606,N_1194);
and U4291 (N_4291,N_46,N_177);
and U4292 (N_4292,N_1179,N_528);
nor U4293 (N_4293,N_1901,N_907);
nor U4294 (N_4294,N_1727,N_2166);
nor U4295 (N_4295,N_1618,N_1807);
nor U4296 (N_4296,N_1952,N_665);
and U4297 (N_4297,N_557,N_496);
or U4298 (N_4298,N_1397,N_197);
or U4299 (N_4299,N_2151,N_1758);
nor U4300 (N_4300,N_102,N_760);
or U4301 (N_4301,N_69,N_186);
and U4302 (N_4302,N_208,N_737);
nand U4303 (N_4303,N_199,N_2123);
nand U4304 (N_4304,N_604,N_2044);
and U4305 (N_4305,N_2384,N_1554);
xnor U4306 (N_4306,N_988,N_2180);
xnor U4307 (N_4307,N_1917,N_455);
or U4308 (N_4308,N_2290,N_1916);
and U4309 (N_4309,N_1220,N_1328);
and U4310 (N_4310,N_295,N_1228);
nand U4311 (N_4311,N_1962,N_1396);
or U4312 (N_4312,N_1006,N_1790);
nand U4313 (N_4313,N_2244,N_2316);
and U4314 (N_4314,N_62,N_1829);
nand U4315 (N_4315,N_1646,N_2208);
nand U4316 (N_4316,N_1910,N_1268);
and U4317 (N_4317,N_1540,N_1108);
and U4318 (N_4318,N_1037,N_1577);
or U4319 (N_4319,N_1925,N_1656);
nor U4320 (N_4320,N_537,N_1391);
nor U4321 (N_4321,N_861,N_1458);
and U4322 (N_4322,N_1834,N_1603);
nand U4323 (N_4323,N_173,N_750);
nand U4324 (N_4324,N_218,N_1712);
or U4325 (N_4325,N_538,N_2429);
xnor U4326 (N_4326,N_1469,N_99);
or U4327 (N_4327,N_1703,N_2444);
and U4328 (N_4328,N_379,N_517);
nor U4329 (N_4329,N_731,N_319);
nand U4330 (N_4330,N_2191,N_993);
nor U4331 (N_4331,N_1492,N_2042);
nor U4332 (N_4332,N_560,N_602);
nand U4333 (N_4333,N_984,N_1850);
or U4334 (N_4334,N_2041,N_1747);
and U4335 (N_4335,N_645,N_2292);
or U4336 (N_4336,N_1240,N_179);
nor U4337 (N_4337,N_2292,N_1648);
and U4338 (N_4338,N_550,N_136);
nand U4339 (N_4339,N_1287,N_1416);
or U4340 (N_4340,N_1647,N_420);
nand U4341 (N_4341,N_1140,N_600);
nor U4342 (N_4342,N_1028,N_2156);
nor U4343 (N_4343,N_2444,N_1849);
nand U4344 (N_4344,N_1573,N_2168);
nand U4345 (N_4345,N_1117,N_1498);
nand U4346 (N_4346,N_2223,N_2297);
and U4347 (N_4347,N_181,N_882);
and U4348 (N_4348,N_2312,N_1133);
and U4349 (N_4349,N_1981,N_1417);
and U4350 (N_4350,N_376,N_272);
and U4351 (N_4351,N_192,N_1897);
or U4352 (N_4352,N_1270,N_2392);
and U4353 (N_4353,N_382,N_1577);
xor U4354 (N_4354,N_604,N_715);
nor U4355 (N_4355,N_2167,N_75);
or U4356 (N_4356,N_1635,N_486);
nand U4357 (N_4357,N_574,N_677);
nor U4358 (N_4358,N_1643,N_2479);
nand U4359 (N_4359,N_631,N_2163);
or U4360 (N_4360,N_1247,N_1901);
nand U4361 (N_4361,N_1283,N_998);
nand U4362 (N_4362,N_85,N_1810);
nand U4363 (N_4363,N_1051,N_1984);
or U4364 (N_4364,N_2014,N_577);
nor U4365 (N_4365,N_2149,N_1150);
nand U4366 (N_4366,N_1391,N_962);
or U4367 (N_4367,N_1355,N_1698);
and U4368 (N_4368,N_1178,N_1671);
xor U4369 (N_4369,N_2244,N_1228);
nand U4370 (N_4370,N_1284,N_646);
xnor U4371 (N_4371,N_2001,N_103);
xor U4372 (N_4372,N_2085,N_12);
nand U4373 (N_4373,N_1664,N_62);
or U4374 (N_4374,N_1197,N_2037);
xnor U4375 (N_4375,N_510,N_2202);
or U4376 (N_4376,N_2469,N_1513);
nand U4377 (N_4377,N_588,N_1742);
and U4378 (N_4378,N_2272,N_1432);
or U4379 (N_4379,N_788,N_929);
nand U4380 (N_4380,N_449,N_251);
and U4381 (N_4381,N_2399,N_1518);
and U4382 (N_4382,N_486,N_1739);
and U4383 (N_4383,N_2496,N_874);
or U4384 (N_4384,N_1260,N_1425);
and U4385 (N_4385,N_1221,N_1811);
and U4386 (N_4386,N_1289,N_947);
nand U4387 (N_4387,N_2348,N_2366);
and U4388 (N_4388,N_339,N_1954);
and U4389 (N_4389,N_308,N_1024);
nor U4390 (N_4390,N_794,N_1425);
xor U4391 (N_4391,N_1319,N_1411);
nand U4392 (N_4392,N_906,N_2330);
and U4393 (N_4393,N_161,N_544);
nand U4394 (N_4394,N_2308,N_973);
nand U4395 (N_4395,N_2494,N_1215);
and U4396 (N_4396,N_2382,N_75);
and U4397 (N_4397,N_2314,N_1740);
nand U4398 (N_4398,N_127,N_104);
and U4399 (N_4399,N_1821,N_1000);
or U4400 (N_4400,N_615,N_1088);
and U4401 (N_4401,N_2234,N_2157);
nor U4402 (N_4402,N_1329,N_240);
nand U4403 (N_4403,N_1378,N_2126);
nor U4404 (N_4404,N_2407,N_1741);
nand U4405 (N_4405,N_2181,N_149);
or U4406 (N_4406,N_2042,N_781);
nor U4407 (N_4407,N_1604,N_2034);
nor U4408 (N_4408,N_1773,N_1669);
nor U4409 (N_4409,N_728,N_646);
or U4410 (N_4410,N_455,N_2064);
nor U4411 (N_4411,N_2480,N_270);
nor U4412 (N_4412,N_2435,N_449);
nor U4413 (N_4413,N_1069,N_2463);
nor U4414 (N_4414,N_723,N_1474);
nand U4415 (N_4415,N_1139,N_1647);
or U4416 (N_4416,N_1060,N_868);
nor U4417 (N_4417,N_922,N_1885);
nand U4418 (N_4418,N_189,N_335);
and U4419 (N_4419,N_2145,N_484);
and U4420 (N_4420,N_967,N_899);
nand U4421 (N_4421,N_2129,N_711);
nor U4422 (N_4422,N_727,N_714);
xnor U4423 (N_4423,N_2017,N_1154);
and U4424 (N_4424,N_958,N_1613);
nor U4425 (N_4425,N_2300,N_98);
nand U4426 (N_4426,N_430,N_2281);
nor U4427 (N_4427,N_209,N_1871);
nor U4428 (N_4428,N_2076,N_66);
nand U4429 (N_4429,N_759,N_1181);
nor U4430 (N_4430,N_1248,N_911);
nor U4431 (N_4431,N_1517,N_768);
and U4432 (N_4432,N_825,N_1014);
or U4433 (N_4433,N_2107,N_568);
nor U4434 (N_4434,N_431,N_388);
and U4435 (N_4435,N_1163,N_1532);
nand U4436 (N_4436,N_249,N_960);
nor U4437 (N_4437,N_635,N_2489);
nor U4438 (N_4438,N_2009,N_1412);
nor U4439 (N_4439,N_77,N_120);
nor U4440 (N_4440,N_1509,N_2415);
and U4441 (N_4441,N_2198,N_2033);
and U4442 (N_4442,N_2223,N_2365);
nor U4443 (N_4443,N_1797,N_2299);
nand U4444 (N_4444,N_1302,N_1285);
or U4445 (N_4445,N_542,N_34);
nand U4446 (N_4446,N_2421,N_1988);
and U4447 (N_4447,N_346,N_532);
or U4448 (N_4448,N_1669,N_1459);
nor U4449 (N_4449,N_2276,N_1626);
nor U4450 (N_4450,N_2179,N_142);
or U4451 (N_4451,N_1178,N_319);
or U4452 (N_4452,N_925,N_83);
or U4453 (N_4453,N_343,N_711);
nor U4454 (N_4454,N_357,N_759);
nor U4455 (N_4455,N_157,N_2153);
or U4456 (N_4456,N_1710,N_2354);
or U4457 (N_4457,N_1316,N_402);
or U4458 (N_4458,N_1707,N_9);
nor U4459 (N_4459,N_1566,N_494);
or U4460 (N_4460,N_1021,N_1528);
nor U4461 (N_4461,N_1851,N_1536);
or U4462 (N_4462,N_968,N_2340);
and U4463 (N_4463,N_2093,N_707);
nor U4464 (N_4464,N_1224,N_274);
nand U4465 (N_4465,N_91,N_1065);
nand U4466 (N_4466,N_1915,N_360);
or U4467 (N_4467,N_353,N_1351);
and U4468 (N_4468,N_783,N_257);
nand U4469 (N_4469,N_594,N_1616);
and U4470 (N_4470,N_238,N_1821);
and U4471 (N_4471,N_2467,N_1708);
nor U4472 (N_4472,N_2212,N_116);
or U4473 (N_4473,N_1852,N_1728);
and U4474 (N_4474,N_760,N_1942);
xor U4475 (N_4475,N_140,N_1926);
and U4476 (N_4476,N_954,N_1627);
nand U4477 (N_4477,N_1026,N_2237);
or U4478 (N_4478,N_2452,N_266);
and U4479 (N_4479,N_1996,N_782);
nor U4480 (N_4480,N_496,N_2148);
or U4481 (N_4481,N_489,N_782);
and U4482 (N_4482,N_1457,N_2179);
and U4483 (N_4483,N_1481,N_541);
nor U4484 (N_4484,N_300,N_2382);
and U4485 (N_4485,N_1327,N_1476);
nor U4486 (N_4486,N_1526,N_870);
and U4487 (N_4487,N_1348,N_377);
nor U4488 (N_4488,N_468,N_114);
nor U4489 (N_4489,N_1333,N_858);
nand U4490 (N_4490,N_1212,N_1133);
or U4491 (N_4491,N_347,N_1867);
and U4492 (N_4492,N_1730,N_306);
and U4493 (N_4493,N_644,N_821);
xor U4494 (N_4494,N_2003,N_2370);
nor U4495 (N_4495,N_1500,N_1164);
nor U4496 (N_4496,N_1440,N_802);
nand U4497 (N_4497,N_1331,N_1478);
nor U4498 (N_4498,N_431,N_1320);
and U4499 (N_4499,N_620,N_1208);
or U4500 (N_4500,N_259,N_2216);
or U4501 (N_4501,N_1962,N_711);
nand U4502 (N_4502,N_1882,N_270);
nand U4503 (N_4503,N_2231,N_920);
nand U4504 (N_4504,N_1113,N_1475);
nor U4505 (N_4505,N_437,N_1952);
and U4506 (N_4506,N_962,N_909);
and U4507 (N_4507,N_1246,N_1957);
nor U4508 (N_4508,N_1722,N_817);
nand U4509 (N_4509,N_168,N_2131);
nand U4510 (N_4510,N_911,N_1801);
nand U4511 (N_4511,N_171,N_2084);
or U4512 (N_4512,N_2259,N_1400);
and U4513 (N_4513,N_364,N_1055);
or U4514 (N_4514,N_1634,N_2439);
nand U4515 (N_4515,N_214,N_1168);
and U4516 (N_4516,N_1813,N_998);
or U4517 (N_4517,N_94,N_2236);
and U4518 (N_4518,N_2449,N_1563);
nand U4519 (N_4519,N_566,N_317);
nor U4520 (N_4520,N_1575,N_242);
xor U4521 (N_4521,N_519,N_1388);
nor U4522 (N_4522,N_1916,N_2204);
or U4523 (N_4523,N_2098,N_67);
nor U4524 (N_4524,N_1984,N_1618);
nand U4525 (N_4525,N_1022,N_354);
nand U4526 (N_4526,N_1080,N_1534);
or U4527 (N_4527,N_1957,N_1752);
nor U4528 (N_4528,N_1384,N_1915);
nor U4529 (N_4529,N_410,N_2129);
nand U4530 (N_4530,N_799,N_608);
nor U4531 (N_4531,N_2385,N_2467);
and U4532 (N_4532,N_1666,N_322);
nor U4533 (N_4533,N_729,N_437);
nand U4534 (N_4534,N_1327,N_2302);
nand U4535 (N_4535,N_405,N_374);
nor U4536 (N_4536,N_893,N_1353);
nor U4537 (N_4537,N_2411,N_2063);
nand U4538 (N_4538,N_1166,N_2310);
nor U4539 (N_4539,N_1070,N_207);
nand U4540 (N_4540,N_138,N_2069);
and U4541 (N_4541,N_130,N_183);
nand U4542 (N_4542,N_2312,N_2287);
or U4543 (N_4543,N_745,N_645);
and U4544 (N_4544,N_1048,N_2053);
nor U4545 (N_4545,N_1772,N_807);
or U4546 (N_4546,N_402,N_384);
nor U4547 (N_4547,N_1636,N_728);
nor U4548 (N_4548,N_2237,N_2169);
and U4549 (N_4549,N_300,N_313);
nand U4550 (N_4550,N_727,N_1701);
or U4551 (N_4551,N_690,N_2224);
nor U4552 (N_4552,N_2224,N_2180);
nand U4553 (N_4553,N_1763,N_2323);
xor U4554 (N_4554,N_1996,N_2358);
and U4555 (N_4555,N_1984,N_1012);
nand U4556 (N_4556,N_943,N_2192);
nand U4557 (N_4557,N_1478,N_210);
nor U4558 (N_4558,N_499,N_148);
nand U4559 (N_4559,N_1285,N_536);
and U4560 (N_4560,N_765,N_2474);
nand U4561 (N_4561,N_1762,N_489);
nor U4562 (N_4562,N_913,N_1395);
nor U4563 (N_4563,N_1184,N_682);
and U4564 (N_4564,N_1280,N_2420);
nand U4565 (N_4565,N_750,N_1046);
and U4566 (N_4566,N_261,N_1478);
nor U4567 (N_4567,N_18,N_688);
and U4568 (N_4568,N_794,N_2129);
or U4569 (N_4569,N_1184,N_1403);
and U4570 (N_4570,N_1375,N_726);
nand U4571 (N_4571,N_1764,N_2374);
nand U4572 (N_4572,N_557,N_265);
nor U4573 (N_4573,N_1780,N_882);
and U4574 (N_4574,N_1755,N_2496);
nand U4575 (N_4575,N_874,N_1681);
and U4576 (N_4576,N_2245,N_606);
nor U4577 (N_4577,N_1966,N_2472);
and U4578 (N_4578,N_2062,N_1758);
or U4579 (N_4579,N_318,N_2200);
xor U4580 (N_4580,N_985,N_164);
nor U4581 (N_4581,N_2017,N_216);
and U4582 (N_4582,N_908,N_518);
nor U4583 (N_4583,N_1950,N_1915);
or U4584 (N_4584,N_1013,N_2384);
nand U4585 (N_4585,N_169,N_1215);
nor U4586 (N_4586,N_408,N_2060);
or U4587 (N_4587,N_661,N_720);
and U4588 (N_4588,N_696,N_1019);
nand U4589 (N_4589,N_1975,N_1125);
nand U4590 (N_4590,N_665,N_729);
and U4591 (N_4591,N_2087,N_2149);
nand U4592 (N_4592,N_2388,N_2337);
xor U4593 (N_4593,N_595,N_1520);
nor U4594 (N_4594,N_2155,N_226);
nand U4595 (N_4595,N_2470,N_228);
nor U4596 (N_4596,N_795,N_1430);
nand U4597 (N_4597,N_459,N_484);
nand U4598 (N_4598,N_1779,N_986);
nand U4599 (N_4599,N_1380,N_339);
xor U4600 (N_4600,N_185,N_976);
nand U4601 (N_4601,N_171,N_733);
and U4602 (N_4602,N_145,N_828);
and U4603 (N_4603,N_1461,N_848);
and U4604 (N_4604,N_958,N_1072);
nor U4605 (N_4605,N_11,N_1815);
nor U4606 (N_4606,N_1831,N_1784);
and U4607 (N_4607,N_1618,N_2395);
and U4608 (N_4608,N_471,N_530);
nor U4609 (N_4609,N_1144,N_1231);
nor U4610 (N_4610,N_1252,N_771);
or U4611 (N_4611,N_56,N_173);
and U4612 (N_4612,N_2024,N_546);
nor U4613 (N_4613,N_1889,N_519);
xnor U4614 (N_4614,N_1622,N_538);
nor U4615 (N_4615,N_1558,N_645);
or U4616 (N_4616,N_299,N_1641);
nand U4617 (N_4617,N_2229,N_1276);
or U4618 (N_4618,N_246,N_1576);
or U4619 (N_4619,N_1565,N_1192);
nand U4620 (N_4620,N_2280,N_685);
nand U4621 (N_4621,N_2406,N_2263);
nand U4622 (N_4622,N_1566,N_1466);
or U4623 (N_4623,N_539,N_1772);
or U4624 (N_4624,N_902,N_371);
or U4625 (N_4625,N_2221,N_182);
nand U4626 (N_4626,N_1516,N_2322);
or U4627 (N_4627,N_1603,N_1171);
nor U4628 (N_4628,N_346,N_798);
and U4629 (N_4629,N_355,N_1118);
or U4630 (N_4630,N_2341,N_1738);
or U4631 (N_4631,N_350,N_691);
nand U4632 (N_4632,N_934,N_244);
nand U4633 (N_4633,N_1130,N_914);
nand U4634 (N_4634,N_22,N_164);
and U4635 (N_4635,N_303,N_66);
or U4636 (N_4636,N_894,N_2328);
nand U4637 (N_4637,N_1019,N_485);
or U4638 (N_4638,N_561,N_1572);
nand U4639 (N_4639,N_1660,N_278);
nor U4640 (N_4640,N_751,N_1676);
nor U4641 (N_4641,N_809,N_2435);
and U4642 (N_4642,N_980,N_2125);
nor U4643 (N_4643,N_2216,N_2376);
and U4644 (N_4644,N_1881,N_432);
or U4645 (N_4645,N_1079,N_2220);
or U4646 (N_4646,N_753,N_1884);
nor U4647 (N_4647,N_1162,N_1462);
nand U4648 (N_4648,N_172,N_1436);
xnor U4649 (N_4649,N_996,N_553);
nand U4650 (N_4650,N_878,N_1653);
or U4651 (N_4651,N_255,N_2005);
nor U4652 (N_4652,N_17,N_782);
and U4653 (N_4653,N_1866,N_1256);
or U4654 (N_4654,N_2122,N_209);
or U4655 (N_4655,N_753,N_809);
nor U4656 (N_4656,N_472,N_651);
or U4657 (N_4657,N_654,N_2036);
or U4658 (N_4658,N_1111,N_275);
nor U4659 (N_4659,N_90,N_2242);
and U4660 (N_4660,N_1943,N_695);
and U4661 (N_4661,N_564,N_547);
nand U4662 (N_4662,N_282,N_493);
nand U4663 (N_4663,N_2032,N_1709);
or U4664 (N_4664,N_2165,N_576);
and U4665 (N_4665,N_2263,N_1246);
nor U4666 (N_4666,N_226,N_311);
and U4667 (N_4667,N_1940,N_2399);
or U4668 (N_4668,N_947,N_1997);
nand U4669 (N_4669,N_742,N_2085);
or U4670 (N_4670,N_1640,N_339);
nor U4671 (N_4671,N_1621,N_1124);
nor U4672 (N_4672,N_1867,N_1009);
nor U4673 (N_4673,N_1900,N_2499);
or U4674 (N_4674,N_2180,N_1659);
or U4675 (N_4675,N_1549,N_2416);
nor U4676 (N_4676,N_1327,N_730);
or U4677 (N_4677,N_73,N_1023);
or U4678 (N_4678,N_1946,N_1728);
nor U4679 (N_4679,N_1167,N_2424);
nand U4680 (N_4680,N_613,N_2253);
or U4681 (N_4681,N_730,N_338);
nand U4682 (N_4682,N_723,N_974);
nand U4683 (N_4683,N_85,N_2013);
nor U4684 (N_4684,N_1172,N_117);
xnor U4685 (N_4685,N_2469,N_258);
nor U4686 (N_4686,N_2189,N_163);
nand U4687 (N_4687,N_139,N_820);
or U4688 (N_4688,N_1747,N_1110);
or U4689 (N_4689,N_1555,N_1527);
nor U4690 (N_4690,N_1753,N_669);
nor U4691 (N_4691,N_2165,N_755);
nor U4692 (N_4692,N_439,N_722);
nor U4693 (N_4693,N_1964,N_591);
xor U4694 (N_4694,N_2459,N_1022);
nor U4695 (N_4695,N_893,N_2416);
and U4696 (N_4696,N_554,N_16);
xor U4697 (N_4697,N_2309,N_1514);
or U4698 (N_4698,N_122,N_304);
nor U4699 (N_4699,N_430,N_2398);
and U4700 (N_4700,N_2041,N_2167);
xor U4701 (N_4701,N_5,N_2213);
nor U4702 (N_4702,N_2386,N_946);
nor U4703 (N_4703,N_2028,N_424);
nor U4704 (N_4704,N_1301,N_414);
or U4705 (N_4705,N_186,N_1366);
nor U4706 (N_4706,N_771,N_524);
or U4707 (N_4707,N_1319,N_1500);
and U4708 (N_4708,N_202,N_330);
nor U4709 (N_4709,N_2373,N_1210);
nor U4710 (N_4710,N_1016,N_593);
nor U4711 (N_4711,N_2147,N_1683);
and U4712 (N_4712,N_836,N_2474);
nand U4713 (N_4713,N_2333,N_1462);
and U4714 (N_4714,N_2192,N_1188);
nand U4715 (N_4715,N_1799,N_100);
xnor U4716 (N_4716,N_2443,N_1369);
nor U4717 (N_4717,N_1905,N_1696);
nand U4718 (N_4718,N_1467,N_337);
nor U4719 (N_4719,N_40,N_844);
nor U4720 (N_4720,N_524,N_1814);
and U4721 (N_4721,N_704,N_2395);
nand U4722 (N_4722,N_1705,N_2059);
nand U4723 (N_4723,N_647,N_1009);
nor U4724 (N_4724,N_433,N_791);
nor U4725 (N_4725,N_551,N_2102);
or U4726 (N_4726,N_2050,N_1441);
nand U4727 (N_4727,N_180,N_2228);
nand U4728 (N_4728,N_572,N_1277);
and U4729 (N_4729,N_1258,N_1408);
nand U4730 (N_4730,N_1834,N_1140);
xor U4731 (N_4731,N_2205,N_652);
or U4732 (N_4732,N_1317,N_1971);
nand U4733 (N_4733,N_962,N_2299);
or U4734 (N_4734,N_1521,N_2035);
and U4735 (N_4735,N_674,N_2433);
or U4736 (N_4736,N_2491,N_92);
nand U4737 (N_4737,N_304,N_1639);
xnor U4738 (N_4738,N_1417,N_801);
nor U4739 (N_4739,N_1317,N_1941);
nand U4740 (N_4740,N_1547,N_1457);
xnor U4741 (N_4741,N_1460,N_1534);
and U4742 (N_4742,N_444,N_325);
or U4743 (N_4743,N_1633,N_434);
or U4744 (N_4744,N_96,N_983);
and U4745 (N_4745,N_1509,N_348);
or U4746 (N_4746,N_1278,N_237);
nand U4747 (N_4747,N_1100,N_1543);
xor U4748 (N_4748,N_870,N_2373);
nor U4749 (N_4749,N_1417,N_1390);
nor U4750 (N_4750,N_169,N_1095);
or U4751 (N_4751,N_930,N_1195);
nor U4752 (N_4752,N_2360,N_476);
nor U4753 (N_4753,N_1175,N_2031);
nor U4754 (N_4754,N_2362,N_580);
nor U4755 (N_4755,N_1584,N_359);
nor U4756 (N_4756,N_2144,N_2066);
and U4757 (N_4757,N_1873,N_2141);
nand U4758 (N_4758,N_2452,N_582);
and U4759 (N_4759,N_2336,N_2127);
nor U4760 (N_4760,N_68,N_79);
nor U4761 (N_4761,N_810,N_1018);
nand U4762 (N_4762,N_605,N_1222);
and U4763 (N_4763,N_486,N_441);
nand U4764 (N_4764,N_1684,N_1683);
or U4765 (N_4765,N_1707,N_731);
nand U4766 (N_4766,N_1286,N_849);
nand U4767 (N_4767,N_1205,N_1237);
and U4768 (N_4768,N_996,N_2329);
and U4769 (N_4769,N_659,N_1753);
or U4770 (N_4770,N_2469,N_1010);
or U4771 (N_4771,N_1771,N_193);
and U4772 (N_4772,N_98,N_1541);
or U4773 (N_4773,N_1069,N_922);
nand U4774 (N_4774,N_2272,N_121);
nand U4775 (N_4775,N_2143,N_2409);
or U4776 (N_4776,N_1545,N_1367);
nor U4777 (N_4777,N_264,N_1891);
and U4778 (N_4778,N_1032,N_1061);
nor U4779 (N_4779,N_410,N_432);
or U4780 (N_4780,N_256,N_1837);
or U4781 (N_4781,N_845,N_567);
nor U4782 (N_4782,N_1121,N_666);
and U4783 (N_4783,N_1666,N_2231);
nand U4784 (N_4784,N_616,N_754);
nand U4785 (N_4785,N_2440,N_488);
and U4786 (N_4786,N_5,N_2275);
nand U4787 (N_4787,N_272,N_1524);
nand U4788 (N_4788,N_264,N_1785);
nand U4789 (N_4789,N_81,N_218);
and U4790 (N_4790,N_75,N_1509);
and U4791 (N_4791,N_822,N_2060);
nor U4792 (N_4792,N_2077,N_2143);
nor U4793 (N_4793,N_1023,N_2289);
xor U4794 (N_4794,N_931,N_2313);
and U4795 (N_4795,N_650,N_1980);
and U4796 (N_4796,N_752,N_278);
and U4797 (N_4797,N_489,N_704);
nand U4798 (N_4798,N_2449,N_967);
nor U4799 (N_4799,N_434,N_1976);
nor U4800 (N_4800,N_2151,N_1026);
or U4801 (N_4801,N_587,N_1347);
nor U4802 (N_4802,N_445,N_1767);
nand U4803 (N_4803,N_939,N_1369);
or U4804 (N_4804,N_2266,N_1409);
nand U4805 (N_4805,N_576,N_827);
nand U4806 (N_4806,N_1492,N_2431);
or U4807 (N_4807,N_1404,N_37);
nor U4808 (N_4808,N_33,N_318);
nand U4809 (N_4809,N_1055,N_2487);
or U4810 (N_4810,N_1293,N_2149);
nor U4811 (N_4811,N_425,N_1173);
or U4812 (N_4812,N_2073,N_1675);
nor U4813 (N_4813,N_419,N_1391);
or U4814 (N_4814,N_710,N_484);
and U4815 (N_4815,N_1369,N_584);
or U4816 (N_4816,N_117,N_238);
nand U4817 (N_4817,N_172,N_1063);
or U4818 (N_4818,N_11,N_2158);
or U4819 (N_4819,N_544,N_1082);
nor U4820 (N_4820,N_838,N_639);
or U4821 (N_4821,N_1315,N_678);
nand U4822 (N_4822,N_1549,N_80);
nor U4823 (N_4823,N_2080,N_125);
and U4824 (N_4824,N_107,N_660);
nand U4825 (N_4825,N_2495,N_1635);
or U4826 (N_4826,N_537,N_2407);
and U4827 (N_4827,N_750,N_1028);
nor U4828 (N_4828,N_1014,N_770);
nand U4829 (N_4829,N_1258,N_2484);
and U4830 (N_4830,N_1105,N_1210);
nand U4831 (N_4831,N_1454,N_1111);
nor U4832 (N_4832,N_511,N_813);
nand U4833 (N_4833,N_468,N_670);
and U4834 (N_4834,N_514,N_341);
nor U4835 (N_4835,N_466,N_1666);
or U4836 (N_4836,N_342,N_416);
nor U4837 (N_4837,N_180,N_294);
nor U4838 (N_4838,N_630,N_1426);
xnor U4839 (N_4839,N_57,N_1929);
nor U4840 (N_4840,N_1342,N_452);
and U4841 (N_4841,N_310,N_42);
and U4842 (N_4842,N_1322,N_1190);
nand U4843 (N_4843,N_2401,N_1014);
and U4844 (N_4844,N_2450,N_81);
or U4845 (N_4845,N_1850,N_42);
or U4846 (N_4846,N_2042,N_968);
or U4847 (N_4847,N_1108,N_1811);
nor U4848 (N_4848,N_1480,N_991);
and U4849 (N_4849,N_1180,N_582);
nand U4850 (N_4850,N_1354,N_945);
nor U4851 (N_4851,N_968,N_1576);
and U4852 (N_4852,N_299,N_1776);
nor U4853 (N_4853,N_2078,N_1860);
or U4854 (N_4854,N_1890,N_803);
nor U4855 (N_4855,N_428,N_1024);
and U4856 (N_4856,N_1461,N_470);
nor U4857 (N_4857,N_2199,N_1572);
or U4858 (N_4858,N_378,N_1201);
nor U4859 (N_4859,N_2242,N_2321);
nor U4860 (N_4860,N_338,N_1339);
nand U4861 (N_4861,N_1799,N_1215);
and U4862 (N_4862,N_1464,N_1390);
or U4863 (N_4863,N_1805,N_2102);
nand U4864 (N_4864,N_1328,N_1399);
nor U4865 (N_4865,N_1476,N_1759);
nand U4866 (N_4866,N_488,N_2142);
or U4867 (N_4867,N_1335,N_1664);
or U4868 (N_4868,N_142,N_2047);
nand U4869 (N_4869,N_1804,N_491);
nand U4870 (N_4870,N_1670,N_1832);
or U4871 (N_4871,N_1603,N_241);
nor U4872 (N_4872,N_642,N_1936);
nand U4873 (N_4873,N_1459,N_1051);
and U4874 (N_4874,N_2375,N_1901);
and U4875 (N_4875,N_1085,N_578);
nor U4876 (N_4876,N_1645,N_164);
xnor U4877 (N_4877,N_1544,N_1701);
or U4878 (N_4878,N_1461,N_1788);
or U4879 (N_4879,N_392,N_1710);
nor U4880 (N_4880,N_385,N_2256);
and U4881 (N_4881,N_1031,N_2011);
or U4882 (N_4882,N_138,N_922);
and U4883 (N_4883,N_2244,N_1728);
or U4884 (N_4884,N_162,N_1104);
and U4885 (N_4885,N_2470,N_1828);
or U4886 (N_4886,N_1300,N_2095);
and U4887 (N_4887,N_946,N_1121);
nor U4888 (N_4888,N_2062,N_1927);
or U4889 (N_4889,N_2291,N_1314);
xor U4890 (N_4890,N_1965,N_379);
or U4891 (N_4891,N_2348,N_1071);
and U4892 (N_4892,N_1005,N_1629);
nor U4893 (N_4893,N_259,N_529);
and U4894 (N_4894,N_2256,N_1510);
nand U4895 (N_4895,N_2036,N_284);
or U4896 (N_4896,N_1122,N_1563);
or U4897 (N_4897,N_1287,N_516);
nand U4898 (N_4898,N_1526,N_1813);
nand U4899 (N_4899,N_11,N_787);
and U4900 (N_4900,N_679,N_705);
and U4901 (N_4901,N_657,N_1045);
nor U4902 (N_4902,N_587,N_249);
nand U4903 (N_4903,N_2319,N_1957);
nand U4904 (N_4904,N_2202,N_1409);
and U4905 (N_4905,N_345,N_1067);
nand U4906 (N_4906,N_2142,N_2494);
nand U4907 (N_4907,N_2318,N_1064);
nor U4908 (N_4908,N_129,N_2286);
and U4909 (N_4909,N_1146,N_1088);
nor U4910 (N_4910,N_2173,N_505);
and U4911 (N_4911,N_1928,N_1740);
nor U4912 (N_4912,N_1033,N_1923);
nand U4913 (N_4913,N_2225,N_2490);
and U4914 (N_4914,N_2177,N_1616);
or U4915 (N_4915,N_612,N_2142);
nor U4916 (N_4916,N_1340,N_1083);
nand U4917 (N_4917,N_1722,N_868);
xnor U4918 (N_4918,N_1335,N_924);
and U4919 (N_4919,N_1488,N_9);
nor U4920 (N_4920,N_1779,N_1463);
nor U4921 (N_4921,N_1070,N_2193);
xnor U4922 (N_4922,N_1586,N_2147);
or U4923 (N_4923,N_1068,N_220);
or U4924 (N_4924,N_1471,N_2353);
or U4925 (N_4925,N_691,N_127);
and U4926 (N_4926,N_1174,N_144);
or U4927 (N_4927,N_2248,N_1754);
and U4928 (N_4928,N_1240,N_106);
nor U4929 (N_4929,N_2019,N_600);
or U4930 (N_4930,N_547,N_70);
or U4931 (N_4931,N_1245,N_925);
or U4932 (N_4932,N_835,N_124);
nor U4933 (N_4933,N_1688,N_159);
or U4934 (N_4934,N_1336,N_2070);
and U4935 (N_4935,N_2386,N_360);
or U4936 (N_4936,N_386,N_956);
or U4937 (N_4937,N_332,N_465);
nand U4938 (N_4938,N_1125,N_614);
nor U4939 (N_4939,N_1914,N_917);
or U4940 (N_4940,N_2345,N_629);
or U4941 (N_4941,N_1034,N_1617);
and U4942 (N_4942,N_625,N_272);
nand U4943 (N_4943,N_1160,N_1955);
nand U4944 (N_4944,N_992,N_2364);
nand U4945 (N_4945,N_264,N_2016);
xnor U4946 (N_4946,N_1774,N_2327);
xnor U4947 (N_4947,N_2036,N_2315);
nand U4948 (N_4948,N_765,N_1243);
or U4949 (N_4949,N_2287,N_2370);
and U4950 (N_4950,N_1509,N_2334);
nor U4951 (N_4951,N_1467,N_2340);
nor U4952 (N_4952,N_2493,N_528);
nand U4953 (N_4953,N_397,N_468);
nor U4954 (N_4954,N_2040,N_925);
nand U4955 (N_4955,N_2234,N_1405);
nand U4956 (N_4956,N_1495,N_876);
and U4957 (N_4957,N_1576,N_2221);
or U4958 (N_4958,N_905,N_1283);
and U4959 (N_4959,N_19,N_2279);
nor U4960 (N_4960,N_2433,N_1442);
or U4961 (N_4961,N_372,N_1890);
nor U4962 (N_4962,N_2313,N_570);
or U4963 (N_4963,N_1558,N_1960);
or U4964 (N_4964,N_374,N_2048);
or U4965 (N_4965,N_1554,N_2206);
nor U4966 (N_4966,N_1183,N_209);
and U4967 (N_4967,N_2285,N_1889);
nor U4968 (N_4968,N_248,N_405);
nor U4969 (N_4969,N_1312,N_1252);
nor U4970 (N_4970,N_1869,N_1097);
or U4971 (N_4971,N_2094,N_1366);
and U4972 (N_4972,N_52,N_2082);
nor U4973 (N_4973,N_2244,N_2466);
and U4974 (N_4974,N_506,N_562);
and U4975 (N_4975,N_2450,N_706);
or U4976 (N_4976,N_251,N_1897);
nor U4977 (N_4977,N_390,N_481);
and U4978 (N_4978,N_1635,N_834);
or U4979 (N_4979,N_2111,N_2141);
and U4980 (N_4980,N_1539,N_2458);
nand U4981 (N_4981,N_698,N_2391);
xnor U4982 (N_4982,N_445,N_2084);
nor U4983 (N_4983,N_1772,N_2242);
or U4984 (N_4984,N_2420,N_527);
nor U4985 (N_4985,N_2168,N_1693);
and U4986 (N_4986,N_1590,N_2375);
nor U4987 (N_4987,N_1476,N_879);
nand U4988 (N_4988,N_2298,N_352);
nor U4989 (N_4989,N_1856,N_953);
and U4990 (N_4990,N_2096,N_529);
nand U4991 (N_4991,N_1484,N_2481);
nand U4992 (N_4992,N_1568,N_2408);
and U4993 (N_4993,N_300,N_564);
nor U4994 (N_4994,N_1099,N_181);
and U4995 (N_4995,N_1034,N_56);
nor U4996 (N_4996,N_1945,N_1523);
nor U4997 (N_4997,N_2199,N_365);
nand U4998 (N_4998,N_1531,N_2263);
or U4999 (N_4999,N_446,N_1713);
or UO_0 (O_0,N_3845,N_4727);
nand UO_1 (O_1,N_4048,N_3936);
and UO_2 (O_2,N_3346,N_3345);
nand UO_3 (O_3,N_3026,N_4180);
or UO_4 (O_4,N_3669,N_2584);
nor UO_5 (O_5,N_3348,N_3312);
nand UO_6 (O_6,N_3298,N_3930);
or UO_7 (O_7,N_3404,N_2793);
or UO_8 (O_8,N_3959,N_3239);
nor UO_9 (O_9,N_3440,N_3178);
or UO_10 (O_10,N_4430,N_3821);
or UO_11 (O_11,N_3851,N_4283);
or UO_12 (O_12,N_2900,N_2760);
xor UO_13 (O_13,N_4312,N_4120);
nor UO_14 (O_14,N_3249,N_2885);
and UO_15 (O_15,N_3644,N_4566);
and UO_16 (O_16,N_4446,N_3882);
nor UO_17 (O_17,N_4227,N_2685);
nand UO_18 (O_18,N_4791,N_2517);
nand UO_19 (O_19,N_3973,N_4493);
nor UO_20 (O_20,N_3451,N_3547);
nor UO_21 (O_21,N_2509,N_2840);
and UO_22 (O_22,N_3187,N_2766);
or UO_23 (O_23,N_3482,N_4220);
or UO_24 (O_24,N_3267,N_4639);
or UO_25 (O_25,N_2617,N_4728);
or UO_26 (O_26,N_4015,N_2985);
nand UO_27 (O_27,N_2571,N_3076);
nand UO_28 (O_28,N_2796,N_3251);
or UO_29 (O_29,N_4000,N_3663);
nand UO_30 (O_30,N_3965,N_4274);
nor UO_31 (O_31,N_4334,N_3607);
nor UO_32 (O_32,N_3981,N_2534);
and UO_33 (O_33,N_3020,N_4801);
nand UO_34 (O_34,N_4861,N_4067);
nor UO_35 (O_35,N_2640,N_3692);
or UO_36 (O_36,N_4780,N_4868);
nor UO_37 (O_37,N_2836,N_2594);
and UO_38 (O_38,N_3854,N_4958);
nand UO_39 (O_39,N_4672,N_3627);
or UO_40 (O_40,N_4191,N_4042);
or UO_41 (O_41,N_3218,N_3562);
nand UO_42 (O_42,N_3002,N_4594);
or UO_43 (O_43,N_3250,N_2950);
and UO_44 (O_44,N_3454,N_4117);
and UO_45 (O_45,N_4578,N_3932);
or UO_46 (O_46,N_3695,N_4087);
nor UO_47 (O_47,N_2965,N_3179);
and UO_48 (O_48,N_3197,N_4556);
xnor UO_49 (O_49,N_4060,N_3637);
nand UO_50 (O_50,N_2955,N_4991);
nor UO_51 (O_51,N_2658,N_3484);
nor UO_52 (O_52,N_3261,N_3158);
nand UO_53 (O_53,N_2986,N_2558);
or UO_54 (O_54,N_4455,N_3150);
or UO_55 (O_55,N_2505,N_4628);
nor UO_56 (O_56,N_2742,N_4416);
or UO_57 (O_57,N_2969,N_4472);
or UO_58 (O_58,N_4950,N_4080);
nor UO_59 (O_59,N_4088,N_4857);
nand UO_60 (O_60,N_4890,N_4581);
or UO_61 (O_61,N_3551,N_2661);
and UO_62 (O_62,N_4997,N_3926);
and UO_63 (O_63,N_2798,N_4613);
or UO_64 (O_64,N_3850,N_3183);
and UO_65 (O_65,N_4111,N_4814);
or UO_66 (O_66,N_3013,N_4383);
and UO_67 (O_67,N_2920,N_3691);
nor UO_68 (O_68,N_2516,N_4644);
and UO_69 (O_69,N_3518,N_3423);
or UO_70 (O_70,N_3489,N_4059);
nor UO_71 (O_71,N_4181,N_4030);
or UO_72 (O_72,N_4620,N_2935);
or UO_73 (O_73,N_2618,N_4586);
and UO_74 (O_74,N_2583,N_4846);
nor UO_75 (O_75,N_3861,N_4209);
and UO_76 (O_76,N_4540,N_2990);
and UO_77 (O_77,N_4364,N_4404);
and UO_78 (O_78,N_2768,N_2753);
and UO_79 (O_79,N_4851,N_3855);
nor UO_80 (O_80,N_3635,N_2549);
nand UO_81 (O_81,N_4725,N_4894);
or UO_82 (O_82,N_3652,N_4520);
nand UO_83 (O_83,N_2645,N_4144);
or UO_84 (O_84,N_4542,N_4172);
nand UO_85 (O_85,N_4391,N_3295);
nor UO_86 (O_86,N_3442,N_3340);
or UO_87 (O_87,N_3420,N_4050);
nand UO_88 (O_88,N_3561,N_2653);
and UO_89 (O_89,N_4585,N_3791);
or UO_90 (O_90,N_4462,N_4577);
or UO_91 (O_91,N_3795,N_4698);
nand UO_92 (O_92,N_4273,N_4864);
or UO_93 (O_93,N_4081,N_4339);
xnor UO_94 (O_94,N_2750,N_2528);
nor UO_95 (O_95,N_3784,N_3928);
nand UO_96 (O_96,N_4233,N_3077);
or UO_97 (O_97,N_4760,N_2731);
or UO_98 (O_98,N_4811,N_2677);
nor UO_99 (O_99,N_3500,N_4847);
or UO_100 (O_100,N_4397,N_4762);
nand UO_101 (O_101,N_2867,N_3583);
or UO_102 (O_102,N_2811,N_3503);
or UO_103 (O_103,N_4980,N_3424);
and UO_104 (O_104,N_4400,N_3598);
nor UO_105 (O_105,N_2657,N_2871);
nor UO_106 (O_106,N_3352,N_3058);
and UO_107 (O_107,N_2575,N_4122);
nand UO_108 (O_108,N_4115,N_3105);
and UO_109 (O_109,N_4982,N_4737);
nand UO_110 (O_110,N_4469,N_3242);
and UO_111 (O_111,N_4041,N_4407);
nor UO_112 (O_112,N_4369,N_3710);
or UO_113 (O_113,N_4975,N_4509);
and UO_114 (O_114,N_4948,N_4051);
or UO_115 (O_115,N_4148,N_2971);
and UO_116 (O_116,N_2684,N_2759);
nor UO_117 (O_117,N_3887,N_3931);
or UO_118 (O_118,N_4477,N_3760);
nor UO_119 (O_119,N_3073,N_4217);
or UO_120 (O_120,N_3045,N_2845);
nand UO_121 (O_121,N_4406,N_4300);
or UO_122 (O_122,N_3875,N_2672);
nor UO_123 (O_123,N_3030,N_3771);
nand UO_124 (O_124,N_3055,N_4827);
or UO_125 (O_125,N_4561,N_3284);
nand UO_126 (O_126,N_3481,N_3409);
nor UO_127 (O_127,N_3773,N_4820);
nor UO_128 (O_128,N_2681,N_4190);
and UO_129 (O_129,N_3210,N_3209);
nor UO_130 (O_130,N_4069,N_4084);
nor UO_131 (O_131,N_3804,N_4086);
nor UO_132 (O_132,N_4686,N_4924);
or UO_133 (O_133,N_2737,N_3883);
nand UO_134 (O_134,N_3703,N_2757);
or UO_135 (O_135,N_3288,N_2665);
xnor UO_136 (O_136,N_2560,N_3745);
nor UO_137 (O_137,N_3343,N_4047);
nor UO_138 (O_138,N_3062,N_3359);
nand UO_139 (O_139,N_3042,N_3180);
nor UO_140 (O_140,N_4337,N_3287);
and UO_141 (O_141,N_4387,N_2582);
or UO_142 (O_142,N_2902,N_3625);
nor UO_143 (O_143,N_4900,N_3617);
and UO_144 (O_144,N_4888,N_3508);
or UO_145 (O_145,N_3240,N_4457);
nand UO_146 (O_146,N_3136,N_2813);
nor UO_147 (O_147,N_4641,N_4216);
nor UO_148 (O_148,N_4451,N_4147);
nor UO_149 (O_149,N_3933,N_4971);
nor UO_150 (O_150,N_4419,N_4351);
and UO_151 (O_151,N_3853,N_4956);
and UO_152 (O_152,N_3093,N_4642);
or UO_153 (O_153,N_2777,N_4913);
or UO_154 (O_154,N_3381,N_3046);
nand UO_155 (O_155,N_4607,N_3107);
nand UO_156 (O_156,N_3106,N_4385);
nand UO_157 (O_157,N_3830,N_4010);
and UO_158 (O_158,N_3266,N_2664);
and UO_159 (O_159,N_3719,N_2843);
and UO_160 (O_160,N_2994,N_2577);
nand UO_161 (O_161,N_4507,N_3734);
and UO_162 (O_162,N_3519,N_2713);
or UO_163 (O_163,N_4770,N_3768);
nor UO_164 (O_164,N_2786,N_2816);
nor UO_165 (O_165,N_2898,N_3716);
and UO_166 (O_166,N_4463,N_4916);
and UO_167 (O_167,N_4331,N_3999);
and UO_168 (O_168,N_2561,N_4837);
nor UO_169 (O_169,N_4210,N_4335);
and UO_170 (O_170,N_3976,N_2634);
nand UO_171 (O_171,N_4141,N_3873);
nand UO_172 (O_172,N_3769,N_4155);
nand UO_173 (O_173,N_2693,N_3004);
nor UO_174 (O_174,N_4878,N_3071);
or UO_175 (O_175,N_3596,N_4710);
or UO_176 (O_176,N_2909,N_3560);
or UO_177 (O_177,N_4867,N_4378);
nor UO_178 (O_178,N_3392,N_4241);
or UO_179 (O_179,N_4207,N_3594);
nor UO_180 (O_180,N_3277,N_4782);
and UO_181 (O_181,N_2879,N_4995);
and UO_182 (O_182,N_4242,N_4872);
nor UO_183 (O_183,N_4546,N_3182);
nand UO_184 (O_184,N_4623,N_3735);
nor UO_185 (O_185,N_2890,N_4899);
nor UO_186 (O_186,N_3238,N_3915);
nand UO_187 (O_187,N_3690,N_3629);
nor UO_188 (O_188,N_3104,N_4550);
and UO_189 (O_189,N_3943,N_2773);
and UO_190 (O_190,N_2968,N_3879);
or UO_191 (O_191,N_4631,N_3957);
and UO_192 (O_192,N_4344,N_4445);
nand UO_193 (O_193,N_3807,N_3796);
nand UO_194 (O_194,N_3382,N_4093);
or UO_195 (O_195,N_3800,N_2774);
and UO_196 (O_196,N_3616,N_4150);
or UO_197 (O_197,N_2784,N_3314);
nand UO_198 (O_198,N_4604,N_3731);
nand UO_199 (O_199,N_4151,N_4277);
nor UO_200 (O_200,N_2578,N_4356);
nor UO_201 (O_201,N_3173,N_2642);
nand UO_202 (O_202,N_3896,N_4448);
or UO_203 (O_203,N_4966,N_3523);
nand UO_204 (O_204,N_3511,N_4254);
nor UO_205 (O_205,N_3953,N_3746);
and UO_206 (O_206,N_2799,N_4286);
nand UO_207 (O_207,N_4146,N_2674);
and UO_208 (O_208,N_3864,N_4315);
nor UO_209 (O_209,N_4943,N_3119);
and UO_210 (O_210,N_4792,N_3488);
or UO_211 (O_211,N_3686,N_4492);
or UO_212 (O_212,N_4929,N_3724);
and UO_213 (O_213,N_4307,N_3418);
and UO_214 (O_214,N_4481,N_4596);
or UO_215 (O_215,N_3836,N_3984);
nor UO_216 (O_216,N_3199,N_4454);
nor UO_217 (O_217,N_3444,N_4701);
nor UO_218 (O_218,N_3743,N_4965);
nor UO_219 (O_219,N_4981,N_4215);
nor UO_220 (O_220,N_2789,N_2779);
and UO_221 (O_221,N_3364,N_3964);
or UO_222 (O_222,N_2883,N_2800);
nor UO_223 (O_223,N_2858,N_2919);
nand UO_224 (O_224,N_4373,N_4841);
nor UO_225 (O_225,N_3164,N_3951);
or UO_226 (O_226,N_2551,N_4771);
or UO_227 (O_227,N_2590,N_4055);
nand UO_228 (O_228,N_3112,N_3799);
nor UO_229 (O_229,N_4402,N_4199);
nand UO_230 (O_230,N_4785,N_2751);
nand UO_231 (O_231,N_2629,N_2592);
or UO_232 (O_232,N_3155,N_4862);
nor UO_233 (O_233,N_3079,N_2601);
and UO_234 (O_234,N_3379,N_4558);
or UO_235 (O_235,N_3262,N_3495);
nor UO_236 (O_236,N_3054,N_4858);
and UO_237 (O_237,N_3475,N_3868);
and UO_238 (O_238,N_3986,N_3610);
and UO_239 (O_239,N_2860,N_4699);
nand UO_240 (O_240,N_2842,N_4333);
nand UO_241 (O_241,N_3016,N_3767);
nand UO_242 (O_242,N_2500,N_3315);
xor UO_243 (O_243,N_4127,N_4590);
nand UO_244 (O_244,N_4753,N_4912);
nor UO_245 (O_245,N_3003,N_3177);
nand UO_246 (O_246,N_3064,N_2988);
nor UO_247 (O_247,N_2704,N_4669);
or UO_248 (O_248,N_4935,N_4228);
or UO_249 (O_249,N_2874,N_3506);
and UO_250 (O_250,N_4797,N_3156);
xor UO_251 (O_251,N_3645,N_3826);
and UO_252 (O_252,N_4922,N_3283);
nand UO_253 (O_253,N_2696,N_2649);
nand UO_254 (O_254,N_2585,N_4034);
nand UO_255 (O_255,N_3914,N_2588);
nor UO_256 (O_256,N_3827,N_3019);
and UO_257 (O_257,N_3968,N_3532);
or UO_258 (O_258,N_3752,N_4420);
and UO_259 (O_259,N_2726,N_4504);
or UO_260 (O_260,N_4626,N_2593);
nor UO_261 (O_261,N_3258,N_3720);
or UO_262 (O_262,N_4389,N_4522);
nor UO_263 (O_263,N_3040,N_4094);
nor UO_264 (O_264,N_3660,N_3318);
nand UO_265 (O_265,N_4382,N_2632);
nor UO_266 (O_266,N_3000,N_4608);
nand UO_267 (O_267,N_2729,N_4361);
and UO_268 (O_268,N_2995,N_4173);
nor UO_269 (O_269,N_3694,N_2984);
or UO_270 (O_270,N_4692,N_2944);
nor UO_271 (O_271,N_3176,N_3033);
nor UO_272 (O_272,N_3022,N_3738);
or UO_273 (O_273,N_3718,N_4292);
and UO_274 (O_274,N_3101,N_2947);
and UO_275 (O_275,N_3670,N_4281);
or UO_276 (O_276,N_3200,N_2695);
nor UO_277 (O_277,N_4214,N_3674);
nor UO_278 (O_278,N_2775,N_4517);
nand UO_279 (O_279,N_4936,N_2848);
and UO_280 (O_280,N_3777,N_4362);
nand UO_281 (O_281,N_2613,N_3036);
xor UO_282 (O_282,N_3917,N_3466);
nand UO_283 (O_283,N_3465,N_3877);
or UO_284 (O_284,N_2720,N_3788);
or UO_285 (O_285,N_3075,N_3858);
nor UO_286 (O_286,N_4880,N_3501);
nor UO_287 (O_287,N_2743,N_3739);
nand UO_288 (O_288,N_4663,N_4011);
nor UO_289 (O_289,N_4587,N_3009);
and UO_290 (O_290,N_4654,N_4942);
nor UO_291 (O_291,N_2612,N_3837);
nand UO_292 (O_292,N_3401,N_3301);
and UO_293 (O_293,N_2916,N_2839);
and UO_294 (O_294,N_4130,N_4290);
nor UO_295 (O_295,N_4129,N_2926);
nand UO_296 (O_296,N_4688,N_4769);
nand UO_297 (O_297,N_3361,N_2795);
and UO_298 (O_298,N_2886,N_2692);
or UO_299 (O_299,N_4836,N_3755);
nor UO_300 (O_300,N_4582,N_3978);
nand UO_301 (O_301,N_3149,N_3437);
nand UO_302 (O_302,N_3162,N_4247);
or UO_303 (O_303,N_2850,N_4551);
and UO_304 (O_304,N_3950,N_2532);
or UO_305 (O_305,N_4225,N_4366);
or UO_306 (O_306,N_4029,N_3111);
nand UO_307 (O_307,N_3567,N_2676);
nand UO_308 (O_308,N_4116,N_3533);
nand UO_309 (O_309,N_3543,N_3166);
or UO_310 (O_310,N_4593,N_4434);
and UO_311 (O_311,N_3434,N_2559);
nor UO_312 (O_312,N_2740,N_2697);
or UO_313 (O_313,N_4140,N_4105);
nand UO_314 (O_314,N_3347,N_4612);
nor UO_315 (O_315,N_3128,N_4321);
nor UO_316 (O_316,N_4275,N_3575);
xnor UO_317 (O_317,N_3292,N_3190);
or UO_318 (O_318,N_3081,N_4224);
and UO_319 (O_319,N_3628,N_3108);
or UO_320 (O_320,N_3386,N_2761);
nand UO_321 (O_321,N_3675,N_4263);
nor UO_322 (O_322,N_3430,N_2863);
or UO_323 (O_323,N_3378,N_4989);
nand UO_324 (O_324,N_3085,N_3473);
or UO_325 (O_325,N_3605,N_3819);
nor UO_326 (O_326,N_4665,N_3702);
nand UO_327 (O_327,N_2818,N_4580);
nand UO_328 (O_328,N_3335,N_3624);
nor UO_329 (O_329,N_4032,N_3127);
and UO_330 (O_330,N_4843,N_4460);
and UO_331 (O_331,N_4365,N_4892);
nor UO_332 (O_332,N_3654,N_4109);
or UO_333 (O_333,N_3168,N_4687);
nor UO_334 (O_334,N_4682,N_3297);
nand UO_335 (O_335,N_2598,N_4573);
or UO_336 (O_336,N_3666,N_4052);
nand UO_337 (O_337,N_2555,N_4204);
nand UO_338 (O_338,N_4835,N_2922);
nand UO_339 (O_339,N_4645,N_3983);
xor UO_340 (O_340,N_3969,N_3816);
and UO_341 (O_341,N_4019,N_4478);
or UO_342 (O_342,N_3846,N_3770);
nand UO_343 (O_343,N_3021,N_2544);
nand UO_344 (O_344,N_4101,N_3833);
nor UO_345 (O_345,N_2691,N_4776);
or UO_346 (O_346,N_3038,N_4376);
nand UO_347 (O_347,N_3142,N_4933);
nor UO_348 (O_348,N_3269,N_3217);
and UO_349 (O_349,N_4486,N_3542);
nor UO_350 (O_350,N_4304,N_3522);
nor UO_351 (O_351,N_3911,N_3758);
nor UO_352 (O_352,N_3165,N_4114);
or UO_353 (O_353,N_2630,N_3649);
or UO_354 (O_354,N_2633,N_4357);
or UO_355 (O_355,N_2894,N_3189);
or UO_356 (O_356,N_4213,N_3711);
or UO_357 (O_357,N_2806,N_4323);
nand UO_358 (O_358,N_3467,N_2893);
nand UO_359 (O_359,N_4166,N_3648);
and UO_360 (O_360,N_2814,N_2828);
or UO_361 (O_361,N_2870,N_3450);
or UO_362 (O_362,N_3416,N_4519);
nand UO_363 (O_363,N_2573,N_4739);
or UO_364 (O_364,N_4901,N_2785);
or UO_365 (O_365,N_3380,N_4394);
nor UO_366 (O_366,N_3774,N_4962);
nor UO_367 (O_367,N_2864,N_3892);
or UO_368 (O_368,N_3387,N_2945);
xor UO_369 (O_369,N_4856,N_3084);
or UO_370 (O_370,N_4360,N_4380);
nor UO_371 (O_371,N_4355,N_4235);
and UO_372 (O_372,N_3222,N_4634);
or UO_373 (O_373,N_2535,N_2989);
and UO_374 (O_374,N_3053,N_3785);
nand UO_375 (O_375,N_2694,N_4296);
nand UO_376 (O_376,N_2749,N_4202);
nor UO_377 (O_377,N_3050,N_3126);
and UO_378 (O_378,N_3052,N_4523);
or UO_379 (O_379,N_2938,N_4656);
or UO_380 (O_380,N_4054,N_4070);
xnor UO_381 (O_381,N_4879,N_3998);
nand UO_382 (O_382,N_3068,N_4735);
and UO_383 (O_383,N_4680,N_3464);
and UO_384 (O_384,N_3570,N_4887);
nor UO_385 (O_385,N_4638,N_4009);
nand UO_386 (O_386,N_4705,N_4045);
or UO_387 (O_387,N_2912,N_3049);
and UO_388 (O_388,N_4489,N_3214);
nand UO_389 (O_389,N_2963,N_3712);
and UO_390 (O_390,N_3714,N_3413);
nor UO_391 (O_391,N_3556,N_4004);
nand UO_392 (O_392,N_4649,N_3923);
nand UO_393 (O_393,N_3375,N_3280);
nor UO_394 (O_394,N_3728,N_4624);
nor UO_395 (O_395,N_3538,N_2838);
nor UO_396 (O_396,N_3171,N_3272);
and UO_397 (O_397,N_3402,N_2735);
nand UO_398 (O_398,N_3606,N_3504);
nor UO_399 (O_399,N_2621,N_4524);
or UO_400 (O_400,N_4066,N_4326);
or UO_401 (O_401,N_4145,N_2576);
and UO_402 (O_402,N_4057,N_3938);
or UO_403 (O_403,N_3227,N_3365);
nor UO_404 (O_404,N_2770,N_4384);
and UO_405 (O_405,N_3034,N_3302);
nor UO_406 (O_406,N_2589,N_2804);
nand UO_407 (O_407,N_4137,N_3920);
nand UO_408 (O_408,N_3157,N_2877);
nand UO_409 (O_409,N_3657,N_2647);
and UO_410 (O_410,N_2736,N_2636);
xnor UO_411 (O_411,N_4164,N_3701);
or UO_412 (O_412,N_4511,N_3895);
or UO_413 (O_413,N_3276,N_4985);
and UO_414 (O_414,N_3462,N_3587);
nor UO_415 (O_415,N_4424,N_2888);
nor UO_416 (O_416,N_4787,N_3757);
and UO_417 (O_417,N_4340,N_2706);
nand UO_418 (O_418,N_4889,N_4317);
or UO_419 (O_419,N_3060,N_4946);
nor UO_420 (O_420,N_3116,N_4502);
and UO_421 (O_421,N_4123,N_3457);
nor UO_422 (O_422,N_4189,N_4614);
nand UO_423 (O_423,N_4249,N_3988);
and UO_424 (O_424,N_3486,N_3993);
nor UO_425 (O_425,N_4849,N_4627);
and UO_426 (O_426,N_2855,N_3775);
or UO_427 (O_427,N_4972,N_4198);
and UO_428 (O_428,N_4866,N_3254);
nand UO_429 (O_429,N_3131,N_3414);
or UO_430 (O_430,N_2891,N_4535);
and UO_431 (O_431,N_4346,N_4919);
nand UO_432 (O_432,N_3281,N_4848);
nand UO_433 (O_433,N_2715,N_4272);
and UO_434 (O_434,N_3505,N_3103);
or UO_435 (O_435,N_4526,N_3507);
or UO_436 (O_436,N_3762,N_3139);
and UO_437 (O_437,N_3460,N_4269);
xor UO_438 (O_438,N_3940,N_3443);
and UO_439 (O_439,N_4999,N_3435);
nand UO_440 (O_440,N_3715,N_4978);
nand UO_441 (O_441,N_4487,N_3445);
and UO_442 (O_442,N_4490,N_4466);
nor UO_443 (O_443,N_4968,N_4957);
and UO_444 (O_444,N_3913,N_2654);
and UO_445 (O_445,N_4883,N_4099);
nand UO_446 (O_446,N_3667,N_4221);
and UO_447 (O_447,N_4533,N_4058);
or UO_448 (O_448,N_4874,N_3067);
nand UO_449 (O_449,N_2846,N_2648);
or UO_450 (O_450,N_3530,N_4259);
xor UO_451 (O_451,N_2959,N_3794);
nor UO_452 (O_452,N_3331,N_3847);
and UO_453 (O_453,N_4470,N_4852);
nand UO_454 (O_454,N_4568,N_3366);
nand UO_455 (O_455,N_4353,N_2718);
or UO_456 (O_456,N_4763,N_2698);
and UO_457 (O_457,N_4098,N_3733);
and UO_458 (O_458,N_4352,N_3664);
or UO_459 (O_459,N_4616,N_4703);
nand UO_460 (O_460,N_4162,N_4393);
or UO_461 (O_461,N_3448,N_2913);
or UO_462 (O_462,N_2527,N_3825);
nand UO_463 (O_463,N_4062,N_2502);
nor UO_464 (O_464,N_4017,N_3955);
nor UO_465 (O_465,N_3480,N_2523);
nor UO_466 (O_466,N_3568,N_4652);
nand UO_467 (O_467,N_3540,N_2831);
nor UO_468 (O_468,N_3193,N_3521);
nand UO_469 (O_469,N_3838,N_3372);
and UO_470 (O_470,N_4421,N_3680);
or UO_471 (O_471,N_4694,N_4882);
nand UO_472 (O_472,N_2880,N_3278);
nand UO_473 (O_473,N_4006,N_4197);
nand UO_474 (O_474,N_2520,N_3544);
or UO_475 (O_475,N_3252,N_3814);
nand UO_476 (O_476,N_3707,N_3351);
nand UO_477 (O_477,N_4374,N_2829);
or UO_478 (O_478,N_4379,N_3922);
and UO_479 (O_479,N_3828,N_3874);
nor UO_480 (O_480,N_3529,N_2597);
or UO_481 (O_481,N_4512,N_4902);
and UO_482 (O_482,N_3520,N_2998);
nand UO_483 (O_483,N_2611,N_4970);
or UO_484 (O_484,N_4726,N_4007);
or UO_485 (O_485,N_3916,N_3289);
and UO_486 (O_486,N_4136,N_3840);
and UO_487 (O_487,N_4169,N_3133);
or UO_488 (O_488,N_4456,N_2610);
and UO_489 (O_489,N_4133,N_2817);
and UO_490 (O_490,N_2518,N_4650);
or UO_491 (O_491,N_2541,N_4266);
and UO_492 (O_492,N_2931,N_4648);
and UO_493 (O_493,N_3808,N_3153);
and UO_494 (O_494,N_2991,N_3952);
or UO_495 (O_495,N_4911,N_4930);
nor UO_496 (O_496,N_4606,N_4951);
nand UO_497 (O_497,N_2703,N_3588);
and UO_498 (O_498,N_4684,N_4767);
nand UO_499 (O_499,N_3643,N_2739);
or UO_500 (O_500,N_3842,N_3862);
or UO_501 (O_501,N_4183,N_4610);
nor UO_502 (O_502,N_4039,N_4609);
nand UO_503 (O_503,N_3994,N_3897);
nor UO_504 (O_504,N_2949,N_4465);
or UO_505 (O_505,N_2788,N_3243);
and UO_506 (O_506,N_3599,N_4530);
and UO_507 (O_507,N_4555,N_3658);
and UO_508 (O_508,N_2972,N_4218);
nand UO_509 (O_509,N_4576,N_4168);
or UO_510 (O_510,N_3592,N_3184);
nand UO_511 (O_511,N_2667,N_2808);
or UO_512 (O_512,N_2526,N_4153);
or UO_513 (O_513,N_4932,N_3264);
or UO_514 (O_514,N_2865,N_3427);
nand UO_515 (O_515,N_2764,N_3783);
nor UO_516 (O_516,N_4396,N_3693);
nand UO_517 (O_517,N_3226,N_4833);
and UO_518 (O_518,N_4256,N_4842);
nor UO_519 (O_519,N_4716,N_3857);
nor UO_520 (O_520,N_3470,N_4031);
nor UO_521 (O_521,N_4876,N_4553);
nor UO_522 (O_522,N_3685,N_2678);
and UO_523 (O_523,N_4370,N_2556);
and UO_524 (O_524,N_4427,N_4994);
or UO_525 (O_525,N_4510,N_4035);
nor UO_526 (O_526,N_4329,N_3782);
or UO_527 (O_527,N_4063,N_4881);
nand UO_528 (O_528,N_3909,N_4818);
or UO_529 (O_529,N_4078,N_4826);
or UO_530 (O_530,N_3270,N_3789);
or UO_531 (O_531,N_3123,N_3221);
and UO_532 (O_532,N_4347,N_4659);
nand UO_533 (O_533,N_3653,N_4024);
or UO_534 (O_534,N_4834,N_2910);
nand UO_535 (O_535,N_3990,N_4237);
or UO_536 (O_536,N_4863,N_4661);
or UO_537 (O_537,N_4496,N_3390);
or UO_538 (O_538,N_4113,N_2564);
and UO_539 (O_539,N_3633,N_4328);
or UO_540 (O_540,N_3322,N_4367);
xnor UO_541 (O_541,N_3793,N_4907);
and UO_542 (O_542,N_3971,N_3072);
and UO_543 (O_543,N_2859,N_3866);
nand UO_544 (O_544,N_2536,N_4128);
or UO_545 (O_545,N_3531,N_4897);
nand UO_546 (O_546,N_3225,N_4761);
or UO_547 (O_547,N_3056,N_3468);
nor UO_548 (O_548,N_3163,N_2805);
or UO_549 (O_549,N_3722,N_2957);
nor UO_550 (O_550,N_4205,N_4158);
and UO_551 (O_551,N_3781,N_3638);
or UO_552 (O_552,N_3859,N_3688);
nor UO_553 (O_553,N_4303,N_4392);
xor UO_554 (O_554,N_4028,N_3485);
or UO_555 (O_555,N_3433,N_4179);
and UO_556 (O_556,N_4655,N_2699);
or UO_557 (O_557,N_3584,N_3776);
or UO_558 (O_558,N_4187,N_2733);
nand UO_559 (O_559,N_3548,N_4092);
and UO_560 (O_560,N_3803,N_3147);
nand UO_561 (O_561,N_4240,N_3399);
nand UO_562 (O_562,N_2689,N_4738);
xor UO_563 (O_563,N_4268,N_4230);
or UO_564 (O_564,N_3047,N_3740);
or UO_565 (O_565,N_3935,N_3391);
nor UO_566 (O_566,N_2605,N_3697);
nand UO_567 (O_567,N_4428,N_4678);
and UO_568 (O_568,N_3031,N_4429);
and UO_569 (O_569,N_4844,N_4773);
xor UO_570 (O_570,N_3082,N_4016);
and UO_571 (O_571,N_3569,N_3905);
nand UO_572 (O_572,N_2540,N_4377);
and UO_573 (O_573,N_2714,N_3809);
nand UO_574 (O_574,N_4765,N_3623);
or UO_575 (O_575,N_2554,N_3383);
nor UO_576 (O_576,N_4513,N_3246);
xnor UO_577 (O_577,N_3344,N_2745);
nand UO_578 (O_578,N_3687,N_3907);
and UO_579 (O_579,N_4601,N_3918);
and UO_580 (O_580,N_4702,N_2550);
nor UO_581 (O_581,N_2682,N_4905);
nand UO_582 (O_582,N_2656,N_4305);
nor UO_583 (O_583,N_4527,N_2790);
or UO_584 (O_584,N_3580,N_3419);
nand UO_585 (O_585,N_3294,N_4819);
and UO_586 (O_586,N_4239,N_4934);
or UO_587 (O_587,N_4839,N_4977);
nand UO_588 (O_588,N_4809,N_2841);
or UO_589 (O_589,N_4417,N_2709);
and UO_590 (O_590,N_4742,N_3245);
nor UO_591 (O_591,N_4721,N_4177);
nand UO_592 (O_592,N_4418,N_4288);
nand UO_593 (O_593,N_4444,N_4040);
and UO_594 (O_594,N_4660,N_4531);
or UO_595 (O_595,N_4845,N_3886);
nor UO_596 (O_596,N_4749,N_2896);
or UO_597 (O_597,N_4562,N_2917);
or UO_598 (O_598,N_4121,N_3871);
and UO_599 (O_599,N_4482,N_4074);
or UO_600 (O_600,N_2680,N_4291);
and UO_601 (O_601,N_3564,N_4043);
and UO_602 (O_602,N_4560,N_3812);
or UO_603 (O_603,N_2942,N_3929);
nor UO_604 (O_604,N_4781,N_3395);
or UO_605 (O_605,N_3211,N_4828);
nand UO_606 (O_606,N_3369,N_2780);
xnor UO_607 (O_607,N_3927,N_4412);
or UO_608 (O_608,N_3829,N_3954);
and UO_609 (O_609,N_3945,N_2710);
and UO_610 (O_610,N_3234,N_3459);
and UO_611 (O_611,N_4789,N_2686);
xor UO_612 (O_612,N_3786,N_4973);
and UO_613 (O_613,N_4222,N_4072);
nand UO_614 (O_614,N_4003,N_4559);
and UO_615 (O_615,N_2504,N_3818);
nor UO_616 (O_616,N_3398,N_3230);
or UO_617 (O_617,N_3140,N_3705);
nor UO_618 (O_618,N_3336,N_4157);
nor UO_619 (O_619,N_4633,N_3400);
nor UO_620 (O_620,N_2809,N_4142);
or UO_621 (O_621,N_4325,N_4910);
and UO_622 (O_622,N_3513,N_4941);
and UO_623 (O_623,N_3491,N_3120);
or UO_624 (O_624,N_2881,N_4823);
nor UO_625 (O_625,N_4134,N_2707);
nor UO_626 (O_626,N_4707,N_3478);
xor UO_627 (O_627,N_3749,N_2889);
and UO_628 (O_628,N_3609,N_2507);
nor UO_629 (O_629,N_4617,N_4371);
and UO_630 (O_630,N_2644,N_4629);
and UO_631 (O_631,N_3354,N_2897);
nor UO_632 (O_632,N_3323,N_3704);
and UO_633 (O_633,N_4651,N_3676);
xor UO_634 (O_634,N_4425,N_3659);
and UO_635 (O_635,N_3349,N_4775);
or UO_636 (O_636,N_3834,N_4061);
or UO_637 (O_637,N_2675,N_4008);
nor UO_638 (O_638,N_2854,N_4673);
and UO_639 (O_639,N_3741,N_4683);
and UO_640 (O_640,N_2537,N_4322);
nand UO_641 (O_641,N_2967,N_3939);
and UO_642 (O_642,N_2997,N_2951);
and UO_643 (O_643,N_4734,N_3196);
and UO_644 (O_644,N_4595,N_4499);
and UO_645 (O_645,N_4805,N_4552);
nand UO_646 (O_646,N_4102,N_2620);
or UO_647 (O_647,N_3982,N_3282);
nand UO_648 (O_648,N_2596,N_3219);
or UO_649 (O_649,N_4744,N_2907);
nand UO_650 (O_650,N_2878,N_4886);
and UO_651 (O_651,N_3397,N_3989);
or UO_652 (O_652,N_4918,N_4548);
or UO_653 (O_653,N_3432,N_4124);
and UO_654 (O_654,N_4817,N_4319);
or UO_655 (O_655,N_3195,N_4637);
nand UO_656 (O_656,N_2562,N_2669);
nor UO_657 (O_657,N_4415,N_4671);
and UO_658 (O_658,N_3074,N_3477);
nand UO_659 (O_659,N_4459,N_3138);
nand UO_660 (O_660,N_2960,N_3937);
xnor UO_661 (O_661,N_4163,N_4597);
or UO_662 (O_662,N_3170,N_4750);
nor UO_663 (O_663,N_2819,N_2587);
and UO_664 (O_664,N_4318,N_4174);
or UO_665 (O_665,N_4717,N_4358);
and UO_666 (O_666,N_3422,N_4494);
nand UO_667 (O_667,N_2567,N_3376);
and UO_668 (O_668,N_4563,N_4875);
and UO_669 (O_669,N_3967,N_3356);
and UO_670 (O_670,N_3593,N_4345);
nor UO_671 (O_671,N_4945,N_3578);
nand UO_672 (O_672,N_3632,N_4161);
nand UO_673 (O_673,N_4297,N_2655);
nand UO_674 (O_674,N_4073,N_3241);
or UO_675 (O_675,N_3132,N_4284);
xor UO_676 (O_676,N_3549,N_4709);
nor UO_677 (O_677,N_2924,N_3602);
and UO_678 (O_678,N_3534,N_3300);
nor UO_679 (O_679,N_3537,N_4988);
nor UO_680 (O_680,N_4013,N_3186);
nand UO_681 (O_681,N_4090,N_2650);
or UO_682 (O_682,N_4250,N_4708);
nand UO_683 (O_683,N_4539,N_2705);
nor UO_684 (O_684,N_4208,N_3035);
and UO_685 (O_685,N_2625,N_4662);
nand UO_686 (O_686,N_4859,N_3385);
or UO_687 (O_687,N_2851,N_3600);
nand UO_688 (O_688,N_4646,N_4302);
nand UO_689 (O_689,N_3872,N_3492);
nor UO_690 (O_690,N_4693,N_3094);
nor UO_691 (O_691,N_3497,N_4575);
nand UO_692 (O_692,N_2533,N_3203);
xor UO_693 (O_693,N_4279,N_2510);
or UO_694 (O_694,N_2717,N_4018);
nand UO_695 (O_695,N_3824,N_4643);
and UO_696 (O_696,N_3090,N_4282);
nand UO_697 (O_697,N_3439,N_4712);
and UO_698 (O_698,N_4772,N_4132);
nor UO_699 (O_699,N_3309,N_4640);
nor UO_700 (O_700,N_3779,N_3188);
nor UO_701 (O_701,N_2666,N_2940);
or UO_702 (O_702,N_4855,N_3512);
and UO_703 (O_703,N_2734,N_2852);
nand UO_704 (O_704,N_3579,N_4056);
nor UO_705 (O_705,N_3801,N_3089);
or UO_706 (O_706,N_3903,N_4953);
nor UO_707 (O_707,N_3005,N_3721);
nand UO_708 (O_708,N_4096,N_4089);
or UO_709 (O_709,N_4375,N_4049);
nand UO_710 (O_710,N_2542,N_4748);
or UO_711 (O_711,N_3975,N_4518);
nor UO_712 (O_712,N_4186,N_4871);
and UO_713 (O_713,N_3679,N_2748);
or UO_714 (O_714,N_3619,N_4423);
and UO_715 (O_715,N_3172,N_4589);
nor UO_716 (O_716,N_2868,N_4537);
or UO_717 (O_717,N_3291,N_2570);
or UO_718 (O_718,N_4484,N_4658);
nand UO_719 (O_719,N_3065,N_3759);
or UO_720 (O_720,N_4790,N_3426);
or UO_721 (O_721,N_3223,N_3516);
nor UO_722 (O_722,N_3729,N_4588);
nand UO_723 (O_723,N_4532,N_3310);
or UO_724 (O_724,N_3048,N_4832);
nand UO_725 (O_725,N_4244,N_3646);
or UO_726 (O_726,N_4246,N_3087);
nor UO_727 (O_727,N_4196,N_3613);
and UO_728 (O_728,N_2929,N_3698);
and UO_729 (O_729,N_3080,N_3947);
nand UO_730 (O_730,N_2982,N_2939);
or UO_731 (O_731,N_3831,N_4768);
nor UO_732 (O_732,N_2607,N_3317);
or UO_733 (O_733,N_3412,N_3338);
and UO_734 (O_734,N_3161,N_3962);
nand UO_735 (O_735,N_4432,N_2565);
nand UO_736 (O_736,N_4248,N_4824);
or UO_737 (O_737,N_4695,N_4257);
or UO_738 (O_738,N_2980,N_2918);
nor UO_739 (O_739,N_4746,N_3748);
nor UO_740 (O_740,N_2801,N_4372);
and UO_741 (O_741,N_3763,N_3061);
or UO_742 (O_742,N_3192,N_3753);
nand UO_743 (O_743,N_4668,N_2659);
nand UO_744 (O_744,N_4433,N_4270);
nand UO_745 (O_745,N_4468,N_3357);
or UO_746 (O_746,N_3682,N_4503);
or UO_747 (O_747,N_4278,N_3949);
and UO_748 (O_748,N_3565,N_4287);
nor UO_749 (O_749,N_4691,N_4625);
nand UO_750 (O_750,N_4755,N_4405);
nor UO_751 (O_751,N_3979,N_3212);
or UO_752 (O_752,N_3410,N_3122);
and UO_753 (O_753,N_3904,N_4354);
nor UO_754 (O_754,N_4311,N_3641);
and UO_755 (O_755,N_3063,N_2937);
and UO_756 (O_756,N_2930,N_3614);
nand UO_757 (O_757,N_3025,N_4395);
nor UO_758 (O_758,N_4622,N_4898);
or UO_759 (O_759,N_3411,N_4853);
nand UO_760 (O_760,N_3232,N_3070);
nor UO_761 (O_761,N_3431,N_2976);
nand UO_762 (O_762,N_4422,N_3236);
or UO_763 (O_763,N_4723,N_2702);
nor UO_764 (O_764,N_4800,N_4294);
and UO_765 (O_765,N_2646,N_4685);
or UO_766 (O_766,N_2701,N_2738);
or UO_767 (O_767,N_3924,N_3761);
and UO_768 (O_768,N_3008,N_2983);
or UO_769 (O_769,N_3191,N_4001);
and UO_770 (O_770,N_3384,N_3350);
nor UO_771 (O_771,N_4998,N_2794);
nor UO_772 (O_772,N_3145,N_2946);
and UO_773 (O_773,N_3327,N_2958);
nand UO_774 (O_774,N_3407,N_4704);
nor UO_775 (O_775,N_4940,N_4348);
or UO_776 (O_776,N_4598,N_2730);
nor UO_777 (O_777,N_4104,N_4083);
nand UO_778 (O_778,N_4632,N_4931);
and UO_779 (O_779,N_2911,N_2756);
nor UO_780 (O_780,N_2727,N_4557);
nand UO_781 (O_781,N_4865,N_4261);
or UO_782 (O_782,N_2668,N_3820);
or UO_783 (O_783,N_4310,N_4774);
nor UO_784 (O_784,N_2832,N_3083);
nor UO_785 (O_785,N_4149,N_4724);
or UO_786 (O_786,N_2519,N_3154);
and UO_787 (O_787,N_3263,N_4075);
nor UO_788 (O_788,N_3324,N_4403);
and UO_789 (O_789,N_2970,N_3438);
xor UO_790 (O_790,N_2823,N_4505);
and UO_791 (O_791,N_3334,N_4944);
and UO_792 (O_792,N_4647,N_4784);
and UO_793 (O_793,N_4778,N_4474);
and UO_794 (O_794,N_4677,N_3612);
nand UO_795 (O_795,N_2747,N_4065);
nor UO_796 (O_796,N_4592,N_3167);
and UO_797 (O_797,N_4741,N_3815);
and UO_798 (O_798,N_3006,N_3091);
and UO_799 (O_799,N_2522,N_3303);
nand UO_800 (O_800,N_3737,N_4184);
nand UO_801 (O_801,N_4491,N_4426);
nor UO_802 (O_802,N_3255,N_3865);
and UO_803 (O_803,N_3421,N_3113);
nand UO_804 (O_804,N_2546,N_4829);
xnor UO_805 (O_805,N_2763,N_2690);
xnor UO_806 (O_806,N_3713,N_4464);
nor UO_807 (O_807,N_3121,N_3946);
nand UO_808 (O_808,N_2708,N_3640);
or UO_809 (O_809,N_3374,N_2956);
nor UO_810 (O_810,N_4271,N_2568);
or UO_811 (O_811,N_3011,N_4138);
or UO_812 (O_812,N_4012,N_2609);
and UO_813 (O_813,N_4458,N_3012);
or UO_814 (O_814,N_4908,N_4745);
or UO_815 (O_815,N_4388,N_3118);
and UO_816 (O_816,N_3273,N_4131);
and UO_817 (O_817,N_3039,N_3517);
or UO_818 (O_818,N_4262,N_3991);
nor UO_819 (O_819,N_2606,N_3764);
or UO_820 (O_820,N_4450,N_4308);
and UO_821 (O_821,N_3388,N_2581);
and UO_822 (O_822,N_3363,N_4565);
and UO_823 (O_823,N_4413,N_2992);
and UO_824 (O_824,N_4156,N_3028);
nor UO_825 (O_825,N_4336,N_3259);
nor UO_826 (O_826,N_3925,N_4926);
nor UO_827 (O_827,N_4176,N_4182);
nor UO_828 (O_828,N_4756,N_4200);
nor UO_829 (O_829,N_4591,N_3898);
nand UO_830 (O_830,N_3980,N_3472);
nor UO_831 (O_831,N_3835,N_3778);
nor UO_832 (O_832,N_3308,N_3095);
nor UO_833 (O_833,N_2771,N_3213);
nor UO_834 (O_834,N_3109,N_4408);
nand UO_835 (O_835,N_2954,N_2671);
or UO_836 (O_836,N_3956,N_4583);
and UO_837 (O_837,N_3525,N_2978);
xor UO_838 (O_838,N_3572,N_3651);
nor UO_839 (O_839,N_3148,N_3966);
nor UO_840 (O_840,N_4330,N_4437);
or UO_841 (O_841,N_4095,N_4231);
or UO_842 (O_842,N_4525,N_4949);
nand UO_843 (O_843,N_4219,N_4483);
and UO_844 (O_844,N_3134,N_4500);
nor UO_845 (O_845,N_3906,N_3736);
nor UO_846 (O_846,N_3856,N_2953);
nand UO_847 (O_847,N_4564,N_3231);
xor UO_848 (O_848,N_4689,N_4327);
and UO_849 (O_849,N_4160,N_4349);
nand UO_850 (O_850,N_3902,N_2525);
and UO_851 (O_851,N_3275,N_2783);
nor UO_852 (O_852,N_3493,N_4674);
nor UO_853 (O_853,N_3811,N_2996);
or UO_854 (O_854,N_4195,N_3017);
and UO_855 (O_855,N_3730,N_4293);
or UO_856 (O_856,N_2932,N_2603);
nor UO_857 (O_857,N_4967,N_2673);
and UO_858 (O_858,N_3207,N_4720);
nor UO_859 (O_859,N_4808,N_2862);
or UO_860 (O_860,N_4332,N_2962);
nand UO_861 (O_861,N_3125,N_4167);
or UO_862 (O_862,N_2769,N_4082);
and UO_863 (O_863,N_2538,N_3742);
and UO_864 (O_864,N_4436,N_3362);
nor UO_865 (O_865,N_4731,N_4796);
nor UO_866 (O_866,N_2776,N_2530);
nor UO_867 (O_867,N_3700,N_3428);
nor UO_868 (O_868,N_3558,N_4341);
nand UO_869 (O_869,N_4026,N_2506);
nand UO_870 (O_870,N_4443,N_4759);
and UO_871 (O_871,N_3326,N_2887);
nor UO_872 (O_872,N_4097,N_4245);
nand UO_873 (O_873,N_3621,N_2543);
or UO_874 (O_874,N_2744,N_4786);
nand UO_875 (O_875,N_4320,N_3110);
nand UO_876 (O_876,N_4758,N_2973);
nand UO_877 (O_877,N_2810,N_4554);
xor UO_878 (O_878,N_3341,N_4171);
nor UO_879 (O_879,N_2964,N_2547);
and UO_880 (O_880,N_3546,N_4501);
nor UO_881 (O_881,N_2732,N_3102);
xor UO_882 (O_882,N_3987,N_3373);
or UO_883 (O_883,N_3325,N_4106);
and UO_884 (O_884,N_3696,N_2857);
or UO_885 (O_885,N_3494,N_4605);
and UO_886 (O_886,N_2892,N_3174);
and UO_887 (O_887,N_3802,N_4821);
and UO_888 (O_888,N_2873,N_4298);
and UO_889 (O_889,N_3456,N_3634);
nand UO_890 (O_890,N_2622,N_3725);
nor UO_891 (O_891,N_4681,N_3247);
or UO_892 (O_892,N_4435,N_2746);
or UO_893 (O_893,N_2824,N_4891);
or UO_894 (O_894,N_3169,N_4584);
nor UO_895 (O_895,N_4449,N_3963);
or UO_896 (O_896,N_2975,N_4830);
nand UO_897 (O_897,N_4529,N_3671);
nor UO_898 (O_898,N_4243,N_3678);
or UO_899 (O_899,N_3394,N_3429);
nand UO_900 (O_900,N_3290,N_2563);
or UO_901 (O_901,N_4545,N_2586);
or UO_902 (O_902,N_3316,N_4342);
nand UO_903 (O_903,N_2638,N_2508);
nand UO_904 (O_904,N_4025,N_3441);
and UO_905 (O_905,N_2501,N_2849);
or UO_906 (O_906,N_4027,N_3124);
nor UO_907 (O_907,N_4267,N_4697);
and UO_908 (O_908,N_3526,N_4100);
or UO_909 (O_909,N_2712,N_3146);
nor UO_910 (O_910,N_4920,N_3894);
nand UO_911 (O_911,N_4937,N_4508);
nor UO_912 (O_912,N_3257,N_2993);
nand UO_913 (O_913,N_3321,N_3224);
nor UO_914 (O_914,N_2875,N_4363);
nor UO_915 (O_915,N_3342,N_2901);
nor UO_916 (O_916,N_3910,N_4265);
and UO_917 (O_917,N_4260,N_4807);
nand UO_918 (O_918,N_4440,N_4906);
nor UO_919 (O_919,N_2866,N_3765);
nor UO_920 (O_920,N_3446,N_4850);
or UO_921 (O_921,N_3114,N_2869);
or UO_922 (O_922,N_3948,N_3502);
or UO_923 (O_923,N_2987,N_4730);
nand UO_924 (O_924,N_3204,N_4696);
nor UO_925 (O_925,N_4927,N_3631);
nand UO_926 (O_926,N_3260,N_3650);
nor UO_927 (O_927,N_3007,N_3810);
nor UO_928 (O_928,N_3958,N_3244);
nor UO_929 (O_929,N_3792,N_3096);
or UO_930 (O_930,N_3550,N_4399);
nor UO_931 (O_931,N_3747,N_3393);
and UO_932 (O_932,N_2683,N_4251);
nand UO_933 (O_933,N_4309,N_3098);
nor UO_934 (O_934,N_2812,N_4925);
or UO_935 (O_935,N_4306,N_3329);
and UO_936 (O_936,N_2952,N_2627);
nor UO_937 (O_937,N_4743,N_4077);
or UO_938 (O_938,N_3332,N_4666);
nand UO_939 (O_939,N_3843,N_4713);
nand UO_940 (O_940,N_4185,N_3469);
nand UO_941 (O_941,N_3844,N_3059);
nand UO_942 (O_942,N_2833,N_3043);
or UO_943 (O_943,N_3890,N_4547);
nor UO_944 (O_944,N_4538,N_4036);
or UO_945 (O_945,N_3175,N_4276);
nand UO_946 (O_946,N_3662,N_3891);
nand UO_947 (O_947,N_4110,N_3683);
nand UO_948 (O_948,N_4414,N_3041);
and UO_949 (O_949,N_3545,N_3636);
or UO_950 (O_950,N_3888,N_2803);
and UO_951 (O_951,N_3220,N_2741);
nor UO_952 (O_952,N_4959,N_2856);
nand UO_953 (O_953,N_4203,N_3689);
or UO_954 (O_954,N_2934,N_3487);
nor UO_955 (O_955,N_2662,N_2830);
nand UO_956 (O_956,N_2923,N_2728);
nand UO_957 (O_957,N_2915,N_3135);
nor UO_958 (O_958,N_3849,N_4223);
and UO_959 (O_959,N_2928,N_3848);
and UO_960 (O_960,N_3285,N_4473);
nand UO_961 (O_961,N_3527,N_3253);
or UO_962 (O_962,N_3582,N_4258);
nor UO_963 (O_963,N_4870,N_2903);
nand UO_964 (O_964,N_3265,N_3618);
and UO_965 (O_965,N_4192,N_4812);
nor UO_966 (O_966,N_3496,N_4635);
nand UO_967 (O_967,N_4923,N_2822);
or UO_968 (O_968,N_3900,N_3941);
nor UO_969 (O_969,N_3893,N_2512);
or UO_970 (O_970,N_3626,N_3305);
nand UO_971 (O_971,N_2591,N_2908);
nand UO_972 (O_972,N_4350,N_3622);
and UO_973 (O_973,N_4021,N_4252);
and UO_974 (O_974,N_4822,N_2599);
nand UO_975 (O_975,N_4014,N_2936);
nand UO_976 (O_976,N_2687,N_2719);
and UO_977 (O_977,N_4236,N_2778);
and UO_978 (O_978,N_2608,N_3256);
or UO_979 (O_979,N_2503,N_3665);
nor UO_980 (O_980,N_4280,N_3772);
xnor UO_981 (O_981,N_4264,N_3559);
nor UO_982 (O_982,N_3630,N_3574);
nand UO_983 (O_983,N_2906,N_3498);
or UO_984 (O_984,N_3010,N_2787);
nor UO_985 (O_985,N_3581,N_3876);
nor UO_986 (O_986,N_3353,N_4234);
nand UO_987 (O_987,N_3396,N_2802);
and UO_988 (O_988,N_3668,N_3037);
nand UO_989 (O_989,N_4992,N_4718);
and UO_990 (O_990,N_3181,N_3370);
nor UO_991 (O_991,N_4700,N_2628);
nor UO_992 (O_992,N_3708,N_2651);
and UO_993 (O_993,N_4740,N_2724);
or UO_994 (O_994,N_4664,N_4194);
nand UO_995 (O_995,N_4914,N_3870);
nor UO_996 (O_996,N_3655,N_4869);
nand UO_997 (O_997,N_3723,N_3601);
and UO_998 (O_998,N_4515,N_4079);
nand UO_999 (O_999,N_4467,N_4112);
endmodule