module basic_1500_15000_2000_15_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_75,In_901);
nor U1 (N_1,In_1182,In_364);
xor U2 (N_2,In_694,In_1377);
xor U3 (N_3,In_197,In_740);
or U4 (N_4,In_351,In_1275);
nor U5 (N_5,In_1080,In_1252);
or U6 (N_6,In_841,In_82);
nor U7 (N_7,In_46,In_398);
and U8 (N_8,In_1142,In_666);
nor U9 (N_9,In_550,In_982);
nand U10 (N_10,In_1257,In_689);
and U11 (N_11,In_1165,In_899);
xor U12 (N_12,In_498,In_1357);
or U13 (N_13,In_566,In_1331);
or U14 (N_14,In_332,In_1179);
xnor U15 (N_15,In_1204,In_97);
nand U16 (N_16,In_80,In_1428);
and U17 (N_17,In_862,In_651);
or U18 (N_18,In_308,In_409);
xor U19 (N_19,In_1405,In_1249);
and U20 (N_20,In_1020,In_174);
nand U21 (N_21,In_630,In_451);
and U22 (N_22,In_372,In_1227);
nand U23 (N_23,In_130,In_1255);
xor U24 (N_24,In_1395,In_1351);
nor U25 (N_25,In_1030,In_1373);
xor U26 (N_26,In_450,In_1430);
or U27 (N_27,In_792,In_500);
nor U28 (N_28,In_229,In_713);
nor U29 (N_29,In_261,In_331);
or U30 (N_30,In_17,In_1233);
and U31 (N_31,In_290,In_1102);
nand U32 (N_32,In_1475,In_449);
or U33 (N_33,In_984,In_262);
nand U34 (N_34,In_503,In_1374);
xor U35 (N_35,In_1322,In_1301);
nand U36 (N_36,In_499,In_359);
nand U37 (N_37,In_416,In_399);
nand U38 (N_38,In_1041,In_947);
nand U39 (N_39,In_1113,In_608);
xnor U40 (N_40,In_168,In_1202);
nor U41 (N_41,In_686,In_246);
nor U42 (N_42,In_1158,In_752);
or U43 (N_43,In_173,In_88);
nor U44 (N_44,In_784,In_693);
nand U45 (N_45,In_1467,In_132);
and U46 (N_46,In_188,In_478);
nor U47 (N_47,In_28,In_487);
or U48 (N_48,In_827,In_417);
nor U49 (N_49,In_1262,In_124);
and U50 (N_50,In_1219,In_381);
nor U51 (N_51,In_18,In_821);
nand U52 (N_52,In_489,In_1008);
and U53 (N_53,In_415,In_1185);
or U54 (N_54,In_454,In_574);
nor U55 (N_55,In_872,In_853);
and U56 (N_56,In_155,In_542);
or U57 (N_57,In_7,In_1332);
nor U58 (N_58,In_881,In_126);
xnor U59 (N_59,In_1250,In_425);
nor U60 (N_60,In_373,In_483);
and U61 (N_61,In_886,In_908);
or U62 (N_62,In_981,In_65);
or U63 (N_63,In_120,In_1366);
or U64 (N_64,In_1324,In_625);
xnor U65 (N_65,In_1263,In_800);
xnor U66 (N_66,In_675,In_996);
nor U67 (N_67,In_1011,In_418);
and U68 (N_68,In_780,In_1264);
and U69 (N_69,In_588,In_851);
xnor U70 (N_70,In_979,In_1378);
and U71 (N_71,In_941,In_723);
xnor U72 (N_72,In_594,In_907);
xnor U73 (N_73,In_997,In_523);
and U74 (N_74,In_179,In_254);
nand U75 (N_75,In_597,In_42);
nand U76 (N_76,In_1025,In_1003);
and U77 (N_77,In_32,In_443);
xnor U78 (N_78,In_718,In_534);
nand U79 (N_79,In_1333,In_1198);
nand U80 (N_80,In_1084,In_255);
nor U81 (N_81,In_1120,In_598);
or U82 (N_82,In_833,In_1069);
or U83 (N_83,In_8,In_115);
or U84 (N_84,In_257,In_1138);
nor U85 (N_85,In_1046,In_730);
or U86 (N_86,In_387,In_1468);
nand U87 (N_87,In_445,In_196);
nor U88 (N_88,In_338,In_326);
nor U89 (N_89,In_864,In_739);
xnor U90 (N_90,In_31,In_61);
or U91 (N_91,In_1319,In_567);
xnor U92 (N_92,In_528,In_538);
xor U93 (N_93,In_1391,In_1444);
and U94 (N_94,In_463,In_1190);
nand U95 (N_95,In_758,In_751);
nor U96 (N_96,In_696,In_754);
and U97 (N_97,In_312,In_43);
nor U98 (N_98,In_81,In_178);
or U99 (N_99,In_1099,In_1037);
nand U100 (N_100,In_295,In_1174);
and U101 (N_101,In_1300,In_1439);
or U102 (N_102,In_47,In_1028);
xor U103 (N_103,In_100,In_735);
xnor U104 (N_104,In_1443,In_1001);
or U105 (N_105,In_223,In_1404);
xor U106 (N_106,In_104,In_1140);
xor U107 (N_107,In_755,In_185);
nand U108 (N_108,In_1387,In_1419);
nor U109 (N_109,In_476,In_243);
and U110 (N_110,In_1336,In_5);
nor U111 (N_111,In_1100,In_339);
nor U112 (N_112,In_45,In_1075);
nor U113 (N_113,In_335,In_1317);
nor U114 (N_114,In_839,In_1045);
nor U115 (N_115,In_12,In_551);
nor U116 (N_116,In_820,In_1335);
xnor U117 (N_117,In_946,In_685);
or U118 (N_118,In_1242,In_1039);
nor U119 (N_119,In_461,In_508);
nor U120 (N_120,In_584,In_1031);
and U121 (N_121,In_1215,In_1464);
or U122 (N_122,In_1083,In_766);
and U123 (N_123,In_802,In_1406);
or U124 (N_124,In_634,In_583);
nand U125 (N_125,In_1426,In_1368);
nor U126 (N_126,In_59,In_638);
nand U127 (N_127,In_1407,In_1296);
and U128 (N_128,In_239,In_627);
nand U129 (N_129,In_281,In_158);
nand U130 (N_130,In_900,In_880);
or U131 (N_131,In_1265,In_562);
nand U132 (N_132,In_378,In_887);
nor U133 (N_133,In_1266,In_55);
or U134 (N_134,In_1445,In_1055);
nand U135 (N_135,In_1048,In_580);
nand U136 (N_136,In_682,In_114);
and U137 (N_137,In_1390,In_96);
nor U138 (N_138,In_218,In_671);
and U139 (N_139,In_1189,In_260);
xor U140 (N_140,In_1306,In_1096);
nor U141 (N_141,In_436,In_960);
nand U142 (N_142,In_324,In_355);
xnor U143 (N_143,In_1431,In_1297);
nand U144 (N_144,In_122,In_1143);
or U145 (N_145,In_533,In_940);
nand U146 (N_146,In_1081,In_863);
or U147 (N_147,In_29,In_605);
and U148 (N_148,In_1343,In_1114);
nand U149 (N_149,In_383,In_1139);
xor U150 (N_150,In_1329,In_1168);
nand U151 (N_151,In_782,In_41);
nand U152 (N_152,In_1375,In_441);
xor U153 (N_153,In_150,In_1002);
nor U154 (N_154,In_1438,In_1471);
nand U155 (N_155,In_184,In_622);
xor U156 (N_156,In_725,In_1454);
nor U157 (N_157,In_456,In_1320);
nand U158 (N_158,In_1321,In_787);
and U159 (N_159,In_1187,In_658);
and U160 (N_160,In_1078,In_560);
and U161 (N_161,In_592,In_1243);
and U162 (N_162,In_433,In_571);
and U163 (N_163,In_1434,In_1289);
nand U164 (N_164,In_706,In_1124);
nor U165 (N_165,In_395,In_657);
or U166 (N_166,In_1062,In_69);
or U167 (N_167,In_294,In_277);
nor U168 (N_168,In_505,In_1010);
or U169 (N_169,In_25,In_288);
or U170 (N_170,In_688,In_3);
nand U171 (N_171,In_342,In_206);
or U172 (N_172,In_585,In_895);
nand U173 (N_173,In_543,In_988);
or U174 (N_174,In_401,In_743);
and U175 (N_175,In_279,In_791);
nor U176 (N_176,In_426,In_1195);
and U177 (N_177,In_147,In_591);
or U178 (N_178,In_545,In_1497);
nor U179 (N_179,In_559,In_926);
or U180 (N_180,In_665,In_64);
nand U181 (N_181,In_131,In_181);
nand U182 (N_182,In_213,In_1276);
or U183 (N_183,In_526,In_889);
xnor U184 (N_184,In_157,In_1261);
xnor U185 (N_185,In_397,In_1418);
xnor U186 (N_186,In_1157,In_1286);
nand U187 (N_187,In_1207,In_840);
or U188 (N_188,In_1298,In_590);
xor U189 (N_189,In_1311,In_1386);
or U190 (N_190,In_1110,In_77);
or U191 (N_191,In_1108,In_1137);
or U192 (N_192,In_323,In_1006);
nand U193 (N_193,In_602,In_63);
xor U194 (N_194,In_492,In_193);
and U195 (N_195,In_915,In_1398);
nand U196 (N_196,In_1441,In_1117);
nand U197 (N_197,In_716,In_637);
and U198 (N_198,In_668,In_394);
nor U199 (N_199,In_662,In_1056);
and U200 (N_200,In_448,In_370);
and U201 (N_201,In_1291,In_452);
or U202 (N_202,In_1044,In_1194);
nor U203 (N_203,In_898,In_149);
nand U204 (N_204,In_1004,In_140);
nor U205 (N_205,In_139,In_110);
nor U206 (N_206,In_432,In_935);
nand U207 (N_207,In_1101,In_1016);
nor U208 (N_208,In_396,In_844);
or U209 (N_209,In_428,In_1068);
and U210 (N_210,In_275,In_764);
xor U211 (N_211,In_67,In_799);
and U212 (N_212,In_507,In_653);
xor U213 (N_213,In_1436,In_164);
nand U214 (N_214,In_530,In_1480);
or U215 (N_215,In_648,In_595);
nor U216 (N_216,In_890,In_210);
and U217 (N_217,In_1367,In_948);
nand U218 (N_218,In_1432,In_402);
nand U219 (N_219,In_965,In_756);
or U220 (N_220,In_111,In_711);
nand U221 (N_221,In_107,In_447);
nand U222 (N_222,In_582,In_1091);
and U223 (N_223,In_138,In_993);
and U224 (N_224,In_883,In_480);
nand U225 (N_225,In_731,In_990);
and U226 (N_226,In_712,In_340);
or U227 (N_227,In_330,In_44);
nor U228 (N_228,In_92,In_250);
nor U229 (N_229,In_525,In_519);
nor U230 (N_230,In_795,In_509);
nand U231 (N_231,In_897,In_116);
nor U232 (N_232,In_994,In_328);
xor U233 (N_233,In_876,In_913);
xnor U234 (N_234,In_976,In_1425);
and U235 (N_235,In_1489,In_23);
xnor U236 (N_236,In_283,In_646);
nor U237 (N_237,In_267,In_1032);
nand U238 (N_238,In_1022,In_609);
nand U239 (N_239,In_258,In_362);
or U240 (N_240,In_209,In_691);
xor U241 (N_241,In_1176,In_462);
or U242 (N_242,In_824,In_917);
or U243 (N_243,In_1036,In_1493);
xnor U244 (N_244,In_527,In_1192);
nor U245 (N_245,In_643,In_1180);
or U246 (N_246,In_143,In_640);
xnor U247 (N_247,In_645,In_217);
xnor U248 (N_248,In_842,In_248);
nor U249 (N_249,In_252,In_1433);
or U250 (N_250,In_199,In_327);
or U251 (N_251,In_1034,In_1244);
and U252 (N_252,In_734,In_785);
nor U253 (N_253,In_78,In_843);
nor U254 (N_254,In_442,In_249);
nand U255 (N_255,In_1225,In_1360);
xnor U256 (N_256,In_522,In_494);
and U257 (N_257,In_1167,In_1392);
xnor U258 (N_258,In_1087,In_977);
and U259 (N_259,In_537,In_1104);
and U260 (N_260,In_49,In_1007);
nand U261 (N_261,In_828,In_1183);
and U262 (N_262,In_269,In_1214);
xnor U263 (N_263,In_79,In_987);
nand U264 (N_264,In_375,In_825);
and U265 (N_265,In_1364,In_431);
and U266 (N_266,In_1248,In_1334);
xor U267 (N_267,In_957,In_729);
nor U268 (N_268,In_486,In_710);
nand U269 (N_269,In_816,In_1231);
nand U270 (N_270,In_105,In_1417);
or U271 (N_271,In_205,In_506);
nor U272 (N_272,In_230,In_763);
and U273 (N_273,In_1452,In_1280);
and U274 (N_274,In_228,In_1494);
and U275 (N_275,In_570,In_297);
nand U276 (N_276,In_667,In_814);
or U277 (N_277,In_177,In_221);
and U278 (N_278,In_967,In_346);
xnor U279 (N_279,In_264,In_893);
nor U280 (N_280,In_350,In_547);
and U281 (N_281,In_921,In_660);
or U282 (N_282,In_892,In_620);
nand U283 (N_283,In_1224,In_72);
xnor U284 (N_284,In_400,In_635);
xor U285 (N_285,In_348,In_1450);
nand U286 (N_286,In_1424,In_161);
or U287 (N_287,In_307,In_1066);
nor U288 (N_288,In_424,In_21);
and U289 (N_289,In_875,In_1388);
nand U290 (N_290,In_203,In_303);
nand U291 (N_291,In_1169,In_51);
xor U292 (N_292,In_1035,In_978);
xnor U293 (N_293,In_769,In_1465);
nand U294 (N_294,In_577,In_834);
nor U295 (N_295,In_84,In_1310);
nand U296 (N_296,In_757,In_391);
nor U297 (N_297,In_699,In_1415);
or U298 (N_298,In_1421,In_1279);
and U299 (N_299,In_903,In_1422);
and U300 (N_300,In_1462,In_1072);
nor U301 (N_301,In_1416,In_1079);
xnor U302 (N_302,In_1213,In_182);
xor U303 (N_303,In_1014,In_936);
xor U304 (N_304,In_1112,In_715);
xnor U305 (N_305,In_475,In_928);
and U306 (N_306,In_1077,In_995);
and U307 (N_307,In_62,In_1402);
xor U308 (N_308,In_1060,In_1043);
and U309 (N_309,In_868,In_720);
or U310 (N_310,In_619,In_1485);
or U311 (N_311,In_33,In_1125);
or U312 (N_312,In_1325,In_623);
nand U313 (N_313,In_244,In_1342);
and U314 (N_314,In_414,In_681);
xor U315 (N_315,In_1199,In_572);
nand U316 (N_316,In_320,In_427);
and U317 (N_317,In_692,In_1477);
and U318 (N_318,In_453,In_541);
or U319 (N_319,In_535,In_1429);
nand U320 (N_320,In_48,In_1299);
nor U321 (N_321,In_194,In_154);
and U322 (N_322,In_1292,In_376);
or U323 (N_323,In_1088,In_1460);
or U324 (N_324,In_200,In_287);
xnor U325 (N_325,In_1328,In_1134);
xor U326 (N_326,In_1063,In_91);
or U327 (N_327,In_263,In_1240);
nor U328 (N_328,In_306,In_937);
or U329 (N_329,In_916,In_1384);
and U330 (N_330,In_1448,In_1021);
xnor U331 (N_331,In_9,In_896);
and U332 (N_332,In_618,In_455);
or U333 (N_333,In_298,In_991);
nand U334 (N_334,In_497,In_628);
and U335 (N_335,In_775,In_736);
nand U336 (N_336,In_808,In_37);
xor U337 (N_337,In_352,In_604);
nor U338 (N_338,In_885,In_274);
nand U339 (N_339,In_1042,In_1197);
or U340 (N_340,In_301,In_515);
nor U341 (N_341,In_971,In_603);
and U342 (N_342,In_1095,In_703);
or U343 (N_343,In_386,In_76);
xnor U344 (N_344,In_801,In_641);
xor U345 (N_345,In_413,In_103);
and U346 (N_346,In_1247,In_569);
and U347 (N_347,In_167,In_974);
and U348 (N_348,In_1272,In_1033);
or U349 (N_349,In_60,In_1074);
nor U350 (N_350,In_655,In_404);
nand U351 (N_351,In_305,In_846);
or U352 (N_352,In_1217,In_810);
and U353 (N_353,In_679,In_134);
xor U354 (N_354,In_961,In_366);
or U355 (N_355,In_1277,In_1040);
or U356 (N_356,In_1018,In_554);
xor U357 (N_357,In_38,In_13);
nand U358 (N_358,In_1123,In_847);
or U359 (N_359,In_1106,In_1057);
or U360 (N_360,In_1193,In_1229);
xnor U361 (N_361,In_68,In_484);
nand U362 (N_362,In_790,In_234);
xnor U363 (N_363,In_353,In_1251);
xor U364 (N_364,In_1293,In_457);
nor U365 (N_365,In_727,In_406);
and U366 (N_366,In_524,In_837);
xnor U367 (N_367,In_16,In_951);
or U368 (N_368,In_11,In_1116);
nor U369 (N_369,In_74,In_1411);
nand U370 (N_370,In_1484,In_204);
or U371 (N_371,In_1050,In_266);
and U372 (N_372,In_1355,In_1282);
xor U373 (N_373,In_70,In_202);
xor U374 (N_374,In_573,In_310);
or U375 (N_375,In_1290,In_322);
and U376 (N_376,In_610,In_1288);
nor U377 (N_377,In_1122,In_1385);
and U378 (N_378,In_614,In_1399);
and U379 (N_379,In_235,In_1254);
xnor U380 (N_380,In_663,In_813);
and U381 (N_381,In_1330,In_356);
nor U382 (N_382,In_855,In_1246);
xor U383 (N_383,In_1323,In_633);
xnor U384 (N_384,In_1029,In_325);
nor U385 (N_385,In_71,In_66);
xnor U386 (N_386,In_664,In_286);
and U387 (N_387,In_869,In_788);
nor U388 (N_388,In_127,In_309);
and U389 (N_389,In_377,In_1408);
xnor U390 (N_390,In_687,In_517);
and U391 (N_391,In_636,In_848);
xnor U392 (N_392,In_721,In_1164);
nor U393 (N_393,In_208,In_1237);
nand U394 (N_394,In_1491,In_293);
or U395 (N_395,In_589,In_201);
nor U396 (N_396,In_1359,In_93);
xor U397 (N_397,In_753,In_985);
or U398 (N_398,In_615,In_1141);
nor U399 (N_399,In_1159,In_190);
xnor U400 (N_400,In_644,In_1175);
xor U401 (N_401,In_1350,In_607);
or U402 (N_402,In_1273,In_379);
nand U403 (N_403,In_302,In_1256);
nand U404 (N_404,In_385,In_884);
nor U405 (N_405,In_944,In_511);
or U406 (N_406,In_1027,In_1208);
and U407 (N_407,In_958,In_1281);
and U408 (N_408,In_1356,In_242);
or U409 (N_409,In_472,In_1064);
nor U410 (N_410,In_1149,In_1352);
nand U411 (N_411,In_905,In_1259);
xor U412 (N_412,In_15,In_1092);
or U413 (N_413,In_1470,In_1369);
and U414 (N_414,In_219,In_600);
nor U415 (N_415,In_118,In_983);
nand U416 (N_416,In_477,In_807);
nand U417 (N_417,In_742,In_969);
or U418 (N_418,In_854,In_1326);
nand U419 (N_419,In_924,In_466);
xnor U420 (N_420,In_793,In_1161);
or U421 (N_421,In_1121,In_914);
xor U422 (N_422,In_256,In_1457);
and U423 (N_423,In_493,In_1241);
nand U424 (N_424,In_112,In_1472);
and U425 (N_425,In_285,In_1235);
or U426 (N_426,In_1476,In_191);
and U427 (N_427,In_467,In_504);
xnor U428 (N_428,In_919,In_358);
or U429 (N_429,In_133,In_1349);
xnor U430 (N_430,In_137,In_783);
xnor U431 (N_431,In_1152,In_101);
nor U432 (N_432,In_280,In_1009);
and U433 (N_433,In_382,In_1059);
nand U434 (N_434,In_1258,In_90);
nor U435 (N_435,In_292,In_867);
nand U436 (N_436,In_39,In_1410);
nand U437 (N_437,In_1371,In_1287);
and U438 (N_438,In_599,In_27);
nand U439 (N_439,In_1314,In_393);
nand U440 (N_440,In_369,In_745);
xor U441 (N_441,In_1362,In_1090);
xor U442 (N_442,In_14,In_337);
and U443 (N_443,In_798,In_1188);
xnor U444 (N_444,In_593,In_1347);
nor U445 (N_445,In_858,In_817);
xor U446 (N_446,In_85,In_1461);
or U447 (N_447,In_232,In_22);
and U448 (N_448,In_52,In_1307);
nor U449 (N_449,In_1365,In_520);
xnor U450 (N_450,In_684,In_945);
nand U451 (N_451,In_1115,In_187);
or U452 (N_452,In_601,In_1107);
nand U453 (N_453,In_514,In_1132);
and U454 (N_454,In_1203,In_624);
and U455 (N_455,In_909,In_271);
xor U456 (N_456,In_704,In_501);
and U457 (N_457,In_586,In_1409);
nand U458 (N_458,In_240,In_1196);
xnor U459 (N_459,In_1054,In_268);
or U460 (N_460,In_561,In_949);
xnor U461 (N_461,In_910,In_1353);
and U462 (N_462,In_170,In_349);
xor U463 (N_463,In_227,In_1383);
nand U464 (N_464,In_849,In_1463);
nor U465 (N_465,In_695,In_1295);
or U466 (N_466,In_35,In_1423);
and U467 (N_467,In_1160,In_1474);
nor U468 (N_468,In_1318,In_726);
nor U469 (N_469,In_932,In_313);
or U470 (N_470,In_888,In_1401);
nand U471 (N_471,In_1304,In_546);
nor U472 (N_472,In_1067,In_1173);
or U473 (N_473,In_776,In_1013);
and U474 (N_474,In_722,In_304);
nand U475 (N_475,In_1397,In_1354);
or U476 (N_476,In_717,In_1481);
xor U477 (N_477,In_1061,In_632);
xnor U478 (N_478,In_761,In_345);
and U479 (N_479,In_56,In_741);
nand U480 (N_480,In_216,In_891);
and U481 (N_481,In_1098,In_224);
or U482 (N_482,In_236,In_160);
or U483 (N_483,In_959,In_803);
and U484 (N_484,In_435,In_1382);
nor U485 (N_485,In_934,In_894);
nand U486 (N_486,In_319,In_108);
nand U487 (N_487,In_491,In_1129);
and U488 (N_488,In_186,In_1228);
and U489 (N_489,In_1151,In_1051);
and U490 (N_490,In_871,In_152);
or U491 (N_491,In_831,In_278);
or U492 (N_492,In_544,In_247);
and U493 (N_493,In_412,In_291);
and U494 (N_494,In_1313,In_119);
and U495 (N_495,In_1205,In_676);
xor U496 (N_496,In_1363,In_789);
nand U497 (N_497,In_568,In_1220);
xor U498 (N_498,In_1146,In_707);
nor U499 (N_499,In_700,In_966);
or U500 (N_500,In_1162,In_1344);
xnor U501 (N_501,In_87,In_1184);
xor U502 (N_502,In_861,In_123);
nor U503 (N_503,In_1130,In_1222);
nor U504 (N_504,In_142,In_95);
and U505 (N_505,In_830,In_94);
or U506 (N_506,In_153,In_141);
and U507 (N_507,In_513,In_672);
nor U508 (N_508,In_1221,In_163);
nor U509 (N_509,In_1109,In_136);
or U510 (N_510,In_1267,In_797);
and U511 (N_511,In_1446,In_1268);
xnor U512 (N_512,In_315,In_963);
or U513 (N_513,In_148,In_1338);
xnor U514 (N_514,In_678,In_631);
and U515 (N_515,In_1412,In_1478);
or U516 (N_516,In_30,In_1019);
nand U517 (N_517,In_804,In_1111);
and U518 (N_518,In_422,In_1260);
nand U519 (N_519,In_744,In_392);
and U520 (N_520,In_576,In_470);
xnor U521 (N_521,In_972,In_459);
or U522 (N_522,In_1346,In_365);
nor U523 (N_523,In_870,In_529);
nor U524 (N_524,In_931,In_1315);
and U525 (N_525,In_380,In_873);
nand U526 (N_526,In_1155,In_1144);
nand U527 (N_527,In_1086,In_171);
xnor U528 (N_528,In_805,In_811);
nor U529 (N_529,In_765,In_24);
nand U530 (N_530,In_222,In_1379);
xnor U531 (N_531,In_420,In_1396);
and U532 (N_532,In_759,In_904);
nor U533 (N_533,In_563,In_272);
xor U534 (N_534,In_1147,In_1119);
nor U535 (N_535,In_99,In_629);
xnor U536 (N_536,In_774,In_474);
xor U537 (N_537,In_768,In_1005);
nand U538 (N_538,In_1283,In_705);
nand U539 (N_539,In_1435,In_1181);
xnor U540 (N_540,In_1,In_368);
or U541 (N_541,In_702,In_473);
nand U542 (N_542,In_857,In_738);
xnor U543 (N_543,In_616,In_1200);
xor U544 (N_544,In_145,In_1490);
nand U545 (N_545,In_749,In_1171);
nand U546 (N_546,In_464,In_1148);
nand U547 (N_547,In_502,In_1105);
or U548 (N_548,In_680,In_19);
and U549 (N_549,In_1453,In_1026);
xnor U550 (N_550,In_1376,In_384);
nand U551 (N_551,In_1177,In_233);
xor U552 (N_552,In_40,In_829);
nor U553 (N_553,In_495,In_1413);
nor U554 (N_554,In_553,In_367);
xnor U555 (N_555,In_859,In_964);
xor U556 (N_556,In_296,In_1053);
xnor U557 (N_557,In_714,In_654);
or U558 (N_558,In_1278,In_1071);
and U559 (N_559,In_439,In_102);
xor U560 (N_560,In_321,In_1458);
nand U561 (N_561,In_612,In_317);
xnor U562 (N_562,In_1482,In_925);
nor U563 (N_563,In_1170,In_106);
nand U564 (N_564,In_558,In_183);
nor U565 (N_565,In_747,In_434);
or U566 (N_566,In_906,In_390);
nor U567 (N_567,In_354,In_933);
nor U568 (N_568,In_329,In_989);
nor U569 (N_569,In_709,In_73);
and U570 (N_570,In_973,In_852);
xor U571 (N_571,In_429,In_98);
nand U572 (N_572,In_929,In_336);
nor U573 (N_573,In_410,In_1498);
nor U574 (N_574,In_1209,In_237);
nand U575 (N_575,In_877,In_955);
nor U576 (N_576,In_1191,In_444);
or U577 (N_577,In_860,In_968);
nor U578 (N_578,In_175,In_215);
or U579 (N_579,In_1269,In_253);
xor U580 (N_580,In_169,In_1223);
or U581 (N_581,In_1271,In_748);
xnor U582 (N_582,In_938,In_245);
xnor U583 (N_583,In_1456,In_942);
xor U584 (N_584,In_724,In_578);
nor U585 (N_585,In_1218,In_683);
and U586 (N_586,In_779,In_1285);
and U587 (N_587,In_611,In_490);
nand U588 (N_588,In_1312,In_117);
nand U589 (N_589,In_374,In_172);
nand U590 (N_590,In_1128,In_1455);
or U591 (N_591,In_316,In_1230);
or U592 (N_592,In_1211,In_673);
nor U593 (N_593,In_531,In_176);
nand U594 (N_594,In_838,In_649);
or U595 (N_595,In_423,In_419);
and U596 (N_596,In_882,In_1118);
or U597 (N_597,In_652,In_701);
xnor U598 (N_598,In_1172,In_1270);
xnor U599 (N_599,In_1437,In_1294);
and U600 (N_600,In_344,In_1210);
nand U601 (N_601,In_225,In_1340);
and U602 (N_602,In_166,In_1447);
or U603 (N_603,In_1308,In_403);
xor U604 (N_604,In_1023,In_83);
xor U605 (N_605,In_129,In_357);
nor U606 (N_606,In_1469,In_581);
xor U607 (N_607,In_939,In_826);
and U608 (N_608,In_677,In_952);
or U609 (N_609,In_1000,In_273);
nand U610 (N_610,In_1049,In_1126);
nand U611 (N_611,In_241,In_962);
or U612 (N_612,In_50,In_879);
or U613 (N_613,In_1400,In_1234);
or U614 (N_614,In_552,In_192);
and U615 (N_615,In_334,In_956);
nor U616 (N_616,In_1136,In_698);
nor U617 (N_617,In_1154,In_954);
nand U618 (N_618,In_289,In_733);
and U619 (N_619,In_1047,In_975);
xnor U620 (N_620,In_1076,In_927);
nand U621 (N_621,In_125,In_845);
nand U622 (N_622,In_819,In_333);
nor U623 (N_623,In_674,In_708);
or U624 (N_624,In_911,In_144);
xnor U625 (N_625,In_361,In_347);
xor U626 (N_626,In_556,In_57);
or U627 (N_627,In_314,In_796);
xor U628 (N_628,In_408,In_180);
nand U629 (N_629,In_53,In_26);
nand U630 (N_630,In_850,In_135);
or U631 (N_631,In_411,In_878);
nand U632 (N_632,In_1492,In_1372);
and U633 (N_633,In_211,In_536);
nand U634 (N_634,In_20,In_516);
and U635 (N_635,In_1393,In_465);
and U636 (N_636,In_251,In_540);
and U637 (N_637,In_284,In_1459);
nor U638 (N_638,In_405,In_86);
nor U639 (N_639,In_430,In_670);
and U640 (N_640,In_58,In_697);
and U641 (N_641,In_438,In_613);
and U642 (N_642,In_771,In_1212);
or U643 (N_643,In_690,In_458);
xnor U644 (N_644,In_1486,In_311);
and U645 (N_645,In_1381,In_389);
nor U646 (N_646,In_1024,In_912);
or U647 (N_647,In_548,In_1358);
and U648 (N_648,In_165,In_1012);
nand U649 (N_649,In_496,In_626);
nand U650 (N_650,In_1380,In_980);
or U651 (N_651,In_809,In_479);
and U652 (N_652,In_835,In_146);
nand U653 (N_653,In_512,In_815);
nand U654 (N_654,In_918,In_772);
or U655 (N_655,In_777,In_446);
xor U656 (N_656,In_2,In_920);
xor U657 (N_657,In_555,In_6);
nand U658 (N_658,In_650,In_1479);
or U659 (N_659,In_1052,In_999);
or U660 (N_660,In_1178,In_10);
nand U661 (N_661,In_659,In_1245);
xnor U662 (N_662,In_468,In_1337);
xnor U663 (N_663,In_943,In_778);
nand U664 (N_664,In_1163,In_1145);
nand U665 (N_665,In_575,In_587);
nor U666 (N_666,In_1361,In_642);
xnor U667 (N_667,In_770,In_794);
xnor U668 (N_668,In_1166,In_198);
and U669 (N_669,In_1127,In_832);
nor U670 (N_670,In_1085,In_1073);
xnor U671 (N_671,In_823,In_121);
nand U672 (N_672,In_300,In_54);
nand U673 (N_673,In_341,In_1440);
xnor U674 (N_674,In_128,In_1302);
and U675 (N_675,In_488,In_1093);
nand U676 (N_676,In_282,In_437);
nand U677 (N_677,In_1156,In_639);
nor U678 (N_678,In_1389,In_532);
or U679 (N_679,In_902,In_1015);
nand U680 (N_680,In_159,In_865);
nor U681 (N_681,In_214,In_89);
nand U682 (N_682,In_1201,In_34);
or U683 (N_683,In_36,In_781);
and U684 (N_684,In_1451,In_113);
and U685 (N_685,In_579,In_737);
and U686 (N_686,In_773,In_1238);
nor U687 (N_687,In_1274,In_1305);
or U688 (N_688,In_1309,In_923);
nand U689 (N_689,In_510,In_1094);
or U690 (N_690,In_1449,In_1065);
xnor U691 (N_691,In_518,In_1316);
and U692 (N_692,In_1135,In_407);
xnor U693 (N_693,In_1150,In_596);
or U694 (N_694,In_0,In_1133);
xor U695 (N_695,In_762,In_371);
and U696 (N_696,In_818,In_1487);
nand U697 (N_697,In_950,In_1420);
xor U698 (N_698,In_4,In_1089);
or U699 (N_699,In_1370,In_856);
nor U700 (N_700,In_156,In_1341);
and U701 (N_701,In_822,In_440);
and U702 (N_702,In_521,In_1097);
and U703 (N_703,In_482,In_259);
nor U704 (N_704,In_669,In_1253);
xor U705 (N_705,In_1483,In_195);
nor U706 (N_706,In_471,In_866);
or U707 (N_707,In_992,In_1303);
or U708 (N_708,In_318,In_970);
and U709 (N_709,In_750,In_1488);
xnor U710 (N_710,In_109,In_1473);
nor U711 (N_711,In_998,In_539);
nor U712 (N_712,In_1339,In_388);
and U713 (N_713,In_1394,In_1082);
nor U714 (N_714,In_299,In_162);
nor U715 (N_715,In_212,In_621);
and U716 (N_716,In_265,In_719);
nand U717 (N_717,In_1017,In_220);
xnor U718 (N_718,In_1058,In_343);
xnor U719 (N_719,In_922,In_986);
nor U720 (N_720,In_767,In_469);
nand U721 (N_721,In_207,In_481);
nor U722 (N_722,In_564,In_1186);
xnor U723 (N_723,In_360,In_1206);
xor U724 (N_724,In_732,In_1496);
nor U725 (N_725,In_953,In_1466);
nand U726 (N_726,In_1495,In_270);
or U727 (N_727,In_189,In_606);
nor U728 (N_728,In_238,In_485);
and U729 (N_729,In_1232,In_746);
nor U730 (N_730,In_1442,In_1327);
nand U731 (N_731,In_1414,In_930);
xnor U732 (N_732,In_1103,In_1070);
or U733 (N_733,In_460,In_231);
and U734 (N_734,In_421,In_874);
nand U735 (N_735,In_363,In_549);
nand U736 (N_736,In_786,In_1239);
xor U737 (N_737,In_1348,In_647);
xor U738 (N_738,In_1153,In_1131);
and U739 (N_739,In_1216,In_1403);
xnor U740 (N_740,In_151,In_1345);
xor U741 (N_741,In_1226,In_760);
xor U742 (N_742,In_1038,In_1236);
or U743 (N_743,In_806,In_812);
nor U744 (N_744,In_617,In_1427);
nand U745 (N_745,In_836,In_557);
nor U746 (N_746,In_565,In_1499);
or U747 (N_747,In_728,In_656);
xor U748 (N_748,In_226,In_1284);
nand U749 (N_749,In_276,In_661);
and U750 (N_750,In_734,In_789);
or U751 (N_751,In_823,In_1144);
and U752 (N_752,In_5,In_965);
nand U753 (N_753,In_547,In_573);
nor U754 (N_754,In_1222,In_1191);
or U755 (N_755,In_1480,In_171);
xnor U756 (N_756,In_1205,In_384);
or U757 (N_757,In_855,In_345);
nand U758 (N_758,In_613,In_1180);
xnor U759 (N_759,In_1459,In_117);
nand U760 (N_760,In_128,In_334);
xnor U761 (N_761,In_1101,In_376);
or U762 (N_762,In_50,In_251);
xor U763 (N_763,In_1248,In_713);
and U764 (N_764,In_849,In_143);
or U765 (N_765,In_128,In_196);
or U766 (N_766,In_55,In_565);
nor U767 (N_767,In_564,In_702);
xor U768 (N_768,In_453,In_821);
or U769 (N_769,In_1384,In_165);
xor U770 (N_770,In_806,In_2);
xnor U771 (N_771,In_760,In_1168);
nor U772 (N_772,In_1240,In_151);
nor U773 (N_773,In_30,In_36);
or U774 (N_774,In_1054,In_1217);
and U775 (N_775,In_1412,In_140);
xor U776 (N_776,In_449,In_1351);
nor U777 (N_777,In_966,In_320);
and U778 (N_778,In_920,In_163);
and U779 (N_779,In_297,In_565);
xnor U780 (N_780,In_1077,In_1126);
xor U781 (N_781,In_1267,In_1402);
nand U782 (N_782,In_346,In_277);
nand U783 (N_783,In_402,In_276);
and U784 (N_784,In_336,In_324);
and U785 (N_785,In_1131,In_500);
nor U786 (N_786,In_474,In_911);
or U787 (N_787,In_1029,In_827);
nand U788 (N_788,In_1055,In_1148);
nand U789 (N_789,In_1146,In_466);
and U790 (N_790,In_737,In_1178);
and U791 (N_791,In_972,In_407);
xnor U792 (N_792,In_1205,In_1100);
xnor U793 (N_793,In_1,In_128);
xnor U794 (N_794,In_1472,In_57);
xor U795 (N_795,In_51,In_129);
nor U796 (N_796,In_1005,In_1268);
and U797 (N_797,In_184,In_1149);
and U798 (N_798,In_544,In_482);
nor U799 (N_799,In_656,In_1171);
nand U800 (N_800,In_412,In_680);
nand U801 (N_801,In_139,In_1046);
xor U802 (N_802,In_6,In_411);
xor U803 (N_803,In_836,In_304);
and U804 (N_804,In_269,In_1078);
nor U805 (N_805,In_343,In_1303);
or U806 (N_806,In_271,In_129);
and U807 (N_807,In_1006,In_1302);
and U808 (N_808,In_635,In_1156);
and U809 (N_809,In_889,In_888);
and U810 (N_810,In_374,In_719);
xor U811 (N_811,In_58,In_1433);
and U812 (N_812,In_909,In_862);
and U813 (N_813,In_48,In_851);
nand U814 (N_814,In_858,In_1112);
nand U815 (N_815,In_1248,In_407);
nor U816 (N_816,In_453,In_756);
nor U817 (N_817,In_1483,In_876);
nor U818 (N_818,In_731,In_237);
xor U819 (N_819,In_15,In_1227);
nor U820 (N_820,In_205,In_102);
nand U821 (N_821,In_1138,In_785);
nand U822 (N_822,In_753,In_18);
xor U823 (N_823,In_797,In_255);
xnor U824 (N_824,In_1270,In_699);
nand U825 (N_825,In_1083,In_705);
nor U826 (N_826,In_674,In_225);
xnor U827 (N_827,In_805,In_1190);
and U828 (N_828,In_54,In_838);
nor U829 (N_829,In_449,In_937);
and U830 (N_830,In_1166,In_1364);
or U831 (N_831,In_1278,In_952);
or U832 (N_832,In_326,In_1316);
nand U833 (N_833,In_1164,In_556);
nor U834 (N_834,In_1293,In_1415);
and U835 (N_835,In_957,In_464);
and U836 (N_836,In_1179,In_671);
or U837 (N_837,In_904,In_37);
and U838 (N_838,In_654,In_961);
nor U839 (N_839,In_57,In_421);
nor U840 (N_840,In_1205,In_661);
nand U841 (N_841,In_208,In_86);
and U842 (N_842,In_1132,In_170);
xor U843 (N_843,In_271,In_936);
and U844 (N_844,In_32,In_181);
nand U845 (N_845,In_194,In_501);
and U846 (N_846,In_807,In_887);
and U847 (N_847,In_233,In_322);
and U848 (N_848,In_305,In_1050);
xor U849 (N_849,In_665,In_325);
nand U850 (N_850,In_28,In_47);
xor U851 (N_851,In_1200,In_123);
nor U852 (N_852,In_52,In_1350);
nand U853 (N_853,In_296,In_1074);
or U854 (N_854,In_1458,In_347);
xnor U855 (N_855,In_405,In_133);
nand U856 (N_856,In_577,In_1499);
xor U857 (N_857,In_1370,In_289);
xnor U858 (N_858,In_471,In_475);
or U859 (N_859,In_1183,In_1111);
xor U860 (N_860,In_231,In_29);
and U861 (N_861,In_1313,In_250);
xnor U862 (N_862,In_905,In_695);
and U863 (N_863,In_1279,In_1008);
xnor U864 (N_864,In_1121,In_889);
and U865 (N_865,In_431,In_667);
and U866 (N_866,In_655,In_1310);
nand U867 (N_867,In_1276,In_1454);
nor U868 (N_868,In_1270,In_635);
and U869 (N_869,In_1039,In_343);
or U870 (N_870,In_265,In_587);
and U871 (N_871,In_92,In_1377);
and U872 (N_872,In_590,In_32);
nand U873 (N_873,In_304,In_133);
xor U874 (N_874,In_546,In_100);
or U875 (N_875,In_1308,In_766);
nand U876 (N_876,In_1211,In_459);
xnor U877 (N_877,In_1053,In_1135);
and U878 (N_878,In_920,In_877);
nor U879 (N_879,In_1455,In_770);
nor U880 (N_880,In_299,In_693);
or U881 (N_881,In_1444,In_940);
or U882 (N_882,In_1259,In_312);
xnor U883 (N_883,In_1102,In_1220);
or U884 (N_884,In_881,In_217);
or U885 (N_885,In_146,In_464);
nand U886 (N_886,In_215,In_1060);
nand U887 (N_887,In_87,In_974);
or U888 (N_888,In_333,In_1261);
or U889 (N_889,In_1202,In_705);
and U890 (N_890,In_1218,In_196);
and U891 (N_891,In_1019,In_889);
xnor U892 (N_892,In_111,In_417);
or U893 (N_893,In_1223,In_1131);
nand U894 (N_894,In_445,In_851);
nand U895 (N_895,In_722,In_809);
xor U896 (N_896,In_274,In_1426);
xor U897 (N_897,In_914,In_353);
or U898 (N_898,In_488,In_404);
and U899 (N_899,In_1085,In_652);
nor U900 (N_900,In_99,In_1444);
xnor U901 (N_901,In_481,In_414);
and U902 (N_902,In_919,In_1160);
xnor U903 (N_903,In_747,In_350);
and U904 (N_904,In_940,In_1158);
xnor U905 (N_905,In_1225,In_608);
xnor U906 (N_906,In_647,In_225);
nor U907 (N_907,In_584,In_459);
or U908 (N_908,In_1257,In_1229);
nor U909 (N_909,In_330,In_163);
or U910 (N_910,In_831,In_775);
xor U911 (N_911,In_1151,In_985);
and U912 (N_912,In_1259,In_1334);
nor U913 (N_913,In_277,In_1069);
xnor U914 (N_914,In_43,In_753);
and U915 (N_915,In_1091,In_1180);
nand U916 (N_916,In_1003,In_1494);
nor U917 (N_917,In_849,In_9);
nand U918 (N_918,In_766,In_620);
nand U919 (N_919,In_328,In_209);
nand U920 (N_920,In_1345,In_242);
xor U921 (N_921,In_1362,In_1055);
or U922 (N_922,In_211,In_341);
and U923 (N_923,In_790,In_1116);
xnor U924 (N_924,In_1086,In_583);
xnor U925 (N_925,In_403,In_1477);
and U926 (N_926,In_113,In_1101);
nand U927 (N_927,In_1045,In_1429);
or U928 (N_928,In_79,In_52);
nor U929 (N_929,In_788,In_286);
nor U930 (N_930,In_1000,In_369);
or U931 (N_931,In_1020,In_714);
and U932 (N_932,In_1357,In_732);
nand U933 (N_933,In_1353,In_895);
or U934 (N_934,In_834,In_140);
or U935 (N_935,In_568,In_1491);
nor U936 (N_936,In_1378,In_693);
or U937 (N_937,In_665,In_178);
xor U938 (N_938,In_759,In_497);
nor U939 (N_939,In_691,In_1099);
and U940 (N_940,In_704,In_1426);
xor U941 (N_941,In_720,In_1468);
nor U942 (N_942,In_371,In_51);
xnor U943 (N_943,In_916,In_573);
xor U944 (N_944,In_633,In_211);
and U945 (N_945,In_41,In_1370);
nor U946 (N_946,In_994,In_244);
nand U947 (N_947,In_515,In_1022);
nor U948 (N_948,In_310,In_230);
and U949 (N_949,In_729,In_1481);
nor U950 (N_950,In_840,In_468);
or U951 (N_951,In_305,In_868);
nand U952 (N_952,In_260,In_936);
nand U953 (N_953,In_990,In_1119);
nand U954 (N_954,In_767,In_157);
or U955 (N_955,In_984,In_1122);
xnor U956 (N_956,In_1350,In_381);
xor U957 (N_957,In_743,In_72);
or U958 (N_958,In_439,In_172);
xor U959 (N_959,In_1383,In_1193);
or U960 (N_960,In_561,In_1161);
nor U961 (N_961,In_1220,In_1003);
nor U962 (N_962,In_536,In_915);
or U963 (N_963,In_1052,In_507);
or U964 (N_964,In_57,In_1428);
nor U965 (N_965,In_1419,In_381);
xnor U966 (N_966,In_732,In_621);
xor U967 (N_967,In_1378,In_1139);
and U968 (N_968,In_429,In_1458);
nand U969 (N_969,In_1491,In_965);
or U970 (N_970,In_1424,In_838);
xnor U971 (N_971,In_648,In_828);
nor U972 (N_972,In_980,In_611);
or U973 (N_973,In_996,In_186);
xor U974 (N_974,In_908,In_589);
nand U975 (N_975,In_571,In_840);
xor U976 (N_976,In_548,In_1233);
or U977 (N_977,In_723,In_91);
xor U978 (N_978,In_915,In_1405);
nor U979 (N_979,In_105,In_635);
xor U980 (N_980,In_421,In_500);
nand U981 (N_981,In_1218,In_68);
or U982 (N_982,In_576,In_996);
nand U983 (N_983,In_166,In_731);
or U984 (N_984,In_72,In_952);
xor U985 (N_985,In_94,In_555);
nor U986 (N_986,In_81,In_670);
xnor U987 (N_987,In_330,In_1399);
nand U988 (N_988,In_236,In_975);
and U989 (N_989,In_1109,In_1115);
and U990 (N_990,In_1065,In_781);
xnor U991 (N_991,In_606,In_20);
xor U992 (N_992,In_758,In_587);
nand U993 (N_993,In_645,In_974);
xor U994 (N_994,In_236,In_389);
nand U995 (N_995,In_1302,In_743);
nand U996 (N_996,In_1010,In_395);
nand U997 (N_997,In_217,In_563);
or U998 (N_998,In_164,In_1331);
nand U999 (N_999,In_1250,In_774);
and U1000 (N_1000,N_641,N_276);
nor U1001 (N_1001,N_927,N_374);
or U1002 (N_1002,N_784,N_421);
and U1003 (N_1003,N_502,N_716);
nor U1004 (N_1004,N_922,N_493);
nor U1005 (N_1005,N_562,N_28);
and U1006 (N_1006,N_742,N_867);
nand U1007 (N_1007,N_692,N_947);
or U1008 (N_1008,N_693,N_843);
and U1009 (N_1009,N_16,N_943);
nand U1010 (N_1010,N_77,N_87);
nand U1011 (N_1011,N_949,N_623);
nand U1012 (N_1012,N_176,N_183);
xnor U1013 (N_1013,N_406,N_361);
or U1014 (N_1014,N_537,N_257);
xor U1015 (N_1015,N_155,N_78);
nor U1016 (N_1016,N_112,N_894);
nand U1017 (N_1017,N_325,N_862);
or U1018 (N_1018,N_69,N_152);
and U1019 (N_1019,N_130,N_431);
xnor U1020 (N_1020,N_428,N_911);
nor U1021 (N_1021,N_929,N_826);
nor U1022 (N_1022,N_430,N_719);
nand U1023 (N_1023,N_665,N_440);
xnor U1024 (N_1024,N_533,N_688);
nand U1025 (N_1025,N_738,N_301);
xor U1026 (N_1026,N_909,N_856);
or U1027 (N_1027,N_48,N_254);
or U1028 (N_1028,N_272,N_504);
and U1029 (N_1029,N_554,N_674);
nor U1030 (N_1030,N_467,N_119);
xor U1031 (N_1031,N_451,N_669);
xnor U1032 (N_1032,N_382,N_633);
nand U1033 (N_1033,N_759,N_445);
and U1034 (N_1034,N_309,N_79);
xor U1035 (N_1035,N_921,N_355);
nor U1036 (N_1036,N_118,N_380);
nand U1037 (N_1037,N_95,N_195);
nor U1038 (N_1038,N_785,N_34);
nand U1039 (N_1039,N_882,N_706);
xor U1040 (N_1040,N_810,N_778);
nand U1041 (N_1041,N_46,N_941);
nand U1042 (N_1042,N_748,N_52);
xnor U1043 (N_1043,N_679,N_164);
nor U1044 (N_1044,N_343,N_967);
or U1045 (N_1045,N_621,N_106);
xor U1046 (N_1046,N_847,N_991);
xor U1047 (N_1047,N_851,N_645);
and U1048 (N_1048,N_455,N_369);
or U1049 (N_1049,N_116,N_629);
xor U1050 (N_1050,N_1,N_626);
and U1051 (N_1051,N_469,N_173);
and U1052 (N_1052,N_560,N_464);
or U1053 (N_1053,N_30,N_558);
xor U1054 (N_1054,N_547,N_391);
or U1055 (N_1055,N_475,N_340);
xor U1056 (N_1056,N_178,N_244);
and U1057 (N_1057,N_267,N_160);
nand U1058 (N_1058,N_830,N_898);
and U1059 (N_1059,N_908,N_162);
xnor U1060 (N_1060,N_494,N_823);
nor U1061 (N_1061,N_584,N_465);
nor U1062 (N_1062,N_189,N_170);
or U1063 (N_1063,N_787,N_161);
and U1064 (N_1064,N_407,N_668);
and U1065 (N_1065,N_275,N_612);
nand U1066 (N_1066,N_920,N_347);
xor U1067 (N_1067,N_43,N_866);
xor U1068 (N_1068,N_655,N_619);
and U1069 (N_1069,N_695,N_863);
nand U1070 (N_1070,N_765,N_757);
and U1071 (N_1071,N_539,N_39);
or U1072 (N_1072,N_875,N_578);
and U1073 (N_1073,N_721,N_594);
or U1074 (N_1074,N_501,N_811);
nor U1075 (N_1075,N_804,N_385);
nor U1076 (N_1076,N_561,N_609);
nand U1077 (N_1077,N_684,N_268);
nor U1078 (N_1078,N_874,N_981);
and U1079 (N_1079,N_315,N_892);
or U1080 (N_1080,N_60,N_559);
or U1081 (N_1081,N_532,N_797);
xnor U1082 (N_1082,N_767,N_148);
nand U1083 (N_1083,N_821,N_958);
nor U1084 (N_1084,N_214,N_435);
nor U1085 (N_1085,N_191,N_53);
nand U1086 (N_1086,N_153,N_128);
nand U1087 (N_1087,N_289,N_915);
and U1088 (N_1088,N_163,N_98);
nand U1089 (N_1089,N_513,N_470);
nor U1090 (N_1090,N_76,N_311);
nand U1091 (N_1091,N_661,N_886);
and U1092 (N_1092,N_528,N_792);
or U1093 (N_1093,N_485,N_381);
nor U1094 (N_1094,N_2,N_703);
xnor U1095 (N_1095,N_263,N_774);
nand U1096 (N_1096,N_47,N_756);
xnor U1097 (N_1097,N_614,N_989);
or U1098 (N_1098,N_322,N_857);
nor U1099 (N_1099,N_646,N_239);
nand U1100 (N_1100,N_243,N_223);
and U1101 (N_1101,N_868,N_218);
and U1102 (N_1102,N_593,N_964);
nor U1103 (N_1103,N_535,N_459);
nor U1104 (N_1104,N_110,N_364);
or U1105 (N_1105,N_67,N_709);
and U1106 (N_1106,N_476,N_8);
xor U1107 (N_1107,N_859,N_417);
and U1108 (N_1108,N_174,N_360);
or U1109 (N_1109,N_832,N_788);
or U1110 (N_1110,N_286,N_251);
nand U1111 (N_1111,N_818,N_509);
xnor U1112 (N_1112,N_26,N_957);
xnor U1113 (N_1113,N_480,N_809);
nor U1114 (N_1114,N_897,N_357);
nor U1115 (N_1115,N_22,N_326);
and U1116 (N_1116,N_534,N_918);
and U1117 (N_1117,N_586,N_350);
nor U1118 (N_1118,N_241,N_20);
or U1119 (N_1119,N_403,N_605);
xor U1120 (N_1120,N_802,N_64);
or U1121 (N_1121,N_68,N_149);
and U1122 (N_1122,N_179,N_583);
nor U1123 (N_1123,N_515,N_763);
nand U1124 (N_1124,N_216,N_849);
nor U1125 (N_1125,N_117,N_966);
or U1126 (N_1126,N_198,N_114);
nand U1127 (N_1127,N_545,N_525);
and U1128 (N_1128,N_105,N_516);
or U1129 (N_1129,N_422,N_491);
or U1130 (N_1130,N_346,N_331);
nor U1131 (N_1131,N_760,N_492);
and U1132 (N_1132,N_600,N_879);
or U1133 (N_1133,N_727,N_202);
or U1134 (N_1134,N_365,N_858);
nand U1135 (N_1135,N_872,N_447);
nand U1136 (N_1136,N_318,N_122);
and U1137 (N_1137,N_711,N_540);
nor U1138 (N_1138,N_154,N_400);
or U1139 (N_1139,N_990,N_676);
xnor U1140 (N_1140,N_429,N_895);
nor U1141 (N_1141,N_893,N_781);
nor U1142 (N_1142,N_671,N_881);
nor U1143 (N_1143,N_25,N_466);
nor U1144 (N_1144,N_187,N_878);
xor U1145 (N_1145,N_889,N_726);
and U1146 (N_1146,N_959,N_635);
and U1147 (N_1147,N_955,N_660);
nand U1148 (N_1148,N_582,N_401);
xnor U1149 (N_1149,N_253,N_463);
and U1150 (N_1150,N_885,N_200);
nor U1151 (N_1151,N_379,N_328);
nor U1152 (N_1152,N_304,N_890);
xnor U1153 (N_1153,N_603,N_490);
nand U1154 (N_1154,N_997,N_975);
nor U1155 (N_1155,N_281,N_770);
nor U1156 (N_1156,N_396,N_731);
nor U1157 (N_1157,N_529,N_324);
xor U1158 (N_1158,N_94,N_415);
and U1159 (N_1159,N_446,N_249);
xnor U1160 (N_1160,N_486,N_739);
nand U1161 (N_1161,N_933,N_245);
nor U1162 (N_1162,N_983,N_852);
or U1163 (N_1163,N_312,N_568);
and U1164 (N_1164,N_702,N_33);
and U1165 (N_1165,N_754,N_632);
nand U1166 (N_1166,N_15,N_722);
nor U1167 (N_1167,N_685,N_83);
or U1168 (N_1168,N_675,N_423);
xnor U1169 (N_1169,N_387,N_375);
or U1170 (N_1170,N_750,N_181);
xnor U1171 (N_1171,N_905,N_377);
or U1172 (N_1172,N_682,N_256);
nor U1173 (N_1173,N_994,N_556);
xnor U1174 (N_1174,N_814,N_631);
or U1175 (N_1175,N_441,N_332);
nor U1176 (N_1176,N_277,N_707);
nand U1177 (N_1177,N_426,N_327);
or U1178 (N_1178,N_691,N_271);
or U1179 (N_1179,N_686,N_371);
xor U1180 (N_1180,N_743,N_55);
or U1181 (N_1181,N_462,N_227);
nor U1182 (N_1182,N_769,N_837);
xnor U1183 (N_1183,N_232,N_523);
nor U1184 (N_1184,N_884,N_12);
and U1185 (N_1185,N_642,N_776);
nand U1186 (N_1186,N_215,N_261);
xor U1187 (N_1187,N_574,N_969);
or U1188 (N_1188,N_71,N_335);
or U1189 (N_1189,N_589,N_799);
or U1190 (N_1190,N_193,N_916);
nor U1191 (N_1191,N_235,N_260);
and U1192 (N_1192,N_590,N_505);
nand U1193 (N_1193,N_530,N_656);
nand U1194 (N_1194,N_511,N_296);
nor U1195 (N_1195,N_390,N_436);
xor U1196 (N_1196,N_13,N_902);
nor U1197 (N_1197,N_820,N_704);
nand U1198 (N_1198,N_433,N_977);
or U1199 (N_1199,N_62,N_771);
nor U1200 (N_1200,N_103,N_993);
and U1201 (N_1201,N_196,N_368);
and U1202 (N_1202,N_229,N_291);
nor U1203 (N_1203,N_316,N_274);
or U1204 (N_1204,N_950,N_376);
or U1205 (N_1205,N_82,N_168);
xor U1206 (N_1206,N_698,N_5);
xnor U1207 (N_1207,N_458,N_735);
or U1208 (N_1208,N_566,N_714);
nand U1209 (N_1209,N_551,N_307);
nand U1210 (N_1210,N_917,N_24);
and U1211 (N_1211,N_487,N_230);
or U1212 (N_1212,N_57,N_14);
or U1213 (N_1213,N_199,N_258);
nand U1214 (N_1214,N_512,N_313);
or U1215 (N_1215,N_388,N_180);
xnor U1216 (N_1216,N_410,N_951);
and U1217 (N_1217,N_109,N_712);
xor U1218 (N_1218,N_579,N_640);
nand U1219 (N_1219,N_65,N_613);
nand U1220 (N_1220,N_54,N_616);
nor U1221 (N_1221,N_352,N_974);
and U1222 (N_1222,N_617,N_45);
or U1223 (N_1223,N_667,N_996);
or U1224 (N_1224,N_982,N_705);
xnor U1225 (N_1225,N_518,N_341);
and U1226 (N_1226,N_987,N_963);
nor U1227 (N_1227,N_782,N_495);
xor U1228 (N_1228,N_454,N_483);
nand U1229 (N_1229,N_777,N_73);
xor U1230 (N_1230,N_194,N_846);
nor U1231 (N_1231,N_489,N_344);
and U1232 (N_1232,N_29,N_132);
nand U1233 (N_1233,N_242,N_126);
xor U1234 (N_1234,N_571,N_337);
nand U1235 (N_1235,N_934,N_452);
xnor U1236 (N_1236,N_803,N_18);
and U1237 (N_1237,N_970,N_753);
nor U1238 (N_1238,N_449,N_165);
and U1239 (N_1239,N_366,N_353);
or U1240 (N_1240,N_510,N_333);
nand U1241 (N_1241,N_177,N_228);
and U1242 (N_1242,N_945,N_143);
xor U1243 (N_1243,N_405,N_740);
nor U1244 (N_1244,N_231,N_737);
nor U1245 (N_1245,N_348,N_443);
xnor U1246 (N_1246,N_808,N_666);
xnor U1247 (N_1247,N_570,N_701);
nor U1248 (N_1248,N_386,N_226);
and U1249 (N_1249,N_358,N_877);
or U1250 (N_1250,N_238,N_651);
xnor U1251 (N_1251,N_795,N_644);
xnor U1252 (N_1252,N_828,N_437);
nand U1253 (N_1253,N_988,N_330);
and U1254 (N_1254,N_891,N_292);
or U1255 (N_1255,N_548,N_936);
or U1256 (N_1256,N_524,N_97);
and U1257 (N_1257,N_608,N_188);
and U1258 (N_1258,N_115,N_624);
nand U1259 (N_1259,N_829,N_157);
xnor U1260 (N_1260,N_473,N_448);
nor U1261 (N_1261,N_92,N_285);
nor U1262 (N_1262,N_323,N_484);
or U1263 (N_1263,N_156,N_456);
or U1264 (N_1264,N_815,N_648);
xor U1265 (N_1265,N_637,N_394);
nand U1266 (N_1266,N_602,N_887);
and U1267 (N_1267,N_10,N_192);
and U1268 (N_1268,N_546,N_497);
xnor U1269 (N_1269,N_869,N_351);
and U1270 (N_1270,N_273,N_555);
nor U1271 (N_1271,N_657,N_710);
and U1272 (N_1272,N_131,N_146);
or U1273 (N_1273,N_827,N_166);
nor U1274 (N_1274,N_72,N_63);
xnor U1275 (N_1275,N_142,N_389);
nand U1276 (N_1276,N_61,N_786);
or U1277 (N_1277,N_506,N_942);
nand U1278 (N_1278,N_32,N_246);
nand U1279 (N_1279,N_734,N_0);
xor U1280 (N_1280,N_222,N_972);
xnor U1281 (N_1281,N_96,N_718);
xnor U1282 (N_1282,N_751,N_564);
xnor U1283 (N_1283,N_549,N_725);
nand U1284 (N_1284,N_101,N_234);
and U1285 (N_1285,N_362,N_658);
xor U1286 (N_1286,N_413,N_461);
and U1287 (N_1287,N_50,N_209);
xor U1288 (N_1288,N_762,N_604);
nand U1289 (N_1289,N_906,N_418);
nor U1290 (N_1290,N_663,N_85);
or U1291 (N_1291,N_597,N_962);
xnor U1292 (N_1292,N_848,N_74);
or U1293 (N_1293,N_80,N_186);
nor U1294 (N_1294,N_393,N_819);
and U1295 (N_1295,N_749,N_690);
and U1296 (N_1296,N_773,N_514);
nand U1297 (N_1297,N_460,N_914);
xor U1298 (N_1298,N_402,N_356);
or U1299 (N_1299,N_172,N_541);
nand U1300 (N_1300,N_806,N_986);
or U1301 (N_1301,N_468,N_184);
and U1302 (N_1302,N_896,N_519);
nor U1303 (N_1303,N_816,N_789);
nand U1304 (N_1304,N_425,N_424);
nor U1305 (N_1305,N_783,N_91);
nor U1306 (N_1306,N_543,N_946);
xnor U1307 (N_1307,N_971,N_766);
or U1308 (N_1308,N_137,N_833);
nor U1309 (N_1309,N_320,N_831);
and U1310 (N_1310,N_221,N_567);
or U1311 (N_1311,N_978,N_290);
or U1312 (N_1312,N_295,N_817);
xnor U1313 (N_1313,N_954,N_610);
xnor U1314 (N_1314,N_84,N_17);
nand U1315 (N_1315,N_19,N_383);
or U1316 (N_1316,N_158,N_683);
nand U1317 (N_1317,N_139,N_659);
and U1318 (N_1318,N_219,N_450);
nand U1319 (N_1319,N_217,N_354);
nand U1320 (N_1320,N_836,N_372);
nor U1321 (N_1321,N_412,N_834);
xor U1322 (N_1322,N_150,N_937);
and U1323 (N_1323,N_520,N_213);
nand U1324 (N_1324,N_81,N_932);
and U1325 (N_1325,N_746,N_888);
nand U1326 (N_1326,N_960,N_27);
and U1327 (N_1327,N_120,N_58);
xor U1328 (N_1328,N_576,N_517);
nor U1329 (N_1329,N_968,N_628);
and U1330 (N_1330,N_167,N_764);
or U1331 (N_1331,N_138,N_907);
or U1332 (N_1332,N_973,N_44);
nor U1333 (N_1333,N_813,N_952);
nor U1334 (N_1334,N_363,N_248);
nand U1335 (N_1335,N_662,N_673);
or U1336 (N_1336,N_419,N_398);
nand U1337 (N_1337,N_596,N_761);
or U1338 (N_1338,N_536,N_100);
and U1339 (N_1339,N_796,N_338);
and U1340 (N_1340,N_930,N_190);
xnor U1341 (N_1341,N_841,N_573);
nand U1342 (N_1342,N_741,N_775);
and U1343 (N_1343,N_845,N_649);
or U1344 (N_1344,N_416,N_636);
and U1345 (N_1345,N_479,N_652);
xnor U1346 (N_1346,N_980,N_538);
and U1347 (N_1347,N_41,N_585);
nand U1348 (N_1348,N_408,N_144);
xnor U1349 (N_1349,N_599,N_399);
nor U1350 (N_1350,N_279,N_317);
and U1351 (N_1351,N_910,N_123);
and U1352 (N_1352,N_850,N_283);
xnor U1353 (N_1353,N_794,N_595);
or U1354 (N_1354,N_38,N_572);
or U1355 (N_1355,N_303,N_42);
and U1356 (N_1356,N_591,N_854);
xnor U1357 (N_1357,N_925,N_370);
and U1358 (N_1358,N_236,N_618);
or U1359 (N_1359,N_615,N_720);
and U1360 (N_1360,N_876,N_6);
and U1361 (N_1361,N_569,N_625);
or U1362 (N_1362,N_284,N_689);
nand U1363 (N_1363,N_713,N_953);
nand U1364 (N_1364,N_21,N_992);
xnor U1365 (N_1365,N_565,N_99);
nor U1366 (N_1366,N_247,N_824);
xor U1367 (N_1367,N_134,N_439);
xnor U1368 (N_1368,N_207,N_210);
nor U1369 (N_1369,N_899,N_171);
nand U1370 (N_1370,N_339,N_308);
and U1371 (N_1371,N_264,N_240);
or U1372 (N_1372,N_125,N_580);
xor U1373 (N_1373,N_627,N_728);
and U1374 (N_1374,N_883,N_36);
or U1375 (N_1375,N_855,N_639);
nand U1376 (N_1376,N_681,N_940);
or U1377 (N_1377,N_880,N_88);
xor U1378 (N_1378,N_453,N_550);
nor U1379 (N_1379,N_444,N_715);
xnor U1380 (N_1380,N_409,N_620);
nor U1381 (N_1381,N_336,N_508);
or U1382 (N_1382,N_938,N_839);
xnor U1383 (N_1383,N_182,N_107);
and U1384 (N_1384,N_758,N_302);
nand U1385 (N_1385,N_287,N_305);
and U1386 (N_1386,N_4,N_237);
or U1387 (N_1387,N_939,N_723);
and U1388 (N_1388,N_844,N_378);
and U1389 (N_1389,N_638,N_384);
or U1390 (N_1390,N_526,N_420);
and U1391 (N_1391,N_86,N_269);
or U1392 (N_1392,N_825,N_800);
nand U1393 (N_1393,N_622,N_768);
or U1394 (N_1394,N_864,N_208);
nor U1395 (N_1395,N_206,N_252);
nor U1396 (N_1396,N_442,N_976);
or U1397 (N_1397,N_211,N_108);
and U1398 (N_1398,N_145,N_745);
and U1399 (N_1399,N_56,N_664);
xnor U1400 (N_1400,N_544,N_643);
and U1401 (N_1401,N_135,N_203);
nor U1402 (N_1402,N_840,N_634);
and U1403 (N_1403,N_871,N_747);
nand U1404 (N_1404,N_127,N_699);
nand U1405 (N_1405,N_300,N_835);
nor U1406 (N_1406,N_220,N_306);
nor U1407 (N_1407,N_791,N_931);
nor U1408 (N_1408,N_488,N_801);
nand U1409 (N_1409,N_204,N_133);
or U1410 (N_1410,N_23,N_581);
or U1411 (N_1411,N_481,N_201);
nor U1412 (N_1412,N_521,N_606);
xor U1413 (N_1413,N_471,N_31);
nor U1414 (N_1414,N_860,N_205);
or U1415 (N_1415,N_553,N_457);
or U1416 (N_1416,N_592,N_861);
nand U1417 (N_1417,N_755,N_70);
and U1418 (N_1418,N_924,N_805);
nor U1419 (N_1419,N_499,N_212);
xnor U1420 (N_1420,N_9,N_140);
nand U1421 (N_1421,N_259,N_552);
and U1422 (N_1422,N_611,N_587);
nand U1423 (N_1423,N_522,N_901);
nand U1424 (N_1424,N_66,N_780);
xnor U1425 (N_1425,N_278,N_531);
xor U1426 (N_1426,N_395,N_224);
nand U1427 (N_1427,N_147,N_527);
or U1428 (N_1428,N_297,N_672);
or U1429 (N_1429,N_225,N_496);
and U1430 (N_1430,N_270,N_601);
nand U1431 (N_1431,N_790,N_752);
and U1432 (N_1432,N_141,N_250);
nor U1433 (N_1433,N_129,N_373);
nand U1434 (N_1434,N_169,N_319);
xnor U1435 (N_1435,N_503,N_233);
nor U1436 (N_1436,N_542,N_11);
and U1437 (N_1437,N_697,N_729);
or U1438 (N_1438,N_3,N_185);
nor U1439 (N_1439,N_507,N_293);
nor U1440 (N_1440,N_434,N_136);
nor U1441 (N_1441,N_575,N_865);
or U1442 (N_1442,N_359,N_49);
xnor U1443 (N_1443,N_37,N_913);
nand U1444 (N_1444,N_255,N_779);
xnor U1445 (N_1445,N_984,N_696);
nor U1446 (N_1446,N_498,N_342);
and U1447 (N_1447,N_104,N_965);
xor U1448 (N_1448,N_102,N_266);
or U1449 (N_1449,N_89,N_822);
and U1450 (N_1450,N_124,N_329);
nor U1451 (N_1451,N_700,N_557);
or U1452 (N_1452,N_7,N_677);
nor U1453 (N_1453,N_51,N_75);
nor U1454 (N_1454,N_923,N_873);
xnor U1455 (N_1455,N_438,N_90);
xnor U1456 (N_1456,N_314,N_310);
or U1457 (N_1457,N_404,N_478);
xor U1458 (N_1458,N_588,N_477);
and U1459 (N_1459,N_197,N_919);
and U1460 (N_1460,N_598,N_630);
or U1461 (N_1461,N_175,N_670);
nand U1462 (N_1462,N_299,N_265);
xnor U1463 (N_1463,N_397,N_321);
nor U1464 (N_1464,N_367,N_956);
or U1465 (N_1465,N_411,N_904);
xnor U1466 (N_1466,N_944,N_708);
nand U1467 (N_1467,N_730,N_912);
xnor U1468 (N_1468,N_647,N_654);
or U1469 (N_1469,N_563,N_653);
nand U1470 (N_1470,N_807,N_853);
and U1471 (N_1471,N_999,N_870);
nor U1472 (N_1472,N_772,N_717);
and U1473 (N_1473,N_472,N_607);
and U1474 (N_1474,N_288,N_694);
nor U1475 (N_1475,N_113,N_432);
or U1476 (N_1476,N_926,N_838);
nor U1477 (N_1477,N_732,N_345);
nand U1478 (N_1478,N_744,N_334);
nor U1479 (N_1479,N_928,N_733);
or U1480 (N_1480,N_724,N_842);
xor U1481 (N_1481,N_793,N_59);
and U1482 (N_1482,N_282,N_680);
xor U1483 (N_1483,N_294,N_414);
nor U1484 (N_1484,N_298,N_900);
nand U1485 (N_1485,N_159,N_474);
or U1486 (N_1486,N_812,N_985);
nand U1487 (N_1487,N_577,N_111);
or U1488 (N_1488,N_151,N_736);
or U1489 (N_1489,N_262,N_979);
nor U1490 (N_1490,N_935,N_280);
or U1491 (N_1491,N_948,N_798);
nand U1492 (N_1492,N_678,N_995);
nor U1493 (N_1493,N_650,N_427);
nor U1494 (N_1494,N_903,N_93);
xor U1495 (N_1495,N_687,N_998);
or U1496 (N_1496,N_35,N_961);
and U1497 (N_1497,N_392,N_482);
nor U1498 (N_1498,N_40,N_500);
or U1499 (N_1499,N_121,N_349);
and U1500 (N_1500,N_437,N_482);
or U1501 (N_1501,N_424,N_413);
nor U1502 (N_1502,N_583,N_669);
or U1503 (N_1503,N_417,N_565);
nand U1504 (N_1504,N_807,N_840);
and U1505 (N_1505,N_477,N_198);
nand U1506 (N_1506,N_995,N_52);
and U1507 (N_1507,N_986,N_948);
xor U1508 (N_1508,N_469,N_391);
or U1509 (N_1509,N_68,N_495);
or U1510 (N_1510,N_376,N_611);
or U1511 (N_1511,N_745,N_225);
nand U1512 (N_1512,N_250,N_609);
xnor U1513 (N_1513,N_811,N_538);
nand U1514 (N_1514,N_967,N_236);
or U1515 (N_1515,N_657,N_882);
or U1516 (N_1516,N_543,N_812);
or U1517 (N_1517,N_706,N_91);
and U1518 (N_1518,N_881,N_583);
or U1519 (N_1519,N_225,N_161);
or U1520 (N_1520,N_957,N_129);
and U1521 (N_1521,N_971,N_312);
xnor U1522 (N_1522,N_78,N_262);
and U1523 (N_1523,N_985,N_806);
nand U1524 (N_1524,N_306,N_809);
nand U1525 (N_1525,N_25,N_886);
or U1526 (N_1526,N_866,N_919);
and U1527 (N_1527,N_751,N_909);
and U1528 (N_1528,N_266,N_339);
and U1529 (N_1529,N_435,N_576);
nand U1530 (N_1530,N_296,N_682);
or U1531 (N_1531,N_990,N_822);
and U1532 (N_1532,N_109,N_80);
xnor U1533 (N_1533,N_377,N_102);
and U1534 (N_1534,N_222,N_886);
and U1535 (N_1535,N_706,N_962);
xor U1536 (N_1536,N_234,N_158);
or U1537 (N_1537,N_849,N_58);
and U1538 (N_1538,N_167,N_777);
or U1539 (N_1539,N_370,N_626);
nand U1540 (N_1540,N_239,N_727);
nand U1541 (N_1541,N_843,N_946);
nand U1542 (N_1542,N_353,N_515);
or U1543 (N_1543,N_640,N_603);
nand U1544 (N_1544,N_450,N_307);
or U1545 (N_1545,N_161,N_584);
and U1546 (N_1546,N_243,N_711);
or U1547 (N_1547,N_858,N_273);
and U1548 (N_1548,N_386,N_893);
and U1549 (N_1549,N_306,N_869);
nor U1550 (N_1550,N_524,N_285);
and U1551 (N_1551,N_931,N_807);
nand U1552 (N_1552,N_316,N_575);
nand U1553 (N_1553,N_651,N_861);
nand U1554 (N_1554,N_581,N_222);
or U1555 (N_1555,N_774,N_509);
nand U1556 (N_1556,N_880,N_302);
nor U1557 (N_1557,N_8,N_919);
nor U1558 (N_1558,N_553,N_111);
and U1559 (N_1559,N_294,N_83);
nor U1560 (N_1560,N_536,N_73);
xnor U1561 (N_1561,N_870,N_968);
nand U1562 (N_1562,N_744,N_642);
nand U1563 (N_1563,N_830,N_961);
nor U1564 (N_1564,N_185,N_126);
xnor U1565 (N_1565,N_757,N_241);
or U1566 (N_1566,N_80,N_610);
nor U1567 (N_1567,N_901,N_873);
nor U1568 (N_1568,N_327,N_248);
nor U1569 (N_1569,N_241,N_729);
nor U1570 (N_1570,N_687,N_510);
xor U1571 (N_1571,N_567,N_26);
nor U1572 (N_1572,N_340,N_9);
nor U1573 (N_1573,N_651,N_709);
nand U1574 (N_1574,N_139,N_87);
nand U1575 (N_1575,N_699,N_16);
nand U1576 (N_1576,N_854,N_755);
or U1577 (N_1577,N_128,N_329);
or U1578 (N_1578,N_716,N_274);
and U1579 (N_1579,N_460,N_489);
and U1580 (N_1580,N_179,N_202);
or U1581 (N_1581,N_944,N_441);
xor U1582 (N_1582,N_62,N_627);
nor U1583 (N_1583,N_971,N_959);
xor U1584 (N_1584,N_477,N_602);
and U1585 (N_1585,N_123,N_834);
nand U1586 (N_1586,N_787,N_788);
xnor U1587 (N_1587,N_606,N_523);
xnor U1588 (N_1588,N_848,N_957);
and U1589 (N_1589,N_54,N_387);
nor U1590 (N_1590,N_60,N_155);
or U1591 (N_1591,N_176,N_507);
or U1592 (N_1592,N_579,N_288);
xor U1593 (N_1593,N_275,N_371);
nand U1594 (N_1594,N_997,N_291);
and U1595 (N_1595,N_1,N_874);
and U1596 (N_1596,N_345,N_524);
nand U1597 (N_1597,N_711,N_302);
xor U1598 (N_1598,N_826,N_915);
xor U1599 (N_1599,N_209,N_23);
and U1600 (N_1600,N_105,N_948);
and U1601 (N_1601,N_626,N_187);
nor U1602 (N_1602,N_487,N_702);
nand U1603 (N_1603,N_577,N_633);
xor U1604 (N_1604,N_481,N_583);
xor U1605 (N_1605,N_571,N_262);
and U1606 (N_1606,N_373,N_212);
nand U1607 (N_1607,N_768,N_295);
and U1608 (N_1608,N_402,N_85);
nand U1609 (N_1609,N_214,N_388);
and U1610 (N_1610,N_430,N_741);
or U1611 (N_1611,N_522,N_541);
or U1612 (N_1612,N_215,N_523);
nand U1613 (N_1613,N_474,N_744);
xor U1614 (N_1614,N_213,N_363);
nand U1615 (N_1615,N_812,N_308);
xnor U1616 (N_1616,N_806,N_731);
and U1617 (N_1617,N_863,N_98);
nor U1618 (N_1618,N_984,N_934);
or U1619 (N_1619,N_727,N_158);
xor U1620 (N_1620,N_45,N_362);
or U1621 (N_1621,N_104,N_300);
nand U1622 (N_1622,N_385,N_951);
and U1623 (N_1623,N_873,N_789);
or U1624 (N_1624,N_551,N_459);
xor U1625 (N_1625,N_454,N_967);
or U1626 (N_1626,N_708,N_2);
or U1627 (N_1627,N_264,N_32);
xor U1628 (N_1628,N_260,N_694);
or U1629 (N_1629,N_560,N_31);
nand U1630 (N_1630,N_529,N_176);
nor U1631 (N_1631,N_19,N_437);
and U1632 (N_1632,N_313,N_7);
nand U1633 (N_1633,N_46,N_420);
and U1634 (N_1634,N_702,N_444);
or U1635 (N_1635,N_423,N_49);
and U1636 (N_1636,N_114,N_438);
or U1637 (N_1637,N_342,N_737);
nand U1638 (N_1638,N_832,N_634);
xnor U1639 (N_1639,N_988,N_232);
and U1640 (N_1640,N_637,N_927);
nand U1641 (N_1641,N_899,N_861);
nand U1642 (N_1642,N_606,N_671);
and U1643 (N_1643,N_782,N_537);
nor U1644 (N_1644,N_762,N_986);
nand U1645 (N_1645,N_858,N_20);
or U1646 (N_1646,N_89,N_775);
xor U1647 (N_1647,N_376,N_864);
or U1648 (N_1648,N_474,N_936);
xor U1649 (N_1649,N_634,N_704);
and U1650 (N_1650,N_456,N_127);
xor U1651 (N_1651,N_219,N_987);
nand U1652 (N_1652,N_466,N_999);
nor U1653 (N_1653,N_472,N_353);
nor U1654 (N_1654,N_339,N_267);
and U1655 (N_1655,N_553,N_431);
xnor U1656 (N_1656,N_43,N_70);
nor U1657 (N_1657,N_228,N_112);
nor U1658 (N_1658,N_125,N_948);
nand U1659 (N_1659,N_589,N_294);
nand U1660 (N_1660,N_729,N_485);
and U1661 (N_1661,N_857,N_386);
or U1662 (N_1662,N_30,N_448);
nand U1663 (N_1663,N_436,N_697);
xor U1664 (N_1664,N_484,N_825);
nand U1665 (N_1665,N_176,N_425);
xnor U1666 (N_1666,N_94,N_23);
or U1667 (N_1667,N_618,N_621);
nor U1668 (N_1668,N_541,N_29);
nor U1669 (N_1669,N_412,N_802);
and U1670 (N_1670,N_180,N_865);
nand U1671 (N_1671,N_973,N_314);
or U1672 (N_1672,N_69,N_12);
and U1673 (N_1673,N_737,N_949);
nand U1674 (N_1674,N_692,N_608);
nand U1675 (N_1675,N_120,N_433);
and U1676 (N_1676,N_866,N_851);
xnor U1677 (N_1677,N_756,N_275);
xor U1678 (N_1678,N_460,N_983);
nor U1679 (N_1679,N_968,N_61);
xnor U1680 (N_1680,N_657,N_896);
xor U1681 (N_1681,N_976,N_465);
nand U1682 (N_1682,N_379,N_858);
xnor U1683 (N_1683,N_191,N_393);
nand U1684 (N_1684,N_106,N_693);
xor U1685 (N_1685,N_31,N_673);
nand U1686 (N_1686,N_636,N_79);
and U1687 (N_1687,N_625,N_123);
xnor U1688 (N_1688,N_237,N_863);
and U1689 (N_1689,N_598,N_992);
or U1690 (N_1690,N_489,N_415);
or U1691 (N_1691,N_309,N_122);
or U1692 (N_1692,N_110,N_480);
nor U1693 (N_1693,N_506,N_663);
and U1694 (N_1694,N_276,N_731);
nor U1695 (N_1695,N_394,N_597);
or U1696 (N_1696,N_263,N_813);
nand U1697 (N_1697,N_778,N_946);
or U1698 (N_1698,N_858,N_391);
nor U1699 (N_1699,N_816,N_111);
nand U1700 (N_1700,N_786,N_578);
xor U1701 (N_1701,N_671,N_316);
xnor U1702 (N_1702,N_602,N_622);
and U1703 (N_1703,N_72,N_421);
xnor U1704 (N_1704,N_962,N_128);
or U1705 (N_1705,N_529,N_173);
and U1706 (N_1706,N_888,N_10);
and U1707 (N_1707,N_100,N_497);
or U1708 (N_1708,N_556,N_817);
and U1709 (N_1709,N_343,N_175);
nand U1710 (N_1710,N_129,N_908);
xor U1711 (N_1711,N_492,N_572);
and U1712 (N_1712,N_909,N_38);
or U1713 (N_1713,N_237,N_834);
and U1714 (N_1714,N_136,N_705);
nor U1715 (N_1715,N_433,N_275);
nor U1716 (N_1716,N_891,N_839);
xor U1717 (N_1717,N_465,N_817);
xnor U1718 (N_1718,N_667,N_474);
nand U1719 (N_1719,N_966,N_679);
nor U1720 (N_1720,N_761,N_368);
xnor U1721 (N_1721,N_240,N_430);
and U1722 (N_1722,N_107,N_431);
nor U1723 (N_1723,N_441,N_791);
nand U1724 (N_1724,N_354,N_300);
and U1725 (N_1725,N_546,N_311);
xor U1726 (N_1726,N_489,N_32);
and U1727 (N_1727,N_814,N_20);
nor U1728 (N_1728,N_479,N_190);
or U1729 (N_1729,N_292,N_348);
nand U1730 (N_1730,N_314,N_64);
nor U1731 (N_1731,N_737,N_685);
nor U1732 (N_1732,N_860,N_690);
nor U1733 (N_1733,N_588,N_967);
or U1734 (N_1734,N_5,N_333);
and U1735 (N_1735,N_639,N_476);
and U1736 (N_1736,N_423,N_33);
xor U1737 (N_1737,N_451,N_461);
and U1738 (N_1738,N_669,N_808);
nor U1739 (N_1739,N_421,N_237);
nor U1740 (N_1740,N_829,N_757);
nand U1741 (N_1741,N_995,N_644);
or U1742 (N_1742,N_28,N_211);
or U1743 (N_1743,N_913,N_387);
nor U1744 (N_1744,N_295,N_344);
and U1745 (N_1745,N_72,N_714);
or U1746 (N_1746,N_321,N_846);
or U1747 (N_1747,N_298,N_73);
nand U1748 (N_1748,N_82,N_755);
xor U1749 (N_1749,N_578,N_122);
nor U1750 (N_1750,N_372,N_678);
and U1751 (N_1751,N_360,N_514);
nand U1752 (N_1752,N_663,N_556);
nor U1753 (N_1753,N_228,N_913);
xnor U1754 (N_1754,N_716,N_869);
nand U1755 (N_1755,N_102,N_708);
nand U1756 (N_1756,N_465,N_388);
xnor U1757 (N_1757,N_690,N_362);
nand U1758 (N_1758,N_753,N_364);
nand U1759 (N_1759,N_45,N_807);
or U1760 (N_1760,N_258,N_235);
nand U1761 (N_1761,N_247,N_394);
xor U1762 (N_1762,N_698,N_319);
nand U1763 (N_1763,N_504,N_315);
nor U1764 (N_1764,N_542,N_916);
nand U1765 (N_1765,N_434,N_779);
and U1766 (N_1766,N_395,N_308);
nor U1767 (N_1767,N_955,N_258);
and U1768 (N_1768,N_570,N_41);
nor U1769 (N_1769,N_340,N_612);
nor U1770 (N_1770,N_475,N_654);
nand U1771 (N_1771,N_21,N_282);
or U1772 (N_1772,N_264,N_9);
xnor U1773 (N_1773,N_931,N_395);
and U1774 (N_1774,N_734,N_872);
or U1775 (N_1775,N_951,N_525);
and U1776 (N_1776,N_585,N_382);
nand U1777 (N_1777,N_850,N_941);
or U1778 (N_1778,N_706,N_773);
nand U1779 (N_1779,N_713,N_733);
xnor U1780 (N_1780,N_968,N_633);
or U1781 (N_1781,N_963,N_636);
xor U1782 (N_1782,N_847,N_574);
nand U1783 (N_1783,N_561,N_14);
nand U1784 (N_1784,N_891,N_572);
nand U1785 (N_1785,N_792,N_251);
and U1786 (N_1786,N_87,N_591);
or U1787 (N_1787,N_398,N_860);
xnor U1788 (N_1788,N_243,N_64);
nor U1789 (N_1789,N_857,N_778);
nor U1790 (N_1790,N_119,N_887);
nand U1791 (N_1791,N_45,N_34);
and U1792 (N_1792,N_474,N_403);
and U1793 (N_1793,N_572,N_642);
and U1794 (N_1794,N_441,N_391);
nand U1795 (N_1795,N_221,N_241);
nand U1796 (N_1796,N_153,N_843);
nor U1797 (N_1797,N_531,N_439);
nand U1798 (N_1798,N_382,N_883);
nor U1799 (N_1799,N_347,N_917);
and U1800 (N_1800,N_391,N_471);
or U1801 (N_1801,N_722,N_537);
nand U1802 (N_1802,N_692,N_613);
xnor U1803 (N_1803,N_622,N_778);
or U1804 (N_1804,N_150,N_669);
xnor U1805 (N_1805,N_475,N_761);
xnor U1806 (N_1806,N_548,N_850);
and U1807 (N_1807,N_750,N_185);
or U1808 (N_1808,N_206,N_299);
or U1809 (N_1809,N_717,N_948);
nor U1810 (N_1810,N_960,N_154);
or U1811 (N_1811,N_618,N_816);
xnor U1812 (N_1812,N_480,N_522);
nor U1813 (N_1813,N_290,N_504);
and U1814 (N_1814,N_179,N_784);
nor U1815 (N_1815,N_0,N_232);
xor U1816 (N_1816,N_409,N_929);
nand U1817 (N_1817,N_453,N_624);
nor U1818 (N_1818,N_866,N_891);
nor U1819 (N_1819,N_512,N_141);
nand U1820 (N_1820,N_436,N_479);
and U1821 (N_1821,N_930,N_628);
nand U1822 (N_1822,N_847,N_818);
nor U1823 (N_1823,N_826,N_64);
nor U1824 (N_1824,N_215,N_237);
and U1825 (N_1825,N_992,N_900);
xnor U1826 (N_1826,N_167,N_625);
nor U1827 (N_1827,N_813,N_828);
nand U1828 (N_1828,N_868,N_960);
or U1829 (N_1829,N_831,N_189);
xnor U1830 (N_1830,N_278,N_829);
nor U1831 (N_1831,N_824,N_285);
and U1832 (N_1832,N_806,N_388);
nand U1833 (N_1833,N_491,N_941);
or U1834 (N_1834,N_170,N_817);
and U1835 (N_1835,N_307,N_554);
xor U1836 (N_1836,N_490,N_556);
nor U1837 (N_1837,N_202,N_587);
and U1838 (N_1838,N_281,N_876);
nor U1839 (N_1839,N_476,N_341);
nand U1840 (N_1840,N_524,N_310);
nand U1841 (N_1841,N_683,N_853);
and U1842 (N_1842,N_433,N_720);
nand U1843 (N_1843,N_271,N_545);
nor U1844 (N_1844,N_166,N_416);
or U1845 (N_1845,N_482,N_756);
and U1846 (N_1846,N_47,N_256);
and U1847 (N_1847,N_285,N_481);
nor U1848 (N_1848,N_904,N_746);
nand U1849 (N_1849,N_944,N_647);
nand U1850 (N_1850,N_242,N_151);
or U1851 (N_1851,N_347,N_158);
or U1852 (N_1852,N_275,N_286);
nor U1853 (N_1853,N_491,N_460);
nand U1854 (N_1854,N_155,N_23);
and U1855 (N_1855,N_404,N_867);
and U1856 (N_1856,N_66,N_672);
and U1857 (N_1857,N_796,N_992);
xor U1858 (N_1858,N_410,N_91);
or U1859 (N_1859,N_122,N_460);
xor U1860 (N_1860,N_959,N_743);
nor U1861 (N_1861,N_483,N_570);
nor U1862 (N_1862,N_369,N_490);
nand U1863 (N_1863,N_143,N_912);
xor U1864 (N_1864,N_595,N_344);
xnor U1865 (N_1865,N_809,N_481);
xor U1866 (N_1866,N_398,N_123);
nand U1867 (N_1867,N_628,N_565);
and U1868 (N_1868,N_359,N_690);
or U1869 (N_1869,N_581,N_446);
or U1870 (N_1870,N_564,N_421);
nand U1871 (N_1871,N_921,N_490);
or U1872 (N_1872,N_124,N_873);
and U1873 (N_1873,N_252,N_943);
nor U1874 (N_1874,N_512,N_467);
or U1875 (N_1875,N_104,N_45);
and U1876 (N_1876,N_764,N_780);
nand U1877 (N_1877,N_404,N_34);
nand U1878 (N_1878,N_265,N_336);
and U1879 (N_1879,N_25,N_990);
nor U1880 (N_1880,N_638,N_972);
nand U1881 (N_1881,N_866,N_854);
nor U1882 (N_1882,N_713,N_753);
or U1883 (N_1883,N_477,N_199);
and U1884 (N_1884,N_603,N_405);
xor U1885 (N_1885,N_825,N_83);
xnor U1886 (N_1886,N_304,N_474);
nor U1887 (N_1887,N_633,N_673);
nor U1888 (N_1888,N_971,N_594);
xnor U1889 (N_1889,N_831,N_935);
and U1890 (N_1890,N_742,N_755);
xnor U1891 (N_1891,N_461,N_52);
and U1892 (N_1892,N_669,N_290);
or U1893 (N_1893,N_559,N_298);
and U1894 (N_1894,N_531,N_443);
xor U1895 (N_1895,N_322,N_443);
nand U1896 (N_1896,N_197,N_689);
and U1897 (N_1897,N_873,N_560);
nand U1898 (N_1898,N_176,N_641);
nand U1899 (N_1899,N_999,N_757);
and U1900 (N_1900,N_590,N_528);
or U1901 (N_1901,N_843,N_46);
xnor U1902 (N_1902,N_815,N_771);
nor U1903 (N_1903,N_125,N_177);
nand U1904 (N_1904,N_148,N_308);
or U1905 (N_1905,N_613,N_489);
or U1906 (N_1906,N_441,N_454);
and U1907 (N_1907,N_986,N_502);
xor U1908 (N_1908,N_604,N_31);
nand U1909 (N_1909,N_273,N_638);
and U1910 (N_1910,N_792,N_498);
nor U1911 (N_1911,N_231,N_613);
xor U1912 (N_1912,N_422,N_837);
and U1913 (N_1913,N_765,N_51);
nand U1914 (N_1914,N_258,N_452);
or U1915 (N_1915,N_828,N_551);
xor U1916 (N_1916,N_715,N_302);
nor U1917 (N_1917,N_368,N_972);
nand U1918 (N_1918,N_460,N_529);
nand U1919 (N_1919,N_725,N_174);
or U1920 (N_1920,N_913,N_293);
nand U1921 (N_1921,N_937,N_437);
and U1922 (N_1922,N_834,N_69);
or U1923 (N_1923,N_199,N_744);
nand U1924 (N_1924,N_373,N_289);
and U1925 (N_1925,N_943,N_279);
or U1926 (N_1926,N_463,N_458);
xnor U1927 (N_1927,N_314,N_301);
or U1928 (N_1928,N_934,N_891);
or U1929 (N_1929,N_963,N_41);
or U1930 (N_1930,N_526,N_839);
xor U1931 (N_1931,N_143,N_107);
or U1932 (N_1932,N_168,N_751);
nand U1933 (N_1933,N_443,N_726);
or U1934 (N_1934,N_414,N_773);
nand U1935 (N_1935,N_242,N_729);
xor U1936 (N_1936,N_901,N_164);
xnor U1937 (N_1937,N_587,N_436);
nand U1938 (N_1938,N_56,N_575);
or U1939 (N_1939,N_798,N_387);
nand U1940 (N_1940,N_353,N_579);
nand U1941 (N_1941,N_552,N_687);
and U1942 (N_1942,N_829,N_630);
and U1943 (N_1943,N_963,N_648);
nor U1944 (N_1944,N_506,N_822);
or U1945 (N_1945,N_749,N_847);
xor U1946 (N_1946,N_980,N_56);
nor U1947 (N_1947,N_107,N_440);
or U1948 (N_1948,N_857,N_811);
or U1949 (N_1949,N_337,N_449);
nor U1950 (N_1950,N_707,N_854);
and U1951 (N_1951,N_411,N_382);
nand U1952 (N_1952,N_406,N_227);
nor U1953 (N_1953,N_838,N_387);
nor U1954 (N_1954,N_417,N_219);
nand U1955 (N_1955,N_141,N_552);
xor U1956 (N_1956,N_739,N_760);
xnor U1957 (N_1957,N_156,N_50);
and U1958 (N_1958,N_924,N_59);
or U1959 (N_1959,N_928,N_773);
xor U1960 (N_1960,N_286,N_365);
and U1961 (N_1961,N_442,N_134);
nand U1962 (N_1962,N_982,N_587);
nor U1963 (N_1963,N_209,N_195);
nor U1964 (N_1964,N_542,N_182);
or U1965 (N_1965,N_508,N_851);
or U1966 (N_1966,N_696,N_626);
xor U1967 (N_1967,N_564,N_581);
nor U1968 (N_1968,N_56,N_75);
nor U1969 (N_1969,N_37,N_276);
or U1970 (N_1970,N_734,N_90);
nor U1971 (N_1971,N_507,N_338);
nand U1972 (N_1972,N_91,N_685);
xor U1973 (N_1973,N_817,N_691);
or U1974 (N_1974,N_299,N_312);
xor U1975 (N_1975,N_434,N_175);
nand U1976 (N_1976,N_145,N_141);
xnor U1977 (N_1977,N_610,N_983);
or U1978 (N_1978,N_230,N_191);
nand U1979 (N_1979,N_606,N_537);
nor U1980 (N_1980,N_11,N_810);
xor U1981 (N_1981,N_388,N_658);
and U1982 (N_1982,N_508,N_625);
nor U1983 (N_1983,N_53,N_143);
and U1984 (N_1984,N_807,N_241);
or U1985 (N_1985,N_858,N_284);
xor U1986 (N_1986,N_926,N_333);
and U1987 (N_1987,N_819,N_435);
xor U1988 (N_1988,N_321,N_155);
nand U1989 (N_1989,N_444,N_316);
and U1990 (N_1990,N_243,N_756);
xor U1991 (N_1991,N_910,N_143);
or U1992 (N_1992,N_108,N_853);
nand U1993 (N_1993,N_558,N_465);
xnor U1994 (N_1994,N_709,N_471);
or U1995 (N_1995,N_245,N_686);
xnor U1996 (N_1996,N_686,N_403);
xor U1997 (N_1997,N_705,N_797);
nor U1998 (N_1998,N_932,N_634);
or U1999 (N_1999,N_641,N_425);
xnor U2000 (N_2000,N_1840,N_1721);
or U2001 (N_2001,N_1901,N_1397);
and U2002 (N_2002,N_1379,N_1073);
and U2003 (N_2003,N_1200,N_1386);
and U2004 (N_2004,N_1712,N_1274);
nor U2005 (N_2005,N_1685,N_1439);
or U2006 (N_2006,N_1490,N_1994);
nand U2007 (N_2007,N_1957,N_1308);
xnor U2008 (N_2008,N_1758,N_1521);
xnor U2009 (N_2009,N_1229,N_1430);
or U2010 (N_2010,N_1411,N_1694);
xor U2011 (N_2011,N_1865,N_1964);
or U2012 (N_2012,N_1236,N_1393);
xor U2013 (N_2013,N_1483,N_1575);
nand U2014 (N_2014,N_1950,N_1226);
or U2015 (N_2015,N_1589,N_1104);
xnor U2016 (N_2016,N_1140,N_1949);
and U2017 (N_2017,N_1193,N_1871);
or U2018 (N_2018,N_1888,N_1674);
or U2019 (N_2019,N_1070,N_1449);
nor U2020 (N_2020,N_1558,N_1458);
nor U2021 (N_2021,N_1807,N_1942);
or U2022 (N_2022,N_1413,N_1195);
nor U2023 (N_2023,N_1680,N_1736);
nor U2024 (N_2024,N_1134,N_1196);
and U2025 (N_2025,N_1216,N_1353);
xor U2026 (N_2026,N_1315,N_1659);
nand U2027 (N_2027,N_1279,N_1813);
or U2028 (N_2028,N_1287,N_1116);
nand U2029 (N_2029,N_1026,N_1811);
nand U2030 (N_2030,N_1552,N_1732);
xor U2031 (N_2031,N_1956,N_1486);
nor U2032 (N_2032,N_1820,N_1730);
and U2033 (N_2033,N_1592,N_1461);
nor U2034 (N_2034,N_1468,N_1317);
and U2035 (N_2035,N_1851,N_1122);
xnor U2036 (N_2036,N_1057,N_1874);
and U2037 (N_2037,N_1645,N_1481);
or U2038 (N_2038,N_1545,N_1740);
and U2039 (N_2039,N_1470,N_1700);
nor U2040 (N_2040,N_1955,N_1288);
or U2041 (N_2041,N_1384,N_1002);
xnor U2042 (N_2042,N_1329,N_1425);
and U2043 (N_2043,N_1444,N_1298);
xnor U2044 (N_2044,N_1445,N_1150);
and U2045 (N_2045,N_1078,N_1414);
xor U2046 (N_2046,N_1107,N_1068);
and U2047 (N_2047,N_1403,N_1181);
and U2048 (N_2048,N_1499,N_1126);
xnor U2049 (N_2049,N_1103,N_1512);
and U2050 (N_2050,N_1669,N_1203);
or U2051 (N_2051,N_1058,N_1176);
nor U2052 (N_2052,N_1014,N_1015);
and U2053 (N_2053,N_1245,N_1451);
or U2054 (N_2054,N_1780,N_1289);
and U2055 (N_2055,N_1997,N_1050);
or U2056 (N_2056,N_1806,N_1038);
nor U2057 (N_2057,N_1812,N_1160);
xnor U2058 (N_2058,N_1460,N_1970);
xor U2059 (N_2059,N_1559,N_1191);
nand U2060 (N_2060,N_1500,N_1830);
nand U2061 (N_2061,N_1376,N_1036);
xnor U2062 (N_2062,N_1961,N_1968);
and U2063 (N_2063,N_1585,N_1642);
or U2064 (N_2064,N_1277,N_1098);
xor U2065 (N_2065,N_1549,N_1695);
and U2066 (N_2066,N_1704,N_1082);
nand U2067 (N_2067,N_1737,N_1377);
nand U2068 (N_2068,N_1917,N_1914);
or U2069 (N_2069,N_1012,N_1013);
xor U2070 (N_2070,N_1782,N_1182);
or U2071 (N_2071,N_1156,N_1869);
and U2072 (N_2072,N_1048,N_1728);
and U2073 (N_2073,N_1554,N_1705);
or U2074 (N_2074,N_1853,N_1819);
or U2075 (N_2075,N_1709,N_1456);
nand U2076 (N_2076,N_1231,N_1551);
and U2077 (N_2077,N_1578,N_1748);
nor U2078 (N_2078,N_1235,N_1804);
nor U2079 (N_2079,N_1305,N_1538);
nand U2080 (N_2080,N_1530,N_1971);
and U2081 (N_2081,N_1518,N_1606);
and U2082 (N_2082,N_1771,N_1412);
and U2083 (N_2083,N_1472,N_1635);
and U2084 (N_2084,N_1844,N_1432);
or U2085 (N_2085,N_1255,N_1332);
nand U2086 (N_2086,N_1357,N_1516);
or U2087 (N_2087,N_1876,N_1212);
nor U2088 (N_2088,N_1524,N_1318);
and U2089 (N_2089,N_1506,N_1570);
xnor U2090 (N_2090,N_1881,N_1679);
and U2091 (N_2091,N_1371,N_1690);
nand U2092 (N_2092,N_1161,N_1568);
xnor U2093 (N_2093,N_1136,N_1110);
or U2094 (N_2094,N_1798,N_1613);
nand U2095 (N_2095,N_1263,N_1459);
nand U2096 (N_2096,N_1701,N_1742);
nor U2097 (N_2097,N_1214,N_1502);
xor U2098 (N_2098,N_1131,N_1598);
or U2099 (N_2099,N_1826,N_1662);
or U2100 (N_2100,N_1375,N_1883);
xnor U2101 (N_2101,N_1610,N_1290);
xor U2102 (N_2102,N_1223,N_1623);
or U2103 (N_2103,N_1567,N_1667);
and U2104 (N_2104,N_1010,N_1462);
xnor U2105 (N_2105,N_1562,N_1640);
nor U2106 (N_2106,N_1841,N_1972);
nor U2107 (N_2107,N_1650,N_1785);
xnor U2108 (N_2108,N_1696,N_1463);
nand U2109 (N_2109,N_1442,N_1842);
nor U2110 (N_2110,N_1920,N_1564);
or U2111 (N_2111,N_1626,N_1615);
nor U2112 (N_2112,N_1147,N_1648);
or U2113 (N_2113,N_1052,N_1275);
nand U2114 (N_2114,N_1396,N_1741);
xor U2115 (N_2115,N_1511,N_1154);
or U2116 (N_2116,N_1508,N_1624);
xnor U2117 (N_2117,N_1781,N_1565);
and U2118 (N_2118,N_1494,N_1264);
or U2119 (N_2119,N_1051,N_1661);
or U2120 (N_2120,N_1049,N_1368);
nand U2121 (N_2121,N_1580,N_1127);
xor U2122 (N_2122,N_1102,N_1985);
or U2123 (N_2123,N_1443,N_1649);
or U2124 (N_2124,N_1911,N_1774);
nor U2125 (N_2125,N_1866,N_1960);
or U2126 (N_2126,N_1039,N_1501);
or U2127 (N_2127,N_1334,N_1984);
xor U2128 (N_2128,N_1145,N_1975);
or U2129 (N_2129,N_1601,N_1827);
nand U2130 (N_2130,N_1587,N_1054);
nand U2131 (N_2131,N_1832,N_1590);
nor U2132 (N_2132,N_1787,N_1707);
nor U2133 (N_2133,N_1055,N_1006);
xnor U2134 (N_2134,N_1687,N_1143);
and U2135 (N_2135,N_1689,N_1810);
or U2136 (N_2136,N_1605,N_1204);
xnor U2137 (N_2137,N_1187,N_1873);
nor U2138 (N_2138,N_1849,N_1333);
and U2139 (N_2139,N_1431,N_1170);
xnor U2140 (N_2140,N_1692,N_1011);
nor U2141 (N_2141,N_1325,N_1388);
nor U2142 (N_2142,N_1285,N_1000);
nor U2143 (N_2143,N_1427,N_1542);
nor U2144 (N_2144,N_1988,N_1335);
nor U2145 (N_2145,N_1703,N_1561);
and U2146 (N_2146,N_1378,N_1752);
nor U2147 (N_2147,N_1789,N_1952);
and U2148 (N_2148,N_1928,N_1850);
and U2149 (N_2149,N_1746,N_1409);
xor U2150 (N_2150,N_1714,N_1165);
xnor U2151 (N_2151,N_1341,N_1278);
or U2152 (N_2152,N_1654,N_1576);
or U2153 (N_2153,N_1360,N_1428);
xnor U2154 (N_2154,N_1517,N_1090);
xnor U2155 (N_2155,N_1373,N_1618);
and U2156 (N_2156,N_1467,N_1025);
or U2157 (N_2157,N_1611,N_1938);
and U2158 (N_2158,N_1905,N_1981);
and U2159 (N_2159,N_1340,N_1089);
and U2160 (N_2160,N_1847,N_1603);
xnor U2161 (N_2161,N_1405,N_1183);
nand U2162 (N_2162,N_1683,N_1254);
or U2163 (N_2163,N_1824,N_1059);
nand U2164 (N_2164,N_1982,N_1722);
xor U2165 (N_2165,N_1902,N_1327);
or U2166 (N_2166,N_1838,N_1673);
xnor U2167 (N_2167,N_1480,N_1908);
nand U2168 (N_2168,N_1529,N_1628);
nor U2169 (N_2169,N_1505,N_1507);
nor U2170 (N_2170,N_1441,N_1056);
or U2171 (N_2171,N_1166,N_1477);
nor U2172 (N_2172,N_1852,N_1138);
or U2173 (N_2173,N_1113,N_1178);
nor U2174 (N_2174,N_1316,N_1205);
nor U2175 (N_2175,N_1239,N_1020);
or U2176 (N_2176,N_1930,N_1915);
and U2177 (N_2177,N_1326,N_1944);
nor U2178 (N_2178,N_1718,N_1794);
nand U2179 (N_2179,N_1488,N_1045);
nor U2180 (N_2180,N_1571,N_1647);
or U2181 (N_2181,N_1632,N_1791);
nand U2182 (N_2182,N_1805,N_1676);
nand U2183 (N_2183,N_1818,N_1410);
nor U2184 (N_2184,N_1756,N_1162);
and U2185 (N_2185,N_1893,N_1111);
xnor U2186 (N_2186,N_1622,N_1969);
nor U2187 (N_2187,N_1777,N_1723);
nand U2188 (N_2188,N_1983,N_1114);
nor U2189 (N_2189,N_1190,N_1872);
nor U2190 (N_2190,N_1243,N_1321);
nor U2191 (N_2191,N_1244,N_1855);
nand U2192 (N_2192,N_1351,N_1836);
and U2193 (N_2193,N_1670,N_1990);
nand U2194 (N_2194,N_1927,N_1715);
nor U2195 (N_2195,N_1485,N_1387);
nand U2196 (N_2196,N_1044,N_1817);
nor U2197 (N_2197,N_1588,N_1475);
xor U2198 (N_2198,N_1929,N_1764);
xnor U2199 (N_2199,N_1232,N_1033);
xnor U2200 (N_2200,N_1260,N_1031);
nand U2201 (N_2201,N_1354,N_1213);
nand U2202 (N_2202,N_1061,N_1312);
and U2203 (N_2203,N_1457,N_1802);
xnor U2204 (N_2204,N_1398,N_1713);
xnor U2205 (N_2205,N_1816,N_1251);
or U2206 (N_2206,N_1133,N_1892);
and U2207 (N_2207,N_1900,N_1967);
nand U2208 (N_2208,N_1407,N_1270);
and U2209 (N_2209,N_1455,N_1898);
xnor U2210 (N_2210,N_1479,N_1656);
nor U2211 (N_2211,N_1537,N_1364);
and U2212 (N_2212,N_1084,N_1450);
or U2213 (N_2213,N_1295,N_1256);
xnor U2214 (N_2214,N_1630,N_1599);
nand U2215 (N_2215,N_1003,N_1751);
nand U2216 (N_2216,N_1418,N_1870);
and U2217 (N_2217,N_1429,N_1207);
or U2218 (N_2218,N_1158,N_1215);
and U2219 (N_2219,N_1658,N_1867);
nor U2220 (N_2220,N_1907,N_1636);
and U2221 (N_2221,N_1725,N_1009);
nand U2222 (N_2222,N_1148,N_1989);
and U2223 (N_2223,N_1421,N_1365);
or U2224 (N_2224,N_1030,N_1453);
nand U2225 (N_2225,N_1047,N_1579);
nor U2226 (N_2226,N_1536,N_1099);
xnor U2227 (N_2227,N_1228,N_1886);
xnor U2228 (N_2228,N_1532,N_1217);
nand U2229 (N_2229,N_1664,N_1064);
and U2230 (N_2230,N_1197,N_1046);
and U2231 (N_2231,N_1541,N_1834);
nor U2232 (N_2232,N_1682,N_1471);
nand U2233 (N_2233,N_1999,N_1300);
nor U2234 (N_2234,N_1080,N_1408);
nand U2235 (N_2235,N_1324,N_1001);
nor U2236 (N_2236,N_1706,N_1271);
or U2237 (N_2237,N_1627,N_1346);
xor U2238 (N_2238,N_1454,N_1916);
or U2239 (N_2239,N_1868,N_1977);
or U2240 (N_2240,N_1426,N_1772);
nand U2241 (N_2241,N_1992,N_1691);
and U2242 (N_2242,N_1302,N_1828);
xor U2243 (N_2243,N_1959,N_1759);
or U2244 (N_2244,N_1864,N_1760);
nor U2245 (N_2245,N_1753,N_1284);
nor U2246 (N_2246,N_1710,N_1222);
nand U2247 (N_2247,N_1209,N_1120);
nand U2248 (N_2248,N_1600,N_1738);
xnor U2249 (N_2249,N_1750,N_1544);
or U2250 (N_2250,N_1037,N_1801);
nand U2251 (N_2251,N_1092,N_1282);
or U2252 (N_2252,N_1087,N_1489);
nor U2253 (N_2253,N_1076,N_1577);
nor U2254 (N_2254,N_1436,N_1607);
nor U2255 (N_2255,N_1109,N_1996);
or U2256 (N_2256,N_1422,N_1124);
nand U2257 (N_2257,N_1677,N_1394);
and U2258 (N_2258,N_1757,N_1616);
nand U2259 (N_2259,N_1857,N_1954);
xnor U2260 (N_2260,N_1447,N_1743);
and U2261 (N_2261,N_1390,N_1581);
nor U2262 (N_2262,N_1185,N_1234);
xor U2263 (N_2263,N_1206,N_1117);
nor U2264 (N_2264,N_1604,N_1392);
or U2265 (N_2265,N_1848,N_1509);
xor U2266 (N_2266,N_1591,N_1169);
or U2267 (N_2267,N_1097,N_1620);
or U2268 (N_2268,N_1446,N_1434);
nor U2269 (N_2269,N_1582,N_1086);
or U2270 (N_2270,N_1720,N_1221);
or U2271 (N_2271,N_1843,N_1478);
and U2272 (N_2272,N_1602,N_1612);
and U2273 (N_2273,N_1947,N_1291);
or U2274 (N_2274,N_1739,N_1912);
nand U2275 (N_2275,N_1194,N_1309);
nor U2276 (N_2276,N_1043,N_1174);
nand U2277 (N_2277,N_1540,N_1168);
and U2278 (N_2278,N_1328,N_1884);
xnor U2279 (N_2279,N_1797,N_1795);
or U2280 (N_2280,N_1527,N_1381);
nor U2281 (N_2281,N_1313,N_1688);
and U2282 (N_2282,N_1246,N_1671);
and U2283 (N_2283,N_1367,N_1889);
and U2284 (N_2284,N_1262,N_1699);
or U2285 (N_2285,N_1796,N_1770);
nor U2286 (N_2286,N_1448,N_1072);
nand U2287 (N_2287,N_1531,N_1171);
or U2288 (N_2288,N_1681,N_1923);
xnor U2289 (N_2289,N_1586,N_1678);
nor U2290 (N_2290,N_1660,N_1331);
nor U2291 (N_2291,N_1583,N_1402);
and U2292 (N_2292,N_1768,N_1619);
nand U2293 (N_2293,N_1273,N_1130);
and U2294 (N_2294,N_1356,N_1909);
and U2295 (N_2295,N_1941,N_1858);
nand U2296 (N_2296,N_1093,N_1067);
xor U2297 (N_2297,N_1032,N_1380);
or U2298 (N_2298,N_1115,N_1355);
nand U2299 (N_2299,N_1361,N_1890);
or U2300 (N_2300,N_1629,N_1281);
or U2301 (N_2301,N_1904,N_1337);
nand U2302 (N_2302,N_1895,N_1118);
nor U2303 (N_2303,N_1711,N_1783);
nor U2304 (N_2304,N_1822,N_1307);
xnor U2305 (N_2305,N_1861,N_1776);
nand U2306 (N_2306,N_1100,N_1137);
or U2307 (N_2307,N_1369,N_1053);
xor U2308 (N_2308,N_1155,N_1135);
xnor U2309 (N_2309,N_1625,N_1153);
xor U2310 (N_2310,N_1762,N_1513);
and U2311 (N_2311,N_1733,N_1250);
and U2312 (N_2312,N_1469,N_1979);
or U2313 (N_2313,N_1555,N_1497);
xnor U2314 (N_2314,N_1966,N_1063);
and U2315 (N_2315,N_1060,N_1062);
nor U2316 (N_2316,N_1877,N_1306);
and U2317 (N_2317,N_1343,N_1350);
nand U2318 (N_2318,N_1347,N_1878);
and U2319 (N_2319,N_1261,N_1765);
and U2320 (N_2320,N_1198,N_1021);
nor U2321 (N_2321,N_1465,N_1790);
xor U2322 (N_2322,N_1083,N_1814);
nor U2323 (N_2323,N_1493,N_1303);
xor U2324 (N_2324,N_1438,N_1069);
nor U2325 (N_2325,N_1077,N_1096);
nand U2326 (N_2326,N_1293,N_1793);
xor U2327 (N_2327,N_1815,N_1906);
nand U2328 (N_2328,N_1514,N_1024);
nor U2329 (N_2329,N_1976,N_1294);
and U2330 (N_2330,N_1833,N_1227);
or U2331 (N_2331,N_1385,N_1731);
xor U2332 (N_2332,N_1775,N_1939);
nor U2333 (N_2333,N_1735,N_1786);
xor U2334 (N_2334,N_1931,N_1440);
and U2335 (N_2335,N_1755,N_1520);
nor U2336 (N_2336,N_1225,N_1141);
and U2337 (N_2337,N_1717,N_1769);
nand U2338 (N_2338,N_1152,N_1320);
nor U2339 (N_2339,N_1835,N_1533);
nor U2340 (N_2340,N_1419,N_1749);
or U2341 (N_2341,N_1362,N_1363);
nand U2342 (N_2342,N_1323,N_1860);
xnor U2343 (N_2343,N_1416,N_1614);
xor U2344 (N_2344,N_1899,N_1885);
nand U2345 (N_2345,N_1473,N_1016);
nand U2346 (N_2346,N_1633,N_1259);
xnor U2347 (N_2347,N_1638,N_1359);
nand U2348 (N_2348,N_1784,N_1747);
nor U2349 (N_2349,N_1823,N_1569);
nand U2350 (N_2350,N_1252,N_1698);
nor U2351 (N_2351,N_1727,N_1167);
or U2352 (N_2352,N_1637,N_1729);
nor U2353 (N_2353,N_1951,N_1437);
and U2354 (N_2354,N_1065,N_1932);
nor U2355 (N_2355,N_1767,N_1593);
xor U2356 (N_2356,N_1267,N_1945);
nand U2357 (N_2357,N_1894,N_1027);
nor U2358 (N_2358,N_1946,N_1401);
and U2359 (N_2359,N_1123,N_1464);
nor U2360 (N_2360,N_1854,N_1404);
xnor U2361 (N_2361,N_1474,N_1184);
and U2362 (N_2362,N_1339,N_1035);
and U2363 (N_2363,N_1066,N_1041);
or U2364 (N_2364,N_1523,N_1879);
or U2365 (N_2365,N_1887,N_1672);
xor U2366 (N_2366,N_1304,N_1655);
nor U2367 (N_2367,N_1292,N_1991);
nor U2368 (N_2368,N_1202,N_1119);
xnor U2369 (N_2369,N_1344,N_1272);
xnor U2370 (N_2370,N_1719,N_1631);
xor U2371 (N_2371,N_1934,N_1744);
and U2372 (N_2372,N_1257,N_1773);
nand U2373 (N_2373,N_1210,N_1374);
and U2374 (N_2374,N_1283,N_1644);
or U2375 (N_2375,N_1132,N_1495);
or U2376 (N_2376,N_1510,N_1745);
xor U2377 (N_2377,N_1597,N_1503);
nor U2378 (N_2378,N_1566,N_1172);
or U2379 (N_2379,N_1803,N_1484);
or U2380 (N_2380,N_1856,N_1233);
xor U2381 (N_2381,N_1336,N_1238);
or U2382 (N_2382,N_1845,N_1543);
xor U2383 (N_2383,N_1891,N_1668);
nor U2384 (N_2384,N_1995,N_1539);
or U2385 (N_2385,N_1573,N_1240);
and U2386 (N_2386,N_1498,N_1417);
or U2387 (N_2387,N_1652,N_1666);
xor U2388 (N_2388,N_1548,N_1296);
or U2389 (N_2389,N_1963,N_1400);
nor U2390 (N_2390,N_1595,N_1547);
nor U2391 (N_2391,N_1253,N_1846);
nand U2392 (N_2392,N_1863,N_1535);
nand U2393 (N_2393,N_1974,N_1121);
and U2394 (N_2394,N_1391,N_1837);
or U2395 (N_2395,N_1125,N_1105);
or U2396 (N_2396,N_1079,N_1268);
nand U2397 (N_2397,N_1761,N_1128);
or U2398 (N_2398,N_1452,N_1247);
nor U2399 (N_2399,N_1903,N_1809);
nand U2400 (N_2400,N_1726,N_1651);
and U2401 (N_2401,N_1189,N_1766);
nand U2402 (N_2402,N_1342,N_1301);
nand U2403 (N_2403,N_1175,N_1617);
nor U2404 (N_2404,N_1896,N_1641);
and U2405 (N_2405,N_1799,N_1962);
nor U2406 (N_2406,N_1504,N_1424);
nand U2407 (N_2407,N_1319,N_1112);
and U2408 (N_2408,N_1926,N_1973);
or U2409 (N_2409,N_1101,N_1609);
and U2410 (N_2410,N_1179,N_1230);
nor U2411 (N_2411,N_1657,N_1875);
xor U2412 (N_2412,N_1399,N_1008);
nand U2413 (N_2413,N_1311,N_1173);
xnor U2414 (N_2414,N_1095,N_1476);
nor U2415 (N_2415,N_1314,N_1146);
xnor U2416 (N_2416,N_1708,N_1734);
nor U2417 (N_2417,N_1919,N_1716);
nand U2418 (N_2418,N_1693,N_1019);
or U2419 (N_2419,N_1349,N_1831);
and U2420 (N_2420,N_1142,N_1792);
nand U2421 (N_2421,N_1151,N_1943);
nand U2422 (N_2422,N_1071,N_1491);
nand U2423 (N_2423,N_1525,N_1897);
nor U2424 (N_2424,N_1022,N_1435);
xor U2425 (N_2425,N_1526,N_1643);
and U2426 (N_2426,N_1201,N_1953);
nand U2427 (N_2427,N_1211,N_1395);
and U2428 (N_2428,N_1348,N_1940);
nand U2429 (N_2429,N_1042,N_1040);
xnor U2430 (N_2430,N_1933,N_1163);
and U2431 (N_2431,N_1948,N_1186);
or U2432 (N_2432,N_1882,N_1675);
and U2433 (N_2433,N_1352,N_1383);
nand U2434 (N_2434,N_1754,N_1998);
or U2435 (N_2435,N_1553,N_1560);
and U2436 (N_2436,N_1515,N_1986);
xnor U2437 (N_2437,N_1023,N_1338);
xnor U2438 (N_2438,N_1965,N_1330);
nand U2439 (N_2439,N_1005,N_1007);
and U2440 (N_2440,N_1653,N_1546);
nand U2441 (N_2441,N_1596,N_1913);
nor U2442 (N_2442,N_1322,N_1249);
xnor U2443 (N_2443,N_1646,N_1594);
or U2444 (N_2444,N_1763,N_1074);
xnor U2445 (N_2445,N_1808,N_1269);
and U2446 (N_2446,N_1534,N_1528);
xor U2447 (N_2447,N_1423,N_1129);
nand U2448 (N_2448,N_1925,N_1094);
and U2449 (N_2449,N_1149,N_1496);
nor U2450 (N_2450,N_1265,N_1788);
and U2451 (N_2451,N_1188,N_1825);
xnor U2452 (N_2452,N_1157,N_1550);
or U2453 (N_2453,N_1563,N_1519);
xnor U2454 (N_2454,N_1993,N_1639);
xor U2455 (N_2455,N_1081,N_1584);
xnor U2456 (N_2456,N_1937,N_1702);
nor U2457 (N_2457,N_1075,N_1034);
or U2458 (N_2458,N_1958,N_1492);
nor U2459 (N_2459,N_1574,N_1139);
or U2460 (N_2460,N_1286,N_1987);
nor U2461 (N_2461,N_1686,N_1415);
and U2462 (N_2462,N_1935,N_1389);
nor U2463 (N_2463,N_1557,N_1663);
nand U2464 (N_2464,N_1220,N_1487);
xor U2465 (N_2465,N_1778,N_1237);
or U2466 (N_2466,N_1004,N_1144);
nor U2467 (N_2467,N_1522,N_1779);
xor U2468 (N_2468,N_1922,N_1108);
and U2469 (N_2469,N_1180,N_1634);
xnor U2470 (N_2470,N_1345,N_1018);
nor U2471 (N_2471,N_1241,N_1106);
xnor U2472 (N_2472,N_1258,N_1088);
or U2473 (N_2473,N_1433,N_1936);
xnor U2474 (N_2474,N_1910,N_1028);
or U2475 (N_2475,N_1420,N_1299);
xor U2476 (N_2476,N_1821,N_1224);
nor U2477 (N_2477,N_1192,N_1370);
nand U2478 (N_2478,N_1310,N_1017);
nor U2479 (N_2479,N_1859,N_1372);
nand U2480 (N_2480,N_1358,N_1621);
xnor U2481 (N_2481,N_1482,N_1572);
nor U2482 (N_2482,N_1164,N_1862);
and U2483 (N_2483,N_1159,N_1091);
nand U2484 (N_2484,N_1366,N_1924);
nand U2485 (N_2485,N_1556,N_1085);
and U2486 (N_2486,N_1829,N_1208);
xnor U2487 (N_2487,N_1029,N_1980);
xor U2488 (N_2488,N_1219,N_1978);
nand U2489 (N_2489,N_1684,N_1724);
xnor U2490 (N_2490,N_1608,N_1800);
xor U2491 (N_2491,N_1665,N_1697);
or U2492 (N_2492,N_1466,N_1177);
nor U2493 (N_2493,N_1297,N_1242);
nor U2494 (N_2494,N_1880,N_1199);
or U2495 (N_2495,N_1280,N_1839);
xor U2496 (N_2496,N_1918,N_1382);
nor U2497 (N_2497,N_1266,N_1248);
xnor U2498 (N_2498,N_1406,N_1276);
nand U2499 (N_2499,N_1921,N_1218);
nand U2500 (N_2500,N_1181,N_1234);
xnor U2501 (N_2501,N_1824,N_1974);
xor U2502 (N_2502,N_1145,N_1157);
nand U2503 (N_2503,N_1606,N_1906);
or U2504 (N_2504,N_1914,N_1220);
nor U2505 (N_2505,N_1866,N_1775);
or U2506 (N_2506,N_1547,N_1216);
nor U2507 (N_2507,N_1018,N_1264);
xor U2508 (N_2508,N_1764,N_1039);
xnor U2509 (N_2509,N_1136,N_1791);
or U2510 (N_2510,N_1323,N_1742);
or U2511 (N_2511,N_1633,N_1531);
and U2512 (N_2512,N_1034,N_1762);
xor U2513 (N_2513,N_1171,N_1444);
nand U2514 (N_2514,N_1852,N_1960);
xnor U2515 (N_2515,N_1751,N_1848);
or U2516 (N_2516,N_1279,N_1305);
nor U2517 (N_2517,N_1249,N_1054);
or U2518 (N_2518,N_1903,N_1402);
and U2519 (N_2519,N_1827,N_1530);
nand U2520 (N_2520,N_1580,N_1573);
nand U2521 (N_2521,N_1048,N_1909);
or U2522 (N_2522,N_1180,N_1145);
and U2523 (N_2523,N_1832,N_1953);
nand U2524 (N_2524,N_1818,N_1931);
xor U2525 (N_2525,N_1793,N_1881);
nor U2526 (N_2526,N_1478,N_1308);
and U2527 (N_2527,N_1163,N_1127);
or U2528 (N_2528,N_1147,N_1971);
nor U2529 (N_2529,N_1914,N_1638);
nand U2530 (N_2530,N_1566,N_1171);
nor U2531 (N_2531,N_1965,N_1138);
and U2532 (N_2532,N_1405,N_1045);
or U2533 (N_2533,N_1158,N_1838);
nor U2534 (N_2534,N_1618,N_1709);
nor U2535 (N_2535,N_1104,N_1622);
and U2536 (N_2536,N_1777,N_1561);
or U2537 (N_2537,N_1689,N_1536);
or U2538 (N_2538,N_1592,N_1853);
xnor U2539 (N_2539,N_1323,N_1854);
nor U2540 (N_2540,N_1443,N_1092);
xor U2541 (N_2541,N_1131,N_1595);
or U2542 (N_2542,N_1704,N_1058);
and U2543 (N_2543,N_1445,N_1024);
nand U2544 (N_2544,N_1097,N_1089);
nand U2545 (N_2545,N_1166,N_1378);
and U2546 (N_2546,N_1431,N_1996);
nor U2547 (N_2547,N_1480,N_1675);
xnor U2548 (N_2548,N_1581,N_1027);
nor U2549 (N_2549,N_1708,N_1536);
nor U2550 (N_2550,N_1336,N_1301);
xor U2551 (N_2551,N_1315,N_1181);
or U2552 (N_2552,N_1266,N_1611);
nor U2553 (N_2553,N_1734,N_1353);
or U2554 (N_2554,N_1235,N_1381);
and U2555 (N_2555,N_1165,N_1319);
nor U2556 (N_2556,N_1712,N_1567);
and U2557 (N_2557,N_1379,N_1206);
nor U2558 (N_2558,N_1361,N_1272);
nor U2559 (N_2559,N_1415,N_1237);
or U2560 (N_2560,N_1346,N_1775);
and U2561 (N_2561,N_1419,N_1280);
nand U2562 (N_2562,N_1104,N_1779);
nor U2563 (N_2563,N_1618,N_1990);
xor U2564 (N_2564,N_1971,N_1816);
nand U2565 (N_2565,N_1656,N_1742);
and U2566 (N_2566,N_1126,N_1287);
xor U2567 (N_2567,N_1493,N_1268);
or U2568 (N_2568,N_1163,N_1780);
xnor U2569 (N_2569,N_1713,N_1547);
nand U2570 (N_2570,N_1364,N_1581);
nor U2571 (N_2571,N_1206,N_1144);
nand U2572 (N_2572,N_1306,N_1950);
nand U2573 (N_2573,N_1195,N_1019);
and U2574 (N_2574,N_1943,N_1541);
xor U2575 (N_2575,N_1626,N_1033);
xor U2576 (N_2576,N_1034,N_1174);
nor U2577 (N_2577,N_1220,N_1637);
nor U2578 (N_2578,N_1222,N_1906);
or U2579 (N_2579,N_1251,N_1580);
nor U2580 (N_2580,N_1353,N_1953);
nor U2581 (N_2581,N_1422,N_1116);
or U2582 (N_2582,N_1029,N_1198);
or U2583 (N_2583,N_1217,N_1004);
xnor U2584 (N_2584,N_1175,N_1713);
nor U2585 (N_2585,N_1537,N_1571);
and U2586 (N_2586,N_1278,N_1287);
xnor U2587 (N_2587,N_1463,N_1432);
and U2588 (N_2588,N_1934,N_1408);
nand U2589 (N_2589,N_1586,N_1831);
or U2590 (N_2590,N_1569,N_1219);
or U2591 (N_2591,N_1011,N_1879);
or U2592 (N_2592,N_1835,N_1559);
or U2593 (N_2593,N_1011,N_1297);
or U2594 (N_2594,N_1896,N_1506);
xor U2595 (N_2595,N_1182,N_1004);
xnor U2596 (N_2596,N_1686,N_1183);
and U2597 (N_2597,N_1148,N_1491);
nor U2598 (N_2598,N_1743,N_1958);
or U2599 (N_2599,N_1368,N_1301);
and U2600 (N_2600,N_1945,N_1330);
xnor U2601 (N_2601,N_1784,N_1631);
nand U2602 (N_2602,N_1369,N_1359);
and U2603 (N_2603,N_1626,N_1262);
or U2604 (N_2604,N_1561,N_1391);
or U2605 (N_2605,N_1825,N_1032);
nor U2606 (N_2606,N_1006,N_1323);
xor U2607 (N_2607,N_1827,N_1990);
or U2608 (N_2608,N_1449,N_1319);
or U2609 (N_2609,N_1734,N_1685);
nand U2610 (N_2610,N_1122,N_1164);
and U2611 (N_2611,N_1112,N_1750);
and U2612 (N_2612,N_1271,N_1088);
nor U2613 (N_2613,N_1943,N_1780);
or U2614 (N_2614,N_1948,N_1610);
nor U2615 (N_2615,N_1041,N_1349);
nand U2616 (N_2616,N_1633,N_1235);
nor U2617 (N_2617,N_1918,N_1609);
xor U2618 (N_2618,N_1125,N_1357);
nor U2619 (N_2619,N_1711,N_1202);
nor U2620 (N_2620,N_1013,N_1405);
nor U2621 (N_2621,N_1741,N_1106);
and U2622 (N_2622,N_1987,N_1239);
xor U2623 (N_2623,N_1967,N_1872);
xor U2624 (N_2624,N_1850,N_1893);
nand U2625 (N_2625,N_1005,N_1187);
xnor U2626 (N_2626,N_1696,N_1205);
nor U2627 (N_2627,N_1415,N_1264);
or U2628 (N_2628,N_1011,N_1625);
xnor U2629 (N_2629,N_1109,N_1826);
xnor U2630 (N_2630,N_1578,N_1935);
xnor U2631 (N_2631,N_1913,N_1678);
and U2632 (N_2632,N_1896,N_1202);
nand U2633 (N_2633,N_1763,N_1902);
or U2634 (N_2634,N_1621,N_1778);
nand U2635 (N_2635,N_1201,N_1718);
nor U2636 (N_2636,N_1676,N_1875);
or U2637 (N_2637,N_1757,N_1014);
and U2638 (N_2638,N_1566,N_1489);
xnor U2639 (N_2639,N_1771,N_1893);
and U2640 (N_2640,N_1119,N_1514);
nor U2641 (N_2641,N_1279,N_1190);
or U2642 (N_2642,N_1353,N_1272);
nand U2643 (N_2643,N_1933,N_1877);
or U2644 (N_2644,N_1692,N_1477);
or U2645 (N_2645,N_1591,N_1618);
or U2646 (N_2646,N_1091,N_1010);
or U2647 (N_2647,N_1026,N_1595);
nand U2648 (N_2648,N_1273,N_1397);
nand U2649 (N_2649,N_1646,N_1012);
nand U2650 (N_2650,N_1033,N_1112);
xor U2651 (N_2651,N_1781,N_1541);
nor U2652 (N_2652,N_1988,N_1914);
nor U2653 (N_2653,N_1948,N_1114);
and U2654 (N_2654,N_1854,N_1223);
xnor U2655 (N_2655,N_1514,N_1262);
nor U2656 (N_2656,N_1394,N_1409);
nand U2657 (N_2657,N_1098,N_1501);
or U2658 (N_2658,N_1559,N_1918);
nand U2659 (N_2659,N_1856,N_1793);
and U2660 (N_2660,N_1796,N_1748);
xor U2661 (N_2661,N_1187,N_1390);
or U2662 (N_2662,N_1609,N_1136);
nand U2663 (N_2663,N_1795,N_1681);
or U2664 (N_2664,N_1956,N_1550);
or U2665 (N_2665,N_1128,N_1649);
xor U2666 (N_2666,N_1463,N_1590);
and U2667 (N_2667,N_1064,N_1462);
nand U2668 (N_2668,N_1844,N_1324);
nand U2669 (N_2669,N_1128,N_1084);
nand U2670 (N_2670,N_1085,N_1547);
nor U2671 (N_2671,N_1375,N_1556);
nand U2672 (N_2672,N_1270,N_1549);
nor U2673 (N_2673,N_1843,N_1273);
xnor U2674 (N_2674,N_1306,N_1710);
xnor U2675 (N_2675,N_1740,N_1994);
nor U2676 (N_2676,N_1954,N_1085);
or U2677 (N_2677,N_1461,N_1495);
nor U2678 (N_2678,N_1590,N_1327);
xor U2679 (N_2679,N_1265,N_1588);
nand U2680 (N_2680,N_1942,N_1609);
or U2681 (N_2681,N_1492,N_1183);
nand U2682 (N_2682,N_1512,N_1180);
nand U2683 (N_2683,N_1368,N_1276);
nand U2684 (N_2684,N_1568,N_1412);
and U2685 (N_2685,N_1056,N_1589);
nand U2686 (N_2686,N_1167,N_1443);
or U2687 (N_2687,N_1925,N_1834);
or U2688 (N_2688,N_1696,N_1146);
or U2689 (N_2689,N_1163,N_1195);
and U2690 (N_2690,N_1566,N_1595);
nand U2691 (N_2691,N_1353,N_1873);
nand U2692 (N_2692,N_1555,N_1768);
xnor U2693 (N_2693,N_1833,N_1086);
and U2694 (N_2694,N_1530,N_1145);
nand U2695 (N_2695,N_1837,N_1456);
and U2696 (N_2696,N_1063,N_1227);
nor U2697 (N_2697,N_1794,N_1358);
nor U2698 (N_2698,N_1256,N_1823);
xnor U2699 (N_2699,N_1915,N_1063);
nand U2700 (N_2700,N_1504,N_1102);
nand U2701 (N_2701,N_1485,N_1200);
or U2702 (N_2702,N_1574,N_1634);
nor U2703 (N_2703,N_1558,N_1547);
or U2704 (N_2704,N_1704,N_1505);
nor U2705 (N_2705,N_1304,N_1188);
or U2706 (N_2706,N_1760,N_1340);
and U2707 (N_2707,N_1520,N_1356);
nand U2708 (N_2708,N_1722,N_1242);
nor U2709 (N_2709,N_1921,N_1901);
and U2710 (N_2710,N_1077,N_1213);
xor U2711 (N_2711,N_1595,N_1253);
or U2712 (N_2712,N_1519,N_1903);
nand U2713 (N_2713,N_1306,N_1407);
or U2714 (N_2714,N_1416,N_1510);
or U2715 (N_2715,N_1379,N_1947);
xnor U2716 (N_2716,N_1671,N_1787);
xnor U2717 (N_2717,N_1137,N_1398);
or U2718 (N_2718,N_1538,N_1342);
xor U2719 (N_2719,N_1924,N_1681);
and U2720 (N_2720,N_1054,N_1694);
or U2721 (N_2721,N_1525,N_1511);
and U2722 (N_2722,N_1666,N_1178);
nor U2723 (N_2723,N_1875,N_1783);
and U2724 (N_2724,N_1278,N_1051);
nand U2725 (N_2725,N_1462,N_1980);
or U2726 (N_2726,N_1571,N_1377);
or U2727 (N_2727,N_1695,N_1112);
nand U2728 (N_2728,N_1248,N_1812);
xnor U2729 (N_2729,N_1867,N_1554);
nor U2730 (N_2730,N_1278,N_1965);
and U2731 (N_2731,N_1182,N_1525);
nor U2732 (N_2732,N_1978,N_1669);
nor U2733 (N_2733,N_1289,N_1727);
nand U2734 (N_2734,N_1711,N_1539);
or U2735 (N_2735,N_1530,N_1265);
xnor U2736 (N_2736,N_1020,N_1465);
nor U2737 (N_2737,N_1040,N_1332);
and U2738 (N_2738,N_1231,N_1820);
and U2739 (N_2739,N_1654,N_1794);
and U2740 (N_2740,N_1105,N_1223);
and U2741 (N_2741,N_1436,N_1348);
or U2742 (N_2742,N_1759,N_1825);
xnor U2743 (N_2743,N_1776,N_1111);
or U2744 (N_2744,N_1963,N_1005);
nor U2745 (N_2745,N_1738,N_1759);
xor U2746 (N_2746,N_1998,N_1892);
and U2747 (N_2747,N_1298,N_1017);
nand U2748 (N_2748,N_1668,N_1275);
or U2749 (N_2749,N_1376,N_1766);
and U2750 (N_2750,N_1440,N_1705);
nand U2751 (N_2751,N_1529,N_1453);
or U2752 (N_2752,N_1076,N_1320);
or U2753 (N_2753,N_1468,N_1598);
xor U2754 (N_2754,N_1276,N_1034);
xor U2755 (N_2755,N_1126,N_1336);
xnor U2756 (N_2756,N_1806,N_1258);
or U2757 (N_2757,N_1450,N_1046);
or U2758 (N_2758,N_1756,N_1577);
xnor U2759 (N_2759,N_1224,N_1988);
or U2760 (N_2760,N_1797,N_1855);
or U2761 (N_2761,N_1837,N_1201);
xor U2762 (N_2762,N_1660,N_1400);
or U2763 (N_2763,N_1058,N_1694);
xor U2764 (N_2764,N_1434,N_1613);
xor U2765 (N_2765,N_1234,N_1649);
nand U2766 (N_2766,N_1759,N_1337);
nor U2767 (N_2767,N_1358,N_1738);
xor U2768 (N_2768,N_1939,N_1179);
xnor U2769 (N_2769,N_1337,N_1160);
nand U2770 (N_2770,N_1727,N_1920);
nand U2771 (N_2771,N_1383,N_1272);
xor U2772 (N_2772,N_1335,N_1631);
and U2773 (N_2773,N_1975,N_1538);
nand U2774 (N_2774,N_1971,N_1939);
xor U2775 (N_2775,N_1662,N_1002);
and U2776 (N_2776,N_1182,N_1447);
or U2777 (N_2777,N_1202,N_1190);
nand U2778 (N_2778,N_1078,N_1278);
and U2779 (N_2779,N_1581,N_1451);
xnor U2780 (N_2780,N_1267,N_1230);
and U2781 (N_2781,N_1480,N_1472);
nor U2782 (N_2782,N_1520,N_1227);
nor U2783 (N_2783,N_1411,N_1337);
or U2784 (N_2784,N_1767,N_1115);
xor U2785 (N_2785,N_1555,N_1144);
nor U2786 (N_2786,N_1669,N_1878);
or U2787 (N_2787,N_1531,N_1779);
xnor U2788 (N_2788,N_1098,N_1086);
and U2789 (N_2789,N_1749,N_1921);
or U2790 (N_2790,N_1676,N_1294);
or U2791 (N_2791,N_1265,N_1969);
nor U2792 (N_2792,N_1229,N_1244);
nand U2793 (N_2793,N_1108,N_1242);
or U2794 (N_2794,N_1250,N_1867);
nand U2795 (N_2795,N_1896,N_1218);
nor U2796 (N_2796,N_1267,N_1618);
xnor U2797 (N_2797,N_1838,N_1321);
xor U2798 (N_2798,N_1075,N_1520);
or U2799 (N_2799,N_1994,N_1246);
nor U2800 (N_2800,N_1016,N_1165);
xnor U2801 (N_2801,N_1795,N_1524);
nand U2802 (N_2802,N_1795,N_1813);
xor U2803 (N_2803,N_1161,N_1473);
xor U2804 (N_2804,N_1628,N_1744);
or U2805 (N_2805,N_1232,N_1636);
or U2806 (N_2806,N_1597,N_1495);
or U2807 (N_2807,N_1947,N_1201);
nand U2808 (N_2808,N_1435,N_1052);
nor U2809 (N_2809,N_1830,N_1266);
xor U2810 (N_2810,N_1715,N_1919);
nor U2811 (N_2811,N_1717,N_1249);
xor U2812 (N_2812,N_1026,N_1004);
or U2813 (N_2813,N_1780,N_1088);
nand U2814 (N_2814,N_1465,N_1304);
xor U2815 (N_2815,N_1218,N_1698);
and U2816 (N_2816,N_1674,N_1824);
and U2817 (N_2817,N_1083,N_1901);
xnor U2818 (N_2818,N_1482,N_1008);
xor U2819 (N_2819,N_1299,N_1865);
nand U2820 (N_2820,N_1105,N_1622);
nor U2821 (N_2821,N_1185,N_1347);
nand U2822 (N_2822,N_1245,N_1026);
xnor U2823 (N_2823,N_1566,N_1785);
and U2824 (N_2824,N_1043,N_1008);
and U2825 (N_2825,N_1242,N_1353);
and U2826 (N_2826,N_1941,N_1658);
xor U2827 (N_2827,N_1380,N_1787);
and U2828 (N_2828,N_1300,N_1368);
nand U2829 (N_2829,N_1346,N_1646);
xnor U2830 (N_2830,N_1477,N_1073);
nand U2831 (N_2831,N_1810,N_1338);
xnor U2832 (N_2832,N_1477,N_1710);
and U2833 (N_2833,N_1866,N_1700);
or U2834 (N_2834,N_1022,N_1401);
and U2835 (N_2835,N_1460,N_1098);
or U2836 (N_2836,N_1208,N_1619);
or U2837 (N_2837,N_1366,N_1002);
and U2838 (N_2838,N_1829,N_1926);
and U2839 (N_2839,N_1938,N_1744);
nor U2840 (N_2840,N_1854,N_1349);
xor U2841 (N_2841,N_1836,N_1169);
or U2842 (N_2842,N_1896,N_1009);
xor U2843 (N_2843,N_1428,N_1041);
or U2844 (N_2844,N_1376,N_1418);
or U2845 (N_2845,N_1459,N_1344);
nor U2846 (N_2846,N_1611,N_1172);
xor U2847 (N_2847,N_1609,N_1850);
nand U2848 (N_2848,N_1531,N_1798);
nor U2849 (N_2849,N_1617,N_1992);
or U2850 (N_2850,N_1015,N_1917);
or U2851 (N_2851,N_1555,N_1191);
nand U2852 (N_2852,N_1228,N_1014);
xnor U2853 (N_2853,N_1958,N_1135);
nand U2854 (N_2854,N_1215,N_1501);
xnor U2855 (N_2855,N_1836,N_1496);
nand U2856 (N_2856,N_1879,N_1928);
and U2857 (N_2857,N_1491,N_1281);
and U2858 (N_2858,N_1976,N_1318);
xor U2859 (N_2859,N_1555,N_1336);
xnor U2860 (N_2860,N_1336,N_1050);
and U2861 (N_2861,N_1073,N_1506);
xor U2862 (N_2862,N_1596,N_1538);
or U2863 (N_2863,N_1298,N_1755);
xor U2864 (N_2864,N_1807,N_1185);
or U2865 (N_2865,N_1708,N_1717);
nand U2866 (N_2866,N_1595,N_1874);
nor U2867 (N_2867,N_1392,N_1945);
or U2868 (N_2868,N_1899,N_1283);
nor U2869 (N_2869,N_1899,N_1711);
and U2870 (N_2870,N_1694,N_1241);
xor U2871 (N_2871,N_1881,N_1572);
nor U2872 (N_2872,N_1272,N_1406);
or U2873 (N_2873,N_1967,N_1853);
nand U2874 (N_2874,N_1409,N_1756);
xor U2875 (N_2875,N_1283,N_1231);
or U2876 (N_2876,N_1098,N_1838);
and U2877 (N_2877,N_1975,N_1772);
xor U2878 (N_2878,N_1487,N_1166);
and U2879 (N_2879,N_1147,N_1697);
nand U2880 (N_2880,N_1614,N_1317);
xor U2881 (N_2881,N_1619,N_1986);
nor U2882 (N_2882,N_1223,N_1981);
nor U2883 (N_2883,N_1552,N_1894);
xor U2884 (N_2884,N_1171,N_1964);
nor U2885 (N_2885,N_1437,N_1324);
and U2886 (N_2886,N_1734,N_1356);
and U2887 (N_2887,N_1651,N_1826);
and U2888 (N_2888,N_1619,N_1552);
or U2889 (N_2889,N_1783,N_1898);
nand U2890 (N_2890,N_1983,N_1949);
nand U2891 (N_2891,N_1263,N_1644);
or U2892 (N_2892,N_1808,N_1200);
and U2893 (N_2893,N_1206,N_1856);
and U2894 (N_2894,N_1198,N_1338);
and U2895 (N_2895,N_1910,N_1550);
nand U2896 (N_2896,N_1239,N_1982);
nor U2897 (N_2897,N_1470,N_1957);
xnor U2898 (N_2898,N_1765,N_1898);
xor U2899 (N_2899,N_1885,N_1799);
xor U2900 (N_2900,N_1691,N_1224);
nor U2901 (N_2901,N_1124,N_1640);
or U2902 (N_2902,N_1888,N_1743);
and U2903 (N_2903,N_1685,N_1731);
or U2904 (N_2904,N_1363,N_1128);
nor U2905 (N_2905,N_1452,N_1004);
nand U2906 (N_2906,N_1262,N_1444);
or U2907 (N_2907,N_1856,N_1903);
and U2908 (N_2908,N_1253,N_1875);
and U2909 (N_2909,N_1989,N_1593);
xor U2910 (N_2910,N_1930,N_1702);
xor U2911 (N_2911,N_1530,N_1567);
or U2912 (N_2912,N_1155,N_1331);
xnor U2913 (N_2913,N_1303,N_1380);
nor U2914 (N_2914,N_1646,N_1616);
xor U2915 (N_2915,N_1592,N_1368);
and U2916 (N_2916,N_1660,N_1168);
or U2917 (N_2917,N_1957,N_1526);
nor U2918 (N_2918,N_1157,N_1652);
nor U2919 (N_2919,N_1743,N_1496);
nor U2920 (N_2920,N_1377,N_1213);
nand U2921 (N_2921,N_1023,N_1707);
nor U2922 (N_2922,N_1811,N_1602);
nor U2923 (N_2923,N_1672,N_1505);
or U2924 (N_2924,N_1047,N_1407);
nor U2925 (N_2925,N_1455,N_1255);
xnor U2926 (N_2926,N_1375,N_1060);
or U2927 (N_2927,N_1948,N_1934);
nand U2928 (N_2928,N_1408,N_1272);
or U2929 (N_2929,N_1807,N_1413);
nor U2930 (N_2930,N_1327,N_1175);
nand U2931 (N_2931,N_1978,N_1976);
nand U2932 (N_2932,N_1104,N_1903);
and U2933 (N_2933,N_1513,N_1080);
or U2934 (N_2934,N_1605,N_1398);
and U2935 (N_2935,N_1788,N_1861);
xnor U2936 (N_2936,N_1104,N_1234);
nand U2937 (N_2937,N_1438,N_1820);
and U2938 (N_2938,N_1534,N_1440);
or U2939 (N_2939,N_1430,N_1761);
nor U2940 (N_2940,N_1547,N_1681);
nor U2941 (N_2941,N_1658,N_1805);
or U2942 (N_2942,N_1116,N_1041);
xnor U2943 (N_2943,N_1726,N_1167);
or U2944 (N_2944,N_1968,N_1857);
xor U2945 (N_2945,N_1725,N_1611);
nor U2946 (N_2946,N_1989,N_1105);
nor U2947 (N_2947,N_1415,N_1258);
xnor U2948 (N_2948,N_1241,N_1437);
xor U2949 (N_2949,N_1040,N_1561);
xnor U2950 (N_2950,N_1136,N_1239);
nand U2951 (N_2951,N_1288,N_1287);
xnor U2952 (N_2952,N_1894,N_1209);
and U2953 (N_2953,N_1157,N_1544);
xnor U2954 (N_2954,N_1385,N_1399);
nand U2955 (N_2955,N_1005,N_1591);
nor U2956 (N_2956,N_1119,N_1658);
nor U2957 (N_2957,N_1106,N_1173);
nand U2958 (N_2958,N_1501,N_1323);
and U2959 (N_2959,N_1888,N_1349);
nor U2960 (N_2960,N_1596,N_1543);
xnor U2961 (N_2961,N_1598,N_1216);
nor U2962 (N_2962,N_1112,N_1278);
and U2963 (N_2963,N_1221,N_1053);
nor U2964 (N_2964,N_1720,N_1531);
xor U2965 (N_2965,N_1429,N_1939);
nor U2966 (N_2966,N_1970,N_1767);
xnor U2967 (N_2967,N_1763,N_1225);
and U2968 (N_2968,N_1105,N_1022);
and U2969 (N_2969,N_1548,N_1239);
or U2970 (N_2970,N_1715,N_1300);
nor U2971 (N_2971,N_1918,N_1924);
or U2972 (N_2972,N_1596,N_1287);
or U2973 (N_2973,N_1347,N_1186);
nor U2974 (N_2974,N_1060,N_1350);
nor U2975 (N_2975,N_1369,N_1836);
nand U2976 (N_2976,N_1807,N_1629);
xnor U2977 (N_2977,N_1635,N_1915);
and U2978 (N_2978,N_1086,N_1535);
nor U2979 (N_2979,N_1947,N_1176);
or U2980 (N_2980,N_1645,N_1468);
and U2981 (N_2981,N_1456,N_1216);
nand U2982 (N_2982,N_1112,N_1712);
nor U2983 (N_2983,N_1236,N_1408);
or U2984 (N_2984,N_1228,N_1423);
and U2985 (N_2985,N_1785,N_1201);
nor U2986 (N_2986,N_1819,N_1593);
xnor U2987 (N_2987,N_1791,N_1677);
nor U2988 (N_2988,N_1961,N_1031);
xnor U2989 (N_2989,N_1428,N_1967);
or U2990 (N_2990,N_1519,N_1039);
or U2991 (N_2991,N_1119,N_1255);
nor U2992 (N_2992,N_1499,N_1996);
and U2993 (N_2993,N_1062,N_1599);
xnor U2994 (N_2994,N_1492,N_1567);
and U2995 (N_2995,N_1510,N_1009);
nor U2996 (N_2996,N_1298,N_1078);
nand U2997 (N_2997,N_1065,N_1133);
nor U2998 (N_2998,N_1059,N_1371);
xor U2999 (N_2999,N_1265,N_1192);
and U3000 (N_3000,N_2012,N_2632);
nor U3001 (N_3001,N_2551,N_2016);
or U3002 (N_3002,N_2333,N_2426);
nor U3003 (N_3003,N_2484,N_2665);
nor U3004 (N_3004,N_2335,N_2981);
xnor U3005 (N_3005,N_2988,N_2510);
and U3006 (N_3006,N_2447,N_2460);
nor U3007 (N_3007,N_2262,N_2050);
and U3008 (N_3008,N_2161,N_2987);
or U3009 (N_3009,N_2656,N_2435);
nor U3010 (N_3010,N_2037,N_2906);
and U3011 (N_3011,N_2862,N_2537);
xnor U3012 (N_3012,N_2894,N_2831);
nor U3013 (N_3013,N_2993,N_2115);
nor U3014 (N_3014,N_2601,N_2373);
nor U3015 (N_3015,N_2807,N_2804);
and U3016 (N_3016,N_2374,N_2899);
nor U3017 (N_3017,N_2554,N_2960);
nor U3018 (N_3018,N_2366,N_2179);
nand U3019 (N_3019,N_2590,N_2642);
xor U3020 (N_3020,N_2901,N_2133);
nor U3021 (N_3021,N_2956,N_2591);
nand U3022 (N_3022,N_2483,N_2748);
nand U3023 (N_3023,N_2886,N_2569);
and U3024 (N_3024,N_2626,N_2630);
nor U3025 (N_3025,N_2280,N_2573);
nand U3026 (N_3026,N_2035,N_2026);
xor U3027 (N_3027,N_2602,N_2568);
nand U3028 (N_3028,N_2726,N_2215);
nand U3029 (N_3029,N_2407,N_2301);
nor U3030 (N_3030,N_2768,N_2648);
or U3031 (N_3031,N_2033,N_2452);
nor U3032 (N_3032,N_2889,N_2455);
nor U3033 (N_3033,N_2297,N_2518);
nor U3034 (N_3034,N_2259,N_2021);
xnor U3035 (N_3035,N_2307,N_2806);
nor U3036 (N_3036,N_2123,N_2370);
nor U3037 (N_3037,N_2681,N_2896);
or U3038 (N_3038,N_2608,N_2060);
or U3039 (N_3039,N_2675,N_2337);
or U3040 (N_3040,N_2405,N_2725);
nor U3041 (N_3041,N_2286,N_2598);
nor U3042 (N_3042,N_2178,N_2345);
or U3043 (N_3043,N_2089,N_2378);
or U3044 (N_3044,N_2176,N_2130);
and U3045 (N_3045,N_2078,N_2134);
or U3046 (N_3046,N_2913,N_2409);
xnor U3047 (N_3047,N_2903,N_2272);
xor U3048 (N_3048,N_2430,N_2266);
xor U3049 (N_3049,N_2369,N_2087);
and U3050 (N_3050,N_2132,N_2287);
nand U3051 (N_3051,N_2208,N_2462);
xnor U3052 (N_3052,N_2047,N_2876);
and U3053 (N_3053,N_2940,N_2222);
nand U3054 (N_3054,N_2186,N_2833);
and U3055 (N_3055,N_2404,N_2531);
nand U3056 (N_3056,N_2613,N_2214);
nand U3057 (N_3057,N_2304,N_2446);
nor U3058 (N_3058,N_2635,N_2224);
or U3059 (N_3059,N_2359,N_2715);
or U3060 (N_3060,N_2197,N_2588);
nor U3061 (N_3061,N_2223,N_2902);
or U3062 (N_3062,N_2283,N_2892);
and U3063 (N_3063,N_2282,N_2014);
or U3064 (N_3064,N_2159,N_2812);
xnor U3065 (N_3065,N_2997,N_2767);
and U3066 (N_3066,N_2924,N_2458);
nor U3067 (N_3067,N_2647,N_2425);
nand U3068 (N_3068,N_2382,N_2189);
xnor U3069 (N_3069,N_2934,N_2929);
nand U3070 (N_3070,N_2488,N_2414);
xor U3071 (N_3071,N_2926,N_2007);
or U3072 (N_3072,N_2508,N_2713);
nor U3073 (N_3073,N_2128,N_2163);
nand U3074 (N_3074,N_2211,N_2803);
or U3075 (N_3075,N_2391,N_2062);
nand U3076 (N_3076,N_2983,N_2503);
nor U3077 (N_3077,N_2645,N_2332);
nor U3078 (N_3078,N_2057,N_2631);
xor U3079 (N_3079,N_2195,N_2381);
or U3080 (N_3080,N_2069,N_2641);
and U3081 (N_3081,N_2238,N_2463);
and U3082 (N_3082,N_2160,N_2908);
nand U3083 (N_3083,N_2196,N_2257);
or U3084 (N_3084,N_2083,N_2486);
nand U3085 (N_3085,N_2158,N_2830);
and U3086 (N_3086,N_2619,N_2148);
nand U3087 (N_3087,N_2730,N_2759);
or U3088 (N_3088,N_2838,N_2239);
xor U3089 (N_3089,N_2342,N_2922);
and U3090 (N_3090,N_2042,N_2618);
and U3091 (N_3091,N_2753,N_2376);
xor U3092 (N_3092,N_2535,N_2315);
and U3093 (N_3093,N_2693,N_2808);
or U3094 (N_3094,N_2689,N_2579);
and U3095 (N_3095,N_2324,N_2822);
and U3096 (N_3096,N_2346,N_2939);
or U3097 (N_3097,N_2390,N_2683);
and U3098 (N_3098,N_2809,N_2989);
xor U3099 (N_3099,N_2005,N_2487);
nor U3100 (N_3100,N_2118,N_2221);
nor U3101 (N_3101,N_2853,N_2536);
or U3102 (N_3102,N_2859,N_2774);
xor U3103 (N_3103,N_2786,N_2230);
or U3104 (N_3104,N_2204,N_2646);
nor U3105 (N_3105,N_2799,N_2321);
xnor U3106 (N_3106,N_2676,N_2972);
nand U3107 (N_3107,N_2720,N_2900);
or U3108 (N_3108,N_2281,N_2246);
nand U3109 (N_3109,N_2098,N_2517);
nand U3110 (N_3110,N_2511,N_2268);
xor U3111 (N_3111,N_2564,N_2560);
xor U3112 (N_3112,N_2493,N_2516);
nor U3113 (N_3113,N_2302,N_2909);
and U3114 (N_3114,N_2476,N_2723);
or U3115 (N_3115,N_2441,N_2780);
or U3116 (N_3116,N_2056,N_2393);
nor U3117 (N_3117,N_2076,N_2457);
nor U3118 (N_3118,N_2314,N_2668);
nand U3119 (N_3119,N_2000,N_2636);
nor U3120 (N_3120,N_2003,N_2750);
or U3121 (N_3121,N_2840,N_2361);
and U3122 (N_3122,N_2942,N_2670);
nor U3123 (N_3123,N_2684,N_2616);
nand U3124 (N_3124,N_2053,N_2582);
nand U3125 (N_3125,N_2193,N_2072);
xor U3126 (N_3126,N_2495,N_2071);
nand U3127 (N_3127,N_2024,N_2592);
nand U3128 (N_3128,N_2261,N_2881);
and U3129 (N_3129,N_2991,N_2164);
or U3130 (N_3130,N_2787,N_2653);
or U3131 (N_3131,N_2250,N_2932);
nand U3132 (N_3132,N_2818,N_2490);
nor U3133 (N_3133,N_2949,N_2334);
nand U3134 (N_3134,N_2336,N_2459);
or U3135 (N_3135,N_2755,N_2930);
xor U3136 (N_3136,N_2309,N_2776);
or U3137 (N_3137,N_2891,N_2984);
nor U3138 (N_3138,N_2088,N_2864);
xnor U3139 (N_3139,N_2200,N_2696);
nand U3140 (N_3140,N_2865,N_2621);
or U3141 (N_3141,N_2437,N_2316);
nand U3142 (N_3142,N_2008,N_2168);
and U3143 (N_3143,N_2883,N_2121);
nor U3144 (N_3144,N_2890,N_2971);
nor U3145 (N_3145,N_2920,N_2917);
and U3146 (N_3146,N_2363,N_2585);
nand U3147 (N_3147,N_2880,N_2350);
xnor U3148 (N_3148,N_2773,N_2438);
or U3149 (N_3149,N_2948,N_2058);
or U3150 (N_3150,N_2769,N_2842);
nand U3151 (N_3151,N_2663,N_2036);
or U3152 (N_3152,N_2629,N_2639);
nor U3153 (N_3153,N_2565,N_2527);
nor U3154 (N_3154,N_2063,N_2563);
nand U3155 (N_3155,N_2789,N_2294);
nor U3156 (N_3156,N_2392,N_2116);
or U3157 (N_3157,N_2513,N_2594);
and U3158 (N_3158,N_2279,N_2443);
nand U3159 (N_3159,N_2338,N_2794);
nand U3160 (N_3160,N_2092,N_2403);
and U3161 (N_3161,N_2276,N_2615);
and U3162 (N_3162,N_2420,N_2846);
and U3163 (N_3163,N_2649,N_2580);
nand U3164 (N_3164,N_2628,N_2874);
or U3165 (N_3165,N_2212,N_2802);
or U3166 (N_3166,N_2686,N_2144);
nor U3167 (N_3167,N_2135,N_2706);
or U3168 (N_3168,N_2567,N_2935);
xnor U3169 (N_3169,N_2104,N_2474);
and U3170 (N_3170,N_2986,N_2109);
nor U3171 (N_3171,N_2293,N_2006);
xnor U3172 (N_3172,N_2423,N_2589);
xor U3173 (N_3173,N_2586,N_2740);
nand U3174 (N_3174,N_2228,N_2959);
and U3175 (N_3175,N_2220,N_2577);
nand U3176 (N_3176,N_2429,N_2442);
nor U3177 (N_3177,N_2235,N_2171);
xnor U3178 (N_3178,N_2013,N_2532);
nand U3179 (N_3179,N_2107,N_2165);
or U3180 (N_3180,N_2152,N_2082);
nor U3181 (N_3181,N_2703,N_2075);
or U3182 (N_3182,N_2002,N_2795);
nand U3183 (N_3183,N_2539,N_2722);
and U3184 (N_3184,N_2739,N_2623);
and U3185 (N_3185,N_2763,N_2432);
xnor U3186 (N_3186,N_2300,N_2733);
nor U3187 (N_3187,N_2182,N_2103);
nor U3188 (N_3188,N_2039,N_2188);
nand U3189 (N_3189,N_2364,N_2718);
or U3190 (N_3190,N_2719,N_2356);
xnor U3191 (N_3191,N_2509,N_2553);
nand U3192 (N_3192,N_2085,N_2368);
nor U3193 (N_3193,N_2701,N_2111);
or U3194 (N_3194,N_2436,N_2660);
and U3195 (N_3195,N_2977,N_2108);
nand U3196 (N_3196,N_2990,N_2669);
or U3197 (N_3197,N_2955,N_2873);
and U3198 (N_3198,N_2832,N_2512);
nand U3199 (N_3199,N_2856,N_2622);
or U3200 (N_3200,N_2729,N_2244);
nand U3201 (N_3201,N_2765,N_2049);
xor U3202 (N_3202,N_2064,N_2785);
nor U3203 (N_3203,N_2844,N_2124);
and U3204 (N_3204,N_2120,N_2581);
or U3205 (N_3205,N_2354,N_2270);
and U3206 (N_3206,N_2925,N_2845);
nor U3207 (N_3207,N_2783,N_2424);
nand U3208 (N_3208,N_2870,N_2600);
nor U3209 (N_3209,N_2728,N_2610);
or U3210 (N_3210,N_2732,N_2814);
nand U3211 (N_3211,N_2471,N_2248);
and U3212 (N_3212,N_2945,N_2073);
and U3213 (N_3213,N_2331,N_2284);
nand U3214 (N_3214,N_2708,N_2947);
xnor U3215 (N_3215,N_2702,N_2371);
xor U3216 (N_3216,N_2792,N_2500);
nor U3217 (N_3217,N_2866,N_2253);
and U3218 (N_3218,N_2348,N_2637);
xor U3219 (N_3219,N_2810,N_2030);
nand U3220 (N_3220,N_2289,N_2587);
nand U3221 (N_3221,N_2805,N_2678);
nand U3222 (N_3222,N_2944,N_2597);
or U3223 (N_3223,N_2943,N_2170);
and U3224 (N_3224,N_2052,N_2218);
xor U3225 (N_3225,N_2032,N_2101);
nor U3226 (N_3226,N_2156,N_2823);
xor U3227 (N_3227,N_2687,N_2698);
nand U3228 (N_3228,N_2966,N_2153);
xnor U3229 (N_3229,N_2341,N_2147);
nand U3230 (N_3230,N_2764,N_2410);
or U3231 (N_3231,N_2923,N_2643);
or U3232 (N_3232,N_2957,N_2682);
nand U3233 (N_3233,N_2916,N_2854);
and U3234 (N_3234,N_2136,N_2735);
or U3235 (N_3235,N_2504,N_2275);
nand U3236 (N_3236,N_2982,N_2263);
nor U3237 (N_3237,N_2761,N_2879);
or U3238 (N_3238,N_2154,N_2209);
nand U3239 (N_3239,N_2482,N_2980);
and U3240 (N_3240,N_2754,N_2146);
and U3241 (N_3241,N_2782,N_2044);
nor U3242 (N_3242,N_2352,N_2548);
xnor U3243 (N_3243,N_2545,N_2968);
and U3244 (N_3244,N_2019,N_2213);
and U3245 (N_3245,N_2367,N_2444);
nand U3246 (N_3246,N_2097,N_2634);
nor U3247 (N_3247,N_2157,N_2743);
or U3248 (N_3248,N_2129,N_2882);
or U3249 (N_3249,N_2766,N_2712);
or U3250 (N_3250,N_2938,N_2907);
nor U3251 (N_3251,N_2954,N_2562);
or U3252 (N_3252,N_2847,N_2408);
nand U3253 (N_3253,N_2251,N_2481);
nor U3254 (N_3254,N_2661,N_2714);
and U3255 (N_3255,N_2625,N_2593);
nor U3256 (N_3256,N_2737,N_2093);
xnor U3257 (N_3257,N_2970,N_2671);
or U3258 (N_3258,N_2100,N_2861);
nand U3259 (N_3259,N_2835,N_2542);
nand U3260 (N_3260,N_2697,N_2177);
or U3261 (N_3261,N_2330,N_2612);
xor U3262 (N_3262,N_2233,N_2340);
and U3263 (N_3263,N_2633,N_2265);
xor U3264 (N_3264,N_2666,N_2237);
nand U3265 (N_3265,N_2815,N_2617);
nor U3266 (N_3266,N_2421,N_2415);
or U3267 (N_3267,N_2974,N_2979);
nor U3268 (N_3268,N_2243,N_2258);
nand U3269 (N_3269,N_2523,N_2095);
or U3270 (N_3270,N_2716,N_2198);
nand U3271 (N_3271,N_2519,N_2395);
or U3272 (N_3272,N_2695,N_2662);
and U3273 (N_3273,N_2738,N_2839);
nor U3274 (N_3274,N_2933,N_2758);
nor U3275 (N_3275,N_2910,N_2175);
or U3276 (N_3276,N_2040,N_2679);
nor U3277 (N_3277,N_2820,N_2267);
nand U3278 (N_3278,N_2143,N_2505);
nor U3279 (N_3279,N_2538,N_2492);
nand U3280 (N_3280,N_2126,N_2973);
or U3281 (N_3281,N_2180,N_2264);
or U3282 (N_3282,N_2606,N_2269);
nand U3283 (N_3283,N_2285,N_2745);
and U3284 (N_3284,N_2796,N_2520);
and U3285 (N_3285,N_2451,N_2790);
and U3286 (N_3286,N_2863,N_2868);
and U3287 (N_3287,N_2306,N_2322);
or U3288 (N_3288,N_2028,N_2313);
xor U3289 (N_3289,N_2234,N_2166);
and U3290 (N_3290,N_2417,N_2034);
nand U3291 (N_3291,N_2245,N_2385);
and U3292 (N_3292,N_2499,N_2657);
or U3293 (N_3293,N_2507,N_2137);
nand U3294 (N_3294,N_2751,N_2066);
nand U3295 (N_3295,N_2172,N_2952);
xor U3296 (N_3296,N_2375,N_2206);
or U3297 (N_3297,N_2688,N_2312);
and U3298 (N_3298,N_2848,N_2122);
or U3299 (N_3299,N_2640,N_2318);
or U3300 (N_3300,N_2529,N_2710);
and U3301 (N_3301,N_2534,N_2936);
xnor U3302 (N_3302,N_2771,N_2961);
and U3303 (N_3303,N_2941,N_2843);
nand U3304 (N_3304,N_2043,N_2018);
or U3305 (N_3305,N_2816,N_2400);
nor U3306 (N_3306,N_2690,N_2469);
nand U3307 (N_3307,N_2788,N_2046);
and U3308 (N_3308,N_2658,N_2439);
nand U3309 (N_3309,N_2192,N_2887);
or U3310 (N_3310,N_2311,N_2976);
nor U3311 (N_3311,N_2699,N_2885);
and U3312 (N_3312,N_2090,N_2320);
nand U3313 (N_3313,N_2819,N_2543);
or U3314 (N_3314,N_2022,N_2607);
nor U3315 (N_3315,N_2328,N_2584);
xor U3316 (N_3316,N_2422,N_2365);
nand U3317 (N_3317,N_2652,N_2999);
xnor U3318 (N_3318,N_2978,N_2967);
and U3319 (N_3319,N_2489,N_2599);
nor U3320 (N_3320,N_2431,N_2604);
xnor U3321 (N_3321,N_2996,N_2691);
nand U3322 (N_3322,N_2260,N_2609);
and U3323 (N_3323,N_2644,N_2216);
nand U3324 (N_3324,N_2247,N_2305);
nand U3325 (N_3325,N_2308,N_2397);
and U3326 (N_3326,N_2841,N_2528);
nor U3327 (N_3327,N_2897,N_2461);
and U3328 (N_3328,N_2398,N_2914);
nor U3329 (N_3329,N_2453,N_2203);
nand U3330 (N_3330,N_2477,N_2800);
nor U3331 (N_3331,N_2888,N_2875);
xnor U3332 (N_3332,N_2672,N_2491);
xnor U3333 (N_3333,N_2544,N_2756);
nand U3334 (N_3334,N_2068,N_2388);
or U3335 (N_3335,N_2394,N_2110);
xnor U3336 (N_3336,N_2498,N_2497);
xnor U3337 (N_3337,N_2406,N_2242);
nor U3338 (N_3338,N_2749,N_2834);
or U3339 (N_3339,N_2347,N_2227);
xor U3340 (N_3340,N_2319,N_2550);
or U3341 (N_3341,N_2918,N_2667);
nand U3342 (N_3342,N_2201,N_2349);
and U3343 (N_3343,N_2558,N_2310);
and U3344 (N_3344,N_2045,N_2029);
and U3345 (N_3345,N_2950,N_2546);
or U3346 (N_3346,N_2290,N_2860);
or U3347 (N_3347,N_2358,N_2775);
or U3348 (N_3348,N_2638,N_2557);
xor U3349 (N_3349,N_2141,N_2241);
nor U3350 (N_3350,N_2798,N_2526);
xor U3351 (N_3351,N_2867,N_2249);
or U3352 (N_3352,N_2998,N_2521);
nor U3353 (N_3353,N_2449,N_2884);
nand U3354 (N_3354,N_2271,N_2065);
nand U3355 (N_3355,N_2454,N_2533);
and U3356 (N_3356,N_2360,N_2086);
xnor U3357 (N_3357,N_2797,N_2556);
nand U3358 (N_3358,N_2210,N_2339);
xnor U3359 (N_3359,N_2694,N_2829);
xnor U3360 (N_3360,N_2292,N_2741);
xor U3361 (N_3361,N_2871,N_2813);
xor U3362 (N_3362,N_2522,N_2202);
nand U3363 (N_3363,N_2023,N_2480);
nand U3364 (N_3364,N_2872,N_2850);
xor U3365 (N_3365,N_2450,N_2205);
xnor U3366 (N_3366,N_2377,N_2836);
nor U3367 (N_3367,N_2174,N_2372);
nor U3368 (N_3368,N_2605,N_2434);
or U3369 (N_3369,N_2811,N_2650);
xnor U3370 (N_3370,N_2139,N_2054);
nand U3371 (N_3371,N_2965,N_2418);
xnor U3372 (N_3372,N_2027,N_2946);
and U3373 (N_3373,N_2145,N_2199);
nand U3374 (N_3374,N_2274,N_2416);
nor U3375 (N_3375,N_2760,N_2167);
and U3376 (N_3376,N_2419,N_2825);
xor U3377 (N_3377,N_2389,N_2399);
or U3378 (N_3378,N_2921,N_2898);
nor U3379 (N_3379,N_2155,N_2817);
nand U3380 (N_3380,N_2576,N_2826);
xor U3381 (N_3381,N_2692,N_2963);
and U3382 (N_3382,N_2067,N_2962);
xor U3383 (N_3383,N_2411,N_2525);
xor U3384 (N_3384,N_2578,N_2895);
and U3385 (N_3385,N_2468,N_2911);
nor U3386 (N_3386,N_2747,N_2327);
xor U3387 (N_3387,N_2080,N_2985);
nor U3388 (N_3388,N_2734,N_2849);
or U3389 (N_3389,N_2478,N_2169);
and U3390 (N_3390,N_2225,N_2323);
and U3391 (N_3391,N_2709,N_2232);
xor U3392 (N_3392,N_2413,N_2278);
and U3393 (N_3393,N_2010,N_2524);
or U3394 (N_3394,N_2295,N_2851);
nor U3395 (N_3395,N_2975,N_2995);
nor U3396 (N_3396,N_2048,N_2721);
nor U3397 (N_3397,N_2705,N_2094);
and U3398 (N_3398,N_2401,N_2680);
nor U3399 (N_3399,N_2717,N_2791);
or U3400 (N_3400,N_2762,N_2298);
and U3401 (N_3401,N_2217,N_2994);
nor U3402 (N_3402,N_2912,N_2479);
nand U3403 (N_3403,N_2904,N_2362);
or U3404 (N_3404,N_2291,N_2931);
or U3405 (N_3405,N_2020,N_2254);
or U3406 (N_3406,N_2757,N_2927);
and U3407 (N_3407,N_2387,N_2878);
or U3408 (N_3408,N_2541,N_2114);
nor U3409 (N_3409,N_2119,N_2770);
xor U3410 (N_3410,N_2704,N_2559);
nand U3411 (N_3411,N_2654,N_2465);
nand U3412 (N_3412,N_2074,N_2547);
xnor U3413 (N_3413,N_2707,N_2583);
or U3414 (N_3414,N_2969,N_2869);
xor U3415 (N_3415,N_2096,N_2219);
nor U3416 (N_3416,N_2099,N_2343);
xor U3417 (N_3417,N_2396,N_2772);
nor U3418 (N_3418,N_2473,N_2549);
xor U3419 (N_3419,N_2501,N_2677);
or U3420 (N_3420,N_2624,N_2236);
xor U3421 (N_3421,N_2659,N_2140);
nor U3422 (N_3422,N_2502,N_2004);
xor U3423 (N_3423,N_2857,N_2744);
nor U3424 (N_3424,N_2781,N_2344);
xor U3425 (N_3425,N_2746,N_2494);
nand U3426 (N_3426,N_2566,N_2038);
nor U3427 (N_3427,N_2784,N_2113);
or U3428 (N_3428,N_2575,N_2127);
xor U3429 (N_3429,N_2651,N_2051);
nand U3430 (N_3430,N_2837,N_2015);
xor U3431 (N_3431,N_2821,N_2112);
nor U3432 (N_3432,N_2685,N_2162);
nand U3433 (N_3433,N_2288,N_2515);
and U3434 (N_3434,N_2540,N_2077);
nand U3435 (N_3435,N_2530,N_2514);
nor U3436 (N_3436,N_2191,N_2596);
or U3437 (N_3437,N_2149,N_2736);
nor U3438 (N_3438,N_2572,N_2017);
and U3439 (N_3439,N_2011,N_2079);
and U3440 (N_3440,N_2142,N_2570);
or U3441 (N_3441,N_2467,N_2059);
nand U3442 (N_3442,N_2448,N_2824);
xnor U3443 (N_3443,N_2855,N_2953);
and U3444 (N_3444,N_2611,N_2778);
and U3445 (N_3445,N_2561,N_2801);
xor U3446 (N_3446,N_2951,N_2464);
or U3447 (N_3447,N_2852,N_2919);
xnor U3448 (N_3448,N_2353,N_2386);
or U3449 (N_3449,N_2355,N_2061);
nor U3450 (N_3450,N_2031,N_2506);
or U3451 (N_3451,N_2777,N_2958);
xor U3452 (N_3452,N_2184,N_2105);
nand U3453 (N_3453,N_2009,N_2470);
xor U3454 (N_3454,N_2964,N_2150);
and U3455 (N_3455,N_2742,N_2384);
nand U3456 (N_3456,N_2383,N_2673);
xnor U3457 (N_3457,N_2380,N_2181);
and U3458 (N_3458,N_2402,N_2711);
nand U3459 (N_3459,N_2858,N_2496);
xnor U3460 (N_3460,N_2229,N_2325);
nor U3461 (N_3461,N_2603,N_2793);
and U3462 (N_3462,N_2252,N_2207);
or U3463 (N_3463,N_2173,N_2937);
or U3464 (N_3464,N_2827,N_2151);
xnor U3465 (N_3465,N_2240,N_2187);
nand U3466 (N_3466,N_2700,N_2779);
xor U3467 (N_3467,N_2574,N_2379);
and U3468 (N_3468,N_2595,N_2485);
or U3469 (N_3469,N_2552,N_2277);
xor U3470 (N_3470,N_2992,N_2231);
nand U3471 (N_3471,N_2877,N_2001);
and U3472 (N_3472,N_2915,N_2724);
or U3473 (N_3473,N_2190,N_2091);
and U3474 (N_3474,N_2433,N_2138);
xor U3475 (N_3475,N_2614,N_2828);
and U3476 (N_3476,N_2674,N_2655);
and U3477 (N_3477,N_2928,N_2117);
nand U3478 (N_3478,N_2456,N_2185);
and U3479 (N_3479,N_2296,N_2025);
and U3480 (N_3480,N_2555,N_2440);
and U3481 (N_3481,N_2412,N_2620);
and U3482 (N_3482,N_2131,N_2329);
nand U3483 (N_3483,N_2255,N_2194);
nand U3484 (N_3484,N_2475,N_2106);
xor U3485 (N_3485,N_2627,N_2428);
nor U3486 (N_3486,N_2466,N_2727);
and U3487 (N_3487,N_2125,N_2351);
nor U3488 (N_3488,N_2299,N_2664);
nand U3489 (N_3489,N_2256,N_2081);
or U3490 (N_3490,N_2102,N_2084);
xnor U3491 (N_3491,N_2055,N_2041);
and U3492 (N_3492,N_2357,N_2731);
and U3493 (N_3493,N_2571,N_2445);
xor U3494 (N_3494,N_2303,N_2472);
or U3495 (N_3495,N_2427,N_2273);
nand U3496 (N_3496,N_2183,N_2317);
nand U3497 (N_3497,N_2326,N_2905);
nand U3498 (N_3498,N_2070,N_2893);
nor U3499 (N_3499,N_2752,N_2226);
nor U3500 (N_3500,N_2537,N_2657);
xnor U3501 (N_3501,N_2037,N_2784);
nor U3502 (N_3502,N_2512,N_2058);
nand U3503 (N_3503,N_2615,N_2379);
or U3504 (N_3504,N_2600,N_2714);
nand U3505 (N_3505,N_2979,N_2193);
xor U3506 (N_3506,N_2553,N_2258);
or U3507 (N_3507,N_2793,N_2630);
and U3508 (N_3508,N_2057,N_2567);
nor U3509 (N_3509,N_2584,N_2890);
or U3510 (N_3510,N_2220,N_2832);
nor U3511 (N_3511,N_2107,N_2069);
nand U3512 (N_3512,N_2621,N_2177);
and U3513 (N_3513,N_2033,N_2711);
and U3514 (N_3514,N_2015,N_2373);
or U3515 (N_3515,N_2104,N_2547);
and U3516 (N_3516,N_2270,N_2768);
or U3517 (N_3517,N_2617,N_2760);
nor U3518 (N_3518,N_2010,N_2931);
or U3519 (N_3519,N_2698,N_2781);
xnor U3520 (N_3520,N_2741,N_2300);
nor U3521 (N_3521,N_2409,N_2773);
xor U3522 (N_3522,N_2261,N_2863);
nor U3523 (N_3523,N_2892,N_2875);
nor U3524 (N_3524,N_2484,N_2554);
xnor U3525 (N_3525,N_2626,N_2066);
nand U3526 (N_3526,N_2952,N_2524);
or U3527 (N_3527,N_2253,N_2682);
and U3528 (N_3528,N_2113,N_2397);
or U3529 (N_3529,N_2248,N_2048);
and U3530 (N_3530,N_2491,N_2274);
or U3531 (N_3531,N_2883,N_2071);
nor U3532 (N_3532,N_2321,N_2195);
nor U3533 (N_3533,N_2857,N_2930);
nand U3534 (N_3534,N_2366,N_2847);
xnor U3535 (N_3535,N_2178,N_2479);
xor U3536 (N_3536,N_2271,N_2556);
nor U3537 (N_3537,N_2094,N_2469);
nand U3538 (N_3538,N_2988,N_2427);
nand U3539 (N_3539,N_2075,N_2450);
nor U3540 (N_3540,N_2277,N_2585);
and U3541 (N_3541,N_2030,N_2388);
nor U3542 (N_3542,N_2747,N_2724);
nor U3543 (N_3543,N_2064,N_2676);
or U3544 (N_3544,N_2584,N_2896);
and U3545 (N_3545,N_2979,N_2782);
nor U3546 (N_3546,N_2241,N_2204);
nand U3547 (N_3547,N_2413,N_2119);
xor U3548 (N_3548,N_2574,N_2810);
nand U3549 (N_3549,N_2928,N_2175);
and U3550 (N_3550,N_2603,N_2357);
nor U3551 (N_3551,N_2654,N_2138);
nor U3552 (N_3552,N_2649,N_2988);
or U3553 (N_3553,N_2358,N_2234);
xnor U3554 (N_3554,N_2060,N_2125);
nand U3555 (N_3555,N_2159,N_2412);
and U3556 (N_3556,N_2864,N_2661);
nor U3557 (N_3557,N_2720,N_2515);
or U3558 (N_3558,N_2988,N_2753);
xnor U3559 (N_3559,N_2437,N_2682);
or U3560 (N_3560,N_2668,N_2909);
nor U3561 (N_3561,N_2927,N_2038);
and U3562 (N_3562,N_2064,N_2202);
nor U3563 (N_3563,N_2046,N_2014);
xnor U3564 (N_3564,N_2570,N_2504);
xor U3565 (N_3565,N_2576,N_2828);
nand U3566 (N_3566,N_2871,N_2625);
or U3567 (N_3567,N_2152,N_2984);
xnor U3568 (N_3568,N_2698,N_2769);
nand U3569 (N_3569,N_2290,N_2545);
nor U3570 (N_3570,N_2950,N_2699);
or U3571 (N_3571,N_2613,N_2218);
xnor U3572 (N_3572,N_2481,N_2596);
nor U3573 (N_3573,N_2430,N_2714);
and U3574 (N_3574,N_2872,N_2453);
nand U3575 (N_3575,N_2667,N_2030);
nor U3576 (N_3576,N_2572,N_2451);
and U3577 (N_3577,N_2213,N_2999);
nand U3578 (N_3578,N_2760,N_2613);
nand U3579 (N_3579,N_2237,N_2874);
xnor U3580 (N_3580,N_2331,N_2519);
and U3581 (N_3581,N_2031,N_2329);
and U3582 (N_3582,N_2965,N_2172);
or U3583 (N_3583,N_2141,N_2224);
nor U3584 (N_3584,N_2690,N_2497);
nand U3585 (N_3585,N_2537,N_2494);
xnor U3586 (N_3586,N_2579,N_2791);
nand U3587 (N_3587,N_2204,N_2857);
nor U3588 (N_3588,N_2581,N_2362);
nand U3589 (N_3589,N_2900,N_2483);
nor U3590 (N_3590,N_2232,N_2989);
nor U3591 (N_3591,N_2967,N_2689);
and U3592 (N_3592,N_2962,N_2201);
xnor U3593 (N_3593,N_2745,N_2485);
xor U3594 (N_3594,N_2515,N_2702);
and U3595 (N_3595,N_2303,N_2425);
or U3596 (N_3596,N_2500,N_2192);
and U3597 (N_3597,N_2034,N_2105);
or U3598 (N_3598,N_2804,N_2878);
and U3599 (N_3599,N_2905,N_2513);
nand U3600 (N_3600,N_2792,N_2656);
xor U3601 (N_3601,N_2790,N_2383);
nor U3602 (N_3602,N_2135,N_2776);
nor U3603 (N_3603,N_2434,N_2946);
or U3604 (N_3604,N_2222,N_2145);
xnor U3605 (N_3605,N_2966,N_2018);
xnor U3606 (N_3606,N_2538,N_2703);
or U3607 (N_3607,N_2249,N_2607);
or U3608 (N_3608,N_2982,N_2320);
xnor U3609 (N_3609,N_2023,N_2394);
nor U3610 (N_3610,N_2396,N_2675);
nor U3611 (N_3611,N_2561,N_2625);
nand U3612 (N_3612,N_2770,N_2903);
xor U3613 (N_3613,N_2135,N_2585);
nand U3614 (N_3614,N_2679,N_2332);
xor U3615 (N_3615,N_2028,N_2152);
nor U3616 (N_3616,N_2556,N_2791);
or U3617 (N_3617,N_2419,N_2702);
and U3618 (N_3618,N_2172,N_2772);
nand U3619 (N_3619,N_2845,N_2261);
and U3620 (N_3620,N_2048,N_2146);
and U3621 (N_3621,N_2154,N_2452);
or U3622 (N_3622,N_2299,N_2658);
xnor U3623 (N_3623,N_2111,N_2848);
or U3624 (N_3624,N_2915,N_2960);
and U3625 (N_3625,N_2147,N_2235);
nor U3626 (N_3626,N_2713,N_2978);
and U3627 (N_3627,N_2257,N_2178);
nor U3628 (N_3628,N_2358,N_2539);
or U3629 (N_3629,N_2542,N_2425);
and U3630 (N_3630,N_2738,N_2939);
xor U3631 (N_3631,N_2814,N_2221);
or U3632 (N_3632,N_2020,N_2832);
and U3633 (N_3633,N_2932,N_2364);
xor U3634 (N_3634,N_2042,N_2873);
and U3635 (N_3635,N_2075,N_2966);
nor U3636 (N_3636,N_2424,N_2821);
nor U3637 (N_3637,N_2738,N_2567);
and U3638 (N_3638,N_2749,N_2767);
xnor U3639 (N_3639,N_2887,N_2247);
and U3640 (N_3640,N_2806,N_2959);
and U3641 (N_3641,N_2762,N_2053);
nor U3642 (N_3642,N_2391,N_2834);
nand U3643 (N_3643,N_2144,N_2543);
and U3644 (N_3644,N_2300,N_2040);
or U3645 (N_3645,N_2863,N_2053);
or U3646 (N_3646,N_2443,N_2565);
or U3647 (N_3647,N_2759,N_2892);
or U3648 (N_3648,N_2847,N_2506);
or U3649 (N_3649,N_2661,N_2170);
or U3650 (N_3650,N_2690,N_2840);
or U3651 (N_3651,N_2106,N_2788);
nor U3652 (N_3652,N_2690,N_2232);
nand U3653 (N_3653,N_2640,N_2325);
or U3654 (N_3654,N_2144,N_2548);
or U3655 (N_3655,N_2949,N_2489);
nor U3656 (N_3656,N_2726,N_2999);
or U3657 (N_3657,N_2775,N_2521);
and U3658 (N_3658,N_2756,N_2389);
nor U3659 (N_3659,N_2073,N_2871);
and U3660 (N_3660,N_2282,N_2314);
or U3661 (N_3661,N_2972,N_2710);
or U3662 (N_3662,N_2425,N_2638);
and U3663 (N_3663,N_2106,N_2136);
nor U3664 (N_3664,N_2198,N_2239);
and U3665 (N_3665,N_2988,N_2572);
and U3666 (N_3666,N_2102,N_2356);
and U3667 (N_3667,N_2915,N_2264);
or U3668 (N_3668,N_2458,N_2389);
nor U3669 (N_3669,N_2014,N_2392);
nor U3670 (N_3670,N_2842,N_2355);
nor U3671 (N_3671,N_2019,N_2253);
xnor U3672 (N_3672,N_2154,N_2239);
nand U3673 (N_3673,N_2278,N_2843);
nand U3674 (N_3674,N_2416,N_2731);
xor U3675 (N_3675,N_2015,N_2832);
xor U3676 (N_3676,N_2629,N_2910);
xnor U3677 (N_3677,N_2109,N_2839);
nor U3678 (N_3678,N_2823,N_2060);
xor U3679 (N_3679,N_2066,N_2499);
nor U3680 (N_3680,N_2356,N_2888);
nor U3681 (N_3681,N_2317,N_2944);
and U3682 (N_3682,N_2918,N_2695);
or U3683 (N_3683,N_2311,N_2535);
xor U3684 (N_3684,N_2591,N_2354);
xnor U3685 (N_3685,N_2383,N_2107);
nor U3686 (N_3686,N_2715,N_2871);
or U3687 (N_3687,N_2760,N_2848);
or U3688 (N_3688,N_2995,N_2507);
nand U3689 (N_3689,N_2655,N_2104);
or U3690 (N_3690,N_2122,N_2033);
nor U3691 (N_3691,N_2321,N_2861);
nand U3692 (N_3692,N_2329,N_2184);
nand U3693 (N_3693,N_2226,N_2888);
or U3694 (N_3694,N_2016,N_2561);
and U3695 (N_3695,N_2071,N_2673);
and U3696 (N_3696,N_2936,N_2481);
nor U3697 (N_3697,N_2850,N_2673);
nor U3698 (N_3698,N_2955,N_2668);
and U3699 (N_3699,N_2829,N_2616);
nor U3700 (N_3700,N_2450,N_2594);
nand U3701 (N_3701,N_2270,N_2042);
nand U3702 (N_3702,N_2292,N_2918);
nor U3703 (N_3703,N_2131,N_2219);
nor U3704 (N_3704,N_2016,N_2898);
nand U3705 (N_3705,N_2495,N_2649);
nor U3706 (N_3706,N_2547,N_2979);
or U3707 (N_3707,N_2476,N_2606);
and U3708 (N_3708,N_2934,N_2362);
nor U3709 (N_3709,N_2801,N_2246);
or U3710 (N_3710,N_2761,N_2551);
or U3711 (N_3711,N_2662,N_2199);
xor U3712 (N_3712,N_2662,N_2973);
and U3713 (N_3713,N_2757,N_2644);
nor U3714 (N_3714,N_2860,N_2171);
and U3715 (N_3715,N_2096,N_2246);
or U3716 (N_3716,N_2507,N_2346);
nor U3717 (N_3717,N_2781,N_2191);
xnor U3718 (N_3718,N_2473,N_2631);
and U3719 (N_3719,N_2974,N_2605);
xnor U3720 (N_3720,N_2938,N_2604);
and U3721 (N_3721,N_2163,N_2106);
nand U3722 (N_3722,N_2105,N_2275);
nor U3723 (N_3723,N_2436,N_2676);
and U3724 (N_3724,N_2063,N_2252);
nand U3725 (N_3725,N_2360,N_2089);
xnor U3726 (N_3726,N_2562,N_2172);
xor U3727 (N_3727,N_2980,N_2705);
or U3728 (N_3728,N_2758,N_2416);
nor U3729 (N_3729,N_2990,N_2817);
nand U3730 (N_3730,N_2401,N_2719);
or U3731 (N_3731,N_2923,N_2893);
nand U3732 (N_3732,N_2327,N_2738);
nand U3733 (N_3733,N_2537,N_2268);
xor U3734 (N_3734,N_2444,N_2798);
nor U3735 (N_3735,N_2732,N_2687);
and U3736 (N_3736,N_2405,N_2542);
xor U3737 (N_3737,N_2328,N_2789);
xnor U3738 (N_3738,N_2545,N_2563);
nand U3739 (N_3739,N_2852,N_2255);
or U3740 (N_3740,N_2980,N_2733);
xor U3741 (N_3741,N_2768,N_2859);
and U3742 (N_3742,N_2817,N_2179);
or U3743 (N_3743,N_2264,N_2408);
xor U3744 (N_3744,N_2574,N_2566);
xnor U3745 (N_3745,N_2968,N_2793);
and U3746 (N_3746,N_2400,N_2894);
xor U3747 (N_3747,N_2088,N_2149);
nor U3748 (N_3748,N_2350,N_2141);
and U3749 (N_3749,N_2993,N_2104);
and U3750 (N_3750,N_2762,N_2107);
and U3751 (N_3751,N_2020,N_2235);
and U3752 (N_3752,N_2912,N_2091);
or U3753 (N_3753,N_2205,N_2378);
and U3754 (N_3754,N_2172,N_2467);
nand U3755 (N_3755,N_2472,N_2412);
and U3756 (N_3756,N_2317,N_2178);
or U3757 (N_3757,N_2432,N_2546);
and U3758 (N_3758,N_2059,N_2234);
or U3759 (N_3759,N_2700,N_2760);
xor U3760 (N_3760,N_2125,N_2488);
nand U3761 (N_3761,N_2580,N_2428);
nor U3762 (N_3762,N_2921,N_2501);
xor U3763 (N_3763,N_2409,N_2075);
or U3764 (N_3764,N_2902,N_2836);
and U3765 (N_3765,N_2559,N_2975);
and U3766 (N_3766,N_2818,N_2066);
nand U3767 (N_3767,N_2418,N_2336);
nand U3768 (N_3768,N_2953,N_2271);
and U3769 (N_3769,N_2743,N_2202);
nor U3770 (N_3770,N_2539,N_2409);
or U3771 (N_3771,N_2147,N_2297);
nand U3772 (N_3772,N_2160,N_2862);
xnor U3773 (N_3773,N_2090,N_2864);
and U3774 (N_3774,N_2091,N_2026);
or U3775 (N_3775,N_2371,N_2439);
xnor U3776 (N_3776,N_2371,N_2981);
nand U3777 (N_3777,N_2560,N_2939);
and U3778 (N_3778,N_2808,N_2624);
nor U3779 (N_3779,N_2566,N_2491);
or U3780 (N_3780,N_2956,N_2121);
nor U3781 (N_3781,N_2013,N_2359);
xor U3782 (N_3782,N_2177,N_2229);
and U3783 (N_3783,N_2471,N_2263);
nand U3784 (N_3784,N_2946,N_2378);
nor U3785 (N_3785,N_2119,N_2405);
xnor U3786 (N_3786,N_2551,N_2292);
or U3787 (N_3787,N_2324,N_2825);
or U3788 (N_3788,N_2059,N_2041);
nand U3789 (N_3789,N_2349,N_2938);
or U3790 (N_3790,N_2499,N_2228);
or U3791 (N_3791,N_2234,N_2147);
nor U3792 (N_3792,N_2918,N_2341);
nor U3793 (N_3793,N_2185,N_2524);
or U3794 (N_3794,N_2730,N_2473);
and U3795 (N_3795,N_2515,N_2255);
nand U3796 (N_3796,N_2547,N_2667);
or U3797 (N_3797,N_2224,N_2882);
nor U3798 (N_3798,N_2490,N_2560);
xnor U3799 (N_3799,N_2581,N_2217);
or U3800 (N_3800,N_2924,N_2814);
or U3801 (N_3801,N_2555,N_2730);
xor U3802 (N_3802,N_2961,N_2960);
nand U3803 (N_3803,N_2914,N_2574);
nor U3804 (N_3804,N_2236,N_2636);
nand U3805 (N_3805,N_2294,N_2424);
nand U3806 (N_3806,N_2157,N_2456);
nand U3807 (N_3807,N_2342,N_2197);
or U3808 (N_3808,N_2110,N_2588);
xnor U3809 (N_3809,N_2941,N_2111);
nor U3810 (N_3810,N_2882,N_2934);
or U3811 (N_3811,N_2847,N_2578);
xor U3812 (N_3812,N_2785,N_2447);
or U3813 (N_3813,N_2658,N_2326);
xnor U3814 (N_3814,N_2090,N_2350);
or U3815 (N_3815,N_2368,N_2113);
and U3816 (N_3816,N_2432,N_2110);
xnor U3817 (N_3817,N_2735,N_2928);
and U3818 (N_3818,N_2014,N_2432);
and U3819 (N_3819,N_2352,N_2222);
and U3820 (N_3820,N_2004,N_2368);
or U3821 (N_3821,N_2844,N_2297);
and U3822 (N_3822,N_2372,N_2630);
xor U3823 (N_3823,N_2049,N_2855);
nor U3824 (N_3824,N_2818,N_2085);
nand U3825 (N_3825,N_2560,N_2187);
or U3826 (N_3826,N_2507,N_2090);
nand U3827 (N_3827,N_2942,N_2237);
xnor U3828 (N_3828,N_2878,N_2877);
and U3829 (N_3829,N_2635,N_2188);
nand U3830 (N_3830,N_2954,N_2593);
nor U3831 (N_3831,N_2825,N_2957);
nand U3832 (N_3832,N_2986,N_2905);
or U3833 (N_3833,N_2061,N_2609);
or U3834 (N_3834,N_2693,N_2445);
nor U3835 (N_3835,N_2079,N_2066);
or U3836 (N_3836,N_2272,N_2650);
xor U3837 (N_3837,N_2931,N_2255);
or U3838 (N_3838,N_2951,N_2091);
and U3839 (N_3839,N_2089,N_2553);
xor U3840 (N_3840,N_2054,N_2189);
or U3841 (N_3841,N_2595,N_2169);
or U3842 (N_3842,N_2898,N_2167);
or U3843 (N_3843,N_2577,N_2795);
or U3844 (N_3844,N_2555,N_2239);
nor U3845 (N_3845,N_2935,N_2333);
xnor U3846 (N_3846,N_2175,N_2158);
nor U3847 (N_3847,N_2411,N_2974);
and U3848 (N_3848,N_2197,N_2311);
nor U3849 (N_3849,N_2257,N_2243);
and U3850 (N_3850,N_2650,N_2146);
nand U3851 (N_3851,N_2525,N_2877);
xor U3852 (N_3852,N_2117,N_2711);
xor U3853 (N_3853,N_2552,N_2309);
or U3854 (N_3854,N_2620,N_2609);
or U3855 (N_3855,N_2276,N_2067);
xor U3856 (N_3856,N_2541,N_2716);
nand U3857 (N_3857,N_2267,N_2682);
nand U3858 (N_3858,N_2982,N_2335);
or U3859 (N_3859,N_2160,N_2442);
or U3860 (N_3860,N_2555,N_2274);
nand U3861 (N_3861,N_2326,N_2557);
xor U3862 (N_3862,N_2782,N_2700);
or U3863 (N_3863,N_2816,N_2851);
and U3864 (N_3864,N_2365,N_2729);
xor U3865 (N_3865,N_2357,N_2558);
xor U3866 (N_3866,N_2912,N_2916);
nand U3867 (N_3867,N_2426,N_2366);
nor U3868 (N_3868,N_2606,N_2823);
xnor U3869 (N_3869,N_2779,N_2648);
or U3870 (N_3870,N_2419,N_2133);
nand U3871 (N_3871,N_2067,N_2037);
or U3872 (N_3872,N_2485,N_2900);
or U3873 (N_3873,N_2702,N_2168);
nand U3874 (N_3874,N_2155,N_2594);
xor U3875 (N_3875,N_2696,N_2599);
xnor U3876 (N_3876,N_2593,N_2517);
xor U3877 (N_3877,N_2047,N_2212);
or U3878 (N_3878,N_2989,N_2213);
nand U3879 (N_3879,N_2654,N_2884);
nor U3880 (N_3880,N_2605,N_2627);
xor U3881 (N_3881,N_2556,N_2009);
xor U3882 (N_3882,N_2628,N_2297);
or U3883 (N_3883,N_2195,N_2988);
xnor U3884 (N_3884,N_2542,N_2745);
or U3885 (N_3885,N_2195,N_2025);
nand U3886 (N_3886,N_2279,N_2258);
nand U3887 (N_3887,N_2247,N_2417);
and U3888 (N_3888,N_2735,N_2993);
and U3889 (N_3889,N_2014,N_2952);
nand U3890 (N_3890,N_2659,N_2263);
or U3891 (N_3891,N_2925,N_2364);
nor U3892 (N_3892,N_2173,N_2256);
and U3893 (N_3893,N_2514,N_2846);
xor U3894 (N_3894,N_2439,N_2637);
nand U3895 (N_3895,N_2401,N_2173);
or U3896 (N_3896,N_2701,N_2643);
or U3897 (N_3897,N_2577,N_2679);
or U3898 (N_3898,N_2721,N_2265);
nand U3899 (N_3899,N_2295,N_2521);
and U3900 (N_3900,N_2280,N_2532);
or U3901 (N_3901,N_2786,N_2347);
and U3902 (N_3902,N_2260,N_2774);
and U3903 (N_3903,N_2003,N_2835);
xnor U3904 (N_3904,N_2961,N_2495);
xor U3905 (N_3905,N_2591,N_2619);
xnor U3906 (N_3906,N_2985,N_2586);
nand U3907 (N_3907,N_2152,N_2873);
nand U3908 (N_3908,N_2920,N_2553);
nand U3909 (N_3909,N_2317,N_2749);
or U3910 (N_3910,N_2765,N_2312);
xor U3911 (N_3911,N_2696,N_2729);
xor U3912 (N_3912,N_2971,N_2111);
nor U3913 (N_3913,N_2251,N_2553);
and U3914 (N_3914,N_2853,N_2582);
nor U3915 (N_3915,N_2846,N_2958);
nor U3916 (N_3916,N_2333,N_2786);
xor U3917 (N_3917,N_2394,N_2798);
and U3918 (N_3918,N_2181,N_2973);
nand U3919 (N_3919,N_2967,N_2423);
nand U3920 (N_3920,N_2571,N_2228);
nor U3921 (N_3921,N_2212,N_2158);
nor U3922 (N_3922,N_2283,N_2626);
xnor U3923 (N_3923,N_2080,N_2295);
and U3924 (N_3924,N_2130,N_2997);
nor U3925 (N_3925,N_2409,N_2006);
nand U3926 (N_3926,N_2954,N_2387);
and U3927 (N_3927,N_2059,N_2475);
xor U3928 (N_3928,N_2296,N_2863);
xor U3929 (N_3929,N_2026,N_2461);
nand U3930 (N_3930,N_2208,N_2434);
or U3931 (N_3931,N_2291,N_2484);
xor U3932 (N_3932,N_2561,N_2295);
xnor U3933 (N_3933,N_2168,N_2478);
xor U3934 (N_3934,N_2172,N_2043);
and U3935 (N_3935,N_2076,N_2135);
nor U3936 (N_3936,N_2177,N_2815);
nand U3937 (N_3937,N_2190,N_2556);
nand U3938 (N_3938,N_2962,N_2145);
nand U3939 (N_3939,N_2318,N_2453);
or U3940 (N_3940,N_2593,N_2527);
xor U3941 (N_3941,N_2889,N_2545);
and U3942 (N_3942,N_2037,N_2220);
xor U3943 (N_3943,N_2162,N_2919);
nor U3944 (N_3944,N_2432,N_2830);
or U3945 (N_3945,N_2069,N_2659);
nor U3946 (N_3946,N_2456,N_2038);
or U3947 (N_3947,N_2360,N_2608);
nor U3948 (N_3948,N_2868,N_2528);
xor U3949 (N_3949,N_2322,N_2943);
xnor U3950 (N_3950,N_2902,N_2571);
or U3951 (N_3951,N_2550,N_2922);
or U3952 (N_3952,N_2236,N_2863);
and U3953 (N_3953,N_2030,N_2328);
nor U3954 (N_3954,N_2257,N_2536);
and U3955 (N_3955,N_2650,N_2843);
or U3956 (N_3956,N_2718,N_2935);
xnor U3957 (N_3957,N_2304,N_2730);
or U3958 (N_3958,N_2625,N_2728);
and U3959 (N_3959,N_2401,N_2904);
or U3960 (N_3960,N_2609,N_2905);
and U3961 (N_3961,N_2419,N_2297);
xnor U3962 (N_3962,N_2534,N_2643);
nand U3963 (N_3963,N_2750,N_2586);
and U3964 (N_3964,N_2057,N_2358);
nor U3965 (N_3965,N_2168,N_2750);
xor U3966 (N_3966,N_2454,N_2595);
and U3967 (N_3967,N_2362,N_2725);
xor U3968 (N_3968,N_2322,N_2854);
xnor U3969 (N_3969,N_2850,N_2790);
xor U3970 (N_3970,N_2754,N_2302);
nand U3971 (N_3971,N_2868,N_2273);
or U3972 (N_3972,N_2855,N_2260);
nor U3973 (N_3973,N_2282,N_2784);
xnor U3974 (N_3974,N_2412,N_2538);
or U3975 (N_3975,N_2906,N_2647);
nand U3976 (N_3976,N_2265,N_2142);
nand U3977 (N_3977,N_2297,N_2252);
xor U3978 (N_3978,N_2368,N_2696);
xor U3979 (N_3979,N_2646,N_2074);
nand U3980 (N_3980,N_2232,N_2322);
nand U3981 (N_3981,N_2652,N_2100);
nor U3982 (N_3982,N_2237,N_2960);
nand U3983 (N_3983,N_2049,N_2031);
xnor U3984 (N_3984,N_2073,N_2622);
xnor U3985 (N_3985,N_2573,N_2283);
and U3986 (N_3986,N_2536,N_2380);
or U3987 (N_3987,N_2323,N_2617);
nor U3988 (N_3988,N_2060,N_2453);
and U3989 (N_3989,N_2326,N_2624);
nand U3990 (N_3990,N_2738,N_2259);
nor U3991 (N_3991,N_2202,N_2082);
nor U3992 (N_3992,N_2453,N_2992);
nor U3993 (N_3993,N_2144,N_2998);
nor U3994 (N_3994,N_2257,N_2915);
or U3995 (N_3995,N_2940,N_2125);
nor U3996 (N_3996,N_2130,N_2462);
xnor U3997 (N_3997,N_2778,N_2168);
nand U3998 (N_3998,N_2146,N_2803);
xor U3999 (N_3999,N_2363,N_2487);
nor U4000 (N_4000,N_3439,N_3209);
xor U4001 (N_4001,N_3879,N_3019);
nand U4002 (N_4002,N_3229,N_3497);
nand U4003 (N_4003,N_3186,N_3381);
nor U4004 (N_4004,N_3899,N_3978);
nand U4005 (N_4005,N_3580,N_3417);
nor U4006 (N_4006,N_3364,N_3976);
xnor U4007 (N_4007,N_3688,N_3956);
nand U4008 (N_4008,N_3441,N_3894);
or U4009 (N_4009,N_3516,N_3246);
and U4010 (N_4010,N_3714,N_3606);
or U4011 (N_4011,N_3507,N_3334);
nor U4012 (N_4012,N_3251,N_3846);
or U4013 (N_4013,N_3578,N_3941);
xnor U4014 (N_4014,N_3601,N_3177);
nor U4015 (N_4015,N_3961,N_3442);
xor U4016 (N_4016,N_3201,N_3313);
nand U4017 (N_4017,N_3066,N_3435);
xor U4018 (N_4018,N_3451,N_3995);
nor U4019 (N_4019,N_3521,N_3621);
or U4020 (N_4020,N_3812,N_3678);
nand U4021 (N_4021,N_3659,N_3002);
and U4022 (N_4022,N_3420,N_3188);
or U4023 (N_4023,N_3958,N_3180);
nor U4024 (N_4024,N_3550,N_3985);
or U4025 (N_4025,N_3199,N_3003);
xnor U4026 (N_4026,N_3144,N_3754);
or U4027 (N_4027,N_3324,N_3522);
nand U4028 (N_4028,N_3134,N_3018);
or U4029 (N_4029,N_3074,N_3977);
nor U4030 (N_4030,N_3486,N_3929);
and U4031 (N_4031,N_3426,N_3783);
xor U4032 (N_4032,N_3132,N_3967);
or U4033 (N_4033,N_3938,N_3106);
and U4034 (N_4034,N_3457,N_3479);
xnor U4035 (N_4035,N_3296,N_3254);
and U4036 (N_4036,N_3576,N_3989);
nor U4037 (N_4037,N_3255,N_3500);
and U4038 (N_4038,N_3205,N_3249);
or U4039 (N_4039,N_3393,N_3087);
xnor U4040 (N_4040,N_3190,N_3449);
nand U4041 (N_4041,N_3660,N_3928);
and U4042 (N_4042,N_3487,N_3666);
nand U4043 (N_4043,N_3921,N_3837);
xnor U4044 (N_4044,N_3102,N_3603);
and U4045 (N_4045,N_3565,N_3962);
xnor U4046 (N_4046,N_3937,N_3480);
nand U4047 (N_4047,N_3670,N_3455);
xor U4048 (N_4048,N_3013,N_3333);
nand U4049 (N_4049,N_3972,N_3337);
xnor U4050 (N_4050,N_3751,N_3129);
nand U4051 (N_4051,N_3234,N_3864);
and U4052 (N_4052,N_3034,N_3467);
xor U4053 (N_4053,N_3966,N_3308);
xor U4054 (N_4054,N_3561,N_3121);
nand U4055 (N_4055,N_3555,N_3734);
xnor U4056 (N_4056,N_3077,N_3007);
or U4057 (N_4057,N_3567,N_3010);
nor U4058 (N_4058,N_3064,N_3287);
nand U4059 (N_4059,N_3429,N_3416);
or U4060 (N_4060,N_3023,N_3244);
nor U4061 (N_4061,N_3338,N_3679);
xnor U4062 (N_4062,N_3725,N_3206);
nor U4063 (N_4063,N_3015,N_3695);
xnor U4064 (N_4064,N_3027,N_3748);
nand U4065 (N_4065,N_3769,N_3892);
nand U4066 (N_4066,N_3707,N_3261);
xor U4067 (N_4067,N_3822,N_3794);
or U4068 (N_4068,N_3264,N_3026);
xor U4069 (N_4069,N_3503,N_3418);
nand U4070 (N_4070,N_3021,N_3908);
xor U4071 (N_4071,N_3991,N_3940);
nand U4072 (N_4072,N_3654,N_3331);
nand U4073 (N_4073,N_3388,N_3906);
or U4074 (N_4074,N_3189,N_3655);
nor U4075 (N_4075,N_3073,N_3422);
or U4076 (N_4076,N_3675,N_3615);
and U4077 (N_4077,N_3971,N_3488);
nand U4078 (N_4078,N_3008,N_3147);
or U4079 (N_4079,N_3665,N_3166);
nor U4080 (N_4080,N_3499,N_3598);
xor U4081 (N_4081,N_3236,N_3932);
or U4082 (N_4082,N_3609,N_3288);
and U4083 (N_4083,N_3881,N_3557);
and U4084 (N_4084,N_3588,N_3385);
and U4085 (N_4085,N_3570,N_3095);
nor U4086 (N_4086,N_3365,N_3515);
xor U4087 (N_4087,N_3523,N_3868);
nor U4088 (N_4088,N_3548,N_3344);
or U4089 (N_4089,N_3415,N_3776);
nand U4090 (N_4090,N_3446,N_3240);
and U4091 (N_4091,N_3512,N_3233);
or U4092 (N_4092,N_3491,N_3610);
nor U4093 (N_4093,N_3283,N_3832);
nand U4094 (N_4094,N_3104,N_3960);
nor U4095 (N_4095,N_3402,N_3247);
nor U4096 (N_4096,N_3726,N_3080);
nand U4097 (N_4097,N_3860,N_3181);
nand U4098 (N_4098,N_3857,N_3524);
xor U4099 (N_4099,N_3278,N_3594);
xnor U4100 (N_4100,N_3505,N_3668);
xnor U4101 (N_4101,N_3401,N_3841);
nor U4102 (N_4102,N_3145,N_3886);
or U4103 (N_4103,N_3819,N_3999);
and U4104 (N_4104,N_3112,N_3099);
nand U4105 (N_4105,N_3183,N_3838);
or U4106 (N_4106,N_3988,N_3445);
or U4107 (N_4107,N_3107,N_3475);
or U4108 (N_4108,N_3825,N_3680);
or U4109 (N_4109,N_3597,N_3810);
nand U4110 (N_4110,N_3872,N_3865);
nand U4111 (N_4111,N_3752,N_3400);
xnor U4112 (N_4112,N_3032,N_3114);
nor U4113 (N_4113,N_3215,N_3624);
nor U4114 (N_4114,N_3849,N_3437);
nor U4115 (N_4115,N_3572,N_3395);
or U4116 (N_4116,N_3788,N_3672);
nor U4117 (N_4117,N_3139,N_3973);
and U4118 (N_4118,N_3438,N_3709);
nor U4119 (N_4119,N_3773,N_3454);
nand U4120 (N_4120,N_3744,N_3760);
or U4121 (N_4121,N_3224,N_3765);
nand U4122 (N_4122,N_3762,N_3544);
and U4123 (N_4123,N_3753,N_3631);
nor U4124 (N_4124,N_3065,N_3697);
and U4125 (N_4125,N_3396,N_3954);
xor U4126 (N_4126,N_3738,N_3489);
and U4127 (N_4127,N_3893,N_3780);
or U4128 (N_4128,N_3115,N_3390);
nand U4129 (N_4129,N_3062,N_3558);
and U4130 (N_4130,N_3270,N_3309);
nand U4131 (N_4131,N_3903,N_3646);
and U4132 (N_4132,N_3399,N_3828);
or U4133 (N_4133,N_3485,N_3377);
and U4134 (N_4134,N_3269,N_3963);
xor U4135 (N_4135,N_3847,N_3593);
nor U4136 (N_4136,N_3855,N_3332);
and U4137 (N_4137,N_3260,N_3817);
xnor U4138 (N_4138,N_3017,N_3133);
xnor U4139 (N_4139,N_3901,N_3407);
nand U4140 (N_4140,N_3252,N_3859);
or U4141 (N_4141,N_3876,N_3771);
nand U4142 (N_4142,N_3952,N_3001);
or U4143 (N_4143,N_3996,N_3258);
or U4144 (N_4144,N_3834,N_3242);
or U4145 (N_4145,N_3858,N_3067);
or U4146 (N_4146,N_3814,N_3203);
nor U4147 (N_4147,N_3174,N_3117);
xnor U4148 (N_4148,N_3361,N_3448);
nand U4149 (N_4149,N_3577,N_3699);
nor U4150 (N_4150,N_3775,N_3232);
or U4151 (N_4151,N_3740,N_3428);
and U4152 (N_4152,N_3757,N_3531);
or U4153 (N_4153,N_3942,N_3343);
xnor U4154 (N_4154,N_3784,N_3118);
nand U4155 (N_4155,N_3267,N_3944);
nor U4156 (N_4156,N_3673,N_3044);
nand U4157 (N_4157,N_3807,N_3824);
nand U4158 (N_4158,N_3727,N_3239);
and U4159 (N_4159,N_3829,N_3998);
and U4160 (N_4160,N_3900,N_3994);
and U4161 (N_4161,N_3347,N_3719);
nor U4162 (N_4162,N_3284,N_3140);
and U4163 (N_4163,N_3421,N_3518);
and U4164 (N_4164,N_3282,N_3669);
nor U4165 (N_4165,N_3579,N_3878);
nor U4166 (N_4166,N_3405,N_3702);
nand U4167 (N_4167,N_3533,N_3854);
xnor U4168 (N_4168,N_3194,N_3667);
nor U4169 (N_4169,N_3919,N_3917);
nor U4170 (N_4170,N_3210,N_3048);
and U4171 (N_4171,N_3185,N_3339);
or U4172 (N_4172,N_3092,N_3148);
nand U4173 (N_4173,N_3465,N_3778);
nor U4174 (N_4174,N_3664,N_3804);
nand U4175 (N_4175,N_3009,N_3161);
nand U4176 (N_4176,N_3294,N_3471);
and U4177 (N_4177,N_3627,N_3110);
or U4178 (N_4178,N_3536,N_3447);
nand U4179 (N_4179,N_3800,N_3717);
nor U4180 (N_4180,N_3649,N_3035);
and U4181 (N_4181,N_3852,N_3947);
nand U4182 (N_4182,N_3196,N_3217);
and U4183 (N_4183,N_3534,N_3028);
and U4184 (N_4184,N_3614,N_3378);
nand U4185 (N_4185,N_3850,N_3770);
xnor U4186 (N_4186,N_3936,N_3453);
or U4187 (N_4187,N_3158,N_3354);
or U4188 (N_4188,N_3081,N_3136);
nor U4189 (N_4189,N_3305,N_3633);
or U4190 (N_4190,N_3352,N_3708);
nor U4191 (N_4191,N_3314,N_3241);
or U4192 (N_4192,N_3359,N_3192);
or U4193 (N_4193,N_3330,N_3861);
xor U4194 (N_4194,N_3526,N_3692);
or U4195 (N_4195,N_3404,N_3358);
and U4196 (N_4196,N_3120,N_3142);
or U4197 (N_4197,N_3295,N_3566);
and U4198 (N_4198,N_3041,N_3289);
xor U4199 (N_4199,N_3355,N_3266);
and U4200 (N_4200,N_3423,N_3443);
nand U4201 (N_4201,N_3513,N_3767);
xnor U4202 (N_4202,N_3583,N_3363);
nand U4203 (N_4203,N_3279,N_3605);
or U4204 (N_4204,N_3732,N_3463);
or U4205 (N_4205,N_3571,N_3406);
or U4206 (N_4206,N_3298,N_3758);
or U4207 (N_4207,N_3974,N_3212);
nand U4208 (N_4208,N_3257,N_3816);
nand U4209 (N_4209,N_3167,N_3641);
or U4210 (N_4210,N_3141,N_3634);
and U4211 (N_4211,N_3712,N_3366);
or U4212 (N_4212,N_3763,N_3096);
xor U4213 (N_4213,N_3651,N_3097);
nor U4214 (N_4214,N_3884,N_3844);
and U4215 (N_4215,N_3663,N_3341);
nand U4216 (N_4216,N_3169,N_3801);
nand U4217 (N_4217,N_3591,N_3535);
or U4218 (N_4218,N_3020,N_3509);
or U4219 (N_4219,N_3173,N_3596);
or U4220 (N_4220,N_3336,N_3731);
nor U4221 (N_4221,N_3179,N_3376);
nor U4222 (N_4222,N_3722,N_3766);
or U4223 (N_4223,N_3030,N_3785);
nand U4224 (N_4224,N_3683,N_3460);
nor U4225 (N_4225,N_3368,N_3642);
nand U4226 (N_4226,N_3885,N_3711);
nor U4227 (N_4227,N_3890,N_3623);
nor U4228 (N_4228,N_3113,N_3170);
nand U4229 (N_4229,N_3587,N_3645);
nor U4230 (N_4230,N_3414,N_3301);
nor U4231 (N_4231,N_3951,N_3316);
nand U4232 (N_4232,N_3078,N_3387);
and U4233 (N_4233,N_3584,N_3302);
nor U4234 (N_4234,N_3383,N_3389);
xor U4235 (N_4235,N_3686,N_3369);
xor U4236 (N_4236,N_3700,N_3052);
or U4237 (N_4237,N_3705,N_3815);
xor U4238 (N_4238,N_3000,N_3060);
nand U4239 (N_4239,N_3636,N_3508);
nand U4240 (N_4240,N_3737,N_3933);
or U4241 (N_4241,N_3853,N_3045);
xor U4242 (N_4242,N_3863,N_3093);
nor U4243 (N_4243,N_3154,N_3650);
or U4244 (N_4244,N_3281,N_3547);
and U4245 (N_4245,N_3831,N_3882);
and U4246 (N_4246,N_3468,N_3756);
and U4247 (N_4247,N_3676,N_3582);
and U4248 (N_4248,N_3345,N_3628);
nor U4249 (N_4249,N_3063,N_3741);
xnor U4250 (N_4250,N_3128,N_3079);
nor U4251 (N_4251,N_3532,N_3564);
nand U4252 (N_4252,N_3806,N_3713);
nor U4253 (N_4253,N_3470,N_3473);
nand U4254 (N_4254,N_3585,N_3721);
nand U4255 (N_4255,N_3682,N_3061);
or U4256 (N_4256,N_3984,N_3303);
or U4257 (N_4257,N_3285,N_3123);
or U4258 (N_4258,N_3743,N_3476);
nand U4259 (N_4259,N_3091,N_3346);
or U4260 (N_4260,N_3716,N_3504);
nand U4261 (N_4261,N_3350,N_3348);
xnor U4262 (N_4262,N_3604,N_3506);
nand U4263 (N_4263,N_3652,N_3552);
xor U4264 (N_4264,N_3216,N_3159);
and U4265 (N_4265,N_3012,N_3862);
nor U4266 (N_4266,N_3790,N_3004);
or U4267 (N_4267,N_3275,N_3360);
nand U4268 (N_4268,N_3306,N_3502);
or U4269 (N_4269,N_3638,N_3452);
xor U4270 (N_4270,N_3704,N_3927);
nand U4271 (N_4271,N_3379,N_3321);
nor U4272 (N_4272,N_3643,N_3171);
xor U4273 (N_4273,N_3342,N_3070);
nor U4274 (N_4274,N_3759,N_3156);
and U4275 (N_4275,N_3193,N_3746);
and U4276 (N_4276,N_3982,N_3461);
or U4277 (N_4277,N_3276,N_3436);
and U4278 (N_4278,N_3225,N_3105);
xnor U4279 (N_4279,N_3075,N_3808);
and U4280 (N_4280,N_3155,N_3701);
or U4281 (N_4281,N_3029,N_3312);
or U4282 (N_4282,N_3510,N_3116);
nand U4283 (N_4283,N_3235,N_3519);
nand U4284 (N_4284,N_3813,N_3291);
or U4285 (N_4285,N_3484,N_3130);
xor U4286 (N_4286,N_3011,N_3057);
and U4287 (N_4287,N_3213,N_3033);
or U4288 (N_4288,N_3979,N_3164);
and U4289 (N_4289,N_3602,N_3540);
nor U4290 (N_4290,N_3218,N_3970);
nor U4291 (N_4291,N_3042,N_3089);
or U4292 (N_4292,N_3419,N_3968);
nor U4293 (N_4293,N_3211,N_3054);
and U4294 (N_4294,N_3595,N_3362);
or U4295 (N_4295,N_3082,N_3589);
nor U4296 (N_4296,N_3798,N_3792);
or U4297 (N_4297,N_3153,N_3883);
xor U4298 (N_4298,N_3072,N_3948);
nand U4299 (N_4299,N_3227,N_3990);
xnor U4300 (N_4300,N_3617,N_3228);
xnor U4301 (N_4301,N_3297,N_3930);
nand U4302 (N_4302,N_3630,N_3411);
xor U4303 (N_4303,N_3736,N_3273);
nand U4304 (N_4304,N_3823,N_3101);
or U4305 (N_4305,N_3049,N_3934);
nand U4306 (N_4306,N_3175,N_3318);
and U4307 (N_4307,N_3924,N_3820);
nor U4308 (N_4308,N_3625,N_3554);
or U4309 (N_4309,N_3277,N_3478);
or U4310 (N_4310,N_3993,N_3237);
nor U4311 (N_4311,N_3922,N_3323);
nor U4312 (N_4312,N_3317,N_3626);
nor U4313 (N_4313,N_3833,N_3613);
nor U4314 (N_4314,N_3710,N_3459);
nand U4315 (N_4315,N_3322,N_3162);
and U4316 (N_4316,N_3644,N_3618);
or U4317 (N_4317,N_3474,N_3867);
nor U4318 (N_4318,N_3047,N_3635);
xor U4319 (N_4319,N_3085,N_3542);
and U4320 (N_4320,N_3843,N_3037);
xor U4321 (N_4321,N_3600,N_3839);
nor U4322 (N_4322,N_3907,N_3747);
or U4323 (N_4323,N_3648,N_3925);
or U4324 (N_4324,N_3926,N_3498);
nand U4325 (N_4325,N_3913,N_3681);
or U4326 (N_4326,N_3492,N_3527);
and U4327 (N_4327,N_3969,N_3517);
xor U4328 (N_4328,N_3469,N_3674);
nor U4329 (N_4329,N_3562,N_3198);
or U4330 (N_4330,N_3184,N_3898);
nor U4331 (N_4331,N_3689,N_3290);
nand U4332 (N_4332,N_3069,N_3611);
xnor U4333 (N_4333,N_3549,N_3202);
nor U4334 (N_4334,N_3458,N_3071);
xnor U4335 (N_4335,N_3911,N_3772);
nor U4336 (N_4336,N_3980,N_3918);
and U4337 (N_4337,N_3799,N_3250);
or U4338 (N_4338,N_3545,N_3653);
or U4339 (N_4339,N_3394,N_3889);
xor U4340 (N_4340,N_3386,N_3300);
or U4341 (N_4341,N_3450,N_3981);
nor U4342 (N_4342,N_3274,N_3887);
or U4343 (N_4343,N_3656,N_3943);
nand U4344 (N_4344,N_3151,N_3373);
xnor U4345 (N_4345,N_3372,N_3735);
and U4346 (N_4346,N_3127,N_3723);
nand U4347 (N_4347,N_3616,N_3214);
nor U4348 (N_4348,N_3100,N_3742);
or U4349 (N_4349,N_3685,N_3088);
and U4350 (N_4350,N_3612,N_3329);
or U4351 (N_4351,N_3511,N_3168);
and U4352 (N_4352,N_3403,N_3891);
or U4353 (N_4353,N_3083,N_3223);
nand U4354 (N_4354,N_3076,N_3146);
and U4355 (N_4355,N_3231,N_3043);
nand U4356 (N_4356,N_3408,N_3207);
or U4357 (N_4357,N_3870,N_3541);
and U4358 (N_4358,N_3357,N_3835);
nand U4359 (N_4359,N_3909,N_3124);
and U4360 (N_4360,N_3326,N_3152);
or U4361 (N_4361,N_3050,N_3764);
xor U4362 (N_4362,N_3456,N_3874);
and U4363 (N_4363,N_3693,N_3657);
and U4364 (N_4364,N_3964,N_3126);
xor U4365 (N_4365,N_3574,N_3219);
and U4366 (N_4366,N_3434,N_3569);
and U4367 (N_4367,N_3483,N_3559);
xor U4368 (N_4368,N_3031,N_3715);
and U4369 (N_4369,N_3975,N_3182);
nand U4370 (N_4370,N_3983,N_3818);
or U4371 (N_4371,N_3265,N_3671);
nor U4372 (N_4372,N_3292,N_3959);
xnor U4373 (N_4373,N_3755,N_3325);
nor U4374 (N_4374,N_3398,N_3382);
or U4375 (N_4375,N_3014,N_3622);
nand U4376 (N_4376,N_3793,N_3157);
and U4377 (N_4377,N_3724,N_3262);
nand U4378 (N_4378,N_3703,N_3094);
xnor U4379 (N_4379,N_3424,N_3084);
nand U4380 (N_4380,N_3840,N_3946);
nand U4381 (N_4381,N_3811,N_3315);
or U4382 (N_4382,N_3912,N_3481);
and U4383 (N_4383,N_3706,N_3789);
or U4384 (N_4384,N_3556,N_3895);
nand U4385 (N_4385,N_3327,N_3586);
nand U4386 (N_4386,N_3135,N_3501);
nand U4387 (N_4387,N_3340,N_3370);
and U4388 (N_4388,N_3953,N_3138);
nand U4389 (N_4389,N_3195,N_3935);
nand U4390 (N_4390,N_3493,N_3068);
or U4391 (N_4391,N_3684,N_3410);
or U4392 (N_4392,N_3514,N_3696);
nand U4393 (N_4393,N_3529,N_3950);
xor U4394 (N_4394,N_3016,N_3902);
or U4395 (N_4395,N_3425,N_3774);
xnor U4396 (N_4396,N_3024,N_3896);
and U4397 (N_4397,N_3607,N_3090);
nor U4398 (N_4398,N_3647,N_3039);
xor U4399 (N_4399,N_3728,N_3022);
nand U4400 (N_4400,N_3871,N_3374);
xor U4401 (N_4401,N_3433,N_3413);
nor U4402 (N_4402,N_3149,N_3494);
xor U4403 (N_4403,N_3304,N_3915);
nand U4404 (N_4404,N_3830,N_3197);
and U4405 (N_4405,N_3055,N_3619);
xnor U4406 (N_4406,N_3351,N_3957);
xnor U4407 (N_4407,N_3786,N_3945);
or U4408 (N_4408,N_3826,N_3581);
nand U4409 (N_4409,N_3640,N_3165);
and U4410 (N_4410,N_3103,N_3280);
xor U4411 (N_4411,N_3477,N_3910);
xnor U4412 (N_4412,N_3472,N_3661);
xnor U4413 (N_4413,N_3006,N_3856);
xnor U4414 (N_4414,N_3191,N_3328);
or U4415 (N_4415,N_3904,N_3923);
nor U4416 (N_4416,N_3310,N_3431);
and U4417 (N_4417,N_3931,N_3495);
and U4418 (N_4418,N_3380,N_3590);
xor U4419 (N_4419,N_3391,N_3543);
nand U4420 (N_4420,N_3525,N_3496);
and U4421 (N_4421,N_3307,N_3538);
nor U4422 (N_4422,N_3761,N_3528);
xor U4423 (N_4423,N_3916,N_3539);
xor U4424 (N_4424,N_3729,N_3848);
or U4425 (N_4425,N_3620,N_3965);
nand U4426 (N_4426,N_3220,N_3230);
or U4427 (N_4427,N_3997,N_3733);
and U4428 (N_4428,N_3877,N_3464);
xor U4429 (N_4429,N_3059,N_3392);
and U4430 (N_4430,N_3178,N_3821);
nand U4431 (N_4431,N_3320,N_3568);
nand U4432 (N_4432,N_3111,N_3311);
nor U4433 (N_4433,N_3200,N_3253);
or U4434 (N_4434,N_3805,N_3880);
or U4435 (N_4435,N_3599,N_3888);
and U4436 (N_4436,N_3873,N_3920);
or U4437 (N_4437,N_3781,N_3384);
and U4438 (N_4438,N_3286,N_3397);
xor U4439 (N_4439,N_3272,N_3795);
nor U4440 (N_4440,N_3036,N_3356);
or U4441 (N_4441,N_3108,N_3551);
and U4442 (N_4442,N_3632,N_3268);
nor U4443 (N_4443,N_3827,N_3629);
xnor U4444 (N_4444,N_3259,N_3639);
nor U4445 (N_4445,N_3745,N_3730);
and U4446 (N_4446,N_3694,N_3739);
nor U4447 (N_4447,N_3086,N_3779);
and U4448 (N_4448,N_3851,N_3546);
nand U4449 (N_4449,N_3119,N_3122);
nor U4450 (N_4450,N_3263,N_3462);
or U4451 (N_4451,N_3005,N_3791);
and U4452 (N_4452,N_3143,N_3271);
nor U4453 (N_4453,N_3208,N_3520);
or U4454 (N_4454,N_3226,N_3248);
xnor U4455 (N_4455,N_3949,N_3750);
and U4456 (N_4456,N_3987,N_3137);
nand U4457 (N_4457,N_3836,N_3537);
nand U4458 (N_4458,N_3046,N_3842);
nor U4459 (N_4459,N_3172,N_3176);
and U4460 (N_4460,N_3299,N_3691);
and U4461 (N_4461,N_3025,N_3809);
xor U4462 (N_4462,N_3677,N_3371);
nand U4463 (N_4463,N_3575,N_3803);
nand U4464 (N_4464,N_3053,N_3637);
xor U4465 (N_4465,N_3845,N_3040);
or U4466 (N_4466,N_3897,N_3427);
nor U4467 (N_4467,N_3440,N_3768);
or U4468 (N_4468,N_3131,N_3658);
nand U4469 (N_4469,N_3690,N_3187);
or U4470 (N_4470,N_3787,N_3430);
nor U4471 (N_4471,N_3125,N_3796);
or U4472 (N_4472,N_3051,N_3992);
and U4473 (N_4473,N_3367,N_3056);
nand U4474 (N_4474,N_3482,N_3245);
or U4475 (N_4475,N_3038,N_3353);
xnor U4476 (N_4476,N_3222,N_3432);
nand U4477 (N_4477,N_3955,N_3238);
xnor U4478 (N_4478,N_3608,N_3058);
nor U4479 (N_4479,N_3720,N_3412);
or U4480 (N_4480,N_3163,N_3150);
or U4481 (N_4481,N_3777,N_3592);
nand U4482 (N_4482,N_3718,N_3098);
or U4483 (N_4483,N_3687,N_3319);
and U4484 (N_4484,N_3782,N_3409);
nor U4485 (N_4485,N_3221,N_3986);
or U4486 (N_4486,N_3905,N_3875);
xor U4487 (N_4487,N_3698,N_3749);
xnor U4488 (N_4488,N_3573,N_3662);
xor U4489 (N_4489,N_3802,N_3204);
nor U4490 (N_4490,N_3293,N_3335);
nor U4491 (N_4491,N_3560,N_3466);
xnor U4492 (N_4492,N_3256,N_3797);
or U4493 (N_4493,N_3160,N_3375);
nor U4494 (N_4494,N_3866,N_3490);
or U4495 (N_4495,N_3869,N_3563);
xnor U4496 (N_4496,N_3914,N_3939);
xnor U4497 (N_4497,N_3109,N_3530);
nand U4498 (N_4498,N_3553,N_3243);
xnor U4499 (N_4499,N_3444,N_3349);
nand U4500 (N_4500,N_3924,N_3045);
xor U4501 (N_4501,N_3541,N_3200);
xnor U4502 (N_4502,N_3879,N_3834);
or U4503 (N_4503,N_3636,N_3156);
and U4504 (N_4504,N_3955,N_3936);
nor U4505 (N_4505,N_3314,N_3378);
xor U4506 (N_4506,N_3590,N_3423);
nor U4507 (N_4507,N_3304,N_3607);
nor U4508 (N_4508,N_3821,N_3166);
nor U4509 (N_4509,N_3546,N_3223);
and U4510 (N_4510,N_3646,N_3824);
and U4511 (N_4511,N_3540,N_3501);
nand U4512 (N_4512,N_3034,N_3575);
or U4513 (N_4513,N_3405,N_3623);
nor U4514 (N_4514,N_3552,N_3166);
nor U4515 (N_4515,N_3597,N_3560);
xor U4516 (N_4516,N_3875,N_3182);
xor U4517 (N_4517,N_3754,N_3605);
or U4518 (N_4518,N_3203,N_3924);
xnor U4519 (N_4519,N_3480,N_3815);
or U4520 (N_4520,N_3327,N_3592);
nand U4521 (N_4521,N_3506,N_3314);
nand U4522 (N_4522,N_3762,N_3411);
or U4523 (N_4523,N_3187,N_3185);
nor U4524 (N_4524,N_3918,N_3731);
or U4525 (N_4525,N_3839,N_3961);
xor U4526 (N_4526,N_3553,N_3132);
and U4527 (N_4527,N_3807,N_3299);
nor U4528 (N_4528,N_3240,N_3629);
or U4529 (N_4529,N_3650,N_3002);
or U4530 (N_4530,N_3740,N_3628);
and U4531 (N_4531,N_3959,N_3562);
and U4532 (N_4532,N_3650,N_3360);
or U4533 (N_4533,N_3417,N_3451);
xor U4534 (N_4534,N_3231,N_3262);
xor U4535 (N_4535,N_3815,N_3392);
xor U4536 (N_4536,N_3126,N_3553);
and U4537 (N_4537,N_3965,N_3606);
nor U4538 (N_4538,N_3824,N_3739);
nand U4539 (N_4539,N_3379,N_3675);
nand U4540 (N_4540,N_3939,N_3520);
or U4541 (N_4541,N_3191,N_3347);
xor U4542 (N_4542,N_3388,N_3831);
nor U4543 (N_4543,N_3835,N_3296);
xnor U4544 (N_4544,N_3606,N_3882);
nand U4545 (N_4545,N_3390,N_3945);
nand U4546 (N_4546,N_3572,N_3223);
xnor U4547 (N_4547,N_3172,N_3591);
and U4548 (N_4548,N_3844,N_3496);
xnor U4549 (N_4549,N_3513,N_3076);
nor U4550 (N_4550,N_3046,N_3570);
nor U4551 (N_4551,N_3652,N_3725);
or U4552 (N_4552,N_3864,N_3848);
and U4553 (N_4553,N_3961,N_3067);
xnor U4554 (N_4554,N_3642,N_3420);
nand U4555 (N_4555,N_3641,N_3652);
nand U4556 (N_4556,N_3217,N_3742);
or U4557 (N_4557,N_3045,N_3619);
and U4558 (N_4558,N_3571,N_3498);
nand U4559 (N_4559,N_3862,N_3567);
or U4560 (N_4560,N_3130,N_3841);
nand U4561 (N_4561,N_3429,N_3679);
nand U4562 (N_4562,N_3465,N_3443);
nand U4563 (N_4563,N_3088,N_3453);
and U4564 (N_4564,N_3158,N_3202);
nand U4565 (N_4565,N_3422,N_3857);
nand U4566 (N_4566,N_3807,N_3518);
nand U4567 (N_4567,N_3425,N_3437);
nand U4568 (N_4568,N_3606,N_3058);
or U4569 (N_4569,N_3780,N_3609);
or U4570 (N_4570,N_3049,N_3545);
xor U4571 (N_4571,N_3583,N_3227);
and U4572 (N_4572,N_3446,N_3970);
nor U4573 (N_4573,N_3206,N_3417);
nand U4574 (N_4574,N_3458,N_3706);
and U4575 (N_4575,N_3286,N_3686);
or U4576 (N_4576,N_3346,N_3867);
and U4577 (N_4577,N_3310,N_3881);
nand U4578 (N_4578,N_3596,N_3948);
nand U4579 (N_4579,N_3414,N_3082);
nor U4580 (N_4580,N_3254,N_3821);
and U4581 (N_4581,N_3057,N_3992);
nor U4582 (N_4582,N_3099,N_3990);
xnor U4583 (N_4583,N_3278,N_3651);
nand U4584 (N_4584,N_3899,N_3513);
xnor U4585 (N_4585,N_3188,N_3336);
or U4586 (N_4586,N_3913,N_3987);
or U4587 (N_4587,N_3908,N_3705);
or U4588 (N_4588,N_3492,N_3334);
nor U4589 (N_4589,N_3049,N_3387);
or U4590 (N_4590,N_3522,N_3299);
and U4591 (N_4591,N_3200,N_3422);
or U4592 (N_4592,N_3376,N_3902);
nor U4593 (N_4593,N_3388,N_3818);
nor U4594 (N_4594,N_3842,N_3261);
nand U4595 (N_4595,N_3965,N_3959);
nand U4596 (N_4596,N_3335,N_3962);
nor U4597 (N_4597,N_3298,N_3047);
xnor U4598 (N_4598,N_3695,N_3771);
xor U4599 (N_4599,N_3555,N_3697);
or U4600 (N_4600,N_3420,N_3437);
and U4601 (N_4601,N_3607,N_3706);
or U4602 (N_4602,N_3041,N_3347);
and U4603 (N_4603,N_3603,N_3133);
and U4604 (N_4604,N_3579,N_3472);
xor U4605 (N_4605,N_3441,N_3671);
xor U4606 (N_4606,N_3966,N_3465);
xnor U4607 (N_4607,N_3933,N_3638);
or U4608 (N_4608,N_3683,N_3951);
and U4609 (N_4609,N_3466,N_3317);
and U4610 (N_4610,N_3593,N_3541);
or U4611 (N_4611,N_3280,N_3010);
or U4612 (N_4612,N_3233,N_3442);
xor U4613 (N_4613,N_3788,N_3963);
xnor U4614 (N_4614,N_3679,N_3393);
xnor U4615 (N_4615,N_3532,N_3595);
or U4616 (N_4616,N_3221,N_3077);
nor U4617 (N_4617,N_3532,N_3316);
or U4618 (N_4618,N_3896,N_3044);
or U4619 (N_4619,N_3327,N_3565);
xnor U4620 (N_4620,N_3926,N_3705);
nand U4621 (N_4621,N_3994,N_3243);
xor U4622 (N_4622,N_3552,N_3117);
nor U4623 (N_4623,N_3082,N_3629);
and U4624 (N_4624,N_3569,N_3633);
nor U4625 (N_4625,N_3694,N_3864);
nor U4626 (N_4626,N_3123,N_3667);
and U4627 (N_4627,N_3685,N_3652);
and U4628 (N_4628,N_3205,N_3383);
and U4629 (N_4629,N_3389,N_3744);
nor U4630 (N_4630,N_3526,N_3838);
nor U4631 (N_4631,N_3706,N_3757);
xor U4632 (N_4632,N_3852,N_3499);
nand U4633 (N_4633,N_3071,N_3203);
nor U4634 (N_4634,N_3289,N_3008);
xnor U4635 (N_4635,N_3246,N_3139);
or U4636 (N_4636,N_3714,N_3755);
and U4637 (N_4637,N_3144,N_3340);
or U4638 (N_4638,N_3406,N_3402);
xor U4639 (N_4639,N_3031,N_3028);
or U4640 (N_4640,N_3706,N_3834);
nor U4641 (N_4641,N_3392,N_3699);
or U4642 (N_4642,N_3008,N_3718);
or U4643 (N_4643,N_3859,N_3391);
nor U4644 (N_4644,N_3630,N_3274);
and U4645 (N_4645,N_3007,N_3624);
nand U4646 (N_4646,N_3851,N_3981);
xnor U4647 (N_4647,N_3619,N_3043);
nand U4648 (N_4648,N_3848,N_3922);
nor U4649 (N_4649,N_3627,N_3312);
or U4650 (N_4650,N_3719,N_3703);
xnor U4651 (N_4651,N_3074,N_3200);
xor U4652 (N_4652,N_3009,N_3298);
and U4653 (N_4653,N_3383,N_3852);
nand U4654 (N_4654,N_3607,N_3543);
nand U4655 (N_4655,N_3024,N_3531);
nand U4656 (N_4656,N_3993,N_3689);
and U4657 (N_4657,N_3759,N_3505);
nor U4658 (N_4658,N_3720,N_3946);
or U4659 (N_4659,N_3053,N_3384);
or U4660 (N_4660,N_3534,N_3928);
nand U4661 (N_4661,N_3110,N_3571);
xnor U4662 (N_4662,N_3873,N_3757);
nor U4663 (N_4663,N_3851,N_3319);
nand U4664 (N_4664,N_3031,N_3956);
nor U4665 (N_4665,N_3415,N_3994);
and U4666 (N_4666,N_3860,N_3252);
nand U4667 (N_4667,N_3350,N_3000);
nand U4668 (N_4668,N_3647,N_3339);
or U4669 (N_4669,N_3665,N_3510);
xor U4670 (N_4670,N_3644,N_3978);
or U4671 (N_4671,N_3919,N_3118);
xor U4672 (N_4672,N_3011,N_3581);
nor U4673 (N_4673,N_3177,N_3032);
xor U4674 (N_4674,N_3144,N_3224);
xor U4675 (N_4675,N_3561,N_3272);
nand U4676 (N_4676,N_3206,N_3703);
and U4677 (N_4677,N_3932,N_3265);
and U4678 (N_4678,N_3069,N_3729);
xor U4679 (N_4679,N_3979,N_3726);
xnor U4680 (N_4680,N_3004,N_3273);
or U4681 (N_4681,N_3976,N_3894);
and U4682 (N_4682,N_3524,N_3227);
or U4683 (N_4683,N_3166,N_3160);
or U4684 (N_4684,N_3054,N_3015);
or U4685 (N_4685,N_3562,N_3123);
xnor U4686 (N_4686,N_3109,N_3292);
nor U4687 (N_4687,N_3793,N_3999);
or U4688 (N_4688,N_3132,N_3960);
or U4689 (N_4689,N_3865,N_3282);
xor U4690 (N_4690,N_3745,N_3239);
nor U4691 (N_4691,N_3662,N_3901);
or U4692 (N_4692,N_3208,N_3567);
nand U4693 (N_4693,N_3690,N_3468);
nor U4694 (N_4694,N_3466,N_3809);
nand U4695 (N_4695,N_3612,N_3955);
or U4696 (N_4696,N_3858,N_3336);
nor U4697 (N_4697,N_3350,N_3129);
nand U4698 (N_4698,N_3478,N_3581);
xor U4699 (N_4699,N_3062,N_3414);
or U4700 (N_4700,N_3721,N_3333);
nand U4701 (N_4701,N_3509,N_3936);
nor U4702 (N_4702,N_3975,N_3454);
and U4703 (N_4703,N_3919,N_3628);
xor U4704 (N_4704,N_3329,N_3270);
xnor U4705 (N_4705,N_3825,N_3401);
nand U4706 (N_4706,N_3461,N_3146);
nor U4707 (N_4707,N_3359,N_3739);
nor U4708 (N_4708,N_3545,N_3331);
or U4709 (N_4709,N_3649,N_3631);
or U4710 (N_4710,N_3095,N_3321);
nor U4711 (N_4711,N_3552,N_3849);
xor U4712 (N_4712,N_3802,N_3992);
or U4713 (N_4713,N_3892,N_3502);
nand U4714 (N_4714,N_3422,N_3153);
nor U4715 (N_4715,N_3468,N_3667);
xnor U4716 (N_4716,N_3758,N_3169);
and U4717 (N_4717,N_3926,N_3774);
and U4718 (N_4718,N_3899,N_3465);
nor U4719 (N_4719,N_3103,N_3277);
or U4720 (N_4720,N_3244,N_3211);
nand U4721 (N_4721,N_3462,N_3529);
xor U4722 (N_4722,N_3712,N_3424);
and U4723 (N_4723,N_3218,N_3954);
nand U4724 (N_4724,N_3136,N_3990);
and U4725 (N_4725,N_3105,N_3261);
xor U4726 (N_4726,N_3813,N_3839);
nand U4727 (N_4727,N_3046,N_3236);
or U4728 (N_4728,N_3045,N_3621);
xnor U4729 (N_4729,N_3649,N_3394);
xor U4730 (N_4730,N_3210,N_3785);
nor U4731 (N_4731,N_3321,N_3117);
nand U4732 (N_4732,N_3871,N_3083);
and U4733 (N_4733,N_3376,N_3480);
xor U4734 (N_4734,N_3004,N_3410);
or U4735 (N_4735,N_3034,N_3360);
xnor U4736 (N_4736,N_3190,N_3922);
nand U4737 (N_4737,N_3597,N_3899);
nand U4738 (N_4738,N_3292,N_3409);
xnor U4739 (N_4739,N_3453,N_3763);
nand U4740 (N_4740,N_3651,N_3758);
or U4741 (N_4741,N_3455,N_3080);
or U4742 (N_4742,N_3403,N_3924);
nand U4743 (N_4743,N_3943,N_3668);
and U4744 (N_4744,N_3474,N_3178);
and U4745 (N_4745,N_3381,N_3151);
or U4746 (N_4746,N_3729,N_3115);
xnor U4747 (N_4747,N_3760,N_3635);
or U4748 (N_4748,N_3636,N_3426);
nor U4749 (N_4749,N_3742,N_3913);
xnor U4750 (N_4750,N_3001,N_3132);
xor U4751 (N_4751,N_3100,N_3153);
and U4752 (N_4752,N_3302,N_3931);
nand U4753 (N_4753,N_3973,N_3011);
nor U4754 (N_4754,N_3292,N_3684);
xor U4755 (N_4755,N_3382,N_3066);
and U4756 (N_4756,N_3462,N_3112);
nand U4757 (N_4757,N_3310,N_3778);
xor U4758 (N_4758,N_3401,N_3862);
nor U4759 (N_4759,N_3396,N_3228);
nand U4760 (N_4760,N_3542,N_3726);
and U4761 (N_4761,N_3213,N_3222);
and U4762 (N_4762,N_3152,N_3124);
and U4763 (N_4763,N_3890,N_3501);
nor U4764 (N_4764,N_3364,N_3620);
nand U4765 (N_4765,N_3744,N_3268);
nor U4766 (N_4766,N_3185,N_3470);
and U4767 (N_4767,N_3655,N_3071);
and U4768 (N_4768,N_3390,N_3642);
or U4769 (N_4769,N_3379,N_3175);
xnor U4770 (N_4770,N_3474,N_3489);
xor U4771 (N_4771,N_3040,N_3325);
and U4772 (N_4772,N_3015,N_3098);
nor U4773 (N_4773,N_3661,N_3473);
nand U4774 (N_4774,N_3866,N_3002);
nor U4775 (N_4775,N_3875,N_3136);
or U4776 (N_4776,N_3428,N_3745);
or U4777 (N_4777,N_3740,N_3779);
or U4778 (N_4778,N_3523,N_3743);
or U4779 (N_4779,N_3747,N_3920);
nor U4780 (N_4780,N_3696,N_3372);
or U4781 (N_4781,N_3961,N_3587);
nor U4782 (N_4782,N_3040,N_3354);
nor U4783 (N_4783,N_3820,N_3784);
xnor U4784 (N_4784,N_3680,N_3419);
nor U4785 (N_4785,N_3886,N_3085);
nor U4786 (N_4786,N_3410,N_3289);
nand U4787 (N_4787,N_3181,N_3296);
or U4788 (N_4788,N_3071,N_3348);
nor U4789 (N_4789,N_3022,N_3785);
and U4790 (N_4790,N_3601,N_3348);
nand U4791 (N_4791,N_3765,N_3878);
and U4792 (N_4792,N_3520,N_3706);
xnor U4793 (N_4793,N_3925,N_3592);
and U4794 (N_4794,N_3556,N_3215);
xor U4795 (N_4795,N_3963,N_3084);
nand U4796 (N_4796,N_3861,N_3885);
xnor U4797 (N_4797,N_3863,N_3962);
and U4798 (N_4798,N_3462,N_3942);
xnor U4799 (N_4799,N_3680,N_3433);
or U4800 (N_4800,N_3844,N_3996);
and U4801 (N_4801,N_3682,N_3089);
nor U4802 (N_4802,N_3619,N_3673);
and U4803 (N_4803,N_3944,N_3888);
nand U4804 (N_4804,N_3717,N_3622);
xnor U4805 (N_4805,N_3578,N_3956);
xnor U4806 (N_4806,N_3516,N_3215);
nor U4807 (N_4807,N_3737,N_3784);
nor U4808 (N_4808,N_3780,N_3098);
or U4809 (N_4809,N_3856,N_3267);
xor U4810 (N_4810,N_3747,N_3451);
xor U4811 (N_4811,N_3021,N_3936);
xnor U4812 (N_4812,N_3170,N_3609);
or U4813 (N_4813,N_3287,N_3117);
or U4814 (N_4814,N_3142,N_3660);
nor U4815 (N_4815,N_3217,N_3049);
nor U4816 (N_4816,N_3728,N_3809);
xnor U4817 (N_4817,N_3006,N_3660);
or U4818 (N_4818,N_3228,N_3173);
or U4819 (N_4819,N_3987,N_3513);
nor U4820 (N_4820,N_3333,N_3042);
xnor U4821 (N_4821,N_3958,N_3274);
xnor U4822 (N_4822,N_3351,N_3144);
xnor U4823 (N_4823,N_3569,N_3414);
nor U4824 (N_4824,N_3799,N_3866);
and U4825 (N_4825,N_3203,N_3190);
and U4826 (N_4826,N_3864,N_3361);
nor U4827 (N_4827,N_3425,N_3059);
nand U4828 (N_4828,N_3807,N_3990);
and U4829 (N_4829,N_3398,N_3117);
or U4830 (N_4830,N_3815,N_3449);
xnor U4831 (N_4831,N_3718,N_3828);
nor U4832 (N_4832,N_3312,N_3817);
nand U4833 (N_4833,N_3312,N_3078);
and U4834 (N_4834,N_3264,N_3765);
nand U4835 (N_4835,N_3096,N_3570);
nor U4836 (N_4836,N_3333,N_3110);
nand U4837 (N_4837,N_3307,N_3682);
nand U4838 (N_4838,N_3045,N_3061);
and U4839 (N_4839,N_3476,N_3993);
nor U4840 (N_4840,N_3360,N_3295);
and U4841 (N_4841,N_3249,N_3922);
or U4842 (N_4842,N_3103,N_3307);
and U4843 (N_4843,N_3745,N_3813);
xor U4844 (N_4844,N_3742,N_3594);
and U4845 (N_4845,N_3507,N_3026);
nor U4846 (N_4846,N_3203,N_3765);
nor U4847 (N_4847,N_3910,N_3479);
and U4848 (N_4848,N_3565,N_3189);
nor U4849 (N_4849,N_3299,N_3047);
or U4850 (N_4850,N_3544,N_3885);
and U4851 (N_4851,N_3310,N_3706);
or U4852 (N_4852,N_3881,N_3050);
xor U4853 (N_4853,N_3492,N_3267);
and U4854 (N_4854,N_3008,N_3431);
nand U4855 (N_4855,N_3608,N_3159);
nor U4856 (N_4856,N_3916,N_3650);
nor U4857 (N_4857,N_3375,N_3577);
nand U4858 (N_4858,N_3310,N_3429);
nand U4859 (N_4859,N_3961,N_3800);
nor U4860 (N_4860,N_3738,N_3729);
nor U4861 (N_4861,N_3233,N_3947);
nor U4862 (N_4862,N_3632,N_3876);
xnor U4863 (N_4863,N_3329,N_3582);
nor U4864 (N_4864,N_3233,N_3635);
nor U4865 (N_4865,N_3267,N_3634);
nand U4866 (N_4866,N_3044,N_3480);
and U4867 (N_4867,N_3736,N_3933);
nor U4868 (N_4868,N_3744,N_3628);
xnor U4869 (N_4869,N_3397,N_3903);
or U4870 (N_4870,N_3631,N_3588);
nor U4871 (N_4871,N_3427,N_3340);
xnor U4872 (N_4872,N_3935,N_3713);
and U4873 (N_4873,N_3881,N_3682);
xor U4874 (N_4874,N_3417,N_3562);
nor U4875 (N_4875,N_3978,N_3556);
nor U4876 (N_4876,N_3243,N_3465);
or U4877 (N_4877,N_3652,N_3565);
xnor U4878 (N_4878,N_3125,N_3323);
and U4879 (N_4879,N_3862,N_3376);
or U4880 (N_4880,N_3070,N_3369);
nand U4881 (N_4881,N_3129,N_3555);
nor U4882 (N_4882,N_3798,N_3476);
or U4883 (N_4883,N_3403,N_3708);
and U4884 (N_4884,N_3942,N_3631);
or U4885 (N_4885,N_3500,N_3147);
or U4886 (N_4886,N_3658,N_3894);
xor U4887 (N_4887,N_3130,N_3806);
or U4888 (N_4888,N_3513,N_3082);
nand U4889 (N_4889,N_3289,N_3786);
nor U4890 (N_4890,N_3927,N_3156);
and U4891 (N_4891,N_3158,N_3970);
nor U4892 (N_4892,N_3946,N_3670);
nor U4893 (N_4893,N_3493,N_3854);
and U4894 (N_4894,N_3460,N_3959);
nor U4895 (N_4895,N_3198,N_3825);
nand U4896 (N_4896,N_3913,N_3896);
nor U4897 (N_4897,N_3936,N_3834);
nand U4898 (N_4898,N_3491,N_3465);
and U4899 (N_4899,N_3810,N_3177);
nand U4900 (N_4900,N_3520,N_3629);
and U4901 (N_4901,N_3605,N_3099);
nor U4902 (N_4902,N_3624,N_3658);
nor U4903 (N_4903,N_3391,N_3642);
nand U4904 (N_4904,N_3855,N_3295);
xor U4905 (N_4905,N_3225,N_3454);
nor U4906 (N_4906,N_3412,N_3433);
or U4907 (N_4907,N_3333,N_3521);
xnor U4908 (N_4908,N_3328,N_3277);
nand U4909 (N_4909,N_3134,N_3815);
and U4910 (N_4910,N_3913,N_3420);
nor U4911 (N_4911,N_3325,N_3811);
or U4912 (N_4912,N_3609,N_3838);
nand U4913 (N_4913,N_3967,N_3656);
xor U4914 (N_4914,N_3310,N_3982);
and U4915 (N_4915,N_3269,N_3577);
or U4916 (N_4916,N_3583,N_3507);
or U4917 (N_4917,N_3510,N_3963);
nor U4918 (N_4918,N_3698,N_3476);
or U4919 (N_4919,N_3330,N_3408);
xnor U4920 (N_4920,N_3735,N_3973);
nand U4921 (N_4921,N_3077,N_3356);
nand U4922 (N_4922,N_3929,N_3935);
or U4923 (N_4923,N_3118,N_3241);
xnor U4924 (N_4924,N_3118,N_3855);
or U4925 (N_4925,N_3423,N_3369);
or U4926 (N_4926,N_3717,N_3399);
and U4927 (N_4927,N_3450,N_3615);
and U4928 (N_4928,N_3147,N_3244);
nor U4929 (N_4929,N_3751,N_3373);
nor U4930 (N_4930,N_3856,N_3366);
or U4931 (N_4931,N_3439,N_3049);
xnor U4932 (N_4932,N_3942,N_3525);
nand U4933 (N_4933,N_3562,N_3590);
nand U4934 (N_4934,N_3314,N_3159);
and U4935 (N_4935,N_3806,N_3812);
and U4936 (N_4936,N_3923,N_3966);
nor U4937 (N_4937,N_3700,N_3642);
xor U4938 (N_4938,N_3460,N_3119);
nand U4939 (N_4939,N_3863,N_3329);
nor U4940 (N_4940,N_3480,N_3026);
nor U4941 (N_4941,N_3450,N_3918);
xor U4942 (N_4942,N_3095,N_3918);
and U4943 (N_4943,N_3280,N_3669);
or U4944 (N_4944,N_3842,N_3888);
nand U4945 (N_4945,N_3421,N_3562);
and U4946 (N_4946,N_3566,N_3177);
and U4947 (N_4947,N_3935,N_3839);
xor U4948 (N_4948,N_3681,N_3130);
or U4949 (N_4949,N_3568,N_3660);
xor U4950 (N_4950,N_3788,N_3911);
or U4951 (N_4951,N_3873,N_3389);
nor U4952 (N_4952,N_3763,N_3995);
nor U4953 (N_4953,N_3991,N_3344);
nor U4954 (N_4954,N_3494,N_3381);
nor U4955 (N_4955,N_3017,N_3665);
nor U4956 (N_4956,N_3318,N_3493);
and U4957 (N_4957,N_3293,N_3170);
nor U4958 (N_4958,N_3873,N_3559);
or U4959 (N_4959,N_3119,N_3653);
xnor U4960 (N_4960,N_3802,N_3042);
nand U4961 (N_4961,N_3009,N_3677);
and U4962 (N_4962,N_3869,N_3436);
and U4963 (N_4963,N_3013,N_3853);
nand U4964 (N_4964,N_3962,N_3738);
or U4965 (N_4965,N_3148,N_3637);
xnor U4966 (N_4966,N_3633,N_3052);
nor U4967 (N_4967,N_3708,N_3642);
xor U4968 (N_4968,N_3622,N_3353);
nor U4969 (N_4969,N_3073,N_3319);
xnor U4970 (N_4970,N_3608,N_3370);
or U4971 (N_4971,N_3530,N_3912);
or U4972 (N_4972,N_3493,N_3843);
nand U4973 (N_4973,N_3017,N_3368);
nand U4974 (N_4974,N_3671,N_3694);
nand U4975 (N_4975,N_3481,N_3712);
xor U4976 (N_4976,N_3842,N_3927);
nand U4977 (N_4977,N_3473,N_3361);
or U4978 (N_4978,N_3284,N_3644);
and U4979 (N_4979,N_3127,N_3513);
and U4980 (N_4980,N_3556,N_3464);
xor U4981 (N_4981,N_3941,N_3795);
or U4982 (N_4982,N_3952,N_3979);
and U4983 (N_4983,N_3981,N_3951);
or U4984 (N_4984,N_3710,N_3680);
or U4985 (N_4985,N_3973,N_3728);
nand U4986 (N_4986,N_3383,N_3679);
nand U4987 (N_4987,N_3359,N_3442);
or U4988 (N_4988,N_3784,N_3201);
nand U4989 (N_4989,N_3346,N_3808);
nor U4990 (N_4990,N_3856,N_3473);
nand U4991 (N_4991,N_3091,N_3141);
xnor U4992 (N_4992,N_3866,N_3296);
or U4993 (N_4993,N_3937,N_3296);
and U4994 (N_4994,N_3389,N_3969);
or U4995 (N_4995,N_3819,N_3787);
xnor U4996 (N_4996,N_3516,N_3434);
or U4997 (N_4997,N_3555,N_3298);
xnor U4998 (N_4998,N_3769,N_3921);
xnor U4999 (N_4999,N_3383,N_3344);
xnor U5000 (N_5000,N_4831,N_4688);
nor U5001 (N_5001,N_4135,N_4145);
nand U5002 (N_5002,N_4327,N_4924);
nor U5003 (N_5003,N_4255,N_4848);
xor U5004 (N_5004,N_4596,N_4203);
xnor U5005 (N_5005,N_4572,N_4120);
nor U5006 (N_5006,N_4598,N_4983);
xnor U5007 (N_5007,N_4495,N_4721);
nor U5008 (N_5008,N_4579,N_4759);
xor U5009 (N_5009,N_4954,N_4814);
and U5010 (N_5010,N_4841,N_4535);
or U5011 (N_5011,N_4909,N_4289);
nand U5012 (N_5012,N_4534,N_4293);
xor U5013 (N_5013,N_4362,N_4118);
xnor U5014 (N_5014,N_4073,N_4714);
and U5015 (N_5015,N_4766,N_4067);
or U5016 (N_5016,N_4190,N_4687);
nor U5017 (N_5017,N_4873,N_4940);
nor U5018 (N_5018,N_4597,N_4884);
or U5019 (N_5019,N_4171,N_4728);
nor U5020 (N_5020,N_4013,N_4823);
xnor U5021 (N_5021,N_4585,N_4191);
and U5022 (N_5022,N_4715,N_4212);
nand U5023 (N_5023,N_4219,N_4718);
nor U5024 (N_5024,N_4244,N_4545);
xnor U5025 (N_5025,N_4961,N_4303);
and U5026 (N_5026,N_4665,N_4425);
nand U5027 (N_5027,N_4394,N_4007);
nand U5028 (N_5028,N_4151,N_4932);
nand U5029 (N_5029,N_4195,N_4971);
and U5030 (N_5030,N_4652,N_4836);
xor U5031 (N_5031,N_4215,N_4323);
nor U5032 (N_5032,N_4374,N_4678);
nor U5033 (N_5033,N_4328,N_4160);
and U5034 (N_5034,N_4381,N_4371);
or U5035 (N_5035,N_4207,N_4651);
or U5036 (N_5036,N_4764,N_4296);
nand U5037 (N_5037,N_4205,N_4737);
xor U5038 (N_5038,N_4262,N_4680);
xor U5039 (N_5039,N_4149,N_4908);
nand U5040 (N_5040,N_4438,N_4870);
nor U5041 (N_5041,N_4866,N_4096);
xnor U5042 (N_5042,N_4020,N_4294);
or U5043 (N_5043,N_4433,N_4268);
or U5044 (N_5044,N_4054,N_4837);
nand U5045 (N_5045,N_4918,N_4095);
nor U5046 (N_5046,N_4101,N_4887);
and U5047 (N_5047,N_4341,N_4157);
or U5048 (N_5048,N_4565,N_4454);
nand U5049 (N_5049,N_4318,N_4339);
and U5050 (N_5050,N_4566,N_4700);
and U5051 (N_5051,N_4458,N_4900);
xnor U5052 (N_5052,N_4933,N_4673);
xnor U5053 (N_5053,N_4635,N_4899);
or U5054 (N_5054,N_4740,N_4326);
nor U5055 (N_5055,N_4178,N_4209);
nand U5056 (N_5056,N_4478,N_4005);
and U5057 (N_5057,N_4291,N_4174);
nor U5058 (N_5058,N_4632,N_4970);
and U5059 (N_5059,N_4965,N_4320);
nand U5060 (N_5060,N_4379,N_4642);
nand U5061 (N_5061,N_4485,N_4507);
nor U5062 (N_5062,N_4310,N_4240);
and U5063 (N_5063,N_4769,N_4509);
xor U5064 (N_5064,N_4134,N_4351);
nor U5065 (N_5065,N_4391,N_4439);
and U5066 (N_5066,N_4524,N_4761);
nand U5067 (N_5067,N_4807,N_4563);
xor U5068 (N_5068,N_4414,N_4558);
and U5069 (N_5069,N_4313,N_4501);
and U5070 (N_5070,N_4650,N_4669);
xor U5071 (N_5071,N_4051,N_4756);
nor U5072 (N_5072,N_4466,N_4591);
nand U5073 (N_5073,N_4399,N_4859);
nor U5074 (N_5074,N_4206,N_4401);
xnor U5075 (N_5075,N_4959,N_4238);
and U5076 (N_5076,N_4987,N_4854);
xnor U5077 (N_5077,N_4931,N_4960);
nand U5078 (N_5078,N_4464,N_4008);
xnor U5079 (N_5079,N_4040,N_4239);
nand U5080 (N_5080,N_4516,N_4062);
or U5081 (N_5081,N_4861,N_4305);
xor U5082 (N_5082,N_4772,N_4702);
nand U5083 (N_5083,N_4985,N_4638);
nor U5084 (N_5084,N_4802,N_4066);
xor U5085 (N_5085,N_4281,N_4350);
or U5086 (N_5086,N_4974,N_4382);
or U5087 (N_5087,N_4139,N_4282);
xor U5088 (N_5088,N_4152,N_4417);
and U5089 (N_5089,N_4408,N_4457);
and U5090 (N_5090,N_4274,N_4886);
xnor U5091 (N_5091,N_4449,N_4666);
xor U5092 (N_5092,N_4016,N_4935);
nand U5093 (N_5093,N_4055,N_4595);
and U5094 (N_5094,N_4947,N_4763);
nor U5095 (N_5095,N_4813,N_4036);
nor U5096 (N_5096,N_4574,N_4695);
or U5097 (N_5097,N_4148,N_4405);
nor U5098 (N_5098,N_4684,N_4636);
xor U5099 (N_5099,N_4277,N_4169);
nand U5100 (N_5100,N_4435,N_4560);
xnor U5101 (N_5101,N_4132,N_4033);
xnor U5102 (N_5102,N_4301,N_4001);
nand U5103 (N_5103,N_4540,N_4470);
or U5104 (N_5104,N_4967,N_4283);
or U5105 (N_5105,N_4156,N_4874);
and U5106 (N_5106,N_4533,N_4634);
nand U5107 (N_5107,N_4388,N_4317);
nand U5108 (N_5108,N_4590,N_4307);
and U5109 (N_5109,N_4819,N_4779);
nand U5110 (N_5110,N_4617,N_4483);
nand U5111 (N_5111,N_4093,N_4757);
and U5112 (N_5112,N_4701,N_4821);
nor U5113 (N_5113,N_4245,N_4357);
xnor U5114 (N_5114,N_4928,N_4696);
xnor U5115 (N_5115,N_4229,N_4988);
and U5116 (N_5116,N_4549,N_4895);
xnor U5117 (N_5117,N_4847,N_4853);
xor U5118 (N_5118,N_4710,N_4923);
or U5119 (N_5119,N_4760,N_4712);
xor U5120 (N_5120,N_4913,N_4131);
xnor U5121 (N_5121,N_4775,N_4522);
xnor U5122 (N_5122,N_4415,N_4811);
nor U5123 (N_5123,N_4529,N_4493);
and U5124 (N_5124,N_4538,N_4746);
or U5125 (N_5125,N_4530,N_4074);
nand U5126 (N_5126,N_4739,N_4738);
and U5127 (N_5127,N_4264,N_4484);
and U5128 (N_5128,N_4898,N_4254);
and U5129 (N_5129,N_4795,N_4041);
nor U5130 (N_5130,N_4850,N_4612);
nor U5131 (N_5131,N_4794,N_4600);
nor U5132 (N_5132,N_4711,N_4774);
and U5133 (N_5133,N_4902,N_4044);
or U5134 (N_5134,N_4561,N_4496);
nand U5135 (N_5135,N_4112,N_4419);
and U5136 (N_5136,N_4885,N_4792);
or U5137 (N_5137,N_4311,N_4542);
xnor U5138 (N_5138,N_4511,N_4919);
xor U5139 (N_5139,N_4355,N_4882);
and U5140 (N_5140,N_4555,N_4499);
and U5141 (N_5141,N_4197,N_4842);
xnor U5142 (N_5142,N_4876,N_4372);
nand U5143 (N_5143,N_4707,N_4298);
or U5144 (N_5144,N_4083,N_4945);
nand U5145 (N_5145,N_4028,N_4914);
nor U5146 (N_5146,N_4984,N_4488);
xor U5147 (N_5147,N_4162,N_4778);
and U5148 (N_5148,N_4183,N_4697);
or U5149 (N_5149,N_4312,N_4990);
and U5150 (N_5150,N_4986,N_4646);
and U5151 (N_5151,N_4531,N_4981);
xor U5152 (N_5152,N_4604,N_4386);
nor U5153 (N_5153,N_4295,N_4510);
xor U5154 (N_5154,N_4235,N_4639);
xor U5155 (N_5155,N_4290,N_4490);
nor U5156 (N_5156,N_4825,N_4605);
xor U5157 (N_5157,N_4578,N_4336);
xor U5158 (N_5158,N_4855,N_4751);
or U5159 (N_5159,N_4453,N_4606);
xnor U5160 (N_5160,N_4237,N_4086);
and U5161 (N_5161,N_4471,N_4640);
and U5162 (N_5162,N_4809,N_4750);
nand U5163 (N_5163,N_4610,N_4552);
xnor U5164 (N_5164,N_4867,N_4691);
xor U5165 (N_5165,N_4690,N_4818);
nand U5166 (N_5166,N_4773,N_4342);
or U5167 (N_5167,N_4991,N_4042);
and U5168 (N_5168,N_4181,N_4300);
nor U5169 (N_5169,N_4359,N_4308);
nand U5170 (N_5170,N_4142,N_4503);
nand U5171 (N_5171,N_4445,N_4827);
and U5172 (N_5172,N_4315,N_4905);
xnor U5173 (N_5173,N_4890,N_4693);
nand U5174 (N_5174,N_4260,N_4978);
nand U5175 (N_5175,N_4976,N_4706);
nand U5176 (N_5176,N_4910,N_4917);
or U5177 (N_5177,N_4892,N_4121);
nor U5178 (N_5178,N_4647,N_4504);
xor U5179 (N_5179,N_4380,N_4888);
and U5180 (N_5180,N_4514,N_4060);
nor U5181 (N_5181,N_4285,N_4973);
or U5182 (N_5182,N_4431,N_4621);
nor U5183 (N_5183,N_4267,N_4799);
or U5184 (N_5184,N_4662,N_4340);
or U5185 (N_5185,N_4094,N_4223);
nand U5186 (N_5186,N_4951,N_4934);
nor U5187 (N_5187,N_4752,N_4172);
or U5188 (N_5188,N_4109,N_4498);
xor U5189 (N_5189,N_4589,N_4188);
nand U5190 (N_5190,N_4024,N_4029);
nor U5191 (N_5191,N_4929,N_4143);
nor U5192 (N_5192,N_4225,N_4879);
nand U5193 (N_5193,N_4655,N_4337);
xor U5194 (N_5194,N_4958,N_4955);
nand U5195 (N_5195,N_4626,N_4480);
xor U5196 (N_5196,N_4402,N_4039);
xor U5197 (N_5197,N_4309,N_4460);
nor U5198 (N_5198,N_4804,N_4852);
nor U5199 (N_5199,N_4835,N_4361);
xnor U5200 (N_5200,N_4059,N_4186);
and U5201 (N_5201,N_4602,N_4047);
or U5202 (N_5202,N_4037,N_4570);
xnor U5203 (N_5203,N_4213,N_4796);
nand U5204 (N_5204,N_4243,N_4941);
and U5205 (N_5205,N_4014,N_4754);
nor U5206 (N_5206,N_4742,N_4812);
nor U5207 (N_5207,N_4091,N_4168);
nand U5208 (N_5208,N_4137,N_4840);
nor U5209 (N_5209,N_4130,N_4393);
nand U5210 (N_5210,N_4576,N_4980);
nand U5211 (N_5211,N_4163,N_4649);
nand U5212 (N_5212,N_4364,N_4184);
nand U5213 (N_5213,N_4758,N_4006);
and U5214 (N_5214,N_4582,N_4127);
and U5215 (N_5215,N_4896,N_4170);
xnor U5216 (N_5216,N_4452,N_4226);
and U5217 (N_5217,N_4875,N_4833);
nor U5218 (N_5218,N_4878,N_4770);
xnor U5219 (N_5219,N_4079,N_4500);
nor U5220 (N_5220,N_4735,N_4858);
and U5221 (N_5221,N_4104,N_4801);
xnor U5222 (N_5222,N_4525,N_4674);
nand U5223 (N_5223,N_4658,N_4656);
nand U5224 (N_5224,N_4147,N_4584);
or U5225 (N_5225,N_4434,N_4894);
nor U5226 (N_5226,N_4231,N_4732);
xnor U5227 (N_5227,N_4546,N_4138);
or U5228 (N_5228,N_4851,N_4273);
xor U5229 (N_5229,N_4302,N_4200);
nand U5230 (N_5230,N_4999,N_4705);
nand U5231 (N_5231,N_4349,N_4553);
or U5232 (N_5232,N_4368,N_4257);
or U5233 (N_5233,N_4920,N_4099);
and U5234 (N_5234,N_4614,N_4193);
and U5235 (N_5235,N_4627,N_4429);
xor U5236 (N_5236,N_4571,N_4616);
nand U5237 (N_5237,N_4410,N_4734);
xnor U5238 (N_5238,N_4948,N_4862);
nor U5239 (N_5239,N_4249,N_4594);
nand U5240 (N_5240,N_4615,N_4263);
nand U5241 (N_5241,N_4520,N_4581);
or U5242 (N_5242,N_4620,N_4297);
xnor U5243 (N_5243,N_4411,N_4428);
nand U5244 (N_5244,N_4962,N_4915);
nand U5245 (N_5245,N_4564,N_4942);
xor U5246 (N_5246,N_4724,N_4664);
nor U5247 (N_5247,N_4343,N_4446);
nand U5248 (N_5248,N_4330,N_4443);
and U5249 (N_5249,N_4776,N_4292);
and U5250 (N_5250,N_4078,N_4893);
xnor U5251 (N_5251,N_4901,N_4528);
and U5252 (N_5252,N_4869,N_4663);
and U5253 (N_5253,N_4420,N_4106);
and U5254 (N_5254,N_4247,N_4881);
and U5255 (N_5255,N_4645,N_4345);
or U5256 (N_5256,N_4708,N_4822);
and U5257 (N_5257,N_4472,N_4783);
nor U5258 (N_5258,N_4385,N_4834);
or U5259 (N_5259,N_4068,N_4736);
nand U5260 (N_5260,N_4084,N_4221);
xnor U5261 (N_5261,N_4994,N_4883);
nand U5262 (N_5262,N_4119,N_4703);
xnor U5263 (N_5263,N_4473,N_4459);
or U5264 (N_5264,N_4196,N_4857);
nor U5265 (N_5265,N_4199,N_4583);
nor U5266 (N_5266,N_4465,N_4421);
nor U5267 (N_5267,N_4304,N_4335);
and U5268 (N_5268,N_4939,N_4166);
nand U5269 (N_5269,N_4798,N_4319);
nor U5270 (N_5270,N_4021,N_4234);
or U5271 (N_5271,N_4092,N_4442);
nand U5272 (N_5272,N_4768,N_4906);
or U5273 (N_5273,N_4032,N_4412);
nor U5274 (N_5274,N_4494,N_4177);
nand U5275 (N_5275,N_4116,N_4027);
xnor U5276 (N_5276,N_4603,N_4233);
nor U5277 (N_5277,N_4676,N_4100);
nor U5278 (N_5278,N_4586,N_4717);
xnor U5279 (N_5279,N_4912,N_4236);
nor U5280 (N_5280,N_4050,N_4916);
xnor U5281 (N_5281,N_4019,N_4220);
xor U5282 (N_5282,N_4911,N_4011);
nor U5283 (N_5283,N_4211,N_4747);
xnor U5284 (N_5284,N_4017,N_4124);
nand U5285 (N_5285,N_4159,N_4165);
and U5286 (N_5286,N_4187,N_4216);
nand U5287 (N_5287,N_4781,N_4679);
xor U5288 (N_5288,N_4550,N_4369);
or U5289 (N_5289,N_4176,N_4539);
xor U5290 (N_5290,N_4506,N_4749);
nand U5291 (N_5291,N_4481,N_4261);
and U5292 (N_5292,N_4424,N_4447);
xor U5293 (N_5293,N_4623,N_4926);
or U5294 (N_5294,N_4765,N_4963);
nor U5295 (N_5295,N_4956,N_4266);
and U5296 (N_5296,N_4720,N_4521);
or U5297 (N_5297,N_4444,N_4826);
nand U5298 (N_5298,N_4629,N_4618);
or U5299 (N_5299,N_4815,N_4643);
nand U5300 (N_5300,N_4133,N_4252);
nand U5301 (N_5301,N_4448,N_4657);
xor U5302 (N_5302,N_4085,N_4271);
and U5303 (N_5303,N_4670,N_4146);
nand U5304 (N_5304,N_4377,N_4845);
and U5305 (N_5305,N_4681,N_4248);
and U5306 (N_5306,N_4175,N_4568);
xnor U5307 (N_5307,N_4398,N_4719);
xor U5308 (N_5308,N_4150,N_4413);
and U5309 (N_5309,N_4167,N_4904);
and U5310 (N_5310,N_4921,N_4153);
xor U5311 (N_5311,N_4659,N_4727);
nand U5312 (N_5312,N_4000,N_4105);
and U5313 (N_5313,N_4416,N_4654);
and U5314 (N_5314,N_4993,N_4467);
or U5315 (N_5315,N_4440,N_4977);
nor U5316 (N_5316,N_4536,N_4155);
nand U5317 (N_5317,N_4547,N_4463);
nor U5318 (N_5318,N_4208,N_4569);
nand U5319 (N_5319,N_4709,N_4087);
xor U5320 (N_5320,N_4637,N_4002);
or U5321 (N_5321,N_4671,N_4076);
xnor U5322 (N_5322,N_4354,N_4276);
nand U5323 (N_5323,N_4513,N_4532);
and U5324 (N_5324,N_4198,N_4686);
or U5325 (N_5325,N_4998,N_4432);
or U5326 (N_5326,N_4406,N_4396);
nor U5327 (N_5327,N_4889,N_4026);
and U5328 (N_5328,N_4061,N_4562);
or U5329 (N_5329,N_4436,N_4048);
nor U5330 (N_5330,N_4389,N_4468);
and U5331 (N_5331,N_4577,N_4046);
xnor U5332 (N_5332,N_4515,N_4609);
and U5333 (N_5333,N_4284,N_4682);
and U5334 (N_5334,N_4789,N_4541);
xnor U5335 (N_5335,N_4730,N_4180);
and U5336 (N_5336,N_4593,N_4242);
and U5337 (N_5337,N_4324,N_4230);
or U5338 (N_5338,N_4097,N_4383);
or U5339 (N_5339,N_4025,N_4832);
nor U5340 (N_5340,N_4699,N_4788);
nor U5341 (N_5341,N_4949,N_4587);
xnor U5342 (N_5342,N_4451,N_4217);
nand U5343 (N_5343,N_4660,N_4376);
or U5344 (N_5344,N_4683,N_4075);
nand U5345 (N_5345,N_4018,N_4373);
xnor U5346 (N_5346,N_4573,N_4430);
xnor U5347 (N_5347,N_4334,N_4628);
nand U5348 (N_5348,N_4797,N_4793);
xor U5349 (N_5349,N_4052,N_4090);
nand U5350 (N_5350,N_4108,N_4519);
nor U5351 (N_5351,N_4755,N_4077);
or U5352 (N_5352,N_4810,N_4397);
or U5353 (N_5353,N_4868,N_4624);
and U5354 (N_5354,N_4404,N_4543);
nand U5355 (N_5355,N_4992,N_4856);
and U5356 (N_5356,N_4395,N_4489);
xnor U5357 (N_5357,N_4968,N_4316);
or U5358 (N_5358,N_4088,N_4009);
or U5359 (N_5359,N_4299,N_4744);
or U5360 (N_5360,N_4482,N_4456);
or U5361 (N_5361,N_4347,N_4422);
or U5362 (N_5362,N_4762,N_4390);
or U5363 (N_5363,N_4502,N_4601);
or U5364 (N_5364,N_4441,N_4677);
nand U5365 (N_5365,N_4479,N_4461);
or U5366 (N_5366,N_4592,N_4588);
nand U5367 (N_5367,N_4462,N_4863);
nor U5368 (N_5368,N_4551,N_4922);
and U5369 (N_5369,N_4829,N_4925);
nand U5370 (N_5370,N_4907,N_4930);
and U5371 (N_5371,N_4491,N_4497);
or U5372 (N_5372,N_4098,N_4426);
nor U5373 (N_5373,N_4250,N_4625);
xor U5374 (N_5374,N_4607,N_4232);
nor U5375 (N_5375,N_4224,N_4648);
nor U5376 (N_5376,N_4580,N_4611);
xor U5377 (N_5377,N_4338,N_4056);
or U5378 (N_5378,N_4204,N_4698);
or U5379 (N_5379,N_4003,N_4979);
and U5380 (N_5380,N_4314,N_4071);
xor U5381 (N_5381,N_4192,N_4475);
nor U5382 (N_5382,N_4838,N_4182);
xnor U5383 (N_5383,N_4222,N_4140);
or U5384 (N_5384,N_4556,N_4820);
xor U5385 (N_5385,N_4741,N_4731);
and U5386 (N_5386,N_4619,N_4816);
nand U5387 (N_5387,N_4070,N_4903);
nor U5388 (N_5388,N_4729,N_4950);
xnor U5389 (N_5389,N_4344,N_4784);
nand U5390 (N_5390,N_4817,N_4953);
or U5391 (N_5391,N_4806,N_4031);
and U5392 (N_5392,N_4034,N_4455);
or U5393 (N_5393,N_4716,N_4270);
and U5394 (N_5394,N_4554,N_4544);
or U5395 (N_5395,N_4871,N_4103);
or U5396 (N_5396,N_4946,N_4957);
xor U5397 (N_5397,N_4865,N_4672);
xnor U5398 (N_5398,N_4286,N_4228);
xnor U5399 (N_5399,N_4241,N_4129);
or U5400 (N_5400,N_4278,N_4189);
xnor U5401 (N_5401,N_4136,N_4653);
nor U5402 (N_5402,N_4423,N_4063);
xor U5403 (N_5403,N_4748,N_4015);
nor U5404 (N_5404,N_4306,N_4777);
and U5405 (N_5405,N_4830,N_4202);
nor U5406 (N_5406,N_4864,N_4358);
xor U5407 (N_5407,N_4370,N_4280);
and U5408 (N_5408,N_4661,N_4843);
and U5409 (N_5409,N_4325,N_4846);
or U5410 (N_5410,N_4474,N_4049);
xnor U5411 (N_5411,N_4427,N_4487);
nand U5412 (N_5412,N_4469,N_4780);
nand U5413 (N_5413,N_4123,N_4694);
nor U5414 (N_5414,N_4743,N_4072);
or U5415 (N_5415,N_4505,N_4733);
and U5416 (N_5416,N_4035,N_4476);
nand U5417 (N_5417,N_4575,N_4782);
or U5418 (N_5418,N_4321,N_4997);
xnor U5419 (N_5419,N_4353,N_4065);
and U5420 (N_5420,N_4348,N_4256);
nand U5421 (N_5421,N_4064,N_4057);
and U5422 (N_5422,N_4378,N_4844);
and U5423 (N_5423,N_4996,N_4808);
or U5424 (N_5424,N_4622,N_4689);
and U5425 (N_5425,N_4692,N_4403);
or U5426 (N_5426,N_4128,N_4275);
nand U5427 (N_5427,N_4322,N_4246);
xor U5428 (N_5428,N_4173,N_4392);
or U5429 (N_5429,N_4849,N_4407);
or U5430 (N_5430,N_4012,N_4966);
xor U5431 (N_5431,N_4214,N_4081);
or U5432 (N_5432,N_4030,N_4667);
or U5433 (N_5433,N_4251,N_4185);
nand U5434 (N_5434,N_4548,N_4644);
nand U5435 (N_5435,N_4989,N_4633);
xor U5436 (N_5436,N_4723,N_4872);
xor U5437 (N_5437,N_4144,N_4725);
or U5438 (N_5438,N_4082,N_4517);
nor U5439 (N_5439,N_4210,N_4080);
and U5440 (N_5440,N_4023,N_4279);
or U5441 (N_5441,N_4333,N_4786);
xnor U5442 (N_5442,N_4771,N_4253);
xor U5443 (N_5443,N_4010,N_4141);
nand U5444 (N_5444,N_4803,N_4559);
nor U5445 (N_5445,N_4179,N_4418);
or U5446 (N_5446,N_4069,N_4877);
nor U5447 (N_5447,N_4114,N_4567);
nand U5448 (N_5448,N_4384,N_4366);
nand U5449 (N_5449,N_4599,N_4258);
and U5450 (N_5450,N_4969,N_4437);
nor U5451 (N_5451,N_4964,N_4972);
xor U5452 (N_5452,N_4022,N_4363);
or U5453 (N_5453,N_4839,N_4492);
nand U5454 (N_5454,N_4880,N_4937);
nand U5455 (N_5455,N_4367,N_4194);
and U5456 (N_5456,N_4043,N_4089);
xor U5457 (N_5457,N_4356,N_4409);
nand U5458 (N_5458,N_4518,N_4995);
nand U5459 (N_5459,N_4346,N_4631);
and U5460 (N_5460,N_4523,N_4287);
or U5461 (N_5461,N_4053,N_4272);
and U5462 (N_5462,N_4800,N_4975);
xor U5463 (N_5463,N_4927,N_4508);
xnor U5464 (N_5464,N_4891,N_4477);
xnor U5465 (N_5465,N_4110,N_4938);
and U5466 (N_5466,N_4161,N_4360);
nor U5467 (N_5467,N_4126,N_4722);
and U5468 (N_5468,N_4753,N_4450);
nor U5469 (N_5469,N_4824,N_4745);
or U5470 (N_5470,N_4668,N_4952);
nand U5471 (N_5471,N_4537,N_4512);
or U5472 (N_5472,N_4164,N_4045);
xor U5473 (N_5473,N_4685,N_4288);
nand U5474 (N_5474,N_4630,N_4641);
nand U5475 (N_5475,N_4218,N_4608);
xor U5476 (N_5476,N_4944,N_4387);
nand U5477 (N_5477,N_4726,N_4943);
and U5478 (N_5478,N_4158,N_4375);
nor U5479 (N_5479,N_4982,N_4767);
nor U5480 (N_5480,N_4400,N_4004);
xnor U5481 (N_5481,N_4125,N_4613);
xor U5482 (N_5482,N_4365,N_4675);
nand U5483 (N_5483,N_4115,N_4936);
nand U5484 (N_5484,N_4704,N_4713);
and U5485 (N_5485,N_4828,N_4331);
nor U5486 (N_5486,N_4117,N_4201);
nand U5487 (N_5487,N_4269,N_4102);
and U5488 (N_5488,N_4557,N_4527);
or U5489 (N_5489,N_4329,N_4897);
xor U5490 (N_5490,N_4122,N_4332);
nand U5491 (N_5491,N_4526,N_4259);
xnor U5492 (N_5492,N_4227,N_4113);
or U5493 (N_5493,N_4787,N_4111);
or U5494 (N_5494,N_4038,N_4352);
and U5495 (N_5495,N_4860,N_4107);
or U5496 (N_5496,N_4805,N_4058);
nor U5497 (N_5497,N_4785,N_4791);
nand U5498 (N_5498,N_4265,N_4486);
xnor U5499 (N_5499,N_4154,N_4790);
or U5500 (N_5500,N_4582,N_4622);
and U5501 (N_5501,N_4414,N_4977);
or U5502 (N_5502,N_4775,N_4621);
nand U5503 (N_5503,N_4111,N_4620);
or U5504 (N_5504,N_4677,N_4986);
nand U5505 (N_5505,N_4766,N_4925);
nand U5506 (N_5506,N_4412,N_4964);
nand U5507 (N_5507,N_4169,N_4303);
nand U5508 (N_5508,N_4025,N_4150);
xnor U5509 (N_5509,N_4629,N_4308);
nor U5510 (N_5510,N_4974,N_4750);
or U5511 (N_5511,N_4534,N_4733);
or U5512 (N_5512,N_4148,N_4905);
or U5513 (N_5513,N_4050,N_4582);
xnor U5514 (N_5514,N_4045,N_4082);
nand U5515 (N_5515,N_4305,N_4595);
nor U5516 (N_5516,N_4365,N_4091);
or U5517 (N_5517,N_4797,N_4515);
nor U5518 (N_5518,N_4637,N_4523);
or U5519 (N_5519,N_4580,N_4817);
or U5520 (N_5520,N_4366,N_4712);
xnor U5521 (N_5521,N_4602,N_4743);
xor U5522 (N_5522,N_4606,N_4666);
nor U5523 (N_5523,N_4881,N_4026);
xnor U5524 (N_5524,N_4688,N_4696);
xnor U5525 (N_5525,N_4169,N_4062);
nand U5526 (N_5526,N_4070,N_4538);
and U5527 (N_5527,N_4963,N_4529);
xor U5528 (N_5528,N_4821,N_4842);
xnor U5529 (N_5529,N_4589,N_4386);
xnor U5530 (N_5530,N_4726,N_4956);
and U5531 (N_5531,N_4739,N_4105);
nor U5532 (N_5532,N_4796,N_4063);
xor U5533 (N_5533,N_4502,N_4125);
or U5534 (N_5534,N_4898,N_4588);
and U5535 (N_5535,N_4918,N_4826);
nor U5536 (N_5536,N_4387,N_4572);
xnor U5537 (N_5537,N_4549,N_4323);
nor U5538 (N_5538,N_4253,N_4072);
or U5539 (N_5539,N_4715,N_4863);
xnor U5540 (N_5540,N_4309,N_4870);
nor U5541 (N_5541,N_4508,N_4086);
or U5542 (N_5542,N_4359,N_4610);
nor U5543 (N_5543,N_4045,N_4243);
and U5544 (N_5544,N_4194,N_4176);
and U5545 (N_5545,N_4630,N_4973);
or U5546 (N_5546,N_4998,N_4695);
xnor U5547 (N_5547,N_4422,N_4267);
and U5548 (N_5548,N_4967,N_4598);
or U5549 (N_5549,N_4852,N_4373);
nand U5550 (N_5550,N_4147,N_4907);
and U5551 (N_5551,N_4484,N_4167);
xnor U5552 (N_5552,N_4977,N_4912);
nand U5553 (N_5553,N_4117,N_4664);
xor U5554 (N_5554,N_4280,N_4569);
nor U5555 (N_5555,N_4074,N_4733);
xor U5556 (N_5556,N_4689,N_4424);
xnor U5557 (N_5557,N_4425,N_4465);
or U5558 (N_5558,N_4135,N_4985);
xnor U5559 (N_5559,N_4523,N_4135);
or U5560 (N_5560,N_4480,N_4917);
or U5561 (N_5561,N_4602,N_4295);
xor U5562 (N_5562,N_4485,N_4375);
or U5563 (N_5563,N_4288,N_4064);
xor U5564 (N_5564,N_4501,N_4033);
or U5565 (N_5565,N_4642,N_4686);
xor U5566 (N_5566,N_4519,N_4312);
and U5567 (N_5567,N_4822,N_4369);
xor U5568 (N_5568,N_4523,N_4742);
and U5569 (N_5569,N_4496,N_4029);
nand U5570 (N_5570,N_4648,N_4709);
or U5571 (N_5571,N_4558,N_4329);
nor U5572 (N_5572,N_4095,N_4098);
or U5573 (N_5573,N_4111,N_4428);
or U5574 (N_5574,N_4191,N_4020);
and U5575 (N_5575,N_4149,N_4114);
xnor U5576 (N_5576,N_4248,N_4858);
or U5577 (N_5577,N_4163,N_4713);
nor U5578 (N_5578,N_4326,N_4666);
nand U5579 (N_5579,N_4999,N_4904);
xnor U5580 (N_5580,N_4196,N_4903);
or U5581 (N_5581,N_4252,N_4869);
nor U5582 (N_5582,N_4998,N_4230);
or U5583 (N_5583,N_4896,N_4587);
or U5584 (N_5584,N_4548,N_4173);
nor U5585 (N_5585,N_4523,N_4952);
nor U5586 (N_5586,N_4888,N_4294);
nor U5587 (N_5587,N_4305,N_4285);
nand U5588 (N_5588,N_4878,N_4917);
xnor U5589 (N_5589,N_4564,N_4672);
nor U5590 (N_5590,N_4329,N_4842);
xor U5591 (N_5591,N_4590,N_4106);
xnor U5592 (N_5592,N_4801,N_4577);
nor U5593 (N_5593,N_4204,N_4823);
or U5594 (N_5594,N_4842,N_4330);
xnor U5595 (N_5595,N_4131,N_4410);
nand U5596 (N_5596,N_4262,N_4647);
xor U5597 (N_5597,N_4866,N_4189);
nor U5598 (N_5598,N_4454,N_4232);
nor U5599 (N_5599,N_4220,N_4815);
and U5600 (N_5600,N_4178,N_4196);
or U5601 (N_5601,N_4246,N_4636);
nand U5602 (N_5602,N_4483,N_4794);
or U5603 (N_5603,N_4527,N_4903);
and U5604 (N_5604,N_4919,N_4658);
xnor U5605 (N_5605,N_4452,N_4446);
nor U5606 (N_5606,N_4326,N_4138);
and U5607 (N_5607,N_4117,N_4170);
xor U5608 (N_5608,N_4407,N_4162);
and U5609 (N_5609,N_4488,N_4952);
nand U5610 (N_5610,N_4029,N_4159);
nand U5611 (N_5611,N_4913,N_4931);
nand U5612 (N_5612,N_4859,N_4545);
xnor U5613 (N_5613,N_4400,N_4926);
nor U5614 (N_5614,N_4318,N_4716);
or U5615 (N_5615,N_4913,N_4581);
or U5616 (N_5616,N_4354,N_4202);
nor U5617 (N_5617,N_4028,N_4501);
or U5618 (N_5618,N_4008,N_4914);
nand U5619 (N_5619,N_4026,N_4951);
nor U5620 (N_5620,N_4345,N_4562);
or U5621 (N_5621,N_4476,N_4073);
nor U5622 (N_5622,N_4472,N_4214);
nor U5623 (N_5623,N_4877,N_4671);
nor U5624 (N_5624,N_4961,N_4879);
nor U5625 (N_5625,N_4048,N_4816);
and U5626 (N_5626,N_4743,N_4425);
or U5627 (N_5627,N_4901,N_4310);
and U5628 (N_5628,N_4611,N_4851);
nor U5629 (N_5629,N_4360,N_4405);
nor U5630 (N_5630,N_4267,N_4089);
and U5631 (N_5631,N_4347,N_4812);
nand U5632 (N_5632,N_4530,N_4088);
nor U5633 (N_5633,N_4953,N_4864);
nor U5634 (N_5634,N_4533,N_4853);
or U5635 (N_5635,N_4049,N_4529);
nand U5636 (N_5636,N_4003,N_4595);
xor U5637 (N_5637,N_4563,N_4152);
and U5638 (N_5638,N_4419,N_4360);
nor U5639 (N_5639,N_4936,N_4536);
or U5640 (N_5640,N_4727,N_4074);
or U5641 (N_5641,N_4589,N_4216);
or U5642 (N_5642,N_4619,N_4923);
nand U5643 (N_5643,N_4176,N_4617);
or U5644 (N_5644,N_4276,N_4931);
nand U5645 (N_5645,N_4964,N_4010);
nand U5646 (N_5646,N_4755,N_4328);
and U5647 (N_5647,N_4686,N_4422);
and U5648 (N_5648,N_4021,N_4367);
and U5649 (N_5649,N_4788,N_4805);
nor U5650 (N_5650,N_4633,N_4896);
nor U5651 (N_5651,N_4282,N_4332);
and U5652 (N_5652,N_4740,N_4271);
and U5653 (N_5653,N_4190,N_4115);
nor U5654 (N_5654,N_4781,N_4722);
and U5655 (N_5655,N_4773,N_4528);
nor U5656 (N_5656,N_4956,N_4931);
and U5657 (N_5657,N_4136,N_4145);
nor U5658 (N_5658,N_4721,N_4484);
xnor U5659 (N_5659,N_4867,N_4686);
nand U5660 (N_5660,N_4695,N_4802);
and U5661 (N_5661,N_4662,N_4553);
xnor U5662 (N_5662,N_4113,N_4383);
xor U5663 (N_5663,N_4934,N_4280);
nand U5664 (N_5664,N_4817,N_4234);
nand U5665 (N_5665,N_4094,N_4960);
xnor U5666 (N_5666,N_4767,N_4586);
nand U5667 (N_5667,N_4115,N_4620);
xnor U5668 (N_5668,N_4135,N_4405);
nor U5669 (N_5669,N_4135,N_4260);
nand U5670 (N_5670,N_4340,N_4577);
xor U5671 (N_5671,N_4919,N_4403);
xor U5672 (N_5672,N_4611,N_4324);
nand U5673 (N_5673,N_4376,N_4475);
and U5674 (N_5674,N_4747,N_4142);
or U5675 (N_5675,N_4744,N_4346);
nand U5676 (N_5676,N_4300,N_4846);
xnor U5677 (N_5677,N_4215,N_4591);
or U5678 (N_5678,N_4370,N_4391);
and U5679 (N_5679,N_4906,N_4102);
or U5680 (N_5680,N_4168,N_4194);
xnor U5681 (N_5681,N_4700,N_4476);
or U5682 (N_5682,N_4230,N_4534);
xnor U5683 (N_5683,N_4548,N_4345);
or U5684 (N_5684,N_4046,N_4526);
xor U5685 (N_5685,N_4595,N_4656);
or U5686 (N_5686,N_4572,N_4879);
nor U5687 (N_5687,N_4022,N_4617);
or U5688 (N_5688,N_4590,N_4005);
or U5689 (N_5689,N_4163,N_4131);
and U5690 (N_5690,N_4186,N_4392);
and U5691 (N_5691,N_4526,N_4230);
xor U5692 (N_5692,N_4898,N_4782);
xor U5693 (N_5693,N_4361,N_4627);
or U5694 (N_5694,N_4321,N_4137);
xor U5695 (N_5695,N_4424,N_4667);
nand U5696 (N_5696,N_4635,N_4797);
or U5697 (N_5697,N_4594,N_4271);
or U5698 (N_5698,N_4305,N_4988);
nand U5699 (N_5699,N_4377,N_4887);
nor U5700 (N_5700,N_4935,N_4405);
xor U5701 (N_5701,N_4542,N_4131);
xor U5702 (N_5702,N_4572,N_4295);
or U5703 (N_5703,N_4437,N_4492);
xor U5704 (N_5704,N_4706,N_4831);
nand U5705 (N_5705,N_4504,N_4528);
nand U5706 (N_5706,N_4591,N_4068);
xor U5707 (N_5707,N_4617,N_4263);
and U5708 (N_5708,N_4061,N_4270);
nor U5709 (N_5709,N_4032,N_4040);
nand U5710 (N_5710,N_4825,N_4760);
xnor U5711 (N_5711,N_4608,N_4715);
or U5712 (N_5712,N_4649,N_4996);
xnor U5713 (N_5713,N_4951,N_4353);
nand U5714 (N_5714,N_4785,N_4939);
xor U5715 (N_5715,N_4007,N_4502);
nand U5716 (N_5716,N_4528,N_4082);
or U5717 (N_5717,N_4895,N_4346);
nand U5718 (N_5718,N_4678,N_4864);
xor U5719 (N_5719,N_4529,N_4742);
or U5720 (N_5720,N_4796,N_4960);
and U5721 (N_5721,N_4440,N_4394);
and U5722 (N_5722,N_4166,N_4606);
nand U5723 (N_5723,N_4429,N_4704);
and U5724 (N_5724,N_4482,N_4305);
and U5725 (N_5725,N_4533,N_4769);
and U5726 (N_5726,N_4954,N_4349);
or U5727 (N_5727,N_4746,N_4160);
xor U5728 (N_5728,N_4117,N_4087);
nand U5729 (N_5729,N_4314,N_4263);
nand U5730 (N_5730,N_4028,N_4252);
xnor U5731 (N_5731,N_4302,N_4573);
nand U5732 (N_5732,N_4030,N_4216);
nor U5733 (N_5733,N_4194,N_4984);
nor U5734 (N_5734,N_4393,N_4837);
and U5735 (N_5735,N_4732,N_4667);
xnor U5736 (N_5736,N_4211,N_4688);
nand U5737 (N_5737,N_4496,N_4855);
and U5738 (N_5738,N_4293,N_4034);
xor U5739 (N_5739,N_4804,N_4566);
nor U5740 (N_5740,N_4425,N_4243);
nor U5741 (N_5741,N_4273,N_4754);
nand U5742 (N_5742,N_4439,N_4529);
and U5743 (N_5743,N_4097,N_4667);
nor U5744 (N_5744,N_4427,N_4588);
or U5745 (N_5745,N_4453,N_4341);
nor U5746 (N_5746,N_4467,N_4480);
or U5747 (N_5747,N_4669,N_4290);
nor U5748 (N_5748,N_4817,N_4131);
and U5749 (N_5749,N_4716,N_4222);
xnor U5750 (N_5750,N_4523,N_4113);
nand U5751 (N_5751,N_4609,N_4334);
nand U5752 (N_5752,N_4455,N_4480);
nand U5753 (N_5753,N_4835,N_4677);
nand U5754 (N_5754,N_4919,N_4724);
xnor U5755 (N_5755,N_4144,N_4909);
or U5756 (N_5756,N_4546,N_4863);
or U5757 (N_5757,N_4340,N_4545);
nor U5758 (N_5758,N_4548,N_4169);
and U5759 (N_5759,N_4962,N_4893);
and U5760 (N_5760,N_4149,N_4577);
nor U5761 (N_5761,N_4256,N_4998);
nor U5762 (N_5762,N_4406,N_4995);
and U5763 (N_5763,N_4734,N_4668);
or U5764 (N_5764,N_4370,N_4980);
nand U5765 (N_5765,N_4144,N_4507);
xor U5766 (N_5766,N_4273,N_4229);
xnor U5767 (N_5767,N_4783,N_4375);
xor U5768 (N_5768,N_4729,N_4758);
or U5769 (N_5769,N_4973,N_4320);
nand U5770 (N_5770,N_4602,N_4179);
nor U5771 (N_5771,N_4819,N_4074);
xnor U5772 (N_5772,N_4990,N_4189);
nand U5773 (N_5773,N_4709,N_4917);
xor U5774 (N_5774,N_4310,N_4587);
xor U5775 (N_5775,N_4913,N_4085);
nand U5776 (N_5776,N_4795,N_4182);
nor U5777 (N_5777,N_4249,N_4616);
and U5778 (N_5778,N_4843,N_4252);
or U5779 (N_5779,N_4147,N_4062);
or U5780 (N_5780,N_4174,N_4321);
nor U5781 (N_5781,N_4157,N_4459);
nor U5782 (N_5782,N_4295,N_4895);
or U5783 (N_5783,N_4003,N_4784);
or U5784 (N_5784,N_4765,N_4018);
and U5785 (N_5785,N_4062,N_4833);
xor U5786 (N_5786,N_4225,N_4041);
nand U5787 (N_5787,N_4169,N_4501);
nor U5788 (N_5788,N_4277,N_4347);
xnor U5789 (N_5789,N_4244,N_4834);
nand U5790 (N_5790,N_4592,N_4446);
nor U5791 (N_5791,N_4497,N_4612);
and U5792 (N_5792,N_4090,N_4077);
and U5793 (N_5793,N_4033,N_4554);
nor U5794 (N_5794,N_4375,N_4474);
nor U5795 (N_5795,N_4681,N_4887);
or U5796 (N_5796,N_4634,N_4791);
or U5797 (N_5797,N_4582,N_4993);
nand U5798 (N_5798,N_4051,N_4717);
or U5799 (N_5799,N_4984,N_4531);
or U5800 (N_5800,N_4266,N_4596);
nor U5801 (N_5801,N_4297,N_4117);
xnor U5802 (N_5802,N_4655,N_4876);
nor U5803 (N_5803,N_4692,N_4977);
nor U5804 (N_5804,N_4689,N_4346);
xnor U5805 (N_5805,N_4821,N_4278);
nor U5806 (N_5806,N_4283,N_4742);
nand U5807 (N_5807,N_4401,N_4590);
nand U5808 (N_5808,N_4283,N_4802);
and U5809 (N_5809,N_4777,N_4129);
and U5810 (N_5810,N_4971,N_4561);
and U5811 (N_5811,N_4801,N_4508);
and U5812 (N_5812,N_4171,N_4558);
or U5813 (N_5813,N_4482,N_4987);
xnor U5814 (N_5814,N_4728,N_4006);
or U5815 (N_5815,N_4612,N_4340);
nor U5816 (N_5816,N_4020,N_4515);
or U5817 (N_5817,N_4373,N_4420);
and U5818 (N_5818,N_4091,N_4842);
xnor U5819 (N_5819,N_4310,N_4198);
xnor U5820 (N_5820,N_4499,N_4463);
nor U5821 (N_5821,N_4426,N_4529);
xor U5822 (N_5822,N_4036,N_4590);
and U5823 (N_5823,N_4597,N_4462);
or U5824 (N_5824,N_4833,N_4798);
xor U5825 (N_5825,N_4166,N_4753);
xnor U5826 (N_5826,N_4942,N_4253);
nand U5827 (N_5827,N_4233,N_4761);
nor U5828 (N_5828,N_4363,N_4276);
nor U5829 (N_5829,N_4336,N_4870);
and U5830 (N_5830,N_4703,N_4860);
and U5831 (N_5831,N_4843,N_4162);
nor U5832 (N_5832,N_4352,N_4197);
and U5833 (N_5833,N_4918,N_4729);
or U5834 (N_5834,N_4802,N_4134);
or U5835 (N_5835,N_4434,N_4863);
and U5836 (N_5836,N_4506,N_4590);
nand U5837 (N_5837,N_4697,N_4973);
xor U5838 (N_5838,N_4621,N_4387);
or U5839 (N_5839,N_4287,N_4820);
xnor U5840 (N_5840,N_4471,N_4151);
and U5841 (N_5841,N_4515,N_4276);
xor U5842 (N_5842,N_4965,N_4978);
nor U5843 (N_5843,N_4879,N_4546);
and U5844 (N_5844,N_4715,N_4186);
nor U5845 (N_5845,N_4856,N_4115);
or U5846 (N_5846,N_4079,N_4159);
nor U5847 (N_5847,N_4913,N_4393);
nor U5848 (N_5848,N_4791,N_4478);
nand U5849 (N_5849,N_4179,N_4343);
nand U5850 (N_5850,N_4730,N_4380);
and U5851 (N_5851,N_4696,N_4071);
nor U5852 (N_5852,N_4974,N_4857);
and U5853 (N_5853,N_4949,N_4775);
xor U5854 (N_5854,N_4946,N_4096);
and U5855 (N_5855,N_4370,N_4288);
xnor U5856 (N_5856,N_4684,N_4053);
or U5857 (N_5857,N_4215,N_4621);
xor U5858 (N_5858,N_4446,N_4248);
nor U5859 (N_5859,N_4116,N_4827);
nand U5860 (N_5860,N_4179,N_4255);
and U5861 (N_5861,N_4440,N_4620);
nor U5862 (N_5862,N_4008,N_4661);
nand U5863 (N_5863,N_4287,N_4328);
nand U5864 (N_5864,N_4585,N_4918);
or U5865 (N_5865,N_4517,N_4914);
nor U5866 (N_5866,N_4765,N_4378);
nand U5867 (N_5867,N_4894,N_4409);
xnor U5868 (N_5868,N_4303,N_4826);
or U5869 (N_5869,N_4392,N_4740);
nand U5870 (N_5870,N_4609,N_4558);
nor U5871 (N_5871,N_4762,N_4313);
or U5872 (N_5872,N_4416,N_4130);
nand U5873 (N_5873,N_4516,N_4352);
xor U5874 (N_5874,N_4497,N_4245);
or U5875 (N_5875,N_4770,N_4884);
xor U5876 (N_5876,N_4323,N_4857);
xor U5877 (N_5877,N_4882,N_4947);
xnor U5878 (N_5878,N_4807,N_4710);
nand U5879 (N_5879,N_4396,N_4444);
xor U5880 (N_5880,N_4117,N_4576);
and U5881 (N_5881,N_4174,N_4920);
or U5882 (N_5882,N_4043,N_4732);
xnor U5883 (N_5883,N_4046,N_4525);
nand U5884 (N_5884,N_4790,N_4596);
nor U5885 (N_5885,N_4884,N_4148);
nor U5886 (N_5886,N_4587,N_4550);
nand U5887 (N_5887,N_4985,N_4463);
or U5888 (N_5888,N_4695,N_4518);
xor U5889 (N_5889,N_4737,N_4224);
nor U5890 (N_5890,N_4164,N_4506);
nor U5891 (N_5891,N_4832,N_4687);
xnor U5892 (N_5892,N_4594,N_4090);
and U5893 (N_5893,N_4805,N_4013);
or U5894 (N_5894,N_4509,N_4595);
nand U5895 (N_5895,N_4818,N_4284);
or U5896 (N_5896,N_4770,N_4576);
nor U5897 (N_5897,N_4743,N_4345);
nand U5898 (N_5898,N_4619,N_4067);
nor U5899 (N_5899,N_4207,N_4389);
xor U5900 (N_5900,N_4954,N_4326);
and U5901 (N_5901,N_4969,N_4104);
nor U5902 (N_5902,N_4781,N_4917);
nor U5903 (N_5903,N_4301,N_4962);
nor U5904 (N_5904,N_4525,N_4684);
or U5905 (N_5905,N_4369,N_4764);
or U5906 (N_5906,N_4023,N_4373);
and U5907 (N_5907,N_4907,N_4727);
nand U5908 (N_5908,N_4977,N_4422);
or U5909 (N_5909,N_4760,N_4845);
xor U5910 (N_5910,N_4884,N_4029);
or U5911 (N_5911,N_4483,N_4742);
and U5912 (N_5912,N_4936,N_4615);
xnor U5913 (N_5913,N_4972,N_4061);
or U5914 (N_5914,N_4876,N_4163);
or U5915 (N_5915,N_4791,N_4628);
and U5916 (N_5916,N_4818,N_4923);
or U5917 (N_5917,N_4254,N_4641);
nor U5918 (N_5918,N_4807,N_4178);
xor U5919 (N_5919,N_4592,N_4022);
nor U5920 (N_5920,N_4387,N_4826);
xor U5921 (N_5921,N_4861,N_4238);
nor U5922 (N_5922,N_4976,N_4055);
nor U5923 (N_5923,N_4203,N_4479);
nand U5924 (N_5924,N_4254,N_4943);
and U5925 (N_5925,N_4024,N_4385);
nand U5926 (N_5926,N_4626,N_4666);
or U5927 (N_5927,N_4349,N_4678);
or U5928 (N_5928,N_4715,N_4267);
nand U5929 (N_5929,N_4727,N_4408);
nor U5930 (N_5930,N_4957,N_4664);
or U5931 (N_5931,N_4099,N_4432);
or U5932 (N_5932,N_4278,N_4689);
or U5933 (N_5933,N_4451,N_4447);
nand U5934 (N_5934,N_4197,N_4928);
and U5935 (N_5935,N_4330,N_4284);
nand U5936 (N_5936,N_4458,N_4488);
nand U5937 (N_5937,N_4308,N_4803);
xnor U5938 (N_5938,N_4176,N_4129);
xnor U5939 (N_5939,N_4923,N_4917);
nand U5940 (N_5940,N_4479,N_4111);
nand U5941 (N_5941,N_4425,N_4045);
nor U5942 (N_5942,N_4206,N_4689);
or U5943 (N_5943,N_4852,N_4854);
nor U5944 (N_5944,N_4236,N_4454);
nand U5945 (N_5945,N_4605,N_4573);
nor U5946 (N_5946,N_4362,N_4551);
nor U5947 (N_5947,N_4587,N_4177);
or U5948 (N_5948,N_4784,N_4490);
nand U5949 (N_5949,N_4744,N_4704);
or U5950 (N_5950,N_4309,N_4663);
xor U5951 (N_5951,N_4257,N_4500);
xor U5952 (N_5952,N_4833,N_4212);
xor U5953 (N_5953,N_4002,N_4834);
xnor U5954 (N_5954,N_4037,N_4207);
and U5955 (N_5955,N_4001,N_4075);
and U5956 (N_5956,N_4571,N_4959);
and U5957 (N_5957,N_4609,N_4418);
and U5958 (N_5958,N_4699,N_4403);
nand U5959 (N_5959,N_4462,N_4443);
nand U5960 (N_5960,N_4617,N_4659);
nand U5961 (N_5961,N_4697,N_4254);
or U5962 (N_5962,N_4074,N_4221);
nand U5963 (N_5963,N_4051,N_4099);
or U5964 (N_5964,N_4030,N_4075);
nor U5965 (N_5965,N_4970,N_4383);
nand U5966 (N_5966,N_4979,N_4858);
and U5967 (N_5967,N_4159,N_4038);
nor U5968 (N_5968,N_4928,N_4386);
or U5969 (N_5969,N_4343,N_4029);
and U5970 (N_5970,N_4314,N_4506);
and U5971 (N_5971,N_4972,N_4128);
xnor U5972 (N_5972,N_4158,N_4516);
nand U5973 (N_5973,N_4473,N_4712);
and U5974 (N_5974,N_4039,N_4501);
or U5975 (N_5975,N_4323,N_4018);
or U5976 (N_5976,N_4707,N_4505);
nor U5977 (N_5977,N_4825,N_4955);
nor U5978 (N_5978,N_4135,N_4942);
nand U5979 (N_5979,N_4254,N_4397);
xor U5980 (N_5980,N_4955,N_4930);
nand U5981 (N_5981,N_4291,N_4452);
nand U5982 (N_5982,N_4014,N_4349);
nand U5983 (N_5983,N_4157,N_4915);
or U5984 (N_5984,N_4756,N_4116);
xnor U5985 (N_5985,N_4858,N_4786);
nand U5986 (N_5986,N_4807,N_4093);
xnor U5987 (N_5987,N_4661,N_4935);
or U5988 (N_5988,N_4333,N_4930);
xor U5989 (N_5989,N_4109,N_4437);
and U5990 (N_5990,N_4769,N_4897);
or U5991 (N_5991,N_4864,N_4599);
xnor U5992 (N_5992,N_4186,N_4504);
nand U5993 (N_5993,N_4424,N_4184);
and U5994 (N_5994,N_4362,N_4530);
nand U5995 (N_5995,N_4461,N_4287);
nor U5996 (N_5996,N_4982,N_4812);
nand U5997 (N_5997,N_4077,N_4093);
nor U5998 (N_5998,N_4616,N_4880);
nor U5999 (N_5999,N_4407,N_4086);
nand U6000 (N_6000,N_5829,N_5888);
or U6001 (N_6001,N_5167,N_5385);
nor U6002 (N_6002,N_5961,N_5636);
nand U6003 (N_6003,N_5699,N_5431);
and U6004 (N_6004,N_5819,N_5512);
or U6005 (N_6005,N_5274,N_5973);
and U6006 (N_6006,N_5059,N_5152);
and U6007 (N_6007,N_5579,N_5088);
and U6008 (N_6008,N_5519,N_5017);
and U6009 (N_6009,N_5104,N_5214);
and U6010 (N_6010,N_5120,N_5731);
nand U6011 (N_6011,N_5720,N_5365);
nor U6012 (N_6012,N_5601,N_5500);
and U6013 (N_6013,N_5798,N_5107);
and U6014 (N_6014,N_5738,N_5140);
nand U6015 (N_6015,N_5981,N_5785);
nand U6016 (N_6016,N_5681,N_5090);
and U6017 (N_6017,N_5928,N_5462);
xnor U6018 (N_6018,N_5389,N_5861);
nand U6019 (N_6019,N_5988,N_5710);
and U6020 (N_6020,N_5357,N_5799);
or U6021 (N_6021,N_5038,N_5895);
nor U6022 (N_6022,N_5644,N_5989);
or U6023 (N_6023,N_5976,N_5905);
xnor U6024 (N_6024,N_5933,N_5084);
or U6025 (N_6025,N_5269,N_5061);
and U6026 (N_6026,N_5493,N_5438);
and U6027 (N_6027,N_5805,N_5137);
xnor U6028 (N_6028,N_5008,N_5787);
nor U6029 (N_6029,N_5974,N_5396);
or U6030 (N_6030,N_5985,N_5771);
nor U6031 (N_6031,N_5245,N_5891);
xor U6032 (N_6032,N_5547,N_5917);
nand U6033 (N_6033,N_5643,N_5066);
or U6034 (N_6034,N_5565,N_5237);
or U6035 (N_6035,N_5837,N_5412);
or U6036 (N_6036,N_5574,N_5662);
xor U6037 (N_6037,N_5646,N_5005);
nand U6038 (N_6038,N_5630,N_5401);
or U6039 (N_6039,N_5901,N_5658);
nor U6040 (N_6040,N_5388,N_5912);
xnor U6041 (N_6041,N_5424,N_5511);
nand U6042 (N_6042,N_5170,N_5617);
nand U6043 (N_6043,N_5822,N_5853);
xnor U6044 (N_6044,N_5289,N_5468);
nor U6045 (N_6045,N_5158,N_5344);
or U6046 (N_6046,N_5508,N_5845);
nand U6047 (N_6047,N_5536,N_5362);
nor U6048 (N_6048,N_5629,N_5095);
nand U6049 (N_6049,N_5665,N_5437);
xor U6050 (N_6050,N_5725,N_5218);
nor U6051 (N_6051,N_5654,N_5071);
and U6052 (N_6052,N_5467,N_5619);
nand U6053 (N_6053,N_5782,N_5872);
nor U6054 (N_6054,N_5865,N_5201);
nand U6055 (N_6055,N_5373,N_5524);
nand U6056 (N_6056,N_5919,N_5906);
nor U6057 (N_6057,N_5937,N_5454);
and U6058 (N_6058,N_5674,N_5657);
or U6059 (N_6059,N_5265,N_5585);
and U6060 (N_6060,N_5719,N_5859);
nand U6061 (N_6061,N_5982,N_5676);
xor U6062 (N_6062,N_5094,N_5737);
nand U6063 (N_6063,N_5768,N_5656);
nand U6064 (N_6064,N_5130,N_5145);
or U6065 (N_6065,N_5439,N_5247);
and U6066 (N_6066,N_5180,N_5118);
nor U6067 (N_6067,N_5641,N_5234);
and U6068 (N_6068,N_5922,N_5826);
xnor U6069 (N_6069,N_5063,N_5885);
nor U6070 (N_6070,N_5211,N_5416);
nor U6071 (N_6071,N_5293,N_5904);
nor U6072 (N_6072,N_5195,N_5591);
xnor U6073 (N_6073,N_5196,N_5542);
nand U6074 (N_6074,N_5428,N_5212);
nand U6075 (N_6075,N_5587,N_5345);
or U6076 (N_6076,N_5242,N_5332);
xnor U6077 (N_6077,N_5229,N_5956);
nand U6078 (N_6078,N_5726,N_5238);
or U6079 (N_6079,N_5372,N_5831);
nand U6080 (N_6080,N_5984,N_5839);
or U6081 (N_6081,N_5426,N_5767);
nand U6082 (N_6082,N_5138,N_5313);
or U6083 (N_6083,N_5147,N_5484);
nor U6084 (N_6084,N_5049,N_5376);
xnor U6085 (N_6085,N_5998,N_5934);
xnor U6086 (N_6086,N_5207,N_5325);
and U6087 (N_6087,N_5036,N_5114);
xor U6088 (N_6088,N_5341,N_5625);
or U6089 (N_6089,N_5999,N_5696);
and U6090 (N_6090,N_5480,N_5323);
nand U6091 (N_6091,N_5046,N_5635);
or U6092 (N_6092,N_5628,N_5442);
xor U6093 (N_6093,N_5538,N_5133);
xor U6094 (N_6094,N_5487,N_5550);
and U6095 (N_6095,N_5975,N_5679);
and U6096 (N_6096,N_5503,N_5203);
xor U6097 (N_6097,N_5276,N_5057);
and U6098 (N_6098,N_5441,N_5987);
xnor U6099 (N_6099,N_5686,N_5391);
nand U6100 (N_6100,N_5097,N_5384);
or U6101 (N_6101,N_5425,N_5564);
nand U6102 (N_6102,N_5667,N_5887);
or U6103 (N_6103,N_5947,N_5551);
or U6104 (N_6104,N_5606,N_5666);
xor U6105 (N_6105,N_5744,N_5330);
and U6106 (N_6106,N_5404,N_5303);
or U6107 (N_6107,N_5312,N_5406);
nor U6108 (N_6108,N_5306,N_5706);
xor U6109 (N_6109,N_5759,N_5777);
and U6110 (N_6110,N_5556,N_5966);
and U6111 (N_6111,N_5205,N_5714);
xnor U6112 (N_6112,N_5364,N_5563);
and U6113 (N_6113,N_5224,N_5623);
nand U6114 (N_6114,N_5311,N_5490);
nor U6115 (N_6115,N_5148,N_5308);
or U6116 (N_6116,N_5285,N_5582);
xnor U6117 (N_6117,N_5459,N_5978);
and U6118 (N_6118,N_5335,N_5117);
nor U6119 (N_6119,N_5031,N_5350);
and U6120 (N_6120,N_5680,N_5788);
or U6121 (N_6121,N_5271,N_5294);
nor U6122 (N_6122,N_5047,N_5122);
and U6123 (N_6123,N_5754,N_5669);
and U6124 (N_6124,N_5422,N_5716);
nor U6125 (N_6125,N_5011,N_5724);
or U6126 (N_6126,N_5544,N_5275);
and U6127 (N_6127,N_5451,N_5883);
nand U6128 (N_6128,N_5263,N_5692);
xor U6129 (N_6129,N_5227,N_5817);
nand U6130 (N_6130,N_5370,N_5160);
nor U6131 (N_6131,N_5394,N_5222);
nand U6132 (N_6132,N_5597,N_5778);
or U6133 (N_6133,N_5295,N_5125);
nand U6134 (N_6134,N_5832,N_5260);
nor U6135 (N_6135,N_5183,N_5034);
and U6136 (N_6136,N_5115,N_5820);
xnor U6137 (N_6137,N_5334,N_5486);
nor U6138 (N_6138,N_5081,N_5175);
or U6139 (N_6139,N_5127,N_5535);
nand U6140 (N_6140,N_5360,N_5124);
nor U6141 (N_6141,N_5419,N_5021);
xnor U6142 (N_6142,N_5531,N_5509);
and U6143 (N_6143,N_5268,N_5809);
or U6144 (N_6144,N_5675,N_5594);
and U6145 (N_6145,N_5811,N_5695);
nand U6146 (N_6146,N_5387,N_5721);
xnor U6147 (N_6147,N_5033,N_5185);
and U6148 (N_6148,N_5326,N_5056);
nor U6149 (N_6149,N_5233,N_5504);
or U6150 (N_6150,N_5445,N_5627);
and U6151 (N_6151,N_5995,N_5209);
xnor U6152 (N_6152,N_5116,N_5371);
or U6153 (N_6153,N_5403,N_5583);
xor U6154 (N_6154,N_5497,N_5640);
nand U6155 (N_6155,N_5801,N_5070);
or U6156 (N_6156,N_5996,N_5913);
or U6157 (N_6157,N_5942,N_5164);
nor U6158 (N_6158,N_5959,N_5123);
xnor U6159 (N_6159,N_5383,N_5397);
and U6160 (N_6160,N_5010,N_5022);
or U6161 (N_6161,N_5409,N_5476);
nand U6162 (N_6162,N_5882,N_5483);
nor U6163 (N_6163,N_5316,N_5711);
and U6164 (N_6164,N_5427,N_5291);
or U6165 (N_6165,N_5050,N_5566);
and U6166 (N_6166,N_5664,N_5529);
nand U6167 (N_6167,N_5267,N_5073);
nand U6168 (N_6168,N_5800,N_5044);
xor U6169 (N_6169,N_5348,N_5660);
and U6170 (N_6170,N_5226,N_5089);
and U6171 (N_6171,N_5062,N_5739);
nor U6172 (N_6172,N_5054,N_5743);
nand U6173 (N_6173,N_5890,N_5834);
and U6174 (N_6174,N_5053,N_5889);
xnor U6175 (N_6175,N_5277,N_5712);
or U6176 (N_6176,N_5361,N_5161);
or U6177 (N_6177,N_5604,N_5560);
nand U6178 (N_6178,N_5596,N_5390);
or U6179 (N_6179,N_5408,N_5842);
xnor U6180 (N_6180,N_5634,N_5900);
nand U6181 (N_6181,N_5707,N_5150);
nand U6182 (N_6182,N_5908,N_5301);
nand U6183 (N_6183,N_5398,N_5824);
nor U6184 (N_6184,N_5399,N_5518);
nor U6185 (N_6185,N_5897,N_5402);
xnor U6186 (N_6186,N_5825,N_5704);
nor U6187 (N_6187,N_5366,N_5249);
nand U6188 (N_6188,N_5894,N_5747);
nand U6189 (N_6189,N_5093,N_5953);
nor U6190 (N_6190,N_5239,N_5698);
nor U6191 (N_6191,N_5331,N_5027);
nor U6192 (N_6192,N_5177,N_5455);
or U6193 (N_6193,N_5156,N_5159);
nor U6194 (N_6194,N_5405,N_5553);
and U6195 (N_6195,N_5914,N_5297);
xnor U6196 (N_6196,N_5697,N_5460);
and U6197 (N_6197,N_5807,N_5279);
or U6198 (N_6198,N_5015,N_5045);
or U6199 (N_6199,N_5652,N_5983);
or U6200 (N_6200,N_5163,N_5713);
xor U6201 (N_6201,N_5270,N_5653);
nand U6202 (N_6202,N_5557,N_5622);
nor U6203 (N_6203,N_5283,N_5745);
xor U6204 (N_6204,N_5085,N_5307);
xor U6205 (N_6205,N_5962,N_5000);
or U6206 (N_6206,N_5154,N_5317);
nor U6207 (N_6207,N_5990,N_5593);
nand U6208 (N_6208,N_5902,N_5337);
or U6209 (N_6209,N_5333,N_5172);
nand U6210 (N_6210,N_5735,N_5608);
or U6211 (N_6211,N_5588,N_5346);
or U6212 (N_6212,N_5816,N_5621);
and U6213 (N_6213,N_5144,N_5936);
nor U6214 (N_6214,N_5539,N_5789);
or U6215 (N_6215,N_5082,N_5461);
nor U6216 (N_6216,N_5775,N_5432);
and U6217 (N_6217,N_5753,N_5616);
nand U6218 (N_6218,N_5377,N_5136);
xnor U6219 (N_6219,N_5932,N_5048);
and U6220 (N_6220,N_5794,N_5857);
and U6221 (N_6221,N_5868,N_5411);
nor U6222 (N_6222,N_5190,N_5258);
nor U6223 (N_6223,N_5494,N_5077);
or U6224 (N_6224,N_5722,N_5573);
nand U6225 (N_6225,N_5304,N_5952);
and U6226 (N_6226,N_5192,N_5182);
and U6227 (N_6227,N_5727,N_5429);
xnor U6228 (N_6228,N_5482,N_5613);
xor U6229 (N_6229,N_5446,N_5687);
xor U6230 (N_6230,N_5491,N_5705);
and U6231 (N_6231,N_5873,N_5068);
nand U6232 (N_6232,N_5945,N_5702);
and U6233 (N_6233,N_5328,N_5909);
or U6234 (N_6234,N_5272,N_5336);
nor U6235 (N_6235,N_5911,N_5774);
nor U6236 (N_6236,N_5729,N_5951);
or U6237 (N_6237,N_5142,N_5450);
xnor U6238 (N_6238,N_5296,N_5521);
and U6239 (N_6239,N_5578,N_5452);
and U6240 (N_6240,N_5067,N_5064);
nor U6241 (N_6241,N_5139,N_5670);
or U6242 (N_6242,N_5540,N_5434);
and U6243 (N_6243,N_5228,N_5112);
nor U6244 (N_6244,N_5079,N_5991);
nand U6245 (N_6245,N_5478,N_5691);
or U6246 (N_6246,N_5121,N_5375);
nor U6247 (N_6247,N_5471,N_5080);
nor U6248 (N_6248,N_5760,N_5672);
nand U6249 (N_6249,N_5523,N_5633);
nand U6250 (N_6250,N_5684,N_5166);
nor U6251 (N_6251,N_5925,N_5580);
xor U6252 (N_6252,N_5605,N_5786);
nand U6253 (N_6253,N_5693,N_5571);
or U6254 (N_6254,N_5287,N_5752);
nor U6255 (N_6255,N_5251,N_5457);
and U6256 (N_6256,N_5614,N_5174);
nor U6257 (N_6257,N_5252,N_5244);
or U6258 (N_6258,N_5972,N_5612);
and U6259 (N_6259,N_5510,N_5410);
nand U6260 (N_6260,N_5321,N_5162);
nor U6261 (N_6261,N_5230,N_5213);
nor U6262 (N_6262,N_5862,N_5165);
nor U6263 (N_6263,N_5382,N_5200);
nand U6264 (N_6264,N_5732,N_5610);
xor U6265 (N_6265,N_5943,N_5818);
nand U6266 (N_6266,N_5474,N_5892);
or U6267 (N_6267,N_5899,N_5266);
nand U6268 (N_6268,N_5042,N_5264);
nor U6269 (N_6269,N_5576,N_5866);
xnor U6270 (N_6270,N_5530,N_5701);
nand U6271 (N_6271,N_5948,N_5023);
nor U6272 (N_6272,N_5545,N_5241);
nand U6273 (N_6273,N_5717,N_5682);
nor U6274 (N_6274,N_5528,N_5537);
nand U6275 (N_6275,N_5004,N_5083);
and U6276 (N_6276,N_5052,N_5099);
nand U6277 (N_6277,N_5111,N_5813);
or U6278 (N_6278,N_5694,N_5690);
and U6279 (N_6279,N_5965,N_5481);
xor U6280 (N_6280,N_5035,N_5920);
nor U6281 (N_6281,N_5864,N_5028);
and U6282 (N_6282,N_5880,N_5135);
and U6283 (N_6283,N_5647,N_5359);
xor U6284 (N_6284,N_5569,N_5969);
and U6285 (N_6285,N_5874,N_5299);
xnor U6286 (N_6286,N_5584,N_5178);
nor U6287 (N_6287,N_5197,N_5848);
and U6288 (N_6288,N_5844,N_5761);
nand U6289 (N_6289,N_5802,N_5639);
nor U6290 (N_6290,N_5992,N_5562);
xor U6291 (N_6291,N_5146,N_5931);
nor U6292 (N_6292,N_5828,N_5907);
nor U6293 (N_6293,N_5833,N_5558);
nand U6294 (N_6294,N_5255,N_5709);
xor U6295 (N_6295,N_5319,N_5339);
and U6296 (N_6296,N_5860,N_5219);
or U6297 (N_6297,N_5413,N_5740);
nand U6298 (N_6298,N_5513,N_5273);
nand U6299 (N_6299,N_5688,N_5204);
and U6300 (N_6300,N_5967,N_5448);
nand U6301 (N_6301,N_5821,N_5921);
xor U6302 (N_6302,N_5443,N_5659);
or U6303 (N_6303,N_5168,N_5058);
nor U6304 (N_6304,N_5220,N_5003);
or U6305 (N_6305,N_5827,N_5193);
xnor U6306 (N_6306,N_5433,N_5091);
and U6307 (N_6307,N_5645,N_5001);
nand U6308 (N_6308,N_5522,N_5343);
nor U6309 (N_6309,N_5997,N_5815);
and U6310 (N_6310,N_5946,N_5626);
nor U6311 (N_6311,N_5869,N_5533);
or U6312 (N_6312,N_5355,N_5347);
nand U6313 (N_6313,N_5783,N_5986);
nor U6314 (N_6314,N_5096,N_5318);
nor U6315 (N_6315,N_5955,N_5856);
xnor U6316 (N_6316,N_5930,N_5843);
and U6317 (N_6317,N_5132,N_5620);
or U6318 (N_6318,N_5552,N_5013);
or U6319 (N_6319,N_5624,N_5225);
or U6320 (N_6320,N_5363,N_5589);
nor U6321 (N_6321,N_5101,N_5208);
nor U6322 (N_6322,N_5290,N_5092);
nor U6323 (N_6323,N_5758,N_5977);
nand U6324 (N_6324,N_5278,N_5473);
xor U6325 (N_6325,N_5126,N_5100);
nor U6326 (N_6326,N_5918,N_5924);
nor U6327 (N_6327,N_5577,N_5803);
and U6328 (N_6328,N_5602,N_5598);
or U6329 (N_6329,N_5407,N_5430);
xnor U6330 (N_6330,N_5309,N_5495);
xor U6331 (N_6331,N_5103,N_5240);
xnor U6332 (N_6332,N_5393,N_5795);
nor U6333 (N_6333,N_5236,N_5029);
or U6334 (N_6334,N_5746,N_5575);
nand U6335 (N_6335,N_5065,N_5060);
nor U6336 (N_6336,N_5543,N_5176);
and U6337 (N_6337,N_5854,N_5302);
nor U6338 (N_6338,N_5736,N_5836);
or U6339 (N_6339,N_5515,N_5051);
nor U6340 (N_6340,N_5850,N_5632);
nor U6341 (N_6341,N_5548,N_5024);
xnor U6342 (N_6342,N_5507,N_5559);
or U6343 (N_6343,N_5179,N_5109);
nor U6344 (N_6344,N_5351,N_5173);
nand U6345 (N_6345,N_5796,N_5926);
nor U6346 (N_6346,N_5730,N_5689);
or U6347 (N_6347,N_5668,N_5810);
xor U6348 (N_6348,N_5835,N_5026);
nor U6349 (N_6349,N_5505,N_5940);
nand U6350 (N_6350,N_5353,N_5581);
nand U6351 (N_6351,N_5465,N_5206);
or U6352 (N_6352,N_5143,N_5534);
nor U6353 (N_6353,N_5751,N_5055);
nand U6354 (N_6354,N_5765,N_5186);
xor U6355 (N_6355,N_5342,N_5655);
nand U6356 (N_6356,N_5119,N_5896);
and U6357 (N_6357,N_5041,N_5916);
nor U6358 (N_6358,N_5650,N_5631);
nand U6359 (N_6359,N_5779,N_5841);
nor U6360 (N_6360,N_5472,N_5106);
or U6361 (N_6361,N_5611,N_5315);
or U6362 (N_6362,N_5131,N_5994);
nand U6363 (N_6363,N_5840,N_5072);
xor U6364 (N_6364,N_5189,N_5806);
or U6365 (N_6365,N_5773,N_5199);
nand U6366 (N_6366,N_5475,N_5567);
xor U6367 (N_6367,N_5546,N_5456);
or U6368 (N_6368,N_5742,N_5979);
xor U6369 (N_6369,N_5780,N_5863);
nor U6370 (N_6370,N_5506,N_5499);
nor U6371 (N_6371,N_5723,N_5440);
nand U6372 (N_6372,N_5804,N_5259);
xnor U6373 (N_6373,N_5025,N_5216);
or U6374 (N_6374,N_5618,N_5678);
and U6375 (N_6375,N_5223,N_5980);
nand U6376 (N_6376,N_5851,N_5141);
xor U6377 (N_6377,N_5436,N_5485);
and U6378 (N_6378,N_5849,N_5210);
and U6379 (N_6379,N_5254,N_5374);
xnor U6380 (N_6380,N_5683,N_5520);
nor U6381 (N_6381,N_5392,N_5338);
xnor U6382 (N_6382,N_5703,N_5250);
or U6383 (N_6383,N_5298,N_5007);
or U6384 (N_6384,N_5221,N_5526);
xnor U6385 (N_6385,N_5086,N_5950);
xor U6386 (N_6386,N_5420,N_5541);
nor U6387 (N_6387,N_5417,N_5903);
xor U6388 (N_6388,N_5184,N_5570);
xor U6389 (N_6389,N_5797,N_5525);
nand U6390 (N_6390,N_5108,N_5600);
nand U6391 (N_6391,N_5489,N_5502);
nor U6392 (N_6392,N_5215,N_5447);
nand U6393 (N_6393,N_5435,N_5322);
or U6394 (N_6394,N_5009,N_5855);
xnor U6395 (N_6395,N_5957,N_5415);
nand U6396 (N_6396,N_5261,N_5352);
xnor U6397 (N_6397,N_5781,N_5069);
xor U6398 (N_6398,N_5970,N_5651);
nand U6399 (N_6399,N_5923,N_5246);
nor U6400 (N_6400,N_5893,N_5414);
or U6401 (N_6401,N_5453,N_5949);
or U6402 (N_6402,N_5418,N_5876);
or U6403 (N_6403,N_5202,N_5286);
or U6404 (N_6404,N_5155,N_5129);
nor U6405 (N_6405,N_5532,N_5592);
xor U6406 (N_6406,N_5040,N_5648);
nand U6407 (N_6407,N_5715,N_5793);
and U6408 (N_6408,N_5615,N_5368);
xnor U6409 (N_6409,N_5232,N_5012);
or U6410 (N_6410,N_5941,N_5595);
nand U6411 (N_6411,N_5354,N_5110);
xnor U6412 (N_6412,N_5479,N_5733);
or U6413 (N_6413,N_5400,N_5728);
or U6414 (N_6414,N_5020,N_5792);
and U6415 (N_6415,N_5938,N_5838);
or U6416 (N_6416,N_5910,N_5762);
or U6417 (N_6417,N_5078,N_5284);
xor U6418 (N_6418,N_5191,N_5944);
nor U6419 (N_6419,N_5380,N_5043);
and U6420 (N_6420,N_5609,N_5935);
or U6421 (N_6421,N_5217,N_5037);
or U6422 (N_6422,N_5750,N_5075);
xnor U6423 (N_6423,N_5741,N_5395);
nand U6424 (N_6424,N_5194,N_5823);
nand U6425 (N_6425,N_5492,N_5749);
xor U6426 (N_6426,N_5881,N_5847);
xor U6427 (N_6427,N_5603,N_5498);
and U6428 (N_6428,N_5993,N_5757);
xor U6429 (N_6429,N_5960,N_5877);
nand U6430 (N_6430,N_5102,N_5327);
and U6431 (N_6431,N_5463,N_5964);
or U6432 (N_6432,N_5663,N_5310);
nor U6433 (N_6433,N_5358,N_5879);
xor U6434 (N_6434,N_5198,N_5590);
nand U6435 (N_6435,N_5763,N_5105);
xor U6436 (N_6436,N_5898,N_5253);
nand U6437 (N_6437,N_5458,N_5549);
or U6438 (N_6438,N_5830,N_5700);
nor U6439 (N_6439,N_5477,N_5846);
nor U6440 (N_6440,N_5867,N_5488);
or U6441 (N_6441,N_5243,N_5280);
or U6442 (N_6442,N_5878,N_5637);
and U6443 (N_6443,N_5748,N_5188);
nor U6444 (N_6444,N_5875,N_5927);
or U6445 (N_6445,N_5087,N_5812);
or U6446 (N_6446,N_5153,N_5006);
or U6447 (N_6447,N_5288,N_5324);
and U6448 (N_6448,N_5181,N_5356);
nor U6449 (N_6449,N_5772,N_5673);
and U6450 (N_6450,N_5386,N_5852);
and U6451 (N_6451,N_5171,N_5858);
nor U6452 (N_6452,N_5231,N_5329);
or U6453 (N_6453,N_5381,N_5367);
and U6454 (N_6454,N_5030,N_5886);
and U6455 (N_6455,N_5677,N_5444);
xnor U6456 (N_6456,N_5708,N_5514);
nor U6457 (N_6457,N_5929,N_5469);
nor U6458 (N_6458,N_5501,N_5555);
and U6459 (N_6459,N_5586,N_5527);
nor U6460 (N_6460,N_5561,N_5349);
or U6461 (N_6461,N_5642,N_5378);
nand U6462 (N_6462,N_5661,N_5128);
nor U6463 (N_6463,N_5002,N_5718);
xor U6464 (N_6464,N_5791,N_5340);
nand U6465 (N_6465,N_5939,N_5808);
or U6466 (N_6466,N_5599,N_5870);
or U6467 (N_6467,N_5282,N_5671);
xnor U6468 (N_6468,N_5516,N_5971);
and U6469 (N_6469,N_5134,N_5320);
and U6470 (N_6470,N_5016,N_5300);
and U6471 (N_6471,N_5784,N_5958);
xor U6472 (N_6472,N_5756,N_5157);
nand U6473 (N_6473,N_5032,N_5305);
nand U6474 (N_6474,N_5151,N_5915);
nor U6475 (N_6475,N_5421,N_5149);
and U6476 (N_6476,N_5466,N_5235);
or U6477 (N_6477,N_5281,N_5113);
nand U6478 (N_6478,N_5770,N_5554);
or U6479 (N_6479,N_5568,N_5187);
and U6480 (N_6480,N_5790,N_5764);
xor U6481 (N_6481,N_5572,N_5968);
nand U6482 (N_6482,N_5517,N_5734);
and U6483 (N_6483,N_5292,N_5871);
nand U6484 (N_6484,N_5496,N_5262);
xnor U6485 (N_6485,N_5449,N_5954);
nand U6486 (N_6486,N_5256,N_5766);
or U6487 (N_6487,N_5649,N_5607);
xor U6488 (N_6488,N_5314,N_5470);
or U6489 (N_6489,N_5248,N_5076);
and U6490 (N_6490,N_5018,N_5257);
or U6491 (N_6491,N_5014,N_5776);
or U6492 (N_6492,N_5464,N_5884);
nor U6493 (N_6493,N_5369,N_5814);
xnor U6494 (N_6494,N_5685,N_5169);
nand U6495 (N_6495,N_5019,N_5755);
nor U6496 (N_6496,N_5963,N_5039);
and U6497 (N_6497,N_5638,N_5074);
and U6498 (N_6498,N_5769,N_5423);
nor U6499 (N_6499,N_5098,N_5379);
and U6500 (N_6500,N_5041,N_5130);
and U6501 (N_6501,N_5847,N_5242);
nor U6502 (N_6502,N_5677,N_5261);
xor U6503 (N_6503,N_5938,N_5771);
nor U6504 (N_6504,N_5394,N_5999);
nor U6505 (N_6505,N_5393,N_5542);
and U6506 (N_6506,N_5107,N_5181);
and U6507 (N_6507,N_5806,N_5064);
and U6508 (N_6508,N_5788,N_5222);
nand U6509 (N_6509,N_5528,N_5806);
xnor U6510 (N_6510,N_5558,N_5610);
and U6511 (N_6511,N_5855,N_5627);
nand U6512 (N_6512,N_5313,N_5153);
nor U6513 (N_6513,N_5582,N_5699);
nand U6514 (N_6514,N_5356,N_5828);
and U6515 (N_6515,N_5412,N_5233);
nand U6516 (N_6516,N_5507,N_5702);
or U6517 (N_6517,N_5469,N_5903);
or U6518 (N_6518,N_5907,N_5971);
nor U6519 (N_6519,N_5504,N_5650);
nor U6520 (N_6520,N_5242,N_5310);
nor U6521 (N_6521,N_5210,N_5870);
nand U6522 (N_6522,N_5113,N_5844);
xor U6523 (N_6523,N_5576,N_5215);
xnor U6524 (N_6524,N_5431,N_5255);
nand U6525 (N_6525,N_5121,N_5202);
and U6526 (N_6526,N_5168,N_5052);
xnor U6527 (N_6527,N_5523,N_5890);
nand U6528 (N_6528,N_5913,N_5291);
nand U6529 (N_6529,N_5691,N_5518);
or U6530 (N_6530,N_5763,N_5648);
nor U6531 (N_6531,N_5012,N_5205);
and U6532 (N_6532,N_5522,N_5988);
nand U6533 (N_6533,N_5730,N_5257);
xor U6534 (N_6534,N_5485,N_5086);
or U6535 (N_6535,N_5280,N_5962);
nor U6536 (N_6536,N_5602,N_5500);
or U6537 (N_6537,N_5422,N_5125);
or U6538 (N_6538,N_5645,N_5780);
nor U6539 (N_6539,N_5301,N_5126);
xor U6540 (N_6540,N_5190,N_5866);
nor U6541 (N_6541,N_5240,N_5485);
or U6542 (N_6542,N_5572,N_5321);
or U6543 (N_6543,N_5430,N_5962);
xnor U6544 (N_6544,N_5375,N_5051);
nor U6545 (N_6545,N_5012,N_5421);
and U6546 (N_6546,N_5596,N_5565);
or U6547 (N_6547,N_5201,N_5738);
nand U6548 (N_6548,N_5088,N_5977);
xnor U6549 (N_6549,N_5231,N_5197);
nand U6550 (N_6550,N_5551,N_5835);
and U6551 (N_6551,N_5923,N_5550);
xor U6552 (N_6552,N_5518,N_5404);
xnor U6553 (N_6553,N_5356,N_5837);
nor U6554 (N_6554,N_5423,N_5905);
nand U6555 (N_6555,N_5410,N_5458);
and U6556 (N_6556,N_5636,N_5754);
or U6557 (N_6557,N_5028,N_5221);
xnor U6558 (N_6558,N_5286,N_5003);
or U6559 (N_6559,N_5747,N_5740);
and U6560 (N_6560,N_5948,N_5350);
xnor U6561 (N_6561,N_5984,N_5737);
nand U6562 (N_6562,N_5026,N_5424);
nand U6563 (N_6563,N_5503,N_5826);
xnor U6564 (N_6564,N_5339,N_5667);
nand U6565 (N_6565,N_5718,N_5991);
or U6566 (N_6566,N_5153,N_5753);
or U6567 (N_6567,N_5456,N_5633);
and U6568 (N_6568,N_5495,N_5186);
xnor U6569 (N_6569,N_5466,N_5971);
nor U6570 (N_6570,N_5217,N_5483);
and U6571 (N_6571,N_5007,N_5831);
or U6572 (N_6572,N_5304,N_5530);
and U6573 (N_6573,N_5958,N_5961);
and U6574 (N_6574,N_5367,N_5818);
nor U6575 (N_6575,N_5320,N_5091);
or U6576 (N_6576,N_5153,N_5987);
or U6577 (N_6577,N_5902,N_5349);
xor U6578 (N_6578,N_5081,N_5177);
or U6579 (N_6579,N_5664,N_5158);
xor U6580 (N_6580,N_5845,N_5496);
and U6581 (N_6581,N_5481,N_5474);
nor U6582 (N_6582,N_5547,N_5113);
xor U6583 (N_6583,N_5632,N_5532);
nor U6584 (N_6584,N_5134,N_5305);
nor U6585 (N_6585,N_5485,N_5210);
or U6586 (N_6586,N_5865,N_5068);
nand U6587 (N_6587,N_5110,N_5054);
xor U6588 (N_6588,N_5628,N_5214);
xor U6589 (N_6589,N_5116,N_5764);
and U6590 (N_6590,N_5700,N_5986);
nor U6591 (N_6591,N_5234,N_5951);
xnor U6592 (N_6592,N_5990,N_5513);
and U6593 (N_6593,N_5590,N_5494);
nor U6594 (N_6594,N_5568,N_5458);
nor U6595 (N_6595,N_5638,N_5796);
nand U6596 (N_6596,N_5987,N_5655);
nand U6597 (N_6597,N_5169,N_5812);
xor U6598 (N_6598,N_5081,N_5716);
nor U6599 (N_6599,N_5368,N_5631);
nor U6600 (N_6600,N_5821,N_5096);
xor U6601 (N_6601,N_5300,N_5218);
and U6602 (N_6602,N_5030,N_5733);
xnor U6603 (N_6603,N_5704,N_5127);
or U6604 (N_6604,N_5083,N_5819);
nand U6605 (N_6605,N_5980,N_5115);
or U6606 (N_6606,N_5331,N_5008);
nor U6607 (N_6607,N_5657,N_5706);
nor U6608 (N_6608,N_5883,N_5008);
and U6609 (N_6609,N_5466,N_5438);
or U6610 (N_6610,N_5398,N_5251);
nor U6611 (N_6611,N_5576,N_5063);
and U6612 (N_6612,N_5792,N_5551);
xor U6613 (N_6613,N_5070,N_5314);
nor U6614 (N_6614,N_5465,N_5877);
or U6615 (N_6615,N_5698,N_5662);
nor U6616 (N_6616,N_5001,N_5912);
xor U6617 (N_6617,N_5004,N_5742);
or U6618 (N_6618,N_5984,N_5954);
xnor U6619 (N_6619,N_5062,N_5065);
nor U6620 (N_6620,N_5491,N_5975);
xor U6621 (N_6621,N_5594,N_5478);
nor U6622 (N_6622,N_5388,N_5858);
and U6623 (N_6623,N_5251,N_5799);
nor U6624 (N_6624,N_5582,N_5396);
or U6625 (N_6625,N_5428,N_5523);
and U6626 (N_6626,N_5365,N_5166);
xnor U6627 (N_6627,N_5814,N_5259);
or U6628 (N_6628,N_5185,N_5895);
and U6629 (N_6629,N_5933,N_5621);
xor U6630 (N_6630,N_5672,N_5114);
and U6631 (N_6631,N_5190,N_5683);
and U6632 (N_6632,N_5362,N_5901);
or U6633 (N_6633,N_5512,N_5892);
nor U6634 (N_6634,N_5801,N_5741);
nor U6635 (N_6635,N_5676,N_5025);
or U6636 (N_6636,N_5582,N_5094);
and U6637 (N_6637,N_5674,N_5858);
xnor U6638 (N_6638,N_5451,N_5773);
nand U6639 (N_6639,N_5613,N_5791);
nor U6640 (N_6640,N_5007,N_5827);
nor U6641 (N_6641,N_5370,N_5465);
or U6642 (N_6642,N_5162,N_5161);
and U6643 (N_6643,N_5692,N_5023);
and U6644 (N_6644,N_5473,N_5003);
and U6645 (N_6645,N_5666,N_5668);
nor U6646 (N_6646,N_5469,N_5074);
or U6647 (N_6647,N_5712,N_5819);
nor U6648 (N_6648,N_5303,N_5152);
nand U6649 (N_6649,N_5329,N_5973);
or U6650 (N_6650,N_5785,N_5856);
nand U6651 (N_6651,N_5268,N_5726);
or U6652 (N_6652,N_5870,N_5658);
nor U6653 (N_6653,N_5948,N_5034);
or U6654 (N_6654,N_5430,N_5487);
nor U6655 (N_6655,N_5418,N_5838);
and U6656 (N_6656,N_5357,N_5928);
nor U6657 (N_6657,N_5982,N_5509);
nor U6658 (N_6658,N_5394,N_5751);
or U6659 (N_6659,N_5020,N_5025);
nor U6660 (N_6660,N_5012,N_5249);
or U6661 (N_6661,N_5645,N_5015);
or U6662 (N_6662,N_5906,N_5723);
nand U6663 (N_6663,N_5864,N_5075);
nand U6664 (N_6664,N_5653,N_5215);
and U6665 (N_6665,N_5933,N_5896);
or U6666 (N_6666,N_5691,N_5576);
or U6667 (N_6667,N_5257,N_5108);
nand U6668 (N_6668,N_5978,N_5316);
and U6669 (N_6669,N_5148,N_5046);
nor U6670 (N_6670,N_5627,N_5095);
xnor U6671 (N_6671,N_5719,N_5121);
xor U6672 (N_6672,N_5810,N_5982);
nor U6673 (N_6673,N_5302,N_5489);
nand U6674 (N_6674,N_5944,N_5228);
and U6675 (N_6675,N_5352,N_5147);
xnor U6676 (N_6676,N_5513,N_5851);
xnor U6677 (N_6677,N_5894,N_5229);
or U6678 (N_6678,N_5882,N_5935);
and U6679 (N_6679,N_5023,N_5485);
and U6680 (N_6680,N_5026,N_5637);
or U6681 (N_6681,N_5417,N_5376);
xnor U6682 (N_6682,N_5655,N_5506);
xor U6683 (N_6683,N_5986,N_5808);
or U6684 (N_6684,N_5277,N_5678);
and U6685 (N_6685,N_5602,N_5161);
or U6686 (N_6686,N_5791,N_5358);
xor U6687 (N_6687,N_5104,N_5427);
and U6688 (N_6688,N_5091,N_5594);
xor U6689 (N_6689,N_5834,N_5973);
and U6690 (N_6690,N_5359,N_5829);
nand U6691 (N_6691,N_5972,N_5188);
nor U6692 (N_6692,N_5775,N_5550);
nor U6693 (N_6693,N_5573,N_5669);
or U6694 (N_6694,N_5668,N_5674);
and U6695 (N_6695,N_5322,N_5120);
and U6696 (N_6696,N_5666,N_5361);
xor U6697 (N_6697,N_5200,N_5733);
xnor U6698 (N_6698,N_5393,N_5626);
or U6699 (N_6699,N_5760,N_5446);
xnor U6700 (N_6700,N_5492,N_5146);
or U6701 (N_6701,N_5480,N_5999);
xor U6702 (N_6702,N_5821,N_5914);
nor U6703 (N_6703,N_5325,N_5898);
or U6704 (N_6704,N_5085,N_5038);
nand U6705 (N_6705,N_5622,N_5815);
or U6706 (N_6706,N_5845,N_5531);
xnor U6707 (N_6707,N_5755,N_5609);
nor U6708 (N_6708,N_5896,N_5197);
or U6709 (N_6709,N_5301,N_5910);
nor U6710 (N_6710,N_5089,N_5774);
nor U6711 (N_6711,N_5306,N_5827);
xnor U6712 (N_6712,N_5922,N_5404);
or U6713 (N_6713,N_5497,N_5235);
nor U6714 (N_6714,N_5825,N_5191);
or U6715 (N_6715,N_5977,N_5736);
or U6716 (N_6716,N_5600,N_5346);
and U6717 (N_6717,N_5938,N_5660);
or U6718 (N_6718,N_5049,N_5172);
xor U6719 (N_6719,N_5755,N_5577);
and U6720 (N_6720,N_5566,N_5427);
or U6721 (N_6721,N_5980,N_5338);
or U6722 (N_6722,N_5526,N_5921);
nor U6723 (N_6723,N_5309,N_5057);
nor U6724 (N_6724,N_5017,N_5544);
nand U6725 (N_6725,N_5494,N_5280);
nand U6726 (N_6726,N_5505,N_5969);
nand U6727 (N_6727,N_5060,N_5130);
or U6728 (N_6728,N_5313,N_5181);
nor U6729 (N_6729,N_5634,N_5345);
nand U6730 (N_6730,N_5690,N_5877);
and U6731 (N_6731,N_5436,N_5659);
and U6732 (N_6732,N_5041,N_5943);
or U6733 (N_6733,N_5815,N_5533);
nor U6734 (N_6734,N_5424,N_5334);
nand U6735 (N_6735,N_5064,N_5208);
nor U6736 (N_6736,N_5300,N_5921);
nand U6737 (N_6737,N_5500,N_5482);
nand U6738 (N_6738,N_5270,N_5949);
xnor U6739 (N_6739,N_5958,N_5246);
and U6740 (N_6740,N_5329,N_5725);
nand U6741 (N_6741,N_5903,N_5284);
nand U6742 (N_6742,N_5138,N_5974);
nor U6743 (N_6743,N_5275,N_5560);
nor U6744 (N_6744,N_5680,N_5067);
and U6745 (N_6745,N_5995,N_5747);
xnor U6746 (N_6746,N_5343,N_5070);
or U6747 (N_6747,N_5255,N_5343);
xnor U6748 (N_6748,N_5406,N_5849);
nand U6749 (N_6749,N_5055,N_5000);
nand U6750 (N_6750,N_5492,N_5024);
and U6751 (N_6751,N_5964,N_5022);
or U6752 (N_6752,N_5236,N_5954);
xor U6753 (N_6753,N_5536,N_5309);
xor U6754 (N_6754,N_5380,N_5828);
and U6755 (N_6755,N_5819,N_5300);
and U6756 (N_6756,N_5083,N_5116);
nor U6757 (N_6757,N_5475,N_5725);
xnor U6758 (N_6758,N_5595,N_5137);
xnor U6759 (N_6759,N_5193,N_5763);
xnor U6760 (N_6760,N_5548,N_5523);
and U6761 (N_6761,N_5172,N_5083);
nand U6762 (N_6762,N_5529,N_5580);
nand U6763 (N_6763,N_5020,N_5757);
xnor U6764 (N_6764,N_5051,N_5852);
nor U6765 (N_6765,N_5952,N_5168);
nand U6766 (N_6766,N_5368,N_5123);
xor U6767 (N_6767,N_5688,N_5595);
nor U6768 (N_6768,N_5558,N_5450);
or U6769 (N_6769,N_5915,N_5425);
nand U6770 (N_6770,N_5038,N_5903);
nor U6771 (N_6771,N_5887,N_5749);
nand U6772 (N_6772,N_5285,N_5604);
xnor U6773 (N_6773,N_5287,N_5827);
and U6774 (N_6774,N_5595,N_5728);
nand U6775 (N_6775,N_5729,N_5296);
nand U6776 (N_6776,N_5336,N_5370);
xor U6777 (N_6777,N_5022,N_5138);
and U6778 (N_6778,N_5171,N_5924);
nand U6779 (N_6779,N_5651,N_5104);
nand U6780 (N_6780,N_5120,N_5082);
and U6781 (N_6781,N_5456,N_5580);
nand U6782 (N_6782,N_5977,N_5488);
nand U6783 (N_6783,N_5884,N_5969);
and U6784 (N_6784,N_5687,N_5624);
nor U6785 (N_6785,N_5210,N_5427);
or U6786 (N_6786,N_5560,N_5462);
and U6787 (N_6787,N_5509,N_5811);
nor U6788 (N_6788,N_5775,N_5530);
nand U6789 (N_6789,N_5349,N_5094);
nand U6790 (N_6790,N_5559,N_5487);
xnor U6791 (N_6791,N_5434,N_5797);
xor U6792 (N_6792,N_5411,N_5859);
or U6793 (N_6793,N_5544,N_5323);
xor U6794 (N_6794,N_5789,N_5530);
nor U6795 (N_6795,N_5550,N_5194);
nand U6796 (N_6796,N_5302,N_5818);
nand U6797 (N_6797,N_5432,N_5623);
and U6798 (N_6798,N_5256,N_5041);
and U6799 (N_6799,N_5734,N_5679);
nand U6800 (N_6800,N_5325,N_5087);
and U6801 (N_6801,N_5246,N_5174);
nor U6802 (N_6802,N_5113,N_5246);
nand U6803 (N_6803,N_5396,N_5182);
nor U6804 (N_6804,N_5302,N_5957);
nor U6805 (N_6805,N_5309,N_5962);
or U6806 (N_6806,N_5289,N_5673);
xnor U6807 (N_6807,N_5503,N_5513);
and U6808 (N_6808,N_5957,N_5373);
or U6809 (N_6809,N_5724,N_5395);
nor U6810 (N_6810,N_5991,N_5393);
nor U6811 (N_6811,N_5567,N_5304);
and U6812 (N_6812,N_5271,N_5968);
nand U6813 (N_6813,N_5157,N_5891);
or U6814 (N_6814,N_5780,N_5101);
nand U6815 (N_6815,N_5299,N_5346);
or U6816 (N_6816,N_5058,N_5305);
xnor U6817 (N_6817,N_5213,N_5954);
xor U6818 (N_6818,N_5570,N_5092);
nor U6819 (N_6819,N_5743,N_5682);
or U6820 (N_6820,N_5316,N_5931);
nand U6821 (N_6821,N_5494,N_5675);
and U6822 (N_6822,N_5954,N_5013);
xnor U6823 (N_6823,N_5426,N_5288);
or U6824 (N_6824,N_5045,N_5784);
xnor U6825 (N_6825,N_5344,N_5146);
or U6826 (N_6826,N_5908,N_5446);
xnor U6827 (N_6827,N_5963,N_5604);
xor U6828 (N_6828,N_5903,N_5515);
xor U6829 (N_6829,N_5197,N_5828);
or U6830 (N_6830,N_5099,N_5399);
xnor U6831 (N_6831,N_5301,N_5383);
nand U6832 (N_6832,N_5881,N_5014);
and U6833 (N_6833,N_5316,N_5716);
nand U6834 (N_6834,N_5692,N_5140);
or U6835 (N_6835,N_5473,N_5981);
nand U6836 (N_6836,N_5934,N_5643);
and U6837 (N_6837,N_5457,N_5806);
xnor U6838 (N_6838,N_5497,N_5611);
nand U6839 (N_6839,N_5653,N_5119);
or U6840 (N_6840,N_5164,N_5455);
nor U6841 (N_6841,N_5740,N_5219);
nor U6842 (N_6842,N_5028,N_5039);
nor U6843 (N_6843,N_5552,N_5803);
nor U6844 (N_6844,N_5098,N_5028);
or U6845 (N_6845,N_5244,N_5522);
nand U6846 (N_6846,N_5620,N_5457);
nand U6847 (N_6847,N_5452,N_5117);
nor U6848 (N_6848,N_5113,N_5849);
and U6849 (N_6849,N_5808,N_5774);
nand U6850 (N_6850,N_5263,N_5936);
xnor U6851 (N_6851,N_5368,N_5488);
nand U6852 (N_6852,N_5887,N_5338);
xnor U6853 (N_6853,N_5351,N_5675);
and U6854 (N_6854,N_5400,N_5885);
xnor U6855 (N_6855,N_5033,N_5833);
or U6856 (N_6856,N_5691,N_5335);
xor U6857 (N_6857,N_5725,N_5724);
nand U6858 (N_6858,N_5710,N_5836);
nand U6859 (N_6859,N_5589,N_5545);
nand U6860 (N_6860,N_5440,N_5918);
or U6861 (N_6861,N_5813,N_5978);
and U6862 (N_6862,N_5868,N_5894);
nor U6863 (N_6863,N_5599,N_5871);
xnor U6864 (N_6864,N_5893,N_5772);
or U6865 (N_6865,N_5491,N_5506);
xnor U6866 (N_6866,N_5962,N_5422);
nand U6867 (N_6867,N_5675,N_5202);
xnor U6868 (N_6868,N_5287,N_5754);
nor U6869 (N_6869,N_5758,N_5572);
or U6870 (N_6870,N_5959,N_5367);
and U6871 (N_6871,N_5985,N_5839);
and U6872 (N_6872,N_5178,N_5982);
xnor U6873 (N_6873,N_5633,N_5922);
or U6874 (N_6874,N_5593,N_5203);
nand U6875 (N_6875,N_5656,N_5791);
nand U6876 (N_6876,N_5543,N_5672);
nor U6877 (N_6877,N_5890,N_5845);
and U6878 (N_6878,N_5120,N_5130);
xor U6879 (N_6879,N_5574,N_5083);
or U6880 (N_6880,N_5968,N_5025);
nand U6881 (N_6881,N_5583,N_5648);
nor U6882 (N_6882,N_5515,N_5092);
nor U6883 (N_6883,N_5744,N_5965);
xor U6884 (N_6884,N_5524,N_5438);
and U6885 (N_6885,N_5643,N_5306);
nor U6886 (N_6886,N_5504,N_5367);
and U6887 (N_6887,N_5748,N_5545);
xnor U6888 (N_6888,N_5034,N_5510);
nor U6889 (N_6889,N_5160,N_5069);
nor U6890 (N_6890,N_5900,N_5283);
nor U6891 (N_6891,N_5149,N_5262);
xor U6892 (N_6892,N_5688,N_5859);
nor U6893 (N_6893,N_5879,N_5912);
or U6894 (N_6894,N_5441,N_5296);
and U6895 (N_6895,N_5626,N_5693);
and U6896 (N_6896,N_5570,N_5327);
nor U6897 (N_6897,N_5372,N_5894);
xor U6898 (N_6898,N_5265,N_5088);
nand U6899 (N_6899,N_5263,N_5626);
and U6900 (N_6900,N_5422,N_5230);
xnor U6901 (N_6901,N_5263,N_5997);
or U6902 (N_6902,N_5993,N_5652);
nor U6903 (N_6903,N_5104,N_5717);
nor U6904 (N_6904,N_5863,N_5251);
nor U6905 (N_6905,N_5227,N_5637);
nor U6906 (N_6906,N_5236,N_5540);
and U6907 (N_6907,N_5047,N_5522);
nand U6908 (N_6908,N_5987,N_5258);
nand U6909 (N_6909,N_5634,N_5225);
xor U6910 (N_6910,N_5395,N_5828);
and U6911 (N_6911,N_5894,N_5213);
nor U6912 (N_6912,N_5139,N_5634);
nand U6913 (N_6913,N_5587,N_5886);
xor U6914 (N_6914,N_5984,N_5694);
nand U6915 (N_6915,N_5805,N_5380);
and U6916 (N_6916,N_5513,N_5419);
nor U6917 (N_6917,N_5423,N_5479);
and U6918 (N_6918,N_5228,N_5189);
and U6919 (N_6919,N_5988,N_5934);
nor U6920 (N_6920,N_5524,N_5156);
xnor U6921 (N_6921,N_5871,N_5121);
nand U6922 (N_6922,N_5637,N_5588);
xnor U6923 (N_6923,N_5820,N_5887);
and U6924 (N_6924,N_5912,N_5881);
nor U6925 (N_6925,N_5885,N_5620);
xnor U6926 (N_6926,N_5108,N_5454);
xnor U6927 (N_6927,N_5465,N_5533);
and U6928 (N_6928,N_5337,N_5382);
and U6929 (N_6929,N_5895,N_5701);
or U6930 (N_6930,N_5860,N_5225);
and U6931 (N_6931,N_5544,N_5104);
xnor U6932 (N_6932,N_5632,N_5013);
and U6933 (N_6933,N_5207,N_5854);
or U6934 (N_6934,N_5923,N_5769);
nand U6935 (N_6935,N_5593,N_5911);
or U6936 (N_6936,N_5803,N_5463);
and U6937 (N_6937,N_5875,N_5609);
nor U6938 (N_6938,N_5861,N_5772);
and U6939 (N_6939,N_5792,N_5053);
or U6940 (N_6940,N_5811,N_5287);
nor U6941 (N_6941,N_5683,N_5678);
nand U6942 (N_6942,N_5210,N_5518);
nand U6943 (N_6943,N_5934,N_5419);
nor U6944 (N_6944,N_5961,N_5002);
xnor U6945 (N_6945,N_5698,N_5513);
xor U6946 (N_6946,N_5362,N_5863);
xnor U6947 (N_6947,N_5753,N_5513);
nand U6948 (N_6948,N_5818,N_5790);
nor U6949 (N_6949,N_5639,N_5262);
xor U6950 (N_6950,N_5872,N_5118);
nor U6951 (N_6951,N_5166,N_5035);
nor U6952 (N_6952,N_5059,N_5779);
xnor U6953 (N_6953,N_5252,N_5573);
nor U6954 (N_6954,N_5800,N_5210);
and U6955 (N_6955,N_5014,N_5798);
xor U6956 (N_6956,N_5211,N_5742);
and U6957 (N_6957,N_5879,N_5656);
and U6958 (N_6958,N_5957,N_5187);
nand U6959 (N_6959,N_5797,N_5748);
and U6960 (N_6960,N_5028,N_5231);
nor U6961 (N_6961,N_5747,N_5573);
nor U6962 (N_6962,N_5035,N_5500);
nand U6963 (N_6963,N_5405,N_5753);
or U6964 (N_6964,N_5664,N_5237);
and U6965 (N_6965,N_5284,N_5633);
and U6966 (N_6966,N_5344,N_5942);
xnor U6967 (N_6967,N_5729,N_5230);
nand U6968 (N_6968,N_5201,N_5743);
nand U6969 (N_6969,N_5455,N_5158);
and U6970 (N_6970,N_5973,N_5426);
and U6971 (N_6971,N_5936,N_5681);
nor U6972 (N_6972,N_5793,N_5712);
nand U6973 (N_6973,N_5555,N_5385);
nor U6974 (N_6974,N_5241,N_5075);
nand U6975 (N_6975,N_5304,N_5817);
nor U6976 (N_6976,N_5930,N_5560);
nand U6977 (N_6977,N_5693,N_5217);
or U6978 (N_6978,N_5139,N_5203);
and U6979 (N_6979,N_5228,N_5214);
xnor U6980 (N_6980,N_5150,N_5828);
or U6981 (N_6981,N_5513,N_5080);
xor U6982 (N_6982,N_5624,N_5325);
and U6983 (N_6983,N_5062,N_5871);
nand U6984 (N_6984,N_5897,N_5670);
nor U6985 (N_6985,N_5546,N_5951);
and U6986 (N_6986,N_5212,N_5977);
and U6987 (N_6987,N_5401,N_5674);
xnor U6988 (N_6988,N_5364,N_5614);
or U6989 (N_6989,N_5011,N_5374);
and U6990 (N_6990,N_5273,N_5267);
and U6991 (N_6991,N_5450,N_5502);
xor U6992 (N_6992,N_5120,N_5395);
nor U6993 (N_6993,N_5862,N_5284);
or U6994 (N_6994,N_5257,N_5691);
xor U6995 (N_6995,N_5368,N_5543);
and U6996 (N_6996,N_5279,N_5999);
nor U6997 (N_6997,N_5962,N_5398);
nand U6998 (N_6998,N_5356,N_5854);
or U6999 (N_6999,N_5930,N_5202);
nor U7000 (N_7000,N_6862,N_6103);
nand U7001 (N_7001,N_6437,N_6373);
nor U7002 (N_7002,N_6704,N_6052);
and U7003 (N_7003,N_6358,N_6520);
and U7004 (N_7004,N_6949,N_6476);
and U7005 (N_7005,N_6564,N_6779);
or U7006 (N_7006,N_6436,N_6843);
and U7007 (N_7007,N_6984,N_6817);
or U7008 (N_7008,N_6709,N_6975);
xnor U7009 (N_7009,N_6488,N_6911);
nor U7010 (N_7010,N_6890,N_6695);
nand U7011 (N_7011,N_6435,N_6896);
nand U7012 (N_7012,N_6874,N_6361);
and U7013 (N_7013,N_6509,N_6357);
nand U7014 (N_7014,N_6586,N_6456);
nor U7015 (N_7015,N_6699,N_6521);
xnor U7016 (N_7016,N_6825,N_6137);
nor U7017 (N_7017,N_6562,N_6302);
nor U7018 (N_7018,N_6875,N_6311);
or U7019 (N_7019,N_6459,N_6215);
and U7020 (N_7020,N_6447,N_6833);
nand U7021 (N_7021,N_6674,N_6517);
nand U7022 (N_7022,N_6392,N_6183);
or U7023 (N_7023,N_6532,N_6180);
and U7024 (N_7024,N_6263,N_6058);
nand U7025 (N_7025,N_6761,N_6479);
and U7026 (N_7026,N_6635,N_6305);
xor U7027 (N_7027,N_6913,N_6427);
or U7028 (N_7028,N_6719,N_6577);
nor U7029 (N_7029,N_6483,N_6527);
and U7030 (N_7030,N_6268,N_6838);
or U7031 (N_7031,N_6953,N_6960);
nand U7032 (N_7032,N_6772,N_6744);
or U7033 (N_7033,N_6248,N_6627);
nor U7034 (N_7034,N_6254,N_6619);
and U7035 (N_7035,N_6714,N_6675);
or U7036 (N_7036,N_6015,N_6548);
or U7037 (N_7037,N_6217,N_6941);
xor U7038 (N_7038,N_6343,N_6687);
nand U7039 (N_7039,N_6725,N_6860);
and U7040 (N_7040,N_6556,N_6579);
nand U7041 (N_7041,N_6482,N_6454);
xor U7042 (N_7042,N_6255,N_6581);
nor U7043 (N_7043,N_6669,N_6227);
or U7044 (N_7044,N_6584,N_6452);
or U7045 (N_7045,N_6059,N_6694);
and U7046 (N_7046,N_6224,N_6603);
xnor U7047 (N_7047,N_6411,N_6750);
or U7048 (N_7048,N_6707,N_6478);
or U7049 (N_7049,N_6800,N_6448);
or U7050 (N_7050,N_6561,N_6028);
nand U7051 (N_7051,N_6464,N_6012);
nand U7052 (N_7052,N_6794,N_6991);
nand U7053 (N_7053,N_6128,N_6956);
or U7054 (N_7054,N_6901,N_6516);
nand U7055 (N_7055,N_6628,N_6943);
nand U7056 (N_7056,N_6216,N_6929);
and U7057 (N_7057,N_6412,N_6904);
xor U7058 (N_7058,N_6115,N_6667);
xor U7059 (N_7059,N_6646,N_6085);
or U7060 (N_7060,N_6283,N_6942);
and U7061 (N_7061,N_6206,N_6125);
and U7062 (N_7062,N_6474,N_6597);
or U7063 (N_7063,N_6848,N_6082);
or U7064 (N_7064,N_6232,N_6788);
xnor U7065 (N_7065,N_6458,N_6225);
or U7066 (N_7066,N_6996,N_6298);
nand U7067 (N_7067,N_6626,N_6193);
xnor U7068 (N_7068,N_6055,N_6442);
and U7069 (N_7069,N_6678,N_6790);
nor U7070 (N_7070,N_6945,N_6202);
xnor U7071 (N_7071,N_6129,N_6332);
nand U7072 (N_7072,N_6401,N_6297);
nand U7073 (N_7073,N_6065,N_6722);
nand U7074 (N_7074,N_6428,N_6054);
and U7075 (N_7075,N_6624,N_6731);
and U7076 (N_7076,N_6819,N_6745);
nand U7077 (N_7077,N_6823,N_6889);
or U7078 (N_7078,N_6824,N_6154);
nor U7079 (N_7079,N_6403,N_6625);
xor U7080 (N_7080,N_6457,N_6831);
nor U7081 (N_7081,N_6952,N_6194);
or U7082 (N_7082,N_6190,N_6106);
or U7083 (N_7083,N_6679,N_6555);
and U7084 (N_7084,N_6023,N_6970);
and U7085 (N_7085,N_6547,N_6680);
xnor U7086 (N_7086,N_6963,N_6449);
nand U7087 (N_7087,N_6024,N_6810);
and U7088 (N_7088,N_6355,N_6208);
nor U7089 (N_7089,N_6124,N_6756);
xor U7090 (N_7090,N_6853,N_6262);
nand U7091 (N_7091,N_6591,N_6836);
nand U7092 (N_7092,N_6220,N_6739);
nor U7093 (N_7093,N_6265,N_6425);
xnor U7094 (N_7094,N_6090,N_6161);
or U7095 (N_7095,N_6391,N_6030);
xnor U7096 (N_7096,N_6347,N_6506);
nor U7097 (N_7097,N_6405,N_6372);
and U7098 (N_7098,N_6293,N_6239);
nor U7099 (N_7099,N_6400,N_6727);
nand U7100 (N_7100,N_6187,N_6368);
or U7101 (N_7101,N_6198,N_6309);
and U7102 (N_7102,N_6152,N_6720);
nor U7103 (N_7103,N_6643,N_6075);
and U7104 (N_7104,N_6869,N_6006);
and U7105 (N_7105,N_6985,N_6267);
nand U7106 (N_7106,N_6191,N_6351);
and U7107 (N_7107,N_6111,N_6087);
and U7108 (N_7108,N_6803,N_6732);
nand U7109 (N_7109,N_6236,N_6431);
and U7110 (N_7110,N_6933,N_6558);
and U7111 (N_7111,N_6492,N_6573);
xnor U7112 (N_7112,N_6374,N_6938);
or U7113 (N_7113,N_6385,N_6326);
nand U7114 (N_7114,N_6257,N_6818);
nor U7115 (N_7115,N_6201,N_6972);
xor U7116 (N_7116,N_6681,N_6529);
and U7117 (N_7117,N_6356,N_6014);
and U7118 (N_7118,N_6086,N_6041);
nor U7119 (N_7119,N_6738,N_6925);
and U7120 (N_7120,N_6341,N_6931);
xor U7121 (N_7121,N_6673,N_6653);
or U7122 (N_7122,N_6246,N_6915);
or U7123 (N_7123,N_6429,N_6583);
and U7124 (N_7124,N_6524,N_6313);
or U7125 (N_7125,N_6852,N_6451);
and U7126 (N_7126,N_6905,N_6621);
xnor U7127 (N_7127,N_6139,N_6753);
or U7128 (N_7128,N_6204,N_6336);
nand U7129 (N_7129,N_6546,N_6430);
nand U7130 (N_7130,N_6001,N_6146);
or U7131 (N_7131,N_6921,N_6671);
xnor U7132 (N_7132,N_6473,N_6064);
or U7133 (N_7133,N_6043,N_6032);
or U7134 (N_7134,N_6820,N_6050);
nand U7135 (N_7135,N_6801,N_6866);
xor U7136 (N_7136,N_6315,N_6652);
or U7137 (N_7137,N_6835,N_6917);
or U7138 (N_7138,N_6544,N_6384);
and U7139 (N_7139,N_6730,N_6636);
or U7140 (N_7140,N_6329,N_6540);
xnor U7141 (N_7141,N_6666,N_6044);
nor U7142 (N_7142,N_6928,N_6763);
nand U7143 (N_7143,N_6986,N_6419);
and U7144 (N_7144,N_6057,N_6640);
xor U7145 (N_7145,N_6535,N_6655);
nor U7146 (N_7146,N_6936,N_6786);
xnor U7147 (N_7147,N_6600,N_6651);
or U7148 (N_7148,N_6770,N_6394);
nor U7149 (N_7149,N_6791,N_6499);
xor U7150 (N_7150,N_6434,N_6560);
nand U7151 (N_7151,N_6379,N_6729);
nor U7152 (N_7152,N_6967,N_6554);
and U7153 (N_7153,N_6229,N_6513);
nor U7154 (N_7154,N_6865,N_6409);
nand U7155 (N_7155,N_6278,N_6117);
nand U7156 (N_7156,N_6290,N_6203);
nand U7157 (N_7157,N_6766,N_6138);
or U7158 (N_7158,N_6010,N_6946);
and U7159 (N_7159,N_6846,N_6701);
nand U7160 (N_7160,N_6842,N_6897);
nor U7161 (N_7161,N_6935,N_6333);
and U7162 (N_7162,N_6370,N_6710);
nand U7163 (N_7163,N_6609,N_6887);
xnor U7164 (N_7164,N_6153,N_6036);
xnor U7165 (N_7165,N_6784,N_6049);
or U7166 (N_7166,N_6839,N_6533);
nand U7167 (N_7167,N_6100,N_6299);
and U7168 (N_7168,N_6330,N_6169);
nand U7169 (N_7169,N_6027,N_6785);
nor U7170 (N_7170,N_6740,N_6205);
or U7171 (N_7171,N_6250,N_6120);
and U7172 (N_7172,N_6119,N_6777);
nand U7173 (N_7173,N_6053,N_6092);
or U7174 (N_7174,N_6498,N_6261);
xor U7175 (N_7175,N_6295,N_6961);
nor U7176 (N_7176,N_6815,N_6570);
xor U7177 (N_7177,N_6172,N_6567);
or U7178 (N_7178,N_6211,N_6654);
and U7179 (N_7179,N_6335,N_6571);
nand U7180 (N_7180,N_6551,N_6622);
nand U7181 (N_7181,N_6408,N_6633);
or U7182 (N_7182,N_6070,N_6608);
and U7183 (N_7183,N_6214,N_6787);
and U7184 (N_7184,N_6317,N_6559);
xnor U7185 (N_7185,N_6510,N_6182);
nand U7186 (N_7186,N_6281,N_6662);
nand U7187 (N_7187,N_6514,N_6795);
or U7188 (N_7188,N_6525,N_6539);
xor U7189 (N_7189,N_6156,N_6926);
nand U7190 (N_7190,N_6883,N_6375);
nor U7191 (N_7191,N_6620,N_6076);
and U7192 (N_7192,N_6410,N_6876);
xor U7193 (N_7193,N_6140,N_6523);
and U7194 (N_7194,N_6614,N_6439);
or U7195 (N_7195,N_6016,N_6098);
nand U7196 (N_7196,N_6512,N_6136);
xnor U7197 (N_7197,N_6197,N_6418);
nand U7198 (N_7198,N_6954,N_6402);
nor U7199 (N_7199,N_6017,N_6645);
and U7200 (N_7200,N_6046,N_6184);
and U7201 (N_7201,N_6390,N_6444);
or U7202 (N_7202,N_6241,N_6980);
nor U7203 (N_7203,N_6094,N_6147);
xnor U7204 (N_7204,N_6804,N_6417);
and U7205 (N_7205,N_6407,N_6207);
nand U7206 (N_7206,N_6465,N_6271);
nor U7207 (N_7207,N_6768,N_6445);
nor U7208 (N_7208,N_6338,N_6007);
nand U7209 (N_7209,N_6462,N_6826);
or U7210 (N_7210,N_6109,N_6966);
and U7211 (N_7211,N_6982,N_6393);
xnor U7212 (N_7212,N_6237,N_6944);
nand U7213 (N_7213,N_6327,N_6045);
nand U7214 (N_7214,N_6420,N_6218);
and U7215 (N_7215,N_6598,N_6829);
or U7216 (N_7216,N_6003,N_6665);
or U7217 (N_7217,N_6808,N_6174);
and U7218 (N_7218,N_6979,N_6081);
and U7219 (N_7219,N_6378,N_6895);
xor U7220 (N_7220,N_6397,N_6095);
xor U7221 (N_7221,N_6747,N_6864);
xnor U7222 (N_7222,N_6580,N_6923);
nor U7223 (N_7223,N_6932,N_6048);
xor U7224 (N_7224,N_6350,N_6371);
nand U7225 (N_7225,N_6515,N_6634);
and U7226 (N_7226,N_6959,N_6582);
nand U7227 (N_7227,N_6256,N_6453);
or U7228 (N_7228,N_6757,N_6748);
nor U7229 (N_7229,N_6596,N_6536);
or U7230 (N_7230,N_6522,N_6133);
nor U7231 (N_7231,N_6888,N_6806);
xnor U7232 (N_7232,N_6123,N_6421);
nand U7233 (N_7233,N_6861,N_6181);
or U7234 (N_7234,N_6530,N_6159);
nor U7235 (N_7235,N_6973,N_6922);
and U7236 (N_7236,N_6863,N_6388);
or U7237 (N_7237,N_6637,N_6735);
or U7238 (N_7238,N_6775,N_6828);
nor U7239 (N_7239,N_6993,N_6303);
nand U7240 (N_7240,N_6067,N_6639);
or U7241 (N_7241,N_6446,N_6000);
or U7242 (N_7242,N_6386,N_6534);
nor U7243 (N_7243,N_6920,N_6228);
or U7244 (N_7244,N_6809,N_6934);
and U7245 (N_7245,N_6300,N_6879);
and U7246 (N_7246,N_6307,N_6778);
nor U7247 (N_7247,N_6294,N_6359);
and U7248 (N_7248,N_6244,N_6649);
and U7249 (N_7249,N_6734,N_6576);
and U7250 (N_7250,N_6565,N_6762);
nor U7251 (N_7251,N_6723,N_6323);
and U7252 (N_7252,N_6691,N_6346);
nand U7253 (N_7253,N_6912,N_6741);
and U7254 (N_7254,N_6189,N_6276);
nand U7255 (N_7255,N_6319,N_6280);
xor U7256 (N_7256,N_6360,N_6965);
and U7257 (N_7257,N_6837,N_6051);
xnor U7258 (N_7258,N_6105,N_6604);
or U7259 (N_7259,N_6886,N_6816);
xnor U7260 (N_7260,N_6321,N_6969);
and U7261 (N_7261,N_6178,N_6957);
and U7262 (N_7262,N_6557,N_6497);
and U7263 (N_7263,N_6716,N_6978);
nand U7264 (N_7264,N_6277,N_6776);
nand U7265 (N_7265,N_6519,N_6441);
xor U7266 (N_7266,N_6663,N_6079);
xor U7267 (N_7267,N_6363,N_6176);
or U7268 (N_7268,N_6251,N_6018);
nor U7269 (N_7269,N_6354,N_6141);
xor U7270 (N_7270,N_6868,N_6706);
or U7271 (N_7271,N_6907,N_6316);
nor U7272 (N_7272,N_6684,N_6061);
nor U7273 (N_7273,N_6164,N_6672);
or U7274 (N_7274,N_6387,N_6767);
nand U7275 (N_7275,N_6998,N_6192);
or U7276 (N_7276,N_6287,N_6011);
xnor U7277 (N_7277,N_6163,N_6171);
nor U7278 (N_7278,N_6881,N_6592);
and U7279 (N_7279,N_6867,N_6502);
xnor U7280 (N_7280,N_6212,N_6078);
or U7281 (N_7281,N_6805,N_6541);
and U7282 (N_7282,N_6234,N_6947);
and U7283 (N_7283,N_6781,N_6145);
nand U7284 (N_7284,N_6508,N_6093);
and U7285 (N_7285,N_6084,N_6252);
nor U7286 (N_7286,N_6495,N_6493);
nand U7287 (N_7287,N_6173,N_6526);
and U7288 (N_7288,N_6366,N_6020);
and U7289 (N_7289,N_6132,N_6623);
nor U7290 (N_7290,N_6274,N_6322);
nor U7291 (N_7291,N_6481,N_6594);
nand U7292 (N_7292,N_6796,N_6091);
and U7293 (N_7293,N_6771,N_6712);
nand U7294 (N_7294,N_6670,N_6542);
nand U7295 (N_7295,N_6398,N_6951);
or U7296 (N_7296,N_6110,N_6035);
xor U7297 (N_7297,N_6339,N_6170);
or U7298 (N_7298,N_6759,N_6312);
or U7299 (N_7299,N_6467,N_6563);
nor U7300 (N_7300,N_6769,N_6369);
xnor U7301 (N_7301,N_6013,N_6149);
nor U7302 (N_7302,N_6331,N_6029);
nor U7303 (N_7303,N_6696,N_6113);
xor U7304 (N_7304,N_6650,N_6642);
nor U7305 (N_7305,N_6977,N_6927);
nand U7306 (N_7306,N_6083,N_6891);
nand U7307 (N_7307,N_6814,N_6974);
or U7308 (N_7308,N_6968,N_6047);
nand U7309 (N_7309,N_6460,N_6210);
nand U7310 (N_7310,N_6328,N_6916);
or U7311 (N_7311,N_6334,N_6792);
nand U7312 (N_7312,N_6721,N_6450);
and U7313 (N_7313,N_6135,N_6549);
nor U7314 (N_7314,N_6504,N_6717);
nand U7315 (N_7315,N_6324,N_6605);
and U7316 (N_7316,N_6746,N_6857);
xnor U7317 (N_7317,N_6406,N_6071);
xor U7318 (N_7318,N_6703,N_6845);
or U7319 (N_7319,N_6475,N_6903);
or U7320 (N_7320,N_6291,N_6258);
or U7321 (N_7321,N_6501,N_6292);
nor U7322 (N_7322,N_6893,N_6711);
or U7323 (N_7323,N_6438,N_6367);
xnor U7324 (N_7324,N_6574,N_6072);
or U7325 (N_7325,N_6325,N_6025);
and U7326 (N_7326,N_6648,N_6569);
or U7327 (N_7327,N_6222,N_6376);
or U7328 (N_7328,N_6894,N_6066);
xor U7329 (N_7329,N_6758,N_6179);
nor U7330 (N_7330,N_6127,N_6689);
nand U7331 (N_7331,N_6199,N_6461);
nor U7332 (N_7332,N_6426,N_6937);
nor U7333 (N_7333,N_6486,N_6260);
xor U7334 (N_7334,N_6518,N_6381);
nor U7335 (N_7335,N_6342,N_6914);
or U7336 (N_7336,N_6349,N_6884);
and U7337 (N_7337,N_6102,N_6380);
xor U7338 (N_7338,N_6296,N_6992);
nor U7339 (N_7339,N_6247,N_6902);
and U7340 (N_7340,N_6273,N_6686);
nand U7341 (N_7341,N_6096,N_6659);
nor U7342 (N_7342,N_6743,N_6807);
or U7343 (N_7343,N_6031,N_6243);
nand U7344 (N_7344,N_6851,N_6601);
nand U7345 (N_7345,N_6314,N_6301);
nand U7346 (N_7346,N_6238,N_6221);
and U7347 (N_7347,N_6455,N_6616);
or U7348 (N_7348,N_6657,N_6069);
nor U7349 (N_7349,N_6566,N_6939);
xnor U7350 (N_7350,N_6976,N_6266);
nor U7351 (N_7351,N_6231,N_6037);
xor U7352 (N_7352,N_6638,N_6858);
nand U7353 (N_7353,N_6760,N_6480);
and U7354 (N_7354,N_6304,N_6543);
nor U7355 (N_7355,N_6463,N_6470);
nand U7356 (N_7356,N_6702,N_6924);
or U7357 (N_7357,N_6150,N_6490);
nor U7358 (N_7358,N_6981,N_6629);
xor U7359 (N_7359,N_6958,N_6423);
nand U7360 (N_7360,N_6872,N_6878);
nand U7361 (N_7361,N_6587,N_6641);
nor U7362 (N_7362,N_6167,N_6588);
nor U7363 (N_7363,N_6811,N_6160);
or U7364 (N_7364,N_6416,N_6578);
xor U7365 (N_7365,N_6726,N_6812);
nand U7366 (N_7366,N_6906,N_6918);
xnor U7367 (N_7367,N_6158,N_6728);
nand U7368 (N_7368,N_6773,N_6797);
or U7369 (N_7369,N_6697,N_6683);
nor U7370 (N_7370,N_6469,N_6821);
and U7371 (N_7371,N_6116,N_6286);
nand U7372 (N_7372,N_6930,N_6955);
and U7373 (N_7373,N_6664,N_6765);
nand U7374 (N_7374,N_6617,N_6834);
nor U7375 (N_7375,N_6004,N_6353);
or U7376 (N_7376,N_6308,N_6404);
xor U7377 (N_7377,N_6854,N_6793);
and U7378 (N_7378,N_6068,N_6155);
nor U7379 (N_7379,N_6080,N_6484);
nor U7380 (N_7380,N_6780,N_6676);
or U7381 (N_7381,N_6724,N_6097);
xnor U7382 (N_7382,N_6337,N_6118);
or U7383 (N_7383,N_6783,N_6382);
or U7384 (N_7384,N_6751,N_6511);
xor U7385 (N_7385,N_6964,N_6994);
or U7386 (N_7386,N_6656,N_6989);
nand U7387 (N_7387,N_6151,N_6713);
nor U7388 (N_7388,N_6162,N_6644);
and U7389 (N_7389,N_6364,N_6200);
nand U7390 (N_7390,N_6545,N_6737);
and U7391 (N_7391,N_6505,N_6682);
xnor U7392 (N_7392,N_6802,N_6107);
nand U7393 (N_7393,N_6249,N_6042);
nor U7394 (N_7394,N_6056,N_6259);
nand U7395 (N_7395,N_6832,N_6088);
or U7396 (N_7396,N_6496,N_6995);
nand U7397 (N_7397,N_6632,N_6971);
nand U7398 (N_7398,N_6755,N_6022);
nor U7399 (N_7399,N_6466,N_6233);
and U7400 (N_7400,N_6752,N_6873);
nor U7401 (N_7401,N_6631,N_6383);
or U7402 (N_7402,N_6840,N_6693);
and U7403 (N_7403,N_6074,N_6063);
nor U7404 (N_7404,N_6395,N_6491);
nor U7405 (N_7405,N_6568,N_6658);
xnor U7406 (N_7406,N_6611,N_6344);
xnor U7407 (N_7407,N_6602,N_6485);
and U7408 (N_7408,N_6122,N_6253);
nand U7409 (N_7409,N_6289,N_6114);
or U7410 (N_7410,N_6223,N_6213);
xor U7411 (N_7411,N_6705,N_6168);
xnor U7412 (N_7412,N_6742,N_6668);
nor U7413 (N_7413,N_6099,N_6472);
and U7414 (N_7414,N_6882,N_6270);
xor U7415 (N_7415,N_6275,N_6073);
xnor U7416 (N_7416,N_6021,N_6552);
nand U7417 (N_7417,N_6789,N_6647);
nand U7418 (N_7418,N_6471,N_6537);
nor U7419 (N_7419,N_6660,N_6477);
or U7420 (N_7420,N_6165,N_6494);
nand U7421 (N_7421,N_6245,N_6708);
and U7422 (N_7422,N_6288,N_6877);
and U7423 (N_7423,N_6618,N_6528);
xor U7424 (N_7424,N_6396,N_6230);
xnor U7425 (N_7425,N_6209,N_6415);
or U7426 (N_7426,N_6910,N_6898);
and U7427 (N_7427,N_6440,N_6500);
and U7428 (N_7428,N_6692,N_6885);
nor U7429 (N_7429,N_6999,N_6607);
and U7430 (N_7430,N_6005,N_6909);
nand U7431 (N_7431,N_6104,N_6610);
and U7432 (N_7432,N_6112,N_6827);
and U7433 (N_7433,N_6688,N_6859);
nor U7434 (N_7434,N_6039,N_6661);
xor U7435 (N_7435,N_6443,N_6130);
nor U7436 (N_7436,N_6900,N_6919);
xor U7437 (N_7437,N_6983,N_6121);
or U7438 (N_7438,N_6143,N_6306);
or U7439 (N_7439,N_6352,N_6089);
nor U7440 (N_7440,N_6715,N_6987);
xor U7441 (N_7441,N_6002,N_6282);
nor U7442 (N_7442,N_6433,N_6855);
xor U7443 (N_7443,N_6997,N_6272);
nand U7444 (N_7444,N_6062,N_6749);
xor U7445 (N_7445,N_6284,N_6468);
or U7446 (N_7446,N_6700,N_6310);
and U7447 (N_7447,N_6948,N_6503);
xor U7448 (N_7448,N_6899,N_6538);
xnor U7449 (N_7449,N_6908,N_6698);
and U7450 (N_7450,N_6148,N_6186);
nand U7451 (N_7451,N_6988,N_6844);
nor U7452 (N_7452,N_6108,N_6799);
or U7453 (N_7453,N_6599,N_6677);
nor U7454 (N_7454,N_6962,N_6377);
or U7455 (N_7455,N_6040,N_6365);
or U7456 (N_7456,N_6166,N_6131);
nand U7457 (N_7457,N_6185,N_6595);
and U7458 (N_7458,N_6142,N_6774);
nand U7459 (N_7459,N_6830,N_6764);
or U7460 (N_7460,N_6019,N_6101);
nand U7461 (N_7461,N_6613,N_6733);
nand U7462 (N_7462,N_6033,N_6060);
and U7463 (N_7463,N_6414,N_6362);
nand U7464 (N_7464,N_6685,N_6340);
nor U7465 (N_7465,N_6871,N_6240);
and U7466 (N_7466,N_6507,N_6606);
xnor U7467 (N_7467,N_6593,N_6034);
and U7468 (N_7468,N_6550,N_6422);
nand U7469 (N_7469,N_6269,N_6038);
xor U7470 (N_7470,N_6615,N_6348);
xnor U7471 (N_7471,N_6553,N_6718);
and U7472 (N_7472,N_6264,N_6389);
xor U7473 (N_7473,N_6009,N_6279);
nor U7474 (N_7474,N_6177,N_6026);
and U7475 (N_7475,N_6612,N_6736);
nor U7476 (N_7476,N_6590,N_6531);
xor U7477 (N_7477,N_6320,N_6196);
and U7478 (N_7478,N_6345,N_6399);
and U7479 (N_7479,N_6870,N_6175);
nor U7480 (N_7480,N_6589,N_6572);
nor U7481 (N_7481,N_6219,N_6188);
or U7482 (N_7482,N_6856,N_6318);
nand U7483 (N_7483,N_6690,N_6134);
nor U7484 (N_7484,N_6242,N_6424);
nor U7485 (N_7485,N_6487,N_6157);
nand U7486 (N_7486,N_6008,N_6990);
and U7487 (N_7487,N_6144,N_6235);
xor U7488 (N_7488,N_6489,N_6841);
nand U7489 (N_7489,N_6226,N_6940);
xnor U7490 (N_7490,N_6950,N_6782);
and U7491 (N_7491,N_6850,N_6880);
and U7492 (N_7492,N_6630,N_6413);
xor U7493 (N_7493,N_6822,N_6847);
nor U7494 (N_7494,N_6126,N_6813);
xnor U7495 (N_7495,N_6285,N_6585);
nand U7496 (N_7496,N_6195,N_6754);
nor U7497 (N_7497,N_6432,N_6892);
nand U7498 (N_7498,N_6575,N_6798);
nand U7499 (N_7499,N_6077,N_6849);
and U7500 (N_7500,N_6986,N_6778);
and U7501 (N_7501,N_6483,N_6619);
nand U7502 (N_7502,N_6615,N_6790);
nand U7503 (N_7503,N_6470,N_6635);
nor U7504 (N_7504,N_6827,N_6282);
and U7505 (N_7505,N_6676,N_6782);
nand U7506 (N_7506,N_6759,N_6906);
or U7507 (N_7507,N_6130,N_6114);
or U7508 (N_7508,N_6417,N_6420);
or U7509 (N_7509,N_6636,N_6491);
nand U7510 (N_7510,N_6157,N_6566);
or U7511 (N_7511,N_6795,N_6027);
xnor U7512 (N_7512,N_6158,N_6008);
xnor U7513 (N_7513,N_6156,N_6196);
nor U7514 (N_7514,N_6391,N_6220);
or U7515 (N_7515,N_6955,N_6762);
nor U7516 (N_7516,N_6048,N_6155);
nand U7517 (N_7517,N_6603,N_6705);
and U7518 (N_7518,N_6737,N_6410);
and U7519 (N_7519,N_6266,N_6747);
xor U7520 (N_7520,N_6780,N_6516);
nor U7521 (N_7521,N_6647,N_6643);
nor U7522 (N_7522,N_6785,N_6023);
xor U7523 (N_7523,N_6677,N_6149);
nand U7524 (N_7524,N_6783,N_6883);
xor U7525 (N_7525,N_6811,N_6406);
and U7526 (N_7526,N_6646,N_6414);
and U7527 (N_7527,N_6448,N_6605);
nand U7528 (N_7528,N_6884,N_6589);
nor U7529 (N_7529,N_6759,N_6659);
xnor U7530 (N_7530,N_6245,N_6074);
or U7531 (N_7531,N_6657,N_6359);
nor U7532 (N_7532,N_6760,N_6385);
nand U7533 (N_7533,N_6502,N_6882);
xor U7534 (N_7534,N_6937,N_6801);
xor U7535 (N_7535,N_6929,N_6716);
and U7536 (N_7536,N_6926,N_6465);
or U7537 (N_7537,N_6871,N_6808);
xor U7538 (N_7538,N_6611,N_6558);
xnor U7539 (N_7539,N_6325,N_6190);
xnor U7540 (N_7540,N_6428,N_6325);
xor U7541 (N_7541,N_6382,N_6662);
nor U7542 (N_7542,N_6237,N_6006);
and U7543 (N_7543,N_6547,N_6662);
nor U7544 (N_7544,N_6113,N_6350);
xor U7545 (N_7545,N_6224,N_6141);
xnor U7546 (N_7546,N_6618,N_6940);
xor U7547 (N_7547,N_6522,N_6407);
nor U7548 (N_7548,N_6093,N_6569);
or U7549 (N_7549,N_6470,N_6703);
nand U7550 (N_7550,N_6103,N_6279);
or U7551 (N_7551,N_6803,N_6841);
nor U7552 (N_7552,N_6000,N_6043);
and U7553 (N_7553,N_6324,N_6067);
xnor U7554 (N_7554,N_6632,N_6183);
xor U7555 (N_7555,N_6692,N_6353);
and U7556 (N_7556,N_6525,N_6745);
and U7557 (N_7557,N_6969,N_6639);
nor U7558 (N_7558,N_6935,N_6585);
xnor U7559 (N_7559,N_6384,N_6323);
nor U7560 (N_7560,N_6665,N_6838);
xor U7561 (N_7561,N_6779,N_6517);
and U7562 (N_7562,N_6936,N_6497);
and U7563 (N_7563,N_6444,N_6128);
and U7564 (N_7564,N_6957,N_6490);
xnor U7565 (N_7565,N_6545,N_6677);
and U7566 (N_7566,N_6489,N_6105);
or U7567 (N_7567,N_6442,N_6949);
or U7568 (N_7568,N_6029,N_6574);
nor U7569 (N_7569,N_6606,N_6491);
nor U7570 (N_7570,N_6998,N_6480);
nand U7571 (N_7571,N_6153,N_6720);
nand U7572 (N_7572,N_6334,N_6366);
or U7573 (N_7573,N_6259,N_6787);
nor U7574 (N_7574,N_6594,N_6984);
xnor U7575 (N_7575,N_6125,N_6958);
and U7576 (N_7576,N_6437,N_6775);
nor U7577 (N_7577,N_6594,N_6566);
nand U7578 (N_7578,N_6090,N_6620);
or U7579 (N_7579,N_6851,N_6139);
nor U7580 (N_7580,N_6234,N_6281);
xor U7581 (N_7581,N_6198,N_6727);
xnor U7582 (N_7582,N_6558,N_6118);
or U7583 (N_7583,N_6364,N_6134);
nor U7584 (N_7584,N_6044,N_6966);
xnor U7585 (N_7585,N_6260,N_6413);
nor U7586 (N_7586,N_6598,N_6670);
or U7587 (N_7587,N_6882,N_6617);
nand U7588 (N_7588,N_6771,N_6615);
nand U7589 (N_7589,N_6606,N_6645);
nand U7590 (N_7590,N_6101,N_6708);
and U7591 (N_7591,N_6294,N_6299);
xnor U7592 (N_7592,N_6860,N_6718);
nor U7593 (N_7593,N_6454,N_6033);
and U7594 (N_7594,N_6118,N_6974);
and U7595 (N_7595,N_6098,N_6296);
and U7596 (N_7596,N_6686,N_6776);
nor U7597 (N_7597,N_6340,N_6896);
nor U7598 (N_7598,N_6837,N_6884);
and U7599 (N_7599,N_6066,N_6559);
xnor U7600 (N_7600,N_6198,N_6413);
xor U7601 (N_7601,N_6685,N_6856);
and U7602 (N_7602,N_6741,N_6810);
nor U7603 (N_7603,N_6818,N_6281);
nor U7604 (N_7604,N_6353,N_6761);
and U7605 (N_7605,N_6802,N_6332);
xor U7606 (N_7606,N_6880,N_6968);
and U7607 (N_7607,N_6450,N_6399);
nor U7608 (N_7608,N_6612,N_6202);
nor U7609 (N_7609,N_6321,N_6905);
xor U7610 (N_7610,N_6212,N_6708);
xnor U7611 (N_7611,N_6034,N_6027);
nand U7612 (N_7612,N_6494,N_6285);
nand U7613 (N_7613,N_6858,N_6678);
nor U7614 (N_7614,N_6863,N_6601);
xnor U7615 (N_7615,N_6599,N_6122);
and U7616 (N_7616,N_6143,N_6991);
and U7617 (N_7617,N_6420,N_6211);
nand U7618 (N_7618,N_6739,N_6806);
nor U7619 (N_7619,N_6252,N_6191);
xor U7620 (N_7620,N_6478,N_6859);
and U7621 (N_7621,N_6357,N_6571);
or U7622 (N_7622,N_6617,N_6087);
nor U7623 (N_7623,N_6744,N_6336);
nand U7624 (N_7624,N_6554,N_6442);
nor U7625 (N_7625,N_6712,N_6192);
nand U7626 (N_7626,N_6612,N_6937);
nand U7627 (N_7627,N_6905,N_6750);
nor U7628 (N_7628,N_6990,N_6932);
or U7629 (N_7629,N_6912,N_6194);
nand U7630 (N_7630,N_6681,N_6024);
nand U7631 (N_7631,N_6048,N_6272);
nand U7632 (N_7632,N_6487,N_6439);
nor U7633 (N_7633,N_6580,N_6209);
or U7634 (N_7634,N_6099,N_6813);
or U7635 (N_7635,N_6392,N_6821);
nand U7636 (N_7636,N_6941,N_6282);
or U7637 (N_7637,N_6041,N_6392);
nor U7638 (N_7638,N_6100,N_6729);
xor U7639 (N_7639,N_6230,N_6884);
xor U7640 (N_7640,N_6685,N_6169);
nand U7641 (N_7641,N_6633,N_6039);
xnor U7642 (N_7642,N_6661,N_6737);
nor U7643 (N_7643,N_6519,N_6551);
xor U7644 (N_7644,N_6609,N_6687);
nor U7645 (N_7645,N_6314,N_6282);
nor U7646 (N_7646,N_6214,N_6835);
nor U7647 (N_7647,N_6834,N_6603);
nor U7648 (N_7648,N_6356,N_6461);
nand U7649 (N_7649,N_6939,N_6610);
nor U7650 (N_7650,N_6490,N_6974);
or U7651 (N_7651,N_6079,N_6642);
nand U7652 (N_7652,N_6079,N_6248);
or U7653 (N_7653,N_6649,N_6932);
or U7654 (N_7654,N_6049,N_6713);
nand U7655 (N_7655,N_6832,N_6063);
and U7656 (N_7656,N_6151,N_6677);
and U7657 (N_7657,N_6035,N_6312);
nand U7658 (N_7658,N_6109,N_6123);
xor U7659 (N_7659,N_6960,N_6977);
nand U7660 (N_7660,N_6054,N_6779);
xnor U7661 (N_7661,N_6677,N_6346);
xor U7662 (N_7662,N_6108,N_6206);
nor U7663 (N_7663,N_6721,N_6017);
and U7664 (N_7664,N_6497,N_6110);
or U7665 (N_7665,N_6459,N_6601);
nand U7666 (N_7666,N_6206,N_6992);
xnor U7667 (N_7667,N_6127,N_6175);
and U7668 (N_7668,N_6598,N_6628);
xor U7669 (N_7669,N_6126,N_6803);
xnor U7670 (N_7670,N_6379,N_6392);
xnor U7671 (N_7671,N_6980,N_6348);
nand U7672 (N_7672,N_6687,N_6940);
or U7673 (N_7673,N_6423,N_6294);
and U7674 (N_7674,N_6455,N_6348);
nor U7675 (N_7675,N_6416,N_6708);
and U7676 (N_7676,N_6361,N_6216);
nand U7677 (N_7677,N_6560,N_6275);
or U7678 (N_7678,N_6247,N_6313);
or U7679 (N_7679,N_6998,N_6808);
xnor U7680 (N_7680,N_6701,N_6613);
or U7681 (N_7681,N_6560,N_6837);
or U7682 (N_7682,N_6858,N_6435);
and U7683 (N_7683,N_6631,N_6520);
xor U7684 (N_7684,N_6851,N_6641);
and U7685 (N_7685,N_6760,N_6800);
or U7686 (N_7686,N_6657,N_6992);
and U7687 (N_7687,N_6971,N_6818);
nor U7688 (N_7688,N_6132,N_6760);
xor U7689 (N_7689,N_6258,N_6835);
nand U7690 (N_7690,N_6731,N_6864);
nor U7691 (N_7691,N_6369,N_6206);
or U7692 (N_7692,N_6987,N_6503);
nand U7693 (N_7693,N_6256,N_6783);
xor U7694 (N_7694,N_6567,N_6201);
nor U7695 (N_7695,N_6483,N_6916);
xnor U7696 (N_7696,N_6926,N_6636);
xor U7697 (N_7697,N_6077,N_6299);
nand U7698 (N_7698,N_6435,N_6883);
nand U7699 (N_7699,N_6694,N_6808);
xnor U7700 (N_7700,N_6329,N_6832);
or U7701 (N_7701,N_6645,N_6597);
nor U7702 (N_7702,N_6765,N_6264);
xnor U7703 (N_7703,N_6664,N_6225);
and U7704 (N_7704,N_6879,N_6669);
or U7705 (N_7705,N_6622,N_6326);
or U7706 (N_7706,N_6706,N_6062);
or U7707 (N_7707,N_6641,N_6527);
xor U7708 (N_7708,N_6719,N_6554);
xor U7709 (N_7709,N_6534,N_6157);
nand U7710 (N_7710,N_6416,N_6874);
and U7711 (N_7711,N_6288,N_6361);
nor U7712 (N_7712,N_6790,N_6137);
nand U7713 (N_7713,N_6811,N_6298);
nor U7714 (N_7714,N_6765,N_6820);
and U7715 (N_7715,N_6542,N_6603);
nor U7716 (N_7716,N_6785,N_6715);
and U7717 (N_7717,N_6990,N_6254);
xnor U7718 (N_7718,N_6261,N_6215);
xor U7719 (N_7719,N_6205,N_6767);
or U7720 (N_7720,N_6768,N_6381);
or U7721 (N_7721,N_6230,N_6714);
and U7722 (N_7722,N_6243,N_6456);
nor U7723 (N_7723,N_6479,N_6385);
and U7724 (N_7724,N_6260,N_6591);
nor U7725 (N_7725,N_6478,N_6778);
or U7726 (N_7726,N_6242,N_6808);
and U7727 (N_7727,N_6895,N_6178);
or U7728 (N_7728,N_6150,N_6721);
and U7729 (N_7729,N_6252,N_6678);
and U7730 (N_7730,N_6990,N_6900);
nor U7731 (N_7731,N_6189,N_6288);
or U7732 (N_7732,N_6220,N_6481);
nand U7733 (N_7733,N_6745,N_6636);
and U7734 (N_7734,N_6376,N_6334);
nand U7735 (N_7735,N_6364,N_6464);
and U7736 (N_7736,N_6869,N_6529);
and U7737 (N_7737,N_6507,N_6146);
xor U7738 (N_7738,N_6287,N_6696);
and U7739 (N_7739,N_6059,N_6274);
nor U7740 (N_7740,N_6754,N_6291);
xor U7741 (N_7741,N_6666,N_6269);
nand U7742 (N_7742,N_6709,N_6999);
nor U7743 (N_7743,N_6409,N_6993);
xnor U7744 (N_7744,N_6236,N_6607);
nand U7745 (N_7745,N_6684,N_6892);
and U7746 (N_7746,N_6235,N_6839);
and U7747 (N_7747,N_6631,N_6651);
nor U7748 (N_7748,N_6426,N_6460);
nand U7749 (N_7749,N_6606,N_6383);
nand U7750 (N_7750,N_6951,N_6227);
and U7751 (N_7751,N_6711,N_6158);
and U7752 (N_7752,N_6872,N_6968);
nor U7753 (N_7753,N_6216,N_6053);
xor U7754 (N_7754,N_6560,N_6946);
or U7755 (N_7755,N_6518,N_6616);
xnor U7756 (N_7756,N_6927,N_6852);
xor U7757 (N_7757,N_6276,N_6316);
or U7758 (N_7758,N_6232,N_6229);
xor U7759 (N_7759,N_6012,N_6349);
or U7760 (N_7760,N_6866,N_6083);
nand U7761 (N_7761,N_6205,N_6090);
or U7762 (N_7762,N_6725,N_6592);
and U7763 (N_7763,N_6705,N_6344);
and U7764 (N_7764,N_6552,N_6915);
nand U7765 (N_7765,N_6854,N_6534);
and U7766 (N_7766,N_6748,N_6431);
and U7767 (N_7767,N_6207,N_6893);
xnor U7768 (N_7768,N_6898,N_6283);
nand U7769 (N_7769,N_6615,N_6428);
or U7770 (N_7770,N_6007,N_6526);
nor U7771 (N_7771,N_6454,N_6408);
and U7772 (N_7772,N_6427,N_6165);
and U7773 (N_7773,N_6627,N_6058);
nor U7774 (N_7774,N_6288,N_6546);
xnor U7775 (N_7775,N_6986,N_6870);
nor U7776 (N_7776,N_6012,N_6905);
nand U7777 (N_7777,N_6745,N_6897);
nor U7778 (N_7778,N_6703,N_6713);
nand U7779 (N_7779,N_6145,N_6681);
nor U7780 (N_7780,N_6131,N_6928);
and U7781 (N_7781,N_6064,N_6011);
nand U7782 (N_7782,N_6894,N_6569);
or U7783 (N_7783,N_6219,N_6746);
xnor U7784 (N_7784,N_6944,N_6752);
or U7785 (N_7785,N_6942,N_6030);
nand U7786 (N_7786,N_6968,N_6957);
nor U7787 (N_7787,N_6775,N_6287);
and U7788 (N_7788,N_6497,N_6383);
and U7789 (N_7789,N_6371,N_6630);
nand U7790 (N_7790,N_6644,N_6490);
or U7791 (N_7791,N_6172,N_6215);
or U7792 (N_7792,N_6422,N_6844);
xnor U7793 (N_7793,N_6285,N_6230);
nor U7794 (N_7794,N_6403,N_6873);
xor U7795 (N_7795,N_6611,N_6064);
and U7796 (N_7796,N_6325,N_6959);
and U7797 (N_7797,N_6616,N_6735);
and U7798 (N_7798,N_6778,N_6129);
nor U7799 (N_7799,N_6037,N_6496);
nor U7800 (N_7800,N_6516,N_6043);
xor U7801 (N_7801,N_6197,N_6285);
xnor U7802 (N_7802,N_6352,N_6525);
xnor U7803 (N_7803,N_6382,N_6216);
nor U7804 (N_7804,N_6380,N_6032);
xnor U7805 (N_7805,N_6567,N_6133);
nand U7806 (N_7806,N_6698,N_6328);
or U7807 (N_7807,N_6291,N_6784);
nand U7808 (N_7808,N_6470,N_6536);
nand U7809 (N_7809,N_6109,N_6931);
or U7810 (N_7810,N_6978,N_6961);
nand U7811 (N_7811,N_6192,N_6620);
nand U7812 (N_7812,N_6814,N_6821);
or U7813 (N_7813,N_6728,N_6234);
xor U7814 (N_7814,N_6548,N_6505);
xor U7815 (N_7815,N_6199,N_6852);
xor U7816 (N_7816,N_6688,N_6712);
nand U7817 (N_7817,N_6667,N_6285);
or U7818 (N_7818,N_6406,N_6025);
or U7819 (N_7819,N_6290,N_6218);
xnor U7820 (N_7820,N_6426,N_6231);
xor U7821 (N_7821,N_6996,N_6385);
or U7822 (N_7822,N_6009,N_6192);
and U7823 (N_7823,N_6056,N_6065);
xor U7824 (N_7824,N_6670,N_6282);
nand U7825 (N_7825,N_6191,N_6477);
and U7826 (N_7826,N_6555,N_6078);
and U7827 (N_7827,N_6346,N_6115);
nand U7828 (N_7828,N_6458,N_6738);
or U7829 (N_7829,N_6847,N_6304);
xnor U7830 (N_7830,N_6102,N_6662);
or U7831 (N_7831,N_6326,N_6641);
xnor U7832 (N_7832,N_6245,N_6317);
or U7833 (N_7833,N_6988,N_6795);
and U7834 (N_7834,N_6018,N_6944);
xnor U7835 (N_7835,N_6941,N_6010);
xnor U7836 (N_7836,N_6229,N_6606);
xnor U7837 (N_7837,N_6207,N_6652);
xnor U7838 (N_7838,N_6437,N_6570);
xor U7839 (N_7839,N_6587,N_6336);
nand U7840 (N_7840,N_6641,N_6896);
and U7841 (N_7841,N_6673,N_6643);
and U7842 (N_7842,N_6140,N_6803);
xor U7843 (N_7843,N_6421,N_6489);
nor U7844 (N_7844,N_6280,N_6241);
and U7845 (N_7845,N_6512,N_6653);
nor U7846 (N_7846,N_6104,N_6680);
or U7847 (N_7847,N_6170,N_6315);
nor U7848 (N_7848,N_6249,N_6853);
or U7849 (N_7849,N_6313,N_6646);
and U7850 (N_7850,N_6460,N_6677);
nor U7851 (N_7851,N_6441,N_6949);
nand U7852 (N_7852,N_6916,N_6709);
xor U7853 (N_7853,N_6608,N_6047);
xor U7854 (N_7854,N_6799,N_6050);
and U7855 (N_7855,N_6585,N_6964);
nor U7856 (N_7856,N_6226,N_6772);
nand U7857 (N_7857,N_6575,N_6394);
xnor U7858 (N_7858,N_6468,N_6729);
nor U7859 (N_7859,N_6284,N_6533);
or U7860 (N_7860,N_6162,N_6902);
xnor U7861 (N_7861,N_6070,N_6142);
xor U7862 (N_7862,N_6206,N_6074);
nor U7863 (N_7863,N_6150,N_6079);
xor U7864 (N_7864,N_6915,N_6885);
nand U7865 (N_7865,N_6500,N_6287);
or U7866 (N_7866,N_6155,N_6106);
or U7867 (N_7867,N_6945,N_6330);
xor U7868 (N_7868,N_6414,N_6855);
and U7869 (N_7869,N_6704,N_6253);
or U7870 (N_7870,N_6116,N_6956);
nand U7871 (N_7871,N_6688,N_6689);
nor U7872 (N_7872,N_6141,N_6683);
xor U7873 (N_7873,N_6816,N_6222);
and U7874 (N_7874,N_6114,N_6342);
or U7875 (N_7875,N_6226,N_6336);
xnor U7876 (N_7876,N_6756,N_6815);
and U7877 (N_7877,N_6505,N_6993);
or U7878 (N_7878,N_6463,N_6113);
nor U7879 (N_7879,N_6583,N_6674);
xnor U7880 (N_7880,N_6378,N_6010);
nand U7881 (N_7881,N_6581,N_6801);
and U7882 (N_7882,N_6825,N_6025);
nand U7883 (N_7883,N_6885,N_6919);
and U7884 (N_7884,N_6635,N_6467);
nor U7885 (N_7885,N_6521,N_6982);
or U7886 (N_7886,N_6649,N_6279);
nand U7887 (N_7887,N_6023,N_6381);
xor U7888 (N_7888,N_6422,N_6047);
and U7889 (N_7889,N_6331,N_6160);
xor U7890 (N_7890,N_6606,N_6265);
xor U7891 (N_7891,N_6096,N_6170);
and U7892 (N_7892,N_6832,N_6816);
nand U7893 (N_7893,N_6834,N_6091);
nand U7894 (N_7894,N_6866,N_6120);
and U7895 (N_7895,N_6216,N_6368);
nor U7896 (N_7896,N_6787,N_6090);
or U7897 (N_7897,N_6281,N_6858);
xor U7898 (N_7898,N_6827,N_6279);
nor U7899 (N_7899,N_6853,N_6490);
and U7900 (N_7900,N_6681,N_6403);
nand U7901 (N_7901,N_6047,N_6347);
nand U7902 (N_7902,N_6719,N_6109);
xnor U7903 (N_7903,N_6058,N_6435);
nand U7904 (N_7904,N_6491,N_6361);
and U7905 (N_7905,N_6536,N_6584);
xor U7906 (N_7906,N_6248,N_6032);
and U7907 (N_7907,N_6600,N_6472);
and U7908 (N_7908,N_6973,N_6598);
nand U7909 (N_7909,N_6657,N_6800);
or U7910 (N_7910,N_6887,N_6200);
nand U7911 (N_7911,N_6447,N_6269);
or U7912 (N_7912,N_6849,N_6688);
nand U7913 (N_7913,N_6066,N_6106);
or U7914 (N_7914,N_6618,N_6085);
nor U7915 (N_7915,N_6020,N_6851);
xnor U7916 (N_7916,N_6538,N_6241);
xnor U7917 (N_7917,N_6865,N_6204);
or U7918 (N_7918,N_6106,N_6609);
and U7919 (N_7919,N_6473,N_6257);
nand U7920 (N_7920,N_6312,N_6149);
nor U7921 (N_7921,N_6882,N_6880);
or U7922 (N_7922,N_6589,N_6960);
and U7923 (N_7923,N_6065,N_6215);
and U7924 (N_7924,N_6621,N_6130);
xor U7925 (N_7925,N_6155,N_6567);
or U7926 (N_7926,N_6131,N_6972);
and U7927 (N_7927,N_6757,N_6536);
or U7928 (N_7928,N_6812,N_6683);
nor U7929 (N_7929,N_6142,N_6862);
and U7930 (N_7930,N_6981,N_6662);
xor U7931 (N_7931,N_6877,N_6607);
xnor U7932 (N_7932,N_6379,N_6053);
nand U7933 (N_7933,N_6288,N_6025);
nand U7934 (N_7934,N_6884,N_6601);
or U7935 (N_7935,N_6828,N_6911);
and U7936 (N_7936,N_6804,N_6591);
xnor U7937 (N_7937,N_6055,N_6719);
nor U7938 (N_7938,N_6746,N_6186);
nor U7939 (N_7939,N_6631,N_6806);
and U7940 (N_7940,N_6123,N_6009);
nand U7941 (N_7941,N_6834,N_6421);
xor U7942 (N_7942,N_6549,N_6459);
xor U7943 (N_7943,N_6944,N_6559);
nor U7944 (N_7944,N_6902,N_6023);
nor U7945 (N_7945,N_6406,N_6492);
and U7946 (N_7946,N_6842,N_6868);
or U7947 (N_7947,N_6527,N_6887);
xnor U7948 (N_7948,N_6668,N_6361);
nand U7949 (N_7949,N_6412,N_6006);
nand U7950 (N_7950,N_6281,N_6226);
nor U7951 (N_7951,N_6711,N_6349);
or U7952 (N_7952,N_6458,N_6000);
nand U7953 (N_7953,N_6388,N_6724);
and U7954 (N_7954,N_6058,N_6407);
nand U7955 (N_7955,N_6732,N_6171);
xor U7956 (N_7956,N_6479,N_6237);
nand U7957 (N_7957,N_6436,N_6604);
nand U7958 (N_7958,N_6897,N_6508);
and U7959 (N_7959,N_6754,N_6864);
or U7960 (N_7960,N_6947,N_6911);
nor U7961 (N_7961,N_6072,N_6248);
or U7962 (N_7962,N_6251,N_6987);
nor U7963 (N_7963,N_6615,N_6140);
and U7964 (N_7964,N_6177,N_6897);
and U7965 (N_7965,N_6125,N_6067);
or U7966 (N_7966,N_6175,N_6905);
nand U7967 (N_7967,N_6464,N_6495);
and U7968 (N_7968,N_6505,N_6915);
xor U7969 (N_7969,N_6477,N_6978);
nor U7970 (N_7970,N_6400,N_6284);
or U7971 (N_7971,N_6795,N_6995);
nand U7972 (N_7972,N_6366,N_6083);
or U7973 (N_7973,N_6873,N_6779);
and U7974 (N_7974,N_6906,N_6559);
or U7975 (N_7975,N_6574,N_6648);
and U7976 (N_7976,N_6078,N_6795);
nand U7977 (N_7977,N_6546,N_6773);
nand U7978 (N_7978,N_6950,N_6319);
nor U7979 (N_7979,N_6961,N_6891);
or U7980 (N_7980,N_6912,N_6472);
nor U7981 (N_7981,N_6884,N_6239);
and U7982 (N_7982,N_6402,N_6162);
or U7983 (N_7983,N_6577,N_6432);
nand U7984 (N_7984,N_6567,N_6174);
nand U7985 (N_7985,N_6852,N_6254);
or U7986 (N_7986,N_6803,N_6821);
or U7987 (N_7987,N_6729,N_6593);
nor U7988 (N_7988,N_6210,N_6937);
xor U7989 (N_7989,N_6472,N_6339);
xor U7990 (N_7990,N_6562,N_6469);
or U7991 (N_7991,N_6050,N_6480);
nor U7992 (N_7992,N_6807,N_6197);
or U7993 (N_7993,N_6147,N_6158);
or U7994 (N_7994,N_6975,N_6864);
nand U7995 (N_7995,N_6945,N_6705);
and U7996 (N_7996,N_6840,N_6445);
xnor U7997 (N_7997,N_6770,N_6638);
and U7998 (N_7998,N_6068,N_6392);
and U7999 (N_7999,N_6617,N_6373);
nor U8000 (N_8000,N_7997,N_7221);
xor U8001 (N_8001,N_7716,N_7601);
xor U8002 (N_8002,N_7846,N_7898);
nand U8003 (N_8003,N_7240,N_7805);
xnor U8004 (N_8004,N_7752,N_7638);
xor U8005 (N_8005,N_7047,N_7529);
xnor U8006 (N_8006,N_7842,N_7011);
nand U8007 (N_8007,N_7644,N_7283);
nand U8008 (N_8008,N_7152,N_7951);
nand U8009 (N_8009,N_7564,N_7282);
nor U8010 (N_8010,N_7099,N_7685);
nand U8011 (N_8011,N_7753,N_7910);
nand U8012 (N_8012,N_7679,N_7612);
and U8013 (N_8013,N_7175,N_7156);
or U8014 (N_8014,N_7378,N_7751);
xnor U8015 (N_8015,N_7520,N_7558);
xnor U8016 (N_8016,N_7195,N_7990);
nor U8017 (N_8017,N_7700,N_7699);
nor U8018 (N_8018,N_7310,N_7109);
or U8019 (N_8019,N_7523,N_7486);
or U8020 (N_8020,N_7643,N_7742);
xnor U8021 (N_8021,N_7784,N_7304);
and U8022 (N_8022,N_7026,N_7423);
or U8023 (N_8023,N_7607,N_7112);
or U8024 (N_8024,N_7447,N_7391);
nand U8025 (N_8025,N_7858,N_7881);
or U8026 (N_8026,N_7978,N_7327);
nand U8027 (N_8027,N_7519,N_7534);
or U8028 (N_8028,N_7479,N_7583);
nand U8029 (N_8029,N_7689,N_7835);
or U8030 (N_8030,N_7884,N_7398);
and U8031 (N_8031,N_7022,N_7771);
nand U8032 (N_8032,N_7560,N_7106);
or U8033 (N_8033,N_7533,N_7933);
and U8034 (N_8034,N_7872,N_7707);
and U8035 (N_8035,N_7646,N_7375);
xnor U8036 (N_8036,N_7308,N_7614);
xor U8037 (N_8037,N_7193,N_7758);
or U8038 (N_8038,N_7900,N_7851);
and U8039 (N_8039,N_7586,N_7796);
nand U8040 (N_8040,N_7738,N_7717);
xor U8041 (N_8041,N_7843,N_7345);
or U8042 (N_8042,N_7130,N_7224);
xor U8043 (N_8043,N_7330,N_7958);
or U8044 (N_8044,N_7902,N_7246);
or U8045 (N_8045,N_7182,N_7979);
nor U8046 (N_8046,N_7487,N_7135);
or U8047 (N_8047,N_7856,N_7788);
or U8048 (N_8048,N_7138,N_7163);
and U8049 (N_8049,N_7128,N_7365);
or U8050 (N_8050,N_7739,N_7190);
and U8051 (N_8051,N_7995,N_7262);
nand U8052 (N_8052,N_7094,N_7342);
xor U8053 (N_8053,N_7313,N_7052);
and U8054 (N_8054,N_7893,N_7053);
nand U8055 (N_8055,N_7671,N_7204);
nor U8056 (N_8056,N_7168,N_7957);
and U8057 (N_8057,N_7018,N_7118);
and U8058 (N_8058,N_7265,N_7062);
nor U8059 (N_8059,N_7206,N_7007);
or U8060 (N_8060,N_7693,N_7343);
xor U8061 (N_8061,N_7129,N_7822);
nor U8062 (N_8062,N_7575,N_7297);
xor U8063 (N_8063,N_7888,N_7244);
and U8064 (N_8064,N_7291,N_7503);
nor U8065 (N_8065,N_7287,N_7861);
and U8066 (N_8066,N_7029,N_7532);
nor U8067 (N_8067,N_7115,N_7696);
and U8068 (N_8068,N_7662,N_7768);
xnor U8069 (N_8069,N_7101,N_7477);
or U8070 (N_8070,N_7478,N_7930);
xor U8071 (N_8071,N_7725,N_7513);
nand U8072 (N_8072,N_7613,N_7603);
and U8073 (N_8073,N_7501,N_7294);
nand U8074 (N_8074,N_7277,N_7966);
nand U8075 (N_8075,N_7780,N_7923);
nand U8076 (N_8076,N_7866,N_7213);
nor U8077 (N_8077,N_7499,N_7985);
nand U8078 (N_8078,N_7008,N_7386);
or U8079 (N_8079,N_7422,N_7599);
xor U8080 (N_8080,N_7453,N_7829);
nand U8081 (N_8081,N_7465,N_7761);
nor U8082 (N_8082,N_7977,N_7050);
nand U8083 (N_8083,N_7431,N_7507);
or U8084 (N_8084,N_7238,N_7383);
and U8085 (N_8085,N_7284,N_7247);
xnor U8086 (N_8086,N_7909,N_7409);
and U8087 (N_8087,N_7218,N_7415);
and U8088 (N_8088,N_7838,N_7546);
xnor U8089 (N_8089,N_7595,N_7493);
and U8090 (N_8090,N_7312,N_7773);
xnor U8091 (N_8091,N_7694,N_7432);
and U8092 (N_8092,N_7661,N_7082);
nand U8093 (N_8093,N_7426,N_7054);
or U8094 (N_8094,N_7496,N_7755);
and U8095 (N_8095,N_7637,N_7307);
and U8096 (N_8096,N_7540,N_7239);
and U8097 (N_8097,N_7719,N_7678);
xnor U8098 (N_8098,N_7883,N_7566);
nand U8099 (N_8099,N_7559,N_7639);
or U8100 (N_8100,N_7037,N_7565);
or U8101 (N_8101,N_7418,N_7046);
and U8102 (N_8102,N_7337,N_7356);
or U8103 (N_8103,N_7947,N_7808);
nand U8104 (N_8104,N_7439,N_7350);
xor U8105 (N_8105,N_7579,N_7876);
nand U8106 (N_8106,N_7381,N_7535);
or U8107 (N_8107,N_7950,N_7165);
or U8108 (N_8108,N_7669,N_7146);
xor U8109 (N_8109,N_7133,N_7681);
nand U8110 (N_8110,N_7114,N_7652);
nand U8111 (N_8111,N_7899,N_7802);
or U8112 (N_8112,N_7830,N_7172);
nor U8113 (N_8113,N_7819,N_7848);
and U8114 (N_8114,N_7061,N_7113);
xnor U8115 (N_8115,N_7056,N_7938);
nor U8116 (N_8116,N_7438,N_7273);
xnor U8117 (N_8117,N_7587,N_7770);
and U8118 (N_8118,N_7711,N_7762);
xor U8119 (N_8119,N_7740,N_7941);
nor U8120 (N_8120,N_7929,N_7927);
nand U8121 (N_8121,N_7654,N_7723);
or U8122 (N_8122,N_7442,N_7572);
nor U8123 (N_8123,N_7640,N_7359);
and U8124 (N_8124,N_7107,N_7470);
nor U8125 (N_8125,N_7994,N_7497);
or U8126 (N_8126,N_7041,N_7473);
and U8127 (N_8127,N_7173,N_7582);
or U8128 (N_8128,N_7076,N_7650);
xor U8129 (N_8129,N_7801,N_7619);
nand U8130 (N_8130,N_7731,N_7389);
and U8131 (N_8131,N_7547,N_7410);
nand U8132 (N_8132,N_7522,N_7824);
nor U8133 (N_8133,N_7746,N_7400);
xor U8134 (N_8134,N_7028,N_7139);
xnor U8135 (N_8135,N_7321,N_7598);
nand U8136 (N_8136,N_7216,N_7364);
nand U8137 (N_8137,N_7073,N_7452);
and U8138 (N_8138,N_7394,N_7539);
nor U8139 (N_8139,N_7401,N_7825);
or U8140 (N_8140,N_7136,N_7664);
and U8141 (N_8141,N_7070,N_7288);
nand U8142 (N_8142,N_7385,N_7285);
nor U8143 (N_8143,N_7594,N_7797);
nor U8144 (N_8144,N_7778,N_7592);
xnor U8145 (N_8145,N_7648,N_7715);
or U8146 (N_8146,N_7220,N_7005);
nand U8147 (N_8147,N_7404,N_7684);
xor U8148 (N_8148,N_7817,N_7406);
nor U8149 (N_8149,N_7266,N_7143);
and U8150 (N_8150,N_7710,N_7955);
nand U8151 (N_8151,N_7346,N_7148);
or U8152 (N_8152,N_7688,N_7417);
nand U8153 (N_8153,N_7176,N_7475);
or U8154 (N_8154,N_7485,N_7430);
nand U8155 (N_8155,N_7369,N_7205);
xnor U8156 (N_8156,N_7180,N_7809);
and U8157 (N_8157,N_7620,N_7363);
or U8158 (N_8158,N_7120,N_7875);
or U8159 (N_8159,N_7074,N_7628);
xnor U8160 (N_8160,N_7286,N_7034);
nand U8161 (N_8161,N_7116,N_7704);
nand U8162 (N_8162,N_7141,N_7818);
nand U8163 (N_8163,N_7948,N_7166);
nand U8164 (N_8164,N_7413,N_7293);
or U8165 (N_8165,N_7724,N_7741);
nand U8166 (N_8166,N_7623,N_7320);
nand U8167 (N_8167,N_7254,N_7090);
and U8168 (N_8168,N_7785,N_7571);
nor U8169 (N_8169,N_7806,N_7207);
nand U8170 (N_8170,N_7167,N_7542);
and U8171 (N_8171,N_7328,N_7508);
nand U8172 (N_8172,N_7014,N_7836);
nor U8173 (N_8173,N_7517,N_7857);
nor U8174 (N_8174,N_7086,N_7358);
nand U8175 (N_8175,N_7488,N_7622);
nor U8176 (N_8176,N_7084,N_7184);
and U8177 (N_8177,N_7965,N_7103);
or U8178 (N_8178,N_7943,N_7879);
nor U8179 (N_8179,N_7604,N_7713);
xor U8180 (N_8180,N_7561,N_7766);
nand U8181 (N_8181,N_7782,N_7827);
nand U8182 (N_8182,N_7241,N_7554);
and U8183 (N_8183,N_7064,N_7436);
and U8184 (N_8184,N_7949,N_7227);
or U8185 (N_8185,N_7886,N_7144);
nand U8186 (N_8186,N_7305,N_7555);
nor U8187 (N_8187,N_7874,N_7088);
xnor U8188 (N_8188,N_7589,N_7382);
xnor U8189 (N_8189,N_7556,N_7521);
nor U8190 (N_8190,N_7306,N_7392);
nand U8191 (N_8191,N_7611,N_7020);
nand U8192 (N_8192,N_7726,N_7325);
xnor U8193 (N_8193,N_7686,N_7170);
and U8194 (N_8194,N_7091,N_7980);
nor U8195 (N_8195,N_7695,N_7464);
or U8196 (N_8196,N_7706,N_7859);
xor U8197 (N_8197,N_7937,N_7961);
nand U8198 (N_8198,N_7189,N_7588);
nand U8199 (N_8199,N_7396,N_7368);
and U8200 (N_8200,N_7631,N_7104);
xnor U8201 (N_8201,N_7407,N_7016);
nor U8202 (N_8202,N_7934,N_7333);
and U8203 (N_8203,N_7576,N_7089);
or U8204 (N_8204,N_7108,N_7009);
nor U8205 (N_8205,N_7270,N_7111);
or U8206 (N_8206,N_7492,N_7887);
nand U8207 (N_8207,N_7720,N_7581);
xnor U8208 (N_8208,N_7869,N_7690);
nor U8209 (N_8209,N_7721,N_7969);
nor U8210 (N_8210,N_7373,N_7121);
and U8211 (N_8211,N_7300,N_7913);
xnor U8212 (N_8212,N_7647,N_7946);
xnor U8213 (N_8213,N_7511,N_7181);
nand U8214 (N_8214,N_7920,N_7259);
and U8215 (N_8215,N_7481,N_7811);
xnor U8216 (N_8216,N_7162,N_7360);
xor U8217 (N_8217,N_7049,N_7624);
xnor U8218 (N_8218,N_7515,N_7362);
or U8219 (N_8219,N_7341,N_7912);
or U8220 (N_8220,N_7408,N_7367);
xor U8221 (N_8221,N_7196,N_7885);
and U8222 (N_8222,N_7211,N_7735);
xnor U8223 (N_8223,N_7975,N_7323);
xnor U8224 (N_8224,N_7126,N_7353);
or U8225 (N_8225,N_7355,N_7187);
nand U8226 (N_8226,N_7380,N_7030);
and U8227 (N_8227,N_7756,N_7701);
xor U8228 (N_8228,N_7919,N_7258);
and U8229 (N_8229,N_7472,N_7440);
or U8230 (N_8230,N_7197,N_7536);
and U8231 (N_8231,N_7469,N_7907);
or U8232 (N_8232,N_7458,N_7461);
and U8233 (N_8233,N_7730,N_7823);
xor U8234 (N_8234,N_7370,N_7468);
or U8235 (N_8235,N_7889,N_7545);
nor U8236 (N_8236,N_7528,N_7970);
nand U8237 (N_8237,N_7202,N_7223);
and U8238 (N_8238,N_7451,N_7010);
and U8239 (N_8239,N_7840,N_7072);
xor U8240 (N_8240,N_7964,N_7659);
or U8241 (N_8241,N_7734,N_7845);
nor U8242 (N_8242,N_7657,N_7460);
or U8243 (N_8243,N_7524,N_7625);
and U8244 (N_8244,N_7925,N_7781);
xnor U8245 (N_8245,N_7999,N_7132);
xnor U8246 (N_8246,N_7063,N_7494);
nand U8247 (N_8247,N_7783,N_7296);
nor U8248 (N_8248,N_7489,N_7526);
nand U8249 (N_8249,N_7066,N_7550);
xor U8250 (N_8250,N_7642,N_7527);
or U8251 (N_8251,N_7618,N_7043);
or U8252 (N_8252,N_7807,N_7810);
nand U8253 (N_8253,N_7892,N_7441);
xor U8254 (N_8254,N_7236,N_7059);
nor U8255 (N_8255,N_7281,N_7656);
xor U8256 (N_8256,N_7864,N_7853);
nor U8257 (N_8257,N_7349,N_7562);
xor U8258 (N_8258,N_7702,N_7402);
or U8259 (N_8259,N_7763,N_7347);
and U8260 (N_8260,N_7931,N_7516);
xor U8261 (N_8261,N_7159,N_7267);
nor U8262 (N_8262,N_7388,N_7023);
or U8263 (N_8263,N_7145,N_7793);
nand U8264 (N_8264,N_7456,N_7484);
or U8265 (N_8265,N_7680,N_7260);
xnor U8266 (N_8266,N_7483,N_7079);
xnor U8267 (N_8267,N_7776,N_7459);
nand U8268 (N_8268,N_7935,N_7667);
nand U8269 (N_8269,N_7253,N_7414);
xnor U8270 (N_8270,N_7687,N_7606);
nand U8271 (N_8271,N_7429,N_7155);
xor U8272 (N_8272,N_7048,N_7004);
nor U8273 (N_8273,N_7655,N_7192);
or U8274 (N_8274,N_7502,N_7316);
or U8275 (N_8275,N_7445,N_7971);
xnor U8276 (N_8276,N_7868,N_7891);
nor U8277 (N_8277,N_7928,N_7901);
and U8278 (N_8278,N_7709,N_7544);
xnor U8279 (N_8279,N_7963,N_7772);
xnor U8280 (N_8280,N_7065,N_7351);
nand U8281 (N_8281,N_7134,N_7672);
and U8282 (N_8282,N_7911,N_7068);
xnor U8283 (N_8283,N_7543,N_7775);
nand U8284 (N_8284,N_7036,N_7127);
nand U8285 (N_8285,N_7003,N_7015);
nor U8286 (N_8286,N_7568,N_7040);
and U8287 (N_8287,N_7191,N_7322);
nand U8288 (N_8288,N_7303,N_7880);
xor U8289 (N_8289,N_7416,N_7377);
nor U8290 (N_8290,N_7153,N_7828);
nor U8291 (N_8291,N_7890,N_7031);
nor U8292 (N_8292,N_7666,N_7905);
xnor U8293 (N_8293,N_7627,N_7779);
nand U8294 (N_8294,N_7837,N_7674);
nand U8295 (N_8295,N_7573,N_7292);
nand U8296 (N_8296,N_7692,N_7676);
nand U8297 (N_8297,N_7530,N_7590);
xor U8298 (N_8298,N_7315,N_7744);
nor U8299 (N_8299,N_7311,N_7177);
nor U8300 (N_8300,N_7754,N_7161);
xor U8301 (N_8301,N_7737,N_7371);
and U8302 (N_8302,N_7991,N_7006);
xnor U8303 (N_8303,N_7097,N_7651);
nor U8304 (N_8304,N_7425,N_7348);
or U8305 (N_8305,N_7615,N_7832);
nor U8306 (N_8306,N_7233,N_7697);
nand U8307 (N_8307,N_7675,N_7329);
nor U8308 (N_8308,N_7448,N_7593);
nand U8309 (N_8309,N_7149,N_7945);
or U8310 (N_8310,N_7922,N_7942);
nand U8311 (N_8311,N_7727,N_7228);
xnor U8312 (N_8312,N_7201,N_7921);
xnor U8313 (N_8313,N_7765,N_7340);
or U8314 (N_8314,N_7421,N_7505);
nand U8315 (N_8315,N_7102,N_7051);
nand U8316 (N_8316,N_7915,N_7335);
nand U8317 (N_8317,N_7044,N_7634);
nand U8318 (N_8318,N_7959,N_7844);
and U8319 (N_8319,N_7736,N_7812);
nor U8320 (N_8320,N_7361,N_7215);
nand U8321 (N_8321,N_7870,N_7256);
xor U8322 (N_8322,N_7462,N_7110);
xor U8323 (N_8323,N_7552,N_7747);
xor U8324 (N_8324,N_7790,N_7854);
nand U8325 (N_8325,N_7171,N_7045);
xor U8326 (N_8326,N_7841,N_7209);
xor U8327 (N_8327,N_7179,N_7142);
nor U8328 (N_8328,N_7446,N_7981);
nand U8329 (N_8329,N_7633,N_7261);
xnor U8330 (N_8330,N_7424,N_7506);
nor U8331 (N_8331,N_7914,N_7509);
nor U8332 (N_8332,N_7903,N_7298);
xor U8333 (N_8333,N_7557,N_7339);
nand U8334 (N_8334,N_7714,N_7279);
and U8335 (N_8335,N_7248,N_7057);
nand U8336 (N_8336,N_7093,N_7140);
or U8337 (N_8337,N_7317,N_7708);
nand U8338 (N_8338,N_7855,N_7466);
and U8339 (N_8339,N_7548,N_7427);
nand U8340 (N_8340,N_7217,N_7989);
nand U8341 (N_8341,N_7663,N_7610);
xor U8342 (N_8342,N_7251,N_7013);
and U8343 (N_8343,N_7896,N_7372);
xnor U8344 (N_8344,N_7984,N_7419);
nor U8345 (N_8345,N_7393,N_7384);
and U8346 (N_8346,N_7231,N_7956);
and U8347 (N_8347,N_7275,N_7750);
and U8348 (N_8348,N_7276,N_7743);
and U8349 (N_8349,N_7636,N_7366);
nand U8350 (N_8350,N_7691,N_7397);
xor U8351 (N_8351,N_7235,N_7100);
nand U8352 (N_8352,N_7833,N_7198);
nor U8353 (N_8353,N_7973,N_7268);
nor U8354 (N_8354,N_7630,N_7147);
xor U8355 (N_8355,N_7665,N_7834);
nor U8356 (N_8356,N_7278,N_7792);
nor U8357 (N_8357,N_7498,N_7125);
xor U8358 (N_8358,N_7376,N_7677);
xnor U8359 (N_8359,N_7096,N_7081);
and U8360 (N_8360,N_7877,N_7972);
nor U8361 (N_8361,N_7718,N_7437);
or U8362 (N_8362,N_7087,N_7993);
or U8363 (N_8363,N_7476,N_7002);
nand U8364 (N_8364,N_7443,N_7490);
or U8365 (N_8365,N_7976,N_7865);
or U8366 (N_8366,N_7060,N_7234);
xor U8367 (N_8367,N_7183,N_7331);
nor U8368 (N_8368,N_7212,N_7480);
xnor U8369 (N_8369,N_7164,N_7255);
nor U8370 (N_8370,N_7174,N_7314);
nand U8371 (N_8371,N_7974,N_7225);
or U8372 (N_8372,N_7795,N_7326);
nor U8373 (N_8373,N_7653,N_7732);
nand U8374 (N_8374,N_7495,N_7577);
or U8375 (N_8375,N_7021,N_7816);
nor U8376 (N_8376,N_7237,N_7541);
or U8377 (N_8377,N_7800,N_7042);
nor U8378 (N_8378,N_7200,N_7435);
nor U8379 (N_8379,N_7878,N_7491);
xor U8380 (N_8380,N_7301,N_7374);
and U8381 (N_8381,N_7563,N_7897);
nor U8382 (N_8382,N_7621,N_7733);
xor U8383 (N_8383,N_7839,N_7597);
or U8384 (N_8384,N_7918,N_7379);
nand U8385 (N_8385,N_7596,N_7154);
and U8386 (N_8386,N_7600,N_7186);
and U8387 (N_8387,N_7185,N_7271);
xnor U8388 (N_8388,N_7789,N_7962);
or U8389 (N_8389,N_7444,N_7629);
and U8390 (N_8390,N_7263,N_7124);
nand U8391 (N_8391,N_7131,N_7119);
nand U8392 (N_8392,N_7357,N_7787);
or U8393 (N_8393,N_7698,N_7078);
or U8394 (N_8394,N_7777,N_7849);
nand U8395 (N_8395,N_7518,N_7745);
nand U8396 (N_8396,N_7616,N_7584);
xor U8397 (N_8397,N_7411,N_7803);
nand U8398 (N_8398,N_7831,N_7035);
xor U8399 (N_8399,N_7214,N_7894);
and U8400 (N_8400,N_7024,N_7757);
or U8401 (N_8401,N_7334,N_7712);
xor U8402 (N_8402,N_7944,N_7500);
or U8403 (N_8403,N_7578,N_7272);
and U8404 (N_8404,N_7525,N_7257);
xor U8405 (N_8405,N_7080,N_7917);
and U8406 (N_8406,N_7160,N_7705);
nor U8407 (N_8407,N_7463,N_7230);
or U8408 (N_8408,N_7826,N_7820);
nand U8409 (N_8409,N_7434,N_7242);
nor U8410 (N_8410,N_7570,N_7992);
xor U8411 (N_8411,N_7151,N_7814);
or U8412 (N_8412,N_7815,N_7531);
or U8413 (N_8413,N_7245,N_7067);
and U8414 (N_8414,N_7988,N_7703);
and U8415 (N_8415,N_7967,N_7908);
xnor U8416 (N_8416,N_7626,N_7774);
nand U8417 (N_8417,N_7454,N_7658);
nand U8418 (N_8418,N_7226,N_7862);
and U8419 (N_8419,N_7336,N_7580);
xnor U8420 (N_8420,N_7924,N_7038);
nor U8421 (N_8421,N_7264,N_7860);
or U8422 (N_8422,N_7998,N_7670);
nand U8423 (N_8423,N_7759,N_7514);
nor U8424 (N_8424,N_7318,N_7032);
xnor U8425 (N_8425,N_7591,N_7504);
or U8426 (N_8426,N_7538,N_7722);
nor U8427 (N_8427,N_7786,N_7605);
xnor U8428 (N_8428,N_7158,N_7055);
or U8429 (N_8429,N_7471,N_7926);
xor U8430 (N_8430,N_7169,N_7039);
xnor U8431 (N_8431,N_7895,N_7123);
xnor U8432 (N_8432,N_7764,N_7940);
xor U8433 (N_8433,N_7474,N_7660);
xnor U8434 (N_8434,N_7399,N_7728);
and U8435 (N_8435,N_7157,N_7450);
nand U8436 (N_8436,N_7309,N_7000);
and U8437 (N_8437,N_7798,N_7682);
nor U8438 (N_8438,N_7428,N_7799);
nand U8439 (N_8439,N_7332,N_7249);
and U8440 (N_8440,N_7274,N_7729);
nor U8441 (N_8441,N_7553,N_7390);
nand U8442 (N_8442,N_7295,N_7344);
nand U8443 (N_8443,N_7122,N_7092);
or U8444 (N_8444,N_7095,N_7012);
nor U8445 (N_8445,N_7512,N_7632);
or U8446 (N_8446,N_7150,N_7645);
and U8447 (N_8447,N_7804,N_7058);
nand U8448 (N_8448,N_7319,N_7290);
or U8449 (N_8449,N_7250,N_7222);
or U8450 (N_8450,N_7467,N_7852);
nor U8451 (N_8451,N_7882,N_7289);
or U8452 (N_8452,N_7210,N_7617);
and U8453 (N_8453,N_7904,N_7668);
and U8454 (N_8454,N_7873,N_7302);
and U8455 (N_8455,N_7352,N_7098);
nor U8456 (N_8456,N_7075,N_7208);
or U8457 (N_8457,N_7847,N_7968);
xor U8458 (N_8458,N_7071,N_7748);
xor U8459 (N_8459,N_7982,N_7403);
nor U8460 (N_8460,N_7791,N_7280);
nor U8461 (N_8461,N_7017,N_7549);
nand U8462 (N_8462,N_7609,N_7641);
and U8463 (N_8463,N_7537,N_7987);
and U8464 (N_8464,N_7025,N_7033);
or U8465 (N_8465,N_7585,N_7354);
nand U8466 (N_8466,N_7683,N_7871);
and U8467 (N_8467,N_7769,N_7996);
and U8468 (N_8468,N_7455,N_7324);
xnor U8469 (N_8469,N_7953,N_7203);
xor U8470 (N_8470,N_7551,N_7299);
xnor U8471 (N_8471,N_7387,N_7001);
xnor U8472 (N_8472,N_7569,N_7867);
nor U8473 (N_8473,N_7952,N_7760);
nor U8474 (N_8474,N_7821,N_7510);
nor U8475 (N_8475,N_7936,N_7960);
or U8476 (N_8476,N_7482,N_7243);
xor U8477 (N_8477,N_7083,N_7457);
and U8478 (N_8478,N_7906,N_7338);
nor U8479 (N_8479,N_7178,N_7954);
or U8480 (N_8480,N_7269,N_7749);
and U8481 (N_8481,N_7405,N_7567);
nor U8482 (N_8482,N_7105,N_7085);
xor U8483 (N_8483,N_7635,N_7449);
nor U8484 (N_8484,N_7199,N_7219);
xnor U8485 (N_8485,N_7939,N_7813);
nor U8486 (N_8486,N_7117,N_7932);
and U8487 (N_8487,N_7232,N_7019);
nand U8488 (N_8488,N_7863,N_7077);
xor U8489 (N_8489,N_7188,N_7420);
nand U8490 (N_8490,N_7850,N_7602);
nand U8491 (N_8491,N_7916,N_7794);
and U8492 (N_8492,N_7252,N_7574);
and U8493 (N_8493,N_7027,N_7069);
nor U8494 (N_8494,N_7983,N_7229);
or U8495 (N_8495,N_7137,N_7986);
nor U8496 (N_8496,N_7433,N_7395);
xnor U8497 (N_8497,N_7767,N_7194);
nor U8498 (N_8498,N_7608,N_7649);
and U8499 (N_8499,N_7412,N_7673);
xnor U8500 (N_8500,N_7505,N_7046);
nor U8501 (N_8501,N_7612,N_7335);
or U8502 (N_8502,N_7118,N_7698);
nor U8503 (N_8503,N_7122,N_7033);
nand U8504 (N_8504,N_7364,N_7538);
xor U8505 (N_8505,N_7128,N_7760);
and U8506 (N_8506,N_7927,N_7993);
xnor U8507 (N_8507,N_7934,N_7367);
nand U8508 (N_8508,N_7278,N_7339);
nor U8509 (N_8509,N_7935,N_7501);
xnor U8510 (N_8510,N_7483,N_7873);
or U8511 (N_8511,N_7349,N_7103);
or U8512 (N_8512,N_7223,N_7586);
or U8513 (N_8513,N_7768,N_7652);
nand U8514 (N_8514,N_7978,N_7923);
nand U8515 (N_8515,N_7785,N_7096);
nor U8516 (N_8516,N_7579,N_7333);
nor U8517 (N_8517,N_7391,N_7980);
or U8518 (N_8518,N_7141,N_7915);
and U8519 (N_8519,N_7887,N_7660);
xor U8520 (N_8520,N_7485,N_7086);
nor U8521 (N_8521,N_7591,N_7889);
and U8522 (N_8522,N_7935,N_7407);
or U8523 (N_8523,N_7293,N_7369);
nor U8524 (N_8524,N_7232,N_7460);
xor U8525 (N_8525,N_7144,N_7344);
nand U8526 (N_8526,N_7687,N_7501);
xor U8527 (N_8527,N_7692,N_7199);
xnor U8528 (N_8528,N_7359,N_7542);
and U8529 (N_8529,N_7426,N_7944);
nor U8530 (N_8530,N_7092,N_7112);
nand U8531 (N_8531,N_7225,N_7319);
xnor U8532 (N_8532,N_7910,N_7429);
nand U8533 (N_8533,N_7097,N_7172);
xnor U8534 (N_8534,N_7741,N_7571);
nor U8535 (N_8535,N_7011,N_7630);
and U8536 (N_8536,N_7545,N_7986);
nand U8537 (N_8537,N_7130,N_7499);
and U8538 (N_8538,N_7075,N_7859);
nor U8539 (N_8539,N_7655,N_7700);
xor U8540 (N_8540,N_7504,N_7756);
nor U8541 (N_8541,N_7459,N_7628);
nor U8542 (N_8542,N_7318,N_7028);
and U8543 (N_8543,N_7619,N_7666);
xor U8544 (N_8544,N_7810,N_7102);
nand U8545 (N_8545,N_7514,N_7167);
and U8546 (N_8546,N_7738,N_7145);
and U8547 (N_8547,N_7274,N_7564);
nor U8548 (N_8548,N_7588,N_7335);
xnor U8549 (N_8549,N_7178,N_7151);
and U8550 (N_8550,N_7258,N_7361);
xor U8551 (N_8551,N_7815,N_7116);
or U8552 (N_8552,N_7715,N_7187);
xor U8553 (N_8553,N_7236,N_7063);
nor U8554 (N_8554,N_7551,N_7302);
xnor U8555 (N_8555,N_7650,N_7073);
and U8556 (N_8556,N_7230,N_7340);
nand U8557 (N_8557,N_7566,N_7457);
or U8558 (N_8558,N_7445,N_7306);
nand U8559 (N_8559,N_7829,N_7999);
and U8560 (N_8560,N_7354,N_7753);
xnor U8561 (N_8561,N_7139,N_7790);
nand U8562 (N_8562,N_7467,N_7555);
nor U8563 (N_8563,N_7446,N_7019);
xor U8564 (N_8564,N_7440,N_7712);
and U8565 (N_8565,N_7415,N_7664);
or U8566 (N_8566,N_7574,N_7467);
and U8567 (N_8567,N_7382,N_7743);
nor U8568 (N_8568,N_7847,N_7407);
or U8569 (N_8569,N_7665,N_7736);
or U8570 (N_8570,N_7072,N_7424);
and U8571 (N_8571,N_7082,N_7702);
nor U8572 (N_8572,N_7965,N_7727);
nor U8573 (N_8573,N_7402,N_7566);
nand U8574 (N_8574,N_7555,N_7246);
nor U8575 (N_8575,N_7293,N_7090);
or U8576 (N_8576,N_7866,N_7586);
nand U8577 (N_8577,N_7611,N_7087);
nand U8578 (N_8578,N_7370,N_7772);
xor U8579 (N_8579,N_7603,N_7748);
and U8580 (N_8580,N_7496,N_7586);
nand U8581 (N_8581,N_7495,N_7543);
nand U8582 (N_8582,N_7368,N_7712);
xor U8583 (N_8583,N_7146,N_7421);
and U8584 (N_8584,N_7315,N_7420);
nand U8585 (N_8585,N_7509,N_7535);
xnor U8586 (N_8586,N_7734,N_7210);
nor U8587 (N_8587,N_7235,N_7081);
or U8588 (N_8588,N_7819,N_7143);
xor U8589 (N_8589,N_7143,N_7098);
nor U8590 (N_8590,N_7252,N_7675);
nand U8591 (N_8591,N_7012,N_7296);
xnor U8592 (N_8592,N_7117,N_7598);
xnor U8593 (N_8593,N_7171,N_7462);
nand U8594 (N_8594,N_7002,N_7560);
xor U8595 (N_8595,N_7303,N_7107);
and U8596 (N_8596,N_7224,N_7189);
xor U8597 (N_8597,N_7249,N_7066);
nor U8598 (N_8598,N_7646,N_7573);
nor U8599 (N_8599,N_7062,N_7093);
and U8600 (N_8600,N_7918,N_7488);
xnor U8601 (N_8601,N_7108,N_7440);
nand U8602 (N_8602,N_7793,N_7269);
nor U8603 (N_8603,N_7295,N_7403);
nor U8604 (N_8604,N_7145,N_7301);
or U8605 (N_8605,N_7898,N_7403);
nor U8606 (N_8606,N_7946,N_7883);
and U8607 (N_8607,N_7863,N_7267);
or U8608 (N_8608,N_7393,N_7923);
and U8609 (N_8609,N_7694,N_7699);
or U8610 (N_8610,N_7138,N_7051);
nor U8611 (N_8611,N_7264,N_7951);
or U8612 (N_8612,N_7824,N_7305);
xor U8613 (N_8613,N_7819,N_7961);
xor U8614 (N_8614,N_7851,N_7451);
or U8615 (N_8615,N_7937,N_7401);
or U8616 (N_8616,N_7388,N_7700);
or U8617 (N_8617,N_7355,N_7259);
nor U8618 (N_8618,N_7435,N_7554);
nor U8619 (N_8619,N_7518,N_7717);
and U8620 (N_8620,N_7733,N_7295);
xor U8621 (N_8621,N_7574,N_7144);
nand U8622 (N_8622,N_7293,N_7957);
nor U8623 (N_8623,N_7507,N_7248);
and U8624 (N_8624,N_7494,N_7169);
xor U8625 (N_8625,N_7412,N_7137);
nand U8626 (N_8626,N_7607,N_7554);
xnor U8627 (N_8627,N_7581,N_7366);
and U8628 (N_8628,N_7569,N_7089);
or U8629 (N_8629,N_7498,N_7088);
and U8630 (N_8630,N_7171,N_7562);
nand U8631 (N_8631,N_7874,N_7143);
and U8632 (N_8632,N_7026,N_7856);
xor U8633 (N_8633,N_7658,N_7057);
and U8634 (N_8634,N_7886,N_7522);
nand U8635 (N_8635,N_7087,N_7501);
nor U8636 (N_8636,N_7181,N_7110);
nor U8637 (N_8637,N_7534,N_7659);
and U8638 (N_8638,N_7655,N_7202);
and U8639 (N_8639,N_7121,N_7850);
nor U8640 (N_8640,N_7227,N_7998);
or U8641 (N_8641,N_7023,N_7212);
and U8642 (N_8642,N_7639,N_7820);
and U8643 (N_8643,N_7036,N_7131);
nor U8644 (N_8644,N_7518,N_7498);
xnor U8645 (N_8645,N_7978,N_7917);
or U8646 (N_8646,N_7823,N_7054);
and U8647 (N_8647,N_7397,N_7514);
nand U8648 (N_8648,N_7313,N_7956);
nand U8649 (N_8649,N_7703,N_7284);
or U8650 (N_8650,N_7328,N_7980);
nand U8651 (N_8651,N_7671,N_7905);
nand U8652 (N_8652,N_7185,N_7134);
and U8653 (N_8653,N_7840,N_7700);
nor U8654 (N_8654,N_7264,N_7751);
nor U8655 (N_8655,N_7571,N_7813);
nor U8656 (N_8656,N_7996,N_7890);
xor U8657 (N_8657,N_7276,N_7062);
nand U8658 (N_8658,N_7099,N_7297);
or U8659 (N_8659,N_7536,N_7769);
or U8660 (N_8660,N_7225,N_7622);
and U8661 (N_8661,N_7118,N_7457);
and U8662 (N_8662,N_7393,N_7974);
nand U8663 (N_8663,N_7704,N_7060);
nand U8664 (N_8664,N_7412,N_7257);
or U8665 (N_8665,N_7180,N_7174);
nor U8666 (N_8666,N_7593,N_7681);
or U8667 (N_8667,N_7154,N_7796);
and U8668 (N_8668,N_7324,N_7981);
nor U8669 (N_8669,N_7029,N_7888);
and U8670 (N_8670,N_7158,N_7977);
and U8671 (N_8671,N_7840,N_7221);
nor U8672 (N_8672,N_7657,N_7189);
xor U8673 (N_8673,N_7542,N_7725);
or U8674 (N_8674,N_7737,N_7137);
and U8675 (N_8675,N_7324,N_7360);
xor U8676 (N_8676,N_7500,N_7278);
xor U8677 (N_8677,N_7174,N_7249);
xnor U8678 (N_8678,N_7176,N_7487);
or U8679 (N_8679,N_7583,N_7222);
or U8680 (N_8680,N_7686,N_7848);
xnor U8681 (N_8681,N_7303,N_7017);
nor U8682 (N_8682,N_7730,N_7122);
or U8683 (N_8683,N_7526,N_7340);
nand U8684 (N_8684,N_7254,N_7311);
xor U8685 (N_8685,N_7636,N_7869);
nand U8686 (N_8686,N_7222,N_7096);
or U8687 (N_8687,N_7840,N_7702);
nor U8688 (N_8688,N_7743,N_7755);
nand U8689 (N_8689,N_7071,N_7954);
nand U8690 (N_8690,N_7785,N_7196);
and U8691 (N_8691,N_7890,N_7311);
nor U8692 (N_8692,N_7928,N_7545);
nor U8693 (N_8693,N_7960,N_7039);
and U8694 (N_8694,N_7818,N_7567);
nor U8695 (N_8695,N_7695,N_7927);
and U8696 (N_8696,N_7064,N_7147);
nor U8697 (N_8697,N_7850,N_7694);
or U8698 (N_8698,N_7006,N_7310);
nand U8699 (N_8699,N_7098,N_7839);
nor U8700 (N_8700,N_7088,N_7624);
nand U8701 (N_8701,N_7444,N_7523);
or U8702 (N_8702,N_7370,N_7686);
xnor U8703 (N_8703,N_7497,N_7356);
xnor U8704 (N_8704,N_7095,N_7398);
and U8705 (N_8705,N_7638,N_7107);
xnor U8706 (N_8706,N_7533,N_7750);
xor U8707 (N_8707,N_7418,N_7473);
nand U8708 (N_8708,N_7604,N_7773);
nand U8709 (N_8709,N_7159,N_7614);
nor U8710 (N_8710,N_7910,N_7018);
and U8711 (N_8711,N_7485,N_7326);
nand U8712 (N_8712,N_7088,N_7288);
nand U8713 (N_8713,N_7367,N_7292);
or U8714 (N_8714,N_7545,N_7279);
or U8715 (N_8715,N_7194,N_7835);
nor U8716 (N_8716,N_7896,N_7654);
or U8717 (N_8717,N_7242,N_7228);
or U8718 (N_8718,N_7545,N_7114);
nor U8719 (N_8719,N_7087,N_7683);
and U8720 (N_8720,N_7689,N_7030);
nand U8721 (N_8721,N_7631,N_7097);
nand U8722 (N_8722,N_7201,N_7669);
and U8723 (N_8723,N_7307,N_7533);
or U8724 (N_8724,N_7814,N_7083);
or U8725 (N_8725,N_7449,N_7687);
nor U8726 (N_8726,N_7937,N_7050);
and U8727 (N_8727,N_7219,N_7564);
or U8728 (N_8728,N_7544,N_7380);
and U8729 (N_8729,N_7843,N_7161);
or U8730 (N_8730,N_7327,N_7370);
nand U8731 (N_8731,N_7320,N_7545);
xor U8732 (N_8732,N_7417,N_7825);
nor U8733 (N_8733,N_7640,N_7242);
or U8734 (N_8734,N_7948,N_7172);
or U8735 (N_8735,N_7466,N_7810);
or U8736 (N_8736,N_7648,N_7516);
nand U8737 (N_8737,N_7633,N_7651);
xnor U8738 (N_8738,N_7747,N_7386);
xor U8739 (N_8739,N_7462,N_7816);
and U8740 (N_8740,N_7152,N_7886);
nand U8741 (N_8741,N_7526,N_7795);
or U8742 (N_8742,N_7928,N_7351);
nor U8743 (N_8743,N_7366,N_7823);
nor U8744 (N_8744,N_7151,N_7643);
nor U8745 (N_8745,N_7783,N_7733);
xor U8746 (N_8746,N_7469,N_7119);
or U8747 (N_8747,N_7688,N_7917);
nor U8748 (N_8748,N_7043,N_7040);
nor U8749 (N_8749,N_7412,N_7762);
and U8750 (N_8750,N_7000,N_7504);
xnor U8751 (N_8751,N_7776,N_7991);
or U8752 (N_8752,N_7550,N_7922);
or U8753 (N_8753,N_7508,N_7573);
xor U8754 (N_8754,N_7126,N_7159);
nor U8755 (N_8755,N_7707,N_7072);
xor U8756 (N_8756,N_7407,N_7112);
and U8757 (N_8757,N_7342,N_7463);
nor U8758 (N_8758,N_7638,N_7501);
xor U8759 (N_8759,N_7958,N_7743);
and U8760 (N_8760,N_7480,N_7113);
and U8761 (N_8761,N_7633,N_7112);
and U8762 (N_8762,N_7196,N_7178);
nor U8763 (N_8763,N_7855,N_7790);
nand U8764 (N_8764,N_7691,N_7303);
or U8765 (N_8765,N_7667,N_7231);
nand U8766 (N_8766,N_7085,N_7158);
nand U8767 (N_8767,N_7411,N_7623);
nor U8768 (N_8768,N_7574,N_7673);
or U8769 (N_8769,N_7090,N_7785);
or U8770 (N_8770,N_7750,N_7718);
and U8771 (N_8771,N_7419,N_7640);
or U8772 (N_8772,N_7845,N_7903);
nor U8773 (N_8773,N_7174,N_7346);
and U8774 (N_8774,N_7825,N_7386);
xnor U8775 (N_8775,N_7835,N_7770);
xnor U8776 (N_8776,N_7823,N_7203);
and U8777 (N_8777,N_7032,N_7523);
and U8778 (N_8778,N_7259,N_7664);
and U8779 (N_8779,N_7871,N_7429);
nor U8780 (N_8780,N_7117,N_7125);
and U8781 (N_8781,N_7798,N_7326);
nand U8782 (N_8782,N_7343,N_7674);
nor U8783 (N_8783,N_7386,N_7173);
xnor U8784 (N_8784,N_7906,N_7727);
nor U8785 (N_8785,N_7413,N_7609);
xnor U8786 (N_8786,N_7555,N_7088);
nand U8787 (N_8787,N_7295,N_7355);
or U8788 (N_8788,N_7398,N_7630);
and U8789 (N_8789,N_7392,N_7354);
and U8790 (N_8790,N_7198,N_7760);
nor U8791 (N_8791,N_7114,N_7309);
nor U8792 (N_8792,N_7226,N_7627);
xor U8793 (N_8793,N_7895,N_7839);
nand U8794 (N_8794,N_7499,N_7107);
and U8795 (N_8795,N_7866,N_7018);
or U8796 (N_8796,N_7314,N_7799);
or U8797 (N_8797,N_7341,N_7818);
or U8798 (N_8798,N_7860,N_7196);
and U8799 (N_8799,N_7747,N_7510);
nor U8800 (N_8800,N_7160,N_7839);
nand U8801 (N_8801,N_7056,N_7213);
and U8802 (N_8802,N_7839,N_7425);
xor U8803 (N_8803,N_7647,N_7153);
nand U8804 (N_8804,N_7406,N_7560);
or U8805 (N_8805,N_7055,N_7872);
xor U8806 (N_8806,N_7621,N_7782);
nor U8807 (N_8807,N_7129,N_7281);
xor U8808 (N_8808,N_7016,N_7553);
nand U8809 (N_8809,N_7365,N_7760);
nand U8810 (N_8810,N_7680,N_7716);
xnor U8811 (N_8811,N_7484,N_7678);
or U8812 (N_8812,N_7020,N_7076);
and U8813 (N_8813,N_7505,N_7122);
xnor U8814 (N_8814,N_7652,N_7950);
nor U8815 (N_8815,N_7068,N_7668);
and U8816 (N_8816,N_7857,N_7364);
xnor U8817 (N_8817,N_7791,N_7234);
nor U8818 (N_8818,N_7081,N_7241);
nand U8819 (N_8819,N_7839,N_7859);
or U8820 (N_8820,N_7522,N_7728);
or U8821 (N_8821,N_7958,N_7593);
nand U8822 (N_8822,N_7677,N_7506);
nor U8823 (N_8823,N_7220,N_7892);
nand U8824 (N_8824,N_7689,N_7177);
xor U8825 (N_8825,N_7267,N_7309);
nor U8826 (N_8826,N_7202,N_7575);
xnor U8827 (N_8827,N_7743,N_7797);
nor U8828 (N_8828,N_7980,N_7361);
and U8829 (N_8829,N_7432,N_7423);
nor U8830 (N_8830,N_7403,N_7369);
nor U8831 (N_8831,N_7057,N_7294);
xor U8832 (N_8832,N_7413,N_7793);
nor U8833 (N_8833,N_7419,N_7139);
nor U8834 (N_8834,N_7799,N_7652);
or U8835 (N_8835,N_7101,N_7281);
xnor U8836 (N_8836,N_7328,N_7218);
and U8837 (N_8837,N_7165,N_7637);
or U8838 (N_8838,N_7115,N_7570);
xnor U8839 (N_8839,N_7146,N_7812);
or U8840 (N_8840,N_7184,N_7832);
nand U8841 (N_8841,N_7970,N_7439);
xnor U8842 (N_8842,N_7007,N_7140);
nor U8843 (N_8843,N_7509,N_7059);
or U8844 (N_8844,N_7904,N_7913);
nor U8845 (N_8845,N_7221,N_7720);
nand U8846 (N_8846,N_7924,N_7855);
or U8847 (N_8847,N_7169,N_7093);
nor U8848 (N_8848,N_7196,N_7984);
nor U8849 (N_8849,N_7905,N_7945);
nand U8850 (N_8850,N_7585,N_7144);
xnor U8851 (N_8851,N_7718,N_7774);
nor U8852 (N_8852,N_7145,N_7851);
nor U8853 (N_8853,N_7674,N_7333);
xnor U8854 (N_8854,N_7303,N_7275);
xnor U8855 (N_8855,N_7043,N_7468);
nand U8856 (N_8856,N_7626,N_7845);
and U8857 (N_8857,N_7761,N_7934);
nand U8858 (N_8858,N_7970,N_7593);
nor U8859 (N_8859,N_7481,N_7757);
nor U8860 (N_8860,N_7951,N_7964);
and U8861 (N_8861,N_7189,N_7878);
xnor U8862 (N_8862,N_7388,N_7547);
and U8863 (N_8863,N_7065,N_7272);
nor U8864 (N_8864,N_7523,N_7383);
nor U8865 (N_8865,N_7146,N_7165);
nand U8866 (N_8866,N_7973,N_7472);
or U8867 (N_8867,N_7154,N_7241);
nor U8868 (N_8868,N_7625,N_7871);
and U8869 (N_8869,N_7361,N_7495);
nor U8870 (N_8870,N_7592,N_7493);
xor U8871 (N_8871,N_7333,N_7670);
nor U8872 (N_8872,N_7712,N_7396);
and U8873 (N_8873,N_7879,N_7891);
xnor U8874 (N_8874,N_7720,N_7762);
and U8875 (N_8875,N_7962,N_7178);
nor U8876 (N_8876,N_7125,N_7824);
xnor U8877 (N_8877,N_7100,N_7993);
and U8878 (N_8878,N_7745,N_7470);
and U8879 (N_8879,N_7555,N_7600);
xor U8880 (N_8880,N_7745,N_7513);
and U8881 (N_8881,N_7257,N_7839);
or U8882 (N_8882,N_7292,N_7463);
and U8883 (N_8883,N_7601,N_7183);
nand U8884 (N_8884,N_7841,N_7856);
and U8885 (N_8885,N_7922,N_7996);
or U8886 (N_8886,N_7002,N_7167);
nor U8887 (N_8887,N_7878,N_7227);
and U8888 (N_8888,N_7504,N_7876);
and U8889 (N_8889,N_7258,N_7922);
nor U8890 (N_8890,N_7179,N_7402);
xor U8891 (N_8891,N_7775,N_7592);
and U8892 (N_8892,N_7774,N_7385);
nor U8893 (N_8893,N_7924,N_7490);
nand U8894 (N_8894,N_7280,N_7443);
nor U8895 (N_8895,N_7000,N_7905);
nand U8896 (N_8896,N_7937,N_7026);
nand U8897 (N_8897,N_7186,N_7593);
nand U8898 (N_8898,N_7041,N_7404);
xnor U8899 (N_8899,N_7904,N_7021);
nand U8900 (N_8900,N_7980,N_7828);
nand U8901 (N_8901,N_7631,N_7861);
nand U8902 (N_8902,N_7135,N_7538);
nand U8903 (N_8903,N_7414,N_7993);
or U8904 (N_8904,N_7626,N_7919);
xnor U8905 (N_8905,N_7792,N_7653);
and U8906 (N_8906,N_7018,N_7270);
xnor U8907 (N_8907,N_7242,N_7589);
nand U8908 (N_8908,N_7954,N_7400);
xnor U8909 (N_8909,N_7056,N_7257);
xnor U8910 (N_8910,N_7272,N_7321);
and U8911 (N_8911,N_7278,N_7831);
nor U8912 (N_8912,N_7041,N_7352);
xor U8913 (N_8913,N_7626,N_7147);
and U8914 (N_8914,N_7907,N_7607);
and U8915 (N_8915,N_7822,N_7582);
nor U8916 (N_8916,N_7340,N_7459);
nand U8917 (N_8917,N_7805,N_7351);
or U8918 (N_8918,N_7031,N_7094);
xnor U8919 (N_8919,N_7268,N_7866);
or U8920 (N_8920,N_7426,N_7741);
nor U8921 (N_8921,N_7131,N_7691);
xnor U8922 (N_8922,N_7189,N_7758);
or U8923 (N_8923,N_7975,N_7151);
nand U8924 (N_8924,N_7902,N_7288);
nor U8925 (N_8925,N_7818,N_7422);
nor U8926 (N_8926,N_7532,N_7617);
nand U8927 (N_8927,N_7659,N_7116);
and U8928 (N_8928,N_7965,N_7589);
xor U8929 (N_8929,N_7847,N_7412);
or U8930 (N_8930,N_7363,N_7770);
nand U8931 (N_8931,N_7832,N_7888);
xor U8932 (N_8932,N_7292,N_7009);
or U8933 (N_8933,N_7102,N_7932);
xor U8934 (N_8934,N_7674,N_7643);
xor U8935 (N_8935,N_7393,N_7435);
and U8936 (N_8936,N_7499,N_7336);
nand U8937 (N_8937,N_7133,N_7542);
and U8938 (N_8938,N_7425,N_7415);
or U8939 (N_8939,N_7970,N_7505);
or U8940 (N_8940,N_7049,N_7346);
nand U8941 (N_8941,N_7610,N_7948);
or U8942 (N_8942,N_7061,N_7231);
or U8943 (N_8943,N_7091,N_7218);
nor U8944 (N_8944,N_7941,N_7149);
or U8945 (N_8945,N_7201,N_7747);
and U8946 (N_8946,N_7609,N_7349);
xnor U8947 (N_8947,N_7321,N_7970);
xnor U8948 (N_8948,N_7977,N_7854);
and U8949 (N_8949,N_7793,N_7536);
nor U8950 (N_8950,N_7738,N_7449);
nor U8951 (N_8951,N_7835,N_7731);
and U8952 (N_8952,N_7041,N_7418);
and U8953 (N_8953,N_7224,N_7079);
or U8954 (N_8954,N_7584,N_7900);
and U8955 (N_8955,N_7804,N_7671);
and U8956 (N_8956,N_7983,N_7360);
xnor U8957 (N_8957,N_7005,N_7962);
nand U8958 (N_8958,N_7953,N_7462);
nand U8959 (N_8959,N_7434,N_7233);
nand U8960 (N_8960,N_7631,N_7675);
nand U8961 (N_8961,N_7459,N_7577);
nand U8962 (N_8962,N_7200,N_7554);
or U8963 (N_8963,N_7799,N_7689);
xnor U8964 (N_8964,N_7328,N_7349);
nor U8965 (N_8965,N_7669,N_7277);
nand U8966 (N_8966,N_7339,N_7675);
nor U8967 (N_8967,N_7035,N_7335);
nand U8968 (N_8968,N_7173,N_7533);
and U8969 (N_8969,N_7898,N_7720);
nand U8970 (N_8970,N_7606,N_7794);
or U8971 (N_8971,N_7508,N_7779);
and U8972 (N_8972,N_7695,N_7297);
or U8973 (N_8973,N_7454,N_7139);
and U8974 (N_8974,N_7873,N_7713);
nand U8975 (N_8975,N_7487,N_7071);
nor U8976 (N_8976,N_7326,N_7418);
nor U8977 (N_8977,N_7704,N_7833);
xnor U8978 (N_8978,N_7966,N_7563);
nor U8979 (N_8979,N_7184,N_7309);
xnor U8980 (N_8980,N_7719,N_7619);
nor U8981 (N_8981,N_7291,N_7837);
xor U8982 (N_8982,N_7400,N_7260);
or U8983 (N_8983,N_7228,N_7142);
xnor U8984 (N_8984,N_7092,N_7986);
xor U8985 (N_8985,N_7791,N_7681);
nand U8986 (N_8986,N_7904,N_7403);
xor U8987 (N_8987,N_7723,N_7381);
nand U8988 (N_8988,N_7825,N_7021);
nand U8989 (N_8989,N_7798,N_7292);
xor U8990 (N_8990,N_7743,N_7777);
or U8991 (N_8991,N_7168,N_7507);
and U8992 (N_8992,N_7313,N_7610);
nand U8993 (N_8993,N_7647,N_7346);
nand U8994 (N_8994,N_7543,N_7392);
nor U8995 (N_8995,N_7997,N_7946);
nand U8996 (N_8996,N_7310,N_7703);
nand U8997 (N_8997,N_7780,N_7589);
nor U8998 (N_8998,N_7924,N_7306);
or U8999 (N_8999,N_7809,N_7103);
nand U9000 (N_9000,N_8258,N_8982);
nand U9001 (N_9001,N_8841,N_8035);
and U9002 (N_9002,N_8657,N_8522);
or U9003 (N_9003,N_8094,N_8741);
nand U9004 (N_9004,N_8224,N_8276);
nor U9005 (N_9005,N_8429,N_8550);
or U9006 (N_9006,N_8484,N_8973);
nor U9007 (N_9007,N_8130,N_8318);
xnor U9008 (N_9008,N_8166,N_8197);
nand U9009 (N_9009,N_8064,N_8553);
xor U9010 (N_9010,N_8976,N_8746);
or U9011 (N_9011,N_8145,N_8005);
nand U9012 (N_9012,N_8415,N_8950);
nor U9013 (N_9013,N_8901,N_8398);
nor U9014 (N_9014,N_8394,N_8709);
xnor U9015 (N_9015,N_8567,N_8155);
or U9016 (N_9016,N_8316,N_8960);
or U9017 (N_9017,N_8821,N_8171);
nand U9018 (N_9018,N_8311,N_8674);
nand U9019 (N_9019,N_8201,N_8246);
and U9020 (N_9020,N_8534,N_8921);
nand U9021 (N_9021,N_8693,N_8981);
nand U9022 (N_9022,N_8274,N_8896);
xor U9023 (N_9023,N_8230,N_8541);
nor U9024 (N_9024,N_8615,N_8302);
nand U9025 (N_9025,N_8334,N_8793);
xnor U9026 (N_9026,N_8372,N_8272);
and U9027 (N_9027,N_8473,N_8235);
xnor U9028 (N_9028,N_8255,N_8962);
xor U9029 (N_9029,N_8771,N_8571);
nor U9030 (N_9030,N_8149,N_8373);
and U9031 (N_9031,N_8468,N_8944);
xor U9032 (N_9032,N_8706,N_8381);
or U9033 (N_9033,N_8117,N_8486);
nand U9034 (N_9034,N_8238,N_8600);
and U9035 (N_9035,N_8937,N_8399);
and U9036 (N_9036,N_8009,N_8996);
and U9037 (N_9037,N_8879,N_8025);
nor U9038 (N_9038,N_8717,N_8384);
and U9039 (N_9039,N_8846,N_8371);
nor U9040 (N_9040,N_8152,N_8379);
and U9041 (N_9041,N_8714,N_8294);
and U9042 (N_9042,N_8237,N_8652);
and U9043 (N_9043,N_8998,N_8927);
nand U9044 (N_9044,N_8199,N_8519);
nor U9045 (N_9045,N_8071,N_8857);
nand U9046 (N_9046,N_8252,N_8408);
nand U9047 (N_9047,N_8417,N_8396);
or U9048 (N_9048,N_8114,N_8864);
and U9049 (N_9049,N_8990,N_8698);
nor U9050 (N_9050,N_8032,N_8491);
or U9051 (N_9051,N_8087,N_8466);
nor U9052 (N_9052,N_8104,N_8858);
or U9053 (N_9053,N_8557,N_8953);
or U9054 (N_9054,N_8301,N_8449);
or U9055 (N_9055,N_8203,N_8605);
nor U9056 (N_9056,N_8556,N_8049);
nor U9057 (N_9057,N_8721,N_8632);
or U9058 (N_9058,N_8216,N_8697);
xor U9059 (N_9059,N_8143,N_8227);
nor U9060 (N_9060,N_8346,N_8897);
or U9061 (N_9061,N_8213,N_8492);
nor U9062 (N_9062,N_8254,N_8456);
nor U9063 (N_9063,N_8343,N_8631);
and U9064 (N_9064,N_8447,N_8759);
or U9065 (N_9065,N_8813,N_8137);
xor U9066 (N_9066,N_8963,N_8552);
nand U9067 (N_9067,N_8917,N_8115);
nor U9068 (N_9068,N_8961,N_8193);
or U9069 (N_9069,N_8423,N_8840);
nand U9070 (N_9070,N_8716,N_8363);
and U9071 (N_9071,N_8367,N_8579);
or U9072 (N_9072,N_8377,N_8044);
xnor U9073 (N_9073,N_8738,N_8414);
nand U9074 (N_9074,N_8477,N_8894);
xnor U9075 (N_9075,N_8956,N_8620);
nor U9076 (N_9076,N_8649,N_8271);
xor U9077 (N_9077,N_8482,N_8058);
and U9078 (N_9078,N_8220,N_8125);
nor U9079 (N_9079,N_8419,N_8782);
or U9080 (N_9080,N_8008,N_8368);
xor U9081 (N_9081,N_8979,N_8562);
and U9082 (N_9082,N_8000,N_8893);
nor U9083 (N_9083,N_8431,N_8899);
nor U9084 (N_9084,N_8861,N_8862);
and U9085 (N_9085,N_8184,N_8083);
nand U9086 (N_9086,N_8845,N_8980);
xor U9087 (N_9087,N_8226,N_8544);
nor U9088 (N_9088,N_8671,N_8450);
nor U9089 (N_9089,N_8779,N_8691);
or U9090 (N_9090,N_8539,N_8860);
or U9091 (N_9091,N_8890,N_8121);
nand U9092 (N_9092,N_8656,N_8867);
nor U9093 (N_9093,N_8364,N_8452);
and U9094 (N_9094,N_8543,N_8688);
xnor U9095 (N_9095,N_8509,N_8554);
and U9096 (N_9096,N_8968,N_8244);
nor U9097 (N_9097,N_8595,N_8403);
and U9098 (N_9098,N_8333,N_8215);
or U9099 (N_9099,N_8922,N_8163);
or U9100 (N_9100,N_8733,N_8358);
or U9101 (N_9101,N_8475,N_8854);
xor U9102 (N_9102,N_8624,N_8514);
or U9103 (N_9103,N_8745,N_8504);
and U9104 (N_9104,N_8382,N_8683);
or U9105 (N_9105,N_8096,N_8353);
nand U9106 (N_9106,N_8167,N_8080);
nand U9107 (N_9107,N_8128,N_8762);
or U9108 (N_9108,N_8843,N_8742);
xor U9109 (N_9109,N_8329,N_8764);
and U9110 (N_9110,N_8587,N_8659);
or U9111 (N_9111,N_8866,N_8014);
nor U9112 (N_9112,N_8200,N_8964);
nand U9113 (N_9113,N_8208,N_8780);
and U9114 (N_9114,N_8040,N_8942);
and U9115 (N_9115,N_8977,N_8725);
nor U9116 (N_9116,N_8261,N_8891);
xor U9117 (N_9117,N_8066,N_8995);
or U9118 (N_9118,N_8033,N_8701);
xor U9119 (N_9119,N_8004,N_8744);
xor U9120 (N_9120,N_8672,N_8202);
xor U9121 (N_9121,N_8775,N_8795);
nand U9122 (N_9122,N_8485,N_8387);
or U9123 (N_9123,N_8880,N_8139);
xnor U9124 (N_9124,N_8703,N_8434);
xor U9125 (N_9125,N_8747,N_8713);
xnor U9126 (N_9126,N_8234,N_8401);
xnor U9127 (N_9127,N_8106,N_8283);
or U9128 (N_9128,N_8676,N_8502);
nor U9129 (N_9129,N_8673,N_8132);
nor U9130 (N_9130,N_8270,N_8259);
nor U9131 (N_9131,N_8530,N_8506);
nand U9132 (N_9132,N_8275,N_8548);
xor U9133 (N_9133,N_8489,N_8832);
or U9134 (N_9134,N_8940,N_8777);
and U9135 (N_9135,N_8931,N_8818);
xnor U9136 (N_9136,N_8889,N_8195);
xnor U9137 (N_9137,N_8680,N_8206);
nor U9138 (N_9138,N_8257,N_8625);
xor U9139 (N_9139,N_8663,N_8116);
or U9140 (N_9140,N_8061,N_8189);
xor U9141 (N_9141,N_8805,N_8919);
xnor U9142 (N_9142,N_8908,N_8952);
and U9143 (N_9143,N_8273,N_8635);
nand U9144 (N_9144,N_8001,N_8490);
and U9145 (N_9145,N_8611,N_8930);
or U9146 (N_9146,N_8729,N_8225);
and U9147 (N_9147,N_8570,N_8397);
and U9148 (N_9148,N_8679,N_8469);
xnor U9149 (N_9149,N_8675,N_8898);
xor U9150 (N_9150,N_8056,N_8198);
nor U9151 (N_9151,N_8465,N_8699);
and U9152 (N_9152,N_8321,N_8036);
nand U9153 (N_9153,N_8427,N_8422);
nand U9154 (N_9154,N_8722,N_8281);
nor U9155 (N_9155,N_8409,N_8822);
xnor U9156 (N_9156,N_8849,N_8402);
or U9157 (N_9157,N_8936,N_8410);
nand U9158 (N_9158,N_8618,N_8268);
nand U9159 (N_9159,N_8161,N_8041);
nor U9160 (N_9160,N_8970,N_8411);
and U9161 (N_9161,N_8480,N_8141);
nor U9162 (N_9162,N_8781,N_8914);
or U9163 (N_9163,N_8053,N_8310);
xnor U9164 (N_9164,N_8778,N_8006);
or U9165 (N_9165,N_8994,N_8516);
and U9166 (N_9166,N_8695,N_8753);
nand U9167 (N_9167,N_8169,N_8178);
and U9168 (N_9168,N_8535,N_8501);
xnor U9169 (N_9169,N_8819,N_8391);
and U9170 (N_9170,N_8007,N_8655);
nor U9171 (N_9171,N_8266,N_8926);
nand U9172 (N_9172,N_8378,N_8694);
xnor U9173 (N_9173,N_8988,N_8075);
nor U9174 (N_9174,N_8023,N_8015);
nand U9175 (N_9175,N_8118,N_8765);
or U9176 (N_9176,N_8324,N_8959);
and U9177 (N_9177,N_8016,N_8205);
nor U9178 (N_9178,N_8702,N_8856);
and U9179 (N_9179,N_8609,N_8574);
nor U9180 (N_9180,N_8907,N_8572);
xnor U9181 (N_9181,N_8873,N_8545);
nand U9182 (N_9182,N_8568,N_8481);
and U9183 (N_9183,N_8325,N_8222);
or U9184 (N_9184,N_8877,N_8135);
and U9185 (N_9185,N_8351,N_8050);
nor U9186 (N_9186,N_8551,N_8507);
nor U9187 (N_9187,N_8223,N_8749);
or U9188 (N_9188,N_8774,N_8677);
xor U9189 (N_9189,N_8724,N_8369);
and U9190 (N_9190,N_8344,N_8278);
xor U9191 (N_9191,N_8499,N_8847);
xnor U9192 (N_9192,N_8848,N_8581);
nand U9193 (N_9193,N_8971,N_8515);
nor U9194 (N_9194,N_8686,N_8194);
or U9195 (N_9195,N_8370,N_8026);
xor U9196 (N_9196,N_8168,N_8298);
and U9197 (N_9197,N_8123,N_8599);
nor U9198 (N_9198,N_8458,N_8374);
xor U9199 (N_9199,N_8425,N_8002);
nand U9200 (N_9200,N_8718,N_8958);
or U9201 (N_9201,N_8186,N_8185);
nor U9202 (N_9202,N_8527,N_8508);
xnor U9203 (N_9203,N_8256,N_8766);
nand U9204 (N_9204,N_8433,N_8196);
xnor U9205 (N_9205,N_8089,N_8662);
nand U9206 (N_9206,N_8459,N_8945);
nand U9207 (N_9207,N_8086,N_8732);
or U9208 (N_9208,N_8210,N_8987);
nor U9209 (N_9209,N_8120,N_8623);
and U9210 (N_9210,N_8380,N_8350);
xor U9211 (N_9211,N_8664,N_8003);
and U9212 (N_9212,N_8560,N_8634);
nand U9213 (N_9213,N_8451,N_8510);
or U9214 (N_9214,N_8838,N_8851);
and U9215 (N_9215,N_8991,N_8156);
and U9216 (N_9216,N_8740,N_8455);
nand U9217 (N_9217,N_8159,N_8192);
and U9218 (N_9218,N_8647,N_8601);
and U9219 (N_9219,N_8020,N_8844);
and U9220 (N_9220,N_8191,N_8101);
or U9221 (N_9221,N_8768,N_8179);
or U9222 (N_9222,N_8021,N_8072);
and U9223 (N_9223,N_8284,N_8412);
or U9224 (N_9224,N_8790,N_8954);
nor U9225 (N_9225,N_8047,N_8886);
or U9226 (N_9226,N_8214,N_8165);
or U9227 (N_9227,N_8517,N_8883);
nor U9228 (N_9228,N_8918,N_8109);
nor U9229 (N_9229,N_8288,N_8591);
nor U9230 (N_9230,N_8669,N_8651);
or U9231 (N_9231,N_8407,N_8144);
or U9232 (N_9232,N_8218,N_8794);
nand U9233 (N_9233,N_8267,N_8339);
or U9234 (N_9234,N_8943,N_8127);
or U9235 (N_9235,N_8063,N_8426);
and U9236 (N_9236,N_8999,N_8293);
xnor U9237 (N_9237,N_8947,N_8354);
or U9238 (N_9238,N_8483,N_8390);
or U9239 (N_9239,N_8682,N_8079);
nand U9240 (N_9240,N_8577,N_8046);
nand U9241 (N_9241,N_8839,N_8934);
or U9242 (N_9242,N_8176,N_8105);
or U9243 (N_9243,N_8816,N_8592);
nor U9244 (N_9244,N_8785,N_8019);
or U9245 (N_9245,N_8984,N_8667);
nor U9246 (N_9246,N_8362,N_8823);
nor U9247 (N_9247,N_8523,N_8102);
nor U9248 (N_9248,N_8707,N_8013);
xor U9249 (N_9249,N_8340,N_8209);
nand U9250 (N_9250,N_8438,N_8457);
nand U9251 (N_9251,N_8436,N_8405);
nor U9252 (N_9252,N_8467,N_8606);
or U9253 (N_9253,N_8935,N_8453);
and U9254 (N_9254,N_8424,N_8232);
nor U9255 (N_9255,N_8309,N_8524);
nor U9256 (N_9256,N_8824,N_8319);
xor U9257 (N_9257,N_8594,N_8685);
nand U9258 (N_9258,N_8582,N_8641);
xor U9259 (N_9259,N_8588,N_8360);
nand U9260 (N_9260,N_8734,N_8151);
nor U9261 (N_9261,N_8913,N_8630);
xnor U9262 (N_9262,N_8231,N_8590);
nor U9263 (N_9263,N_8797,N_8689);
nor U9264 (N_9264,N_8498,N_8924);
nand U9265 (N_9265,N_8332,N_8241);
nand U9266 (N_9266,N_8126,N_8039);
or U9267 (N_9267,N_8090,N_8787);
xor U9268 (N_9268,N_8286,N_8077);
nor U9269 (N_9269,N_8204,N_8737);
nor U9270 (N_9270,N_8989,N_8831);
nand U9271 (N_9271,N_8906,N_8487);
xor U9272 (N_9272,N_8726,N_8900);
and U9273 (N_9273,N_8603,N_8108);
and U9274 (N_9274,N_8700,N_8948);
and U9275 (N_9275,N_8463,N_8495);
xor U9276 (N_9276,N_8345,N_8388);
and U9277 (N_9277,N_8692,N_8376);
xor U9278 (N_9278,N_8583,N_8789);
xnor U9279 (N_9279,N_8538,N_8140);
xor U9280 (N_9280,N_8068,N_8060);
nand U9281 (N_9281,N_8826,N_8095);
or U9282 (N_9282,N_8796,N_8251);
and U9283 (N_9283,N_8070,N_8113);
or U9284 (N_9284,N_8142,N_8758);
xor U9285 (N_9285,N_8313,N_8555);
xor U9286 (N_9286,N_8250,N_8341);
and U9287 (N_9287,N_8828,N_8735);
nor U9288 (N_9288,N_8312,N_8347);
and U9289 (N_9289,N_8925,N_8279);
and U9290 (N_9290,N_8532,N_8331);
and U9291 (N_9291,N_8157,N_8756);
and U9292 (N_9292,N_8119,N_8236);
or U9293 (N_9293,N_8442,N_8057);
or U9294 (N_9294,N_8177,N_8661);
xnor U9295 (N_9295,N_8690,N_8091);
nand U9296 (N_9296,N_8640,N_8598);
and U9297 (N_9297,N_8616,N_8285);
nor U9298 (N_9298,N_8349,N_8696);
and U9299 (N_9299,N_8739,N_8932);
nand U9300 (N_9300,N_8359,N_8802);
xnor U9301 (N_9301,N_8027,N_8134);
nor U9302 (N_9302,N_8546,N_8180);
nand U9303 (N_9303,N_8472,N_8011);
nor U9304 (N_9304,N_8646,N_8761);
xor U9305 (N_9305,N_8129,N_8645);
xor U9306 (N_9306,N_8814,N_8566);
xnor U9307 (N_9307,N_8642,N_8788);
or U9308 (N_9308,N_8299,N_8972);
or U9309 (N_9309,N_8949,N_8051);
xor U9310 (N_9310,N_8065,N_8540);
nand U9311 (N_9311,N_8076,N_8461);
nand U9312 (N_9312,N_8708,N_8307);
nor U9313 (N_9313,N_8911,N_8978);
nand U9314 (N_9314,N_8607,N_8470);
nor U9315 (N_9315,N_8356,N_8799);
nor U9316 (N_9316,N_8637,N_8355);
and U9317 (N_9317,N_8443,N_8092);
and U9318 (N_9318,N_8772,N_8705);
nor U9319 (N_9319,N_8786,N_8993);
xor U9320 (N_9320,N_8808,N_8612);
and U9321 (N_9321,N_8903,N_8062);
nand U9322 (N_9322,N_8967,N_8245);
nor U9323 (N_9323,N_8892,N_8549);
and U9324 (N_9324,N_8803,N_8493);
xnor U9325 (N_9325,N_8448,N_8392);
xnor U9326 (N_9326,N_8029,N_8754);
or U9327 (N_9327,N_8228,N_8097);
nand U9328 (N_9328,N_8093,N_8289);
and U9329 (N_9329,N_8654,N_8136);
nor U9330 (N_9330,N_8253,N_8357);
or U9331 (N_9331,N_8648,N_8160);
nor U9332 (N_9332,N_8174,N_8644);
or U9333 (N_9333,N_8314,N_8593);
xor U9334 (N_9334,N_8247,N_8017);
nor U9335 (N_9335,N_8670,N_8336);
nor U9336 (N_9336,N_8404,N_8773);
nor U9337 (N_9337,N_8445,N_8511);
xor U9338 (N_9338,N_8992,N_8711);
xor U9339 (N_9339,N_8327,N_8084);
nand U9340 (N_9340,N_8505,N_8798);
and U9341 (N_9341,N_8526,N_8100);
nor U9342 (N_9342,N_8454,N_8054);
or U9343 (N_9343,N_8352,N_8164);
nor U9344 (N_9344,N_8939,N_8441);
and U9345 (N_9345,N_8881,N_8986);
xnor U9346 (N_9346,N_8815,N_8966);
nor U9347 (N_9347,N_8767,N_8052);
or U9348 (N_9348,N_8763,N_8525);
and U9349 (N_9349,N_8059,N_8938);
nor U9350 (N_9350,N_8290,N_8030);
nand U9351 (N_9351,N_8326,N_8162);
and U9352 (N_9352,N_8099,N_8969);
nor U9353 (N_9353,N_8619,N_8338);
xnor U9354 (N_9354,N_8576,N_8531);
nor U9355 (N_9355,N_8811,N_8175);
and U9356 (N_9356,N_8687,N_8211);
xor U9357 (N_9357,N_8809,N_8723);
or U9358 (N_9358,N_8614,N_8478);
or U9359 (N_9359,N_8704,N_8865);
xnor U9360 (N_9360,N_8869,N_8138);
nor U9361 (N_9361,N_8946,N_8666);
nor U9362 (N_9362,N_8172,N_8416);
nand U9363 (N_9363,N_8081,N_8277);
xor U9364 (N_9364,N_8755,N_8905);
nand U9365 (N_9365,N_8750,N_8916);
or U9366 (N_9366,N_8018,N_8190);
nor U9367 (N_9367,N_8269,N_8784);
nand U9368 (N_9368,N_8112,N_8024);
nor U9369 (N_9369,N_8439,N_8400);
xnor U9370 (N_9370,N_8678,N_8280);
and U9371 (N_9371,N_8150,N_8503);
xnor U9372 (N_9372,N_8558,N_8859);
or U9373 (N_9373,N_8428,N_8533);
nor U9374 (N_9374,N_8348,N_8320);
xnor U9375 (N_9375,N_8010,N_8863);
and U9376 (N_9376,N_8884,N_8957);
and U9377 (N_9377,N_8330,N_8833);
nand U9378 (N_9378,N_8770,N_8807);
nand U9379 (N_9379,N_8148,N_8328);
nand U9380 (N_9380,N_8836,N_8188);
or U9381 (N_9381,N_8520,N_8835);
nor U9382 (N_9382,N_8239,N_8496);
and U9383 (N_9383,N_8263,N_8103);
nor U9384 (N_9384,N_8069,N_8233);
nor U9385 (N_9385,N_8633,N_8107);
or U9386 (N_9386,N_8791,N_8752);
nand U9387 (N_9387,N_8306,N_8537);
and U9388 (N_9388,N_8170,N_8181);
and U9389 (N_9389,N_8585,N_8643);
xor U9390 (N_9390,N_8034,N_8604);
xnor U9391 (N_9391,N_8561,N_8776);
or U9392 (N_9392,N_8668,N_8337);
and U9393 (N_9393,N_8375,N_8660);
and U9394 (N_9394,N_8296,N_8406);
xor U9395 (N_9395,N_8923,N_8315);
nor U9396 (N_9396,N_8710,N_8929);
nand U9397 (N_9397,N_8420,N_8748);
nand U9398 (N_9398,N_8085,N_8596);
nand U9399 (N_9399,N_8915,N_8751);
nand U9400 (N_9400,N_8681,N_8440);
xor U9401 (N_9401,N_8389,N_8575);
and U9402 (N_9402,N_8626,N_8810);
xnor U9403 (N_9403,N_8622,N_8804);
nor U9404 (N_9404,N_8872,N_8565);
nand U9405 (N_9405,N_8757,N_8895);
nand U9406 (N_9406,N_8719,N_8262);
or U9407 (N_9407,N_8146,N_8037);
xnor U9408 (N_9408,N_8240,N_8042);
nor U9409 (N_9409,N_8207,N_8650);
and U9410 (N_9410,N_8882,N_8476);
and U9411 (N_9411,N_8852,N_8413);
nand U9412 (N_9412,N_8529,N_8474);
and U9413 (N_9413,N_8303,N_8249);
and U9414 (N_9414,N_8528,N_8855);
and U9415 (N_9415,N_8665,N_8088);
or U9416 (N_9416,N_8627,N_8183);
nor U9417 (N_9417,N_8243,N_8124);
and U9418 (N_9418,N_8743,N_8783);
and U9419 (N_9419,N_8361,N_8073);
xor U9420 (N_9420,N_8653,N_8827);
xnor U9421 (N_9421,N_8038,N_8928);
and U9422 (N_9422,N_8820,N_8264);
or U9423 (N_9423,N_8153,N_8837);
xnor U9424 (N_9424,N_8613,N_8830);
nor U9425 (N_9425,N_8715,N_8887);
and U9426 (N_9426,N_8658,N_8187);
nand U9427 (N_9427,N_8573,N_8684);
xnor U9428 (N_9428,N_8727,N_8983);
nand U9429 (N_9429,N_8217,N_8536);
nand U9430 (N_9430,N_8421,N_8385);
xnor U9431 (N_9431,N_8965,N_8974);
nand U9432 (N_9432,N_8817,N_8564);
nand U9433 (N_9433,N_8559,N_8728);
and U9434 (N_9434,N_8850,N_8444);
xor U9435 (N_9435,N_8464,N_8806);
or U9436 (N_9436,N_8513,N_8242);
nand U9437 (N_9437,N_8586,N_8610);
nor U9438 (N_9438,N_8323,N_8386);
xor U9439 (N_9439,N_8497,N_8292);
nor U9440 (N_9440,N_8304,N_8951);
nor U9441 (N_9441,N_8910,N_8074);
nor U9442 (N_9442,N_8584,N_8874);
and U9443 (N_9443,N_8342,N_8393);
xnor U9444 (N_9444,N_8888,N_8048);
nand U9445 (N_9445,N_8580,N_8569);
nand U9446 (N_9446,N_8521,N_8801);
xor U9447 (N_9447,N_8933,N_8628);
or U9448 (N_9448,N_8997,N_8825);
nand U9449 (N_9449,N_8909,N_8043);
xnor U9450 (N_9450,N_8300,N_8158);
nor U9451 (N_9451,N_8985,N_8173);
xnor U9452 (N_9452,N_8366,N_8078);
and U9453 (N_9453,N_8031,N_8853);
or U9454 (N_9454,N_8287,N_8547);
or U9455 (N_9455,N_8730,N_8110);
or U9456 (N_9456,N_8720,N_8395);
nand U9457 (N_9457,N_8518,N_8608);
nand U9458 (N_9458,N_8941,N_8418);
or U9459 (N_9459,N_8902,N_8636);
nor U9460 (N_9460,N_8028,N_8920);
and U9461 (N_9461,N_8563,N_8462);
xor U9462 (N_9462,N_8597,N_8868);
and U9463 (N_9463,N_8870,N_8512);
nor U9464 (N_9464,N_8383,N_8067);
xnor U9465 (N_9465,N_8842,N_8147);
or U9466 (N_9466,N_8297,N_8494);
and U9467 (N_9467,N_8308,N_8871);
nor U9468 (N_9468,N_8133,N_8446);
or U9469 (N_9469,N_8365,N_8282);
or U9470 (N_9470,N_8955,N_8212);
and U9471 (N_9471,N_8435,N_8479);
nor U9472 (N_9472,N_8229,N_8792);
or U9473 (N_9473,N_8639,N_8432);
nor U9474 (N_9474,N_8437,N_8834);
and U9475 (N_9475,N_8430,N_8295);
or U9476 (N_9476,N_8221,N_8800);
or U9477 (N_9477,N_8317,N_8736);
nand U9478 (N_9478,N_8975,N_8602);
nor U9479 (N_9479,N_8291,N_8878);
nor U9480 (N_9480,N_8629,N_8621);
xor U9481 (N_9481,N_8912,N_8638);
xor U9482 (N_9482,N_8885,N_8022);
nor U9483 (N_9483,N_8322,N_8012);
or U9484 (N_9484,N_8248,N_8617);
nand U9485 (N_9485,N_8578,N_8904);
and U9486 (N_9486,N_8111,N_8098);
and U9487 (N_9487,N_8812,N_8876);
xor U9488 (N_9488,N_8712,N_8335);
or U9489 (N_9489,N_8875,N_8260);
xor U9490 (N_9490,N_8829,N_8219);
and U9491 (N_9491,N_8769,N_8082);
and U9492 (N_9492,N_8488,N_8265);
and U9493 (N_9493,N_8154,N_8045);
nand U9494 (N_9494,N_8471,N_8305);
nor U9495 (N_9495,N_8760,N_8182);
and U9496 (N_9496,N_8122,N_8500);
or U9497 (N_9497,N_8055,N_8731);
and U9498 (N_9498,N_8542,N_8460);
nor U9499 (N_9499,N_8589,N_8131);
nor U9500 (N_9500,N_8871,N_8682);
and U9501 (N_9501,N_8478,N_8677);
or U9502 (N_9502,N_8456,N_8725);
xor U9503 (N_9503,N_8801,N_8334);
xor U9504 (N_9504,N_8469,N_8481);
or U9505 (N_9505,N_8103,N_8670);
or U9506 (N_9506,N_8483,N_8896);
or U9507 (N_9507,N_8116,N_8247);
and U9508 (N_9508,N_8576,N_8079);
xor U9509 (N_9509,N_8823,N_8506);
and U9510 (N_9510,N_8769,N_8623);
xor U9511 (N_9511,N_8642,N_8723);
or U9512 (N_9512,N_8929,N_8063);
nor U9513 (N_9513,N_8799,N_8958);
nand U9514 (N_9514,N_8614,N_8183);
or U9515 (N_9515,N_8616,N_8840);
nand U9516 (N_9516,N_8152,N_8965);
xnor U9517 (N_9517,N_8257,N_8769);
nor U9518 (N_9518,N_8219,N_8256);
nor U9519 (N_9519,N_8752,N_8647);
xor U9520 (N_9520,N_8171,N_8240);
or U9521 (N_9521,N_8371,N_8650);
xor U9522 (N_9522,N_8275,N_8243);
nand U9523 (N_9523,N_8631,N_8409);
xnor U9524 (N_9524,N_8585,N_8484);
or U9525 (N_9525,N_8316,N_8146);
nor U9526 (N_9526,N_8460,N_8198);
and U9527 (N_9527,N_8795,N_8038);
nand U9528 (N_9528,N_8276,N_8910);
xor U9529 (N_9529,N_8072,N_8536);
xnor U9530 (N_9530,N_8831,N_8437);
and U9531 (N_9531,N_8809,N_8248);
or U9532 (N_9532,N_8596,N_8333);
xor U9533 (N_9533,N_8452,N_8013);
nor U9534 (N_9534,N_8511,N_8382);
nor U9535 (N_9535,N_8766,N_8009);
and U9536 (N_9536,N_8820,N_8028);
nor U9537 (N_9537,N_8057,N_8654);
nand U9538 (N_9538,N_8684,N_8259);
and U9539 (N_9539,N_8374,N_8936);
and U9540 (N_9540,N_8300,N_8615);
nand U9541 (N_9541,N_8124,N_8301);
or U9542 (N_9542,N_8032,N_8634);
xnor U9543 (N_9543,N_8086,N_8197);
and U9544 (N_9544,N_8463,N_8535);
and U9545 (N_9545,N_8528,N_8567);
nor U9546 (N_9546,N_8095,N_8972);
and U9547 (N_9547,N_8673,N_8909);
and U9548 (N_9548,N_8332,N_8773);
and U9549 (N_9549,N_8547,N_8203);
nor U9550 (N_9550,N_8046,N_8852);
xnor U9551 (N_9551,N_8567,N_8363);
and U9552 (N_9552,N_8281,N_8770);
xnor U9553 (N_9553,N_8564,N_8504);
nand U9554 (N_9554,N_8833,N_8983);
nor U9555 (N_9555,N_8455,N_8424);
and U9556 (N_9556,N_8686,N_8237);
or U9557 (N_9557,N_8467,N_8991);
nand U9558 (N_9558,N_8324,N_8641);
xor U9559 (N_9559,N_8547,N_8564);
xnor U9560 (N_9560,N_8642,N_8698);
xor U9561 (N_9561,N_8501,N_8872);
nand U9562 (N_9562,N_8485,N_8913);
nand U9563 (N_9563,N_8331,N_8436);
nand U9564 (N_9564,N_8380,N_8348);
nor U9565 (N_9565,N_8320,N_8276);
nand U9566 (N_9566,N_8077,N_8432);
and U9567 (N_9567,N_8492,N_8999);
and U9568 (N_9568,N_8455,N_8553);
nand U9569 (N_9569,N_8025,N_8413);
nand U9570 (N_9570,N_8417,N_8884);
and U9571 (N_9571,N_8442,N_8761);
xnor U9572 (N_9572,N_8137,N_8669);
or U9573 (N_9573,N_8171,N_8572);
or U9574 (N_9574,N_8060,N_8152);
nor U9575 (N_9575,N_8419,N_8647);
xnor U9576 (N_9576,N_8637,N_8668);
xor U9577 (N_9577,N_8713,N_8704);
nand U9578 (N_9578,N_8403,N_8334);
nor U9579 (N_9579,N_8122,N_8388);
and U9580 (N_9580,N_8933,N_8673);
nor U9581 (N_9581,N_8556,N_8070);
and U9582 (N_9582,N_8565,N_8989);
or U9583 (N_9583,N_8483,N_8106);
nand U9584 (N_9584,N_8435,N_8004);
xor U9585 (N_9585,N_8015,N_8712);
or U9586 (N_9586,N_8589,N_8166);
and U9587 (N_9587,N_8924,N_8653);
or U9588 (N_9588,N_8706,N_8497);
xnor U9589 (N_9589,N_8989,N_8327);
nor U9590 (N_9590,N_8406,N_8386);
nor U9591 (N_9591,N_8830,N_8521);
and U9592 (N_9592,N_8184,N_8622);
nor U9593 (N_9593,N_8011,N_8021);
nand U9594 (N_9594,N_8129,N_8236);
or U9595 (N_9595,N_8032,N_8802);
or U9596 (N_9596,N_8641,N_8960);
xnor U9597 (N_9597,N_8817,N_8472);
xor U9598 (N_9598,N_8115,N_8759);
and U9599 (N_9599,N_8532,N_8023);
nand U9600 (N_9600,N_8114,N_8667);
nand U9601 (N_9601,N_8215,N_8756);
nand U9602 (N_9602,N_8534,N_8018);
and U9603 (N_9603,N_8315,N_8373);
nand U9604 (N_9604,N_8790,N_8599);
nand U9605 (N_9605,N_8918,N_8102);
or U9606 (N_9606,N_8209,N_8756);
nand U9607 (N_9607,N_8226,N_8716);
nor U9608 (N_9608,N_8898,N_8329);
and U9609 (N_9609,N_8327,N_8447);
nor U9610 (N_9610,N_8770,N_8701);
and U9611 (N_9611,N_8032,N_8642);
nor U9612 (N_9612,N_8639,N_8864);
or U9613 (N_9613,N_8070,N_8723);
xnor U9614 (N_9614,N_8842,N_8665);
nand U9615 (N_9615,N_8011,N_8532);
nor U9616 (N_9616,N_8803,N_8210);
or U9617 (N_9617,N_8806,N_8765);
and U9618 (N_9618,N_8691,N_8585);
nand U9619 (N_9619,N_8473,N_8942);
and U9620 (N_9620,N_8122,N_8499);
or U9621 (N_9621,N_8228,N_8415);
or U9622 (N_9622,N_8368,N_8672);
and U9623 (N_9623,N_8777,N_8938);
nand U9624 (N_9624,N_8688,N_8888);
or U9625 (N_9625,N_8418,N_8498);
nand U9626 (N_9626,N_8935,N_8784);
xnor U9627 (N_9627,N_8636,N_8961);
or U9628 (N_9628,N_8875,N_8438);
xnor U9629 (N_9629,N_8585,N_8775);
xnor U9630 (N_9630,N_8459,N_8075);
nand U9631 (N_9631,N_8764,N_8158);
nor U9632 (N_9632,N_8784,N_8417);
or U9633 (N_9633,N_8645,N_8387);
nand U9634 (N_9634,N_8293,N_8802);
and U9635 (N_9635,N_8859,N_8129);
and U9636 (N_9636,N_8682,N_8844);
and U9637 (N_9637,N_8156,N_8196);
nor U9638 (N_9638,N_8995,N_8114);
and U9639 (N_9639,N_8532,N_8354);
xnor U9640 (N_9640,N_8484,N_8390);
or U9641 (N_9641,N_8375,N_8625);
nor U9642 (N_9642,N_8469,N_8964);
xnor U9643 (N_9643,N_8761,N_8239);
and U9644 (N_9644,N_8006,N_8905);
and U9645 (N_9645,N_8131,N_8695);
nor U9646 (N_9646,N_8518,N_8029);
and U9647 (N_9647,N_8383,N_8969);
or U9648 (N_9648,N_8771,N_8878);
or U9649 (N_9649,N_8764,N_8150);
and U9650 (N_9650,N_8317,N_8755);
and U9651 (N_9651,N_8616,N_8224);
nor U9652 (N_9652,N_8040,N_8547);
or U9653 (N_9653,N_8885,N_8928);
or U9654 (N_9654,N_8215,N_8954);
nand U9655 (N_9655,N_8076,N_8734);
and U9656 (N_9656,N_8426,N_8390);
xor U9657 (N_9657,N_8110,N_8457);
nor U9658 (N_9658,N_8549,N_8915);
nor U9659 (N_9659,N_8338,N_8785);
and U9660 (N_9660,N_8435,N_8283);
or U9661 (N_9661,N_8179,N_8625);
or U9662 (N_9662,N_8480,N_8670);
nor U9663 (N_9663,N_8067,N_8464);
nor U9664 (N_9664,N_8239,N_8098);
nor U9665 (N_9665,N_8629,N_8246);
nand U9666 (N_9666,N_8614,N_8413);
nor U9667 (N_9667,N_8726,N_8268);
and U9668 (N_9668,N_8686,N_8584);
or U9669 (N_9669,N_8601,N_8758);
and U9670 (N_9670,N_8181,N_8876);
and U9671 (N_9671,N_8651,N_8955);
or U9672 (N_9672,N_8931,N_8353);
nand U9673 (N_9673,N_8321,N_8265);
or U9674 (N_9674,N_8575,N_8374);
or U9675 (N_9675,N_8308,N_8931);
or U9676 (N_9676,N_8368,N_8946);
nand U9677 (N_9677,N_8214,N_8570);
xor U9678 (N_9678,N_8812,N_8218);
or U9679 (N_9679,N_8350,N_8343);
or U9680 (N_9680,N_8356,N_8954);
nor U9681 (N_9681,N_8464,N_8980);
and U9682 (N_9682,N_8367,N_8500);
nor U9683 (N_9683,N_8276,N_8959);
xor U9684 (N_9684,N_8738,N_8157);
xnor U9685 (N_9685,N_8930,N_8385);
or U9686 (N_9686,N_8486,N_8283);
and U9687 (N_9687,N_8729,N_8810);
xor U9688 (N_9688,N_8042,N_8554);
xnor U9689 (N_9689,N_8666,N_8691);
xor U9690 (N_9690,N_8933,N_8097);
or U9691 (N_9691,N_8992,N_8969);
or U9692 (N_9692,N_8641,N_8543);
and U9693 (N_9693,N_8107,N_8526);
nor U9694 (N_9694,N_8886,N_8032);
or U9695 (N_9695,N_8794,N_8156);
nand U9696 (N_9696,N_8272,N_8999);
and U9697 (N_9697,N_8574,N_8613);
nor U9698 (N_9698,N_8578,N_8399);
and U9699 (N_9699,N_8390,N_8626);
and U9700 (N_9700,N_8304,N_8827);
nand U9701 (N_9701,N_8627,N_8690);
and U9702 (N_9702,N_8875,N_8995);
xor U9703 (N_9703,N_8049,N_8131);
or U9704 (N_9704,N_8884,N_8922);
xnor U9705 (N_9705,N_8406,N_8323);
or U9706 (N_9706,N_8416,N_8701);
nand U9707 (N_9707,N_8304,N_8588);
nand U9708 (N_9708,N_8707,N_8381);
xor U9709 (N_9709,N_8883,N_8051);
and U9710 (N_9710,N_8931,N_8076);
and U9711 (N_9711,N_8219,N_8583);
nand U9712 (N_9712,N_8831,N_8372);
or U9713 (N_9713,N_8622,N_8407);
or U9714 (N_9714,N_8453,N_8732);
and U9715 (N_9715,N_8601,N_8155);
nor U9716 (N_9716,N_8219,N_8393);
nand U9717 (N_9717,N_8057,N_8567);
or U9718 (N_9718,N_8819,N_8577);
and U9719 (N_9719,N_8567,N_8407);
nand U9720 (N_9720,N_8927,N_8658);
xor U9721 (N_9721,N_8458,N_8912);
nor U9722 (N_9722,N_8822,N_8753);
xor U9723 (N_9723,N_8287,N_8899);
and U9724 (N_9724,N_8087,N_8720);
nand U9725 (N_9725,N_8994,N_8251);
nand U9726 (N_9726,N_8113,N_8857);
nor U9727 (N_9727,N_8187,N_8455);
xnor U9728 (N_9728,N_8549,N_8873);
nor U9729 (N_9729,N_8324,N_8765);
or U9730 (N_9730,N_8355,N_8795);
nor U9731 (N_9731,N_8677,N_8959);
and U9732 (N_9732,N_8026,N_8166);
xnor U9733 (N_9733,N_8627,N_8804);
nand U9734 (N_9734,N_8515,N_8757);
or U9735 (N_9735,N_8755,N_8011);
nand U9736 (N_9736,N_8584,N_8915);
xor U9737 (N_9737,N_8248,N_8586);
nand U9738 (N_9738,N_8362,N_8875);
nand U9739 (N_9739,N_8630,N_8118);
nor U9740 (N_9740,N_8468,N_8630);
or U9741 (N_9741,N_8220,N_8273);
or U9742 (N_9742,N_8899,N_8224);
or U9743 (N_9743,N_8542,N_8820);
xnor U9744 (N_9744,N_8590,N_8809);
and U9745 (N_9745,N_8350,N_8480);
and U9746 (N_9746,N_8028,N_8974);
nor U9747 (N_9747,N_8679,N_8717);
nand U9748 (N_9748,N_8124,N_8708);
nand U9749 (N_9749,N_8791,N_8238);
nor U9750 (N_9750,N_8418,N_8403);
or U9751 (N_9751,N_8693,N_8866);
nor U9752 (N_9752,N_8136,N_8343);
nor U9753 (N_9753,N_8805,N_8290);
and U9754 (N_9754,N_8853,N_8923);
or U9755 (N_9755,N_8928,N_8849);
nor U9756 (N_9756,N_8165,N_8537);
or U9757 (N_9757,N_8678,N_8680);
or U9758 (N_9758,N_8861,N_8540);
and U9759 (N_9759,N_8009,N_8286);
nor U9760 (N_9760,N_8402,N_8524);
or U9761 (N_9761,N_8984,N_8264);
nand U9762 (N_9762,N_8687,N_8353);
nor U9763 (N_9763,N_8090,N_8667);
nand U9764 (N_9764,N_8858,N_8427);
nand U9765 (N_9765,N_8024,N_8584);
xnor U9766 (N_9766,N_8215,N_8266);
nor U9767 (N_9767,N_8554,N_8320);
nor U9768 (N_9768,N_8780,N_8774);
nor U9769 (N_9769,N_8503,N_8481);
nor U9770 (N_9770,N_8149,N_8252);
xnor U9771 (N_9771,N_8981,N_8998);
xor U9772 (N_9772,N_8070,N_8601);
xor U9773 (N_9773,N_8111,N_8496);
or U9774 (N_9774,N_8693,N_8280);
xor U9775 (N_9775,N_8229,N_8819);
xnor U9776 (N_9776,N_8654,N_8630);
and U9777 (N_9777,N_8926,N_8352);
nor U9778 (N_9778,N_8533,N_8712);
or U9779 (N_9779,N_8951,N_8223);
nor U9780 (N_9780,N_8508,N_8350);
or U9781 (N_9781,N_8746,N_8361);
xnor U9782 (N_9782,N_8030,N_8213);
nand U9783 (N_9783,N_8712,N_8478);
or U9784 (N_9784,N_8035,N_8133);
xnor U9785 (N_9785,N_8966,N_8711);
nand U9786 (N_9786,N_8742,N_8701);
nand U9787 (N_9787,N_8986,N_8666);
and U9788 (N_9788,N_8384,N_8450);
and U9789 (N_9789,N_8291,N_8225);
nor U9790 (N_9790,N_8721,N_8143);
xor U9791 (N_9791,N_8457,N_8914);
nand U9792 (N_9792,N_8815,N_8527);
and U9793 (N_9793,N_8949,N_8193);
or U9794 (N_9794,N_8220,N_8487);
or U9795 (N_9795,N_8978,N_8946);
or U9796 (N_9796,N_8084,N_8492);
nand U9797 (N_9797,N_8741,N_8281);
nor U9798 (N_9798,N_8816,N_8649);
nand U9799 (N_9799,N_8934,N_8462);
and U9800 (N_9800,N_8825,N_8381);
and U9801 (N_9801,N_8501,N_8668);
nor U9802 (N_9802,N_8663,N_8061);
or U9803 (N_9803,N_8918,N_8549);
nand U9804 (N_9804,N_8857,N_8282);
nand U9805 (N_9805,N_8441,N_8566);
nand U9806 (N_9806,N_8449,N_8615);
or U9807 (N_9807,N_8949,N_8002);
and U9808 (N_9808,N_8129,N_8529);
nand U9809 (N_9809,N_8819,N_8698);
nand U9810 (N_9810,N_8278,N_8581);
nor U9811 (N_9811,N_8288,N_8743);
or U9812 (N_9812,N_8994,N_8381);
nand U9813 (N_9813,N_8713,N_8267);
xnor U9814 (N_9814,N_8726,N_8609);
and U9815 (N_9815,N_8267,N_8122);
nor U9816 (N_9816,N_8566,N_8986);
nor U9817 (N_9817,N_8852,N_8206);
and U9818 (N_9818,N_8853,N_8206);
nand U9819 (N_9819,N_8868,N_8461);
nand U9820 (N_9820,N_8470,N_8669);
nand U9821 (N_9821,N_8971,N_8770);
xor U9822 (N_9822,N_8142,N_8864);
xnor U9823 (N_9823,N_8270,N_8613);
nor U9824 (N_9824,N_8204,N_8325);
xnor U9825 (N_9825,N_8391,N_8885);
nand U9826 (N_9826,N_8843,N_8837);
nand U9827 (N_9827,N_8909,N_8260);
and U9828 (N_9828,N_8066,N_8263);
nor U9829 (N_9829,N_8214,N_8699);
nand U9830 (N_9830,N_8220,N_8056);
or U9831 (N_9831,N_8610,N_8092);
or U9832 (N_9832,N_8876,N_8452);
xnor U9833 (N_9833,N_8487,N_8403);
xnor U9834 (N_9834,N_8373,N_8712);
or U9835 (N_9835,N_8591,N_8480);
or U9836 (N_9836,N_8736,N_8610);
xor U9837 (N_9837,N_8694,N_8965);
or U9838 (N_9838,N_8154,N_8883);
xor U9839 (N_9839,N_8591,N_8132);
xor U9840 (N_9840,N_8546,N_8129);
or U9841 (N_9841,N_8346,N_8994);
and U9842 (N_9842,N_8727,N_8360);
nand U9843 (N_9843,N_8858,N_8822);
xor U9844 (N_9844,N_8256,N_8875);
nand U9845 (N_9845,N_8116,N_8165);
xor U9846 (N_9846,N_8362,N_8423);
and U9847 (N_9847,N_8763,N_8337);
and U9848 (N_9848,N_8985,N_8296);
or U9849 (N_9849,N_8357,N_8422);
and U9850 (N_9850,N_8369,N_8426);
or U9851 (N_9851,N_8566,N_8420);
nor U9852 (N_9852,N_8119,N_8375);
nand U9853 (N_9853,N_8339,N_8177);
nand U9854 (N_9854,N_8370,N_8630);
nand U9855 (N_9855,N_8694,N_8549);
nand U9856 (N_9856,N_8551,N_8940);
or U9857 (N_9857,N_8101,N_8854);
nor U9858 (N_9858,N_8394,N_8260);
xnor U9859 (N_9859,N_8987,N_8209);
nor U9860 (N_9860,N_8201,N_8305);
nand U9861 (N_9861,N_8861,N_8175);
nand U9862 (N_9862,N_8084,N_8349);
and U9863 (N_9863,N_8752,N_8952);
or U9864 (N_9864,N_8586,N_8630);
and U9865 (N_9865,N_8761,N_8064);
nand U9866 (N_9866,N_8286,N_8357);
and U9867 (N_9867,N_8659,N_8497);
nand U9868 (N_9868,N_8091,N_8365);
nand U9869 (N_9869,N_8460,N_8092);
xor U9870 (N_9870,N_8783,N_8770);
and U9871 (N_9871,N_8094,N_8598);
xor U9872 (N_9872,N_8824,N_8842);
or U9873 (N_9873,N_8109,N_8348);
nand U9874 (N_9874,N_8428,N_8350);
nor U9875 (N_9875,N_8186,N_8721);
nand U9876 (N_9876,N_8872,N_8558);
xor U9877 (N_9877,N_8341,N_8578);
nand U9878 (N_9878,N_8968,N_8351);
and U9879 (N_9879,N_8341,N_8060);
nand U9880 (N_9880,N_8137,N_8204);
and U9881 (N_9881,N_8407,N_8101);
nor U9882 (N_9882,N_8786,N_8230);
nand U9883 (N_9883,N_8367,N_8451);
nand U9884 (N_9884,N_8776,N_8184);
and U9885 (N_9885,N_8666,N_8166);
xnor U9886 (N_9886,N_8131,N_8819);
or U9887 (N_9887,N_8438,N_8686);
nand U9888 (N_9888,N_8514,N_8178);
or U9889 (N_9889,N_8714,N_8084);
nand U9890 (N_9890,N_8306,N_8451);
xor U9891 (N_9891,N_8156,N_8042);
nor U9892 (N_9892,N_8870,N_8916);
xnor U9893 (N_9893,N_8025,N_8756);
and U9894 (N_9894,N_8082,N_8059);
xor U9895 (N_9895,N_8058,N_8911);
nand U9896 (N_9896,N_8176,N_8376);
xor U9897 (N_9897,N_8156,N_8858);
nand U9898 (N_9898,N_8989,N_8002);
nand U9899 (N_9899,N_8679,N_8130);
nor U9900 (N_9900,N_8157,N_8547);
nand U9901 (N_9901,N_8626,N_8850);
and U9902 (N_9902,N_8552,N_8254);
nand U9903 (N_9903,N_8286,N_8729);
nor U9904 (N_9904,N_8394,N_8462);
or U9905 (N_9905,N_8323,N_8724);
nand U9906 (N_9906,N_8607,N_8696);
xor U9907 (N_9907,N_8420,N_8297);
xor U9908 (N_9908,N_8674,N_8030);
nor U9909 (N_9909,N_8358,N_8493);
nand U9910 (N_9910,N_8327,N_8899);
xnor U9911 (N_9911,N_8362,N_8224);
nor U9912 (N_9912,N_8422,N_8355);
nand U9913 (N_9913,N_8662,N_8729);
nand U9914 (N_9914,N_8338,N_8068);
nor U9915 (N_9915,N_8770,N_8031);
nor U9916 (N_9916,N_8115,N_8702);
and U9917 (N_9917,N_8588,N_8621);
nand U9918 (N_9918,N_8413,N_8796);
xnor U9919 (N_9919,N_8634,N_8358);
or U9920 (N_9920,N_8166,N_8357);
xnor U9921 (N_9921,N_8581,N_8444);
xnor U9922 (N_9922,N_8386,N_8555);
xnor U9923 (N_9923,N_8597,N_8962);
xor U9924 (N_9924,N_8090,N_8342);
nand U9925 (N_9925,N_8233,N_8863);
or U9926 (N_9926,N_8053,N_8209);
nor U9927 (N_9927,N_8271,N_8614);
nand U9928 (N_9928,N_8392,N_8933);
nand U9929 (N_9929,N_8462,N_8308);
or U9930 (N_9930,N_8368,N_8436);
or U9931 (N_9931,N_8711,N_8722);
nand U9932 (N_9932,N_8499,N_8224);
and U9933 (N_9933,N_8254,N_8928);
xor U9934 (N_9934,N_8828,N_8931);
nor U9935 (N_9935,N_8039,N_8153);
xor U9936 (N_9936,N_8016,N_8705);
nor U9937 (N_9937,N_8737,N_8165);
nor U9938 (N_9938,N_8357,N_8295);
nand U9939 (N_9939,N_8560,N_8111);
and U9940 (N_9940,N_8487,N_8451);
nor U9941 (N_9941,N_8868,N_8093);
and U9942 (N_9942,N_8397,N_8884);
and U9943 (N_9943,N_8468,N_8795);
xnor U9944 (N_9944,N_8572,N_8050);
and U9945 (N_9945,N_8757,N_8267);
xnor U9946 (N_9946,N_8626,N_8953);
nand U9947 (N_9947,N_8059,N_8856);
xnor U9948 (N_9948,N_8595,N_8100);
nand U9949 (N_9949,N_8072,N_8332);
and U9950 (N_9950,N_8296,N_8731);
xnor U9951 (N_9951,N_8989,N_8721);
and U9952 (N_9952,N_8182,N_8632);
nor U9953 (N_9953,N_8180,N_8933);
and U9954 (N_9954,N_8222,N_8108);
or U9955 (N_9955,N_8094,N_8257);
or U9956 (N_9956,N_8315,N_8692);
nand U9957 (N_9957,N_8787,N_8194);
xnor U9958 (N_9958,N_8967,N_8244);
or U9959 (N_9959,N_8776,N_8826);
and U9960 (N_9960,N_8248,N_8087);
nor U9961 (N_9961,N_8325,N_8054);
or U9962 (N_9962,N_8938,N_8782);
and U9963 (N_9963,N_8677,N_8340);
and U9964 (N_9964,N_8033,N_8453);
nand U9965 (N_9965,N_8240,N_8211);
and U9966 (N_9966,N_8477,N_8008);
nor U9967 (N_9967,N_8460,N_8140);
xor U9968 (N_9968,N_8401,N_8930);
nor U9969 (N_9969,N_8199,N_8138);
nand U9970 (N_9970,N_8751,N_8204);
nor U9971 (N_9971,N_8939,N_8701);
nor U9972 (N_9972,N_8993,N_8401);
or U9973 (N_9973,N_8352,N_8371);
or U9974 (N_9974,N_8300,N_8258);
xnor U9975 (N_9975,N_8846,N_8011);
nand U9976 (N_9976,N_8903,N_8130);
or U9977 (N_9977,N_8804,N_8523);
xor U9978 (N_9978,N_8713,N_8537);
nand U9979 (N_9979,N_8481,N_8255);
nand U9980 (N_9980,N_8373,N_8683);
xnor U9981 (N_9981,N_8785,N_8153);
nand U9982 (N_9982,N_8218,N_8431);
nand U9983 (N_9983,N_8504,N_8824);
or U9984 (N_9984,N_8806,N_8203);
xor U9985 (N_9985,N_8122,N_8843);
nand U9986 (N_9986,N_8008,N_8241);
or U9987 (N_9987,N_8053,N_8765);
xnor U9988 (N_9988,N_8177,N_8241);
and U9989 (N_9989,N_8387,N_8404);
nor U9990 (N_9990,N_8066,N_8145);
nor U9991 (N_9991,N_8856,N_8466);
or U9992 (N_9992,N_8086,N_8399);
nor U9993 (N_9993,N_8679,N_8511);
xor U9994 (N_9994,N_8169,N_8214);
nor U9995 (N_9995,N_8098,N_8758);
and U9996 (N_9996,N_8448,N_8037);
nand U9997 (N_9997,N_8134,N_8249);
and U9998 (N_9998,N_8479,N_8321);
and U9999 (N_9999,N_8066,N_8094);
nand U10000 (N_10000,N_9929,N_9725);
xor U10001 (N_10001,N_9705,N_9057);
nand U10002 (N_10002,N_9569,N_9495);
nor U10003 (N_10003,N_9861,N_9145);
xor U10004 (N_10004,N_9825,N_9496);
or U10005 (N_10005,N_9524,N_9322);
nand U10006 (N_10006,N_9081,N_9656);
or U10007 (N_10007,N_9367,N_9455);
nor U10008 (N_10008,N_9125,N_9253);
nor U10009 (N_10009,N_9022,N_9532);
or U10010 (N_10010,N_9719,N_9465);
nor U10011 (N_10011,N_9781,N_9264);
and U10012 (N_10012,N_9324,N_9634);
xnor U10013 (N_10013,N_9297,N_9257);
and U10014 (N_10014,N_9333,N_9796);
and U10015 (N_10015,N_9903,N_9062);
and U10016 (N_10016,N_9748,N_9700);
or U10017 (N_10017,N_9543,N_9564);
and U10018 (N_10018,N_9577,N_9588);
and U10019 (N_10019,N_9172,N_9271);
nor U10020 (N_10020,N_9169,N_9614);
and U10021 (N_10021,N_9316,N_9514);
nand U10022 (N_10022,N_9811,N_9278);
nand U10023 (N_10023,N_9896,N_9262);
and U10024 (N_10024,N_9727,N_9444);
or U10025 (N_10025,N_9506,N_9296);
nor U10026 (N_10026,N_9010,N_9193);
and U10027 (N_10027,N_9866,N_9124);
xnor U10028 (N_10028,N_9395,N_9752);
nor U10029 (N_10029,N_9376,N_9621);
nand U10030 (N_10030,N_9663,N_9282);
and U10031 (N_10031,N_9292,N_9391);
xor U10032 (N_10032,N_9049,N_9187);
xor U10033 (N_10033,N_9398,N_9552);
and U10034 (N_10034,N_9168,N_9142);
nor U10035 (N_10035,N_9009,N_9823);
nor U10036 (N_10036,N_9947,N_9005);
and U10037 (N_10037,N_9043,N_9094);
nor U10038 (N_10038,N_9403,N_9387);
nand U10039 (N_10039,N_9042,N_9404);
nor U10040 (N_10040,N_9438,N_9161);
xnor U10041 (N_10041,N_9131,N_9858);
nor U10042 (N_10042,N_9978,N_9706);
nand U10043 (N_10043,N_9595,N_9639);
or U10044 (N_10044,N_9097,N_9284);
or U10045 (N_10045,N_9312,N_9907);
nand U10046 (N_10046,N_9689,N_9283);
nand U10047 (N_10047,N_9030,N_9237);
nand U10048 (N_10048,N_9270,N_9078);
nor U10049 (N_10049,N_9002,N_9520);
nand U10050 (N_10050,N_9303,N_9860);
nand U10051 (N_10051,N_9613,N_9068);
xnor U10052 (N_10052,N_9905,N_9191);
nor U10053 (N_10053,N_9383,N_9892);
or U10054 (N_10054,N_9247,N_9509);
xor U10055 (N_10055,N_9609,N_9900);
xor U10056 (N_10056,N_9790,N_9968);
and U10057 (N_10057,N_9450,N_9176);
nor U10058 (N_10058,N_9763,N_9877);
nor U10059 (N_10059,N_9849,N_9460);
nand U10060 (N_10060,N_9904,N_9315);
nand U10061 (N_10061,N_9225,N_9654);
nor U10062 (N_10062,N_9684,N_9065);
and U10063 (N_10063,N_9932,N_9650);
or U10064 (N_10064,N_9734,N_9294);
nand U10065 (N_10065,N_9083,N_9227);
nand U10066 (N_10066,N_9546,N_9000);
or U10067 (N_10067,N_9409,N_9522);
and U10068 (N_10068,N_9863,N_9682);
nand U10069 (N_10069,N_9276,N_9224);
nor U10070 (N_10070,N_9573,N_9580);
and U10071 (N_10071,N_9565,N_9024);
nand U10072 (N_10072,N_9659,N_9649);
nand U10073 (N_10073,N_9795,N_9017);
or U10074 (N_10074,N_9412,N_9587);
nor U10075 (N_10075,N_9310,N_9025);
or U10076 (N_10076,N_9973,N_9109);
or U10077 (N_10077,N_9707,N_9267);
xnor U10078 (N_10078,N_9545,N_9553);
nor U10079 (N_10079,N_9711,N_9602);
nor U10080 (N_10080,N_9640,N_9846);
nand U10081 (N_10081,N_9513,N_9632);
and U10082 (N_10082,N_9536,N_9328);
nand U10083 (N_10083,N_9056,N_9058);
xnor U10084 (N_10084,N_9319,N_9320);
xnor U10085 (N_10085,N_9933,N_9851);
or U10086 (N_10086,N_9867,N_9365);
and U10087 (N_10087,N_9622,N_9472);
nand U10088 (N_10088,N_9060,N_9133);
nand U10089 (N_10089,N_9447,N_9433);
xor U10090 (N_10090,N_9642,N_9802);
and U10091 (N_10091,N_9666,N_9072);
nand U10092 (N_10092,N_9054,N_9742);
nor U10093 (N_10093,N_9493,N_9576);
xor U10094 (N_10094,N_9794,N_9202);
xor U10095 (N_10095,N_9070,N_9150);
and U10096 (N_10096,N_9199,N_9188);
xor U10097 (N_10097,N_9361,N_9336);
nor U10098 (N_10098,N_9345,N_9901);
nand U10099 (N_10099,N_9680,N_9250);
nand U10100 (N_10100,N_9557,N_9853);
or U10101 (N_10101,N_9414,N_9881);
and U10102 (N_10102,N_9130,N_9601);
nand U10103 (N_10103,N_9606,N_9562);
or U10104 (N_10104,N_9985,N_9212);
xnor U10105 (N_10105,N_9817,N_9530);
nand U10106 (N_10106,N_9313,N_9647);
or U10107 (N_10107,N_9952,N_9218);
and U10108 (N_10108,N_9041,N_9677);
and U10109 (N_10109,N_9652,N_9238);
xor U10110 (N_10110,N_9789,N_9996);
and U10111 (N_10111,N_9750,N_9340);
or U10112 (N_10112,N_9827,N_9626);
xor U10113 (N_10113,N_9101,N_9048);
nor U10114 (N_10114,N_9113,N_9887);
or U10115 (N_10115,N_9873,N_9665);
xnor U10116 (N_10116,N_9174,N_9852);
nand U10117 (N_10117,N_9772,N_9126);
xor U10118 (N_10118,N_9798,N_9965);
and U10119 (N_10119,N_9026,N_9209);
xnor U10120 (N_10120,N_9696,N_9175);
xnor U10121 (N_10121,N_9200,N_9137);
nand U10122 (N_10122,N_9631,N_9233);
xnor U10123 (N_10123,N_9329,N_9138);
xnor U10124 (N_10124,N_9816,N_9627);
xnor U10125 (N_10125,N_9053,N_9793);
or U10126 (N_10126,N_9069,N_9239);
nor U10127 (N_10127,N_9366,N_9071);
nand U10128 (N_10128,N_9641,N_9628);
nand U10129 (N_10129,N_9957,N_9693);
or U10130 (N_10130,N_9585,N_9882);
nand U10131 (N_10131,N_9857,N_9568);
or U10132 (N_10132,N_9122,N_9166);
and U10133 (N_10133,N_9676,N_9660);
and U10134 (N_10134,N_9898,N_9268);
xor U10135 (N_10135,N_9945,N_9716);
and U10136 (N_10136,N_9314,N_9301);
nand U10137 (N_10137,N_9219,N_9098);
and U10138 (N_10138,N_9426,N_9938);
nor U10139 (N_10139,N_9321,N_9624);
or U10140 (N_10140,N_9061,N_9103);
nand U10141 (N_10141,N_9141,N_9087);
and U10142 (N_10142,N_9761,N_9721);
or U10143 (N_10143,N_9291,N_9067);
or U10144 (N_10144,N_9159,N_9765);
nor U10145 (N_10145,N_9555,N_9106);
or U10146 (N_10146,N_9948,N_9077);
and U10147 (N_10147,N_9116,N_9423);
and U10148 (N_10148,N_9425,N_9604);
nor U10149 (N_10149,N_9389,N_9779);
xor U10150 (N_10150,N_9306,N_9453);
xor U10151 (N_10151,N_9507,N_9217);
and U10152 (N_10152,N_9038,N_9512);
and U10153 (N_10153,N_9277,N_9379);
xor U10154 (N_10154,N_9348,N_9739);
nor U10155 (N_10155,N_9201,N_9894);
xor U10156 (N_10156,N_9986,N_9347);
nand U10157 (N_10157,N_9807,N_9363);
nand U10158 (N_10158,N_9095,N_9865);
or U10159 (N_10159,N_9050,N_9223);
nor U10160 (N_10160,N_9713,N_9788);
nor U10161 (N_10161,N_9970,N_9534);
nor U10162 (N_10162,N_9105,N_9740);
nor U10163 (N_10163,N_9988,N_9619);
nand U10164 (N_10164,N_9027,N_9623);
nor U10165 (N_10165,N_9667,N_9484);
nand U10166 (N_10166,N_9670,N_9474);
nor U10167 (N_10167,N_9246,N_9864);
xor U10168 (N_10168,N_9886,N_9850);
nand U10169 (N_10169,N_9066,N_9777);
or U10170 (N_10170,N_9556,N_9353);
nand U10171 (N_10171,N_9868,N_9951);
or U10172 (N_10172,N_9279,N_9298);
xor U10173 (N_10173,N_9597,N_9251);
nor U10174 (N_10174,N_9773,N_9355);
nand U10175 (N_10175,N_9288,N_9746);
and U10176 (N_10176,N_9419,N_9697);
xor U10177 (N_10177,N_9936,N_9003);
nand U10178 (N_10178,N_9729,N_9813);
xor U10179 (N_10179,N_9551,N_9749);
nor U10180 (N_10180,N_9369,N_9299);
xor U10181 (N_10181,N_9921,N_9452);
nor U10182 (N_10182,N_9954,N_9229);
nor U10183 (N_10183,N_9525,N_9107);
xnor U10184 (N_10184,N_9844,N_9089);
or U10185 (N_10185,N_9144,N_9004);
nand U10186 (N_10186,N_9511,N_9737);
or U10187 (N_10187,N_9554,N_9346);
or U10188 (N_10188,N_9959,N_9088);
nand U10189 (N_10189,N_9280,N_9531);
nor U10190 (N_10190,N_9692,N_9982);
nand U10191 (N_10191,N_9173,N_9931);
or U10192 (N_10192,N_9386,N_9494);
nor U10193 (N_10193,N_9032,N_9093);
or U10194 (N_10194,N_9302,N_9350);
or U10195 (N_10195,N_9994,N_9800);
nor U10196 (N_10196,N_9194,N_9774);
nor U10197 (N_10197,N_9498,N_9709);
nor U10198 (N_10198,N_9051,N_9728);
xor U10199 (N_10199,N_9987,N_9610);
xnor U10200 (N_10200,N_9307,N_9690);
or U10201 (N_10201,N_9919,N_9388);
and U10202 (N_10202,N_9012,N_9318);
and U10203 (N_10203,N_9528,N_9084);
nand U10204 (N_10204,N_9243,N_9521);
nand U10205 (N_10205,N_9226,N_9178);
and U10206 (N_10206,N_9019,N_9152);
and U10207 (N_10207,N_9992,N_9074);
nand U10208 (N_10208,N_9177,N_9869);
xnor U10209 (N_10209,N_9879,N_9338);
xor U10210 (N_10210,N_9162,N_9216);
nand U10211 (N_10211,N_9838,N_9782);
nand U10212 (N_10212,N_9293,N_9439);
and U10213 (N_10213,N_9206,N_9547);
nand U10214 (N_10214,N_9819,N_9821);
and U10215 (N_10215,N_9544,N_9134);
nand U10216 (N_10216,N_9842,N_9421);
nor U10217 (N_10217,N_9598,N_9469);
and U10218 (N_10218,N_9617,N_9516);
nor U10219 (N_10219,N_9435,N_9636);
and U10220 (N_10220,N_9625,N_9490);
nand U10221 (N_10221,N_9741,N_9228);
or U10222 (N_10222,N_9232,N_9723);
or U10223 (N_10223,N_9029,N_9462);
xnor U10224 (N_10224,N_9091,N_9648);
and U10225 (N_10225,N_9230,N_9908);
nor U10226 (N_10226,N_9550,N_9977);
nand U10227 (N_10227,N_9756,N_9934);
or U10228 (N_10228,N_9123,N_9526);
nor U10229 (N_10229,N_9840,N_9016);
xnor U10230 (N_10230,N_9717,N_9578);
or U10231 (N_10231,N_9859,N_9111);
and U10232 (N_10232,N_9377,N_9099);
xor U10233 (N_10233,N_9018,N_9778);
nor U10234 (N_10234,N_9561,N_9160);
nand U10235 (N_10235,N_9235,N_9359);
or U10236 (N_10236,N_9997,N_9681);
nor U10237 (N_10237,N_9411,N_9664);
nand U10238 (N_10238,N_9382,N_9920);
nand U10239 (N_10239,N_9487,N_9834);
nor U10240 (N_10240,N_9086,N_9630);
xnor U10241 (N_10241,N_9593,N_9192);
nor U10242 (N_10242,N_9913,N_9402);
nor U10243 (N_10243,N_9658,N_9431);
and U10244 (N_10244,N_9922,N_9683);
and U10245 (N_10245,N_9703,N_9325);
xnor U10246 (N_10246,N_9535,N_9211);
nor U10247 (N_10247,N_9822,N_9405);
or U10248 (N_10248,N_9135,N_9236);
nor U10249 (N_10249,N_9644,N_9466);
and U10250 (N_10250,N_9184,N_9889);
nor U10251 (N_10251,N_9575,N_9941);
or U10252 (N_10252,N_9810,N_9833);
or U10253 (N_10253,N_9245,N_9620);
and U10254 (N_10254,N_9416,N_9021);
and U10255 (N_10255,N_9286,N_9394);
or U10256 (N_10256,N_9738,N_9946);
or U10257 (N_10257,N_9744,N_9549);
or U10258 (N_10258,N_9927,N_9510);
nand U10259 (N_10259,N_9372,N_9991);
nor U10260 (N_10260,N_9566,N_9427);
nand U10261 (N_10261,N_9758,N_9736);
nor U10262 (N_10262,N_9743,N_9539);
or U10263 (N_10263,N_9502,N_9888);
and U10264 (N_10264,N_9437,N_9776);
nor U10265 (N_10265,N_9352,N_9914);
or U10266 (N_10266,N_9430,N_9208);
nor U10267 (N_10267,N_9167,N_9845);
and U10268 (N_10268,N_9616,N_9847);
nor U10269 (N_10269,N_9001,N_9269);
xor U10270 (N_10270,N_9059,N_9317);
or U10271 (N_10271,N_9085,N_9836);
nor U10272 (N_10272,N_9967,N_9373);
nand U10273 (N_10273,N_9818,N_9963);
nand U10274 (N_10274,N_9221,N_9031);
xor U10275 (N_10275,N_9909,N_9586);
and U10276 (N_10276,N_9615,N_9289);
and U10277 (N_10277,N_9413,N_9481);
nand U10278 (N_10278,N_9529,N_9770);
and U10279 (N_10279,N_9454,N_9491);
and U10280 (N_10280,N_9210,N_9792);
xor U10281 (N_10281,N_9203,N_9344);
and U10282 (N_10282,N_9691,N_9784);
nand U10283 (N_10283,N_9397,N_9256);
nand U10284 (N_10284,N_9582,N_9542);
or U10285 (N_10285,N_9139,N_9249);
nand U10286 (N_10286,N_9831,N_9429);
or U10287 (N_10287,N_9891,N_9854);
nor U10288 (N_10288,N_9244,N_9768);
and U10289 (N_10289,N_9020,N_9600);
nand U10290 (N_10290,N_9733,N_9114);
or U10291 (N_10291,N_9645,N_9517);
xor U10292 (N_10292,N_9183,N_9182);
and U10293 (N_10293,N_9198,N_9505);
xor U10294 (N_10294,N_9343,N_9753);
xor U10295 (N_10295,N_9754,N_9220);
or U10296 (N_10296,N_9540,N_9956);
xnor U10297 (N_10297,N_9976,N_9163);
or U10298 (N_10298,N_9214,N_9839);
and U10299 (N_10299,N_9856,N_9266);
nand U10300 (N_10300,N_9441,N_9400);
xor U10301 (N_10301,N_9806,N_9783);
nor U10302 (N_10302,N_9767,N_9272);
nand U10303 (N_10303,N_9331,N_9942);
or U10304 (N_10304,N_9351,N_9953);
and U10305 (N_10305,N_9456,N_9273);
nand U10306 (N_10306,N_9108,N_9895);
or U10307 (N_10307,N_9492,N_9570);
nor U10308 (N_10308,N_9558,N_9368);
nand U10309 (N_10309,N_9591,N_9969);
or U10310 (N_10310,N_9911,N_9357);
xnor U10311 (N_10311,N_9102,N_9702);
xnor U10312 (N_10312,N_9463,N_9747);
and U10313 (N_10313,N_9799,N_9028);
nor U10314 (N_10314,N_9483,N_9899);
or U10315 (N_10315,N_9263,N_9979);
nor U10316 (N_10316,N_9829,N_9828);
nor U10317 (N_10317,N_9950,N_9949);
or U10318 (N_10318,N_9944,N_9805);
nor U10319 (N_10319,N_9791,N_9637);
nor U10320 (N_10320,N_9657,N_9519);
nor U10321 (N_10321,N_9843,N_9801);
xor U10322 (N_10322,N_9440,N_9073);
and U10323 (N_10323,N_9508,N_9714);
nor U10324 (N_10324,N_9999,N_9457);
nand U10325 (N_10325,N_9234,N_9672);
and U10326 (N_10326,N_9915,N_9390);
nor U10327 (N_10327,N_9170,N_9308);
or U10328 (N_10328,N_9158,N_9764);
or U10329 (N_10329,N_9448,N_9704);
and U10330 (N_10330,N_9605,N_9478);
or U10331 (N_10331,N_9824,N_9735);
nand U10332 (N_10332,N_9486,N_9092);
xnor U10333 (N_10333,N_9629,N_9745);
xor U10334 (N_10334,N_9396,N_9104);
xor U10335 (N_10335,N_9153,N_9036);
nand U10336 (N_10336,N_9603,N_9354);
nand U10337 (N_10337,N_9830,N_9146);
xor U10338 (N_10338,N_9964,N_9724);
nand U10339 (N_10339,N_9730,N_9285);
nand U10340 (N_10340,N_9436,N_9884);
nor U10341 (N_10341,N_9718,N_9918);
nor U10342 (N_10342,N_9890,N_9916);
xnor U10343 (N_10343,N_9592,N_9548);
nand U10344 (N_10344,N_9295,N_9937);
xnor U10345 (N_10345,N_9148,N_9538);
xor U10346 (N_10346,N_9132,N_9215);
nand U10347 (N_10347,N_9668,N_9712);
nand U10348 (N_10348,N_9014,N_9254);
nand U10349 (N_10349,N_9207,N_9883);
nor U10350 (N_10350,N_9780,N_9559);
or U10351 (N_10351,N_9785,N_9826);
and U10352 (N_10352,N_9503,N_9928);
xnor U10353 (N_10353,N_9815,N_9446);
xor U10354 (N_10354,N_9480,N_9181);
and U10355 (N_10355,N_9797,N_9241);
xnor U10356 (N_10356,N_9477,N_9461);
or U10357 (N_10357,N_9820,N_9926);
and U10358 (N_10358,N_9541,N_9485);
xor U10359 (N_10359,N_9100,N_9878);
nor U10360 (N_10360,N_9533,N_9924);
xnor U10361 (N_10361,N_9341,N_9897);
nor U10362 (N_10362,N_9034,N_9339);
or U10363 (N_10363,N_9330,N_9458);
or U10364 (N_10364,N_9118,N_9143);
or U10365 (N_10365,N_9990,N_9653);
xor U10366 (N_10366,N_9076,N_9504);
or U10367 (N_10367,N_9082,N_9121);
xor U10368 (N_10368,N_9305,N_9468);
or U10369 (N_10369,N_9055,N_9874);
nor U10370 (N_10370,N_9304,N_9470);
xnor U10371 (N_10371,N_9309,N_9196);
or U10372 (N_10372,N_9581,N_9044);
nand U10373 (N_10373,N_9923,N_9925);
xnor U10374 (N_10374,N_9686,N_9120);
xnor U10375 (N_10375,N_9832,N_9993);
nand U10376 (N_10376,N_9471,N_9079);
nand U10377 (N_10377,N_9418,N_9190);
nor U10378 (N_10378,N_9489,N_9646);
nand U10379 (N_10379,N_9281,N_9335);
xor U10380 (N_10380,N_9961,N_9231);
or U10381 (N_10381,N_9612,N_9981);
or U10382 (N_10382,N_9407,N_9110);
xor U10383 (N_10383,N_9803,N_9876);
or U10384 (N_10384,N_9180,N_9769);
or U10385 (N_10385,N_9064,N_9370);
nand U10386 (N_10386,N_9323,N_9378);
nand U10387 (N_10387,N_9259,N_9290);
xor U10388 (N_10388,N_9523,N_9119);
nor U10389 (N_10389,N_9424,N_9204);
and U10390 (N_10390,N_9731,N_9422);
xor U10391 (N_10391,N_9935,N_9205);
nor U10392 (N_10392,N_9910,N_9687);
xnor U10393 (N_10393,N_9755,N_9147);
and U10394 (N_10394,N_9045,N_9443);
nor U10395 (N_10395,N_9837,N_9757);
or U10396 (N_10396,N_9760,N_9635);
or U10397 (N_10397,N_9701,N_9155);
nand U10398 (N_10398,N_9432,N_9574);
or U10399 (N_10399,N_9673,N_9955);
nand U10400 (N_10400,N_9611,N_9035);
and U10401 (N_10401,N_9771,N_9699);
nand U10402 (N_10402,N_9618,N_9011);
nor U10403 (N_10403,N_9579,N_9875);
or U10404 (N_10404,N_9381,N_9675);
xnor U10405 (N_10405,N_9384,N_9274);
or U10406 (N_10406,N_9589,N_9408);
and U10407 (N_10407,N_9459,N_9972);
nor U10408 (N_10408,N_9651,N_9287);
nor U10409 (N_10409,N_9410,N_9063);
or U10410 (N_10410,N_9688,N_9371);
nand U10411 (N_10411,N_9497,N_9638);
xor U10412 (N_10412,N_9848,N_9962);
or U10413 (N_10413,N_9488,N_9362);
nand U10414 (N_10414,N_9715,N_9608);
nor U10415 (N_10415,N_9171,N_9872);
nand U10416 (N_10416,N_9136,N_9537);
nand U10417 (N_10417,N_9360,N_9499);
or U10418 (N_10418,N_9033,N_9090);
or U10419 (N_10419,N_9189,N_9240);
nor U10420 (N_10420,N_9157,N_9300);
nand U10421 (N_10421,N_9417,N_9096);
or U10422 (N_10422,N_9720,N_9893);
and U10423 (N_10423,N_9392,N_9871);
or U10424 (N_10424,N_9671,N_9195);
nor U10425 (N_10425,N_9710,N_9129);
and U10426 (N_10426,N_9766,N_9841);
nand U10427 (N_10427,N_9334,N_9870);
nor U10428 (N_10428,N_9902,N_9385);
nor U10429 (N_10429,N_9258,N_9007);
nand U10430 (N_10430,N_9607,N_9475);
xor U10431 (N_10431,N_9563,N_9662);
xnor U10432 (N_10432,N_9008,N_9804);
nand U10433 (N_10433,N_9751,N_9179);
nor U10434 (N_10434,N_9560,N_9265);
xnor U10435 (N_10435,N_9349,N_9974);
nor U10436 (N_10436,N_9698,N_9327);
nand U10437 (N_10437,N_9222,N_9482);
or U10438 (N_10438,N_9584,N_9685);
and U10439 (N_10439,N_9260,N_9275);
nor U10440 (N_10440,N_9943,N_9787);
and U10441 (N_10441,N_9995,N_9140);
nor U10442 (N_10442,N_9694,N_9467);
nor U10443 (N_10443,N_9775,N_9013);
nor U10444 (N_10444,N_9399,N_9364);
and U10445 (N_10445,N_9197,N_9661);
and U10446 (N_10446,N_9023,N_9572);
nand U10447 (N_10447,N_9464,N_9583);
nand U10448 (N_10448,N_9358,N_9998);
xnor U10449 (N_10449,N_9984,N_9980);
or U10450 (N_10450,N_9880,N_9479);
or U10451 (N_10451,N_9814,N_9248);
and U10452 (N_10452,N_9151,N_9401);
or U10453 (N_10453,N_9006,N_9040);
or U10454 (N_10454,N_9906,N_9940);
xnor U10455 (N_10455,N_9311,N_9326);
and U10456 (N_10456,N_9835,N_9451);
nand U10457 (N_10457,N_9434,N_9655);
xor U10458 (N_10458,N_9255,N_9633);
and U10459 (N_10459,N_9669,N_9476);
xor U10460 (N_10460,N_9930,N_9242);
xor U10461 (N_10461,N_9812,N_9406);
xnor U10462 (N_10462,N_9449,N_9808);
xnor U10463 (N_10463,N_9599,N_9643);
nor U10464 (N_10464,N_9117,N_9571);
or U10465 (N_10465,N_9695,N_9052);
nand U10466 (N_10466,N_9374,N_9975);
xor U10467 (N_10467,N_9380,N_9958);
or U10468 (N_10468,N_9356,N_9261);
or U10469 (N_10469,N_9445,N_9075);
nor U10470 (N_10470,N_9809,N_9678);
nor U10471 (N_10471,N_9185,N_9722);
nor U10472 (N_10472,N_9037,N_9393);
or U10473 (N_10473,N_9165,N_9115);
nor U10474 (N_10474,N_9989,N_9442);
xor U10475 (N_10475,N_9500,N_9759);
xor U10476 (N_10476,N_9046,N_9939);
nor U10477 (N_10477,N_9518,N_9375);
and U10478 (N_10478,N_9679,N_9156);
or U10479 (N_10479,N_9515,N_9332);
and U10480 (N_10480,N_9960,N_9420);
xor U10481 (N_10481,N_9501,N_9154);
or U10482 (N_10482,N_9786,N_9732);
nand U10483 (N_10483,N_9337,N_9971);
nor U10484 (N_10484,N_9983,N_9428);
or U10485 (N_10485,N_9473,N_9252);
or U10486 (N_10486,N_9596,N_9047);
nor U10487 (N_10487,N_9762,N_9149);
and U10488 (N_10488,N_9015,N_9080);
or U10489 (N_10489,N_9966,N_9912);
and U10490 (N_10490,N_9862,N_9112);
or U10491 (N_10491,N_9567,N_9674);
nor U10492 (N_10492,N_9885,N_9128);
or U10493 (N_10493,N_9164,N_9342);
or U10494 (N_10494,N_9855,N_9726);
or U10495 (N_10495,N_9186,N_9917);
nand U10496 (N_10496,N_9527,N_9127);
and U10497 (N_10497,N_9590,N_9213);
and U10498 (N_10498,N_9708,N_9039);
and U10499 (N_10499,N_9594,N_9415);
or U10500 (N_10500,N_9272,N_9020);
and U10501 (N_10501,N_9697,N_9700);
and U10502 (N_10502,N_9910,N_9019);
or U10503 (N_10503,N_9531,N_9585);
and U10504 (N_10504,N_9670,N_9336);
xor U10505 (N_10505,N_9080,N_9987);
and U10506 (N_10506,N_9518,N_9737);
or U10507 (N_10507,N_9776,N_9418);
nand U10508 (N_10508,N_9458,N_9569);
nand U10509 (N_10509,N_9168,N_9159);
nand U10510 (N_10510,N_9815,N_9818);
nand U10511 (N_10511,N_9002,N_9511);
nand U10512 (N_10512,N_9801,N_9103);
nand U10513 (N_10513,N_9420,N_9228);
nor U10514 (N_10514,N_9654,N_9738);
and U10515 (N_10515,N_9863,N_9771);
and U10516 (N_10516,N_9630,N_9473);
or U10517 (N_10517,N_9414,N_9257);
xnor U10518 (N_10518,N_9971,N_9291);
and U10519 (N_10519,N_9542,N_9554);
xor U10520 (N_10520,N_9102,N_9620);
and U10521 (N_10521,N_9151,N_9495);
nor U10522 (N_10522,N_9857,N_9870);
nand U10523 (N_10523,N_9797,N_9551);
and U10524 (N_10524,N_9461,N_9178);
nor U10525 (N_10525,N_9738,N_9645);
and U10526 (N_10526,N_9257,N_9003);
nand U10527 (N_10527,N_9651,N_9161);
or U10528 (N_10528,N_9774,N_9173);
xor U10529 (N_10529,N_9333,N_9538);
nor U10530 (N_10530,N_9024,N_9893);
or U10531 (N_10531,N_9506,N_9372);
and U10532 (N_10532,N_9043,N_9975);
and U10533 (N_10533,N_9013,N_9909);
or U10534 (N_10534,N_9105,N_9575);
xor U10535 (N_10535,N_9414,N_9697);
and U10536 (N_10536,N_9866,N_9780);
xnor U10537 (N_10537,N_9050,N_9668);
nand U10538 (N_10538,N_9745,N_9228);
nand U10539 (N_10539,N_9679,N_9260);
or U10540 (N_10540,N_9226,N_9089);
and U10541 (N_10541,N_9513,N_9292);
nand U10542 (N_10542,N_9070,N_9679);
or U10543 (N_10543,N_9124,N_9259);
and U10544 (N_10544,N_9226,N_9416);
nand U10545 (N_10545,N_9495,N_9555);
and U10546 (N_10546,N_9829,N_9536);
or U10547 (N_10547,N_9899,N_9028);
xnor U10548 (N_10548,N_9419,N_9932);
xor U10549 (N_10549,N_9917,N_9737);
and U10550 (N_10550,N_9871,N_9535);
xor U10551 (N_10551,N_9538,N_9784);
nand U10552 (N_10552,N_9814,N_9947);
and U10553 (N_10553,N_9180,N_9577);
nand U10554 (N_10554,N_9974,N_9929);
or U10555 (N_10555,N_9375,N_9503);
or U10556 (N_10556,N_9701,N_9970);
nor U10557 (N_10557,N_9921,N_9666);
nor U10558 (N_10558,N_9795,N_9324);
and U10559 (N_10559,N_9240,N_9396);
and U10560 (N_10560,N_9713,N_9869);
nor U10561 (N_10561,N_9856,N_9200);
and U10562 (N_10562,N_9589,N_9869);
and U10563 (N_10563,N_9556,N_9178);
or U10564 (N_10564,N_9654,N_9082);
nand U10565 (N_10565,N_9795,N_9719);
nand U10566 (N_10566,N_9341,N_9526);
nor U10567 (N_10567,N_9442,N_9287);
nand U10568 (N_10568,N_9333,N_9428);
and U10569 (N_10569,N_9573,N_9834);
xnor U10570 (N_10570,N_9815,N_9509);
xor U10571 (N_10571,N_9080,N_9543);
or U10572 (N_10572,N_9821,N_9994);
and U10573 (N_10573,N_9300,N_9224);
xor U10574 (N_10574,N_9807,N_9190);
nor U10575 (N_10575,N_9172,N_9104);
xnor U10576 (N_10576,N_9673,N_9850);
nand U10577 (N_10577,N_9590,N_9666);
and U10578 (N_10578,N_9251,N_9678);
xor U10579 (N_10579,N_9752,N_9089);
nor U10580 (N_10580,N_9511,N_9619);
xor U10581 (N_10581,N_9932,N_9778);
xor U10582 (N_10582,N_9816,N_9319);
nand U10583 (N_10583,N_9524,N_9019);
and U10584 (N_10584,N_9508,N_9686);
nand U10585 (N_10585,N_9907,N_9731);
nand U10586 (N_10586,N_9693,N_9154);
nand U10587 (N_10587,N_9364,N_9545);
nand U10588 (N_10588,N_9856,N_9237);
xnor U10589 (N_10589,N_9003,N_9231);
and U10590 (N_10590,N_9776,N_9128);
or U10591 (N_10591,N_9044,N_9052);
nand U10592 (N_10592,N_9971,N_9168);
or U10593 (N_10593,N_9364,N_9082);
xor U10594 (N_10594,N_9771,N_9786);
nand U10595 (N_10595,N_9979,N_9361);
or U10596 (N_10596,N_9291,N_9805);
and U10597 (N_10597,N_9716,N_9304);
nand U10598 (N_10598,N_9209,N_9140);
and U10599 (N_10599,N_9508,N_9178);
nor U10600 (N_10600,N_9539,N_9952);
or U10601 (N_10601,N_9692,N_9832);
or U10602 (N_10602,N_9765,N_9405);
or U10603 (N_10603,N_9972,N_9046);
xor U10604 (N_10604,N_9455,N_9581);
and U10605 (N_10605,N_9564,N_9895);
nor U10606 (N_10606,N_9780,N_9411);
nor U10607 (N_10607,N_9894,N_9499);
nand U10608 (N_10608,N_9108,N_9795);
nor U10609 (N_10609,N_9312,N_9781);
xor U10610 (N_10610,N_9920,N_9809);
or U10611 (N_10611,N_9801,N_9960);
and U10612 (N_10612,N_9546,N_9317);
xor U10613 (N_10613,N_9301,N_9234);
or U10614 (N_10614,N_9638,N_9093);
and U10615 (N_10615,N_9965,N_9354);
and U10616 (N_10616,N_9858,N_9868);
nand U10617 (N_10617,N_9563,N_9130);
and U10618 (N_10618,N_9323,N_9630);
nand U10619 (N_10619,N_9693,N_9797);
and U10620 (N_10620,N_9010,N_9572);
or U10621 (N_10621,N_9892,N_9567);
or U10622 (N_10622,N_9939,N_9864);
and U10623 (N_10623,N_9107,N_9552);
xor U10624 (N_10624,N_9599,N_9866);
nand U10625 (N_10625,N_9522,N_9538);
nand U10626 (N_10626,N_9491,N_9368);
nand U10627 (N_10627,N_9476,N_9770);
xor U10628 (N_10628,N_9011,N_9268);
nor U10629 (N_10629,N_9683,N_9828);
and U10630 (N_10630,N_9723,N_9958);
nand U10631 (N_10631,N_9707,N_9895);
nor U10632 (N_10632,N_9766,N_9931);
and U10633 (N_10633,N_9051,N_9099);
nor U10634 (N_10634,N_9414,N_9434);
and U10635 (N_10635,N_9918,N_9030);
or U10636 (N_10636,N_9862,N_9087);
xor U10637 (N_10637,N_9791,N_9778);
and U10638 (N_10638,N_9042,N_9031);
and U10639 (N_10639,N_9346,N_9399);
nand U10640 (N_10640,N_9402,N_9384);
or U10641 (N_10641,N_9964,N_9281);
or U10642 (N_10642,N_9411,N_9596);
and U10643 (N_10643,N_9188,N_9444);
nand U10644 (N_10644,N_9059,N_9795);
and U10645 (N_10645,N_9033,N_9808);
or U10646 (N_10646,N_9656,N_9915);
xor U10647 (N_10647,N_9694,N_9487);
nand U10648 (N_10648,N_9244,N_9756);
xor U10649 (N_10649,N_9196,N_9036);
nor U10650 (N_10650,N_9518,N_9344);
and U10651 (N_10651,N_9481,N_9800);
and U10652 (N_10652,N_9324,N_9330);
xnor U10653 (N_10653,N_9662,N_9781);
nand U10654 (N_10654,N_9952,N_9366);
and U10655 (N_10655,N_9593,N_9352);
or U10656 (N_10656,N_9272,N_9371);
xnor U10657 (N_10657,N_9102,N_9591);
xor U10658 (N_10658,N_9422,N_9746);
xor U10659 (N_10659,N_9866,N_9263);
nand U10660 (N_10660,N_9000,N_9957);
or U10661 (N_10661,N_9930,N_9443);
xor U10662 (N_10662,N_9666,N_9385);
xor U10663 (N_10663,N_9776,N_9471);
nor U10664 (N_10664,N_9516,N_9801);
or U10665 (N_10665,N_9024,N_9367);
and U10666 (N_10666,N_9644,N_9719);
xor U10667 (N_10667,N_9189,N_9746);
xnor U10668 (N_10668,N_9687,N_9760);
and U10669 (N_10669,N_9325,N_9273);
and U10670 (N_10670,N_9079,N_9736);
xnor U10671 (N_10671,N_9355,N_9849);
and U10672 (N_10672,N_9767,N_9007);
nor U10673 (N_10673,N_9551,N_9245);
xnor U10674 (N_10674,N_9717,N_9678);
and U10675 (N_10675,N_9911,N_9276);
nor U10676 (N_10676,N_9443,N_9537);
nand U10677 (N_10677,N_9229,N_9010);
or U10678 (N_10678,N_9399,N_9103);
nor U10679 (N_10679,N_9414,N_9274);
xnor U10680 (N_10680,N_9190,N_9351);
and U10681 (N_10681,N_9211,N_9732);
and U10682 (N_10682,N_9618,N_9835);
and U10683 (N_10683,N_9284,N_9165);
and U10684 (N_10684,N_9911,N_9800);
xnor U10685 (N_10685,N_9914,N_9833);
or U10686 (N_10686,N_9877,N_9428);
or U10687 (N_10687,N_9987,N_9224);
nand U10688 (N_10688,N_9801,N_9675);
nor U10689 (N_10689,N_9496,N_9559);
xor U10690 (N_10690,N_9539,N_9290);
or U10691 (N_10691,N_9259,N_9808);
xnor U10692 (N_10692,N_9379,N_9753);
nand U10693 (N_10693,N_9872,N_9591);
xor U10694 (N_10694,N_9965,N_9836);
xnor U10695 (N_10695,N_9774,N_9380);
nand U10696 (N_10696,N_9990,N_9316);
xor U10697 (N_10697,N_9183,N_9629);
or U10698 (N_10698,N_9449,N_9980);
nand U10699 (N_10699,N_9730,N_9452);
xnor U10700 (N_10700,N_9013,N_9055);
xnor U10701 (N_10701,N_9002,N_9287);
nand U10702 (N_10702,N_9944,N_9453);
or U10703 (N_10703,N_9539,N_9473);
nand U10704 (N_10704,N_9400,N_9857);
xnor U10705 (N_10705,N_9479,N_9593);
nand U10706 (N_10706,N_9197,N_9826);
xnor U10707 (N_10707,N_9236,N_9957);
and U10708 (N_10708,N_9904,N_9960);
or U10709 (N_10709,N_9395,N_9638);
or U10710 (N_10710,N_9907,N_9158);
nand U10711 (N_10711,N_9342,N_9326);
and U10712 (N_10712,N_9410,N_9821);
and U10713 (N_10713,N_9416,N_9365);
or U10714 (N_10714,N_9647,N_9873);
and U10715 (N_10715,N_9482,N_9172);
nand U10716 (N_10716,N_9715,N_9473);
nor U10717 (N_10717,N_9829,N_9575);
xor U10718 (N_10718,N_9026,N_9742);
nand U10719 (N_10719,N_9225,N_9702);
or U10720 (N_10720,N_9368,N_9970);
and U10721 (N_10721,N_9390,N_9576);
or U10722 (N_10722,N_9134,N_9874);
and U10723 (N_10723,N_9957,N_9160);
nand U10724 (N_10724,N_9259,N_9791);
xnor U10725 (N_10725,N_9231,N_9871);
nand U10726 (N_10726,N_9297,N_9167);
or U10727 (N_10727,N_9634,N_9212);
nor U10728 (N_10728,N_9333,N_9465);
and U10729 (N_10729,N_9659,N_9179);
nor U10730 (N_10730,N_9566,N_9368);
and U10731 (N_10731,N_9854,N_9117);
xnor U10732 (N_10732,N_9714,N_9385);
xor U10733 (N_10733,N_9828,N_9570);
and U10734 (N_10734,N_9527,N_9959);
xnor U10735 (N_10735,N_9623,N_9856);
nand U10736 (N_10736,N_9087,N_9054);
or U10737 (N_10737,N_9745,N_9576);
nor U10738 (N_10738,N_9705,N_9416);
xor U10739 (N_10739,N_9840,N_9751);
and U10740 (N_10740,N_9530,N_9288);
xor U10741 (N_10741,N_9884,N_9998);
and U10742 (N_10742,N_9149,N_9480);
xor U10743 (N_10743,N_9466,N_9996);
or U10744 (N_10744,N_9633,N_9295);
or U10745 (N_10745,N_9309,N_9197);
nand U10746 (N_10746,N_9709,N_9993);
and U10747 (N_10747,N_9341,N_9519);
nand U10748 (N_10748,N_9829,N_9095);
nor U10749 (N_10749,N_9855,N_9935);
nand U10750 (N_10750,N_9859,N_9267);
nor U10751 (N_10751,N_9865,N_9448);
nor U10752 (N_10752,N_9751,N_9127);
and U10753 (N_10753,N_9613,N_9465);
nand U10754 (N_10754,N_9391,N_9093);
nor U10755 (N_10755,N_9238,N_9185);
or U10756 (N_10756,N_9390,N_9497);
and U10757 (N_10757,N_9634,N_9935);
nand U10758 (N_10758,N_9552,N_9201);
xnor U10759 (N_10759,N_9494,N_9916);
xnor U10760 (N_10760,N_9857,N_9644);
and U10761 (N_10761,N_9329,N_9444);
or U10762 (N_10762,N_9545,N_9259);
nand U10763 (N_10763,N_9538,N_9716);
nor U10764 (N_10764,N_9521,N_9036);
or U10765 (N_10765,N_9534,N_9736);
nor U10766 (N_10766,N_9978,N_9123);
nand U10767 (N_10767,N_9350,N_9234);
and U10768 (N_10768,N_9590,N_9512);
nand U10769 (N_10769,N_9172,N_9825);
xor U10770 (N_10770,N_9442,N_9099);
nor U10771 (N_10771,N_9478,N_9576);
nand U10772 (N_10772,N_9513,N_9055);
nor U10773 (N_10773,N_9510,N_9537);
and U10774 (N_10774,N_9992,N_9897);
nor U10775 (N_10775,N_9919,N_9763);
xnor U10776 (N_10776,N_9014,N_9453);
or U10777 (N_10777,N_9527,N_9376);
nor U10778 (N_10778,N_9252,N_9189);
nand U10779 (N_10779,N_9321,N_9060);
nor U10780 (N_10780,N_9268,N_9764);
xnor U10781 (N_10781,N_9863,N_9033);
nand U10782 (N_10782,N_9291,N_9501);
nand U10783 (N_10783,N_9963,N_9994);
and U10784 (N_10784,N_9536,N_9225);
and U10785 (N_10785,N_9213,N_9412);
nor U10786 (N_10786,N_9291,N_9253);
or U10787 (N_10787,N_9996,N_9397);
and U10788 (N_10788,N_9475,N_9925);
or U10789 (N_10789,N_9624,N_9094);
nand U10790 (N_10790,N_9111,N_9696);
nand U10791 (N_10791,N_9423,N_9907);
or U10792 (N_10792,N_9746,N_9556);
xnor U10793 (N_10793,N_9819,N_9205);
and U10794 (N_10794,N_9159,N_9583);
nor U10795 (N_10795,N_9201,N_9788);
nor U10796 (N_10796,N_9166,N_9913);
or U10797 (N_10797,N_9268,N_9466);
and U10798 (N_10798,N_9066,N_9724);
and U10799 (N_10799,N_9227,N_9511);
nand U10800 (N_10800,N_9450,N_9670);
xnor U10801 (N_10801,N_9102,N_9172);
nand U10802 (N_10802,N_9147,N_9974);
xor U10803 (N_10803,N_9742,N_9010);
xor U10804 (N_10804,N_9401,N_9422);
nand U10805 (N_10805,N_9672,N_9333);
xor U10806 (N_10806,N_9594,N_9399);
and U10807 (N_10807,N_9371,N_9355);
nor U10808 (N_10808,N_9647,N_9525);
or U10809 (N_10809,N_9437,N_9902);
nand U10810 (N_10810,N_9780,N_9260);
nand U10811 (N_10811,N_9116,N_9353);
and U10812 (N_10812,N_9083,N_9185);
xnor U10813 (N_10813,N_9060,N_9140);
xnor U10814 (N_10814,N_9050,N_9832);
nand U10815 (N_10815,N_9222,N_9776);
and U10816 (N_10816,N_9007,N_9243);
nand U10817 (N_10817,N_9279,N_9373);
nand U10818 (N_10818,N_9658,N_9983);
or U10819 (N_10819,N_9651,N_9506);
and U10820 (N_10820,N_9787,N_9979);
and U10821 (N_10821,N_9363,N_9915);
nand U10822 (N_10822,N_9819,N_9775);
or U10823 (N_10823,N_9568,N_9695);
xnor U10824 (N_10824,N_9366,N_9248);
or U10825 (N_10825,N_9715,N_9541);
xor U10826 (N_10826,N_9756,N_9066);
and U10827 (N_10827,N_9875,N_9634);
nand U10828 (N_10828,N_9630,N_9123);
nand U10829 (N_10829,N_9040,N_9450);
or U10830 (N_10830,N_9667,N_9163);
nor U10831 (N_10831,N_9520,N_9813);
or U10832 (N_10832,N_9312,N_9631);
nor U10833 (N_10833,N_9964,N_9215);
xnor U10834 (N_10834,N_9189,N_9875);
or U10835 (N_10835,N_9965,N_9135);
nand U10836 (N_10836,N_9695,N_9703);
and U10837 (N_10837,N_9184,N_9027);
nor U10838 (N_10838,N_9542,N_9563);
nor U10839 (N_10839,N_9455,N_9826);
xor U10840 (N_10840,N_9351,N_9875);
and U10841 (N_10841,N_9551,N_9342);
or U10842 (N_10842,N_9327,N_9788);
nand U10843 (N_10843,N_9979,N_9341);
or U10844 (N_10844,N_9101,N_9807);
or U10845 (N_10845,N_9983,N_9169);
and U10846 (N_10846,N_9816,N_9230);
or U10847 (N_10847,N_9549,N_9352);
nor U10848 (N_10848,N_9583,N_9407);
nor U10849 (N_10849,N_9937,N_9577);
or U10850 (N_10850,N_9020,N_9081);
and U10851 (N_10851,N_9167,N_9116);
and U10852 (N_10852,N_9988,N_9042);
nor U10853 (N_10853,N_9532,N_9124);
nor U10854 (N_10854,N_9849,N_9871);
nor U10855 (N_10855,N_9579,N_9521);
or U10856 (N_10856,N_9690,N_9253);
and U10857 (N_10857,N_9626,N_9563);
xnor U10858 (N_10858,N_9422,N_9266);
or U10859 (N_10859,N_9769,N_9406);
or U10860 (N_10860,N_9323,N_9099);
xnor U10861 (N_10861,N_9920,N_9452);
or U10862 (N_10862,N_9064,N_9580);
xnor U10863 (N_10863,N_9672,N_9925);
nand U10864 (N_10864,N_9702,N_9846);
or U10865 (N_10865,N_9883,N_9018);
xor U10866 (N_10866,N_9883,N_9497);
or U10867 (N_10867,N_9903,N_9575);
and U10868 (N_10868,N_9358,N_9970);
xnor U10869 (N_10869,N_9892,N_9090);
nand U10870 (N_10870,N_9025,N_9950);
nand U10871 (N_10871,N_9394,N_9517);
nor U10872 (N_10872,N_9872,N_9979);
and U10873 (N_10873,N_9198,N_9519);
and U10874 (N_10874,N_9451,N_9228);
and U10875 (N_10875,N_9750,N_9890);
nand U10876 (N_10876,N_9109,N_9413);
nor U10877 (N_10877,N_9193,N_9544);
nor U10878 (N_10878,N_9900,N_9736);
xor U10879 (N_10879,N_9823,N_9689);
or U10880 (N_10880,N_9678,N_9011);
and U10881 (N_10881,N_9829,N_9823);
nand U10882 (N_10882,N_9844,N_9828);
nand U10883 (N_10883,N_9885,N_9567);
nor U10884 (N_10884,N_9759,N_9823);
nand U10885 (N_10885,N_9215,N_9078);
or U10886 (N_10886,N_9906,N_9173);
or U10887 (N_10887,N_9122,N_9369);
xor U10888 (N_10888,N_9980,N_9577);
xor U10889 (N_10889,N_9122,N_9159);
nor U10890 (N_10890,N_9760,N_9856);
and U10891 (N_10891,N_9898,N_9610);
nor U10892 (N_10892,N_9947,N_9599);
and U10893 (N_10893,N_9824,N_9543);
nor U10894 (N_10894,N_9824,N_9610);
or U10895 (N_10895,N_9009,N_9771);
nand U10896 (N_10896,N_9165,N_9695);
and U10897 (N_10897,N_9295,N_9761);
nand U10898 (N_10898,N_9294,N_9736);
nand U10899 (N_10899,N_9100,N_9992);
nor U10900 (N_10900,N_9860,N_9589);
or U10901 (N_10901,N_9715,N_9612);
xor U10902 (N_10902,N_9295,N_9729);
and U10903 (N_10903,N_9111,N_9481);
and U10904 (N_10904,N_9812,N_9485);
and U10905 (N_10905,N_9580,N_9806);
or U10906 (N_10906,N_9995,N_9590);
xor U10907 (N_10907,N_9771,N_9125);
xnor U10908 (N_10908,N_9149,N_9651);
nor U10909 (N_10909,N_9123,N_9389);
xnor U10910 (N_10910,N_9592,N_9578);
and U10911 (N_10911,N_9047,N_9543);
or U10912 (N_10912,N_9013,N_9290);
and U10913 (N_10913,N_9615,N_9778);
nand U10914 (N_10914,N_9371,N_9274);
or U10915 (N_10915,N_9296,N_9688);
xor U10916 (N_10916,N_9627,N_9760);
nand U10917 (N_10917,N_9378,N_9878);
or U10918 (N_10918,N_9901,N_9512);
xnor U10919 (N_10919,N_9569,N_9412);
and U10920 (N_10920,N_9078,N_9665);
nand U10921 (N_10921,N_9365,N_9410);
nor U10922 (N_10922,N_9461,N_9007);
or U10923 (N_10923,N_9850,N_9126);
and U10924 (N_10924,N_9005,N_9398);
nand U10925 (N_10925,N_9480,N_9803);
and U10926 (N_10926,N_9336,N_9992);
nand U10927 (N_10927,N_9869,N_9728);
nor U10928 (N_10928,N_9272,N_9910);
and U10929 (N_10929,N_9189,N_9335);
xnor U10930 (N_10930,N_9208,N_9314);
xor U10931 (N_10931,N_9308,N_9147);
nand U10932 (N_10932,N_9982,N_9301);
nor U10933 (N_10933,N_9385,N_9467);
and U10934 (N_10934,N_9124,N_9401);
nor U10935 (N_10935,N_9193,N_9443);
nor U10936 (N_10936,N_9559,N_9937);
nand U10937 (N_10937,N_9281,N_9004);
nor U10938 (N_10938,N_9973,N_9794);
nand U10939 (N_10939,N_9309,N_9252);
or U10940 (N_10940,N_9735,N_9391);
or U10941 (N_10941,N_9511,N_9500);
xnor U10942 (N_10942,N_9978,N_9406);
or U10943 (N_10943,N_9013,N_9441);
nand U10944 (N_10944,N_9293,N_9487);
nand U10945 (N_10945,N_9986,N_9176);
and U10946 (N_10946,N_9938,N_9302);
nor U10947 (N_10947,N_9862,N_9897);
and U10948 (N_10948,N_9941,N_9539);
nor U10949 (N_10949,N_9566,N_9983);
and U10950 (N_10950,N_9250,N_9538);
and U10951 (N_10951,N_9014,N_9522);
nand U10952 (N_10952,N_9331,N_9857);
nand U10953 (N_10953,N_9713,N_9418);
nor U10954 (N_10954,N_9751,N_9158);
nand U10955 (N_10955,N_9681,N_9799);
nand U10956 (N_10956,N_9121,N_9191);
or U10957 (N_10957,N_9150,N_9471);
and U10958 (N_10958,N_9454,N_9169);
nand U10959 (N_10959,N_9054,N_9576);
nor U10960 (N_10960,N_9525,N_9482);
nand U10961 (N_10961,N_9291,N_9524);
nand U10962 (N_10962,N_9107,N_9882);
nor U10963 (N_10963,N_9304,N_9733);
nand U10964 (N_10964,N_9546,N_9610);
or U10965 (N_10965,N_9668,N_9588);
or U10966 (N_10966,N_9567,N_9028);
xor U10967 (N_10967,N_9682,N_9019);
nor U10968 (N_10968,N_9372,N_9522);
nand U10969 (N_10969,N_9798,N_9581);
nor U10970 (N_10970,N_9652,N_9628);
nor U10971 (N_10971,N_9230,N_9631);
xor U10972 (N_10972,N_9340,N_9130);
xnor U10973 (N_10973,N_9392,N_9462);
or U10974 (N_10974,N_9865,N_9629);
or U10975 (N_10975,N_9185,N_9586);
nor U10976 (N_10976,N_9883,N_9255);
xor U10977 (N_10977,N_9263,N_9585);
or U10978 (N_10978,N_9752,N_9717);
or U10979 (N_10979,N_9268,N_9409);
xnor U10980 (N_10980,N_9687,N_9660);
nand U10981 (N_10981,N_9102,N_9082);
nor U10982 (N_10982,N_9542,N_9068);
xor U10983 (N_10983,N_9696,N_9671);
nor U10984 (N_10984,N_9279,N_9371);
and U10985 (N_10985,N_9520,N_9361);
nor U10986 (N_10986,N_9435,N_9633);
and U10987 (N_10987,N_9150,N_9083);
nand U10988 (N_10988,N_9191,N_9571);
nor U10989 (N_10989,N_9298,N_9477);
nor U10990 (N_10990,N_9269,N_9511);
and U10991 (N_10991,N_9116,N_9327);
and U10992 (N_10992,N_9774,N_9429);
and U10993 (N_10993,N_9570,N_9779);
or U10994 (N_10994,N_9295,N_9752);
or U10995 (N_10995,N_9300,N_9161);
and U10996 (N_10996,N_9293,N_9658);
xnor U10997 (N_10997,N_9255,N_9866);
xnor U10998 (N_10998,N_9913,N_9444);
and U10999 (N_10999,N_9304,N_9330);
or U11000 (N_11000,N_10057,N_10297);
or U11001 (N_11001,N_10402,N_10673);
or U11002 (N_11002,N_10375,N_10382);
or U11003 (N_11003,N_10159,N_10488);
and U11004 (N_11004,N_10181,N_10048);
nand U11005 (N_11005,N_10182,N_10022);
or U11006 (N_11006,N_10459,N_10859);
nor U11007 (N_11007,N_10699,N_10656);
xnor U11008 (N_11008,N_10323,N_10098);
xor U11009 (N_11009,N_10068,N_10661);
and U11010 (N_11010,N_10192,N_10920);
xor U11011 (N_11011,N_10506,N_10671);
nand U11012 (N_11012,N_10863,N_10199);
nand U11013 (N_11013,N_10019,N_10039);
and U11014 (N_11014,N_10038,N_10064);
or U11015 (N_11015,N_10964,N_10231);
and U11016 (N_11016,N_10155,N_10870);
nor U11017 (N_11017,N_10094,N_10585);
xor U11018 (N_11018,N_10701,N_10813);
nor U11019 (N_11019,N_10886,N_10674);
or U11020 (N_11020,N_10309,N_10467);
and U11021 (N_11021,N_10812,N_10534);
xor U11022 (N_11022,N_10493,N_10634);
or U11023 (N_11023,N_10911,N_10184);
xnor U11024 (N_11024,N_10356,N_10728);
nor U11025 (N_11025,N_10448,N_10265);
nand U11026 (N_11026,N_10059,N_10591);
or U11027 (N_11027,N_10500,N_10716);
or U11028 (N_11028,N_10945,N_10706);
xor U11029 (N_11029,N_10616,N_10052);
nor U11030 (N_11030,N_10028,N_10427);
xnor U11031 (N_11031,N_10594,N_10835);
and U11032 (N_11032,N_10403,N_10602);
nor U11033 (N_11033,N_10082,N_10274);
or U11034 (N_11034,N_10447,N_10625);
or U11035 (N_11035,N_10056,N_10487);
and U11036 (N_11036,N_10332,N_10775);
and U11037 (N_11037,N_10531,N_10908);
nor U11038 (N_11038,N_10814,N_10243);
xnor U11039 (N_11039,N_10700,N_10419);
nor U11040 (N_11040,N_10769,N_10593);
xor U11041 (N_11041,N_10313,N_10854);
and U11042 (N_11042,N_10472,N_10643);
xor U11043 (N_11043,N_10917,N_10832);
xnor U11044 (N_11044,N_10906,N_10826);
nor U11045 (N_11045,N_10977,N_10874);
or U11046 (N_11046,N_10357,N_10291);
nor U11047 (N_11047,N_10363,N_10605);
and U11048 (N_11048,N_10404,N_10724);
xor U11049 (N_11049,N_10330,N_10202);
and U11050 (N_11050,N_10810,N_10709);
nor U11051 (N_11051,N_10461,N_10954);
or U11052 (N_11052,N_10370,N_10936);
and U11053 (N_11053,N_10926,N_10049);
or U11054 (N_11054,N_10755,N_10040);
nand U11055 (N_11055,N_10899,N_10209);
and U11056 (N_11056,N_10953,N_10512);
xnor U11057 (N_11057,N_10617,N_10836);
and U11058 (N_11058,N_10136,N_10258);
or U11059 (N_11059,N_10409,N_10688);
nand U11060 (N_11060,N_10973,N_10750);
and U11061 (N_11061,N_10205,N_10253);
or U11062 (N_11062,N_10008,N_10823);
nand U11063 (N_11063,N_10766,N_10023);
or U11064 (N_11064,N_10809,N_10799);
nor U11065 (N_11065,N_10140,N_10930);
nand U11066 (N_11066,N_10387,N_10690);
nor U11067 (N_11067,N_10508,N_10934);
and U11068 (N_11068,N_10635,N_10360);
nand U11069 (N_11069,N_10212,N_10221);
or U11070 (N_11070,N_10322,N_10670);
xor U11071 (N_11071,N_10552,N_10760);
nand U11072 (N_11072,N_10123,N_10443);
or U11073 (N_11073,N_10245,N_10583);
or U11074 (N_11074,N_10905,N_10868);
or U11075 (N_11075,N_10751,N_10565);
and U11076 (N_11076,N_10173,N_10203);
xnor U11077 (N_11077,N_10511,N_10818);
or U11078 (N_11078,N_10691,N_10067);
and U11079 (N_11079,N_10757,N_10302);
nor U11080 (N_11080,N_10385,N_10948);
nor U11081 (N_11081,N_10995,N_10311);
nand U11082 (N_11082,N_10228,N_10090);
or U11083 (N_11083,N_10430,N_10984);
and U11084 (N_11084,N_10767,N_10485);
nand U11085 (N_11085,N_10029,N_10846);
nand U11086 (N_11086,N_10949,N_10933);
nand U11087 (N_11087,N_10986,N_10663);
xor U11088 (N_11088,N_10218,N_10097);
and U11089 (N_11089,N_10131,N_10120);
or U11090 (N_11090,N_10147,N_10841);
and U11091 (N_11091,N_10843,N_10058);
or U11092 (N_11092,N_10020,N_10395);
nand U11093 (N_11093,N_10907,N_10478);
nor U11094 (N_11094,N_10093,N_10392);
xnor U11095 (N_11095,N_10269,N_10237);
and U11096 (N_11096,N_10225,N_10574);
nand U11097 (N_11097,N_10236,N_10561);
or U11098 (N_11098,N_10956,N_10655);
and U11099 (N_11099,N_10983,N_10080);
nor U11100 (N_11100,N_10334,N_10994);
and U11101 (N_11101,N_10250,N_10292);
xnor U11102 (N_11102,N_10287,N_10925);
and U11103 (N_11103,N_10801,N_10808);
or U11104 (N_11104,N_10341,N_10503);
nand U11105 (N_11105,N_10185,N_10220);
nor U11106 (N_11106,N_10733,N_10646);
or U11107 (N_11107,N_10614,N_10328);
nand U11108 (N_11108,N_10527,N_10229);
nor U11109 (N_11109,N_10932,N_10647);
or U11110 (N_11110,N_10086,N_10743);
nor U11111 (N_11111,N_10279,N_10371);
xor U11112 (N_11112,N_10536,N_10969);
nand U11113 (N_11113,N_10825,N_10036);
and U11114 (N_11114,N_10103,N_10677);
and U11115 (N_11115,N_10833,N_10262);
or U11116 (N_11116,N_10777,N_10384);
or U11117 (N_11117,N_10460,N_10439);
xnor U11118 (N_11118,N_10303,N_10551);
nand U11119 (N_11119,N_10543,N_10003);
xnor U11120 (N_11120,N_10620,N_10352);
xnor U11121 (N_11121,N_10422,N_10014);
xnor U11122 (N_11122,N_10495,N_10326);
or U11123 (N_11123,N_10180,N_10072);
nand U11124 (N_11124,N_10590,N_10013);
or U11125 (N_11125,N_10861,N_10877);
xnor U11126 (N_11126,N_10227,N_10687);
or U11127 (N_11127,N_10464,N_10664);
xor U11128 (N_11128,N_10268,N_10373);
or U11129 (N_11129,N_10164,N_10248);
xor U11130 (N_11130,N_10501,N_10062);
nor U11131 (N_11131,N_10657,N_10736);
nor U11132 (N_11132,N_10931,N_10424);
and U11133 (N_11133,N_10061,N_10758);
nand U11134 (N_11134,N_10756,N_10803);
nand U11135 (N_11135,N_10607,N_10214);
and U11136 (N_11136,N_10513,N_10923);
and U11137 (N_11137,N_10742,N_10662);
xor U11138 (N_11138,N_10586,N_10577);
nor U11139 (N_11139,N_10596,N_10009);
or U11140 (N_11140,N_10284,N_10329);
xor U11141 (N_11141,N_10075,N_10668);
nand U11142 (N_11142,N_10368,N_10795);
nor U11143 (N_11143,N_10183,N_10918);
nor U11144 (N_11144,N_10108,N_10942);
nor U11145 (N_11145,N_10532,N_10649);
xor U11146 (N_11146,N_10016,N_10894);
nand U11147 (N_11147,N_10796,N_10871);
nor U11148 (N_11148,N_10723,N_10989);
or U11149 (N_11149,N_10007,N_10615);
nand U11150 (N_11150,N_10622,N_10981);
and U11151 (N_11151,N_10520,N_10266);
xor U11152 (N_11152,N_10978,N_10828);
or U11153 (N_11153,N_10276,N_10790);
nor U11154 (N_11154,N_10083,N_10963);
and U11155 (N_11155,N_10654,N_10378);
nand U11156 (N_11156,N_10119,N_10141);
or U11157 (N_11157,N_10216,N_10955);
and U11158 (N_11158,N_10484,N_10428);
and U11159 (N_11159,N_10372,N_10351);
xor U11160 (N_11160,N_10912,N_10738);
and U11161 (N_11161,N_10537,N_10306);
nor U11162 (N_11162,N_10299,N_10466);
and U11163 (N_11163,N_10629,N_10554);
nand U11164 (N_11164,N_10000,N_10698);
xor U11165 (N_11165,N_10126,N_10914);
or U11166 (N_11166,N_10928,N_10047);
nor U11167 (N_11167,N_10314,N_10881);
nand U11168 (N_11168,N_10974,N_10855);
nand U11169 (N_11169,N_10754,N_10869);
xor U11170 (N_11170,N_10471,N_10584);
and U11171 (N_11171,N_10707,N_10713);
xor U11172 (N_11172,N_10711,N_10374);
xor U11173 (N_11173,N_10272,N_10325);
or U11174 (N_11174,N_10158,N_10473);
nand U11175 (N_11175,N_10415,N_10421);
nor U11176 (N_11176,N_10069,N_10800);
or U11177 (N_11177,N_10337,N_10358);
xor U11178 (N_11178,N_10442,N_10134);
xor U11179 (N_11179,N_10437,N_10475);
nand U11180 (N_11180,N_10633,N_10542);
nand U11181 (N_11181,N_10689,N_10702);
nand U11182 (N_11182,N_10129,N_10436);
and U11183 (N_11183,N_10568,N_10027);
or U11184 (N_11184,N_10021,N_10610);
and U11185 (N_11185,N_10477,N_10504);
nor U11186 (N_11186,N_10658,N_10366);
nor U11187 (N_11187,N_10365,N_10910);
nor U11188 (N_11188,N_10919,N_10962);
xnor U11189 (N_11189,N_10765,N_10230);
nor U11190 (N_11190,N_10850,N_10667);
nand U11191 (N_11191,N_10544,N_10324);
or U11192 (N_11192,N_10211,N_10012);
nand U11193 (N_11193,N_10940,N_10458);
nand U11194 (N_11194,N_10349,N_10010);
xor U11195 (N_11195,N_10883,N_10223);
xor U11196 (N_11196,N_10939,N_10148);
and U11197 (N_11197,N_10256,N_10824);
nor U11198 (N_11198,N_10556,N_10408);
and U11199 (N_11199,N_10597,N_10224);
nor U11200 (N_11200,N_10496,N_10417);
nor U11201 (N_11201,N_10451,N_10891);
and U11202 (N_11202,N_10095,N_10065);
and U11203 (N_11203,N_10096,N_10710);
nand U11204 (N_11204,N_10522,N_10239);
and U11205 (N_11205,N_10102,N_10416);
nor U11206 (N_11206,N_10867,N_10927);
or U11207 (N_11207,N_10862,N_10222);
or U11208 (N_11208,N_10582,N_10063);
nor U11209 (N_11209,N_10452,N_10393);
nand U11210 (N_11210,N_10208,N_10996);
nor U11211 (N_11211,N_10566,N_10077);
or U11212 (N_11212,N_10347,N_10720);
nor U11213 (N_11213,N_10569,N_10839);
nor U11214 (N_11214,N_10971,N_10830);
nand U11215 (N_11215,N_10338,N_10696);
and U11216 (N_11216,N_10780,N_10559);
nand U11217 (N_11217,N_10457,N_10619);
and U11218 (N_11218,N_10054,N_10335);
and U11219 (N_11219,N_10860,N_10275);
and U11220 (N_11220,N_10315,N_10191);
nand U11221 (N_11221,N_10290,N_10686);
and U11222 (N_11222,N_10684,N_10845);
nor U11223 (N_11223,N_10345,N_10423);
nand U11224 (N_11224,N_10987,N_10492);
nand U11225 (N_11225,N_10782,N_10893);
and U11226 (N_11226,N_10748,N_10901);
or U11227 (N_11227,N_10336,N_10429);
or U11228 (N_11228,N_10331,N_10557);
and U11229 (N_11229,N_10154,N_10186);
or U11230 (N_11230,N_10412,N_10637);
nand U11231 (N_11231,N_10613,N_10172);
and U11232 (N_11232,N_10916,N_10241);
nand U11233 (N_11233,N_10787,N_10117);
or U11234 (N_11234,N_10529,N_10175);
and U11235 (N_11235,N_10353,N_10676);
xor U11236 (N_11236,N_10091,N_10957);
and U11237 (N_11237,N_10618,N_10641);
or U11238 (N_11238,N_10035,N_10648);
nor U11239 (N_11239,N_10479,N_10571);
and U11240 (N_11240,N_10263,N_10609);
xor U11241 (N_11241,N_10307,N_10132);
xnor U11242 (N_11242,N_10727,N_10514);
or U11243 (N_11243,N_10252,N_10006);
nand U11244 (N_11244,N_10895,N_10340);
and U11245 (N_11245,N_10805,N_10078);
and U11246 (N_11246,N_10163,N_10296);
xor U11247 (N_11247,N_10398,N_10197);
xnor U11248 (N_11248,N_10864,N_10413);
and U11249 (N_11249,N_10234,N_10695);
xnor U11250 (N_11250,N_10773,N_10903);
nand U11251 (N_11251,N_10201,N_10762);
xor U11252 (N_11252,N_10545,N_10187);
nor U11253 (N_11253,N_10226,N_10866);
or U11254 (N_11254,N_10879,N_10246);
nand U11255 (N_11255,N_10456,N_10819);
or U11256 (N_11256,N_10207,N_10139);
xnor U11257 (N_11257,N_10792,N_10420);
nand U11258 (N_11258,N_10763,N_10547);
nor U11259 (N_11259,N_10261,N_10213);
and U11260 (N_11260,N_10235,N_10922);
nand U11261 (N_11261,N_10505,N_10741);
nand U11262 (N_11262,N_10632,N_10746);
nor U11263 (N_11263,N_10037,N_10364);
xnor U11264 (N_11264,N_10270,N_10215);
and U11265 (N_11265,N_10138,N_10887);
or U11266 (N_11266,N_10242,N_10598);
nand U11267 (N_11267,N_10359,N_10576);
and U11268 (N_11268,N_10652,N_10101);
or U11269 (N_11269,N_10462,N_10238);
nand U11270 (N_11270,N_10752,N_10169);
nor U11271 (N_11271,N_10998,N_10200);
xor U11272 (N_11272,N_10829,N_10606);
nor U11273 (N_11273,N_10526,N_10703);
and U11274 (N_11274,N_10491,N_10642);
or U11275 (N_11275,N_10286,N_10749);
nand U11276 (N_11276,N_10721,N_10951);
nand U11277 (N_11277,N_10289,N_10950);
xor U11278 (N_11278,N_10188,N_10502);
xnor U11279 (N_11279,N_10446,N_10118);
nand U11280 (N_11280,N_10143,N_10761);
nor U11281 (N_11281,N_10560,N_10152);
nor U11282 (N_11282,N_10444,N_10601);
and U11283 (N_11283,N_10426,N_10960);
and U11284 (N_11284,N_10383,N_10251);
or U11285 (N_11285,N_10639,N_10588);
and U11286 (N_11286,N_10876,N_10320);
and U11287 (N_11287,N_10438,N_10515);
nand U11288 (N_11288,N_10898,N_10913);
xnor U11289 (N_11289,N_10778,N_10644);
xor U11290 (N_11290,N_10011,N_10627);
xor U11291 (N_11291,N_10549,N_10849);
nor U11292 (N_11292,N_10562,N_10030);
nand U11293 (N_11293,N_10482,N_10445);
xor U11294 (N_11294,N_10784,N_10575);
nand U11295 (N_11295,N_10257,N_10573);
xnor U11296 (N_11296,N_10342,N_10033);
nor U11297 (N_11297,N_10198,N_10628);
xor U11298 (N_11298,N_10425,N_10807);
and U11299 (N_11299,N_10831,N_10285);
nor U11300 (N_11300,N_10947,N_10481);
nand U11301 (N_11301,N_10785,N_10781);
nor U11302 (N_11302,N_10463,N_10317);
nand U11303 (N_11303,N_10050,N_10171);
nor U11304 (N_11304,N_10516,N_10278);
nor U11305 (N_11305,N_10400,N_10685);
and U11306 (N_11306,N_10024,N_10260);
and U11307 (N_11307,N_10675,N_10450);
nor U11308 (N_11308,N_10937,N_10961);
or U11309 (N_11309,N_10985,N_10494);
and U11310 (N_11310,N_10884,N_10717);
and U11311 (N_11311,N_10089,N_10600);
nand U11312 (N_11312,N_10546,N_10381);
and U11313 (N_11313,N_10653,N_10092);
xnor U11314 (N_11314,N_10776,N_10411);
xor U11315 (N_11315,N_10110,N_10247);
xnor U11316 (N_11316,N_10672,N_10681);
and U11317 (N_11317,N_10354,N_10592);
and U11318 (N_11318,N_10853,N_10683);
nor U11319 (N_11319,N_10017,N_10298);
xor U11320 (N_11320,N_10304,N_10764);
or U11321 (N_11321,N_10194,N_10921);
xor U11322 (N_11322,N_10145,N_10004);
or U11323 (N_11323,N_10572,N_10390);
nand U11324 (N_11324,N_10770,N_10844);
and U11325 (N_11325,N_10924,N_10518);
nor U11326 (N_11326,N_10791,N_10031);
xor U11327 (N_11327,N_10348,N_10783);
xnor U11328 (N_11328,N_10878,N_10680);
and U11329 (N_11329,N_10204,N_10517);
nor U11330 (N_11330,N_10970,N_10233);
xnor U11331 (N_11331,N_10431,N_10734);
and U11332 (N_11332,N_10693,N_10705);
or U11333 (N_11333,N_10465,N_10165);
nand U11334 (N_11334,N_10255,N_10449);
nand U11335 (N_11335,N_10088,N_10885);
xor U11336 (N_11336,N_10277,N_10470);
nand U11337 (N_11337,N_10333,N_10564);
nand U11338 (N_11338,N_10660,N_10509);
nand U11339 (N_11339,N_10640,N_10821);
xor U11340 (N_11340,N_10168,N_10608);
xnor U11341 (N_11341,N_10650,N_10367);
and U11342 (N_11342,N_10730,N_10966);
and U11343 (N_11343,N_10087,N_10704);
or U11344 (N_11344,N_10414,N_10872);
and U11345 (N_11345,N_10774,N_10135);
xnor U11346 (N_11346,N_10838,N_10679);
and U11347 (N_11347,N_10745,N_10909);
xnor U11348 (N_11348,N_10682,N_10972);
nand U11349 (N_11349,N_10167,N_10666);
xor U11350 (N_11350,N_10490,N_10889);
and U11351 (N_11351,N_10271,N_10521);
xor U11352 (N_11352,N_10935,N_10308);
or U11353 (N_11353,N_10399,N_10100);
and U11354 (N_11354,N_10070,N_10476);
and U11355 (N_11355,N_10651,N_10160);
or U11356 (N_11356,N_10804,N_10524);
nand U11357 (N_11357,N_10283,N_10162);
xor U11358 (N_11358,N_10580,N_10817);
nand U11359 (N_11359,N_10697,N_10993);
nor U11360 (N_11360,N_10979,N_10759);
nor U11361 (N_11361,N_10708,N_10997);
xor U11362 (N_11362,N_10469,N_10725);
xnor U11363 (N_11363,N_10210,N_10567);
nor U11364 (N_11364,N_10944,N_10820);
nand U11365 (N_11365,N_10842,N_10380);
nand U11366 (N_11366,N_10361,N_10873);
nor U11367 (N_11367,N_10797,N_10386);
and U11368 (N_11368,N_10599,N_10137);
nor U11369 (N_11369,N_10788,N_10176);
xor U11370 (N_11370,N_10896,N_10305);
nor U11371 (N_11371,N_10786,N_10888);
nor U11372 (N_11372,N_10046,N_10249);
xnor U11373 (N_11373,N_10975,N_10281);
and U11374 (N_11374,N_10455,N_10043);
and U11375 (N_11375,N_10857,N_10530);
or U11376 (N_11376,N_10025,N_10959);
xor U11377 (N_11377,N_10179,N_10045);
or U11378 (N_11378,N_10254,N_10486);
and U11379 (N_11379,N_10579,N_10771);
or U11380 (N_11380,N_10865,N_10106);
xor U11381 (N_11381,N_10938,N_10161);
nand U11382 (N_11382,N_10541,N_10636);
nand U11383 (N_11383,N_10692,N_10915);
and U11384 (N_11384,N_10084,N_10044);
nor U11385 (N_11385,N_10312,N_10121);
nor U11386 (N_11386,N_10992,N_10267);
nand U11387 (N_11387,N_10999,N_10005);
nor U11388 (N_11388,N_10779,N_10076);
or U11389 (N_11389,N_10377,N_10193);
and U11390 (N_11390,N_10578,N_10976);
or U11391 (N_11391,N_10041,N_10405);
and U11392 (N_11392,N_10104,N_10410);
nand U11393 (N_11393,N_10474,N_10125);
nor U11394 (N_11394,N_10714,N_10499);
nor U11395 (N_11395,N_10665,N_10669);
nand U11396 (N_11396,N_10032,N_10418);
or U11397 (N_11397,N_10264,N_10540);
or U11398 (N_11398,N_10510,N_10074);
or U11399 (N_11399,N_10638,N_10166);
or U11400 (N_11400,N_10150,N_10107);
xor U11401 (N_11401,N_10882,N_10880);
nand U11402 (N_11402,N_10834,N_10624);
nor U11403 (N_11403,N_10732,N_10127);
and U11404 (N_11404,N_10454,N_10406);
nor U11405 (N_11405,N_10929,N_10719);
xnor U11406 (N_11406,N_10114,N_10369);
and U11407 (N_11407,N_10611,N_10435);
and U11408 (N_11408,N_10153,N_10806);
nor U11409 (N_11409,N_10051,N_10827);
or U11410 (N_11410,N_10060,N_10316);
xor U11411 (N_11411,N_10965,N_10982);
and U11412 (N_11412,N_10645,N_10768);
or U11413 (N_11413,N_10079,N_10396);
nor U11414 (N_11414,N_10388,N_10301);
or U11415 (N_11415,N_10802,N_10563);
nand U11416 (N_11416,N_10122,N_10085);
nand U11417 (N_11417,N_10968,N_10282);
and U11418 (N_11418,N_10897,N_10798);
and U11419 (N_11419,N_10731,N_10071);
nor U11420 (N_11420,N_10902,N_10026);
and U11421 (N_11421,N_10535,N_10310);
or U11422 (N_11422,N_10538,N_10124);
and U11423 (N_11423,N_10837,N_10659);
xnor U11424 (N_11424,N_10507,N_10389);
and U11425 (N_11425,N_10144,N_10177);
or U11426 (N_11426,N_10811,N_10483);
xor U11427 (N_11427,N_10295,N_10497);
nand U11428 (N_11428,N_10397,N_10190);
and U11429 (N_11429,N_10753,N_10852);
and U11430 (N_11430,N_10001,N_10815);
and U11431 (N_11431,N_10189,N_10816);
nor U11432 (N_11432,N_10848,N_10595);
nand U11433 (N_11433,N_10990,N_10892);
xnor U11434 (N_11434,N_10339,N_10018);
and U11435 (N_11435,N_10081,N_10300);
or U11436 (N_11436,N_10318,N_10772);
nor U11437 (N_11437,N_10142,N_10875);
nor U11438 (N_11438,N_10157,N_10480);
and U11439 (N_11439,N_10581,N_10943);
xnor U11440 (N_11440,N_10346,N_10146);
or U11441 (N_11441,N_10498,N_10321);
or U11442 (N_11442,N_10362,N_10539);
nand U11443 (N_11443,N_10712,N_10055);
nand U11444 (N_11444,N_10468,N_10991);
xnor U11445 (N_11445,N_10739,N_10570);
or U11446 (N_11446,N_10678,N_10952);
xnor U11447 (N_11447,N_10343,N_10206);
nor U11448 (N_11448,N_10988,N_10111);
and U11449 (N_11449,N_10822,N_10735);
and U11450 (N_11450,N_10128,N_10550);
xnor U11451 (N_11451,N_10626,N_10453);
nor U11452 (N_11452,N_10623,N_10604);
and U11453 (N_11453,N_10718,N_10273);
nor U11454 (N_11454,N_10244,N_10904);
xnor U11455 (N_11455,N_10015,N_10528);
or U11456 (N_11456,N_10099,N_10113);
xor U11457 (N_11457,N_10066,N_10433);
or U11458 (N_11458,N_10553,N_10344);
nor U11459 (N_11459,N_10555,N_10280);
and U11460 (N_11460,N_10151,N_10432);
xor U11461 (N_11461,N_10109,N_10196);
or U11462 (N_11462,N_10407,N_10630);
nand U11463 (N_11463,N_10747,N_10694);
nand U11464 (N_11464,N_10533,N_10350);
xnor U11465 (N_11465,N_10858,N_10401);
xor U11466 (N_11466,N_10294,N_10073);
nor U11467 (N_11467,N_10523,N_10105);
nor U11468 (N_11468,N_10946,N_10489);
xnor U11469 (N_11469,N_10729,N_10737);
and U11470 (N_11470,N_10548,N_10441);
nand U11471 (N_11471,N_10112,N_10434);
and U11472 (N_11472,N_10980,N_10034);
nor U11473 (N_11473,N_10133,N_10293);
nand U11474 (N_11474,N_10631,N_10195);
nor U11475 (N_11475,N_10890,N_10900);
nor U11476 (N_11476,N_10603,N_10587);
nand U11477 (N_11477,N_10440,N_10319);
xor U11478 (N_11478,N_10219,N_10130);
nor U11479 (N_11479,N_10232,N_10170);
nor U11480 (N_11480,N_10793,N_10217);
or U11481 (N_11481,N_10840,N_10856);
or U11482 (N_11482,N_10847,N_10053);
or U11483 (N_11483,N_10391,N_10394);
nand U11484 (N_11484,N_10740,N_10715);
nand U11485 (N_11485,N_10288,N_10355);
nand U11486 (N_11486,N_10744,N_10149);
nor U11487 (N_11487,N_10794,N_10851);
nand U11488 (N_11488,N_10958,N_10002);
nand U11489 (N_11489,N_10941,N_10376);
nand U11490 (N_11490,N_10259,N_10558);
or U11491 (N_11491,N_10612,N_10156);
nand U11492 (N_11492,N_10589,N_10327);
xnor U11493 (N_11493,N_10519,N_10726);
or U11494 (N_11494,N_10789,N_10115);
nor U11495 (N_11495,N_10379,N_10042);
nand U11496 (N_11496,N_10240,N_10525);
nand U11497 (N_11497,N_10722,N_10178);
and U11498 (N_11498,N_10621,N_10174);
nand U11499 (N_11499,N_10116,N_10967);
xnor U11500 (N_11500,N_10947,N_10952);
or U11501 (N_11501,N_10776,N_10443);
nand U11502 (N_11502,N_10602,N_10775);
nor U11503 (N_11503,N_10640,N_10544);
or U11504 (N_11504,N_10144,N_10783);
or U11505 (N_11505,N_10306,N_10270);
nand U11506 (N_11506,N_10990,N_10615);
nand U11507 (N_11507,N_10818,N_10388);
nand U11508 (N_11508,N_10742,N_10100);
or U11509 (N_11509,N_10676,N_10072);
nand U11510 (N_11510,N_10636,N_10312);
nand U11511 (N_11511,N_10832,N_10289);
xor U11512 (N_11512,N_10631,N_10705);
and U11513 (N_11513,N_10088,N_10930);
xor U11514 (N_11514,N_10742,N_10361);
nand U11515 (N_11515,N_10191,N_10631);
and U11516 (N_11516,N_10105,N_10081);
nor U11517 (N_11517,N_10629,N_10770);
or U11518 (N_11518,N_10313,N_10672);
xnor U11519 (N_11519,N_10035,N_10697);
xor U11520 (N_11520,N_10011,N_10972);
nand U11521 (N_11521,N_10063,N_10021);
or U11522 (N_11522,N_10914,N_10810);
nor U11523 (N_11523,N_10776,N_10267);
and U11524 (N_11524,N_10560,N_10947);
nor U11525 (N_11525,N_10836,N_10793);
nor U11526 (N_11526,N_10795,N_10269);
nor U11527 (N_11527,N_10735,N_10464);
nand U11528 (N_11528,N_10949,N_10450);
nand U11529 (N_11529,N_10806,N_10979);
nor U11530 (N_11530,N_10697,N_10257);
xnor U11531 (N_11531,N_10820,N_10634);
and U11532 (N_11532,N_10337,N_10653);
nand U11533 (N_11533,N_10806,N_10901);
and U11534 (N_11534,N_10030,N_10684);
and U11535 (N_11535,N_10962,N_10659);
and U11536 (N_11536,N_10098,N_10560);
nor U11537 (N_11537,N_10967,N_10017);
nand U11538 (N_11538,N_10916,N_10743);
and U11539 (N_11539,N_10124,N_10618);
nand U11540 (N_11540,N_10486,N_10805);
and U11541 (N_11541,N_10394,N_10548);
nor U11542 (N_11542,N_10737,N_10668);
nor U11543 (N_11543,N_10956,N_10959);
or U11544 (N_11544,N_10701,N_10097);
or U11545 (N_11545,N_10661,N_10434);
nor U11546 (N_11546,N_10377,N_10907);
or U11547 (N_11547,N_10856,N_10083);
and U11548 (N_11548,N_10900,N_10748);
and U11549 (N_11549,N_10315,N_10046);
and U11550 (N_11550,N_10957,N_10180);
nor U11551 (N_11551,N_10075,N_10791);
nand U11552 (N_11552,N_10050,N_10834);
nor U11553 (N_11553,N_10269,N_10303);
nor U11554 (N_11554,N_10049,N_10914);
or U11555 (N_11555,N_10210,N_10291);
nand U11556 (N_11556,N_10191,N_10296);
nor U11557 (N_11557,N_10894,N_10243);
xor U11558 (N_11558,N_10182,N_10513);
and U11559 (N_11559,N_10473,N_10544);
nor U11560 (N_11560,N_10482,N_10986);
and U11561 (N_11561,N_10944,N_10584);
xnor U11562 (N_11562,N_10244,N_10806);
and U11563 (N_11563,N_10110,N_10524);
xor U11564 (N_11564,N_10083,N_10972);
nand U11565 (N_11565,N_10588,N_10537);
nand U11566 (N_11566,N_10721,N_10368);
nand U11567 (N_11567,N_10490,N_10627);
or U11568 (N_11568,N_10710,N_10506);
xnor U11569 (N_11569,N_10579,N_10799);
nor U11570 (N_11570,N_10307,N_10017);
xnor U11571 (N_11571,N_10570,N_10886);
and U11572 (N_11572,N_10771,N_10526);
or U11573 (N_11573,N_10374,N_10665);
and U11574 (N_11574,N_10923,N_10847);
or U11575 (N_11575,N_10127,N_10171);
nor U11576 (N_11576,N_10378,N_10728);
nand U11577 (N_11577,N_10158,N_10796);
or U11578 (N_11578,N_10365,N_10876);
and U11579 (N_11579,N_10363,N_10796);
nor U11580 (N_11580,N_10961,N_10734);
xnor U11581 (N_11581,N_10946,N_10428);
nor U11582 (N_11582,N_10944,N_10508);
or U11583 (N_11583,N_10464,N_10632);
or U11584 (N_11584,N_10682,N_10286);
nand U11585 (N_11585,N_10584,N_10808);
or U11586 (N_11586,N_10845,N_10004);
xnor U11587 (N_11587,N_10955,N_10694);
xnor U11588 (N_11588,N_10200,N_10907);
and U11589 (N_11589,N_10283,N_10131);
and U11590 (N_11590,N_10910,N_10465);
nor U11591 (N_11591,N_10834,N_10399);
xnor U11592 (N_11592,N_10779,N_10146);
and U11593 (N_11593,N_10088,N_10684);
or U11594 (N_11594,N_10071,N_10820);
xor U11595 (N_11595,N_10989,N_10629);
xnor U11596 (N_11596,N_10883,N_10444);
and U11597 (N_11597,N_10307,N_10473);
nand U11598 (N_11598,N_10253,N_10911);
or U11599 (N_11599,N_10566,N_10639);
nor U11600 (N_11600,N_10782,N_10294);
xnor U11601 (N_11601,N_10501,N_10679);
nand U11602 (N_11602,N_10383,N_10896);
and U11603 (N_11603,N_10945,N_10830);
nor U11604 (N_11604,N_10238,N_10753);
nand U11605 (N_11605,N_10730,N_10398);
xor U11606 (N_11606,N_10543,N_10643);
nand U11607 (N_11607,N_10309,N_10702);
xnor U11608 (N_11608,N_10326,N_10164);
or U11609 (N_11609,N_10224,N_10872);
nand U11610 (N_11610,N_10572,N_10557);
and U11611 (N_11611,N_10748,N_10701);
nand U11612 (N_11612,N_10193,N_10558);
or U11613 (N_11613,N_10350,N_10209);
nand U11614 (N_11614,N_10503,N_10278);
or U11615 (N_11615,N_10269,N_10415);
xor U11616 (N_11616,N_10484,N_10593);
nand U11617 (N_11617,N_10930,N_10564);
or U11618 (N_11618,N_10112,N_10911);
nor U11619 (N_11619,N_10439,N_10347);
nor U11620 (N_11620,N_10098,N_10883);
nor U11621 (N_11621,N_10669,N_10431);
xor U11622 (N_11622,N_10511,N_10622);
and U11623 (N_11623,N_10935,N_10154);
or U11624 (N_11624,N_10284,N_10702);
or U11625 (N_11625,N_10293,N_10507);
or U11626 (N_11626,N_10853,N_10883);
nand U11627 (N_11627,N_10635,N_10852);
and U11628 (N_11628,N_10577,N_10798);
xnor U11629 (N_11629,N_10460,N_10856);
nand U11630 (N_11630,N_10463,N_10153);
nor U11631 (N_11631,N_10825,N_10076);
xnor U11632 (N_11632,N_10454,N_10581);
nor U11633 (N_11633,N_10780,N_10526);
nor U11634 (N_11634,N_10233,N_10810);
or U11635 (N_11635,N_10754,N_10506);
nor U11636 (N_11636,N_10677,N_10723);
or U11637 (N_11637,N_10181,N_10589);
nand U11638 (N_11638,N_10181,N_10628);
xor U11639 (N_11639,N_10916,N_10541);
nand U11640 (N_11640,N_10072,N_10437);
nor U11641 (N_11641,N_10449,N_10552);
nor U11642 (N_11642,N_10531,N_10592);
and U11643 (N_11643,N_10341,N_10388);
nor U11644 (N_11644,N_10781,N_10990);
xor U11645 (N_11645,N_10675,N_10443);
nand U11646 (N_11646,N_10881,N_10952);
nor U11647 (N_11647,N_10600,N_10014);
and U11648 (N_11648,N_10841,N_10605);
xnor U11649 (N_11649,N_10068,N_10428);
or U11650 (N_11650,N_10247,N_10040);
nand U11651 (N_11651,N_10928,N_10582);
nand U11652 (N_11652,N_10650,N_10998);
and U11653 (N_11653,N_10784,N_10702);
nand U11654 (N_11654,N_10610,N_10853);
xor U11655 (N_11655,N_10375,N_10603);
nor U11656 (N_11656,N_10220,N_10299);
nand U11657 (N_11657,N_10028,N_10099);
or U11658 (N_11658,N_10697,N_10738);
and U11659 (N_11659,N_10229,N_10951);
nand U11660 (N_11660,N_10884,N_10289);
xor U11661 (N_11661,N_10932,N_10384);
or U11662 (N_11662,N_10864,N_10486);
and U11663 (N_11663,N_10949,N_10391);
and U11664 (N_11664,N_10408,N_10212);
xnor U11665 (N_11665,N_10786,N_10299);
and U11666 (N_11666,N_10973,N_10125);
nand U11667 (N_11667,N_10372,N_10976);
nand U11668 (N_11668,N_10940,N_10669);
or U11669 (N_11669,N_10861,N_10277);
and U11670 (N_11670,N_10350,N_10813);
and U11671 (N_11671,N_10081,N_10035);
or U11672 (N_11672,N_10579,N_10795);
xnor U11673 (N_11673,N_10676,N_10110);
nand U11674 (N_11674,N_10939,N_10317);
and U11675 (N_11675,N_10093,N_10572);
or U11676 (N_11676,N_10104,N_10235);
or U11677 (N_11677,N_10712,N_10718);
or U11678 (N_11678,N_10552,N_10890);
nor U11679 (N_11679,N_10431,N_10783);
nor U11680 (N_11680,N_10153,N_10700);
or U11681 (N_11681,N_10060,N_10241);
nand U11682 (N_11682,N_10109,N_10166);
and U11683 (N_11683,N_10262,N_10585);
or U11684 (N_11684,N_10964,N_10836);
and U11685 (N_11685,N_10847,N_10982);
and U11686 (N_11686,N_10143,N_10989);
nor U11687 (N_11687,N_10623,N_10508);
and U11688 (N_11688,N_10844,N_10843);
nand U11689 (N_11689,N_10860,N_10835);
nand U11690 (N_11690,N_10582,N_10532);
or U11691 (N_11691,N_10825,N_10810);
or U11692 (N_11692,N_10512,N_10994);
or U11693 (N_11693,N_10420,N_10190);
nor U11694 (N_11694,N_10355,N_10290);
nand U11695 (N_11695,N_10220,N_10026);
and U11696 (N_11696,N_10324,N_10767);
xor U11697 (N_11697,N_10683,N_10960);
and U11698 (N_11698,N_10911,N_10607);
nor U11699 (N_11699,N_10542,N_10568);
and U11700 (N_11700,N_10901,N_10844);
xnor U11701 (N_11701,N_10540,N_10082);
or U11702 (N_11702,N_10180,N_10493);
and U11703 (N_11703,N_10037,N_10394);
nor U11704 (N_11704,N_10789,N_10119);
nor U11705 (N_11705,N_10263,N_10753);
nor U11706 (N_11706,N_10449,N_10851);
xnor U11707 (N_11707,N_10477,N_10468);
or U11708 (N_11708,N_10179,N_10507);
nand U11709 (N_11709,N_10289,N_10139);
and U11710 (N_11710,N_10102,N_10851);
and U11711 (N_11711,N_10559,N_10894);
or U11712 (N_11712,N_10001,N_10966);
nand U11713 (N_11713,N_10844,N_10188);
nand U11714 (N_11714,N_10330,N_10447);
xor U11715 (N_11715,N_10435,N_10685);
and U11716 (N_11716,N_10763,N_10430);
nand U11717 (N_11717,N_10904,N_10359);
xor U11718 (N_11718,N_10770,N_10851);
and U11719 (N_11719,N_10982,N_10731);
or U11720 (N_11720,N_10893,N_10140);
and U11721 (N_11721,N_10577,N_10974);
or U11722 (N_11722,N_10241,N_10776);
and U11723 (N_11723,N_10246,N_10108);
or U11724 (N_11724,N_10619,N_10387);
xor U11725 (N_11725,N_10263,N_10906);
nor U11726 (N_11726,N_10337,N_10731);
xor U11727 (N_11727,N_10933,N_10544);
nand U11728 (N_11728,N_10234,N_10624);
and U11729 (N_11729,N_10944,N_10925);
xnor U11730 (N_11730,N_10054,N_10513);
nand U11731 (N_11731,N_10405,N_10959);
or U11732 (N_11732,N_10711,N_10257);
and U11733 (N_11733,N_10358,N_10866);
or U11734 (N_11734,N_10049,N_10630);
nand U11735 (N_11735,N_10283,N_10760);
nor U11736 (N_11736,N_10478,N_10372);
or U11737 (N_11737,N_10438,N_10861);
xnor U11738 (N_11738,N_10529,N_10873);
and U11739 (N_11739,N_10839,N_10653);
nand U11740 (N_11740,N_10715,N_10809);
or U11741 (N_11741,N_10246,N_10091);
or U11742 (N_11742,N_10097,N_10843);
and U11743 (N_11743,N_10138,N_10141);
and U11744 (N_11744,N_10088,N_10201);
nand U11745 (N_11745,N_10302,N_10283);
nor U11746 (N_11746,N_10639,N_10194);
and U11747 (N_11747,N_10964,N_10015);
or U11748 (N_11748,N_10267,N_10105);
nand U11749 (N_11749,N_10609,N_10021);
nor U11750 (N_11750,N_10387,N_10488);
nor U11751 (N_11751,N_10592,N_10310);
nor U11752 (N_11752,N_10704,N_10397);
and U11753 (N_11753,N_10897,N_10161);
and U11754 (N_11754,N_10958,N_10786);
or U11755 (N_11755,N_10819,N_10994);
or U11756 (N_11756,N_10618,N_10157);
xor U11757 (N_11757,N_10330,N_10523);
and U11758 (N_11758,N_10464,N_10856);
nor U11759 (N_11759,N_10613,N_10240);
nor U11760 (N_11760,N_10898,N_10583);
or U11761 (N_11761,N_10323,N_10455);
xor U11762 (N_11762,N_10862,N_10818);
nand U11763 (N_11763,N_10959,N_10392);
nand U11764 (N_11764,N_10060,N_10855);
xor U11765 (N_11765,N_10783,N_10043);
or U11766 (N_11766,N_10858,N_10811);
or U11767 (N_11767,N_10497,N_10583);
nor U11768 (N_11768,N_10042,N_10208);
nand U11769 (N_11769,N_10465,N_10739);
nor U11770 (N_11770,N_10573,N_10644);
or U11771 (N_11771,N_10308,N_10795);
xor U11772 (N_11772,N_10608,N_10745);
or U11773 (N_11773,N_10376,N_10587);
nor U11774 (N_11774,N_10476,N_10775);
nand U11775 (N_11775,N_10665,N_10293);
and U11776 (N_11776,N_10076,N_10715);
xnor U11777 (N_11777,N_10944,N_10380);
and U11778 (N_11778,N_10781,N_10943);
or U11779 (N_11779,N_10334,N_10520);
and U11780 (N_11780,N_10189,N_10289);
or U11781 (N_11781,N_10916,N_10885);
xnor U11782 (N_11782,N_10847,N_10754);
and U11783 (N_11783,N_10715,N_10867);
nor U11784 (N_11784,N_10345,N_10347);
or U11785 (N_11785,N_10239,N_10362);
or U11786 (N_11786,N_10619,N_10695);
and U11787 (N_11787,N_10471,N_10065);
nor U11788 (N_11788,N_10424,N_10369);
or U11789 (N_11789,N_10408,N_10309);
xnor U11790 (N_11790,N_10026,N_10396);
nand U11791 (N_11791,N_10031,N_10760);
nand U11792 (N_11792,N_10304,N_10029);
nand U11793 (N_11793,N_10195,N_10642);
nand U11794 (N_11794,N_10486,N_10803);
nand U11795 (N_11795,N_10827,N_10362);
nor U11796 (N_11796,N_10616,N_10708);
or U11797 (N_11797,N_10760,N_10717);
xnor U11798 (N_11798,N_10597,N_10739);
and U11799 (N_11799,N_10442,N_10294);
nor U11800 (N_11800,N_10696,N_10760);
nand U11801 (N_11801,N_10080,N_10501);
nor U11802 (N_11802,N_10747,N_10077);
nand U11803 (N_11803,N_10729,N_10756);
and U11804 (N_11804,N_10837,N_10873);
nand U11805 (N_11805,N_10344,N_10198);
nand U11806 (N_11806,N_10781,N_10270);
and U11807 (N_11807,N_10805,N_10422);
nor U11808 (N_11808,N_10119,N_10331);
xor U11809 (N_11809,N_10117,N_10769);
xor U11810 (N_11810,N_10584,N_10302);
nor U11811 (N_11811,N_10898,N_10881);
and U11812 (N_11812,N_10989,N_10761);
nand U11813 (N_11813,N_10304,N_10549);
nand U11814 (N_11814,N_10718,N_10256);
xor U11815 (N_11815,N_10505,N_10805);
nand U11816 (N_11816,N_10401,N_10746);
nor U11817 (N_11817,N_10031,N_10951);
nand U11818 (N_11818,N_10221,N_10069);
and U11819 (N_11819,N_10792,N_10852);
and U11820 (N_11820,N_10221,N_10343);
and U11821 (N_11821,N_10974,N_10306);
nor U11822 (N_11822,N_10405,N_10541);
or U11823 (N_11823,N_10792,N_10546);
nand U11824 (N_11824,N_10985,N_10117);
nand U11825 (N_11825,N_10096,N_10189);
or U11826 (N_11826,N_10605,N_10610);
xnor U11827 (N_11827,N_10971,N_10847);
and U11828 (N_11828,N_10095,N_10666);
and U11829 (N_11829,N_10655,N_10741);
nor U11830 (N_11830,N_10349,N_10357);
nor U11831 (N_11831,N_10010,N_10138);
and U11832 (N_11832,N_10390,N_10446);
nand U11833 (N_11833,N_10849,N_10906);
nor U11834 (N_11834,N_10588,N_10924);
or U11835 (N_11835,N_10587,N_10818);
or U11836 (N_11836,N_10388,N_10063);
xnor U11837 (N_11837,N_10012,N_10530);
nor U11838 (N_11838,N_10286,N_10083);
xnor U11839 (N_11839,N_10239,N_10703);
and U11840 (N_11840,N_10761,N_10401);
nor U11841 (N_11841,N_10668,N_10377);
nand U11842 (N_11842,N_10904,N_10875);
xnor U11843 (N_11843,N_10928,N_10636);
or U11844 (N_11844,N_10572,N_10358);
xor U11845 (N_11845,N_10544,N_10494);
or U11846 (N_11846,N_10178,N_10493);
nor U11847 (N_11847,N_10015,N_10989);
and U11848 (N_11848,N_10332,N_10484);
xor U11849 (N_11849,N_10859,N_10311);
xor U11850 (N_11850,N_10533,N_10975);
and U11851 (N_11851,N_10038,N_10149);
nor U11852 (N_11852,N_10005,N_10775);
and U11853 (N_11853,N_10895,N_10790);
xnor U11854 (N_11854,N_10537,N_10672);
xor U11855 (N_11855,N_10275,N_10991);
nand U11856 (N_11856,N_10848,N_10188);
nand U11857 (N_11857,N_10738,N_10691);
and U11858 (N_11858,N_10159,N_10692);
nand U11859 (N_11859,N_10217,N_10436);
or U11860 (N_11860,N_10290,N_10888);
or U11861 (N_11861,N_10407,N_10408);
or U11862 (N_11862,N_10228,N_10328);
nor U11863 (N_11863,N_10378,N_10352);
nand U11864 (N_11864,N_10397,N_10038);
nand U11865 (N_11865,N_10015,N_10780);
and U11866 (N_11866,N_10915,N_10093);
nor U11867 (N_11867,N_10001,N_10301);
nor U11868 (N_11868,N_10857,N_10172);
and U11869 (N_11869,N_10495,N_10982);
or U11870 (N_11870,N_10887,N_10312);
and U11871 (N_11871,N_10208,N_10679);
nor U11872 (N_11872,N_10770,N_10633);
xnor U11873 (N_11873,N_10832,N_10666);
and U11874 (N_11874,N_10468,N_10083);
and U11875 (N_11875,N_10480,N_10626);
or U11876 (N_11876,N_10954,N_10425);
nand U11877 (N_11877,N_10200,N_10828);
xor U11878 (N_11878,N_10185,N_10321);
and U11879 (N_11879,N_10612,N_10606);
xor U11880 (N_11880,N_10157,N_10905);
and U11881 (N_11881,N_10338,N_10972);
and U11882 (N_11882,N_10015,N_10217);
and U11883 (N_11883,N_10508,N_10692);
and U11884 (N_11884,N_10246,N_10732);
or U11885 (N_11885,N_10061,N_10624);
and U11886 (N_11886,N_10478,N_10189);
or U11887 (N_11887,N_10185,N_10107);
nor U11888 (N_11888,N_10981,N_10400);
and U11889 (N_11889,N_10130,N_10535);
xor U11890 (N_11890,N_10837,N_10603);
nor U11891 (N_11891,N_10077,N_10638);
nor U11892 (N_11892,N_10868,N_10001);
and U11893 (N_11893,N_10897,N_10900);
and U11894 (N_11894,N_10558,N_10076);
nor U11895 (N_11895,N_10719,N_10278);
nor U11896 (N_11896,N_10776,N_10033);
or U11897 (N_11897,N_10497,N_10387);
xor U11898 (N_11898,N_10817,N_10710);
or U11899 (N_11899,N_10559,N_10632);
and U11900 (N_11900,N_10862,N_10042);
nor U11901 (N_11901,N_10899,N_10098);
and U11902 (N_11902,N_10341,N_10559);
and U11903 (N_11903,N_10071,N_10292);
xor U11904 (N_11904,N_10935,N_10844);
and U11905 (N_11905,N_10108,N_10286);
nor U11906 (N_11906,N_10362,N_10057);
nand U11907 (N_11907,N_10668,N_10107);
or U11908 (N_11908,N_10218,N_10172);
and U11909 (N_11909,N_10138,N_10016);
and U11910 (N_11910,N_10901,N_10304);
or U11911 (N_11911,N_10928,N_10630);
xor U11912 (N_11912,N_10296,N_10227);
and U11913 (N_11913,N_10064,N_10339);
nand U11914 (N_11914,N_10887,N_10046);
nor U11915 (N_11915,N_10010,N_10373);
or U11916 (N_11916,N_10534,N_10305);
xor U11917 (N_11917,N_10009,N_10627);
or U11918 (N_11918,N_10018,N_10606);
xor U11919 (N_11919,N_10282,N_10787);
nor U11920 (N_11920,N_10421,N_10170);
and U11921 (N_11921,N_10132,N_10877);
xnor U11922 (N_11922,N_10579,N_10627);
nand U11923 (N_11923,N_10106,N_10583);
xnor U11924 (N_11924,N_10368,N_10998);
or U11925 (N_11925,N_10812,N_10385);
or U11926 (N_11926,N_10908,N_10485);
nor U11927 (N_11927,N_10437,N_10280);
nor U11928 (N_11928,N_10706,N_10307);
nand U11929 (N_11929,N_10278,N_10340);
nand U11930 (N_11930,N_10222,N_10113);
nand U11931 (N_11931,N_10536,N_10278);
xor U11932 (N_11932,N_10146,N_10882);
nor U11933 (N_11933,N_10584,N_10684);
nand U11934 (N_11934,N_10937,N_10475);
and U11935 (N_11935,N_10974,N_10178);
or U11936 (N_11936,N_10737,N_10387);
or U11937 (N_11937,N_10976,N_10260);
xnor U11938 (N_11938,N_10683,N_10267);
nand U11939 (N_11939,N_10384,N_10105);
nor U11940 (N_11940,N_10944,N_10182);
nor U11941 (N_11941,N_10021,N_10991);
nand U11942 (N_11942,N_10534,N_10302);
or U11943 (N_11943,N_10489,N_10801);
xor U11944 (N_11944,N_10533,N_10399);
or U11945 (N_11945,N_10939,N_10542);
nand U11946 (N_11946,N_10215,N_10329);
nor U11947 (N_11947,N_10642,N_10746);
xnor U11948 (N_11948,N_10323,N_10297);
nor U11949 (N_11949,N_10877,N_10054);
nand U11950 (N_11950,N_10898,N_10058);
or U11951 (N_11951,N_10353,N_10708);
nand U11952 (N_11952,N_10893,N_10037);
nand U11953 (N_11953,N_10126,N_10636);
nand U11954 (N_11954,N_10770,N_10418);
and U11955 (N_11955,N_10904,N_10413);
xnor U11956 (N_11956,N_10519,N_10872);
nand U11957 (N_11957,N_10103,N_10281);
nor U11958 (N_11958,N_10790,N_10215);
and U11959 (N_11959,N_10789,N_10606);
nor U11960 (N_11960,N_10664,N_10705);
nand U11961 (N_11961,N_10640,N_10785);
nand U11962 (N_11962,N_10098,N_10246);
nor U11963 (N_11963,N_10618,N_10938);
nand U11964 (N_11964,N_10168,N_10845);
or U11965 (N_11965,N_10467,N_10887);
nand U11966 (N_11966,N_10091,N_10070);
nor U11967 (N_11967,N_10111,N_10816);
and U11968 (N_11968,N_10809,N_10300);
and U11969 (N_11969,N_10556,N_10498);
nor U11970 (N_11970,N_10261,N_10995);
nand U11971 (N_11971,N_10610,N_10300);
nor U11972 (N_11972,N_10350,N_10356);
or U11973 (N_11973,N_10061,N_10629);
and U11974 (N_11974,N_10392,N_10808);
xnor U11975 (N_11975,N_10075,N_10253);
nor U11976 (N_11976,N_10883,N_10561);
nor U11977 (N_11977,N_10708,N_10575);
nor U11978 (N_11978,N_10264,N_10627);
and U11979 (N_11979,N_10575,N_10551);
and U11980 (N_11980,N_10569,N_10295);
xor U11981 (N_11981,N_10431,N_10918);
nand U11982 (N_11982,N_10464,N_10667);
nor U11983 (N_11983,N_10996,N_10590);
nor U11984 (N_11984,N_10898,N_10737);
and U11985 (N_11985,N_10005,N_10080);
and U11986 (N_11986,N_10818,N_10808);
xor U11987 (N_11987,N_10166,N_10328);
and U11988 (N_11988,N_10150,N_10621);
nor U11989 (N_11989,N_10781,N_10059);
nand U11990 (N_11990,N_10890,N_10034);
nand U11991 (N_11991,N_10735,N_10277);
and U11992 (N_11992,N_10998,N_10172);
nand U11993 (N_11993,N_10962,N_10323);
nand U11994 (N_11994,N_10514,N_10551);
nor U11995 (N_11995,N_10163,N_10841);
or U11996 (N_11996,N_10726,N_10528);
and U11997 (N_11997,N_10014,N_10837);
or U11998 (N_11998,N_10915,N_10770);
or U11999 (N_11999,N_10195,N_10480);
xor U12000 (N_12000,N_11526,N_11764);
or U12001 (N_12001,N_11018,N_11354);
nand U12002 (N_12002,N_11810,N_11772);
nor U12003 (N_12003,N_11224,N_11799);
or U12004 (N_12004,N_11157,N_11501);
nor U12005 (N_12005,N_11162,N_11840);
nor U12006 (N_12006,N_11707,N_11051);
nor U12007 (N_12007,N_11771,N_11201);
nor U12008 (N_12008,N_11305,N_11386);
or U12009 (N_12009,N_11598,N_11984);
nor U12010 (N_12010,N_11602,N_11639);
or U12011 (N_12011,N_11829,N_11798);
nand U12012 (N_12012,N_11301,N_11485);
nand U12013 (N_12013,N_11628,N_11704);
xor U12014 (N_12014,N_11728,N_11767);
and U12015 (N_12015,N_11716,N_11642);
and U12016 (N_12016,N_11696,N_11794);
nor U12017 (N_12017,N_11076,N_11288);
or U12018 (N_12018,N_11291,N_11713);
and U12019 (N_12019,N_11721,N_11368);
or U12020 (N_12020,N_11872,N_11242);
nand U12021 (N_12021,N_11653,N_11910);
nor U12022 (N_12022,N_11035,N_11762);
or U12023 (N_12023,N_11117,N_11662);
or U12024 (N_12024,N_11650,N_11318);
nand U12025 (N_12025,N_11532,N_11904);
xor U12026 (N_12026,N_11362,N_11401);
nor U12027 (N_12027,N_11128,N_11583);
xnor U12028 (N_12028,N_11865,N_11766);
xnor U12029 (N_12029,N_11940,N_11471);
nor U12030 (N_12030,N_11922,N_11360);
or U12031 (N_12031,N_11751,N_11785);
xnor U12032 (N_12032,N_11547,N_11601);
or U12033 (N_12033,N_11879,N_11148);
xnor U12034 (N_12034,N_11052,N_11350);
and U12035 (N_12035,N_11021,N_11186);
or U12036 (N_12036,N_11392,N_11604);
nand U12037 (N_12037,N_11327,N_11285);
nor U12038 (N_12038,N_11325,N_11273);
or U12039 (N_12039,N_11137,N_11041);
nor U12040 (N_12040,N_11376,N_11197);
nand U12041 (N_12041,N_11786,N_11027);
or U12042 (N_12042,N_11812,N_11973);
xor U12043 (N_12043,N_11903,N_11050);
or U12044 (N_12044,N_11811,N_11093);
nand U12045 (N_12045,N_11830,N_11243);
nor U12046 (N_12046,N_11516,N_11121);
or U12047 (N_12047,N_11874,N_11080);
nand U12048 (N_12048,N_11723,N_11784);
xnor U12049 (N_12049,N_11249,N_11511);
or U12050 (N_12050,N_11993,N_11441);
and U12051 (N_12051,N_11084,N_11387);
nor U12052 (N_12052,N_11759,N_11096);
nand U12053 (N_12053,N_11010,N_11057);
and U12054 (N_12054,N_11695,N_11502);
or U12055 (N_12055,N_11341,N_11995);
nand U12056 (N_12056,N_11636,N_11232);
and U12057 (N_12057,N_11528,N_11176);
nand U12058 (N_12058,N_11374,N_11476);
or U12059 (N_12059,N_11550,N_11773);
xor U12060 (N_12060,N_11338,N_11870);
nand U12061 (N_12061,N_11311,N_11275);
nand U12062 (N_12062,N_11733,N_11355);
or U12063 (N_12063,N_11774,N_11174);
or U12064 (N_12064,N_11299,N_11134);
xor U12065 (N_12065,N_11692,N_11433);
nor U12066 (N_12066,N_11490,N_11573);
nand U12067 (N_12067,N_11103,N_11409);
nand U12068 (N_12068,N_11272,N_11938);
nand U12069 (N_12069,N_11383,N_11458);
nor U12070 (N_12070,N_11902,N_11506);
or U12071 (N_12071,N_11289,N_11730);
and U12072 (N_12072,N_11464,N_11608);
nor U12073 (N_12073,N_11711,N_11866);
nor U12074 (N_12074,N_11454,N_11564);
xor U12075 (N_12075,N_11935,N_11058);
nand U12076 (N_12076,N_11257,N_11722);
nand U12077 (N_12077,N_11167,N_11150);
xor U12078 (N_12078,N_11625,N_11432);
nor U12079 (N_12079,N_11655,N_11907);
nand U12080 (N_12080,N_11890,N_11312);
xor U12081 (N_12081,N_11620,N_11496);
nand U12082 (N_12082,N_11286,N_11385);
or U12083 (N_12083,N_11720,N_11482);
xor U12084 (N_12084,N_11280,N_11924);
and U12085 (N_12085,N_11859,N_11581);
nand U12086 (N_12086,N_11609,N_11748);
and U12087 (N_12087,N_11529,N_11073);
and U12088 (N_12088,N_11384,N_11406);
or U12089 (N_12089,N_11541,N_11893);
nand U12090 (N_12090,N_11947,N_11135);
or U12091 (N_12091,N_11488,N_11954);
nor U12092 (N_12092,N_11175,N_11576);
nand U12093 (N_12093,N_11146,N_11672);
nand U12094 (N_12094,N_11558,N_11208);
or U12095 (N_12095,N_11612,N_11055);
or U12096 (N_12096,N_11061,N_11792);
or U12097 (N_12097,N_11348,N_11323);
and U12098 (N_12098,N_11309,N_11365);
xor U12099 (N_12099,N_11965,N_11161);
and U12100 (N_12100,N_11104,N_11423);
nand U12101 (N_12101,N_11807,N_11349);
nor U12102 (N_12102,N_11220,N_11689);
nand U12103 (N_12103,N_11295,N_11132);
nor U12104 (N_12104,N_11140,N_11259);
and U12105 (N_12105,N_11415,N_11127);
and U12106 (N_12106,N_11330,N_11411);
and U12107 (N_12107,N_11382,N_11222);
and U12108 (N_12108,N_11531,N_11557);
or U12109 (N_12109,N_11952,N_11329);
nor U12110 (N_12110,N_11075,N_11871);
or U12111 (N_12111,N_11019,N_11123);
nand U12112 (N_12112,N_11824,N_11231);
or U12113 (N_12113,N_11535,N_11152);
nand U12114 (N_12114,N_11905,N_11580);
or U12115 (N_12115,N_11097,N_11168);
nor U12116 (N_12116,N_11976,N_11473);
xor U12117 (N_12117,N_11837,N_11988);
or U12118 (N_12118,N_11219,N_11202);
and U12119 (N_12119,N_11508,N_11344);
or U12120 (N_12120,N_11548,N_11897);
or U12121 (N_12121,N_11500,N_11586);
or U12122 (N_12122,N_11192,N_11900);
xor U12123 (N_12123,N_11802,N_11841);
nand U12124 (N_12124,N_11153,N_11481);
nand U12125 (N_12125,N_11521,N_11574);
and U12126 (N_12126,N_11142,N_11974);
nand U12127 (N_12127,N_11405,N_11563);
xnor U12128 (N_12128,N_11185,N_11263);
or U12129 (N_12129,N_11334,N_11336);
xor U12130 (N_12130,N_11951,N_11617);
or U12131 (N_12131,N_11795,N_11750);
and U12132 (N_12132,N_11226,N_11765);
and U12133 (N_12133,N_11959,N_11190);
or U12134 (N_12134,N_11063,N_11331);
nand U12135 (N_12135,N_11460,N_11882);
nand U12136 (N_12136,N_11513,N_11844);
nand U12137 (N_12137,N_11948,N_11560);
nor U12138 (N_12138,N_11813,N_11332);
xnor U12139 (N_12139,N_11588,N_11209);
nor U12140 (N_12140,N_11120,N_11943);
xor U12141 (N_12141,N_11568,N_11498);
nor U12142 (N_12142,N_11678,N_11591);
nor U12143 (N_12143,N_11199,N_11915);
or U12144 (N_12144,N_11698,N_11964);
or U12145 (N_12145,N_11503,N_11000);
and U12146 (N_12146,N_11221,N_11358);
and U12147 (N_12147,N_11677,N_11920);
and U12148 (N_12148,N_11863,N_11987);
xor U12149 (N_12149,N_11213,N_11624);
and U12150 (N_12150,N_11530,N_11074);
nand U12151 (N_12151,N_11319,N_11757);
and U12152 (N_12152,N_11394,N_11719);
xor U12153 (N_12153,N_11293,N_11717);
or U12154 (N_12154,N_11651,N_11676);
nor U12155 (N_12155,N_11960,N_11685);
nor U12156 (N_12156,N_11887,N_11925);
or U12157 (N_12157,N_11969,N_11725);
and U12158 (N_12158,N_11026,N_11930);
xnor U12159 (N_12159,N_11489,N_11936);
nand U12160 (N_12160,N_11679,N_11644);
or U12161 (N_12161,N_11281,N_11261);
nor U12162 (N_12162,N_11427,N_11517);
or U12163 (N_12163,N_11129,N_11524);
nand U12164 (N_12164,N_11986,N_11214);
and U12165 (N_12165,N_11047,N_11726);
xnor U12166 (N_12166,N_11040,N_11569);
nor U12167 (N_12167,N_11443,N_11504);
nor U12168 (N_12168,N_11408,N_11067);
xor U12169 (N_12169,N_11928,N_11983);
nand U12170 (N_12170,N_11593,N_11953);
xnor U12171 (N_12171,N_11552,N_11693);
or U12172 (N_12172,N_11042,N_11977);
xnor U12173 (N_12173,N_11838,N_11999);
nor U12174 (N_12174,N_11356,N_11637);
nand U12175 (N_12175,N_11572,N_11596);
or U12176 (N_12176,N_11235,N_11889);
xor U12177 (N_12177,N_11515,N_11687);
or U12178 (N_12178,N_11287,N_11324);
or U12179 (N_12179,N_11089,N_11619);
xnor U12180 (N_12180,N_11206,N_11011);
and U12181 (N_12181,N_11520,N_11949);
nor U12182 (N_12182,N_11234,N_11675);
nor U12183 (N_12183,N_11594,N_11715);
nor U12184 (N_12184,N_11227,N_11378);
nor U12185 (N_12185,N_11701,N_11610);
and U12186 (N_12186,N_11094,N_11975);
and U12187 (N_12187,N_11763,N_11122);
nor U12188 (N_12188,N_11453,N_11429);
or U12189 (N_12189,N_11193,N_11298);
nor U12190 (N_12190,N_11370,N_11156);
or U12191 (N_12191,N_11247,N_11211);
nor U12192 (N_12192,N_11923,N_11934);
xor U12193 (N_12193,N_11125,N_11032);
nor U12194 (N_12194,N_11337,N_11085);
nand U12195 (N_12195,N_11112,N_11787);
and U12196 (N_12196,N_11098,N_11095);
nand U12197 (N_12197,N_11570,N_11809);
nor U12198 (N_12198,N_11407,N_11431);
xor U12199 (N_12199,N_11171,N_11665);
and U12200 (N_12200,N_11523,N_11734);
or U12201 (N_12201,N_11631,N_11945);
and U12202 (N_12202,N_11699,N_11107);
nand U12203 (N_12203,N_11166,N_11419);
xnor U12204 (N_12204,N_11016,N_11700);
or U12205 (N_12205,N_11267,N_11046);
nand U12206 (N_12206,N_11493,N_11484);
xnor U12207 (N_12207,N_11996,N_11937);
nor U12208 (N_12208,N_11860,N_11836);
or U12209 (N_12209,N_11417,N_11422);
nand U12210 (N_12210,N_11194,N_11469);
or U12211 (N_12211,N_11006,N_11169);
xor U12212 (N_12212,N_11566,N_11933);
xnor U12213 (N_12213,N_11816,N_11522);
or U12214 (N_12214,N_11896,N_11605);
nor U12215 (N_12215,N_11187,N_11848);
nand U12216 (N_12216,N_11321,N_11806);
and U12217 (N_12217,N_11709,N_11155);
nor U12218 (N_12218,N_11590,N_11180);
nand U12219 (N_12219,N_11039,N_11845);
and U12220 (N_12220,N_11509,N_11022);
or U12221 (N_12221,N_11549,N_11705);
or U12222 (N_12222,N_11173,N_11236);
nand U12223 (N_12223,N_11462,N_11410);
xor U12224 (N_12224,N_11306,N_11065);
xnor U12225 (N_12225,N_11931,N_11359);
nor U12226 (N_12226,N_11217,N_11111);
or U12227 (N_12227,N_11589,N_11315);
or U12228 (N_12228,N_11487,N_11858);
nand U12229 (N_12229,N_11012,N_11446);
and U12230 (N_12230,N_11126,N_11627);
or U12231 (N_12231,N_11346,N_11989);
or U12232 (N_12232,N_11225,N_11029);
nor U12233 (N_12233,N_11718,N_11649);
or U12234 (N_12234,N_11659,N_11966);
and U12235 (N_12235,N_11316,N_11363);
and U12236 (N_12236,N_11366,N_11512);
or U12237 (N_12237,N_11825,N_11780);
xnor U12238 (N_12238,N_11793,N_11507);
nor U12239 (N_12239,N_11119,N_11702);
nor U12240 (N_12240,N_11543,N_11674);
nand U12241 (N_12241,N_11025,N_11274);
nand U12242 (N_12242,N_11491,N_11664);
xnor U12243 (N_12243,N_11451,N_11198);
nand U12244 (N_12244,N_11205,N_11661);
and U12245 (N_12245,N_11744,N_11308);
and U12246 (N_12246,N_11472,N_11195);
and U12247 (N_12247,N_11447,N_11265);
and U12248 (N_12248,N_11790,N_11823);
nor U12249 (N_12249,N_11929,N_11537);
xnor U12250 (N_12250,N_11303,N_11072);
and U12251 (N_12251,N_11867,N_11048);
xnor U12252 (N_12252,N_11906,N_11375);
xor U12253 (N_12253,N_11483,N_11037);
and U12254 (N_12254,N_11749,N_11536);
or U12255 (N_12255,N_11054,N_11919);
nor U12256 (N_12256,N_11950,N_11390);
xor U12257 (N_12257,N_11779,N_11448);
nand U12258 (N_12258,N_11851,N_11034);
and U12259 (N_12259,N_11847,N_11114);
and U12260 (N_12260,N_11154,N_11898);
nand U12261 (N_12261,N_11562,N_11494);
nor U12262 (N_12262,N_11559,N_11732);
xor U12263 (N_12263,N_11078,N_11635);
nor U12264 (N_12264,N_11138,N_11183);
or U12265 (N_12265,N_11781,N_11099);
nor U12266 (N_12266,N_11478,N_11538);
or U12267 (N_12267,N_11147,N_11708);
or U12268 (N_12268,N_11023,N_11284);
or U12269 (N_12269,N_11783,N_11258);
xnor U12270 (N_12270,N_11626,N_11005);
nor U12271 (N_12271,N_11377,N_11403);
and U12272 (N_12272,N_11342,N_11188);
nand U12273 (N_12273,N_11292,N_11452);
and U12274 (N_12274,N_11361,N_11418);
nand U12275 (N_12275,N_11149,N_11683);
nor U12276 (N_12276,N_11439,N_11527);
nor U12277 (N_12277,N_11020,N_11492);
xor U12278 (N_12278,N_11486,N_11990);
and U12279 (N_12279,N_11690,N_11002);
and U12280 (N_12280,N_11962,N_11395);
and U12281 (N_12281,N_11364,N_11320);
xnor U12282 (N_12282,N_11671,N_11761);
xnor U12283 (N_12283,N_11632,N_11667);
nand U12284 (N_12284,N_11852,N_11615);
or U12285 (N_12285,N_11389,N_11101);
xor U12286 (N_12286,N_11001,N_11455);
and U12287 (N_12287,N_11071,N_11421);
xnor U12288 (N_12288,N_11420,N_11868);
and U12289 (N_12289,N_11139,N_11062);
xnor U12290 (N_12290,N_11282,N_11070);
nor U12291 (N_12291,N_11317,N_11710);
nor U12292 (N_12292,N_11857,N_11087);
nor U12293 (N_12293,N_11004,N_11467);
nor U12294 (N_12294,N_11477,N_11616);
or U12295 (N_12295,N_11100,N_11033);
and U12296 (N_12296,N_11163,N_11880);
nand U12297 (N_12297,N_11461,N_11248);
xor U12298 (N_12298,N_11821,N_11669);
and U12299 (N_12299,N_11963,N_11752);
xnor U12300 (N_12300,N_11077,N_11102);
and U12301 (N_12301,N_11038,N_11831);
nor U12302 (N_12302,N_11641,N_11003);
and U12303 (N_12303,N_11241,N_11200);
xnor U12304 (N_12304,N_11944,N_11981);
nand U12305 (N_12305,N_11459,N_11926);
or U12306 (N_12306,N_11534,N_11393);
xnor U12307 (N_12307,N_11782,N_11505);
nor U12308 (N_12308,N_11172,N_11207);
and U12309 (N_12309,N_11735,N_11917);
or U12310 (N_12310,N_11724,N_11985);
or U12311 (N_12311,N_11328,N_11714);
or U12312 (N_12312,N_11666,N_11108);
nor U12313 (N_12313,N_11706,N_11729);
and U12314 (N_12314,N_11160,N_11131);
and U12315 (N_12315,N_11141,N_11820);
and U12316 (N_12316,N_11045,N_11998);
or U12317 (N_12317,N_11109,N_11565);
xnor U12318 (N_12318,N_11426,N_11068);
xnor U12319 (N_12319,N_11296,N_11412);
nor U12320 (N_12320,N_11776,N_11143);
nand U12321 (N_12321,N_11391,N_11294);
or U12322 (N_12322,N_11450,N_11577);
and U12323 (N_12323,N_11245,N_11850);
or U12324 (N_12324,N_11885,N_11178);
nand U12325 (N_12325,N_11497,N_11083);
and U12326 (N_12326,N_11081,N_11088);
nand U12327 (N_12327,N_11414,N_11133);
nand U12328 (N_12328,N_11253,N_11218);
or U12329 (N_12329,N_11396,N_11579);
or U12330 (N_12330,N_11059,N_11056);
nand U12331 (N_12331,N_11369,N_11353);
and U12332 (N_12332,N_11647,N_11191);
or U12333 (N_12333,N_11252,N_11629);
or U12334 (N_12334,N_11480,N_11430);
xnor U12335 (N_12335,N_11017,N_11351);
xor U12336 (N_12336,N_11290,N_11597);
and U12337 (N_12337,N_11266,N_11404);
nand U12338 (N_12338,N_11712,N_11803);
or U12339 (N_12339,N_11839,N_11468);
xnor U12340 (N_12340,N_11982,N_11340);
nand U12341 (N_12341,N_11886,N_11592);
or U12342 (N_12342,N_11814,N_11682);
xnor U12343 (N_12343,N_11595,N_11630);
and U12344 (N_12344,N_11130,N_11797);
and U12345 (N_12345,N_11908,N_11643);
nor U12346 (N_12346,N_11942,N_11875);
nand U12347 (N_12347,N_11546,N_11972);
nor U12348 (N_12348,N_11028,N_11788);
xnor U12349 (N_12349,N_11397,N_11633);
xnor U12350 (N_12350,N_11738,N_11043);
nand U12351 (N_12351,N_11158,N_11518);
nand U12352 (N_12352,N_11313,N_11778);
nand U12353 (N_12353,N_11145,N_11533);
xnor U12354 (N_12354,N_11648,N_11694);
xor U12355 (N_12355,N_11556,N_11737);
nand U12356 (N_12356,N_11402,N_11115);
and U12357 (N_12357,N_11939,N_11888);
xor U12358 (N_12358,N_11251,N_11189);
nor U12359 (N_12359,N_11053,N_11118);
and U12360 (N_12360,N_11849,N_11381);
nand U12361 (N_12361,N_11442,N_11269);
nand U12362 (N_12362,N_11184,N_11283);
or U12363 (N_12363,N_11606,N_11049);
or U12364 (N_12364,N_11413,N_11638);
nor U12365 (N_12365,N_11449,N_11621);
or U12366 (N_12366,N_11036,N_11876);
xnor U12367 (N_12367,N_11542,N_11181);
and U12368 (N_12368,N_11587,N_11555);
and U12369 (N_12369,N_11691,N_11177);
nor U12370 (N_12370,N_11623,N_11770);
nor U12371 (N_12371,N_11525,N_11571);
and U12372 (N_12372,N_11519,N_11827);
or U12373 (N_12373,N_11646,N_11731);
nor U12374 (N_12374,N_11399,N_11254);
or U12375 (N_12375,N_11540,N_11739);
or U12376 (N_12376,N_11657,N_11400);
nand U12377 (N_12377,N_11203,N_11246);
nand U12378 (N_12378,N_11310,N_11136);
or U12379 (N_12379,N_11970,N_11090);
or U12380 (N_12380,N_11968,N_11333);
nor U12381 (N_12381,N_11585,N_11179);
or U12382 (N_12382,N_11436,N_11918);
xnor U12383 (N_12383,N_11212,N_11474);
nand U12384 (N_12384,N_11278,N_11681);
or U12385 (N_12385,N_11233,N_11456);
and U12386 (N_12386,N_11688,N_11470);
and U12387 (N_12387,N_11553,N_11326);
or U12388 (N_12388,N_11645,N_11240);
and U12389 (N_12389,N_11743,N_11300);
or U12390 (N_12390,N_11881,N_11066);
nor U12391 (N_12391,N_11438,N_11237);
nor U12392 (N_12392,N_11499,N_11092);
nand U12393 (N_12393,N_11684,N_11561);
xnor U12394 (N_12394,N_11544,N_11031);
or U12395 (N_12395,N_11164,N_11854);
xor U12396 (N_12396,N_11668,N_11958);
xnor U12397 (N_12397,N_11204,N_11994);
nor U12398 (N_12398,N_11371,N_11891);
xnor U12399 (N_12399,N_11658,N_11834);
nand U12400 (N_12400,N_11941,N_11804);
xnor U12401 (N_12401,N_11277,N_11869);
nand U12402 (N_12402,N_11894,N_11828);
xnor U12403 (N_12403,N_11105,N_11554);
and U12404 (N_12404,N_11914,N_11791);
or U12405 (N_12405,N_11760,N_11216);
nand U12406 (N_12406,N_11884,N_11013);
nor U12407 (N_12407,N_11086,N_11946);
nor U12408 (N_12408,N_11256,N_11727);
or U12409 (N_12409,N_11611,N_11475);
nand U12410 (N_12410,N_11634,N_11895);
and U12411 (N_12411,N_11742,N_11769);
nand U12412 (N_12412,N_11276,N_11069);
nor U12413 (N_12413,N_11113,N_11991);
xnor U12414 (N_12414,N_11479,N_11613);
or U12415 (N_12415,N_11015,N_11746);
nor U12416 (N_12416,N_11304,N_11777);
nor U12417 (N_12417,N_11575,N_11457);
nand U12418 (N_12418,N_11182,N_11260);
xnor U12419 (N_12419,N_11747,N_11335);
nor U12420 (N_12420,N_11064,N_11736);
or U12421 (N_12421,N_11921,N_11817);
nor U12422 (N_12422,N_11878,N_11927);
nand U12423 (N_12423,N_11789,N_11912);
nand U12424 (N_12424,N_11843,N_11607);
nor U12425 (N_12425,N_11545,N_11345);
nand U12426 (N_12426,N_11466,N_11367);
or U12427 (N_12427,N_11756,N_11796);
nor U12428 (N_12428,N_11911,N_11079);
xor U12429 (N_12429,N_11957,N_11435);
nor U12430 (N_12430,N_11997,N_11398);
xnor U12431 (N_12431,N_11339,N_11883);
xnor U12432 (N_12432,N_11322,N_11992);
nand U12433 (N_12433,N_11916,N_11703);
and U12434 (N_12434,N_11670,N_11229);
xnor U12435 (N_12435,N_11428,N_11864);
nand U12436 (N_12436,N_11082,N_11060);
and U12437 (N_12437,N_11264,N_11663);
and U12438 (N_12438,N_11978,N_11603);
and U12439 (N_12439,N_11116,N_11357);
or U12440 (N_12440,N_11307,N_11230);
and U12441 (N_12441,N_11656,N_11801);
xor U12442 (N_12442,N_11892,N_11239);
xor U12443 (N_12443,N_11955,N_11270);
nor U12444 (N_12444,N_11372,N_11463);
nand U12445 (N_12445,N_11913,N_11856);
nor U12446 (N_12446,N_11215,N_11584);
or U12447 (N_12447,N_11151,N_11618);
nand U12448 (N_12448,N_11855,N_11380);
xor U12449 (N_12449,N_11024,N_11822);
nor U12450 (N_12450,N_11932,N_11800);
nand U12451 (N_12451,N_11510,N_11343);
xor U12452 (N_12452,N_11165,N_11600);
nor U12453 (N_12453,N_11861,N_11818);
nand U12454 (N_12454,N_11445,N_11091);
nand U12455 (N_12455,N_11551,N_11444);
or U12456 (N_12456,N_11862,N_11622);
nor U12457 (N_12457,N_11210,N_11440);
nor U12458 (N_12458,N_11223,N_11654);
nor U12459 (N_12459,N_11578,N_11826);
and U12460 (N_12460,N_11673,N_11238);
and U12461 (N_12461,N_11495,N_11416);
and U12462 (N_12462,N_11971,N_11250);
nand U12463 (N_12463,N_11753,N_11302);
nor U12464 (N_12464,N_11660,N_11044);
and U12465 (N_12465,N_11352,N_11961);
nor U12466 (N_12466,N_11775,N_11567);
or U12467 (N_12467,N_11425,N_11347);
nor U12468 (N_12468,N_11159,N_11686);
or U12469 (N_12469,N_11379,N_11388);
and U12470 (N_12470,N_11899,N_11373);
or U12471 (N_12471,N_11255,N_11808);
and U12472 (N_12472,N_11740,N_11901);
nand U12473 (N_12473,N_11262,N_11819);
or U12474 (N_12474,N_11110,N_11853);
nor U12475 (N_12475,N_11755,N_11614);
nor U12476 (N_12476,N_11196,N_11279);
or U12477 (N_12477,N_11007,N_11741);
and U12478 (N_12478,N_11877,N_11745);
xor U12479 (N_12479,N_11124,N_11754);
nand U12480 (N_12480,N_11008,N_11268);
or U12481 (N_12481,N_11805,N_11244);
nand U12482 (N_12482,N_11170,N_11539);
xnor U12483 (N_12483,N_11228,N_11582);
or U12484 (N_12484,N_11967,N_11271);
or U12485 (N_12485,N_11014,N_11835);
xor U12486 (N_12486,N_11640,N_11030);
or U12487 (N_12487,N_11680,N_11815);
nand U12488 (N_12488,N_11424,N_11842);
xnor U12489 (N_12489,N_11144,N_11832);
xor U12490 (N_12490,N_11697,N_11465);
nor U12491 (N_12491,N_11297,N_11599);
nor U12492 (N_12492,N_11846,N_11980);
and U12493 (N_12493,N_11833,N_11956);
or U12494 (N_12494,N_11009,N_11314);
xnor U12495 (N_12495,N_11437,N_11768);
or U12496 (N_12496,N_11758,N_11434);
nor U12497 (N_12497,N_11873,N_11652);
xnor U12498 (N_12498,N_11979,N_11514);
or U12499 (N_12499,N_11909,N_11106);
nor U12500 (N_12500,N_11966,N_11200);
or U12501 (N_12501,N_11237,N_11888);
and U12502 (N_12502,N_11661,N_11073);
nor U12503 (N_12503,N_11953,N_11305);
nand U12504 (N_12504,N_11226,N_11104);
nor U12505 (N_12505,N_11803,N_11939);
and U12506 (N_12506,N_11594,N_11665);
nand U12507 (N_12507,N_11864,N_11566);
or U12508 (N_12508,N_11242,N_11504);
nor U12509 (N_12509,N_11182,N_11842);
or U12510 (N_12510,N_11727,N_11566);
xnor U12511 (N_12511,N_11578,N_11119);
and U12512 (N_12512,N_11849,N_11860);
and U12513 (N_12513,N_11893,N_11693);
xor U12514 (N_12514,N_11572,N_11617);
nand U12515 (N_12515,N_11240,N_11043);
nand U12516 (N_12516,N_11253,N_11689);
nor U12517 (N_12517,N_11682,N_11201);
xnor U12518 (N_12518,N_11890,N_11426);
xnor U12519 (N_12519,N_11726,N_11031);
or U12520 (N_12520,N_11788,N_11196);
xor U12521 (N_12521,N_11387,N_11686);
and U12522 (N_12522,N_11345,N_11855);
or U12523 (N_12523,N_11356,N_11475);
and U12524 (N_12524,N_11275,N_11183);
nand U12525 (N_12525,N_11718,N_11256);
nor U12526 (N_12526,N_11352,N_11815);
or U12527 (N_12527,N_11860,N_11616);
xor U12528 (N_12528,N_11550,N_11395);
and U12529 (N_12529,N_11682,N_11545);
xor U12530 (N_12530,N_11271,N_11956);
xnor U12531 (N_12531,N_11124,N_11483);
nor U12532 (N_12532,N_11932,N_11305);
xor U12533 (N_12533,N_11811,N_11890);
xor U12534 (N_12534,N_11954,N_11914);
nand U12535 (N_12535,N_11781,N_11308);
and U12536 (N_12536,N_11470,N_11716);
or U12537 (N_12537,N_11351,N_11711);
nand U12538 (N_12538,N_11775,N_11703);
or U12539 (N_12539,N_11020,N_11889);
xor U12540 (N_12540,N_11579,N_11668);
xnor U12541 (N_12541,N_11547,N_11701);
and U12542 (N_12542,N_11625,N_11182);
or U12543 (N_12543,N_11991,N_11155);
and U12544 (N_12544,N_11566,N_11601);
xor U12545 (N_12545,N_11614,N_11573);
or U12546 (N_12546,N_11180,N_11533);
and U12547 (N_12547,N_11909,N_11649);
xor U12548 (N_12548,N_11435,N_11405);
or U12549 (N_12549,N_11797,N_11127);
and U12550 (N_12550,N_11410,N_11894);
xor U12551 (N_12551,N_11923,N_11691);
nand U12552 (N_12552,N_11884,N_11428);
nand U12553 (N_12553,N_11758,N_11739);
or U12554 (N_12554,N_11758,N_11460);
xnor U12555 (N_12555,N_11535,N_11194);
nor U12556 (N_12556,N_11147,N_11383);
nor U12557 (N_12557,N_11901,N_11202);
or U12558 (N_12558,N_11998,N_11088);
or U12559 (N_12559,N_11049,N_11398);
nor U12560 (N_12560,N_11963,N_11182);
xor U12561 (N_12561,N_11257,N_11243);
xor U12562 (N_12562,N_11307,N_11998);
nand U12563 (N_12563,N_11205,N_11209);
xnor U12564 (N_12564,N_11702,N_11069);
nand U12565 (N_12565,N_11987,N_11377);
xor U12566 (N_12566,N_11840,N_11015);
or U12567 (N_12567,N_11993,N_11096);
and U12568 (N_12568,N_11654,N_11322);
nor U12569 (N_12569,N_11860,N_11962);
and U12570 (N_12570,N_11778,N_11141);
xor U12571 (N_12571,N_11892,N_11033);
nand U12572 (N_12572,N_11192,N_11277);
and U12573 (N_12573,N_11711,N_11344);
xnor U12574 (N_12574,N_11497,N_11727);
nor U12575 (N_12575,N_11502,N_11380);
and U12576 (N_12576,N_11612,N_11477);
nor U12577 (N_12577,N_11853,N_11776);
nor U12578 (N_12578,N_11560,N_11203);
xnor U12579 (N_12579,N_11537,N_11923);
xnor U12580 (N_12580,N_11741,N_11084);
and U12581 (N_12581,N_11895,N_11089);
and U12582 (N_12582,N_11458,N_11641);
xor U12583 (N_12583,N_11052,N_11948);
and U12584 (N_12584,N_11584,N_11175);
and U12585 (N_12585,N_11045,N_11295);
and U12586 (N_12586,N_11659,N_11511);
xor U12587 (N_12587,N_11577,N_11127);
or U12588 (N_12588,N_11039,N_11697);
nand U12589 (N_12589,N_11434,N_11929);
xnor U12590 (N_12590,N_11400,N_11268);
nor U12591 (N_12591,N_11051,N_11101);
xor U12592 (N_12592,N_11608,N_11505);
xor U12593 (N_12593,N_11373,N_11207);
nand U12594 (N_12594,N_11105,N_11948);
and U12595 (N_12595,N_11171,N_11468);
nor U12596 (N_12596,N_11992,N_11110);
xnor U12597 (N_12597,N_11829,N_11284);
and U12598 (N_12598,N_11478,N_11612);
or U12599 (N_12599,N_11121,N_11697);
or U12600 (N_12600,N_11291,N_11976);
xor U12601 (N_12601,N_11909,N_11112);
nand U12602 (N_12602,N_11012,N_11695);
or U12603 (N_12603,N_11600,N_11166);
xnor U12604 (N_12604,N_11792,N_11121);
nor U12605 (N_12605,N_11699,N_11047);
xnor U12606 (N_12606,N_11290,N_11869);
nand U12607 (N_12607,N_11261,N_11170);
and U12608 (N_12608,N_11034,N_11867);
and U12609 (N_12609,N_11781,N_11927);
xor U12610 (N_12610,N_11253,N_11958);
nand U12611 (N_12611,N_11733,N_11225);
nand U12612 (N_12612,N_11929,N_11141);
or U12613 (N_12613,N_11257,N_11713);
nor U12614 (N_12614,N_11945,N_11152);
nor U12615 (N_12615,N_11854,N_11397);
nand U12616 (N_12616,N_11865,N_11435);
xor U12617 (N_12617,N_11663,N_11134);
or U12618 (N_12618,N_11039,N_11024);
and U12619 (N_12619,N_11916,N_11631);
xnor U12620 (N_12620,N_11903,N_11613);
nor U12621 (N_12621,N_11251,N_11426);
or U12622 (N_12622,N_11053,N_11319);
and U12623 (N_12623,N_11007,N_11713);
or U12624 (N_12624,N_11922,N_11107);
xor U12625 (N_12625,N_11430,N_11832);
and U12626 (N_12626,N_11122,N_11927);
nor U12627 (N_12627,N_11916,N_11230);
or U12628 (N_12628,N_11787,N_11371);
nor U12629 (N_12629,N_11263,N_11190);
or U12630 (N_12630,N_11267,N_11655);
or U12631 (N_12631,N_11732,N_11677);
xnor U12632 (N_12632,N_11474,N_11105);
xor U12633 (N_12633,N_11519,N_11008);
nor U12634 (N_12634,N_11389,N_11930);
and U12635 (N_12635,N_11386,N_11775);
or U12636 (N_12636,N_11879,N_11611);
and U12637 (N_12637,N_11777,N_11471);
nor U12638 (N_12638,N_11320,N_11491);
nand U12639 (N_12639,N_11362,N_11011);
nand U12640 (N_12640,N_11271,N_11517);
or U12641 (N_12641,N_11928,N_11847);
nor U12642 (N_12642,N_11785,N_11583);
nand U12643 (N_12643,N_11417,N_11766);
and U12644 (N_12644,N_11079,N_11786);
or U12645 (N_12645,N_11405,N_11932);
or U12646 (N_12646,N_11020,N_11542);
nand U12647 (N_12647,N_11833,N_11423);
nor U12648 (N_12648,N_11754,N_11563);
or U12649 (N_12649,N_11479,N_11541);
xor U12650 (N_12650,N_11306,N_11710);
and U12651 (N_12651,N_11953,N_11629);
xnor U12652 (N_12652,N_11825,N_11540);
and U12653 (N_12653,N_11384,N_11908);
xnor U12654 (N_12654,N_11701,N_11511);
nand U12655 (N_12655,N_11421,N_11843);
xor U12656 (N_12656,N_11885,N_11344);
and U12657 (N_12657,N_11628,N_11967);
nand U12658 (N_12658,N_11716,N_11592);
xnor U12659 (N_12659,N_11634,N_11236);
and U12660 (N_12660,N_11383,N_11533);
or U12661 (N_12661,N_11528,N_11827);
and U12662 (N_12662,N_11814,N_11711);
or U12663 (N_12663,N_11432,N_11492);
nand U12664 (N_12664,N_11271,N_11438);
nor U12665 (N_12665,N_11461,N_11311);
or U12666 (N_12666,N_11299,N_11296);
nor U12667 (N_12667,N_11798,N_11449);
xor U12668 (N_12668,N_11911,N_11620);
nand U12669 (N_12669,N_11091,N_11398);
nand U12670 (N_12670,N_11365,N_11611);
xor U12671 (N_12671,N_11082,N_11462);
or U12672 (N_12672,N_11203,N_11578);
nand U12673 (N_12673,N_11054,N_11359);
or U12674 (N_12674,N_11506,N_11090);
and U12675 (N_12675,N_11422,N_11501);
nor U12676 (N_12676,N_11284,N_11220);
or U12677 (N_12677,N_11397,N_11555);
nor U12678 (N_12678,N_11616,N_11695);
or U12679 (N_12679,N_11320,N_11600);
nand U12680 (N_12680,N_11352,N_11194);
xnor U12681 (N_12681,N_11241,N_11778);
nor U12682 (N_12682,N_11417,N_11611);
nand U12683 (N_12683,N_11099,N_11867);
or U12684 (N_12684,N_11178,N_11700);
and U12685 (N_12685,N_11520,N_11616);
nand U12686 (N_12686,N_11273,N_11171);
or U12687 (N_12687,N_11402,N_11063);
xnor U12688 (N_12688,N_11745,N_11347);
and U12689 (N_12689,N_11403,N_11193);
and U12690 (N_12690,N_11541,N_11768);
nand U12691 (N_12691,N_11862,N_11833);
and U12692 (N_12692,N_11173,N_11563);
xnor U12693 (N_12693,N_11359,N_11977);
or U12694 (N_12694,N_11535,N_11569);
xnor U12695 (N_12695,N_11940,N_11981);
nor U12696 (N_12696,N_11355,N_11914);
nor U12697 (N_12697,N_11349,N_11511);
and U12698 (N_12698,N_11270,N_11070);
nand U12699 (N_12699,N_11381,N_11341);
xor U12700 (N_12700,N_11929,N_11173);
nor U12701 (N_12701,N_11526,N_11660);
nor U12702 (N_12702,N_11890,N_11241);
nand U12703 (N_12703,N_11819,N_11336);
xor U12704 (N_12704,N_11005,N_11492);
and U12705 (N_12705,N_11585,N_11353);
nand U12706 (N_12706,N_11741,N_11643);
nor U12707 (N_12707,N_11767,N_11362);
xor U12708 (N_12708,N_11237,N_11060);
or U12709 (N_12709,N_11040,N_11975);
or U12710 (N_12710,N_11982,N_11129);
xnor U12711 (N_12711,N_11667,N_11096);
xnor U12712 (N_12712,N_11259,N_11890);
xor U12713 (N_12713,N_11929,N_11579);
nand U12714 (N_12714,N_11230,N_11463);
or U12715 (N_12715,N_11426,N_11339);
nand U12716 (N_12716,N_11357,N_11630);
nand U12717 (N_12717,N_11858,N_11579);
and U12718 (N_12718,N_11656,N_11318);
xnor U12719 (N_12719,N_11814,N_11601);
nand U12720 (N_12720,N_11379,N_11635);
and U12721 (N_12721,N_11522,N_11212);
and U12722 (N_12722,N_11384,N_11581);
xnor U12723 (N_12723,N_11303,N_11648);
nor U12724 (N_12724,N_11949,N_11663);
nor U12725 (N_12725,N_11114,N_11830);
and U12726 (N_12726,N_11138,N_11371);
nor U12727 (N_12727,N_11591,N_11847);
or U12728 (N_12728,N_11277,N_11805);
and U12729 (N_12729,N_11819,N_11408);
and U12730 (N_12730,N_11236,N_11705);
nand U12731 (N_12731,N_11662,N_11142);
or U12732 (N_12732,N_11276,N_11006);
nand U12733 (N_12733,N_11686,N_11295);
or U12734 (N_12734,N_11894,N_11444);
nor U12735 (N_12735,N_11108,N_11559);
nand U12736 (N_12736,N_11645,N_11601);
and U12737 (N_12737,N_11253,N_11939);
and U12738 (N_12738,N_11404,N_11214);
or U12739 (N_12739,N_11818,N_11799);
nand U12740 (N_12740,N_11961,N_11093);
and U12741 (N_12741,N_11898,N_11959);
xnor U12742 (N_12742,N_11421,N_11670);
or U12743 (N_12743,N_11530,N_11887);
and U12744 (N_12744,N_11015,N_11907);
nand U12745 (N_12745,N_11185,N_11008);
nor U12746 (N_12746,N_11438,N_11933);
xor U12747 (N_12747,N_11151,N_11299);
nand U12748 (N_12748,N_11483,N_11923);
nand U12749 (N_12749,N_11583,N_11804);
nor U12750 (N_12750,N_11789,N_11507);
nor U12751 (N_12751,N_11013,N_11574);
or U12752 (N_12752,N_11091,N_11582);
xor U12753 (N_12753,N_11602,N_11482);
or U12754 (N_12754,N_11269,N_11433);
nor U12755 (N_12755,N_11568,N_11910);
or U12756 (N_12756,N_11587,N_11677);
nor U12757 (N_12757,N_11690,N_11006);
nor U12758 (N_12758,N_11896,N_11627);
nor U12759 (N_12759,N_11914,N_11315);
or U12760 (N_12760,N_11465,N_11764);
and U12761 (N_12761,N_11117,N_11151);
xnor U12762 (N_12762,N_11688,N_11405);
nand U12763 (N_12763,N_11597,N_11232);
nand U12764 (N_12764,N_11212,N_11031);
nand U12765 (N_12765,N_11356,N_11903);
and U12766 (N_12766,N_11965,N_11760);
and U12767 (N_12767,N_11304,N_11749);
nor U12768 (N_12768,N_11026,N_11456);
or U12769 (N_12769,N_11175,N_11097);
and U12770 (N_12770,N_11520,N_11672);
xnor U12771 (N_12771,N_11779,N_11096);
or U12772 (N_12772,N_11162,N_11440);
or U12773 (N_12773,N_11250,N_11658);
nand U12774 (N_12774,N_11213,N_11957);
nor U12775 (N_12775,N_11352,N_11904);
and U12776 (N_12776,N_11911,N_11123);
or U12777 (N_12777,N_11783,N_11497);
and U12778 (N_12778,N_11961,N_11553);
xnor U12779 (N_12779,N_11897,N_11449);
and U12780 (N_12780,N_11128,N_11860);
xnor U12781 (N_12781,N_11488,N_11421);
xnor U12782 (N_12782,N_11604,N_11784);
and U12783 (N_12783,N_11130,N_11276);
nor U12784 (N_12784,N_11019,N_11455);
nand U12785 (N_12785,N_11934,N_11759);
or U12786 (N_12786,N_11592,N_11165);
nand U12787 (N_12787,N_11288,N_11520);
xnor U12788 (N_12788,N_11424,N_11931);
xor U12789 (N_12789,N_11428,N_11677);
and U12790 (N_12790,N_11334,N_11380);
nor U12791 (N_12791,N_11179,N_11644);
xnor U12792 (N_12792,N_11872,N_11544);
nor U12793 (N_12793,N_11744,N_11866);
and U12794 (N_12794,N_11898,N_11253);
nand U12795 (N_12795,N_11539,N_11090);
or U12796 (N_12796,N_11272,N_11736);
or U12797 (N_12797,N_11400,N_11545);
nand U12798 (N_12798,N_11658,N_11335);
or U12799 (N_12799,N_11326,N_11595);
nor U12800 (N_12800,N_11274,N_11234);
nor U12801 (N_12801,N_11204,N_11178);
xor U12802 (N_12802,N_11617,N_11389);
and U12803 (N_12803,N_11874,N_11861);
or U12804 (N_12804,N_11736,N_11697);
and U12805 (N_12805,N_11999,N_11868);
xnor U12806 (N_12806,N_11132,N_11211);
nor U12807 (N_12807,N_11322,N_11558);
nand U12808 (N_12808,N_11049,N_11402);
nand U12809 (N_12809,N_11715,N_11013);
nand U12810 (N_12810,N_11556,N_11107);
nand U12811 (N_12811,N_11886,N_11394);
and U12812 (N_12812,N_11544,N_11182);
nand U12813 (N_12813,N_11154,N_11599);
or U12814 (N_12814,N_11263,N_11810);
and U12815 (N_12815,N_11203,N_11752);
and U12816 (N_12816,N_11478,N_11766);
nand U12817 (N_12817,N_11393,N_11978);
and U12818 (N_12818,N_11657,N_11943);
nor U12819 (N_12819,N_11630,N_11258);
nand U12820 (N_12820,N_11306,N_11828);
nor U12821 (N_12821,N_11794,N_11955);
or U12822 (N_12822,N_11255,N_11793);
nand U12823 (N_12823,N_11721,N_11110);
nand U12824 (N_12824,N_11541,N_11401);
nand U12825 (N_12825,N_11035,N_11587);
and U12826 (N_12826,N_11094,N_11105);
nand U12827 (N_12827,N_11257,N_11428);
and U12828 (N_12828,N_11328,N_11298);
nand U12829 (N_12829,N_11343,N_11625);
nor U12830 (N_12830,N_11031,N_11785);
or U12831 (N_12831,N_11662,N_11678);
or U12832 (N_12832,N_11282,N_11431);
nor U12833 (N_12833,N_11582,N_11547);
nand U12834 (N_12834,N_11319,N_11129);
and U12835 (N_12835,N_11487,N_11550);
or U12836 (N_12836,N_11099,N_11165);
or U12837 (N_12837,N_11788,N_11558);
nor U12838 (N_12838,N_11217,N_11694);
xor U12839 (N_12839,N_11264,N_11516);
or U12840 (N_12840,N_11430,N_11555);
nand U12841 (N_12841,N_11463,N_11944);
nand U12842 (N_12842,N_11949,N_11322);
xnor U12843 (N_12843,N_11298,N_11946);
and U12844 (N_12844,N_11523,N_11770);
nor U12845 (N_12845,N_11898,N_11303);
nor U12846 (N_12846,N_11199,N_11475);
nand U12847 (N_12847,N_11481,N_11532);
xor U12848 (N_12848,N_11519,N_11997);
nand U12849 (N_12849,N_11783,N_11335);
or U12850 (N_12850,N_11249,N_11951);
nand U12851 (N_12851,N_11243,N_11863);
or U12852 (N_12852,N_11488,N_11412);
xnor U12853 (N_12853,N_11314,N_11819);
or U12854 (N_12854,N_11523,N_11260);
and U12855 (N_12855,N_11579,N_11684);
or U12856 (N_12856,N_11837,N_11054);
nand U12857 (N_12857,N_11930,N_11282);
xor U12858 (N_12858,N_11107,N_11713);
and U12859 (N_12859,N_11023,N_11956);
nor U12860 (N_12860,N_11636,N_11142);
and U12861 (N_12861,N_11797,N_11213);
or U12862 (N_12862,N_11973,N_11529);
xor U12863 (N_12863,N_11398,N_11466);
and U12864 (N_12864,N_11272,N_11780);
nor U12865 (N_12865,N_11427,N_11348);
nand U12866 (N_12866,N_11006,N_11823);
nor U12867 (N_12867,N_11943,N_11438);
nor U12868 (N_12868,N_11285,N_11186);
or U12869 (N_12869,N_11955,N_11186);
or U12870 (N_12870,N_11800,N_11093);
and U12871 (N_12871,N_11659,N_11723);
xor U12872 (N_12872,N_11309,N_11968);
xor U12873 (N_12873,N_11168,N_11171);
nor U12874 (N_12874,N_11221,N_11144);
and U12875 (N_12875,N_11832,N_11976);
nor U12876 (N_12876,N_11611,N_11749);
or U12877 (N_12877,N_11676,N_11639);
nor U12878 (N_12878,N_11471,N_11457);
xor U12879 (N_12879,N_11540,N_11710);
nand U12880 (N_12880,N_11607,N_11074);
nor U12881 (N_12881,N_11792,N_11702);
nor U12882 (N_12882,N_11603,N_11159);
nand U12883 (N_12883,N_11029,N_11156);
or U12884 (N_12884,N_11673,N_11979);
nand U12885 (N_12885,N_11331,N_11422);
and U12886 (N_12886,N_11204,N_11082);
xnor U12887 (N_12887,N_11721,N_11036);
or U12888 (N_12888,N_11714,N_11944);
nor U12889 (N_12889,N_11134,N_11623);
and U12890 (N_12890,N_11513,N_11239);
and U12891 (N_12891,N_11044,N_11279);
xor U12892 (N_12892,N_11243,N_11288);
nand U12893 (N_12893,N_11655,N_11648);
xnor U12894 (N_12894,N_11721,N_11506);
nand U12895 (N_12895,N_11111,N_11766);
and U12896 (N_12896,N_11202,N_11248);
or U12897 (N_12897,N_11763,N_11232);
and U12898 (N_12898,N_11805,N_11315);
nand U12899 (N_12899,N_11660,N_11822);
or U12900 (N_12900,N_11870,N_11346);
and U12901 (N_12901,N_11435,N_11093);
nor U12902 (N_12902,N_11954,N_11982);
xnor U12903 (N_12903,N_11176,N_11418);
nand U12904 (N_12904,N_11529,N_11430);
nor U12905 (N_12905,N_11252,N_11663);
and U12906 (N_12906,N_11386,N_11615);
xnor U12907 (N_12907,N_11262,N_11162);
and U12908 (N_12908,N_11623,N_11189);
and U12909 (N_12909,N_11984,N_11464);
nand U12910 (N_12910,N_11755,N_11063);
nand U12911 (N_12911,N_11986,N_11257);
nor U12912 (N_12912,N_11776,N_11156);
or U12913 (N_12913,N_11790,N_11452);
nor U12914 (N_12914,N_11153,N_11625);
nor U12915 (N_12915,N_11347,N_11957);
and U12916 (N_12916,N_11737,N_11152);
nor U12917 (N_12917,N_11505,N_11076);
or U12918 (N_12918,N_11031,N_11800);
nor U12919 (N_12919,N_11830,N_11711);
xnor U12920 (N_12920,N_11339,N_11856);
xor U12921 (N_12921,N_11959,N_11334);
nand U12922 (N_12922,N_11556,N_11190);
or U12923 (N_12923,N_11926,N_11191);
or U12924 (N_12924,N_11823,N_11422);
nor U12925 (N_12925,N_11951,N_11065);
and U12926 (N_12926,N_11636,N_11525);
nand U12927 (N_12927,N_11267,N_11167);
and U12928 (N_12928,N_11279,N_11013);
and U12929 (N_12929,N_11821,N_11837);
xnor U12930 (N_12930,N_11987,N_11920);
or U12931 (N_12931,N_11989,N_11193);
nand U12932 (N_12932,N_11497,N_11395);
nor U12933 (N_12933,N_11167,N_11905);
nand U12934 (N_12934,N_11141,N_11931);
nor U12935 (N_12935,N_11215,N_11800);
xnor U12936 (N_12936,N_11024,N_11980);
and U12937 (N_12937,N_11950,N_11520);
and U12938 (N_12938,N_11400,N_11471);
nor U12939 (N_12939,N_11498,N_11260);
or U12940 (N_12940,N_11131,N_11127);
xor U12941 (N_12941,N_11060,N_11416);
xor U12942 (N_12942,N_11330,N_11219);
xnor U12943 (N_12943,N_11993,N_11919);
nand U12944 (N_12944,N_11220,N_11305);
nand U12945 (N_12945,N_11081,N_11862);
nand U12946 (N_12946,N_11297,N_11357);
nand U12947 (N_12947,N_11373,N_11404);
nand U12948 (N_12948,N_11047,N_11692);
nand U12949 (N_12949,N_11992,N_11482);
nor U12950 (N_12950,N_11188,N_11532);
nor U12951 (N_12951,N_11370,N_11914);
and U12952 (N_12952,N_11493,N_11167);
xor U12953 (N_12953,N_11552,N_11767);
or U12954 (N_12954,N_11277,N_11517);
xor U12955 (N_12955,N_11046,N_11463);
and U12956 (N_12956,N_11387,N_11441);
nand U12957 (N_12957,N_11264,N_11407);
xnor U12958 (N_12958,N_11706,N_11852);
and U12959 (N_12959,N_11112,N_11542);
or U12960 (N_12960,N_11855,N_11518);
or U12961 (N_12961,N_11758,N_11005);
or U12962 (N_12962,N_11904,N_11823);
nor U12963 (N_12963,N_11808,N_11036);
xor U12964 (N_12964,N_11711,N_11781);
nor U12965 (N_12965,N_11842,N_11323);
or U12966 (N_12966,N_11950,N_11572);
nor U12967 (N_12967,N_11381,N_11160);
xor U12968 (N_12968,N_11456,N_11229);
xnor U12969 (N_12969,N_11257,N_11963);
xnor U12970 (N_12970,N_11136,N_11026);
xnor U12971 (N_12971,N_11057,N_11870);
nand U12972 (N_12972,N_11258,N_11217);
nand U12973 (N_12973,N_11276,N_11224);
nand U12974 (N_12974,N_11922,N_11355);
and U12975 (N_12975,N_11820,N_11494);
xnor U12976 (N_12976,N_11821,N_11960);
xor U12977 (N_12977,N_11994,N_11547);
nor U12978 (N_12978,N_11206,N_11180);
and U12979 (N_12979,N_11624,N_11882);
xnor U12980 (N_12980,N_11538,N_11609);
or U12981 (N_12981,N_11292,N_11192);
and U12982 (N_12982,N_11717,N_11426);
or U12983 (N_12983,N_11354,N_11866);
and U12984 (N_12984,N_11083,N_11002);
and U12985 (N_12985,N_11640,N_11083);
nor U12986 (N_12986,N_11313,N_11884);
nor U12987 (N_12987,N_11160,N_11073);
xnor U12988 (N_12988,N_11404,N_11038);
nand U12989 (N_12989,N_11179,N_11796);
xor U12990 (N_12990,N_11986,N_11081);
and U12991 (N_12991,N_11900,N_11559);
nor U12992 (N_12992,N_11331,N_11280);
or U12993 (N_12993,N_11034,N_11279);
nor U12994 (N_12994,N_11657,N_11418);
nand U12995 (N_12995,N_11466,N_11567);
xor U12996 (N_12996,N_11697,N_11543);
xnor U12997 (N_12997,N_11886,N_11331);
and U12998 (N_12998,N_11717,N_11896);
nand U12999 (N_12999,N_11990,N_11655);
and U13000 (N_13000,N_12379,N_12690);
xor U13001 (N_13001,N_12122,N_12175);
and U13002 (N_13002,N_12244,N_12697);
nand U13003 (N_13003,N_12142,N_12202);
nor U13004 (N_13004,N_12651,N_12861);
nor U13005 (N_13005,N_12024,N_12281);
nand U13006 (N_13006,N_12787,N_12738);
xnor U13007 (N_13007,N_12101,N_12856);
or U13008 (N_13008,N_12286,N_12884);
and U13009 (N_13009,N_12640,N_12868);
xor U13010 (N_13010,N_12305,N_12616);
and U13011 (N_13011,N_12888,N_12415);
or U13012 (N_13012,N_12693,N_12176);
nand U13013 (N_13013,N_12980,N_12784);
and U13014 (N_13014,N_12205,N_12493);
nor U13015 (N_13015,N_12181,N_12094);
and U13016 (N_13016,N_12902,N_12439);
nor U13017 (N_13017,N_12885,N_12847);
nand U13018 (N_13018,N_12157,N_12354);
or U13019 (N_13019,N_12214,N_12832);
xor U13020 (N_13020,N_12546,N_12645);
nand U13021 (N_13021,N_12454,N_12704);
nand U13022 (N_13022,N_12227,N_12150);
nand U13023 (N_13023,N_12029,N_12539);
xnor U13024 (N_13024,N_12541,N_12488);
nor U13025 (N_13025,N_12427,N_12880);
xor U13026 (N_13026,N_12449,N_12419);
nor U13027 (N_13027,N_12610,N_12696);
xor U13028 (N_13028,N_12742,N_12702);
and U13029 (N_13029,N_12271,N_12987);
xor U13030 (N_13030,N_12353,N_12525);
and U13031 (N_13031,N_12978,N_12332);
nor U13032 (N_13032,N_12947,N_12827);
or U13033 (N_13033,N_12807,N_12977);
or U13034 (N_13034,N_12422,N_12088);
nand U13035 (N_13035,N_12303,N_12191);
nand U13036 (N_13036,N_12877,N_12802);
and U13037 (N_13037,N_12083,N_12186);
and U13038 (N_13038,N_12786,N_12357);
and U13039 (N_13039,N_12416,N_12195);
nor U13040 (N_13040,N_12243,N_12912);
or U13041 (N_13041,N_12636,N_12476);
or U13042 (N_13042,N_12780,N_12594);
and U13043 (N_13043,N_12665,N_12025);
or U13044 (N_13044,N_12952,N_12925);
nand U13045 (N_13045,N_12405,N_12208);
or U13046 (N_13046,N_12626,N_12344);
and U13047 (N_13047,N_12051,N_12433);
nor U13048 (N_13048,N_12896,N_12089);
nor U13049 (N_13049,N_12413,N_12641);
nor U13050 (N_13050,N_12260,N_12699);
nor U13051 (N_13051,N_12826,N_12921);
nand U13052 (N_13052,N_12076,N_12735);
xor U13053 (N_13053,N_12572,N_12283);
or U13054 (N_13054,N_12772,N_12964);
nand U13055 (N_13055,N_12069,N_12124);
xnor U13056 (N_13056,N_12196,N_12408);
xor U13057 (N_13057,N_12540,N_12324);
nor U13058 (N_13058,N_12732,N_12642);
nor U13059 (N_13059,N_12275,N_12679);
and U13060 (N_13060,N_12431,N_12246);
nand U13061 (N_13061,N_12803,N_12333);
and U13062 (N_13062,N_12755,N_12494);
nand U13063 (N_13063,N_12864,N_12562);
xor U13064 (N_13064,N_12535,N_12597);
and U13065 (N_13065,N_12972,N_12748);
or U13066 (N_13066,N_12652,N_12976);
and U13067 (N_13067,N_12646,N_12458);
nor U13068 (N_13068,N_12653,N_12691);
or U13069 (N_13069,N_12619,N_12355);
and U13070 (N_13070,N_12147,N_12919);
or U13071 (N_13071,N_12436,N_12841);
and U13072 (N_13072,N_12187,N_12666);
or U13073 (N_13073,N_12484,N_12907);
xnor U13074 (N_13074,N_12139,N_12682);
or U13075 (N_13075,N_12614,N_12366);
nand U13076 (N_13076,N_12737,N_12032);
and U13077 (N_13077,N_12339,N_12725);
or U13078 (N_13078,N_12602,N_12517);
nand U13079 (N_13079,N_12277,N_12348);
nor U13080 (N_13080,N_12331,N_12995);
or U13081 (N_13081,N_12292,N_12820);
xnor U13082 (N_13082,N_12064,N_12059);
or U13083 (N_13083,N_12599,N_12204);
xnor U13084 (N_13084,N_12924,N_12960);
nand U13085 (N_13085,N_12074,N_12334);
nand U13086 (N_13086,N_12085,N_12138);
or U13087 (N_13087,N_12844,N_12903);
and U13088 (N_13088,N_12722,N_12643);
or U13089 (N_13089,N_12165,N_12385);
or U13090 (N_13090,N_12050,N_12487);
nor U13091 (N_13091,N_12233,N_12467);
xor U13092 (N_13092,N_12711,N_12582);
and U13093 (N_13093,N_12648,N_12273);
nor U13094 (N_13094,N_12095,N_12628);
nor U13095 (N_13095,N_12021,N_12272);
xnor U13096 (N_13096,N_12097,N_12612);
nand U13097 (N_13097,N_12701,N_12776);
and U13098 (N_13098,N_12609,N_12015);
nand U13099 (N_13099,N_12402,N_12515);
xor U13100 (N_13100,N_12664,N_12683);
nor U13101 (N_13101,N_12749,N_12293);
nor U13102 (N_13102,N_12909,N_12325);
nor U13103 (N_13103,N_12571,N_12881);
or U13104 (N_13104,N_12060,N_12278);
nand U13105 (N_13105,N_12751,N_12151);
nand U13106 (N_13106,N_12632,N_12931);
and U13107 (N_13107,N_12116,N_12489);
xnor U13108 (N_13108,N_12161,N_12045);
xor U13109 (N_13109,N_12115,N_12320);
nor U13110 (N_13110,N_12554,N_12983);
nor U13111 (N_13111,N_12508,N_12680);
nand U13112 (N_13112,N_12058,N_12241);
nor U13113 (N_13113,N_12308,N_12084);
and U13114 (N_13114,N_12746,N_12212);
and U13115 (N_13115,N_12893,N_12438);
nand U13116 (N_13116,N_12812,N_12849);
nand U13117 (N_13117,N_12577,N_12087);
and U13118 (N_13118,N_12140,N_12997);
or U13119 (N_13119,N_12499,N_12403);
nand U13120 (N_13120,N_12253,N_12012);
and U13121 (N_13121,N_12189,N_12791);
xnor U13122 (N_13122,N_12117,N_12713);
nor U13123 (N_13123,N_12676,N_12998);
or U13124 (N_13124,N_12839,N_12011);
nand U13125 (N_13125,N_12444,N_12475);
nand U13126 (N_13126,N_12975,N_12932);
xnor U13127 (N_13127,N_12689,N_12078);
nor U13128 (N_13128,N_12280,N_12586);
xor U13129 (N_13129,N_12093,N_12461);
nor U13130 (N_13130,N_12411,N_12407);
xnor U13131 (N_13131,N_12583,N_12209);
xnor U13132 (N_13132,N_12686,N_12048);
and U13133 (N_13133,N_12179,N_12591);
nand U13134 (N_13134,N_12613,N_12873);
and U13135 (N_13135,N_12125,N_12381);
or U13136 (N_13136,N_12622,N_12347);
and U13137 (N_13137,N_12834,N_12266);
nor U13138 (N_13138,N_12900,N_12930);
nor U13139 (N_13139,N_12647,N_12836);
nand U13140 (N_13140,N_12287,N_12598);
and U13141 (N_13141,N_12245,N_12669);
nor U13142 (N_13142,N_12235,N_12513);
and U13143 (N_13143,N_12443,N_12634);
or U13144 (N_13144,N_12731,N_12466);
or U13145 (N_13145,N_12869,N_12556);
nand U13146 (N_13146,N_12231,N_12670);
or U13147 (N_13147,N_12020,N_12349);
xor U13148 (N_13148,N_12172,N_12961);
xnor U13149 (N_13149,N_12741,N_12703);
xnor U13150 (N_13150,N_12234,N_12080);
nor U13151 (N_13151,N_12967,N_12870);
nor U13152 (N_13152,N_12144,N_12823);
or U13153 (N_13153,N_12090,N_12524);
nor U13154 (N_13154,N_12848,N_12340);
or U13155 (N_13155,N_12863,N_12657);
and U13156 (N_13156,N_12398,N_12430);
nand U13157 (N_13157,N_12254,N_12336);
or U13158 (N_13158,N_12829,N_12809);
nand U13159 (N_13159,N_12534,N_12585);
xor U13160 (N_13160,N_12224,N_12852);
xnor U13161 (N_13161,N_12004,N_12518);
xnor U13162 (N_13162,N_12215,N_12798);
xnor U13163 (N_13163,N_12067,N_12174);
and U13164 (N_13164,N_12356,N_12053);
xor U13165 (N_13165,N_12981,N_12171);
and U13166 (N_13166,N_12092,N_12744);
nor U13167 (N_13167,N_12070,N_12633);
nor U13168 (N_13168,N_12182,N_12386);
nand U13169 (N_13169,N_12491,N_12566);
and U13170 (N_13170,N_12351,N_12740);
nand U13171 (N_13171,N_12459,N_12133);
and U13172 (N_13172,N_12958,N_12079);
and U13173 (N_13173,N_12446,N_12859);
nand U13174 (N_13174,N_12238,N_12581);
nand U13175 (N_13175,N_12230,N_12939);
nor U13176 (N_13176,N_12569,N_12056);
or U13177 (N_13177,N_12804,N_12428);
nand U13178 (N_13178,N_12377,N_12482);
and U13179 (N_13179,N_12259,N_12604);
and U13180 (N_13180,N_12368,N_12014);
nor U13181 (N_13181,N_12201,N_12250);
nor U13182 (N_13182,N_12304,N_12143);
nand U13183 (N_13183,N_12156,N_12999);
xor U13184 (N_13184,N_12000,N_12335);
xor U13185 (N_13185,N_12282,N_12249);
xor U13186 (N_13186,N_12685,N_12075);
and U13187 (N_13187,N_12542,N_12327);
or U13188 (N_13188,N_12871,N_12592);
xor U13189 (N_13189,N_12183,N_12745);
nor U13190 (N_13190,N_12442,N_12522);
or U13191 (N_13191,N_12370,N_12547);
or U13192 (N_13192,N_12892,N_12982);
or U13193 (N_13193,N_12450,N_12031);
xor U13194 (N_13194,N_12166,N_12262);
nor U13195 (N_13195,N_12136,N_12825);
or U13196 (N_13196,N_12432,N_12922);
nand U13197 (N_13197,N_12593,N_12728);
and U13198 (N_13198,N_12644,N_12480);
and U13199 (N_13199,N_12949,N_12086);
nand U13200 (N_13200,N_12677,N_12270);
nand U13201 (N_13201,N_12322,N_12035);
xnor U13202 (N_13202,N_12039,N_12178);
and U13203 (N_13203,N_12984,N_12096);
nand U13204 (N_13204,N_12512,N_12126);
xnor U13205 (N_13205,N_12527,N_12727);
or U13206 (N_13206,N_12624,N_12396);
nand U13207 (N_13207,N_12106,N_12724);
nor U13208 (N_13208,N_12523,N_12605);
and U13209 (N_13209,N_12774,N_12412);
and U13210 (N_13210,N_12188,N_12862);
xnor U13211 (N_13211,N_12681,N_12710);
or U13212 (N_13212,N_12817,N_12819);
xnor U13213 (N_13213,N_12769,N_12107);
nand U13214 (N_13214,N_12955,N_12248);
nand U13215 (N_13215,N_12255,N_12658);
and U13216 (N_13216,N_12137,N_12113);
xnor U13217 (N_13217,N_12928,N_12917);
nor U13218 (N_13218,N_12575,N_12801);
nor U13219 (N_13219,N_12816,N_12994);
and U13220 (N_13220,N_12455,N_12543);
nand U13221 (N_13221,N_12199,N_12574);
or U13222 (N_13222,N_12800,N_12109);
or U13223 (N_13223,N_12152,N_12545);
xnor U13224 (N_13224,N_12164,N_12082);
and U13225 (N_13225,N_12009,N_12914);
and U13226 (N_13226,N_12497,N_12601);
nor U13227 (N_13227,N_12618,N_12034);
or U13228 (N_13228,N_12717,N_12211);
nand U13229 (N_13229,N_12226,N_12714);
and U13230 (N_13230,N_12496,N_12661);
nand U13231 (N_13231,N_12328,N_12429);
and U13232 (N_13232,N_12425,N_12589);
or U13233 (N_13233,N_12018,N_12252);
nand U13234 (N_13234,N_12962,N_12514);
nand U13235 (N_13235,N_12507,N_12898);
or U13236 (N_13236,N_12563,N_12625);
nor U13237 (N_13237,N_12447,N_12756);
nand U13238 (N_13238,N_12951,N_12206);
and U13239 (N_13239,N_12213,N_12342);
xor U13240 (N_13240,N_12923,N_12654);
xnor U13241 (N_13241,N_12072,N_12837);
or U13242 (N_13242,N_12406,N_12110);
or U13243 (N_13243,N_12440,N_12108);
or U13244 (N_13244,N_12926,N_12607);
nand U13245 (N_13245,N_12570,N_12920);
nand U13246 (N_13246,N_12306,N_12378);
nand U13247 (N_13247,N_12777,N_12695);
and U13248 (N_13248,N_12953,N_12806);
nor U13249 (N_13249,N_12866,N_12423);
or U13250 (N_13250,N_12519,N_12276);
and U13251 (N_13251,N_12568,N_12295);
xnor U13252 (N_13252,N_12565,N_12390);
nand U13253 (N_13253,N_12840,N_12875);
or U13254 (N_13254,N_12173,N_12767);
nand U13255 (N_13255,N_12558,N_12391);
or U13256 (N_13256,N_12662,N_12307);
nand U13257 (N_13257,N_12003,N_12845);
nand U13258 (N_13258,N_12452,N_12268);
nand U13259 (N_13259,N_12846,N_12300);
or U13260 (N_13260,N_12030,N_12621);
xor U13261 (N_13261,N_12752,N_12946);
nand U13262 (N_13262,N_12730,N_12131);
and U13263 (N_13263,N_12114,N_12770);
xor U13264 (N_13264,N_12822,N_12285);
and U13265 (N_13265,N_12828,N_12872);
nand U13266 (N_13266,N_12529,N_12672);
xor U13267 (N_13267,N_12036,N_12154);
xor U13268 (N_13268,N_12965,N_12623);
and U13269 (N_13269,N_12037,N_12057);
and U13270 (N_13270,N_12897,N_12323);
or U13271 (N_13271,N_12127,N_12103);
nor U13272 (N_13272,N_12916,N_12158);
or U13273 (N_13273,N_12874,N_12986);
and U13274 (N_13274,N_12155,N_12301);
xor U13275 (N_13275,N_12950,N_12134);
nor U13276 (N_13276,N_12971,N_12890);
nor U13277 (N_13277,N_12838,N_12936);
and U13278 (N_13278,N_12240,N_12105);
nand U13279 (N_13279,N_12477,N_12399);
or U13280 (N_13280,N_12966,N_12296);
and U13281 (N_13281,N_12445,N_12584);
xnor U13282 (N_13282,N_12371,N_12194);
xor U13283 (N_13283,N_12638,N_12375);
xor U13284 (N_13284,N_12933,N_12521);
nor U13285 (N_13285,N_12894,N_12042);
nand U13286 (N_13286,N_12705,N_12185);
or U13287 (N_13287,N_12062,N_12954);
or U13288 (N_13288,N_12790,N_12317);
xor U13289 (N_13289,N_12945,N_12659);
and U13290 (N_13290,N_12899,N_12046);
and U13291 (N_13291,N_12720,N_12363);
or U13292 (N_13292,N_12146,N_12373);
or U13293 (N_13293,N_12941,N_12678);
nor U13294 (N_13294,N_12792,N_12374);
xor U13295 (N_13295,N_12462,N_12942);
and U13296 (N_13296,N_12576,N_12660);
or U13297 (N_13297,N_12123,N_12564);
and U13298 (N_13298,N_12401,N_12441);
and U13299 (N_13299,N_12559,N_12232);
nand U13300 (N_13300,N_12162,N_12537);
nand U13301 (N_13301,N_12511,N_12734);
xor U13302 (N_13302,N_12805,N_12797);
and U13303 (N_13303,N_12198,N_12785);
xor U13304 (N_13304,N_12509,N_12153);
nor U13305 (N_13305,N_12148,N_12367);
nand U13306 (N_13306,N_12973,N_12553);
xor U13307 (N_13307,N_12434,N_12516);
and U13308 (N_13308,N_12560,N_12310);
or U13309 (N_13309,N_12747,N_12895);
nor U13310 (N_13310,N_12901,N_12810);
xnor U13311 (N_13311,N_12383,N_12974);
and U13312 (N_13312,N_12393,N_12218);
nor U13313 (N_13313,N_12929,N_12288);
nand U13314 (N_13314,N_12099,N_12073);
and U13315 (N_13315,N_12044,N_12478);
or U13316 (N_13316,N_12261,N_12066);
or U13317 (N_13317,N_12927,N_12091);
or U13318 (N_13318,N_12457,N_12400);
and U13319 (N_13319,N_12587,N_12674);
xor U13320 (N_13320,N_12128,N_12169);
and U13321 (N_13321,N_12055,N_12754);
or U13322 (N_13322,N_12361,N_12026);
xor U13323 (N_13323,N_12297,N_12799);
xnor U13324 (N_13324,N_12326,N_12555);
nand U13325 (N_13325,N_12733,N_12765);
and U13326 (N_13326,N_12708,N_12318);
xnor U13327 (N_13327,N_12520,N_12149);
or U13328 (N_13328,N_12192,N_12485);
and U13329 (N_13329,N_12236,N_12620);
nand U13330 (N_13330,N_12883,N_12460);
nor U13331 (N_13331,N_12397,N_12414);
nand U13332 (N_13332,N_12061,N_12163);
nand U13333 (N_13333,N_12779,N_12968);
nand U13334 (N_13334,N_12047,N_12410);
nor U13335 (N_13335,N_12160,N_12321);
xnor U13336 (N_13336,N_12309,N_12763);
and U13337 (N_13337,N_12963,N_12913);
nand U13338 (N_13338,N_12985,N_12193);
and U13339 (N_13339,N_12904,N_12854);
nand U13340 (N_13340,N_12650,N_12596);
nor U13341 (N_13341,N_12098,N_12019);
or U13342 (N_13342,N_12343,N_12630);
nor U13343 (N_13343,N_12121,N_12465);
nor U13344 (N_13344,N_12313,N_12842);
nor U13345 (N_13345,N_12530,N_12615);
nor U13346 (N_13346,N_12420,N_12448);
xnor U13347 (N_13347,N_12879,N_12022);
nor U13348 (N_13348,N_12228,N_12041);
nor U13349 (N_13349,N_12145,N_12969);
nor U13350 (N_13350,N_12510,N_12242);
nor U13351 (N_13351,N_12700,N_12207);
nor U13352 (N_13352,N_12435,N_12129);
xor U13353 (N_13353,N_12038,N_12492);
xnor U13354 (N_13354,N_12040,N_12365);
xor U13355 (N_13355,N_12017,N_12023);
or U13356 (N_13356,N_12284,N_12990);
nor U13357 (N_13357,N_12130,N_12891);
and U13358 (N_13358,N_12504,N_12081);
nor U13359 (N_13359,N_12119,N_12384);
nor U13360 (N_13360,N_12418,N_12906);
and U13361 (N_13361,N_12736,N_12346);
nor U13362 (N_13362,N_12389,N_12337);
nand U13363 (N_13363,N_12013,N_12993);
and U13364 (N_13364,N_12818,N_12168);
nand U13365 (N_13365,N_12635,N_12350);
or U13366 (N_13366,N_12684,N_12865);
or U13367 (N_13367,N_12008,N_12256);
and U13368 (N_13368,N_12766,N_12395);
nor U13369 (N_13369,N_12170,N_12549);
or U13370 (N_13370,N_12314,N_12750);
nand U13371 (N_13371,N_12716,N_12793);
and U13372 (N_13372,N_12908,N_12706);
nor U13373 (N_13373,N_12469,N_12608);
or U13374 (N_13374,N_12267,N_12225);
and U13375 (N_13375,N_12360,N_12421);
and U13376 (N_13376,N_12989,N_12426);
xor U13377 (N_13377,N_12220,N_12617);
nand U13378 (N_13378,N_12590,N_12120);
xnor U13379 (N_13379,N_12159,N_12637);
and U13380 (N_13380,N_12100,N_12782);
and U13381 (N_13381,N_12409,N_12001);
and U13382 (N_13382,N_12027,N_12698);
and U13383 (N_13383,N_12312,N_12723);
xor U13384 (N_13384,N_12831,N_12417);
nand U13385 (N_13385,N_12788,N_12758);
or U13386 (N_13386,N_12501,N_12289);
xor U13387 (N_13387,N_12552,N_12112);
nand U13388 (N_13388,N_12006,N_12505);
xnor U13389 (N_13389,N_12490,N_12404);
nor U13390 (N_13390,N_12824,N_12265);
xor U13391 (N_13391,N_12358,N_12821);
xor U13392 (N_13392,N_12111,N_12935);
and U13393 (N_13393,N_12005,N_12860);
xnor U13394 (N_13394,N_12239,N_12671);
nor U13395 (N_13395,N_12551,N_12264);
and U13396 (N_13396,N_12463,N_12269);
xor U13397 (N_13397,N_12392,N_12655);
xor U13398 (N_13398,N_12943,N_12707);
nand U13399 (N_13399,N_12453,N_12210);
or U13400 (N_13400,N_12719,N_12813);
nor U13401 (N_13401,N_12757,N_12851);
xnor U13402 (N_13402,N_12481,N_12667);
or U13403 (N_13403,N_12388,N_12544);
and U13404 (N_13404,N_12369,N_12474);
xnor U13405 (N_13405,N_12996,N_12694);
or U13406 (N_13406,N_12197,N_12850);
and U13407 (N_13407,N_12715,N_12726);
or U13408 (N_13408,N_12663,N_12135);
xor U13409 (N_13409,N_12071,N_12216);
nand U13410 (N_13410,N_12470,N_12251);
nand U13411 (N_13411,N_12815,N_12795);
xor U13412 (N_13412,N_12498,N_12010);
nor U13413 (N_13413,N_12376,N_12988);
nand U13414 (N_13414,N_12471,N_12603);
or U13415 (N_13415,N_12867,N_12203);
nor U13416 (N_13416,N_12611,N_12473);
or U13417 (N_13417,N_12506,N_12948);
xnor U13418 (N_13418,N_12007,N_12561);
or U13419 (N_13419,N_12102,N_12991);
and U13420 (N_13420,N_12631,N_12557);
xor U13421 (N_13421,N_12315,N_12104);
nand U13422 (N_13422,N_12709,N_12712);
and U13423 (N_13423,N_12762,N_12944);
xnor U13424 (N_13424,N_12299,N_12580);
nor U13425 (N_13425,N_12132,N_12673);
xnor U13426 (N_13426,N_12578,N_12219);
nand U13427 (N_13427,N_12853,N_12533);
or U13428 (N_13428,N_12302,N_12217);
nor U13429 (N_13429,N_12595,N_12649);
xor U13430 (N_13430,N_12796,N_12451);
and U13431 (N_13431,N_12294,N_12464);
nand U13432 (N_13432,N_12759,N_12486);
nand U13433 (N_13433,N_12258,N_12789);
and U13434 (N_13434,N_12316,N_12257);
nor U13435 (N_13435,N_12629,N_12915);
and U13436 (N_13436,N_12830,N_12808);
xor U13437 (N_13437,N_12910,N_12743);
nor U13438 (N_13438,N_12424,N_12500);
and U13439 (N_13439,N_12054,N_12052);
and U13440 (N_13440,N_12739,N_12675);
nor U13441 (N_13441,N_12319,N_12721);
nor U13442 (N_13442,N_12298,N_12959);
nand U13443 (N_13443,N_12532,N_12043);
or U13444 (N_13444,N_12550,N_12177);
nand U13445 (N_13445,N_12878,N_12503);
xnor U13446 (N_13446,N_12049,N_12833);
or U13447 (N_13447,N_12065,N_12068);
nor U13448 (N_13448,N_12141,N_12843);
or U13449 (N_13449,N_12934,N_12783);
xnor U13450 (N_13450,N_12876,N_12184);
xor U13451 (N_13451,N_12773,N_12362);
nand U13452 (N_13452,N_12905,N_12033);
nand U13453 (N_13453,N_12528,N_12588);
and U13454 (N_13454,N_12200,N_12814);
nand U13455 (N_13455,N_12345,N_12077);
nand U13456 (N_13456,N_12495,N_12190);
nor U13457 (N_13457,N_12468,N_12341);
and U13458 (N_13458,N_12483,N_12979);
and U13459 (N_13459,N_12918,N_12002);
nor U13460 (N_13460,N_12692,N_12600);
and U13461 (N_13461,N_12263,N_12531);
or U13462 (N_13462,N_12222,N_12394);
xor U13463 (N_13463,N_12279,N_12882);
and U13464 (N_13464,N_12237,N_12794);
xnor U13465 (N_13465,N_12771,N_12380);
xor U13466 (N_13466,N_12956,N_12639);
and U13467 (N_13467,N_12223,N_12548);
or U13468 (N_13468,N_12761,N_12311);
or U13469 (N_13469,N_12536,N_12889);
and U13470 (N_13470,N_12937,N_12437);
nand U13471 (N_13471,N_12502,N_12858);
and U13472 (N_13472,N_12247,N_12329);
nand U13473 (N_13473,N_12372,N_12764);
xor U13474 (N_13474,N_12456,N_12835);
or U13475 (N_13475,N_12718,N_12167);
or U13476 (N_13476,N_12330,N_12992);
or U13477 (N_13477,N_12778,N_12606);
xnor U13478 (N_13478,N_12180,N_12479);
nor U13479 (N_13479,N_12364,N_12538);
nand U13480 (N_13480,N_12627,N_12656);
or U13481 (N_13481,N_12775,N_12359);
or U13482 (N_13482,N_12028,N_12886);
xnor U13483 (N_13483,N_12688,N_12668);
nand U13484 (N_13484,N_12911,N_12938);
and U13485 (N_13485,N_12957,N_12352);
and U13486 (N_13486,N_12940,N_12857);
nand U13487 (N_13487,N_12567,N_12382);
xor U13488 (N_13488,N_12526,N_12729);
nor U13489 (N_13489,N_12016,N_12781);
and U13490 (N_13490,N_12855,N_12811);
nor U13491 (N_13491,N_12472,N_12768);
nor U13492 (N_13492,N_12970,N_12887);
or U13493 (N_13493,N_12229,N_12291);
nor U13494 (N_13494,N_12118,N_12063);
nor U13495 (N_13495,N_12753,N_12338);
nor U13496 (N_13496,N_12760,N_12573);
xnor U13497 (N_13497,N_12579,N_12687);
nor U13498 (N_13498,N_12274,N_12387);
and U13499 (N_13499,N_12221,N_12290);
xnor U13500 (N_13500,N_12602,N_12830);
or U13501 (N_13501,N_12794,N_12914);
xnor U13502 (N_13502,N_12385,N_12939);
nor U13503 (N_13503,N_12191,N_12377);
and U13504 (N_13504,N_12751,N_12899);
or U13505 (N_13505,N_12946,N_12075);
xor U13506 (N_13506,N_12032,N_12866);
nand U13507 (N_13507,N_12854,N_12322);
xnor U13508 (N_13508,N_12428,N_12193);
or U13509 (N_13509,N_12180,N_12197);
and U13510 (N_13510,N_12717,N_12419);
nand U13511 (N_13511,N_12200,N_12802);
nand U13512 (N_13512,N_12109,N_12697);
nand U13513 (N_13513,N_12370,N_12567);
or U13514 (N_13514,N_12602,N_12310);
and U13515 (N_13515,N_12381,N_12796);
nand U13516 (N_13516,N_12942,N_12693);
nor U13517 (N_13517,N_12313,N_12520);
or U13518 (N_13518,N_12837,N_12621);
or U13519 (N_13519,N_12343,N_12163);
nor U13520 (N_13520,N_12076,N_12380);
or U13521 (N_13521,N_12605,N_12000);
nand U13522 (N_13522,N_12595,N_12869);
or U13523 (N_13523,N_12200,N_12097);
xnor U13524 (N_13524,N_12910,N_12374);
and U13525 (N_13525,N_12039,N_12408);
xor U13526 (N_13526,N_12143,N_12467);
nand U13527 (N_13527,N_12881,N_12482);
xor U13528 (N_13528,N_12477,N_12460);
xnor U13529 (N_13529,N_12846,N_12996);
nand U13530 (N_13530,N_12959,N_12978);
or U13531 (N_13531,N_12851,N_12180);
nor U13532 (N_13532,N_12802,N_12989);
or U13533 (N_13533,N_12642,N_12068);
nor U13534 (N_13534,N_12178,N_12754);
and U13535 (N_13535,N_12119,N_12593);
or U13536 (N_13536,N_12444,N_12788);
xnor U13537 (N_13537,N_12210,N_12194);
or U13538 (N_13538,N_12586,N_12549);
and U13539 (N_13539,N_12788,N_12486);
or U13540 (N_13540,N_12502,N_12462);
or U13541 (N_13541,N_12149,N_12901);
or U13542 (N_13542,N_12026,N_12258);
xnor U13543 (N_13543,N_12027,N_12413);
and U13544 (N_13544,N_12057,N_12313);
nand U13545 (N_13545,N_12581,N_12871);
nor U13546 (N_13546,N_12890,N_12572);
or U13547 (N_13547,N_12307,N_12173);
xnor U13548 (N_13548,N_12547,N_12516);
nand U13549 (N_13549,N_12360,N_12127);
nor U13550 (N_13550,N_12913,N_12132);
nor U13551 (N_13551,N_12695,N_12020);
or U13552 (N_13552,N_12800,N_12360);
nor U13553 (N_13553,N_12457,N_12244);
nand U13554 (N_13554,N_12134,N_12338);
nor U13555 (N_13555,N_12225,N_12197);
or U13556 (N_13556,N_12338,N_12415);
nor U13557 (N_13557,N_12074,N_12018);
and U13558 (N_13558,N_12144,N_12059);
nor U13559 (N_13559,N_12488,N_12896);
xor U13560 (N_13560,N_12328,N_12407);
or U13561 (N_13561,N_12101,N_12928);
xor U13562 (N_13562,N_12463,N_12323);
nand U13563 (N_13563,N_12525,N_12401);
xnor U13564 (N_13564,N_12328,N_12338);
nor U13565 (N_13565,N_12151,N_12153);
xnor U13566 (N_13566,N_12363,N_12539);
and U13567 (N_13567,N_12448,N_12692);
nand U13568 (N_13568,N_12587,N_12453);
nand U13569 (N_13569,N_12272,N_12908);
nand U13570 (N_13570,N_12017,N_12350);
xor U13571 (N_13571,N_12306,N_12009);
xnor U13572 (N_13572,N_12939,N_12483);
xor U13573 (N_13573,N_12684,N_12265);
xnor U13574 (N_13574,N_12183,N_12737);
and U13575 (N_13575,N_12490,N_12686);
xor U13576 (N_13576,N_12196,N_12108);
and U13577 (N_13577,N_12565,N_12596);
and U13578 (N_13578,N_12184,N_12077);
xor U13579 (N_13579,N_12155,N_12400);
or U13580 (N_13580,N_12979,N_12339);
and U13581 (N_13581,N_12790,N_12144);
nor U13582 (N_13582,N_12654,N_12402);
xor U13583 (N_13583,N_12265,N_12967);
nand U13584 (N_13584,N_12503,N_12071);
xnor U13585 (N_13585,N_12875,N_12785);
or U13586 (N_13586,N_12168,N_12401);
nand U13587 (N_13587,N_12282,N_12299);
nor U13588 (N_13588,N_12522,N_12541);
or U13589 (N_13589,N_12052,N_12356);
xor U13590 (N_13590,N_12798,N_12773);
nand U13591 (N_13591,N_12312,N_12860);
nor U13592 (N_13592,N_12618,N_12817);
nand U13593 (N_13593,N_12098,N_12525);
and U13594 (N_13594,N_12264,N_12289);
xnor U13595 (N_13595,N_12624,N_12299);
xor U13596 (N_13596,N_12959,N_12615);
nand U13597 (N_13597,N_12058,N_12627);
xnor U13598 (N_13598,N_12994,N_12760);
and U13599 (N_13599,N_12441,N_12354);
or U13600 (N_13600,N_12822,N_12462);
nor U13601 (N_13601,N_12240,N_12159);
and U13602 (N_13602,N_12169,N_12601);
nor U13603 (N_13603,N_12113,N_12375);
or U13604 (N_13604,N_12180,N_12605);
xnor U13605 (N_13605,N_12447,N_12973);
nor U13606 (N_13606,N_12571,N_12930);
xnor U13607 (N_13607,N_12297,N_12449);
xnor U13608 (N_13608,N_12751,N_12082);
nor U13609 (N_13609,N_12207,N_12011);
nor U13610 (N_13610,N_12366,N_12244);
xor U13611 (N_13611,N_12188,N_12821);
xnor U13612 (N_13612,N_12553,N_12199);
nand U13613 (N_13613,N_12664,N_12007);
nand U13614 (N_13614,N_12787,N_12795);
or U13615 (N_13615,N_12584,N_12050);
nand U13616 (N_13616,N_12156,N_12412);
xnor U13617 (N_13617,N_12326,N_12474);
xor U13618 (N_13618,N_12495,N_12461);
nand U13619 (N_13619,N_12255,N_12097);
and U13620 (N_13620,N_12861,N_12149);
xnor U13621 (N_13621,N_12228,N_12546);
nand U13622 (N_13622,N_12562,N_12406);
and U13623 (N_13623,N_12180,N_12269);
nor U13624 (N_13624,N_12763,N_12162);
nor U13625 (N_13625,N_12187,N_12689);
xnor U13626 (N_13626,N_12786,N_12938);
and U13627 (N_13627,N_12434,N_12033);
nand U13628 (N_13628,N_12864,N_12418);
xor U13629 (N_13629,N_12523,N_12228);
or U13630 (N_13630,N_12994,N_12540);
nand U13631 (N_13631,N_12204,N_12647);
nor U13632 (N_13632,N_12651,N_12468);
xor U13633 (N_13633,N_12820,N_12214);
nor U13634 (N_13634,N_12967,N_12358);
nand U13635 (N_13635,N_12507,N_12387);
or U13636 (N_13636,N_12385,N_12584);
and U13637 (N_13637,N_12123,N_12234);
nand U13638 (N_13638,N_12017,N_12385);
and U13639 (N_13639,N_12182,N_12557);
or U13640 (N_13640,N_12005,N_12573);
or U13641 (N_13641,N_12310,N_12497);
nor U13642 (N_13642,N_12215,N_12726);
nor U13643 (N_13643,N_12855,N_12089);
nand U13644 (N_13644,N_12277,N_12119);
and U13645 (N_13645,N_12445,N_12765);
and U13646 (N_13646,N_12095,N_12252);
or U13647 (N_13647,N_12699,N_12858);
nand U13648 (N_13648,N_12992,N_12174);
nor U13649 (N_13649,N_12960,N_12489);
and U13650 (N_13650,N_12367,N_12879);
xor U13651 (N_13651,N_12177,N_12484);
nor U13652 (N_13652,N_12720,N_12355);
nor U13653 (N_13653,N_12415,N_12251);
nand U13654 (N_13654,N_12890,N_12937);
xnor U13655 (N_13655,N_12148,N_12415);
nand U13656 (N_13656,N_12661,N_12883);
and U13657 (N_13657,N_12040,N_12297);
nand U13658 (N_13658,N_12760,N_12804);
xnor U13659 (N_13659,N_12618,N_12109);
or U13660 (N_13660,N_12045,N_12627);
and U13661 (N_13661,N_12965,N_12917);
and U13662 (N_13662,N_12779,N_12324);
and U13663 (N_13663,N_12034,N_12251);
and U13664 (N_13664,N_12477,N_12358);
xor U13665 (N_13665,N_12111,N_12900);
nor U13666 (N_13666,N_12115,N_12855);
nor U13667 (N_13667,N_12173,N_12584);
or U13668 (N_13668,N_12989,N_12135);
nor U13669 (N_13669,N_12286,N_12795);
and U13670 (N_13670,N_12983,N_12242);
or U13671 (N_13671,N_12025,N_12274);
nand U13672 (N_13672,N_12562,N_12074);
and U13673 (N_13673,N_12428,N_12621);
xor U13674 (N_13674,N_12856,N_12766);
nor U13675 (N_13675,N_12627,N_12946);
or U13676 (N_13676,N_12760,N_12981);
or U13677 (N_13677,N_12322,N_12725);
xor U13678 (N_13678,N_12290,N_12507);
xnor U13679 (N_13679,N_12384,N_12650);
and U13680 (N_13680,N_12800,N_12133);
nand U13681 (N_13681,N_12383,N_12709);
and U13682 (N_13682,N_12950,N_12401);
nand U13683 (N_13683,N_12190,N_12423);
and U13684 (N_13684,N_12463,N_12022);
or U13685 (N_13685,N_12041,N_12495);
nand U13686 (N_13686,N_12728,N_12067);
and U13687 (N_13687,N_12123,N_12962);
nand U13688 (N_13688,N_12311,N_12236);
and U13689 (N_13689,N_12302,N_12152);
nor U13690 (N_13690,N_12132,N_12674);
nand U13691 (N_13691,N_12051,N_12369);
xnor U13692 (N_13692,N_12415,N_12416);
xor U13693 (N_13693,N_12423,N_12660);
xnor U13694 (N_13694,N_12909,N_12279);
nor U13695 (N_13695,N_12107,N_12699);
and U13696 (N_13696,N_12920,N_12343);
xor U13697 (N_13697,N_12213,N_12922);
or U13698 (N_13698,N_12890,N_12686);
nand U13699 (N_13699,N_12310,N_12951);
or U13700 (N_13700,N_12469,N_12326);
xor U13701 (N_13701,N_12948,N_12703);
xor U13702 (N_13702,N_12264,N_12111);
or U13703 (N_13703,N_12721,N_12513);
nand U13704 (N_13704,N_12474,N_12453);
nand U13705 (N_13705,N_12463,N_12306);
xnor U13706 (N_13706,N_12093,N_12549);
and U13707 (N_13707,N_12563,N_12184);
nand U13708 (N_13708,N_12653,N_12843);
xnor U13709 (N_13709,N_12358,N_12504);
nor U13710 (N_13710,N_12547,N_12243);
nor U13711 (N_13711,N_12468,N_12493);
nand U13712 (N_13712,N_12289,N_12333);
xor U13713 (N_13713,N_12597,N_12411);
or U13714 (N_13714,N_12971,N_12504);
nor U13715 (N_13715,N_12701,N_12281);
xnor U13716 (N_13716,N_12197,N_12685);
nand U13717 (N_13717,N_12006,N_12598);
or U13718 (N_13718,N_12887,N_12203);
nor U13719 (N_13719,N_12804,N_12988);
xnor U13720 (N_13720,N_12775,N_12481);
and U13721 (N_13721,N_12511,N_12292);
and U13722 (N_13722,N_12033,N_12946);
or U13723 (N_13723,N_12126,N_12907);
or U13724 (N_13724,N_12393,N_12986);
xor U13725 (N_13725,N_12407,N_12717);
nand U13726 (N_13726,N_12099,N_12368);
nand U13727 (N_13727,N_12961,N_12242);
and U13728 (N_13728,N_12823,N_12519);
or U13729 (N_13729,N_12920,N_12705);
xor U13730 (N_13730,N_12274,N_12352);
or U13731 (N_13731,N_12121,N_12905);
and U13732 (N_13732,N_12465,N_12185);
nand U13733 (N_13733,N_12921,N_12539);
nor U13734 (N_13734,N_12921,N_12271);
xnor U13735 (N_13735,N_12092,N_12577);
nor U13736 (N_13736,N_12176,N_12041);
nand U13737 (N_13737,N_12784,N_12893);
or U13738 (N_13738,N_12553,N_12074);
or U13739 (N_13739,N_12659,N_12917);
xnor U13740 (N_13740,N_12787,N_12059);
nor U13741 (N_13741,N_12808,N_12242);
xor U13742 (N_13742,N_12464,N_12552);
and U13743 (N_13743,N_12454,N_12971);
xor U13744 (N_13744,N_12278,N_12650);
nand U13745 (N_13745,N_12666,N_12914);
or U13746 (N_13746,N_12286,N_12124);
nand U13747 (N_13747,N_12998,N_12809);
and U13748 (N_13748,N_12052,N_12535);
nand U13749 (N_13749,N_12821,N_12577);
and U13750 (N_13750,N_12898,N_12993);
and U13751 (N_13751,N_12873,N_12533);
nor U13752 (N_13752,N_12768,N_12619);
or U13753 (N_13753,N_12257,N_12347);
nand U13754 (N_13754,N_12711,N_12957);
nor U13755 (N_13755,N_12687,N_12699);
nor U13756 (N_13756,N_12763,N_12853);
xnor U13757 (N_13757,N_12769,N_12638);
nand U13758 (N_13758,N_12722,N_12397);
and U13759 (N_13759,N_12892,N_12688);
nand U13760 (N_13760,N_12493,N_12959);
nand U13761 (N_13761,N_12722,N_12684);
or U13762 (N_13762,N_12093,N_12546);
nor U13763 (N_13763,N_12475,N_12092);
nand U13764 (N_13764,N_12942,N_12934);
xnor U13765 (N_13765,N_12727,N_12198);
xor U13766 (N_13766,N_12198,N_12937);
and U13767 (N_13767,N_12649,N_12100);
xor U13768 (N_13768,N_12639,N_12361);
or U13769 (N_13769,N_12717,N_12223);
xnor U13770 (N_13770,N_12286,N_12835);
xor U13771 (N_13771,N_12865,N_12593);
xnor U13772 (N_13772,N_12960,N_12461);
nor U13773 (N_13773,N_12781,N_12027);
nor U13774 (N_13774,N_12342,N_12945);
and U13775 (N_13775,N_12157,N_12692);
or U13776 (N_13776,N_12774,N_12711);
or U13777 (N_13777,N_12756,N_12579);
xor U13778 (N_13778,N_12947,N_12708);
nor U13779 (N_13779,N_12376,N_12925);
and U13780 (N_13780,N_12302,N_12361);
or U13781 (N_13781,N_12083,N_12959);
or U13782 (N_13782,N_12733,N_12622);
xor U13783 (N_13783,N_12785,N_12798);
nand U13784 (N_13784,N_12292,N_12124);
nand U13785 (N_13785,N_12381,N_12033);
or U13786 (N_13786,N_12935,N_12394);
nor U13787 (N_13787,N_12226,N_12555);
nor U13788 (N_13788,N_12841,N_12781);
or U13789 (N_13789,N_12593,N_12710);
and U13790 (N_13790,N_12703,N_12566);
nor U13791 (N_13791,N_12729,N_12906);
and U13792 (N_13792,N_12497,N_12053);
and U13793 (N_13793,N_12628,N_12631);
xor U13794 (N_13794,N_12067,N_12872);
xnor U13795 (N_13795,N_12694,N_12349);
xnor U13796 (N_13796,N_12025,N_12941);
nor U13797 (N_13797,N_12900,N_12802);
nor U13798 (N_13798,N_12371,N_12206);
and U13799 (N_13799,N_12252,N_12668);
nor U13800 (N_13800,N_12509,N_12367);
or U13801 (N_13801,N_12536,N_12357);
nand U13802 (N_13802,N_12502,N_12856);
nand U13803 (N_13803,N_12896,N_12640);
or U13804 (N_13804,N_12248,N_12556);
nor U13805 (N_13805,N_12705,N_12269);
or U13806 (N_13806,N_12650,N_12125);
nor U13807 (N_13807,N_12518,N_12993);
nor U13808 (N_13808,N_12541,N_12799);
xnor U13809 (N_13809,N_12799,N_12222);
nand U13810 (N_13810,N_12368,N_12293);
or U13811 (N_13811,N_12207,N_12052);
and U13812 (N_13812,N_12357,N_12359);
nand U13813 (N_13813,N_12136,N_12293);
nor U13814 (N_13814,N_12165,N_12371);
xor U13815 (N_13815,N_12809,N_12136);
and U13816 (N_13816,N_12388,N_12040);
or U13817 (N_13817,N_12530,N_12478);
xnor U13818 (N_13818,N_12276,N_12479);
and U13819 (N_13819,N_12704,N_12432);
xnor U13820 (N_13820,N_12950,N_12718);
or U13821 (N_13821,N_12086,N_12240);
or U13822 (N_13822,N_12226,N_12761);
nand U13823 (N_13823,N_12441,N_12906);
and U13824 (N_13824,N_12846,N_12347);
or U13825 (N_13825,N_12369,N_12486);
nand U13826 (N_13826,N_12598,N_12051);
nor U13827 (N_13827,N_12275,N_12877);
nand U13828 (N_13828,N_12643,N_12857);
and U13829 (N_13829,N_12436,N_12658);
nand U13830 (N_13830,N_12727,N_12043);
or U13831 (N_13831,N_12430,N_12838);
nand U13832 (N_13832,N_12274,N_12497);
xnor U13833 (N_13833,N_12876,N_12146);
and U13834 (N_13834,N_12760,N_12797);
and U13835 (N_13835,N_12333,N_12080);
nor U13836 (N_13836,N_12161,N_12790);
and U13837 (N_13837,N_12827,N_12474);
and U13838 (N_13838,N_12531,N_12710);
xnor U13839 (N_13839,N_12970,N_12956);
nand U13840 (N_13840,N_12381,N_12830);
or U13841 (N_13841,N_12072,N_12043);
nand U13842 (N_13842,N_12377,N_12188);
and U13843 (N_13843,N_12690,N_12321);
nand U13844 (N_13844,N_12476,N_12697);
nor U13845 (N_13845,N_12431,N_12496);
nor U13846 (N_13846,N_12954,N_12915);
xnor U13847 (N_13847,N_12212,N_12485);
xor U13848 (N_13848,N_12084,N_12332);
nand U13849 (N_13849,N_12627,N_12587);
nand U13850 (N_13850,N_12638,N_12331);
xor U13851 (N_13851,N_12644,N_12153);
or U13852 (N_13852,N_12836,N_12944);
nand U13853 (N_13853,N_12674,N_12805);
nand U13854 (N_13854,N_12015,N_12656);
nor U13855 (N_13855,N_12565,N_12010);
nor U13856 (N_13856,N_12269,N_12893);
or U13857 (N_13857,N_12874,N_12757);
and U13858 (N_13858,N_12258,N_12979);
nand U13859 (N_13859,N_12803,N_12112);
nand U13860 (N_13860,N_12925,N_12928);
and U13861 (N_13861,N_12461,N_12400);
xor U13862 (N_13862,N_12543,N_12468);
nand U13863 (N_13863,N_12810,N_12691);
nand U13864 (N_13864,N_12630,N_12362);
and U13865 (N_13865,N_12849,N_12566);
and U13866 (N_13866,N_12604,N_12070);
nand U13867 (N_13867,N_12295,N_12274);
nand U13868 (N_13868,N_12317,N_12883);
nand U13869 (N_13869,N_12250,N_12322);
or U13870 (N_13870,N_12309,N_12877);
nor U13871 (N_13871,N_12883,N_12226);
xor U13872 (N_13872,N_12126,N_12728);
xor U13873 (N_13873,N_12909,N_12357);
xnor U13874 (N_13874,N_12743,N_12349);
nor U13875 (N_13875,N_12392,N_12630);
nand U13876 (N_13876,N_12028,N_12470);
nand U13877 (N_13877,N_12266,N_12907);
and U13878 (N_13878,N_12519,N_12283);
or U13879 (N_13879,N_12498,N_12078);
or U13880 (N_13880,N_12507,N_12835);
xnor U13881 (N_13881,N_12651,N_12510);
nor U13882 (N_13882,N_12349,N_12885);
or U13883 (N_13883,N_12950,N_12392);
and U13884 (N_13884,N_12905,N_12044);
xnor U13885 (N_13885,N_12771,N_12265);
and U13886 (N_13886,N_12338,N_12824);
nand U13887 (N_13887,N_12173,N_12306);
or U13888 (N_13888,N_12890,N_12770);
nor U13889 (N_13889,N_12142,N_12927);
or U13890 (N_13890,N_12160,N_12827);
nand U13891 (N_13891,N_12277,N_12534);
nand U13892 (N_13892,N_12310,N_12142);
and U13893 (N_13893,N_12885,N_12442);
or U13894 (N_13894,N_12396,N_12802);
or U13895 (N_13895,N_12896,N_12297);
nand U13896 (N_13896,N_12584,N_12280);
or U13897 (N_13897,N_12646,N_12883);
nor U13898 (N_13898,N_12699,N_12325);
and U13899 (N_13899,N_12637,N_12848);
nor U13900 (N_13900,N_12571,N_12816);
or U13901 (N_13901,N_12928,N_12794);
nor U13902 (N_13902,N_12751,N_12893);
xnor U13903 (N_13903,N_12952,N_12601);
xnor U13904 (N_13904,N_12731,N_12107);
and U13905 (N_13905,N_12460,N_12703);
nand U13906 (N_13906,N_12997,N_12665);
and U13907 (N_13907,N_12013,N_12367);
and U13908 (N_13908,N_12706,N_12617);
xnor U13909 (N_13909,N_12246,N_12331);
nor U13910 (N_13910,N_12956,N_12545);
and U13911 (N_13911,N_12534,N_12502);
nand U13912 (N_13912,N_12845,N_12415);
nor U13913 (N_13913,N_12759,N_12701);
and U13914 (N_13914,N_12706,N_12588);
and U13915 (N_13915,N_12010,N_12695);
xnor U13916 (N_13916,N_12816,N_12631);
xnor U13917 (N_13917,N_12679,N_12089);
and U13918 (N_13918,N_12541,N_12994);
nor U13919 (N_13919,N_12743,N_12978);
nand U13920 (N_13920,N_12349,N_12499);
nor U13921 (N_13921,N_12829,N_12978);
nand U13922 (N_13922,N_12749,N_12277);
or U13923 (N_13923,N_12608,N_12007);
and U13924 (N_13924,N_12805,N_12803);
and U13925 (N_13925,N_12569,N_12079);
nor U13926 (N_13926,N_12024,N_12267);
xnor U13927 (N_13927,N_12492,N_12706);
nor U13928 (N_13928,N_12948,N_12995);
xor U13929 (N_13929,N_12834,N_12599);
and U13930 (N_13930,N_12419,N_12122);
nor U13931 (N_13931,N_12940,N_12860);
nand U13932 (N_13932,N_12722,N_12051);
xnor U13933 (N_13933,N_12866,N_12748);
nand U13934 (N_13934,N_12333,N_12124);
xnor U13935 (N_13935,N_12635,N_12392);
xnor U13936 (N_13936,N_12115,N_12923);
nor U13937 (N_13937,N_12928,N_12111);
nor U13938 (N_13938,N_12391,N_12171);
nand U13939 (N_13939,N_12357,N_12041);
nand U13940 (N_13940,N_12183,N_12700);
nand U13941 (N_13941,N_12199,N_12242);
nor U13942 (N_13942,N_12484,N_12532);
or U13943 (N_13943,N_12843,N_12034);
xnor U13944 (N_13944,N_12323,N_12910);
nor U13945 (N_13945,N_12956,N_12006);
xnor U13946 (N_13946,N_12014,N_12042);
xnor U13947 (N_13947,N_12975,N_12740);
nand U13948 (N_13948,N_12200,N_12942);
nand U13949 (N_13949,N_12631,N_12379);
xor U13950 (N_13950,N_12743,N_12635);
or U13951 (N_13951,N_12013,N_12983);
xor U13952 (N_13952,N_12555,N_12554);
nand U13953 (N_13953,N_12862,N_12717);
nor U13954 (N_13954,N_12227,N_12440);
nand U13955 (N_13955,N_12235,N_12532);
and U13956 (N_13956,N_12192,N_12441);
nor U13957 (N_13957,N_12521,N_12342);
nand U13958 (N_13958,N_12720,N_12049);
and U13959 (N_13959,N_12755,N_12133);
nor U13960 (N_13960,N_12485,N_12446);
or U13961 (N_13961,N_12083,N_12970);
nor U13962 (N_13962,N_12466,N_12610);
xnor U13963 (N_13963,N_12035,N_12779);
or U13964 (N_13964,N_12392,N_12278);
xor U13965 (N_13965,N_12400,N_12999);
or U13966 (N_13966,N_12420,N_12715);
or U13967 (N_13967,N_12547,N_12987);
or U13968 (N_13968,N_12793,N_12157);
and U13969 (N_13969,N_12874,N_12313);
nand U13970 (N_13970,N_12712,N_12065);
nor U13971 (N_13971,N_12877,N_12207);
and U13972 (N_13972,N_12997,N_12024);
or U13973 (N_13973,N_12665,N_12999);
or U13974 (N_13974,N_12960,N_12786);
nor U13975 (N_13975,N_12135,N_12389);
or U13976 (N_13976,N_12951,N_12367);
nand U13977 (N_13977,N_12719,N_12570);
or U13978 (N_13978,N_12659,N_12507);
xnor U13979 (N_13979,N_12820,N_12440);
nor U13980 (N_13980,N_12595,N_12094);
nand U13981 (N_13981,N_12779,N_12392);
xor U13982 (N_13982,N_12632,N_12099);
or U13983 (N_13983,N_12081,N_12573);
xor U13984 (N_13984,N_12367,N_12010);
or U13985 (N_13985,N_12903,N_12824);
or U13986 (N_13986,N_12697,N_12946);
and U13987 (N_13987,N_12358,N_12902);
nor U13988 (N_13988,N_12400,N_12525);
or U13989 (N_13989,N_12717,N_12567);
nor U13990 (N_13990,N_12500,N_12060);
and U13991 (N_13991,N_12610,N_12491);
xnor U13992 (N_13992,N_12848,N_12089);
xor U13993 (N_13993,N_12363,N_12733);
nand U13994 (N_13994,N_12248,N_12243);
xnor U13995 (N_13995,N_12353,N_12238);
xor U13996 (N_13996,N_12636,N_12699);
and U13997 (N_13997,N_12595,N_12975);
and U13998 (N_13998,N_12987,N_12828);
nand U13999 (N_13999,N_12197,N_12792);
nor U14000 (N_14000,N_13559,N_13404);
and U14001 (N_14001,N_13117,N_13978);
xor U14002 (N_14002,N_13202,N_13287);
or U14003 (N_14003,N_13188,N_13821);
nand U14004 (N_14004,N_13132,N_13000);
nand U14005 (N_14005,N_13951,N_13517);
or U14006 (N_14006,N_13244,N_13363);
or U14007 (N_14007,N_13221,N_13159);
and U14008 (N_14008,N_13151,N_13591);
nand U14009 (N_14009,N_13901,N_13937);
nand U14010 (N_14010,N_13759,N_13869);
nor U14011 (N_14011,N_13085,N_13386);
or U14012 (N_14012,N_13375,N_13235);
nor U14013 (N_14013,N_13447,N_13825);
or U14014 (N_14014,N_13499,N_13753);
or U14015 (N_14015,N_13190,N_13277);
nor U14016 (N_14016,N_13627,N_13981);
nand U14017 (N_14017,N_13785,N_13053);
or U14018 (N_14018,N_13963,N_13373);
nand U14019 (N_14019,N_13947,N_13959);
xor U14020 (N_14020,N_13899,N_13016);
nand U14021 (N_14021,N_13693,N_13496);
and U14022 (N_14022,N_13193,N_13838);
and U14023 (N_14023,N_13628,N_13859);
nor U14024 (N_14024,N_13040,N_13397);
and U14025 (N_14025,N_13174,N_13676);
and U14026 (N_14026,N_13433,N_13633);
nand U14027 (N_14027,N_13649,N_13605);
and U14028 (N_14028,N_13906,N_13957);
nand U14029 (N_14029,N_13055,N_13894);
xor U14030 (N_14030,N_13695,N_13086);
and U14031 (N_14031,N_13245,N_13511);
nor U14032 (N_14032,N_13538,N_13673);
xnor U14033 (N_14033,N_13961,N_13357);
and U14034 (N_14034,N_13896,N_13301);
or U14035 (N_14035,N_13791,N_13032);
xnor U14036 (N_14036,N_13989,N_13781);
nor U14037 (N_14037,N_13598,N_13294);
or U14038 (N_14038,N_13914,N_13281);
nand U14039 (N_14039,N_13526,N_13630);
and U14040 (N_14040,N_13109,N_13594);
and U14041 (N_14041,N_13694,N_13900);
nor U14042 (N_14042,N_13350,N_13782);
nand U14043 (N_14043,N_13269,N_13824);
nand U14044 (N_14044,N_13437,N_13565);
or U14045 (N_14045,N_13846,N_13420);
xnor U14046 (N_14046,N_13201,N_13005);
and U14047 (N_14047,N_13442,N_13857);
xor U14048 (N_14048,N_13060,N_13495);
nor U14049 (N_14049,N_13296,N_13042);
or U14050 (N_14050,N_13012,N_13931);
nand U14051 (N_14051,N_13264,N_13586);
nor U14052 (N_14052,N_13096,N_13196);
nor U14053 (N_14053,N_13229,N_13471);
nor U14054 (N_14054,N_13584,N_13094);
and U14055 (N_14055,N_13172,N_13661);
nor U14056 (N_14056,N_13431,N_13122);
and U14057 (N_14057,N_13432,N_13529);
xnor U14058 (N_14058,N_13589,N_13226);
nor U14059 (N_14059,N_13275,N_13473);
nor U14060 (N_14060,N_13276,N_13504);
or U14061 (N_14061,N_13465,N_13166);
or U14062 (N_14062,N_13116,N_13257);
or U14063 (N_14063,N_13212,N_13622);
and U14064 (N_14064,N_13091,N_13470);
or U14065 (N_14065,N_13002,N_13474);
xnor U14066 (N_14066,N_13514,N_13087);
nand U14067 (N_14067,N_13610,N_13968);
xnor U14068 (N_14068,N_13788,N_13183);
nand U14069 (N_14069,N_13532,N_13810);
xor U14070 (N_14070,N_13969,N_13789);
and U14071 (N_14071,N_13688,N_13831);
and U14072 (N_14072,N_13485,N_13322);
xor U14073 (N_14073,N_13058,N_13929);
or U14074 (N_14074,N_13369,N_13658);
and U14075 (N_14075,N_13065,N_13463);
or U14076 (N_14076,N_13480,N_13338);
nor U14077 (N_14077,N_13068,N_13080);
xnor U14078 (N_14078,N_13483,N_13127);
and U14079 (N_14079,N_13282,N_13569);
nor U14080 (N_14080,N_13644,N_13876);
nand U14081 (N_14081,N_13452,N_13618);
xnor U14082 (N_14082,N_13045,N_13925);
nor U14083 (N_14083,N_13858,N_13601);
nand U14084 (N_14084,N_13550,N_13629);
nor U14085 (N_14085,N_13332,N_13027);
and U14086 (N_14086,N_13198,N_13039);
xnor U14087 (N_14087,N_13572,N_13881);
and U14088 (N_14088,N_13371,N_13641);
nor U14089 (N_14089,N_13067,N_13703);
or U14090 (N_14090,N_13599,N_13152);
nor U14091 (N_14091,N_13977,N_13098);
nor U14092 (N_14092,N_13797,N_13682);
and U14093 (N_14093,N_13317,N_13761);
nand U14094 (N_14094,N_13555,N_13501);
nand U14095 (N_14095,N_13185,N_13835);
nand U14096 (N_14096,N_13554,N_13128);
nand U14097 (N_14097,N_13795,N_13613);
nor U14098 (N_14098,N_13467,N_13998);
nor U14099 (N_14099,N_13587,N_13670);
or U14100 (N_14100,N_13010,N_13953);
or U14101 (N_14101,N_13230,N_13041);
and U14102 (N_14102,N_13216,N_13393);
nand U14103 (N_14103,N_13355,N_13135);
xnor U14104 (N_14104,N_13099,N_13110);
xnor U14105 (N_14105,N_13104,N_13144);
nand U14106 (N_14106,N_13241,N_13402);
and U14107 (N_14107,N_13581,N_13302);
or U14108 (N_14108,N_13879,N_13505);
nor U14109 (N_14109,N_13935,N_13081);
nor U14110 (N_14110,N_13739,N_13379);
nand U14111 (N_14111,N_13069,N_13121);
or U14112 (N_14112,N_13597,N_13033);
or U14113 (N_14113,N_13074,N_13571);
nor U14114 (N_14114,N_13698,N_13583);
or U14115 (N_14115,N_13763,N_13239);
xor U14116 (N_14116,N_13092,N_13286);
and U14117 (N_14117,N_13510,N_13667);
xor U14118 (N_14118,N_13029,N_13263);
xor U14119 (N_14119,N_13671,N_13856);
xnor U14120 (N_14120,N_13840,N_13708);
nor U14121 (N_14121,N_13460,N_13380);
nor U14122 (N_14122,N_13986,N_13639);
nand U14123 (N_14123,N_13478,N_13818);
or U14124 (N_14124,N_13391,N_13819);
and U14125 (N_14125,N_13129,N_13714);
nor U14126 (N_14126,N_13268,N_13751);
or U14127 (N_14127,N_13361,N_13026);
xor U14128 (N_14128,N_13414,N_13038);
and U14129 (N_14129,N_13251,N_13521);
or U14130 (N_14130,N_13036,N_13930);
nand U14131 (N_14131,N_13567,N_13533);
and U14132 (N_14132,N_13164,N_13535);
nor U14133 (N_14133,N_13204,N_13868);
xnor U14134 (N_14134,N_13907,N_13443);
nor U14135 (N_14135,N_13733,N_13617);
xnor U14136 (N_14136,N_13266,N_13035);
xnor U14137 (N_14137,N_13424,N_13063);
xnor U14138 (N_14138,N_13158,N_13209);
or U14139 (N_14139,N_13731,N_13250);
nand U14140 (N_14140,N_13412,N_13330);
nor U14141 (N_14141,N_13400,N_13342);
and U14142 (N_14142,N_13214,N_13738);
nor U14143 (N_14143,N_13323,N_13523);
or U14144 (N_14144,N_13918,N_13179);
or U14145 (N_14145,N_13832,N_13666);
nand U14146 (N_14146,N_13413,N_13562);
xor U14147 (N_14147,N_13839,N_13321);
nor U14148 (N_14148,N_13515,N_13882);
nor U14149 (N_14149,N_13927,N_13451);
and U14150 (N_14150,N_13457,N_13222);
xnor U14151 (N_14151,N_13199,N_13609);
nor U14152 (N_14152,N_13700,N_13362);
nor U14153 (N_14153,N_13624,N_13057);
or U14154 (N_14154,N_13574,N_13636);
nor U14155 (N_14155,N_13246,N_13097);
nor U14156 (N_14156,N_13590,N_13477);
or U14157 (N_14157,N_13249,N_13217);
nand U14158 (N_14158,N_13557,N_13125);
xnor U14159 (N_14159,N_13274,N_13425);
nor U14160 (N_14160,N_13952,N_13461);
xor U14161 (N_14161,N_13255,N_13181);
or U14162 (N_14162,N_13207,N_13180);
nor U14163 (N_14163,N_13909,N_13506);
xnor U14164 (N_14164,N_13724,N_13398);
xor U14165 (N_14165,N_13691,N_13748);
nor U14166 (N_14166,N_13253,N_13975);
xor U14167 (N_14167,N_13189,N_13407);
or U14168 (N_14168,N_13084,N_13101);
or U14169 (N_14169,N_13983,N_13933);
xor U14170 (N_14170,N_13861,N_13757);
or U14171 (N_14171,N_13034,N_13236);
and U14172 (N_14172,N_13006,N_13704);
xor U14173 (N_14173,N_13866,N_13867);
xor U14174 (N_14174,N_13392,N_13976);
and U14175 (N_14175,N_13416,N_13401);
nor U14176 (N_14176,N_13448,N_13928);
and U14177 (N_14177,N_13718,N_13306);
nor U14178 (N_14178,N_13494,N_13349);
or U14179 (N_14179,N_13820,N_13772);
xnor U14180 (N_14180,N_13887,N_13643);
or U14181 (N_14181,N_13359,N_13427);
or U14182 (N_14182,N_13540,N_13408);
and U14183 (N_14183,N_13758,N_13607);
xor U14184 (N_14184,N_13191,N_13133);
and U14185 (N_14185,N_13762,N_13019);
nor U14186 (N_14186,N_13974,N_13844);
nor U14187 (N_14187,N_13187,N_13148);
nand U14188 (N_14188,N_13260,N_13944);
or U14189 (N_14189,N_13114,N_13279);
and U14190 (N_14190,N_13075,N_13542);
nor U14191 (N_14191,N_13439,N_13271);
or U14192 (N_14192,N_13213,N_13806);
nor U14193 (N_14193,N_13942,N_13360);
or U14194 (N_14194,N_13211,N_13549);
nor U14195 (N_14195,N_13653,N_13365);
or U14196 (N_14196,N_13950,N_13728);
xor U14197 (N_14197,N_13220,N_13256);
or U14198 (N_14198,N_13706,N_13366);
nor U14199 (N_14199,N_13145,N_13801);
nor U14200 (N_14200,N_13674,N_13696);
and U14201 (N_14201,N_13812,N_13842);
nor U14202 (N_14202,N_13786,N_13377);
and U14203 (N_14203,N_13507,N_13247);
nor U14204 (N_14204,N_13082,N_13054);
xor U14205 (N_14205,N_13606,N_13774);
xnor U14206 (N_14206,N_13476,N_13358);
and U14207 (N_14207,N_13615,N_13556);
nor U14208 (N_14208,N_13740,N_13156);
or U14209 (N_14209,N_13775,N_13654);
xnor U14210 (N_14210,N_13710,N_13167);
or U14211 (N_14211,N_13875,N_13988);
and U14212 (N_14212,N_13194,N_13422);
nor U14213 (N_14213,N_13307,N_13223);
xor U14214 (N_14214,N_13699,N_13642);
nand U14215 (N_14215,N_13013,N_13771);
and U14216 (N_14216,N_13131,N_13971);
or U14217 (N_14217,N_13095,N_13059);
xor U14218 (N_14218,N_13536,N_13466);
or U14219 (N_14219,N_13309,N_13750);
xnor U14220 (N_14220,N_13999,N_13804);
or U14221 (N_14221,N_13853,N_13237);
and U14222 (N_14222,N_13531,N_13378);
nor U14223 (N_14223,N_13955,N_13090);
or U14224 (N_14224,N_13376,N_13972);
nor U14225 (N_14225,N_13356,N_13954);
xor U14226 (N_14226,N_13182,N_13721);
or U14227 (N_14227,N_13663,N_13770);
or U14228 (N_14228,N_13192,N_13206);
or U14229 (N_14229,N_13387,N_13421);
or U14230 (N_14230,N_13920,N_13348);
or U14231 (N_14231,N_13512,N_13298);
nand U14232 (N_14232,N_13031,N_13836);
xor U14233 (N_14233,N_13243,N_13530);
nor U14234 (N_14234,N_13650,N_13066);
nand U14235 (N_14235,N_13915,N_13585);
and U14236 (N_14236,N_13884,N_13007);
or U14237 (N_14237,N_13534,N_13300);
and U14238 (N_14238,N_13637,N_13056);
xnor U14239 (N_14239,N_13807,N_13735);
and U14240 (N_14240,N_13823,N_13508);
or U14241 (N_14241,N_13527,N_13697);
and U14242 (N_14242,N_13030,N_13525);
nor U14243 (N_14243,N_13280,N_13205);
nand U14244 (N_14244,N_13524,N_13516);
or U14245 (N_14245,N_13488,N_13811);
nand U14246 (N_14246,N_13747,N_13327);
or U14247 (N_14247,N_13903,N_13984);
or U14248 (N_14248,N_13326,N_13766);
nand U14249 (N_14249,N_13502,N_13108);
nor U14250 (N_14250,N_13612,N_13960);
xnor U14251 (N_14251,N_13614,N_13715);
and U14252 (N_14252,N_13454,N_13566);
nand U14253 (N_14253,N_13111,N_13105);
or U14254 (N_14254,N_13816,N_13655);
and U14255 (N_14255,N_13860,N_13712);
or U14256 (N_14256,N_13353,N_13292);
nor U14257 (N_14257,N_13498,N_13102);
and U14258 (N_14258,N_13817,N_13238);
nor U14259 (N_14259,N_13631,N_13956);
nand U14260 (N_14260,N_13345,N_13616);
xnor U14261 (N_14261,N_13992,N_13430);
nor U14262 (N_14262,N_13891,N_13720);
and U14263 (N_14263,N_13050,N_13173);
nand U14264 (N_14264,N_13689,N_13681);
nand U14265 (N_14265,N_13374,N_13796);
nor U14266 (N_14266,N_13814,N_13749);
and U14267 (N_14267,N_13278,N_13225);
nor U14268 (N_14268,N_13500,N_13295);
xor U14269 (N_14269,N_13620,N_13343);
xor U14270 (N_14270,N_13593,N_13004);
xor U14271 (N_14271,N_13822,N_13169);
nor U14272 (N_14272,N_13203,N_13850);
and U14273 (N_14273,N_13608,N_13197);
nor U14274 (N_14274,N_13305,N_13828);
nand U14275 (N_14275,N_13848,N_13503);
and U14276 (N_14276,N_13418,N_13910);
nor U14277 (N_14277,N_13964,N_13215);
or U14278 (N_14278,N_13634,N_13233);
xnor U14279 (N_14279,N_13603,N_13568);
nand U14280 (N_14280,N_13845,N_13446);
or U14281 (N_14281,N_13851,N_13665);
xnor U14282 (N_14282,N_13760,N_13134);
and U14283 (N_14283,N_13551,N_13318);
or U14284 (N_14284,N_13938,N_13472);
nor U14285 (N_14285,N_13445,N_13120);
and U14286 (N_14286,N_13224,N_13254);
nor U14287 (N_14287,N_13578,N_13573);
or U14288 (N_14288,N_13259,N_13790);
nor U14289 (N_14289,N_13570,N_13315);
nand U14290 (N_14290,N_13991,N_13464);
nor U14291 (N_14291,N_13827,N_13178);
or U14292 (N_14292,N_13395,N_13672);
xor U14293 (N_14293,N_13619,N_13547);
nor U14294 (N_14294,N_13023,N_13779);
nor U14295 (N_14295,N_13438,N_13742);
xor U14296 (N_14296,N_13025,N_13484);
nand U14297 (N_14297,N_13519,N_13686);
and U14298 (N_14298,N_13146,N_13898);
and U14299 (N_14299,N_13171,N_13219);
and U14300 (N_14300,N_13435,N_13890);
nand U14301 (N_14301,N_13112,N_13932);
nor U14302 (N_14302,N_13052,N_13662);
nand U14303 (N_14303,N_13061,N_13683);
and U14304 (N_14304,N_13440,N_13563);
or U14305 (N_14305,N_13768,N_13047);
xnor U14306 (N_14306,N_13518,N_13389);
or U14307 (N_14307,N_13635,N_13908);
or U14308 (N_14308,N_13001,N_13680);
nor U14309 (N_14309,N_13450,N_13911);
and U14310 (N_14310,N_13847,N_13668);
nand U14311 (N_14311,N_13626,N_13163);
or U14312 (N_14312,N_13623,N_13079);
and U14313 (N_14313,N_13577,N_13491);
nand U14314 (N_14314,N_13656,N_13647);
or U14315 (N_14315,N_13267,N_13154);
and U14316 (N_14316,N_13258,N_13885);
nand U14317 (N_14317,N_13877,N_13709);
xnor U14318 (N_14318,N_13015,N_13548);
nand U14319 (N_14319,N_13854,N_13793);
nor U14320 (N_14320,N_13429,N_13764);
nor U14321 (N_14321,N_13492,N_13100);
or U14322 (N_14322,N_13829,N_13982);
or U14323 (N_14323,N_13388,N_13544);
xor U14324 (N_14324,N_13741,N_13149);
or U14325 (N_14325,N_13895,N_13985);
nor U14326 (N_14326,N_13331,N_13396);
nor U14327 (N_14327,N_13917,N_13337);
and U14328 (N_14328,N_13611,N_13685);
xnor U14329 (N_14329,N_13073,N_13024);
nand U14330 (N_14330,N_13313,N_13946);
nand U14331 (N_14331,N_13329,N_13048);
nand U14332 (N_14332,N_13692,N_13705);
or U14333 (N_14333,N_13837,N_13973);
nor U14334 (N_14334,N_13826,N_13561);
or U14335 (N_14335,N_13902,N_13924);
nor U14336 (N_14336,N_13419,N_13176);
xnor U14337 (N_14337,N_13690,N_13479);
or U14338 (N_14338,N_13003,N_13072);
xnor U14339 (N_14339,N_13444,N_13730);
and U14340 (N_14340,N_13449,N_13897);
nor U14341 (N_14341,N_13743,N_13778);
xor U14342 (N_14342,N_13883,N_13273);
nor U14343 (N_14343,N_13528,N_13979);
nor U14344 (N_14344,N_13773,N_13904);
xor U14345 (N_14345,N_13888,N_13459);
nor U14346 (N_14346,N_13659,N_13341);
nand U14347 (N_14347,N_13874,N_13600);
or U14348 (N_14348,N_13384,N_13462);
or U14349 (N_14349,N_13399,N_13385);
and U14350 (N_14350,N_13299,N_13049);
nor U14351 (N_14351,N_13161,N_13892);
xor U14352 (N_14352,N_13310,N_13803);
or U14353 (N_14353,N_13147,N_13943);
and U14354 (N_14354,N_13621,N_13162);
nor U14355 (N_14355,N_13651,N_13783);
nor U14356 (N_14356,N_13014,N_13370);
nand U14357 (N_14357,N_13037,N_13736);
or U14358 (N_14358,N_13335,N_13423);
nor U14359 (N_14359,N_13405,N_13428);
nand U14360 (N_14360,N_13546,N_13453);
and U14361 (N_14361,N_13727,N_13234);
and U14362 (N_14362,N_13311,N_13021);
nand U14363 (N_14363,N_13046,N_13936);
and U14364 (N_14364,N_13325,N_13076);
xnor U14365 (N_14365,N_13678,N_13394);
nand U14366 (N_14366,N_13648,N_13308);
or U14367 (N_14367,N_13415,N_13752);
nor U14368 (N_14368,N_13228,N_13833);
nand U14369 (N_14369,N_13140,N_13070);
and U14370 (N_14370,N_13284,N_13262);
xnor U14371 (N_14371,N_13018,N_13071);
xor U14372 (N_14372,N_13130,N_13990);
nand U14373 (N_14373,N_13119,N_13713);
or U14374 (N_14374,N_13490,N_13123);
xor U14375 (N_14375,N_13290,N_13855);
or U14376 (N_14376,N_13722,N_13093);
or U14377 (N_14377,N_13945,N_13020);
or U14378 (N_14378,N_13304,N_13732);
nor U14379 (N_14379,N_13716,N_13410);
or U14380 (N_14380,N_13905,N_13717);
nor U14381 (N_14381,N_13113,N_13138);
and U14382 (N_14382,N_13602,N_13208);
xor U14383 (N_14383,N_13372,N_13289);
and U14384 (N_14384,N_13339,N_13809);
xor U14385 (N_14385,N_13168,N_13077);
and U14386 (N_14386,N_13124,N_13746);
nor U14387 (N_14387,N_13340,N_13261);
and U14388 (N_14388,N_13141,N_13575);
and U14389 (N_14389,N_13165,N_13558);
nand U14390 (N_14390,N_13381,N_13582);
nor U14391 (N_14391,N_13596,N_13800);
xnor U14392 (N_14392,N_13486,N_13878);
nor U14393 (N_14393,N_13687,N_13064);
and U14394 (N_14394,N_13580,N_13592);
nor U14395 (N_14395,N_13303,N_13588);
xnor U14396 (N_14396,N_13880,N_13155);
nand U14397 (N_14397,N_13137,N_13316);
nor U14398 (N_14398,N_13939,N_13638);
nor U14399 (N_14399,N_13351,N_13830);
or U14400 (N_14400,N_13940,N_13934);
nor U14401 (N_14401,N_13889,N_13011);
xnor U14402 (N_14402,N_13767,N_13863);
nand U14403 (N_14403,N_13184,N_13232);
or U14404 (N_14404,N_13106,N_13652);
nor U14405 (N_14405,N_13994,N_13997);
or U14406 (N_14406,N_13513,N_13948);
nor U14407 (N_14407,N_13677,N_13017);
and U14408 (N_14408,N_13734,N_13043);
and U14409 (N_14409,N_13702,N_13965);
nor U14410 (N_14410,N_13493,N_13022);
nor U14411 (N_14411,N_13283,N_13645);
or U14412 (N_14412,N_13725,N_13560);
nor U14413 (N_14413,N_13252,N_13364);
or U14414 (N_14414,N_13949,N_13009);
or U14415 (N_14415,N_13729,N_13765);
nor U14416 (N_14416,N_13669,N_13813);
nand U14417 (N_14417,N_13383,N_13537);
and U14418 (N_14418,N_13792,N_13333);
or U14419 (N_14419,N_13579,N_13871);
and U14420 (N_14420,N_13805,N_13170);
nand U14421 (N_14421,N_13143,N_13595);
nand U14422 (N_14422,N_13509,N_13336);
nand U14423 (N_14423,N_13872,N_13660);
or U14424 (N_14424,N_13139,N_13270);
or U14425 (N_14425,N_13684,N_13089);
nand U14426 (N_14426,N_13707,N_13862);
or U14427 (N_14427,N_13497,N_13469);
nand U14428 (N_14428,N_13324,N_13967);
nor U14429 (N_14429,N_13227,N_13921);
or U14430 (N_14430,N_13328,N_13417);
xnor U14431 (N_14431,N_13726,N_13980);
or U14432 (N_14432,N_13312,N_13923);
or U14433 (N_14433,N_13153,N_13970);
and U14434 (N_14434,N_13776,N_13754);
nor U14435 (N_14435,N_13711,N_13553);
and U14436 (N_14436,N_13798,N_13966);
or U14437 (N_14437,N_13288,N_13787);
nand U14438 (N_14438,N_13865,N_13657);
nand U14439 (N_14439,N_13995,N_13701);
or U14440 (N_14440,N_13426,N_13719);
xnor U14441 (N_14441,N_13334,N_13922);
or U14442 (N_14442,N_13352,N_13354);
xnor U14443 (N_14443,N_13802,N_13675);
xor U14444 (N_14444,N_13320,N_13314);
and U14445 (N_14445,N_13240,N_13541);
and U14446 (N_14446,N_13347,N_13744);
or U14447 (N_14447,N_13679,N_13777);
nor U14448 (N_14448,N_13150,N_13873);
xnor U14449 (N_14449,N_13489,N_13231);
or U14450 (N_14450,N_13769,N_13368);
nor U14451 (N_14451,N_13297,N_13051);
nand U14452 (N_14452,N_13916,N_13993);
and U14453 (N_14453,N_13265,N_13367);
or U14454 (N_14454,N_13436,N_13996);
nand U14455 (N_14455,N_13481,N_13411);
xnor U14456 (N_14456,N_13406,N_13088);
nand U14457 (N_14457,N_13640,N_13319);
xor U14458 (N_14458,N_13755,N_13160);
xor U14459 (N_14459,N_13218,N_13543);
xor U14460 (N_14460,N_13382,N_13409);
or U14461 (N_14461,N_13962,N_13941);
xor U14462 (N_14462,N_13664,N_13177);
nor U14463 (N_14463,N_13456,N_13195);
and U14464 (N_14464,N_13886,N_13815);
nand U14465 (N_14465,N_13799,N_13293);
nand U14466 (N_14466,N_13539,N_13632);
or U14467 (N_14467,N_13912,N_13078);
and U14468 (N_14468,N_13118,N_13248);
or U14469 (N_14469,N_13455,N_13576);
xor U14470 (N_14470,N_13285,N_13987);
xnor U14471 (N_14471,N_13390,N_13646);
xnor U14472 (N_14472,N_13468,N_13115);
or U14473 (N_14473,N_13522,N_13044);
or U14474 (N_14474,N_13864,N_13564);
nor U14475 (N_14475,N_13843,N_13893);
nand U14476 (N_14476,N_13545,N_13604);
or U14477 (N_14477,N_13028,N_13107);
xor U14478 (N_14478,N_13552,N_13958);
and U14479 (N_14479,N_13157,N_13458);
nand U14480 (N_14480,N_13852,N_13142);
xnor U14481 (N_14481,N_13487,N_13475);
and U14482 (N_14482,N_13870,N_13083);
nor U14483 (N_14483,N_13834,N_13200);
nor U14484 (N_14484,N_13062,N_13913);
or U14485 (N_14485,N_13403,N_13841);
xor U14486 (N_14486,N_13186,N_13136);
or U14487 (N_14487,N_13625,N_13126);
xor U14488 (N_14488,N_13808,N_13780);
nor U14489 (N_14489,N_13346,N_13756);
nand U14490 (N_14490,N_13434,N_13784);
or U14491 (N_14491,N_13737,N_13008);
or U14492 (N_14492,N_13745,N_13919);
xor U14493 (N_14493,N_13242,N_13291);
nor U14494 (N_14494,N_13344,N_13849);
or U14495 (N_14495,N_13926,N_13794);
nand U14496 (N_14496,N_13723,N_13520);
xnor U14497 (N_14497,N_13441,N_13482);
nand U14498 (N_14498,N_13210,N_13272);
nor U14499 (N_14499,N_13103,N_13175);
nand U14500 (N_14500,N_13535,N_13084);
nor U14501 (N_14501,N_13487,N_13583);
xor U14502 (N_14502,N_13721,N_13367);
and U14503 (N_14503,N_13822,N_13820);
and U14504 (N_14504,N_13391,N_13772);
and U14505 (N_14505,N_13083,N_13126);
xnor U14506 (N_14506,N_13012,N_13710);
nor U14507 (N_14507,N_13449,N_13338);
nor U14508 (N_14508,N_13465,N_13593);
xor U14509 (N_14509,N_13239,N_13122);
and U14510 (N_14510,N_13745,N_13679);
nand U14511 (N_14511,N_13888,N_13989);
xnor U14512 (N_14512,N_13669,N_13003);
and U14513 (N_14513,N_13489,N_13122);
nor U14514 (N_14514,N_13932,N_13533);
nor U14515 (N_14515,N_13491,N_13225);
nor U14516 (N_14516,N_13860,N_13763);
nand U14517 (N_14517,N_13341,N_13628);
and U14518 (N_14518,N_13099,N_13565);
nor U14519 (N_14519,N_13005,N_13213);
or U14520 (N_14520,N_13912,N_13399);
xnor U14521 (N_14521,N_13688,N_13702);
nand U14522 (N_14522,N_13637,N_13325);
xor U14523 (N_14523,N_13336,N_13256);
xor U14524 (N_14524,N_13443,N_13783);
or U14525 (N_14525,N_13796,N_13818);
and U14526 (N_14526,N_13813,N_13304);
or U14527 (N_14527,N_13924,N_13100);
or U14528 (N_14528,N_13448,N_13125);
nand U14529 (N_14529,N_13567,N_13554);
nor U14530 (N_14530,N_13740,N_13936);
nand U14531 (N_14531,N_13873,N_13529);
xor U14532 (N_14532,N_13690,N_13521);
or U14533 (N_14533,N_13855,N_13298);
nor U14534 (N_14534,N_13857,N_13838);
nand U14535 (N_14535,N_13320,N_13996);
or U14536 (N_14536,N_13379,N_13696);
and U14537 (N_14537,N_13989,N_13590);
or U14538 (N_14538,N_13594,N_13223);
or U14539 (N_14539,N_13387,N_13116);
nand U14540 (N_14540,N_13374,N_13451);
nand U14541 (N_14541,N_13672,N_13763);
or U14542 (N_14542,N_13488,N_13986);
nor U14543 (N_14543,N_13404,N_13402);
and U14544 (N_14544,N_13388,N_13271);
and U14545 (N_14545,N_13024,N_13276);
and U14546 (N_14546,N_13060,N_13772);
nand U14547 (N_14547,N_13871,N_13905);
nand U14548 (N_14548,N_13251,N_13983);
xnor U14549 (N_14549,N_13317,N_13720);
and U14550 (N_14550,N_13204,N_13655);
nor U14551 (N_14551,N_13342,N_13846);
and U14552 (N_14552,N_13091,N_13269);
or U14553 (N_14553,N_13826,N_13691);
and U14554 (N_14554,N_13217,N_13743);
xor U14555 (N_14555,N_13683,N_13021);
nand U14556 (N_14556,N_13805,N_13075);
xor U14557 (N_14557,N_13411,N_13560);
nand U14558 (N_14558,N_13022,N_13070);
xor U14559 (N_14559,N_13973,N_13495);
xnor U14560 (N_14560,N_13194,N_13885);
xnor U14561 (N_14561,N_13300,N_13082);
or U14562 (N_14562,N_13607,N_13823);
nand U14563 (N_14563,N_13718,N_13961);
xor U14564 (N_14564,N_13932,N_13977);
xnor U14565 (N_14565,N_13546,N_13979);
nor U14566 (N_14566,N_13879,N_13064);
and U14567 (N_14567,N_13154,N_13387);
or U14568 (N_14568,N_13413,N_13612);
or U14569 (N_14569,N_13781,N_13436);
or U14570 (N_14570,N_13081,N_13320);
nand U14571 (N_14571,N_13508,N_13329);
and U14572 (N_14572,N_13270,N_13932);
nand U14573 (N_14573,N_13592,N_13088);
and U14574 (N_14574,N_13024,N_13899);
or U14575 (N_14575,N_13445,N_13002);
or U14576 (N_14576,N_13438,N_13984);
or U14577 (N_14577,N_13348,N_13306);
xnor U14578 (N_14578,N_13198,N_13425);
and U14579 (N_14579,N_13158,N_13727);
nand U14580 (N_14580,N_13640,N_13423);
and U14581 (N_14581,N_13966,N_13665);
xor U14582 (N_14582,N_13684,N_13177);
and U14583 (N_14583,N_13616,N_13434);
nand U14584 (N_14584,N_13733,N_13156);
xor U14585 (N_14585,N_13680,N_13253);
xnor U14586 (N_14586,N_13722,N_13357);
and U14587 (N_14587,N_13985,N_13161);
and U14588 (N_14588,N_13536,N_13924);
nand U14589 (N_14589,N_13194,N_13894);
nand U14590 (N_14590,N_13165,N_13915);
and U14591 (N_14591,N_13313,N_13654);
or U14592 (N_14592,N_13067,N_13347);
and U14593 (N_14593,N_13110,N_13377);
nand U14594 (N_14594,N_13763,N_13587);
xor U14595 (N_14595,N_13668,N_13089);
and U14596 (N_14596,N_13061,N_13331);
xnor U14597 (N_14597,N_13992,N_13146);
nand U14598 (N_14598,N_13757,N_13462);
xor U14599 (N_14599,N_13096,N_13119);
nand U14600 (N_14600,N_13726,N_13702);
xor U14601 (N_14601,N_13221,N_13518);
and U14602 (N_14602,N_13955,N_13066);
xnor U14603 (N_14603,N_13433,N_13224);
and U14604 (N_14604,N_13251,N_13604);
or U14605 (N_14605,N_13983,N_13291);
nand U14606 (N_14606,N_13117,N_13444);
nor U14607 (N_14607,N_13896,N_13620);
xnor U14608 (N_14608,N_13302,N_13945);
and U14609 (N_14609,N_13660,N_13022);
or U14610 (N_14610,N_13695,N_13060);
and U14611 (N_14611,N_13483,N_13336);
or U14612 (N_14612,N_13055,N_13292);
nand U14613 (N_14613,N_13342,N_13535);
xnor U14614 (N_14614,N_13589,N_13789);
xor U14615 (N_14615,N_13855,N_13707);
and U14616 (N_14616,N_13323,N_13977);
xnor U14617 (N_14617,N_13735,N_13025);
and U14618 (N_14618,N_13603,N_13575);
nor U14619 (N_14619,N_13339,N_13905);
and U14620 (N_14620,N_13281,N_13182);
or U14621 (N_14621,N_13643,N_13591);
xnor U14622 (N_14622,N_13525,N_13385);
nand U14623 (N_14623,N_13201,N_13985);
or U14624 (N_14624,N_13186,N_13999);
nor U14625 (N_14625,N_13456,N_13582);
or U14626 (N_14626,N_13418,N_13759);
or U14627 (N_14627,N_13207,N_13587);
and U14628 (N_14628,N_13575,N_13531);
nor U14629 (N_14629,N_13952,N_13237);
xor U14630 (N_14630,N_13991,N_13598);
xor U14631 (N_14631,N_13048,N_13277);
nor U14632 (N_14632,N_13033,N_13959);
nand U14633 (N_14633,N_13969,N_13429);
xor U14634 (N_14634,N_13443,N_13851);
or U14635 (N_14635,N_13871,N_13660);
and U14636 (N_14636,N_13755,N_13492);
xor U14637 (N_14637,N_13674,N_13189);
nor U14638 (N_14638,N_13771,N_13958);
xor U14639 (N_14639,N_13377,N_13229);
nand U14640 (N_14640,N_13180,N_13873);
and U14641 (N_14641,N_13066,N_13022);
xor U14642 (N_14642,N_13841,N_13500);
xnor U14643 (N_14643,N_13972,N_13964);
nand U14644 (N_14644,N_13262,N_13398);
nand U14645 (N_14645,N_13991,N_13237);
and U14646 (N_14646,N_13083,N_13404);
nand U14647 (N_14647,N_13091,N_13590);
nand U14648 (N_14648,N_13987,N_13740);
or U14649 (N_14649,N_13360,N_13349);
nor U14650 (N_14650,N_13940,N_13425);
xor U14651 (N_14651,N_13726,N_13056);
nor U14652 (N_14652,N_13928,N_13549);
or U14653 (N_14653,N_13897,N_13580);
and U14654 (N_14654,N_13404,N_13483);
xor U14655 (N_14655,N_13092,N_13240);
or U14656 (N_14656,N_13920,N_13650);
xor U14657 (N_14657,N_13100,N_13137);
xnor U14658 (N_14658,N_13672,N_13373);
xnor U14659 (N_14659,N_13733,N_13357);
nor U14660 (N_14660,N_13444,N_13702);
nor U14661 (N_14661,N_13180,N_13480);
or U14662 (N_14662,N_13149,N_13580);
or U14663 (N_14663,N_13174,N_13823);
or U14664 (N_14664,N_13929,N_13054);
nand U14665 (N_14665,N_13917,N_13325);
nor U14666 (N_14666,N_13359,N_13311);
and U14667 (N_14667,N_13625,N_13755);
nand U14668 (N_14668,N_13799,N_13622);
xor U14669 (N_14669,N_13797,N_13937);
nand U14670 (N_14670,N_13388,N_13236);
xor U14671 (N_14671,N_13786,N_13484);
or U14672 (N_14672,N_13461,N_13829);
nor U14673 (N_14673,N_13061,N_13177);
xor U14674 (N_14674,N_13971,N_13179);
and U14675 (N_14675,N_13140,N_13183);
nand U14676 (N_14676,N_13903,N_13155);
or U14677 (N_14677,N_13048,N_13187);
or U14678 (N_14678,N_13154,N_13945);
and U14679 (N_14679,N_13764,N_13405);
xor U14680 (N_14680,N_13384,N_13953);
xnor U14681 (N_14681,N_13924,N_13465);
nor U14682 (N_14682,N_13551,N_13522);
nor U14683 (N_14683,N_13266,N_13205);
nand U14684 (N_14684,N_13490,N_13625);
or U14685 (N_14685,N_13500,N_13579);
nand U14686 (N_14686,N_13384,N_13758);
nand U14687 (N_14687,N_13523,N_13224);
nor U14688 (N_14688,N_13057,N_13159);
nand U14689 (N_14689,N_13196,N_13137);
nor U14690 (N_14690,N_13738,N_13725);
and U14691 (N_14691,N_13802,N_13138);
xnor U14692 (N_14692,N_13037,N_13973);
or U14693 (N_14693,N_13074,N_13902);
xnor U14694 (N_14694,N_13524,N_13321);
nand U14695 (N_14695,N_13839,N_13672);
or U14696 (N_14696,N_13053,N_13932);
nand U14697 (N_14697,N_13728,N_13183);
or U14698 (N_14698,N_13906,N_13639);
and U14699 (N_14699,N_13088,N_13838);
nor U14700 (N_14700,N_13660,N_13553);
and U14701 (N_14701,N_13834,N_13807);
or U14702 (N_14702,N_13379,N_13764);
nand U14703 (N_14703,N_13043,N_13074);
and U14704 (N_14704,N_13318,N_13458);
and U14705 (N_14705,N_13859,N_13000);
and U14706 (N_14706,N_13990,N_13327);
nor U14707 (N_14707,N_13216,N_13052);
nor U14708 (N_14708,N_13862,N_13095);
and U14709 (N_14709,N_13055,N_13338);
or U14710 (N_14710,N_13214,N_13132);
xnor U14711 (N_14711,N_13147,N_13176);
or U14712 (N_14712,N_13656,N_13129);
xor U14713 (N_14713,N_13536,N_13723);
nor U14714 (N_14714,N_13655,N_13375);
or U14715 (N_14715,N_13071,N_13597);
or U14716 (N_14716,N_13228,N_13400);
xor U14717 (N_14717,N_13141,N_13443);
or U14718 (N_14718,N_13238,N_13933);
and U14719 (N_14719,N_13113,N_13533);
nand U14720 (N_14720,N_13783,N_13744);
and U14721 (N_14721,N_13313,N_13757);
and U14722 (N_14722,N_13134,N_13831);
nor U14723 (N_14723,N_13322,N_13625);
and U14724 (N_14724,N_13498,N_13784);
nor U14725 (N_14725,N_13404,N_13825);
nand U14726 (N_14726,N_13761,N_13260);
xnor U14727 (N_14727,N_13540,N_13121);
or U14728 (N_14728,N_13684,N_13087);
nor U14729 (N_14729,N_13828,N_13910);
or U14730 (N_14730,N_13743,N_13139);
nor U14731 (N_14731,N_13426,N_13068);
and U14732 (N_14732,N_13542,N_13089);
or U14733 (N_14733,N_13273,N_13968);
nand U14734 (N_14734,N_13983,N_13739);
nand U14735 (N_14735,N_13863,N_13438);
xnor U14736 (N_14736,N_13520,N_13574);
xor U14737 (N_14737,N_13928,N_13345);
xor U14738 (N_14738,N_13680,N_13470);
nand U14739 (N_14739,N_13948,N_13635);
xor U14740 (N_14740,N_13155,N_13026);
or U14741 (N_14741,N_13914,N_13299);
and U14742 (N_14742,N_13688,N_13108);
or U14743 (N_14743,N_13056,N_13666);
xnor U14744 (N_14744,N_13881,N_13366);
or U14745 (N_14745,N_13977,N_13618);
xor U14746 (N_14746,N_13457,N_13381);
nor U14747 (N_14747,N_13774,N_13423);
nand U14748 (N_14748,N_13022,N_13646);
nor U14749 (N_14749,N_13715,N_13450);
nand U14750 (N_14750,N_13270,N_13817);
and U14751 (N_14751,N_13579,N_13167);
nand U14752 (N_14752,N_13412,N_13842);
nand U14753 (N_14753,N_13872,N_13766);
nor U14754 (N_14754,N_13551,N_13785);
and U14755 (N_14755,N_13059,N_13753);
and U14756 (N_14756,N_13258,N_13714);
or U14757 (N_14757,N_13336,N_13700);
nand U14758 (N_14758,N_13617,N_13952);
xor U14759 (N_14759,N_13247,N_13846);
nor U14760 (N_14760,N_13797,N_13502);
nor U14761 (N_14761,N_13403,N_13077);
nand U14762 (N_14762,N_13945,N_13798);
nand U14763 (N_14763,N_13066,N_13427);
xnor U14764 (N_14764,N_13257,N_13618);
nor U14765 (N_14765,N_13923,N_13782);
and U14766 (N_14766,N_13238,N_13267);
nand U14767 (N_14767,N_13697,N_13009);
nand U14768 (N_14768,N_13157,N_13207);
xnor U14769 (N_14769,N_13608,N_13322);
or U14770 (N_14770,N_13217,N_13459);
xor U14771 (N_14771,N_13171,N_13144);
xnor U14772 (N_14772,N_13108,N_13748);
nand U14773 (N_14773,N_13659,N_13795);
xnor U14774 (N_14774,N_13568,N_13725);
nor U14775 (N_14775,N_13250,N_13884);
nor U14776 (N_14776,N_13671,N_13021);
xor U14777 (N_14777,N_13619,N_13676);
nor U14778 (N_14778,N_13695,N_13488);
xor U14779 (N_14779,N_13289,N_13023);
nor U14780 (N_14780,N_13594,N_13158);
nor U14781 (N_14781,N_13728,N_13032);
xor U14782 (N_14782,N_13570,N_13916);
xnor U14783 (N_14783,N_13607,N_13228);
and U14784 (N_14784,N_13777,N_13477);
and U14785 (N_14785,N_13000,N_13952);
xor U14786 (N_14786,N_13809,N_13195);
and U14787 (N_14787,N_13089,N_13605);
nand U14788 (N_14788,N_13607,N_13437);
nand U14789 (N_14789,N_13058,N_13951);
nor U14790 (N_14790,N_13830,N_13511);
nor U14791 (N_14791,N_13984,N_13584);
nor U14792 (N_14792,N_13738,N_13580);
or U14793 (N_14793,N_13407,N_13901);
nand U14794 (N_14794,N_13406,N_13839);
or U14795 (N_14795,N_13880,N_13048);
xnor U14796 (N_14796,N_13302,N_13757);
and U14797 (N_14797,N_13866,N_13288);
or U14798 (N_14798,N_13635,N_13967);
nor U14799 (N_14799,N_13434,N_13624);
nor U14800 (N_14800,N_13845,N_13689);
xor U14801 (N_14801,N_13776,N_13689);
nor U14802 (N_14802,N_13272,N_13610);
xor U14803 (N_14803,N_13188,N_13537);
nand U14804 (N_14804,N_13371,N_13056);
xnor U14805 (N_14805,N_13410,N_13292);
xor U14806 (N_14806,N_13755,N_13490);
nand U14807 (N_14807,N_13556,N_13048);
or U14808 (N_14808,N_13543,N_13794);
nor U14809 (N_14809,N_13767,N_13012);
nor U14810 (N_14810,N_13068,N_13479);
nand U14811 (N_14811,N_13147,N_13572);
xnor U14812 (N_14812,N_13729,N_13380);
and U14813 (N_14813,N_13655,N_13299);
or U14814 (N_14814,N_13574,N_13307);
nor U14815 (N_14815,N_13183,N_13048);
nor U14816 (N_14816,N_13245,N_13958);
xor U14817 (N_14817,N_13254,N_13813);
or U14818 (N_14818,N_13298,N_13661);
nor U14819 (N_14819,N_13455,N_13306);
nand U14820 (N_14820,N_13303,N_13402);
and U14821 (N_14821,N_13958,N_13691);
nor U14822 (N_14822,N_13182,N_13383);
nor U14823 (N_14823,N_13128,N_13550);
or U14824 (N_14824,N_13473,N_13293);
or U14825 (N_14825,N_13167,N_13227);
and U14826 (N_14826,N_13845,N_13386);
or U14827 (N_14827,N_13867,N_13687);
and U14828 (N_14828,N_13262,N_13533);
nor U14829 (N_14829,N_13528,N_13379);
nand U14830 (N_14830,N_13308,N_13351);
or U14831 (N_14831,N_13721,N_13273);
nor U14832 (N_14832,N_13494,N_13893);
and U14833 (N_14833,N_13176,N_13388);
and U14834 (N_14834,N_13973,N_13741);
nor U14835 (N_14835,N_13404,N_13166);
xnor U14836 (N_14836,N_13851,N_13878);
nand U14837 (N_14837,N_13869,N_13705);
nand U14838 (N_14838,N_13122,N_13115);
nand U14839 (N_14839,N_13751,N_13096);
and U14840 (N_14840,N_13887,N_13349);
nor U14841 (N_14841,N_13838,N_13636);
or U14842 (N_14842,N_13872,N_13979);
and U14843 (N_14843,N_13779,N_13052);
nor U14844 (N_14844,N_13412,N_13408);
or U14845 (N_14845,N_13681,N_13637);
xor U14846 (N_14846,N_13159,N_13860);
nor U14847 (N_14847,N_13203,N_13935);
or U14848 (N_14848,N_13765,N_13016);
or U14849 (N_14849,N_13880,N_13060);
and U14850 (N_14850,N_13413,N_13185);
nor U14851 (N_14851,N_13931,N_13679);
or U14852 (N_14852,N_13441,N_13011);
nor U14853 (N_14853,N_13426,N_13439);
nand U14854 (N_14854,N_13818,N_13877);
nor U14855 (N_14855,N_13896,N_13374);
or U14856 (N_14856,N_13280,N_13265);
nand U14857 (N_14857,N_13993,N_13934);
or U14858 (N_14858,N_13343,N_13258);
nand U14859 (N_14859,N_13246,N_13606);
xor U14860 (N_14860,N_13464,N_13866);
nor U14861 (N_14861,N_13672,N_13357);
nand U14862 (N_14862,N_13950,N_13135);
xnor U14863 (N_14863,N_13298,N_13588);
nand U14864 (N_14864,N_13260,N_13482);
nand U14865 (N_14865,N_13645,N_13589);
or U14866 (N_14866,N_13135,N_13019);
xor U14867 (N_14867,N_13255,N_13538);
xor U14868 (N_14868,N_13092,N_13728);
xor U14869 (N_14869,N_13977,N_13519);
xor U14870 (N_14870,N_13995,N_13504);
xnor U14871 (N_14871,N_13332,N_13495);
nand U14872 (N_14872,N_13607,N_13162);
xor U14873 (N_14873,N_13262,N_13832);
xnor U14874 (N_14874,N_13823,N_13771);
nand U14875 (N_14875,N_13269,N_13113);
and U14876 (N_14876,N_13791,N_13705);
and U14877 (N_14877,N_13415,N_13903);
and U14878 (N_14878,N_13451,N_13615);
xor U14879 (N_14879,N_13520,N_13104);
and U14880 (N_14880,N_13382,N_13042);
and U14881 (N_14881,N_13931,N_13746);
xor U14882 (N_14882,N_13358,N_13669);
or U14883 (N_14883,N_13026,N_13315);
nor U14884 (N_14884,N_13064,N_13371);
nor U14885 (N_14885,N_13411,N_13629);
or U14886 (N_14886,N_13478,N_13483);
or U14887 (N_14887,N_13668,N_13716);
xnor U14888 (N_14888,N_13189,N_13997);
nand U14889 (N_14889,N_13750,N_13131);
nor U14890 (N_14890,N_13395,N_13625);
xnor U14891 (N_14891,N_13385,N_13962);
xor U14892 (N_14892,N_13541,N_13131);
and U14893 (N_14893,N_13840,N_13307);
and U14894 (N_14894,N_13110,N_13518);
nand U14895 (N_14895,N_13594,N_13744);
nand U14896 (N_14896,N_13988,N_13456);
xnor U14897 (N_14897,N_13894,N_13206);
xor U14898 (N_14898,N_13093,N_13183);
and U14899 (N_14899,N_13868,N_13399);
nor U14900 (N_14900,N_13128,N_13041);
nand U14901 (N_14901,N_13359,N_13840);
or U14902 (N_14902,N_13532,N_13668);
and U14903 (N_14903,N_13672,N_13090);
xor U14904 (N_14904,N_13298,N_13687);
nand U14905 (N_14905,N_13317,N_13067);
or U14906 (N_14906,N_13465,N_13699);
nand U14907 (N_14907,N_13713,N_13164);
and U14908 (N_14908,N_13193,N_13551);
xnor U14909 (N_14909,N_13365,N_13282);
or U14910 (N_14910,N_13178,N_13251);
and U14911 (N_14911,N_13353,N_13885);
xnor U14912 (N_14912,N_13371,N_13817);
nand U14913 (N_14913,N_13428,N_13827);
xor U14914 (N_14914,N_13496,N_13859);
nand U14915 (N_14915,N_13441,N_13487);
or U14916 (N_14916,N_13611,N_13816);
or U14917 (N_14917,N_13314,N_13433);
nor U14918 (N_14918,N_13523,N_13039);
xnor U14919 (N_14919,N_13179,N_13821);
or U14920 (N_14920,N_13229,N_13747);
or U14921 (N_14921,N_13520,N_13597);
xor U14922 (N_14922,N_13980,N_13648);
xnor U14923 (N_14923,N_13408,N_13469);
and U14924 (N_14924,N_13824,N_13295);
and U14925 (N_14925,N_13872,N_13963);
nor U14926 (N_14926,N_13412,N_13240);
and U14927 (N_14927,N_13276,N_13517);
nand U14928 (N_14928,N_13677,N_13460);
or U14929 (N_14929,N_13504,N_13821);
or U14930 (N_14930,N_13602,N_13253);
or U14931 (N_14931,N_13888,N_13284);
and U14932 (N_14932,N_13663,N_13189);
nor U14933 (N_14933,N_13311,N_13061);
xnor U14934 (N_14934,N_13811,N_13050);
xor U14935 (N_14935,N_13018,N_13721);
nand U14936 (N_14936,N_13830,N_13212);
and U14937 (N_14937,N_13447,N_13024);
nand U14938 (N_14938,N_13958,N_13932);
nand U14939 (N_14939,N_13135,N_13207);
or U14940 (N_14940,N_13809,N_13949);
nand U14941 (N_14941,N_13796,N_13096);
xor U14942 (N_14942,N_13090,N_13255);
xor U14943 (N_14943,N_13695,N_13388);
or U14944 (N_14944,N_13680,N_13554);
xnor U14945 (N_14945,N_13800,N_13092);
nand U14946 (N_14946,N_13203,N_13832);
nand U14947 (N_14947,N_13984,N_13694);
or U14948 (N_14948,N_13986,N_13225);
nor U14949 (N_14949,N_13434,N_13642);
or U14950 (N_14950,N_13344,N_13821);
nand U14951 (N_14951,N_13527,N_13613);
or U14952 (N_14952,N_13772,N_13116);
xnor U14953 (N_14953,N_13878,N_13536);
xnor U14954 (N_14954,N_13881,N_13154);
or U14955 (N_14955,N_13925,N_13064);
xor U14956 (N_14956,N_13627,N_13970);
and U14957 (N_14957,N_13180,N_13087);
nand U14958 (N_14958,N_13378,N_13404);
nand U14959 (N_14959,N_13496,N_13541);
xor U14960 (N_14960,N_13510,N_13312);
xor U14961 (N_14961,N_13621,N_13159);
xor U14962 (N_14962,N_13882,N_13430);
nor U14963 (N_14963,N_13483,N_13879);
nor U14964 (N_14964,N_13653,N_13994);
nor U14965 (N_14965,N_13153,N_13030);
nand U14966 (N_14966,N_13515,N_13181);
or U14967 (N_14967,N_13737,N_13974);
xor U14968 (N_14968,N_13100,N_13409);
xnor U14969 (N_14969,N_13184,N_13611);
or U14970 (N_14970,N_13543,N_13564);
nand U14971 (N_14971,N_13040,N_13823);
or U14972 (N_14972,N_13944,N_13347);
nand U14973 (N_14973,N_13755,N_13880);
and U14974 (N_14974,N_13886,N_13428);
nor U14975 (N_14975,N_13288,N_13849);
and U14976 (N_14976,N_13678,N_13151);
xnor U14977 (N_14977,N_13658,N_13059);
or U14978 (N_14978,N_13605,N_13579);
nor U14979 (N_14979,N_13851,N_13413);
nand U14980 (N_14980,N_13450,N_13271);
and U14981 (N_14981,N_13371,N_13382);
xor U14982 (N_14982,N_13502,N_13770);
xor U14983 (N_14983,N_13751,N_13072);
or U14984 (N_14984,N_13678,N_13931);
and U14985 (N_14985,N_13446,N_13176);
or U14986 (N_14986,N_13306,N_13072);
or U14987 (N_14987,N_13426,N_13484);
xnor U14988 (N_14988,N_13452,N_13577);
or U14989 (N_14989,N_13267,N_13743);
nor U14990 (N_14990,N_13819,N_13390);
nand U14991 (N_14991,N_13817,N_13062);
nand U14992 (N_14992,N_13980,N_13243);
or U14993 (N_14993,N_13166,N_13227);
nor U14994 (N_14994,N_13360,N_13561);
nand U14995 (N_14995,N_13531,N_13044);
and U14996 (N_14996,N_13485,N_13859);
nor U14997 (N_14997,N_13593,N_13921);
nand U14998 (N_14998,N_13258,N_13106);
nor U14999 (N_14999,N_13651,N_13085);
or UO_0 (O_0,N_14801,N_14153);
and UO_1 (O_1,N_14635,N_14857);
and UO_2 (O_2,N_14957,N_14575);
or UO_3 (O_3,N_14713,N_14441);
and UO_4 (O_4,N_14506,N_14346);
nor UO_5 (O_5,N_14901,N_14401);
xor UO_6 (O_6,N_14837,N_14912);
or UO_7 (O_7,N_14526,N_14974);
and UO_8 (O_8,N_14085,N_14019);
xor UO_9 (O_9,N_14330,N_14774);
nor UO_10 (O_10,N_14318,N_14761);
nand UO_11 (O_11,N_14354,N_14934);
nor UO_12 (O_12,N_14914,N_14012);
nand UO_13 (O_13,N_14237,N_14843);
nor UO_14 (O_14,N_14953,N_14543);
nor UO_15 (O_15,N_14663,N_14715);
nor UO_16 (O_16,N_14223,N_14764);
or UO_17 (O_17,N_14336,N_14870);
and UO_18 (O_18,N_14042,N_14721);
nand UO_19 (O_19,N_14396,N_14786);
xor UO_20 (O_20,N_14779,N_14530);
nand UO_21 (O_21,N_14355,N_14768);
and UO_22 (O_22,N_14325,N_14694);
and UO_23 (O_23,N_14995,N_14275);
xnor UO_24 (O_24,N_14752,N_14625);
nor UO_25 (O_25,N_14736,N_14051);
nand UO_26 (O_26,N_14047,N_14645);
or UO_27 (O_27,N_14861,N_14831);
xnor UO_28 (O_28,N_14028,N_14658);
nor UO_29 (O_29,N_14821,N_14281);
or UO_30 (O_30,N_14608,N_14502);
nor UO_31 (O_31,N_14911,N_14812);
xor UO_32 (O_32,N_14586,N_14046);
or UO_33 (O_33,N_14943,N_14392);
or UO_34 (O_34,N_14202,N_14698);
nor UO_35 (O_35,N_14522,N_14574);
nor UO_36 (O_36,N_14660,N_14924);
xor UO_37 (O_37,N_14039,N_14100);
nand UO_38 (O_38,N_14387,N_14717);
and UO_39 (O_39,N_14689,N_14650);
nor UO_40 (O_40,N_14862,N_14619);
and UO_41 (O_41,N_14015,N_14675);
and UO_42 (O_42,N_14427,N_14554);
xor UO_43 (O_43,N_14632,N_14144);
xor UO_44 (O_44,N_14101,N_14602);
and UO_45 (O_45,N_14013,N_14527);
nor UO_46 (O_46,N_14380,N_14002);
and UO_47 (O_47,N_14403,N_14139);
nor UO_48 (O_48,N_14183,N_14755);
or UO_49 (O_49,N_14127,N_14391);
nand UO_50 (O_50,N_14769,N_14804);
and UO_51 (O_51,N_14517,N_14647);
and UO_52 (O_52,N_14307,N_14657);
xor UO_53 (O_53,N_14900,N_14731);
and UO_54 (O_54,N_14984,N_14618);
or UO_55 (O_55,N_14567,N_14165);
nand UO_56 (O_56,N_14573,N_14890);
nor UO_57 (O_57,N_14309,N_14669);
nand UO_58 (O_58,N_14808,N_14927);
xnor UO_59 (O_59,N_14584,N_14010);
nand UO_60 (O_60,N_14347,N_14320);
or UO_61 (O_61,N_14117,N_14803);
nand UO_62 (O_62,N_14269,N_14218);
xnor UO_63 (O_63,N_14132,N_14609);
nor UO_64 (O_64,N_14031,N_14288);
xnor UO_65 (O_65,N_14313,N_14692);
or UO_66 (O_66,N_14216,N_14162);
or UO_67 (O_67,N_14287,N_14140);
nand UO_68 (O_68,N_14003,N_14653);
nand UO_69 (O_69,N_14533,N_14091);
nand UO_70 (O_70,N_14185,N_14671);
and UO_71 (O_71,N_14148,N_14365);
nor UO_72 (O_72,N_14025,N_14300);
xnor UO_73 (O_73,N_14680,N_14245);
nand UO_74 (O_74,N_14756,N_14276);
and UO_75 (O_75,N_14058,N_14503);
nor UO_76 (O_76,N_14899,N_14741);
or UO_77 (O_77,N_14036,N_14295);
or UO_78 (O_78,N_14151,N_14119);
nor UO_79 (O_79,N_14024,N_14122);
nor UO_80 (O_80,N_14604,N_14367);
nand UO_81 (O_81,N_14997,N_14677);
or UO_82 (O_82,N_14941,N_14027);
and UO_83 (O_83,N_14490,N_14023);
and UO_84 (O_84,N_14585,N_14145);
xor UO_85 (O_85,N_14215,N_14963);
or UO_86 (O_86,N_14572,N_14563);
and UO_87 (O_87,N_14676,N_14809);
xnor UO_88 (O_88,N_14435,N_14932);
xor UO_89 (O_89,N_14737,N_14534);
and UO_90 (O_90,N_14322,N_14846);
or UO_91 (O_91,N_14884,N_14780);
nand UO_92 (O_92,N_14279,N_14931);
xor UO_93 (O_93,N_14558,N_14221);
nand UO_94 (O_94,N_14952,N_14964);
nor UO_95 (O_95,N_14610,N_14478);
nor UO_96 (O_96,N_14935,N_14008);
xor UO_97 (O_97,N_14455,N_14087);
nor UO_98 (O_98,N_14795,N_14777);
nand UO_99 (O_99,N_14179,N_14277);
nor UO_100 (O_100,N_14972,N_14486);
nand UO_101 (O_101,N_14836,N_14507);
xor UO_102 (O_102,N_14589,N_14746);
nor UO_103 (O_103,N_14516,N_14826);
xor UO_104 (O_104,N_14246,N_14535);
nor UO_105 (O_105,N_14848,N_14686);
or UO_106 (O_106,N_14434,N_14461);
nor UO_107 (O_107,N_14508,N_14829);
nand UO_108 (O_108,N_14975,N_14753);
or UO_109 (O_109,N_14967,N_14334);
nand UO_110 (O_110,N_14099,N_14171);
nor UO_111 (O_111,N_14767,N_14001);
nor UO_112 (O_112,N_14086,N_14388);
nor UO_113 (O_113,N_14893,N_14284);
or UO_114 (O_114,N_14587,N_14670);
xnor UO_115 (O_115,N_14298,N_14371);
xor UO_116 (O_116,N_14882,N_14342);
or UO_117 (O_117,N_14407,N_14173);
nand UO_118 (O_118,N_14982,N_14249);
nand UO_119 (O_119,N_14550,N_14552);
nor UO_120 (O_120,N_14946,N_14523);
or UO_121 (O_121,N_14070,N_14176);
xor UO_122 (O_122,N_14885,N_14131);
or UO_123 (O_123,N_14521,N_14059);
xnor UO_124 (O_124,N_14564,N_14851);
or UO_125 (O_125,N_14049,N_14847);
or UO_126 (O_126,N_14339,N_14240);
xor UO_127 (O_127,N_14887,N_14638);
xnor UO_128 (O_128,N_14005,N_14592);
nor UO_129 (O_129,N_14348,N_14103);
nor UO_130 (O_130,N_14524,N_14616);
or UO_131 (O_131,N_14942,N_14199);
and UO_132 (O_132,N_14303,N_14655);
nand UO_133 (O_133,N_14599,N_14370);
xnor UO_134 (O_134,N_14238,N_14703);
or UO_135 (O_135,N_14394,N_14372);
xnor UO_136 (O_136,N_14965,N_14278);
and UO_137 (O_137,N_14282,N_14204);
nand UO_138 (O_138,N_14440,N_14109);
and UO_139 (O_139,N_14125,N_14557);
xnor UO_140 (O_140,N_14302,N_14673);
xnor UO_141 (O_141,N_14004,N_14402);
xnor UO_142 (O_142,N_14160,N_14494);
and UO_143 (O_143,N_14709,N_14954);
nor UO_144 (O_144,N_14580,N_14636);
or UO_145 (O_145,N_14405,N_14878);
and UO_146 (O_146,N_14877,N_14695);
and UO_147 (O_147,N_14323,N_14227);
nor UO_148 (O_148,N_14343,N_14710);
and UO_149 (O_149,N_14359,N_14189);
nor UO_150 (O_150,N_14373,N_14922);
and UO_151 (O_151,N_14327,N_14470);
nand UO_152 (O_152,N_14788,N_14850);
nand UO_153 (O_153,N_14771,N_14286);
or UO_154 (O_154,N_14224,N_14789);
and UO_155 (O_155,N_14576,N_14785);
or UO_156 (O_156,N_14633,N_14228);
and UO_157 (O_157,N_14696,N_14193);
or UO_158 (O_158,N_14773,N_14560);
or UO_159 (O_159,N_14067,N_14232);
nand UO_160 (O_160,N_14697,N_14351);
and UO_161 (O_161,N_14460,N_14089);
xnor UO_162 (O_162,N_14467,N_14271);
nand UO_163 (O_163,N_14649,N_14104);
nand UO_164 (O_164,N_14601,N_14577);
and UO_165 (O_165,N_14852,N_14541);
or UO_166 (O_166,N_14422,N_14652);
and UO_167 (O_167,N_14762,N_14272);
and UO_168 (O_168,N_14823,N_14389);
nand UO_169 (O_169,N_14687,N_14090);
and UO_170 (O_170,N_14404,N_14811);
and UO_171 (O_171,N_14433,N_14398);
and UO_172 (O_172,N_14429,N_14439);
nand UO_173 (O_173,N_14518,N_14376);
or UO_174 (O_174,N_14681,N_14725);
and UO_175 (O_175,N_14462,N_14138);
nor UO_176 (O_176,N_14594,N_14234);
nand UO_177 (O_177,N_14629,N_14688);
and UO_178 (O_178,N_14068,N_14274);
or UO_179 (O_179,N_14740,N_14763);
xnor UO_180 (O_180,N_14949,N_14532);
or UO_181 (O_181,N_14191,N_14711);
nand UO_182 (O_182,N_14385,N_14312);
or UO_183 (O_183,N_14037,N_14600);
nand UO_184 (O_184,N_14329,N_14416);
or UO_185 (O_185,N_14446,N_14464);
xor UO_186 (O_186,N_14048,N_14016);
or UO_187 (O_187,N_14095,N_14748);
xnor UO_188 (O_188,N_14944,N_14744);
and UO_189 (O_189,N_14475,N_14822);
nand UO_190 (O_190,N_14981,N_14590);
and UO_191 (O_191,N_14693,N_14168);
xor UO_192 (O_192,N_14854,N_14743);
or UO_193 (O_193,N_14319,N_14116);
nor UO_194 (O_194,N_14468,N_14834);
xnor UO_195 (O_195,N_14570,N_14268);
xnor UO_196 (O_196,N_14783,N_14026);
xnor UO_197 (O_197,N_14181,N_14393);
or UO_198 (O_198,N_14328,N_14993);
or UO_199 (O_199,N_14615,N_14933);
or UO_200 (O_200,N_14583,N_14666);
and UO_201 (O_201,N_14641,N_14332);
nand UO_202 (O_202,N_14712,N_14369);
nand UO_203 (O_203,N_14340,N_14252);
xnor UO_204 (O_204,N_14180,N_14169);
or UO_205 (O_205,N_14936,N_14961);
nor UO_206 (O_206,N_14888,N_14793);
nor UO_207 (O_207,N_14297,N_14050);
nor UO_208 (O_208,N_14661,N_14726);
nor UO_209 (O_209,N_14654,N_14990);
nor UO_210 (O_210,N_14118,N_14172);
nand UO_211 (O_211,N_14137,N_14408);
nor UO_212 (O_212,N_14844,N_14057);
xnor UO_213 (O_213,N_14529,N_14738);
nor UO_214 (O_214,N_14285,N_14679);
xor UO_215 (O_215,N_14722,N_14948);
xnor UO_216 (O_216,N_14161,N_14871);
xnor UO_217 (O_217,N_14352,N_14620);
and UO_218 (O_218,N_14656,N_14891);
xor UO_219 (O_219,N_14668,N_14383);
nor UO_220 (O_220,N_14951,N_14164);
xnor UO_221 (O_221,N_14452,N_14420);
nand UO_222 (O_222,N_14859,N_14971);
or UO_223 (O_223,N_14500,N_14749);
nand UO_224 (O_224,N_14923,N_14582);
or UO_225 (O_225,N_14634,N_14730);
nand UO_226 (O_226,N_14056,N_14849);
or UO_227 (O_227,N_14958,N_14614);
nor UO_228 (O_228,N_14106,N_14643);
or UO_229 (O_229,N_14869,N_14874);
nor UO_230 (O_230,N_14640,N_14747);
and UO_231 (O_231,N_14471,N_14515);
and UO_232 (O_232,N_14399,N_14919);
nand UO_233 (O_233,N_14233,N_14421);
and UO_234 (O_234,N_14044,N_14627);
or UO_235 (O_235,N_14551,N_14561);
nand UO_236 (O_236,N_14504,N_14400);
xor UO_237 (O_237,N_14338,N_14546);
or UO_238 (O_238,N_14136,N_14497);
xor UO_239 (O_239,N_14112,N_14978);
nor UO_240 (O_240,N_14644,N_14501);
nor UO_241 (O_241,N_14624,N_14706);
or UO_242 (O_242,N_14187,N_14966);
and UO_243 (O_243,N_14538,N_14875);
and UO_244 (O_244,N_14157,N_14092);
nor UO_245 (O_245,N_14622,N_14236);
nor UO_246 (O_246,N_14796,N_14714);
nor UO_247 (O_247,N_14315,N_14438);
nand UO_248 (O_248,N_14220,N_14815);
or UO_249 (O_249,N_14553,N_14222);
nor UO_250 (O_250,N_14472,N_14835);
xor UO_251 (O_251,N_14055,N_14321);
nor UO_252 (O_252,N_14838,N_14775);
nor UO_253 (O_253,N_14628,N_14491);
or UO_254 (O_254,N_14253,N_14256);
nand UO_255 (O_255,N_14902,N_14559);
or UO_256 (O_256,N_14977,N_14007);
nand UO_257 (O_257,N_14895,N_14667);
nand UO_258 (O_258,N_14682,N_14121);
xor UO_259 (O_259,N_14214,N_14390);
nor UO_260 (O_260,N_14908,N_14998);
and UO_261 (O_261,N_14243,N_14913);
xnor UO_262 (O_262,N_14152,N_14631);
nand UO_263 (O_263,N_14781,N_14605);
and UO_264 (O_264,N_14805,N_14291);
and UO_265 (O_265,N_14498,N_14356);
nand UO_266 (O_266,N_14979,N_14606);
or UO_267 (O_267,N_14537,N_14239);
and UO_268 (O_268,N_14444,N_14866);
and UO_269 (O_269,N_14562,N_14474);
xnor UO_270 (O_270,N_14797,N_14203);
xor UO_271 (O_271,N_14487,N_14456);
and UO_272 (O_272,N_14581,N_14445);
xor UO_273 (O_273,N_14150,N_14034);
nand UO_274 (O_274,N_14443,N_14833);
nor UO_275 (O_275,N_14428,N_14178);
or UO_276 (O_276,N_14873,N_14579);
xor UO_277 (O_277,N_14415,N_14915);
and UO_278 (O_278,N_14333,N_14230);
and UO_279 (O_279,N_14244,N_14108);
and UO_280 (O_280,N_14410,N_14156);
or UO_281 (O_281,N_14344,N_14229);
nor UO_282 (O_282,N_14045,N_14386);
nand UO_283 (O_283,N_14702,N_14621);
xor UO_284 (O_284,N_14910,N_14685);
nand UO_285 (O_285,N_14817,N_14200);
and UO_286 (O_286,N_14166,N_14845);
xnor UO_287 (O_287,N_14480,N_14928);
or UO_288 (O_288,N_14375,N_14970);
nor UO_289 (O_289,N_14335,N_14197);
or UO_290 (O_290,N_14513,N_14798);
and UO_291 (O_291,N_14409,N_14906);
xnor UO_292 (O_292,N_14299,N_14742);
nand UO_293 (O_293,N_14810,N_14465);
or UO_294 (O_294,N_14863,N_14029);
or UO_295 (O_295,N_14384,N_14613);
and UO_296 (O_296,N_14603,N_14192);
or UO_297 (O_297,N_14417,N_14947);
nand UO_298 (O_298,N_14664,N_14186);
nand UO_299 (O_299,N_14489,N_14626);
or UO_300 (O_300,N_14937,N_14700);
nor UO_301 (O_301,N_14418,N_14270);
xor UO_302 (O_302,N_14038,N_14081);
nor UO_303 (O_303,N_14310,N_14041);
nand UO_304 (O_304,N_14733,N_14473);
or UO_305 (O_305,N_14110,N_14976);
or UO_306 (O_306,N_14426,N_14907);
xor UO_307 (O_307,N_14280,N_14242);
xor UO_308 (O_308,N_14536,N_14651);
nand UO_309 (O_309,N_14053,N_14930);
and UO_310 (O_310,N_14163,N_14219);
xor UO_311 (O_311,N_14720,N_14133);
nand UO_312 (O_312,N_14377,N_14481);
nor UO_313 (O_313,N_14510,N_14814);
or UO_314 (O_314,N_14894,N_14305);
nor UO_315 (O_315,N_14991,N_14531);
or UO_316 (O_316,N_14107,N_14544);
nor UO_317 (O_317,N_14672,N_14458);
and UO_318 (O_318,N_14141,N_14381);
xor UO_319 (O_319,N_14378,N_14565);
nor UO_320 (O_320,N_14453,N_14985);
nor UO_321 (O_321,N_14262,N_14765);
nand UO_322 (O_322,N_14331,N_14751);
xor UO_323 (O_323,N_14612,N_14018);
or UO_324 (O_324,N_14938,N_14987);
or UO_325 (O_325,N_14147,N_14159);
nand UO_326 (O_326,N_14595,N_14827);
nor UO_327 (O_327,N_14959,N_14754);
and UO_328 (O_328,N_14520,N_14030);
nor UO_329 (O_329,N_14469,N_14425);
and UO_330 (O_330,N_14054,N_14512);
nor UO_331 (O_331,N_14729,N_14674);
or UO_332 (O_332,N_14865,N_14593);
or UO_333 (O_333,N_14032,N_14542);
nor UO_334 (O_334,N_14155,N_14892);
or UO_335 (O_335,N_14799,N_14898);
xor UO_336 (O_336,N_14170,N_14555);
nand UO_337 (O_337,N_14828,N_14258);
nand UO_338 (O_338,N_14263,N_14662);
and UO_339 (O_339,N_14918,N_14842);
and UO_340 (O_340,N_14317,N_14397);
xnor UO_341 (O_341,N_14926,N_14855);
xor UO_342 (O_342,N_14492,N_14813);
or UO_343 (O_343,N_14825,N_14363);
xor UO_344 (O_344,N_14424,N_14146);
nor UO_345 (O_345,N_14250,N_14301);
nor UO_346 (O_346,N_14881,N_14167);
and UO_347 (O_347,N_14868,N_14361);
and UO_348 (O_348,N_14353,N_14254);
xnor UO_349 (O_349,N_14648,N_14128);
xnor UO_350 (O_350,N_14800,N_14360);
and UO_351 (O_351,N_14925,N_14547);
or UO_352 (O_352,N_14872,N_14097);
nand UO_353 (O_353,N_14758,N_14776);
and UO_354 (O_354,N_14265,N_14337);
nand UO_355 (O_355,N_14566,N_14980);
and UO_356 (O_356,N_14569,N_14113);
xnor UO_357 (O_357,N_14052,N_14528);
nand UO_358 (O_358,N_14296,N_14072);
nor UO_359 (O_359,N_14525,N_14430);
or UO_360 (O_360,N_14886,N_14973);
or UO_361 (O_361,N_14787,N_14314);
and UO_362 (O_362,N_14450,N_14904);
xor UO_363 (O_363,N_14940,N_14519);
xnor UO_364 (O_364,N_14665,N_14316);
and UO_365 (O_365,N_14956,N_14174);
nor UO_366 (O_366,N_14637,N_14540);
xnor UO_367 (O_367,N_14611,N_14734);
and UO_368 (O_368,N_14723,N_14009);
or UO_369 (O_369,N_14324,N_14630);
xor UO_370 (O_370,N_14304,N_14206);
or UO_371 (O_371,N_14929,N_14488);
nor UO_372 (O_372,N_14207,N_14366);
xor UO_373 (O_373,N_14950,N_14905);
or UO_374 (O_374,N_14718,N_14719);
nand UO_375 (O_375,N_14006,N_14463);
nand UO_376 (O_376,N_14413,N_14080);
xor UO_377 (O_377,N_14077,N_14063);
nand UO_378 (O_378,N_14597,N_14511);
nand UO_379 (O_379,N_14556,N_14545);
nand UO_380 (O_380,N_14194,N_14466);
and UO_381 (O_381,N_14791,N_14437);
nor UO_382 (O_382,N_14123,N_14824);
or UO_383 (O_383,N_14225,N_14096);
nand UO_384 (O_384,N_14772,N_14917);
xnor UO_385 (O_385,N_14382,N_14114);
nand UO_386 (O_386,N_14061,N_14617);
and UO_387 (O_387,N_14790,N_14289);
xnor UO_388 (O_388,N_14701,N_14205);
nand UO_389 (O_389,N_14105,N_14739);
nand UO_390 (O_390,N_14832,N_14920);
or UO_391 (O_391,N_14707,N_14839);
or UO_392 (O_392,N_14442,N_14406);
nand UO_393 (O_393,N_14955,N_14358);
xnor UO_394 (O_394,N_14476,N_14345);
nand UO_395 (O_395,N_14142,N_14724);
nor UO_396 (O_396,N_14094,N_14248);
or UO_397 (O_397,N_14571,N_14000);
nor UO_398 (O_398,N_14646,N_14357);
or UO_399 (O_399,N_14195,N_14853);
and UO_400 (O_400,N_14578,N_14479);
or UO_401 (O_401,N_14454,N_14182);
nor UO_402 (O_402,N_14022,N_14130);
or UO_403 (O_403,N_14308,N_14945);
xor UO_404 (O_404,N_14678,N_14499);
or UO_405 (O_405,N_14414,N_14259);
or UO_406 (O_406,N_14154,N_14266);
or UO_407 (O_407,N_14992,N_14766);
nor UO_408 (O_408,N_14184,N_14436);
or UO_409 (O_409,N_14782,N_14568);
nor UO_410 (O_410,N_14889,N_14257);
xor UO_411 (O_411,N_14423,N_14379);
nand UO_412 (O_412,N_14264,N_14075);
xnor UO_413 (O_413,N_14903,N_14960);
or UO_414 (O_414,N_14759,N_14120);
and UO_415 (O_415,N_14292,N_14778);
xor UO_416 (O_416,N_14261,N_14989);
and UO_417 (O_417,N_14231,N_14124);
or UO_418 (O_418,N_14419,N_14149);
and UO_419 (O_419,N_14395,N_14750);
and UO_420 (O_420,N_14447,N_14212);
xnor UO_421 (O_421,N_14247,N_14642);
nor UO_422 (O_422,N_14806,N_14830);
and UO_423 (O_423,N_14065,N_14607);
nand UO_424 (O_424,N_14098,N_14111);
xor UO_425 (O_425,N_14209,N_14457);
and UO_426 (O_426,N_14014,N_14691);
nand UO_427 (O_427,N_14040,N_14374);
xnor UO_428 (O_428,N_14158,N_14073);
nor UO_429 (O_429,N_14349,N_14760);
or UO_430 (O_430,N_14708,N_14598);
nand UO_431 (O_431,N_14482,N_14876);
and UO_432 (O_432,N_14011,N_14062);
nor UO_433 (O_433,N_14735,N_14596);
or UO_434 (O_434,N_14076,N_14083);
nor UO_435 (O_435,N_14818,N_14794);
and UO_436 (O_436,N_14273,N_14241);
or UO_437 (O_437,N_14188,N_14745);
xor UO_438 (O_438,N_14326,N_14177);
and UO_439 (O_439,N_14290,N_14448);
and UO_440 (O_440,N_14548,N_14549);
nand UO_441 (O_441,N_14088,N_14411);
xor UO_442 (O_442,N_14260,N_14883);
nor UO_443 (O_443,N_14858,N_14477);
nor UO_444 (O_444,N_14115,N_14896);
xor UO_445 (O_445,N_14770,N_14210);
nand UO_446 (O_446,N_14432,N_14867);
xor UO_447 (O_447,N_14784,N_14968);
and UO_448 (O_448,N_14840,N_14539);
or UO_449 (O_449,N_14939,N_14306);
nand UO_450 (O_450,N_14451,N_14060);
or UO_451 (O_451,N_14017,N_14683);
nor UO_452 (O_452,N_14064,N_14716);
or UO_453 (O_453,N_14364,N_14082);
xnor UO_454 (O_454,N_14921,N_14485);
xnor UO_455 (O_455,N_14879,N_14659);
nand UO_456 (O_456,N_14493,N_14093);
nor UO_457 (O_457,N_14213,N_14591);
nand UO_458 (O_458,N_14728,N_14020);
or UO_459 (O_459,N_14514,N_14690);
and UO_460 (O_460,N_14033,N_14988);
and UO_461 (O_461,N_14459,N_14996);
nor UO_462 (O_462,N_14079,N_14819);
or UO_463 (O_463,N_14283,N_14757);
or UO_464 (O_464,N_14196,N_14293);
nor UO_465 (O_465,N_14484,N_14129);
nand UO_466 (O_466,N_14208,N_14368);
nand UO_467 (O_467,N_14986,N_14126);
nand UO_468 (O_468,N_14135,N_14880);
nor UO_469 (O_469,N_14198,N_14134);
nor UO_470 (O_470,N_14431,N_14732);
xor UO_471 (O_471,N_14175,N_14916);
and UO_472 (O_472,N_14069,N_14509);
xor UO_473 (O_473,N_14699,N_14983);
or UO_474 (O_474,N_14897,N_14909);
nand UO_475 (O_475,N_14727,N_14496);
or UO_476 (O_476,N_14860,N_14705);
xnor UO_477 (O_477,N_14802,N_14341);
or UO_478 (O_478,N_14820,N_14999);
nor UO_479 (O_479,N_14792,N_14807);
nor UO_480 (O_480,N_14035,N_14864);
and UO_481 (O_481,N_14201,N_14994);
and UO_482 (O_482,N_14211,N_14969);
and UO_483 (O_483,N_14226,N_14684);
xor UO_484 (O_484,N_14505,N_14495);
nand UO_485 (O_485,N_14704,N_14066);
nor UO_486 (O_486,N_14255,N_14235);
nand UO_487 (O_487,N_14362,N_14071);
and UO_488 (O_488,N_14084,N_14143);
and UO_489 (O_489,N_14841,N_14074);
or UO_490 (O_490,N_14816,N_14078);
xor UO_491 (O_491,N_14311,N_14294);
xnor UO_492 (O_492,N_14190,N_14483);
nand UO_493 (O_493,N_14623,N_14267);
nor UO_494 (O_494,N_14350,N_14043);
or UO_495 (O_495,N_14449,N_14639);
nor UO_496 (O_496,N_14856,N_14251);
nor UO_497 (O_497,N_14412,N_14217);
nand UO_498 (O_498,N_14588,N_14102);
and UO_499 (O_499,N_14021,N_14962);
xor UO_500 (O_500,N_14103,N_14938);
nor UO_501 (O_501,N_14840,N_14941);
or UO_502 (O_502,N_14348,N_14429);
and UO_503 (O_503,N_14909,N_14165);
nor UO_504 (O_504,N_14792,N_14553);
nor UO_505 (O_505,N_14744,N_14571);
xor UO_506 (O_506,N_14940,N_14926);
nor UO_507 (O_507,N_14463,N_14262);
xnor UO_508 (O_508,N_14139,N_14028);
nor UO_509 (O_509,N_14664,N_14144);
and UO_510 (O_510,N_14622,N_14367);
and UO_511 (O_511,N_14329,N_14737);
nor UO_512 (O_512,N_14058,N_14961);
and UO_513 (O_513,N_14404,N_14891);
xnor UO_514 (O_514,N_14382,N_14123);
nor UO_515 (O_515,N_14024,N_14272);
xor UO_516 (O_516,N_14708,N_14845);
xnor UO_517 (O_517,N_14411,N_14405);
xnor UO_518 (O_518,N_14834,N_14252);
nand UO_519 (O_519,N_14226,N_14549);
xor UO_520 (O_520,N_14967,N_14199);
or UO_521 (O_521,N_14468,N_14295);
or UO_522 (O_522,N_14005,N_14172);
nor UO_523 (O_523,N_14322,N_14521);
and UO_524 (O_524,N_14532,N_14491);
nor UO_525 (O_525,N_14317,N_14309);
or UO_526 (O_526,N_14377,N_14058);
or UO_527 (O_527,N_14036,N_14133);
nor UO_528 (O_528,N_14751,N_14087);
nor UO_529 (O_529,N_14656,N_14715);
nor UO_530 (O_530,N_14329,N_14991);
nor UO_531 (O_531,N_14570,N_14751);
nand UO_532 (O_532,N_14273,N_14527);
or UO_533 (O_533,N_14855,N_14133);
nor UO_534 (O_534,N_14614,N_14574);
xor UO_535 (O_535,N_14282,N_14087);
nand UO_536 (O_536,N_14820,N_14956);
nor UO_537 (O_537,N_14469,N_14170);
nand UO_538 (O_538,N_14790,N_14925);
or UO_539 (O_539,N_14690,N_14081);
xnor UO_540 (O_540,N_14059,N_14410);
xnor UO_541 (O_541,N_14060,N_14368);
and UO_542 (O_542,N_14853,N_14998);
xnor UO_543 (O_543,N_14836,N_14742);
xnor UO_544 (O_544,N_14191,N_14863);
nor UO_545 (O_545,N_14856,N_14753);
nand UO_546 (O_546,N_14937,N_14527);
xnor UO_547 (O_547,N_14128,N_14051);
nand UO_548 (O_548,N_14639,N_14128);
xor UO_549 (O_549,N_14429,N_14656);
and UO_550 (O_550,N_14041,N_14568);
xnor UO_551 (O_551,N_14186,N_14380);
nor UO_552 (O_552,N_14574,N_14676);
or UO_553 (O_553,N_14037,N_14198);
nor UO_554 (O_554,N_14233,N_14109);
and UO_555 (O_555,N_14723,N_14669);
xor UO_556 (O_556,N_14474,N_14053);
nand UO_557 (O_557,N_14362,N_14631);
and UO_558 (O_558,N_14136,N_14158);
nand UO_559 (O_559,N_14085,N_14230);
and UO_560 (O_560,N_14668,N_14789);
nand UO_561 (O_561,N_14481,N_14830);
nand UO_562 (O_562,N_14576,N_14524);
or UO_563 (O_563,N_14661,N_14650);
xor UO_564 (O_564,N_14291,N_14173);
nor UO_565 (O_565,N_14006,N_14000);
nand UO_566 (O_566,N_14275,N_14951);
nand UO_567 (O_567,N_14361,N_14376);
xor UO_568 (O_568,N_14224,N_14321);
nor UO_569 (O_569,N_14310,N_14123);
xnor UO_570 (O_570,N_14872,N_14379);
nand UO_571 (O_571,N_14727,N_14583);
nor UO_572 (O_572,N_14129,N_14131);
nor UO_573 (O_573,N_14197,N_14807);
nor UO_574 (O_574,N_14509,N_14520);
and UO_575 (O_575,N_14802,N_14994);
and UO_576 (O_576,N_14017,N_14332);
and UO_577 (O_577,N_14051,N_14104);
nor UO_578 (O_578,N_14495,N_14950);
xor UO_579 (O_579,N_14176,N_14656);
nand UO_580 (O_580,N_14640,N_14698);
or UO_581 (O_581,N_14567,N_14752);
xnor UO_582 (O_582,N_14349,N_14258);
nor UO_583 (O_583,N_14078,N_14858);
nand UO_584 (O_584,N_14456,N_14781);
and UO_585 (O_585,N_14697,N_14861);
xnor UO_586 (O_586,N_14621,N_14458);
nor UO_587 (O_587,N_14778,N_14207);
xor UO_588 (O_588,N_14752,N_14689);
and UO_589 (O_589,N_14158,N_14176);
and UO_590 (O_590,N_14282,N_14837);
and UO_591 (O_591,N_14985,N_14122);
or UO_592 (O_592,N_14325,N_14431);
nor UO_593 (O_593,N_14520,N_14230);
and UO_594 (O_594,N_14882,N_14716);
or UO_595 (O_595,N_14165,N_14182);
xor UO_596 (O_596,N_14109,N_14611);
nor UO_597 (O_597,N_14757,N_14013);
nor UO_598 (O_598,N_14573,N_14343);
or UO_599 (O_599,N_14094,N_14327);
xnor UO_600 (O_600,N_14377,N_14620);
nand UO_601 (O_601,N_14875,N_14404);
or UO_602 (O_602,N_14780,N_14537);
nor UO_603 (O_603,N_14692,N_14564);
nand UO_604 (O_604,N_14417,N_14569);
or UO_605 (O_605,N_14240,N_14145);
or UO_606 (O_606,N_14493,N_14345);
xor UO_607 (O_607,N_14699,N_14373);
and UO_608 (O_608,N_14064,N_14080);
nor UO_609 (O_609,N_14655,N_14984);
nand UO_610 (O_610,N_14184,N_14433);
and UO_611 (O_611,N_14036,N_14517);
nor UO_612 (O_612,N_14040,N_14593);
or UO_613 (O_613,N_14333,N_14092);
or UO_614 (O_614,N_14015,N_14169);
nor UO_615 (O_615,N_14407,N_14830);
or UO_616 (O_616,N_14559,N_14143);
and UO_617 (O_617,N_14730,N_14221);
or UO_618 (O_618,N_14443,N_14858);
xnor UO_619 (O_619,N_14165,N_14687);
and UO_620 (O_620,N_14461,N_14776);
and UO_621 (O_621,N_14983,N_14590);
or UO_622 (O_622,N_14041,N_14624);
or UO_623 (O_623,N_14426,N_14918);
nand UO_624 (O_624,N_14783,N_14954);
and UO_625 (O_625,N_14113,N_14508);
nor UO_626 (O_626,N_14351,N_14703);
xnor UO_627 (O_627,N_14058,N_14356);
nand UO_628 (O_628,N_14024,N_14462);
nor UO_629 (O_629,N_14261,N_14772);
xnor UO_630 (O_630,N_14605,N_14945);
xor UO_631 (O_631,N_14735,N_14378);
or UO_632 (O_632,N_14348,N_14290);
or UO_633 (O_633,N_14029,N_14779);
and UO_634 (O_634,N_14888,N_14186);
and UO_635 (O_635,N_14131,N_14648);
or UO_636 (O_636,N_14567,N_14461);
or UO_637 (O_637,N_14581,N_14011);
xnor UO_638 (O_638,N_14824,N_14334);
nor UO_639 (O_639,N_14468,N_14904);
xnor UO_640 (O_640,N_14081,N_14128);
or UO_641 (O_641,N_14710,N_14344);
nand UO_642 (O_642,N_14918,N_14412);
nor UO_643 (O_643,N_14684,N_14390);
nor UO_644 (O_644,N_14044,N_14441);
or UO_645 (O_645,N_14016,N_14698);
nand UO_646 (O_646,N_14197,N_14581);
or UO_647 (O_647,N_14576,N_14801);
nand UO_648 (O_648,N_14526,N_14183);
nor UO_649 (O_649,N_14282,N_14255);
nand UO_650 (O_650,N_14362,N_14496);
or UO_651 (O_651,N_14973,N_14141);
nor UO_652 (O_652,N_14189,N_14074);
or UO_653 (O_653,N_14735,N_14062);
xor UO_654 (O_654,N_14203,N_14750);
and UO_655 (O_655,N_14769,N_14144);
and UO_656 (O_656,N_14539,N_14083);
xor UO_657 (O_657,N_14090,N_14706);
and UO_658 (O_658,N_14740,N_14989);
nand UO_659 (O_659,N_14769,N_14297);
and UO_660 (O_660,N_14025,N_14346);
xnor UO_661 (O_661,N_14482,N_14642);
nand UO_662 (O_662,N_14393,N_14862);
xnor UO_663 (O_663,N_14814,N_14775);
and UO_664 (O_664,N_14225,N_14752);
nand UO_665 (O_665,N_14489,N_14388);
or UO_666 (O_666,N_14165,N_14593);
nor UO_667 (O_667,N_14068,N_14958);
nor UO_668 (O_668,N_14776,N_14443);
nand UO_669 (O_669,N_14761,N_14885);
and UO_670 (O_670,N_14260,N_14045);
or UO_671 (O_671,N_14314,N_14041);
nand UO_672 (O_672,N_14593,N_14630);
and UO_673 (O_673,N_14252,N_14085);
nand UO_674 (O_674,N_14241,N_14187);
nor UO_675 (O_675,N_14228,N_14187);
and UO_676 (O_676,N_14413,N_14933);
or UO_677 (O_677,N_14002,N_14051);
and UO_678 (O_678,N_14984,N_14788);
nor UO_679 (O_679,N_14755,N_14274);
or UO_680 (O_680,N_14202,N_14337);
xor UO_681 (O_681,N_14696,N_14620);
xor UO_682 (O_682,N_14617,N_14908);
or UO_683 (O_683,N_14031,N_14713);
or UO_684 (O_684,N_14064,N_14876);
or UO_685 (O_685,N_14972,N_14322);
or UO_686 (O_686,N_14305,N_14057);
nor UO_687 (O_687,N_14426,N_14625);
and UO_688 (O_688,N_14169,N_14824);
nor UO_689 (O_689,N_14922,N_14187);
nand UO_690 (O_690,N_14097,N_14403);
and UO_691 (O_691,N_14905,N_14290);
or UO_692 (O_692,N_14410,N_14200);
nand UO_693 (O_693,N_14055,N_14713);
nor UO_694 (O_694,N_14316,N_14367);
nand UO_695 (O_695,N_14018,N_14435);
xor UO_696 (O_696,N_14804,N_14530);
and UO_697 (O_697,N_14997,N_14695);
nor UO_698 (O_698,N_14347,N_14511);
or UO_699 (O_699,N_14921,N_14019);
or UO_700 (O_700,N_14301,N_14731);
xnor UO_701 (O_701,N_14558,N_14706);
and UO_702 (O_702,N_14901,N_14045);
and UO_703 (O_703,N_14274,N_14809);
nand UO_704 (O_704,N_14193,N_14135);
and UO_705 (O_705,N_14732,N_14825);
and UO_706 (O_706,N_14620,N_14968);
xnor UO_707 (O_707,N_14479,N_14541);
nand UO_708 (O_708,N_14123,N_14687);
xnor UO_709 (O_709,N_14464,N_14486);
nand UO_710 (O_710,N_14899,N_14487);
and UO_711 (O_711,N_14460,N_14216);
nor UO_712 (O_712,N_14473,N_14041);
or UO_713 (O_713,N_14163,N_14846);
nand UO_714 (O_714,N_14056,N_14431);
xnor UO_715 (O_715,N_14689,N_14157);
nor UO_716 (O_716,N_14411,N_14658);
or UO_717 (O_717,N_14174,N_14830);
or UO_718 (O_718,N_14382,N_14921);
xnor UO_719 (O_719,N_14175,N_14639);
xor UO_720 (O_720,N_14271,N_14273);
nand UO_721 (O_721,N_14425,N_14848);
or UO_722 (O_722,N_14240,N_14336);
xor UO_723 (O_723,N_14972,N_14243);
nor UO_724 (O_724,N_14191,N_14008);
nand UO_725 (O_725,N_14992,N_14119);
xor UO_726 (O_726,N_14783,N_14670);
xor UO_727 (O_727,N_14060,N_14895);
or UO_728 (O_728,N_14988,N_14288);
or UO_729 (O_729,N_14167,N_14527);
nor UO_730 (O_730,N_14404,N_14577);
nand UO_731 (O_731,N_14755,N_14146);
nand UO_732 (O_732,N_14518,N_14147);
and UO_733 (O_733,N_14062,N_14766);
or UO_734 (O_734,N_14282,N_14706);
and UO_735 (O_735,N_14086,N_14658);
and UO_736 (O_736,N_14927,N_14233);
nand UO_737 (O_737,N_14425,N_14696);
or UO_738 (O_738,N_14674,N_14093);
nand UO_739 (O_739,N_14745,N_14896);
and UO_740 (O_740,N_14273,N_14755);
and UO_741 (O_741,N_14078,N_14483);
and UO_742 (O_742,N_14888,N_14536);
xor UO_743 (O_743,N_14937,N_14211);
or UO_744 (O_744,N_14916,N_14102);
xnor UO_745 (O_745,N_14505,N_14086);
xnor UO_746 (O_746,N_14787,N_14559);
and UO_747 (O_747,N_14510,N_14697);
xnor UO_748 (O_748,N_14387,N_14865);
or UO_749 (O_749,N_14515,N_14943);
nor UO_750 (O_750,N_14567,N_14761);
nor UO_751 (O_751,N_14402,N_14204);
nor UO_752 (O_752,N_14920,N_14815);
or UO_753 (O_753,N_14022,N_14412);
xor UO_754 (O_754,N_14719,N_14709);
nor UO_755 (O_755,N_14930,N_14455);
or UO_756 (O_756,N_14538,N_14320);
or UO_757 (O_757,N_14176,N_14035);
nand UO_758 (O_758,N_14511,N_14081);
nor UO_759 (O_759,N_14855,N_14436);
or UO_760 (O_760,N_14641,N_14534);
nand UO_761 (O_761,N_14963,N_14312);
xor UO_762 (O_762,N_14572,N_14644);
nand UO_763 (O_763,N_14665,N_14453);
xor UO_764 (O_764,N_14818,N_14326);
nor UO_765 (O_765,N_14831,N_14615);
nor UO_766 (O_766,N_14806,N_14116);
nand UO_767 (O_767,N_14739,N_14124);
and UO_768 (O_768,N_14636,N_14434);
xor UO_769 (O_769,N_14641,N_14158);
or UO_770 (O_770,N_14346,N_14071);
nand UO_771 (O_771,N_14319,N_14573);
or UO_772 (O_772,N_14114,N_14386);
and UO_773 (O_773,N_14947,N_14582);
nand UO_774 (O_774,N_14037,N_14338);
and UO_775 (O_775,N_14554,N_14968);
and UO_776 (O_776,N_14956,N_14451);
nor UO_777 (O_777,N_14987,N_14720);
xor UO_778 (O_778,N_14803,N_14394);
nor UO_779 (O_779,N_14573,N_14193);
or UO_780 (O_780,N_14831,N_14927);
xor UO_781 (O_781,N_14955,N_14824);
and UO_782 (O_782,N_14994,N_14967);
nor UO_783 (O_783,N_14881,N_14898);
and UO_784 (O_784,N_14984,N_14594);
and UO_785 (O_785,N_14268,N_14799);
or UO_786 (O_786,N_14311,N_14354);
nand UO_787 (O_787,N_14640,N_14285);
nand UO_788 (O_788,N_14715,N_14044);
and UO_789 (O_789,N_14680,N_14852);
nand UO_790 (O_790,N_14735,N_14416);
and UO_791 (O_791,N_14990,N_14543);
xor UO_792 (O_792,N_14516,N_14879);
nor UO_793 (O_793,N_14608,N_14450);
nor UO_794 (O_794,N_14618,N_14932);
and UO_795 (O_795,N_14317,N_14819);
xnor UO_796 (O_796,N_14811,N_14009);
nand UO_797 (O_797,N_14977,N_14883);
nor UO_798 (O_798,N_14905,N_14812);
and UO_799 (O_799,N_14769,N_14865);
and UO_800 (O_800,N_14128,N_14359);
xnor UO_801 (O_801,N_14732,N_14601);
and UO_802 (O_802,N_14477,N_14423);
or UO_803 (O_803,N_14811,N_14148);
or UO_804 (O_804,N_14443,N_14003);
or UO_805 (O_805,N_14239,N_14018);
and UO_806 (O_806,N_14328,N_14592);
nor UO_807 (O_807,N_14415,N_14424);
nand UO_808 (O_808,N_14192,N_14076);
xnor UO_809 (O_809,N_14557,N_14725);
nand UO_810 (O_810,N_14651,N_14521);
and UO_811 (O_811,N_14514,N_14195);
nor UO_812 (O_812,N_14590,N_14149);
xnor UO_813 (O_813,N_14102,N_14618);
and UO_814 (O_814,N_14596,N_14729);
nand UO_815 (O_815,N_14969,N_14045);
xor UO_816 (O_816,N_14345,N_14149);
nor UO_817 (O_817,N_14144,N_14581);
nand UO_818 (O_818,N_14838,N_14780);
or UO_819 (O_819,N_14231,N_14799);
and UO_820 (O_820,N_14046,N_14920);
or UO_821 (O_821,N_14770,N_14735);
nand UO_822 (O_822,N_14806,N_14296);
and UO_823 (O_823,N_14962,N_14773);
nand UO_824 (O_824,N_14834,N_14321);
or UO_825 (O_825,N_14374,N_14701);
or UO_826 (O_826,N_14900,N_14274);
xnor UO_827 (O_827,N_14388,N_14060);
or UO_828 (O_828,N_14388,N_14168);
nand UO_829 (O_829,N_14333,N_14275);
nor UO_830 (O_830,N_14784,N_14534);
or UO_831 (O_831,N_14209,N_14158);
xnor UO_832 (O_832,N_14506,N_14980);
nor UO_833 (O_833,N_14774,N_14481);
xor UO_834 (O_834,N_14681,N_14809);
xnor UO_835 (O_835,N_14405,N_14351);
or UO_836 (O_836,N_14634,N_14108);
nor UO_837 (O_837,N_14313,N_14278);
nor UO_838 (O_838,N_14192,N_14522);
nand UO_839 (O_839,N_14482,N_14945);
nand UO_840 (O_840,N_14607,N_14293);
nor UO_841 (O_841,N_14944,N_14937);
and UO_842 (O_842,N_14255,N_14995);
and UO_843 (O_843,N_14731,N_14961);
or UO_844 (O_844,N_14674,N_14323);
nand UO_845 (O_845,N_14976,N_14586);
xnor UO_846 (O_846,N_14088,N_14366);
nand UO_847 (O_847,N_14755,N_14703);
nand UO_848 (O_848,N_14333,N_14052);
nor UO_849 (O_849,N_14102,N_14453);
nor UO_850 (O_850,N_14776,N_14398);
or UO_851 (O_851,N_14242,N_14748);
or UO_852 (O_852,N_14759,N_14251);
nor UO_853 (O_853,N_14108,N_14848);
or UO_854 (O_854,N_14257,N_14301);
or UO_855 (O_855,N_14262,N_14711);
and UO_856 (O_856,N_14260,N_14554);
nand UO_857 (O_857,N_14521,N_14355);
and UO_858 (O_858,N_14353,N_14218);
nor UO_859 (O_859,N_14631,N_14459);
and UO_860 (O_860,N_14416,N_14623);
xor UO_861 (O_861,N_14346,N_14309);
nor UO_862 (O_862,N_14850,N_14291);
nand UO_863 (O_863,N_14555,N_14064);
nor UO_864 (O_864,N_14622,N_14366);
nor UO_865 (O_865,N_14985,N_14513);
nor UO_866 (O_866,N_14852,N_14003);
and UO_867 (O_867,N_14282,N_14774);
or UO_868 (O_868,N_14309,N_14205);
xnor UO_869 (O_869,N_14074,N_14434);
nor UO_870 (O_870,N_14477,N_14300);
and UO_871 (O_871,N_14290,N_14883);
nor UO_872 (O_872,N_14221,N_14172);
xor UO_873 (O_873,N_14010,N_14353);
xnor UO_874 (O_874,N_14938,N_14504);
xor UO_875 (O_875,N_14175,N_14628);
nand UO_876 (O_876,N_14326,N_14155);
nand UO_877 (O_877,N_14570,N_14234);
and UO_878 (O_878,N_14419,N_14682);
nand UO_879 (O_879,N_14063,N_14712);
or UO_880 (O_880,N_14137,N_14282);
and UO_881 (O_881,N_14672,N_14253);
xor UO_882 (O_882,N_14390,N_14343);
and UO_883 (O_883,N_14845,N_14989);
xnor UO_884 (O_884,N_14525,N_14056);
nand UO_885 (O_885,N_14801,N_14001);
xnor UO_886 (O_886,N_14097,N_14791);
or UO_887 (O_887,N_14207,N_14417);
nor UO_888 (O_888,N_14233,N_14294);
and UO_889 (O_889,N_14349,N_14670);
nand UO_890 (O_890,N_14473,N_14228);
and UO_891 (O_891,N_14004,N_14531);
nand UO_892 (O_892,N_14398,N_14856);
xor UO_893 (O_893,N_14130,N_14533);
and UO_894 (O_894,N_14345,N_14438);
xnor UO_895 (O_895,N_14862,N_14404);
nor UO_896 (O_896,N_14424,N_14620);
and UO_897 (O_897,N_14406,N_14198);
or UO_898 (O_898,N_14858,N_14239);
nand UO_899 (O_899,N_14939,N_14280);
nand UO_900 (O_900,N_14193,N_14960);
or UO_901 (O_901,N_14682,N_14899);
nor UO_902 (O_902,N_14856,N_14308);
or UO_903 (O_903,N_14938,N_14382);
nand UO_904 (O_904,N_14726,N_14372);
or UO_905 (O_905,N_14289,N_14515);
nor UO_906 (O_906,N_14133,N_14492);
and UO_907 (O_907,N_14377,N_14386);
xor UO_908 (O_908,N_14449,N_14001);
nand UO_909 (O_909,N_14899,N_14389);
xor UO_910 (O_910,N_14174,N_14050);
xor UO_911 (O_911,N_14304,N_14570);
and UO_912 (O_912,N_14883,N_14906);
xnor UO_913 (O_913,N_14007,N_14561);
or UO_914 (O_914,N_14590,N_14559);
nand UO_915 (O_915,N_14329,N_14728);
nor UO_916 (O_916,N_14750,N_14129);
xor UO_917 (O_917,N_14424,N_14144);
nor UO_918 (O_918,N_14010,N_14077);
nor UO_919 (O_919,N_14036,N_14997);
or UO_920 (O_920,N_14276,N_14665);
nor UO_921 (O_921,N_14793,N_14703);
nand UO_922 (O_922,N_14050,N_14153);
nor UO_923 (O_923,N_14316,N_14675);
and UO_924 (O_924,N_14010,N_14368);
or UO_925 (O_925,N_14541,N_14240);
nand UO_926 (O_926,N_14097,N_14441);
nor UO_927 (O_927,N_14220,N_14974);
xor UO_928 (O_928,N_14526,N_14240);
nor UO_929 (O_929,N_14622,N_14493);
nand UO_930 (O_930,N_14585,N_14406);
or UO_931 (O_931,N_14897,N_14193);
and UO_932 (O_932,N_14218,N_14719);
nor UO_933 (O_933,N_14130,N_14033);
nor UO_934 (O_934,N_14612,N_14714);
or UO_935 (O_935,N_14640,N_14089);
and UO_936 (O_936,N_14293,N_14279);
or UO_937 (O_937,N_14646,N_14092);
and UO_938 (O_938,N_14924,N_14793);
or UO_939 (O_939,N_14497,N_14662);
nor UO_940 (O_940,N_14565,N_14468);
xor UO_941 (O_941,N_14927,N_14561);
or UO_942 (O_942,N_14695,N_14437);
or UO_943 (O_943,N_14740,N_14896);
nor UO_944 (O_944,N_14461,N_14571);
or UO_945 (O_945,N_14683,N_14078);
and UO_946 (O_946,N_14994,N_14986);
nand UO_947 (O_947,N_14925,N_14227);
nand UO_948 (O_948,N_14178,N_14058);
or UO_949 (O_949,N_14554,N_14105);
xor UO_950 (O_950,N_14025,N_14800);
nand UO_951 (O_951,N_14889,N_14518);
nand UO_952 (O_952,N_14500,N_14954);
nand UO_953 (O_953,N_14974,N_14329);
and UO_954 (O_954,N_14619,N_14004);
xor UO_955 (O_955,N_14239,N_14043);
nor UO_956 (O_956,N_14691,N_14864);
and UO_957 (O_957,N_14950,N_14829);
nand UO_958 (O_958,N_14411,N_14248);
or UO_959 (O_959,N_14999,N_14920);
and UO_960 (O_960,N_14300,N_14554);
or UO_961 (O_961,N_14607,N_14083);
and UO_962 (O_962,N_14679,N_14619);
xor UO_963 (O_963,N_14756,N_14838);
and UO_964 (O_964,N_14362,N_14391);
nor UO_965 (O_965,N_14280,N_14935);
and UO_966 (O_966,N_14608,N_14859);
nand UO_967 (O_967,N_14440,N_14915);
nor UO_968 (O_968,N_14293,N_14725);
nor UO_969 (O_969,N_14070,N_14408);
nor UO_970 (O_970,N_14140,N_14346);
nor UO_971 (O_971,N_14655,N_14271);
xor UO_972 (O_972,N_14951,N_14021);
xnor UO_973 (O_973,N_14141,N_14247);
nand UO_974 (O_974,N_14749,N_14439);
xnor UO_975 (O_975,N_14528,N_14702);
and UO_976 (O_976,N_14612,N_14709);
or UO_977 (O_977,N_14298,N_14698);
nor UO_978 (O_978,N_14688,N_14180);
and UO_979 (O_979,N_14815,N_14408);
and UO_980 (O_980,N_14243,N_14719);
xnor UO_981 (O_981,N_14264,N_14405);
and UO_982 (O_982,N_14310,N_14084);
nor UO_983 (O_983,N_14044,N_14075);
or UO_984 (O_984,N_14841,N_14578);
and UO_985 (O_985,N_14716,N_14261);
or UO_986 (O_986,N_14456,N_14836);
or UO_987 (O_987,N_14895,N_14402);
and UO_988 (O_988,N_14950,N_14625);
or UO_989 (O_989,N_14151,N_14779);
and UO_990 (O_990,N_14634,N_14523);
xor UO_991 (O_991,N_14650,N_14691);
nand UO_992 (O_992,N_14916,N_14154);
or UO_993 (O_993,N_14411,N_14044);
nor UO_994 (O_994,N_14131,N_14061);
nand UO_995 (O_995,N_14945,N_14838);
nand UO_996 (O_996,N_14983,N_14530);
nor UO_997 (O_997,N_14366,N_14987);
and UO_998 (O_998,N_14467,N_14808);
xor UO_999 (O_999,N_14657,N_14780);
xor UO_1000 (O_1000,N_14309,N_14838);
nor UO_1001 (O_1001,N_14893,N_14595);
nor UO_1002 (O_1002,N_14500,N_14975);
xor UO_1003 (O_1003,N_14488,N_14928);
or UO_1004 (O_1004,N_14145,N_14082);
nor UO_1005 (O_1005,N_14432,N_14725);
nor UO_1006 (O_1006,N_14264,N_14051);
nor UO_1007 (O_1007,N_14748,N_14747);
nand UO_1008 (O_1008,N_14787,N_14763);
nor UO_1009 (O_1009,N_14867,N_14689);
xor UO_1010 (O_1010,N_14560,N_14973);
or UO_1011 (O_1011,N_14962,N_14297);
or UO_1012 (O_1012,N_14957,N_14637);
xnor UO_1013 (O_1013,N_14363,N_14872);
xor UO_1014 (O_1014,N_14516,N_14001);
and UO_1015 (O_1015,N_14597,N_14636);
and UO_1016 (O_1016,N_14950,N_14861);
or UO_1017 (O_1017,N_14521,N_14588);
and UO_1018 (O_1018,N_14131,N_14516);
nor UO_1019 (O_1019,N_14276,N_14348);
or UO_1020 (O_1020,N_14966,N_14450);
xor UO_1021 (O_1021,N_14794,N_14386);
and UO_1022 (O_1022,N_14251,N_14884);
or UO_1023 (O_1023,N_14091,N_14663);
xor UO_1024 (O_1024,N_14707,N_14054);
or UO_1025 (O_1025,N_14423,N_14633);
nor UO_1026 (O_1026,N_14021,N_14481);
xor UO_1027 (O_1027,N_14976,N_14862);
and UO_1028 (O_1028,N_14410,N_14351);
and UO_1029 (O_1029,N_14405,N_14796);
nor UO_1030 (O_1030,N_14081,N_14817);
xnor UO_1031 (O_1031,N_14318,N_14366);
nand UO_1032 (O_1032,N_14338,N_14158);
or UO_1033 (O_1033,N_14528,N_14274);
xnor UO_1034 (O_1034,N_14251,N_14766);
and UO_1035 (O_1035,N_14449,N_14052);
xnor UO_1036 (O_1036,N_14728,N_14558);
xnor UO_1037 (O_1037,N_14774,N_14883);
xnor UO_1038 (O_1038,N_14564,N_14555);
and UO_1039 (O_1039,N_14185,N_14850);
and UO_1040 (O_1040,N_14539,N_14457);
nand UO_1041 (O_1041,N_14694,N_14105);
and UO_1042 (O_1042,N_14723,N_14040);
and UO_1043 (O_1043,N_14481,N_14698);
xor UO_1044 (O_1044,N_14666,N_14804);
or UO_1045 (O_1045,N_14260,N_14988);
and UO_1046 (O_1046,N_14298,N_14575);
xnor UO_1047 (O_1047,N_14319,N_14820);
or UO_1048 (O_1048,N_14975,N_14209);
xnor UO_1049 (O_1049,N_14434,N_14291);
or UO_1050 (O_1050,N_14355,N_14551);
and UO_1051 (O_1051,N_14345,N_14953);
xnor UO_1052 (O_1052,N_14326,N_14011);
nor UO_1053 (O_1053,N_14117,N_14885);
or UO_1054 (O_1054,N_14773,N_14570);
and UO_1055 (O_1055,N_14507,N_14990);
nand UO_1056 (O_1056,N_14894,N_14952);
nand UO_1057 (O_1057,N_14952,N_14018);
and UO_1058 (O_1058,N_14236,N_14373);
xnor UO_1059 (O_1059,N_14400,N_14146);
xnor UO_1060 (O_1060,N_14556,N_14304);
and UO_1061 (O_1061,N_14317,N_14147);
and UO_1062 (O_1062,N_14228,N_14560);
xor UO_1063 (O_1063,N_14612,N_14481);
and UO_1064 (O_1064,N_14336,N_14332);
or UO_1065 (O_1065,N_14893,N_14040);
nand UO_1066 (O_1066,N_14532,N_14827);
xnor UO_1067 (O_1067,N_14961,N_14743);
nor UO_1068 (O_1068,N_14857,N_14052);
xor UO_1069 (O_1069,N_14628,N_14239);
xnor UO_1070 (O_1070,N_14031,N_14421);
nand UO_1071 (O_1071,N_14830,N_14726);
nor UO_1072 (O_1072,N_14249,N_14888);
or UO_1073 (O_1073,N_14284,N_14453);
xnor UO_1074 (O_1074,N_14366,N_14539);
nor UO_1075 (O_1075,N_14178,N_14990);
and UO_1076 (O_1076,N_14549,N_14809);
nand UO_1077 (O_1077,N_14444,N_14526);
and UO_1078 (O_1078,N_14426,N_14978);
nand UO_1079 (O_1079,N_14989,N_14569);
nand UO_1080 (O_1080,N_14227,N_14689);
or UO_1081 (O_1081,N_14111,N_14954);
xnor UO_1082 (O_1082,N_14071,N_14391);
xor UO_1083 (O_1083,N_14618,N_14368);
and UO_1084 (O_1084,N_14850,N_14103);
and UO_1085 (O_1085,N_14642,N_14748);
nand UO_1086 (O_1086,N_14980,N_14971);
nor UO_1087 (O_1087,N_14692,N_14841);
nand UO_1088 (O_1088,N_14846,N_14883);
and UO_1089 (O_1089,N_14364,N_14133);
xnor UO_1090 (O_1090,N_14337,N_14046);
and UO_1091 (O_1091,N_14324,N_14960);
xor UO_1092 (O_1092,N_14407,N_14012);
nor UO_1093 (O_1093,N_14895,N_14951);
nand UO_1094 (O_1094,N_14729,N_14336);
xor UO_1095 (O_1095,N_14551,N_14122);
nor UO_1096 (O_1096,N_14241,N_14053);
nor UO_1097 (O_1097,N_14402,N_14151);
and UO_1098 (O_1098,N_14852,N_14904);
nand UO_1099 (O_1099,N_14072,N_14405);
nand UO_1100 (O_1100,N_14963,N_14324);
nand UO_1101 (O_1101,N_14537,N_14297);
or UO_1102 (O_1102,N_14824,N_14590);
xnor UO_1103 (O_1103,N_14483,N_14150);
and UO_1104 (O_1104,N_14124,N_14043);
or UO_1105 (O_1105,N_14321,N_14047);
or UO_1106 (O_1106,N_14944,N_14018);
nor UO_1107 (O_1107,N_14657,N_14671);
and UO_1108 (O_1108,N_14253,N_14737);
or UO_1109 (O_1109,N_14956,N_14665);
or UO_1110 (O_1110,N_14933,N_14492);
nor UO_1111 (O_1111,N_14006,N_14700);
xnor UO_1112 (O_1112,N_14348,N_14708);
nor UO_1113 (O_1113,N_14796,N_14285);
nand UO_1114 (O_1114,N_14642,N_14198);
and UO_1115 (O_1115,N_14828,N_14931);
nor UO_1116 (O_1116,N_14442,N_14873);
or UO_1117 (O_1117,N_14403,N_14986);
xor UO_1118 (O_1118,N_14964,N_14216);
nor UO_1119 (O_1119,N_14187,N_14026);
and UO_1120 (O_1120,N_14380,N_14115);
or UO_1121 (O_1121,N_14343,N_14679);
xnor UO_1122 (O_1122,N_14055,N_14756);
xor UO_1123 (O_1123,N_14225,N_14627);
or UO_1124 (O_1124,N_14725,N_14010);
nand UO_1125 (O_1125,N_14785,N_14427);
nand UO_1126 (O_1126,N_14224,N_14296);
and UO_1127 (O_1127,N_14669,N_14421);
xnor UO_1128 (O_1128,N_14853,N_14710);
and UO_1129 (O_1129,N_14876,N_14800);
nor UO_1130 (O_1130,N_14838,N_14406);
xor UO_1131 (O_1131,N_14256,N_14447);
xnor UO_1132 (O_1132,N_14711,N_14267);
xnor UO_1133 (O_1133,N_14749,N_14973);
or UO_1134 (O_1134,N_14933,N_14205);
nor UO_1135 (O_1135,N_14125,N_14938);
xnor UO_1136 (O_1136,N_14057,N_14296);
xnor UO_1137 (O_1137,N_14380,N_14895);
xor UO_1138 (O_1138,N_14713,N_14046);
xnor UO_1139 (O_1139,N_14284,N_14791);
xor UO_1140 (O_1140,N_14981,N_14280);
or UO_1141 (O_1141,N_14564,N_14027);
or UO_1142 (O_1142,N_14737,N_14677);
and UO_1143 (O_1143,N_14150,N_14524);
nand UO_1144 (O_1144,N_14894,N_14792);
nor UO_1145 (O_1145,N_14538,N_14154);
nand UO_1146 (O_1146,N_14958,N_14223);
xor UO_1147 (O_1147,N_14694,N_14395);
and UO_1148 (O_1148,N_14647,N_14115);
and UO_1149 (O_1149,N_14474,N_14671);
nand UO_1150 (O_1150,N_14327,N_14096);
nand UO_1151 (O_1151,N_14232,N_14116);
or UO_1152 (O_1152,N_14769,N_14391);
and UO_1153 (O_1153,N_14309,N_14162);
xnor UO_1154 (O_1154,N_14483,N_14140);
xnor UO_1155 (O_1155,N_14374,N_14971);
and UO_1156 (O_1156,N_14515,N_14680);
or UO_1157 (O_1157,N_14691,N_14840);
nand UO_1158 (O_1158,N_14913,N_14646);
or UO_1159 (O_1159,N_14804,N_14954);
nor UO_1160 (O_1160,N_14990,N_14960);
xnor UO_1161 (O_1161,N_14869,N_14124);
nand UO_1162 (O_1162,N_14466,N_14057);
nand UO_1163 (O_1163,N_14861,N_14781);
nand UO_1164 (O_1164,N_14833,N_14438);
nor UO_1165 (O_1165,N_14108,N_14027);
nor UO_1166 (O_1166,N_14079,N_14210);
or UO_1167 (O_1167,N_14734,N_14621);
nand UO_1168 (O_1168,N_14330,N_14249);
and UO_1169 (O_1169,N_14082,N_14347);
xnor UO_1170 (O_1170,N_14836,N_14154);
or UO_1171 (O_1171,N_14504,N_14727);
nand UO_1172 (O_1172,N_14910,N_14547);
nand UO_1173 (O_1173,N_14756,N_14313);
and UO_1174 (O_1174,N_14803,N_14173);
nand UO_1175 (O_1175,N_14647,N_14949);
and UO_1176 (O_1176,N_14028,N_14827);
xor UO_1177 (O_1177,N_14544,N_14680);
nand UO_1178 (O_1178,N_14844,N_14863);
or UO_1179 (O_1179,N_14347,N_14308);
or UO_1180 (O_1180,N_14606,N_14623);
and UO_1181 (O_1181,N_14284,N_14866);
nor UO_1182 (O_1182,N_14381,N_14814);
and UO_1183 (O_1183,N_14784,N_14884);
xor UO_1184 (O_1184,N_14477,N_14073);
nand UO_1185 (O_1185,N_14376,N_14816);
or UO_1186 (O_1186,N_14177,N_14100);
nor UO_1187 (O_1187,N_14701,N_14813);
or UO_1188 (O_1188,N_14063,N_14169);
nand UO_1189 (O_1189,N_14332,N_14021);
nand UO_1190 (O_1190,N_14311,N_14304);
nand UO_1191 (O_1191,N_14232,N_14844);
nor UO_1192 (O_1192,N_14148,N_14374);
nand UO_1193 (O_1193,N_14722,N_14503);
and UO_1194 (O_1194,N_14706,N_14443);
or UO_1195 (O_1195,N_14294,N_14114);
and UO_1196 (O_1196,N_14206,N_14257);
nand UO_1197 (O_1197,N_14234,N_14364);
xnor UO_1198 (O_1198,N_14315,N_14487);
nand UO_1199 (O_1199,N_14289,N_14551);
nor UO_1200 (O_1200,N_14234,N_14104);
nor UO_1201 (O_1201,N_14552,N_14848);
xor UO_1202 (O_1202,N_14653,N_14582);
and UO_1203 (O_1203,N_14627,N_14521);
nor UO_1204 (O_1204,N_14928,N_14478);
nand UO_1205 (O_1205,N_14472,N_14595);
and UO_1206 (O_1206,N_14338,N_14922);
nor UO_1207 (O_1207,N_14320,N_14571);
xnor UO_1208 (O_1208,N_14640,N_14151);
or UO_1209 (O_1209,N_14979,N_14346);
xnor UO_1210 (O_1210,N_14743,N_14756);
nor UO_1211 (O_1211,N_14822,N_14736);
nor UO_1212 (O_1212,N_14188,N_14438);
xor UO_1213 (O_1213,N_14673,N_14083);
nand UO_1214 (O_1214,N_14403,N_14088);
or UO_1215 (O_1215,N_14906,N_14361);
xor UO_1216 (O_1216,N_14778,N_14589);
xor UO_1217 (O_1217,N_14111,N_14329);
nand UO_1218 (O_1218,N_14504,N_14680);
or UO_1219 (O_1219,N_14688,N_14345);
xnor UO_1220 (O_1220,N_14146,N_14322);
or UO_1221 (O_1221,N_14958,N_14194);
nand UO_1222 (O_1222,N_14969,N_14359);
nor UO_1223 (O_1223,N_14536,N_14406);
or UO_1224 (O_1224,N_14931,N_14046);
nand UO_1225 (O_1225,N_14622,N_14877);
nor UO_1226 (O_1226,N_14303,N_14537);
and UO_1227 (O_1227,N_14710,N_14886);
xnor UO_1228 (O_1228,N_14553,N_14141);
or UO_1229 (O_1229,N_14404,N_14908);
nand UO_1230 (O_1230,N_14948,N_14459);
xor UO_1231 (O_1231,N_14596,N_14521);
xnor UO_1232 (O_1232,N_14754,N_14745);
nand UO_1233 (O_1233,N_14591,N_14172);
or UO_1234 (O_1234,N_14775,N_14632);
and UO_1235 (O_1235,N_14110,N_14920);
nand UO_1236 (O_1236,N_14737,N_14517);
or UO_1237 (O_1237,N_14385,N_14569);
nand UO_1238 (O_1238,N_14425,N_14338);
nand UO_1239 (O_1239,N_14590,N_14311);
or UO_1240 (O_1240,N_14783,N_14168);
and UO_1241 (O_1241,N_14872,N_14993);
xor UO_1242 (O_1242,N_14322,N_14355);
or UO_1243 (O_1243,N_14265,N_14306);
nor UO_1244 (O_1244,N_14668,N_14120);
and UO_1245 (O_1245,N_14602,N_14594);
nor UO_1246 (O_1246,N_14372,N_14184);
and UO_1247 (O_1247,N_14603,N_14253);
nand UO_1248 (O_1248,N_14851,N_14152);
or UO_1249 (O_1249,N_14544,N_14446);
and UO_1250 (O_1250,N_14915,N_14258);
or UO_1251 (O_1251,N_14986,N_14867);
or UO_1252 (O_1252,N_14045,N_14117);
and UO_1253 (O_1253,N_14396,N_14500);
nor UO_1254 (O_1254,N_14081,N_14838);
or UO_1255 (O_1255,N_14026,N_14224);
or UO_1256 (O_1256,N_14175,N_14760);
or UO_1257 (O_1257,N_14929,N_14605);
nor UO_1258 (O_1258,N_14885,N_14130);
or UO_1259 (O_1259,N_14184,N_14207);
nor UO_1260 (O_1260,N_14174,N_14525);
and UO_1261 (O_1261,N_14903,N_14021);
nand UO_1262 (O_1262,N_14788,N_14805);
nand UO_1263 (O_1263,N_14127,N_14529);
nor UO_1264 (O_1264,N_14688,N_14304);
and UO_1265 (O_1265,N_14661,N_14332);
nand UO_1266 (O_1266,N_14808,N_14718);
or UO_1267 (O_1267,N_14653,N_14832);
nor UO_1268 (O_1268,N_14293,N_14034);
or UO_1269 (O_1269,N_14307,N_14852);
nand UO_1270 (O_1270,N_14684,N_14691);
xnor UO_1271 (O_1271,N_14622,N_14439);
nor UO_1272 (O_1272,N_14016,N_14977);
and UO_1273 (O_1273,N_14905,N_14870);
xor UO_1274 (O_1274,N_14719,N_14161);
and UO_1275 (O_1275,N_14165,N_14048);
or UO_1276 (O_1276,N_14709,N_14791);
xnor UO_1277 (O_1277,N_14661,N_14495);
nor UO_1278 (O_1278,N_14317,N_14813);
and UO_1279 (O_1279,N_14656,N_14505);
and UO_1280 (O_1280,N_14286,N_14674);
xor UO_1281 (O_1281,N_14641,N_14117);
nand UO_1282 (O_1282,N_14735,N_14798);
or UO_1283 (O_1283,N_14866,N_14671);
nand UO_1284 (O_1284,N_14006,N_14940);
xnor UO_1285 (O_1285,N_14665,N_14896);
or UO_1286 (O_1286,N_14002,N_14718);
nand UO_1287 (O_1287,N_14370,N_14059);
nor UO_1288 (O_1288,N_14324,N_14173);
nand UO_1289 (O_1289,N_14998,N_14939);
nor UO_1290 (O_1290,N_14626,N_14766);
or UO_1291 (O_1291,N_14819,N_14694);
nand UO_1292 (O_1292,N_14609,N_14891);
nand UO_1293 (O_1293,N_14456,N_14379);
or UO_1294 (O_1294,N_14581,N_14904);
and UO_1295 (O_1295,N_14340,N_14668);
and UO_1296 (O_1296,N_14878,N_14786);
xor UO_1297 (O_1297,N_14653,N_14283);
nand UO_1298 (O_1298,N_14964,N_14561);
nor UO_1299 (O_1299,N_14726,N_14734);
nor UO_1300 (O_1300,N_14682,N_14309);
nor UO_1301 (O_1301,N_14903,N_14861);
xnor UO_1302 (O_1302,N_14706,N_14599);
nor UO_1303 (O_1303,N_14979,N_14963);
nand UO_1304 (O_1304,N_14391,N_14822);
nand UO_1305 (O_1305,N_14080,N_14528);
nand UO_1306 (O_1306,N_14768,N_14711);
nor UO_1307 (O_1307,N_14933,N_14935);
xnor UO_1308 (O_1308,N_14258,N_14707);
nor UO_1309 (O_1309,N_14439,N_14789);
xor UO_1310 (O_1310,N_14312,N_14875);
xor UO_1311 (O_1311,N_14802,N_14104);
and UO_1312 (O_1312,N_14385,N_14513);
and UO_1313 (O_1313,N_14136,N_14351);
or UO_1314 (O_1314,N_14006,N_14290);
nor UO_1315 (O_1315,N_14433,N_14672);
or UO_1316 (O_1316,N_14736,N_14538);
xnor UO_1317 (O_1317,N_14181,N_14857);
and UO_1318 (O_1318,N_14223,N_14362);
nand UO_1319 (O_1319,N_14799,N_14157);
xor UO_1320 (O_1320,N_14124,N_14650);
xor UO_1321 (O_1321,N_14231,N_14726);
nand UO_1322 (O_1322,N_14733,N_14766);
nand UO_1323 (O_1323,N_14741,N_14451);
nand UO_1324 (O_1324,N_14857,N_14109);
xnor UO_1325 (O_1325,N_14325,N_14672);
or UO_1326 (O_1326,N_14484,N_14339);
xor UO_1327 (O_1327,N_14576,N_14079);
and UO_1328 (O_1328,N_14672,N_14618);
nand UO_1329 (O_1329,N_14839,N_14969);
nor UO_1330 (O_1330,N_14313,N_14133);
or UO_1331 (O_1331,N_14266,N_14363);
or UO_1332 (O_1332,N_14891,N_14467);
xnor UO_1333 (O_1333,N_14308,N_14996);
nor UO_1334 (O_1334,N_14431,N_14137);
or UO_1335 (O_1335,N_14253,N_14398);
or UO_1336 (O_1336,N_14039,N_14033);
and UO_1337 (O_1337,N_14685,N_14010);
or UO_1338 (O_1338,N_14462,N_14778);
xnor UO_1339 (O_1339,N_14320,N_14595);
nand UO_1340 (O_1340,N_14888,N_14404);
or UO_1341 (O_1341,N_14886,N_14564);
nand UO_1342 (O_1342,N_14134,N_14792);
xnor UO_1343 (O_1343,N_14220,N_14972);
nor UO_1344 (O_1344,N_14428,N_14407);
nor UO_1345 (O_1345,N_14058,N_14316);
nor UO_1346 (O_1346,N_14127,N_14627);
and UO_1347 (O_1347,N_14098,N_14801);
and UO_1348 (O_1348,N_14596,N_14699);
nand UO_1349 (O_1349,N_14850,N_14354);
or UO_1350 (O_1350,N_14957,N_14259);
nor UO_1351 (O_1351,N_14042,N_14560);
and UO_1352 (O_1352,N_14444,N_14080);
nor UO_1353 (O_1353,N_14171,N_14173);
xnor UO_1354 (O_1354,N_14821,N_14178);
or UO_1355 (O_1355,N_14750,N_14504);
or UO_1356 (O_1356,N_14388,N_14279);
xor UO_1357 (O_1357,N_14523,N_14001);
or UO_1358 (O_1358,N_14355,N_14888);
nor UO_1359 (O_1359,N_14023,N_14432);
nand UO_1360 (O_1360,N_14173,N_14110);
nor UO_1361 (O_1361,N_14232,N_14503);
nand UO_1362 (O_1362,N_14338,N_14673);
and UO_1363 (O_1363,N_14437,N_14070);
xor UO_1364 (O_1364,N_14382,N_14793);
nor UO_1365 (O_1365,N_14728,N_14005);
and UO_1366 (O_1366,N_14155,N_14384);
nand UO_1367 (O_1367,N_14958,N_14818);
nand UO_1368 (O_1368,N_14298,N_14225);
or UO_1369 (O_1369,N_14680,N_14283);
or UO_1370 (O_1370,N_14406,N_14444);
nand UO_1371 (O_1371,N_14421,N_14282);
or UO_1372 (O_1372,N_14384,N_14083);
and UO_1373 (O_1373,N_14546,N_14057);
xnor UO_1374 (O_1374,N_14484,N_14476);
nor UO_1375 (O_1375,N_14019,N_14784);
and UO_1376 (O_1376,N_14556,N_14323);
nor UO_1377 (O_1377,N_14917,N_14337);
nor UO_1378 (O_1378,N_14937,N_14234);
nand UO_1379 (O_1379,N_14386,N_14148);
and UO_1380 (O_1380,N_14418,N_14028);
nor UO_1381 (O_1381,N_14999,N_14866);
nand UO_1382 (O_1382,N_14134,N_14609);
or UO_1383 (O_1383,N_14727,N_14345);
nand UO_1384 (O_1384,N_14518,N_14587);
nor UO_1385 (O_1385,N_14072,N_14233);
nor UO_1386 (O_1386,N_14804,N_14849);
nand UO_1387 (O_1387,N_14160,N_14595);
nor UO_1388 (O_1388,N_14728,N_14832);
nand UO_1389 (O_1389,N_14860,N_14540);
and UO_1390 (O_1390,N_14192,N_14333);
and UO_1391 (O_1391,N_14217,N_14572);
nand UO_1392 (O_1392,N_14116,N_14886);
nand UO_1393 (O_1393,N_14877,N_14786);
or UO_1394 (O_1394,N_14380,N_14577);
and UO_1395 (O_1395,N_14292,N_14411);
or UO_1396 (O_1396,N_14162,N_14477);
xor UO_1397 (O_1397,N_14340,N_14171);
and UO_1398 (O_1398,N_14800,N_14831);
nand UO_1399 (O_1399,N_14039,N_14261);
nor UO_1400 (O_1400,N_14632,N_14828);
xnor UO_1401 (O_1401,N_14558,N_14254);
and UO_1402 (O_1402,N_14692,N_14658);
nor UO_1403 (O_1403,N_14826,N_14938);
and UO_1404 (O_1404,N_14889,N_14945);
and UO_1405 (O_1405,N_14902,N_14785);
nor UO_1406 (O_1406,N_14913,N_14016);
nor UO_1407 (O_1407,N_14534,N_14828);
and UO_1408 (O_1408,N_14738,N_14622);
nand UO_1409 (O_1409,N_14192,N_14478);
nor UO_1410 (O_1410,N_14416,N_14502);
nand UO_1411 (O_1411,N_14514,N_14390);
or UO_1412 (O_1412,N_14619,N_14930);
nor UO_1413 (O_1413,N_14025,N_14222);
or UO_1414 (O_1414,N_14274,N_14210);
and UO_1415 (O_1415,N_14477,N_14728);
or UO_1416 (O_1416,N_14787,N_14880);
xor UO_1417 (O_1417,N_14464,N_14587);
nor UO_1418 (O_1418,N_14104,N_14246);
nand UO_1419 (O_1419,N_14982,N_14278);
and UO_1420 (O_1420,N_14355,N_14361);
nand UO_1421 (O_1421,N_14120,N_14739);
and UO_1422 (O_1422,N_14618,N_14033);
xnor UO_1423 (O_1423,N_14731,N_14366);
nand UO_1424 (O_1424,N_14105,N_14355);
or UO_1425 (O_1425,N_14568,N_14029);
nand UO_1426 (O_1426,N_14953,N_14752);
nor UO_1427 (O_1427,N_14688,N_14878);
and UO_1428 (O_1428,N_14544,N_14335);
nor UO_1429 (O_1429,N_14497,N_14440);
nand UO_1430 (O_1430,N_14921,N_14750);
or UO_1431 (O_1431,N_14547,N_14525);
or UO_1432 (O_1432,N_14420,N_14609);
xnor UO_1433 (O_1433,N_14285,N_14897);
nor UO_1434 (O_1434,N_14211,N_14701);
or UO_1435 (O_1435,N_14971,N_14037);
and UO_1436 (O_1436,N_14447,N_14368);
xor UO_1437 (O_1437,N_14901,N_14953);
nor UO_1438 (O_1438,N_14043,N_14516);
and UO_1439 (O_1439,N_14476,N_14309);
xnor UO_1440 (O_1440,N_14525,N_14822);
nor UO_1441 (O_1441,N_14213,N_14793);
xor UO_1442 (O_1442,N_14760,N_14213);
nand UO_1443 (O_1443,N_14656,N_14412);
xnor UO_1444 (O_1444,N_14194,N_14243);
nor UO_1445 (O_1445,N_14015,N_14269);
nor UO_1446 (O_1446,N_14773,N_14768);
nor UO_1447 (O_1447,N_14516,N_14108);
and UO_1448 (O_1448,N_14485,N_14716);
nor UO_1449 (O_1449,N_14261,N_14747);
or UO_1450 (O_1450,N_14019,N_14087);
and UO_1451 (O_1451,N_14580,N_14560);
nand UO_1452 (O_1452,N_14912,N_14477);
nor UO_1453 (O_1453,N_14518,N_14074);
nor UO_1454 (O_1454,N_14218,N_14580);
nor UO_1455 (O_1455,N_14343,N_14307);
xor UO_1456 (O_1456,N_14451,N_14724);
nor UO_1457 (O_1457,N_14960,N_14489);
nand UO_1458 (O_1458,N_14352,N_14421);
or UO_1459 (O_1459,N_14957,N_14750);
or UO_1460 (O_1460,N_14788,N_14333);
xor UO_1461 (O_1461,N_14865,N_14198);
xor UO_1462 (O_1462,N_14151,N_14260);
xnor UO_1463 (O_1463,N_14955,N_14774);
xor UO_1464 (O_1464,N_14652,N_14832);
nand UO_1465 (O_1465,N_14520,N_14313);
and UO_1466 (O_1466,N_14187,N_14501);
nor UO_1467 (O_1467,N_14450,N_14205);
xor UO_1468 (O_1468,N_14526,N_14474);
nand UO_1469 (O_1469,N_14255,N_14788);
nor UO_1470 (O_1470,N_14149,N_14392);
nor UO_1471 (O_1471,N_14580,N_14386);
nor UO_1472 (O_1472,N_14930,N_14438);
xnor UO_1473 (O_1473,N_14161,N_14818);
and UO_1474 (O_1474,N_14248,N_14831);
or UO_1475 (O_1475,N_14237,N_14085);
and UO_1476 (O_1476,N_14802,N_14417);
nand UO_1477 (O_1477,N_14986,N_14127);
or UO_1478 (O_1478,N_14653,N_14350);
xor UO_1479 (O_1479,N_14906,N_14230);
nand UO_1480 (O_1480,N_14293,N_14493);
nor UO_1481 (O_1481,N_14885,N_14066);
nand UO_1482 (O_1482,N_14178,N_14686);
and UO_1483 (O_1483,N_14167,N_14160);
xor UO_1484 (O_1484,N_14357,N_14092);
xor UO_1485 (O_1485,N_14388,N_14375);
xor UO_1486 (O_1486,N_14329,N_14904);
nor UO_1487 (O_1487,N_14293,N_14280);
nor UO_1488 (O_1488,N_14167,N_14040);
nand UO_1489 (O_1489,N_14787,N_14943);
and UO_1490 (O_1490,N_14534,N_14540);
nand UO_1491 (O_1491,N_14861,N_14665);
xor UO_1492 (O_1492,N_14908,N_14368);
or UO_1493 (O_1493,N_14002,N_14793);
xor UO_1494 (O_1494,N_14488,N_14282);
and UO_1495 (O_1495,N_14243,N_14224);
xnor UO_1496 (O_1496,N_14345,N_14129);
and UO_1497 (O_1497,N_14613,N_14689);
or UO_1498 (O_1498,N_14701,N_14669);
nor UO_1499 (O_1499,N_14636,N_14457);
xor UO_1500 (O_1500,N_14722,N_14633);
xor UO_1501 (O_1501,N_14329,N_14170);
or UO_1502 (O_1502,N_14422,N_14575);
or UO_1503 (O_1503,N_14907,N_14516);
or UO_1504 (O_1504,N_14270,N_14674);
nand UO_1505 (O_1505,N_14735,N_14064);
nand UO_1506 (O_1506,N_14970,N_14822);
or UO_1507 (O_1507,N_14166,N_14784);
xor UO_1508 (O_1508,N_14602,N_14895);
nand UO_1509 (O_1509,N_14436,N_14543);
nor UO_1510 (O_1510,N_14435,N_14846);
nor UO_1511 (O_1511,N_14869,N_14149);
xnor UO_1512 (O_1512,N_14611,N_14668);
and UO_1513 (O_1513,N_14999,N_14163);
nor UO_1514 (O_1514,N_14737,N_14146);
nor UO_1515 (O_1515,N_14493,N_14486);
or UO_1516 (O_1516,N_14718,N_14715);
nand UO_1517 (O_1517,N_14592,N_14848);
xor UO_1518 (O_1518,N_14105,N_14715);
and UO_1519 (O_1519,N_14351,N_14683);
nand UO_1520 (O_1520,N_14124,N_14169);
and UO_1521 (O_1521,N_14956,N_14544);
nor UO_1522 (O_1522,N_14306,N_14491);
or UO_1523 (O_1523,N_14829,N_14557);
xnor UO_1524 (O_1524,N_14795,N_14094);
xnor UO_1525 (O_1525,N_14941,N_14040);
nor UO_1526 (O_1526,N_14531,N_14062);
and UO_1527 (O_1527,N_14678,N_14751);
nor UO_1528 (O_1528,N_14459,N_14387);
nand UO_1529 (O_1529,N_14648,N_14532);
nand UO_1530 (O_1530,N_14366,N_14342);
nand UO_1531 (O_1531,N_14354,N_14439);
nand UO_1532 (O_1532,N_14167,N_14860);
xnor UO_1533 (O_1533,N_14418,N_14194);
nand UO_1534 (O_1534,N_14919,N_14952);
and UO_1535 (O_1535,N_14592,N_14590);
or UO_1536 (O_1536,N_14394,N_14474);
or UO_1537 (O_1537,N_14070,N_14246);
or UO_1538 (O_1538,N_14587,N_14611);
xnor UO_1539 (O_1539,N_14798,N_14057);
nand UO_1540 (O_1540,N_14083,N_14248);
and UO_1541 (O_1541,N_14705,N_14532);
nand UO_1542 (O_1542,N_14493,N_14286);
and UO_1543 (O_1543,N_14765,N_14425);
or UO_1544 (O_1544,N_14311,N_14060);
nand UO_1545 (O_1545,N_14566,N_14755);
and UO_1546 (O_1546,N_14816,N_14040);
and UO_1547 (O_1547,N_14256,N_14439);
or UO_1548 (O_1548,N_14320,N_14478);
nand UO_1549 (O_1549,N_14905,N_14996);
and UO_1550 (O_1550,N_14209,N_14932);
xnor UO_1551 (O_1551,N_14552,N_14348);
xnor UO_1552 (O_1552,N_14070,N_14844);
xnor UO_1553 (O_1553,N_14959,N_14354);
xor UO_1554 (O_1554,N_14385,N_14988);
and UO_1555 (O_1555,N_14362,N_14294);
and UO_1556 (O_1556,N_14397,N_14143);
nor UO_1557 (O_1557,N_14408,N_14117);
xnor UO_1558 (O_1558,N_14914,N_14949);
nand UO_1559 (O_1559,N_14045,N_14088);
nand UO_1560 (O_1560,N_14691,N_14660);
xor UO_1561 (O_1561,N_14401,N_14055);
nor UO_1562 (O_1562,N_14418,N_14942);
xnor UO_1563 (O_1563,N_14817,N_14062);
xor UO_1564 (O_1564,N_14882,N_14068);
or UO_1565 (O_1565,N_14287,N_14529);
and UO_1566 (O_1566,N_14424,N_14524);
nand UO_1567 (O_1567,N_14963,N_14354);
nor UO_1568 (O_1568,N_14904,N_14864);
nand UO_1569 (O_1569,N_14785,N_14046);
or UO_1570 (O_1570,N_14402,N_14304);
xor UO_1571 (O_1571,N_14187,N_14815);
or UO_1572 (O_1572,N_14259,N_14335);
and UO_1573 (O_1573,N_14959,N_14662);
nor UO_1574 (O_1574,N_14164,N_14461);
or UO_1575 (O_1575,N_14320,N_14194);
xor UO_1576 (O_1576,N_14755,N_14642);
and UO_1577 (O_1577,N_14882,N_14178);
or UO_1578 (O_1578,N_14982,N_14484);
nand UO_1579 (O_1579,N_14324,N_14519);
xnor UO_1580 (O_1580,N_14656,N_14069);
nand UO_1581 (O_1581,N_14522,N_14406);
xnor UO_1582 (O_1582,N_14046,N_14746);
and UO_1583 (O_1583,N_14163,N_14588);
nand UO_1584 (O_1584,N_14613,N_14085);
xor UO_1585 (O_1585,N_14448,N_14760);
xnor UO_1586 (O_1586,N_14107,N_14224);
xnor UO_1587 (O_1587,N_14669,N_14227);
nor UO_1588 (O_1588,N_14450,N_14469);
nand UO_1589 (O_1589,N_14521,N_14327);
and UO_1590 (O_1590,N_14144,N_14642);
nor UO_1591 (O_1591,N_14836,N_14886);
nor UO_1592 (O_1592,N_14338,N_14068);
and UO_1593 (O_1593,N_14767,N_14567);
or UO_1594 (O_1594,N_14079,N_14689);
xor UO_1595 (O_1595,N_14261,N_14529);
nand UO_1596 (O_1596,N_14104,N_14731);
xor UO_1597 (O_1597,N_14746,N_14343);
nand UO_1598 (O_1598,N_14206,N_14458);
nand UO_1599 (O_1599,N_14310,N_14062);
or UO_1600 (O_1600,N_14250,N_14995);
and UO_1601 (O_1601,N_14978,N_14275);
or UO_1602 (O_1602,N_14092,N_14027);
nor UO_1603 (O_1603,N_14919,N_14713);
or UO_1604 (O_1604,N_14286,N_14621);
xnor UO_1605 (O_1605,N_14773,N_14113);
nor UO_1606 (O_1606,N_14012,N_14677);
or UO_1607 (O_1607,N_14001,N_14377);
or UO_1608 (O_1608,N_14035,N_14343);
nor UO_1609 (O_1609,N_14963,N_14533);
and UO_1610 (O_1610,N_14735,N_14748);
xnor UO_1611 (O_1611,N_14879,N_14003);
nor UO_1612 (O_1612,N_14790,N_14484);
nor UO_1613 (O_1613,N_14713,N_14135);
or UO_1614 (O_1614,N_14493,N_14009);
and UO_1615 (O_1615,N_14593,N_14098);
xor UO_1616 (O_1616,N_14591,N_14518);
or UO_1617 (O_1617,N_14868,N_14135);
and UO_1618 (O_1618,N_14190,N_14602);
xor UO_1619 (O_1619,N_14525,N_14421);
nand UO_1620 (O_1620,N_14267,N_14132);
nand UO_1621 (O_1621,N_14555,N_14502);
nor UO_1622 (O_1622,N_14354,N_14153);
or UO_1623 (O_1623,N_14947,N_14292);
xnor UO_1624 (O_1624,N_14679,N_14613);
or UO_1625 (O_1625,N_14431,N_14541);
nand UO_1626 (O_1626,N_14206,N_14548);
nor UO_1627 (O_1627,N_14674,N_14411);
and UO_1628 (O_1628,N_14267,N_14760);
nand UO_1629 (O_1629,N_14479,N_14299);
xor UO_1630 (O_1630,N_14015,N_14865);
and UO_1631 (O_1631,N_14427,N_14642);
nor UO_1632 (O_1632,N_14633,N_14836);
nor UO_1633 (O_1633,N_14072,N_14420);
nor UO_1634 (O_1634,N_14701,N_14618);
nand UO_1635 (O_1635,N_14333,N_14743);
nand UO_1636 (O_1636,N_14724,N_14720);
xnor UO_1637 (O_1637,N_14869,N_14038);
and UO_1638 (O_1638,N_14026,N_14273);
and UO_1639 (O_1639,N_14736,N_14484);
xor UO_1640 (O_1640,N_14855,N_14916);
nand UO_1641 (O_1641,N_14533,N_14983);
nand UO_1642 (O_1642,N_14599,N_14787);
nor UO_1643 (O_1643,N_14433,N_14860);
or UO_1644 (O_1644,N_14088,N_14149);
nand UO_1645 (O_1645,N_14108,N_14234);
nor UO_1646 (O_1646,N_14781,N_14120);
or UO_1647 (O_1647,N_14341,N_14760);
and UO_1648 (O_1648,N_14213,N_14739);
nand UO_1649 (O_1649,N_14794,N_14733);
nor UO_1650 (O_1650,N_14686,N_14783);
or UO_1651 (O_1651,N_14314,N_14716);
nand UO_1652 (O_1652,N_14554,N_14710);
or UO_1653 (O_1653,N_14081,N_14868);
xnor UO_1654 (O_1654,N_14522,N_14948);
or UO_1655 (O_1655,N_14168,N_14161);
and UO_1656 (O_1656,N_14761,N_14321);
nand UO_1657 (O_1657,N_14409,N_14496);
nor UO_1658 (O_1658,N_14228,N_14461);
xor UO_1659 (O_1659,N_14261,N_14998);
or UO_1660 (O_1660,N_14409,N_14898);
nand UO_1661 (O_1661,N_14214,N_14937);
xor UO_1662 (O_1662,N_14618,N_14295);
nand UO_1663 (O_1663,N_14207,N_14498);
nand UO_1664 (O_1664,N_14313,N_14533);
nor UO_1665 (O_1665,N_14330,N_14630);
xnor UO_1666 (O_1666,N_14200,N_14939);
nor UO_1667 (O_1667,N_14616,N_14494);
nand UO_1668 (O_1668,N_14319,N_14454);
nor UO_1669 (O_1669,N_14678,N_14692);
nor UO_1670 (O_1670,N_14031,N_14183);
or UO_1671 (O_1671,N_14935,N_14963);
xor UO_1672 (O_1672,N_14534,N_14845);
or UO_1673 (O_1673,N_14353,N_14688);
nor UO_1674 (O_1674,N_14504,N_14521);
nor UO_1675 (O_1675,N_14230,N_14000);
or UO_1676 (O_1676,N_14657,N_14824);
xor UO_1677 (O_1677,N_14772,N_14004);
nor UO_1678 (O_1678,N_14208,N_14943);
xnor UO_1679 (O_1679,N_14652,N_14048);
and UO_1680 (O_1680,N_14632,N_14279);
or UO_1681 (O_1681,N_14343,N_14173);
nor UO_1682 (O_1682,N_14094,N_14680);
nand UO_1683 (O_1683,N_14781,N_14430);
xnor UO_1684 (O_1684,N_14298,N_14643);
xnor UO_1685 (O_1685,N_14405,N_14964);
xnor UO_1686 (O_1686,N_14576,N_14024);
or UO_1687 (O_1687,N_14215,N_14892);
xnor UO_1688 (O_1688,N_14953,N_14630);
nor UO_1689 (O_1689,N_14389,N_14888);
xor UO_1690 (O_1690,N_14686,N_14485);
nor UO_1691 (O_1691,N_14941,N_14009);
nand UO_1692 (O_1692,N_14999,N_14286);
or UO_1693 (O_1693,N_14495,N_14069);
and UO_1694 (O_1694,N_14469,N_14088);
xor UO_1695 (O_1695,N_14490,N_14327);
nand UO_1696 (O_1696,N_14972,N_14988);
xor UO_1697 (O_1697,N_14429,N_14855);
nor UO_1698 (O_1698,N_14454,N_14471);
and UO_1699 (O_1699,N_14231,N_14268);
xnor UO_1700 (O_1700,N_14491,N_14448);
or UO_1701 (O_1701,N_14262,N_14665);
xor UO_1702 (O_1702,N_14369,N_14133);
or UO_1703 (O_1703,N_14221,N_14207);
xnor UO_1704 (O_1704,N_14172,N_14220);
and UO_1705 (O_1705,N_14783,N_14450);
xnor UO_1706 (O_1706,N_14478,N_14071);
and UO_1707 (O_1707,N_14261,N_14138);
or UO_1708 (O_1708,N_14822,N_14755);
nand UO_1709 (O_1709,N_14511,N_14292);
nand UO_1710 (O_1710,N_14005,N_14471);
xor UO_1711 (O_1711,N_14217,N_14943);
and UO_1712 (O_1712,N_14746,N_14559);
or UO_1713 (O_1713,N_14168,N_14635);
xor UO_1714 (O_1714,N_14903,N_14441);
nor UO_1715 (O_1715,N_14764,N_14840);
or UO_1716 (O_1716,N_14995,N_14459);
xor UO_1717 (O_1717,N_14352,N_14211);
or UO_1718 (O_1718,N_14896,N_14037);
or UO_1719 (O_1719,N_14473,N_14496);
nor UO_1720 (O_1720,N_14377,N_14490);
and UO_1721 (O_1721,N_14103,N_14581);
nor UO_1722 (O_1722,N_14381,N_14017);
xnor UO_1723 (O_1723,N_14314,N_14334);
or UO_1724 (O_1724,N_14448,N_14877);
nor UO_1725 (O_1725,N_14958,N_14240);
xnor UO_1726 (O_1726,N_14064,N_14408);
or UO_1727 (O_1727,N_14205,N_14266);
or UO_1728 (O_1728,N_14420,N_14005);
and UO_1729 (O_1729,N_14902,N_14149);
nor UO_1730 (O_1730,N_14875,N_14909);
nand UO_1731 (O_1731,N_14874,N_14040);
xnor UO_1732 (O_1732,N_14708,N_14815);
or UO_1733 (O_1733,N_14375,N_14642);
or UO_1734 (O_1734,N_14965,N_14460);
nor UO_1735 (O_1735,N_14163,N_14403);
or UO_1736 (O_1736,N_14637,N_14144);
and UO_1737 (O_1737,N_14646,N_14264);
xnor UO_1738 (O_1738,N_14095,N_14237);
and UO_1739 (O_1739,N_14870,N_14623);
or UO_1740 (O_1740,N_14843,N_14251);
xnor UO_1741 (O_1741,N_14402,N_14710);
nand UO_1742 (O_1742,N_14222,N_14609);
xor UO_1743 (O_1743,N_14318,N_14923);
nand UO_1744 (O_1744,N_14016,N_14988);
xnor UO_1745 (O_1745,N_14913,N_14728);
and UO_1746 (O_1746,N_14801,N_14794);
or UO_1747 (O_1747,N_14002,N_14743);
or UO_1748 (O_1748,N_14624,N_14433);
nor UO_1749 (O_1749,N_14057,N_14739);
xnor UO_1750 (O_1750,N_14265,N_14154);
and UO_1751 (O_1751,N_14152,N_14055);
nand UO_1752 (O_1752,N_14061,N_14588);
nand UO_1753 (O_1753,N_14645,N_14920);
nor UO_1754 (O_1754,N_14017,N_14051);
or UO_1755 (O_1755,N_14614,N_14484);
xor UO_1756 (O_1756,N_14863,N_14091);
nor UO_1757 (O_1757,N_14185,N_14500);
and UO_1758 (O_1758,N_14594,N_14923);
nor UO_1759 (O_1759,N_14133,N_14665);
or UO_1760 (O_1760,N_14934,N_14529);
or UO_1761 (O_1761,N_14231,N_14303);
nand UO_1762 (O_1762,N_14973,N_14231);
or UO_1763 (O_1763,N_14572,N_14367);
xnor UO_1764 (O_1764,N_14645,N_14268);
xnor UO_1765 (O_1765,N_14602,N_14513);
or UO_1766 (O_1766,N_14091,N_14894);
nand UO_1767 (O_1767,N_14302,N_14613);
nand UO_1768 (O_1768,N_14325,N_14181);
and UO_1769 (O_1769,N_14985,N_14103);
and UO_1770 (O_1770,N_14219,N_14568);
or UO_1771 (O_1771,N_14095,N_14295);
nor UO_1772 (O_1772,N_14523,N_14199);
nor UO_1773 (O_1773,N_14744,N_14790);
nand UO_1774 (O_1774,N_14634,N_14063);
xnor UO_1775 (O_1775,N_14783,N_14965);
nor UO_1776 (O_1776,N_14216,N_14292);
nand UO_1777 (O_1777,N_14228,N_14531);
nor UO_1778 (O_1778,N_14768,N_14862);
and UO_1779 (O_1779,N_14173,N_14704);
nand UO_1780 (O_1780,N_14351,N_14644);
nand UO_1781 (O_1781,N_14795,N_14611);
xor UO_1782 (O_1782,N_14632,N_14291);
nor UO_1783 (O_1783,N_14384,N_14179);
and UO_1784 (O_1784,N_14524,N_14941);
and UO_1785 (O_1785,N_14729,N_14861);
xor UO_1786 (O_1786,N_14646,N_14990);
nand UO_1787 (O_1787,N_14087,N_14440);
nor UO_1788 (O_1788,N_14012,N_14669);
nand UO_1789 (O_1789,N_14846,N_14827);
and UO_1790 (O_1790,N_14443,N_14467);
or UO_1791 (O_1791,N_14182,N_14225);
and UO_1792 (O_1792,N_14269,N_14001);
and UO_1793 (O_1793,N_14625,N_14826);
or UO_1794 (O_1794,N_14667,N_14644);
and UO_1795 (O_1795,N_14246,N_14076);
xor UO_1796 (O_1796,N_14205,N_14247);
nand UO_1797 (O_1797,N_14760,N_14520);
or UO_1798 (O_1798,N_14720,N_14287);
nand UO_1799 (O_1799,N_14772,N_14263);
and UO_1800 (O_1800,N_14816,N_14989);
nand UO_1801 (O_1801,N_14796,N_14116);
xor UO_1802 (O_1802,N_14898,N_14868);
xnor UO_1803 (O_1803,N_14996,N_14696);
or UO_1804 (O_1804,N_14877,N_14740);
and UO_1805 (O_1805,N_14091,N_14539);
nand UO_1806 (O_1806,N_14292,N_14373);
xnor UO_1807 (O_1807,N_14609,N_14838);
and UO_1808 (O_1808,N_14939,N_14919);
or UO_1809 (O_1809,N_14545,N_14201);
or UO_1810 (O_1810,N_14743,N_14919);
or UO_1811 (O_1811,N_14222,N_14185);
nand UO_1812 (O_1812,N_14890,N_14330);
nand UO_1813 (O_1813,N_14008,N_14718);
or UO_1814 (O_1814,N_14997,N_14552);
xnor UO_1815 (O_1815,N_14557,N_14500);
nand UO_1816 (O_1816,N_14312,N_14163);
and UO_1817 (O_1817,N_14319,N_14658);
or UO_1818 (O_1818,N_14243,N_14088);
or UO_1819 (O_1819,N_14147,N_14731);
and UO_1820 (O_1820,N_14996,N_14552);
and UO_1821 (O_1821,N_14010,N_14283);
or UO_1822 (O_1822,N_14985,N_14965);
nand UO_1823 (O_1823,N_14705,N_14361);
or UO_1824 (O_1824,N_14550,N_14336);
nor UO_1825 (O_1825,N_14242,N_14946);
or UO_1826 (O_1826,N_14118,N_14893);
nor UO_1827 (O_1827,N_14879,N_14657);
xnor UO_1828 (O_1828,N_14231,N_14242);
and UO_1829 (O_1829,N_14263,N_14229);
nor UO_1830 (O_1830,N_14021,N_14022);
or UO_1831 (O_1831,N_14743,N_14582);
xnor UO_1832 (O_1832,N_14927,N_14786);
xnor UO_1833 (O_1833,N_14332,N_14062);
xnor UO_1834 (O_1834,N_14106,N_14740);
nand UO_1835 (O_1835,N_14982,N_14644);
xnor UO_1836 (O_1836,N_14541,N_14659);
nand UO_1837 (O_1837,N_14991,N_14089);
and UO_1838 (O_1838,N_14653,N_14619);
and UO_1839 (O_1839,N_14193,N_14372);
nand UO_1840 (O_1840,N_14857,N_14678);
and UO_1841 (O_1841,N_14494,N_14282);
nor UO_1842 (O_1842,N_14458,N_14890);
nor UO_1843 (O_1843,N_14565,N_14267);
xor UO_1844 (O_1844,N_14989,N_14987);
nand UO_1845 (O_1845,N_14258,N_14257);
nor UO_1846 (O_1846,N_14890,N_14428);
nor UO_1847 (O_1847,N_14311,N_14727);
or UO_1848 (O_1848,N_14654,N_14133);
nand UO_1849 (O_1849,N_14906,N_14843);
xor UO_1850 (O_1850,N_14160,N_14327);
and UO_1851 (O_1851,N_14909,N_14728);
xor UO_1852 (O_1852,N_14139,N_14790);
and UO_1853 (O_1853,N_14018,N_14566);
nor UO_1854 (O_1854,N_14040,N_14352);
or UO_1855 (O_1855,N_14721,N_14795);
or UO_1856 (O_1856,N_14585,N_14345);
or UO_1857 (O_1857,N_14561,N_14711);
or UO_1858 (O_1858,N_14770,N_14625);
or UO_1859 (O_1859,N_14030,N_14598);
xnor UO_1860 (O_1860,N_14328,N_14738);
nor UO_1861 (O_1861,N_14685,N_14474);
xnor UO_1862 (O_1862,N_14584,N_14708);
or UO_1863 (O_1863,N_14822,N_14343);
or UO_1864 (O_1864,N_14042,N_14212);
xnor UO_1865 (O_1865,N_14772,N_14977);
nand UO_1866 (O_1866,N_14194,N_14999);
nor UO_1867 (O_1867,N_14752,N_14248);
and UO_1868 (O_1868,N_14000,N_14752);
or UO_1869 (O_1869,N_14047,N_14498);
or UO_1870 (O_1870,N_14896,N_14347);
nor UO_1871 (O_1871,N_14394,N_14053);
and UO_1872 (O_1872,N_14577,N_14596);
nor UO_1873 (O_1873,N_14350,N_14984);
or UO_1874 (O_1874,N_14864,N_14253);
and UO_1875 (O_1875,N_14094,N_14767);
nor UO_1876 (O_1876,N_14947,N_14011);
nand UO_1877 (O_1877,N_14600,N_14331);
xnor UO_1878 (O_1878,N_14509,N_14036);
xnor UO_1879 (O_1879,N_14531,N_14543);
nand UO_1880 (O_1880,N_14298,N_14495);
or UO_1881 (O_1881,N_14610,N_14978);
nand UO_1882 (O_1882,N_14268,N_14436);
nand UO_1883 (O_1883,N_14897,N_14769);
and UO_1884 (O_1884,N_14762,N_14541);
xnor UO_1885 (O_1885,N_14599,N_14136);
and UO_1886 (O_1886,N_14239,N_14465);
xnor UO_1887 (O_1887,N_14620,N_14279);
and UO_1888 (O_1888,N_14929,N_14215);
and UO_1889 (O_1889,N_14238,N_14944);
or UO_1890 (O_1890,N_14254,N_14187);
xnor UO_1891 (O_1891,N_14321,N_14559);
nor UO_1892 (O_1892,N_14731,N_14258);
xnor UO_1893 (O_1893,N_14765,N_14774);
and UO_1894 (O_1894,N_14800,N_14906);
or UO_1895 (O_1895,N_14939,N_14095);
or UO_1896 (O_1896,N_14738,N_14285);
nor UO_1897 (O_1897,N_14710,N_14349);
nor UO_1898 (O_1898,N_14411,N_14014);
nand UO_1899 (O_1899,N_14174,N_14781);
or UO_1900 (O_1900,N_14129,N_14087);
nor UO_1901 (O_1901,N_14131,N_14854);
nor UO_1902 (O_1902,N_14676,N_14356);
xnor UO_1903 (O_1903,N_14804,N_14004);
nand UO_1904 (O_1904,N_14469,N_14693);
xor UO_1905 (O_1905,N_14957,N_14563);
xor UO_1906 (O_1906,N_14264,N_14269);
and UO_1907 (O_1907,N_14973,N_14635);
nor UO_1908 (O_1908,N_14142,N_14786);
xor UO_1909 (O_1909,N_14933,N_14606);
xor UO_1910 (O_1910,N_14950,N_14936);
nor UO_1911 (O_1911,N_14472,N_14622);
or UO_1912 (O_1912,N_14435,N_14444);
or UO_1913 (O_1913,N_14763,N_14859);
nand UO_1914 (O_1914,N_14655,N_14242);
xor UO_1915 (O_1915,N_14604,N_14293);
xor UO_1916 (O_1916,N_14934,N_14089);
or UO_1917 (O_1917,N_14244,N_14653);
or UO_1918 (O_1918,N_14548,N_14505);
nand UO_1919 (O_1919,N_14001,N_14170);
and UO_1920 (O_1920,N_14558,N_14435);
or UO_1921 (O_1921,N_14723,N_14619);
xnor UO_1922 (O_1922,N_14920,N_14903);
nand UO_1923 (O_1923,N_14376,N_14995);
or UO_1924 (O_1924,N_14523,N_14011);
nand UO_1925 (O_1925,N_14034,N_14346);
nand UO_1926 (O_1926,N_14219,N_14731);
nor UO_1927 (O_1927,N_14685,N_14532);
or UO_1928 (O_1928,N_14858,N_14895);
and UO_1929 (O_1929,N_14757,N_14646);
or UO_1930 (O_1930,N_14955,N_14554);
or UO_1931 (O_1931,N_14813,N_14261);
xor UO_1932 (O_1932,N_14939,N_14577);
nand UO_1933 (O_1933,N_14422,N_14824);
nand UO_1934 (O_1934,N_14932,N_14604);
nand UO_1935 (O_1935,N_14435,N_14373);
nor UO_1936 (O_1936,N_14349,N_14048);
and UO_1937 (O_1937,N_14663,N_14937);
or UO_1938 (O_1938,N_14461,N_14376);
nor UO_1939 (O_1939,N_14053,N_14124);
nand UO_1940 (O_1940,N_14357,N_14236);
or UO_1941 (O_1941,N_14857,N_14373);
nand UO_1942 (O_1942,N_14672,N_14549);
nor UO_1943 (O_1943,N_14640,N_14570);
nand UO_1944 (O_1944,N_14834,N_14138);
and UO_1945 (O_1945,N_14988,N_14796);
xor UO_1946 (O_1946,N_14919,N_14593);
nor UO_1947 (O_1947,N_14120,N_14883);
and UO_1948 (O_1948,N_14843,N_14416);
nand UO_1949 (O_1949,N_14739,N_14152);
or UO_1950 (O_1950,N_14333,N_14269);
xnor UO_1951 (O_1951,N_14802,N_14819);
nand UO_1952 (O_1952,N_14232,N_14280);
xnor UO_1953 (O_1953,N_14443,N_14126);
nand UO_1954 (O_1954,N_14790,N_14164);
xor UO_1955 (O_1955,N_14374,N_14622);
nor UO_1956 (O_1956,N_14294,N_14202);
or UO_1957 (O_1957,N_14339,N_14137);
xnor UO_1958 (O_1958,N_14687,N_14728);
xor UO_1959 (O_1959,N_14553,N_14306);
nor UO_1960 (O_1960,N_14283,N_14881);
nand UO_1961 (O_1961,N_14386,N_14479);
nand UO_1962 (O_1962,N_14560,N_14118);
and UO_1963 (O_1963,N_14673,N_14506);
xnor UO_1964 (O_1964,N_14308,N_14060);
nor UO_1965 (O_1965,N_14006,N_14695);
nor UO_1966 (O_1966,N_14707,N_14962);
and UO_1967 (O_1967,N_14630,N_14364);
xor UO_1968 (O_1968,N_14014,N_14959);
nand UO_1969 (O_1969,N_14960,N_14910);
nor UO_1970 (O_1970,N_14449,N_14030);
and UO_1971 (O_1971,N_14440,N_14654);
nor UO_1972 (O_1972,N_14107,N_14295);
nor UO_1973 (O_1973,N_14712,N_14190);
or UO_1974 (O_1974,N_14121,N_14152);
and UO_1975 (O_1975,N_14925,N_14644);
xnor UO_1976 (O_1976,N_14799,N_14846);
and UO_1977 (O_1977,N_14446,N_14241);
xnor UO_1978 (O_1978,N_14038,N_14699);
and UO_1979 (O_1979,N_14311,N_14096);
nor UO_1980 (O_1980,N_14585,N_14758);
nor UO_1981 (O_1981,N_14074,N_14171);
or UO_1982 (O_1982,N_14209,N_14110);
xor UO_1983 (O_1983,N_14900,N_14201);
nand UO_1984 (O_1984,N_14588,N_14571);
xor UO_1985 (O_1985,N_14517,N_14535);
or UO_1986 (O_1986,N_14880,N_14552);
nor UO_1987 (O_1987,N_14620,N_14328);
and UO_1988 (O_1988,N_14411,N_14593);
nor UO_1989 (O_1989,N_14713,N_14231);
and UO_1990 (O_1990,N_14288,N_14630);
or UO_1991 (O_1991,N_14863,N_14890);
nand UO_1992 (O_1992,N_14994,N_14377);
xnor UO_1993 (O_1993,N_14085,N_14282);
xnor UO_1994 (O_1994,N_14352,N_14685);
xor UO_1995 (O_1995,N_14077,N_14215);
or UO_1996 (O_1996,N_14944,N_14846);
nor UO_1997 (O_1997,N_14423,N_14948);
xor UO_1998 (O_1998,N_14649,N_14075);
xnor UO_1999 (O_1999,N_14151,N_14921);
endmodule