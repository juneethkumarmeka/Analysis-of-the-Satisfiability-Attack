module basic_3000_30000_3500_60_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2946,In_2942);
nand U1 (N_1,In_814,In_1894);
and U2 (N_2,In_1457,In_139);
nand U3 (N_3,In_1020,In_623);
and U4 (N_4,In_2290,In_1587);
and U5 (N_5,In_2828,In_1550);
nor U6 (N_6,In_997,In_2575);
xnor U7 (N_7,In_772,In_1104);
nor U8 (N_8,In_2721,In_425);
nand U9 (N_9,In_829,In_1694);
nor U10 (N_10,In_1732,In_2028);
or U11 (N_11,In_2604,In_991);
or U12 (N_12,In_2882,In_2117);
and U13 (N_13,In_2211,In_608);
or U14 (N_14,In_1613,In_118);
and U15 (N_15,In_577,In_190);
and U16 (N_16,In_1944,In_638);
nor U17 (N_17,In_2042,In_1171);
or U18 (N_18,In_2159,In_1836);
or U19 (N_19,In_2876,In_2519);
nor U20 (N_20,In_1692,In_2657);
nor U21 (N_21,In_2983,In_1452);
and U22 (N_22,In_2294,In_2223);
and U23 (N_23,In_539,In_2201);
nor U24 (N_24,In_2792,In_169);
nand U25 (N_25,In_1342,In_1699);
nand U26 (N_26,In_2491,In_2477);
and U27 (N_27,In_1958,In_1541);
xor U28 (N_28,In_2600,In_360);
xor U29 (N_29,In_1771,In_1775);
and U30 (N_30,In_2923,In_74);
nor U31 (N_31,In_2426,In_1562);
and U32 (N_32,In_1768,In_2394);
or U33 (N_33,In_1461,In_2191);
and U34 (N_34,In_1950,In_2265);
nand U35 (N_35,In_602,In_1546);
nor U36 (N_36,In_150,In_1834);
xnor U37 (N_37,In_2027,In_678);
nand U38 (N_38,In_2267,In_610);
xor U39 (N_39,In_2398,In_2659);
nand U40 (N_40,In_1917,In_2019);
or U41 (N_41,In_36,In_1920);
nand U42 (N_42,In_2249,In_902);
nand U43 (N_43,In_2741,In_653);
nor U44 (N_44,In_1513,In_254);
nor U45 (N_45,In_69,In_498);
nor U46 (N_46,In_2081,In_1900);
and U47 (N_47,In_2718,In_667);
nor U48 (N_48,In_1828,In_2002);
or U49 (N_49,In_1747,In_480);
or U50 (N_50,In_2054,In_822);
and U51 (N_51,In_890,In_559);
nand U52 (N_52,In_2569,In_1782);
and U53 (N_53,In_1156,In_1510);
and U54 (N_54,In_2000,In_2768);
xor U55 (N_55,In_2092,In_905);
or U56 (N_56,In_2835,In_28);
and U57 (N_57,In_2839,In_2136);
nor U58 (N_58,In_1762,In_216);
and U59 (N_59,In_1619,In_736);
xnor U60 (N_60,In_2952,In_1890);
and U61 (N_61,In_2958,In_1903);
xnor U62 (N_62,In_1312,In_523);
xor U63 (N_63,In_2617,In_362);
nor U64 (N_64,In_1646,In_461);
xnor U65 (N_65,In_513,In_242);
and U66 (N_66,In_1435,In_2545);
or U67 (N_67,In_495,In_1751);
nor U68 (N_68,In_2816,In_2486);
xnor U69 (N_69,In_2182,In_1637);
nor U70 (N_70,In_131,In_1235);
nand U71 (N_71,In_2607,In_1796);
and U72 (N_72,In_1552,In_339);
xor U73 (N_73,In_1757,In_1942);
xnor U74 (N_74,In_1639,In_570);
and U75 (N_75,In_977,In_1412);
nand U76 (N_76,In_1248,In_2503);
xnor U77 (N_77,In_2367,In_1257);
nand U78 (N_78,In_89,In_2689);
nor U79 (N_79,In_2484,In_591);
xnor U80 (N_80,In_2467,In_200);
nand U81 (N_81,In_2628,In_2955);
nand U82 (N_82,In_21,In_1082);
or U83 (N_83,In_2242,In_961);
and U84 (N_84,In_2760,In_132);
xnor U85 (N_85,In_1889,In_1251);
and U86 (N_86,In_368,In_606);
or U87 (N_87,In_2720,In_2485);
nor U88 (N_88,In_527,In_2761);
and U89 (N_89,In_558,In_1945);
or U90 (N_90,In_1464,In_1309);
or U91 (N_91,In_301,In_2245);
or U92 (N_92,In_2570,In_1738);
nor U93 (N_93,In_2993,In_1574);
xor U94 (N_94,In_2091,In_1878);
nand U95 (N_95,In_1924,In_1350);
xnor U96 (N_96,In_913,In_1451);
nand U97 (N_97,In_705,In_2927);
xor U98 (N_98,In_1238,In_91);
nor U99 (N_99,In_1634,In_850);
nand U100 (N_100,In_2407,In_198);
nand U101 (N_101,In_2779,In_740);
nand U102 (N_102,In_304,In_411);
and U103 (N_103,In_128,In_928);
xor U104 (N_104,In_939,In_827);
nand U105 (N_105,In_552,In_77);
or U106 (N_106,In_2315,In_2547);
and U107 (N_107,In_792,In_1223);
or U108 (N_108,In_2346,In_2590);
nor U109 (N_109,In_2082,In_689);
and U110 (N_110,In_1706,In_371);
nand U111 (N_111,In_397,In_2125);
nor U112 (N_112,In_340,In_885);
nor U113 (N_113,In_1861,In_1946);
xor U114 (N_114,In_2798,In_2293);
nor U115 (N_115,In_1013,In_2241);
and U116 (N_116,In_2668,In_910);
and U117 (N_117,In_1977,In_305);
nor U118 (N_118,In_2038,In_1124);
nor U119 (N_119,In_1403,In_1315);
or U120 (N_120,In_2285,In_2014);
xor U121 (N_121,In_1602,In_2957);
nand U122 (N_122,In_2013,In_1860);
and U123 (N_123,In_988,In_1724);
nor U124 (N_124,In_572,In_2253);
or U125 (N_125,In_1839,In_1061);
nand U126 (N_126,In_289,In_2871);
nand U127 (N_127,In_1449,In_457);
nand U128 (N_128,In_2645,In_1189);
nor U129 (N_129,In_1126,In_2968);
and U130 (N_130,In_1794,In_2530);
xor U131 (N_131,In_418,In_993);
xor U132 (N_132,In_2465,In_1200);
nor U133 (N_133,In_1108,In_1532);
and U134 (N_134,In_2744,In_1190);
or U135 (N_135,In_807,In_497);
nor U136 (N_136,In_1623,In_1489);
or U137 (N_137,In_2234,In_2387);
or U138 (N_138,In_2115,In_1310);
xor U139 (N_139,In_847,In_1756);
or U140 (N_140,In_370,In_1129);
nor U141 (N_141,In_2279,In_1676);
nand U142 (N_142,In_1687,In_1501);
nor U143 (N_143,In_2706,In_2304);
nor U144 (N_144,In_982,In_2419);
nor U145 (N_145,In_600,In_87);
and U146 (N_146,In_2552,In_2655);
xnor U147 (N_147,In_920,In_1908);
and U148 (N_148,In_141,In_1499);
xor U149 (N_149,In_701,In_2787);
and U150 (N_150,In_126,In_2554);
xnor U151 (N_151,In_421,In_2155);
nor U152 (N_152,In_1640,In_1769);
nand U153 (N_153,In_1181,In_954);
nor U154 (N_154,In_1143,In_2749);
nand U155 (N_155,In_2203,In_679);
nand U156 (N_156,In_2624,In_180);
nand U157 (N_157,In_1659,In_1644);
and U158 (N_158,In_70,In_1657);
or U159 (N_159,In_2940,In_1853);
nor U160 (N_160,In_1217,In_1795);
or U161 (N_161,In_1130,In_2746);
nor U162 (N_162,In_2856,In_1247);
or U163 (N_163,In_1666,In_1517);
xor U164 (N_164,In_579,In_2058);
and U165 (N_165,In_2813,In_854);
nor U166 (N_166,In_2928,In_60);
or U167 (N_167,In_757,In_2152);
nand U168 (N_168,In_294,In_2646);
nor U169 (N_169,In_587,In_1547);
and U170 (N_170,In_2085,In_359);
or U171 (N_171,In_963,In_2239);
xor U172 (N_172,In_1231,In_2272);
nand U173 (N_173,In_1997,In_1446);
or U174 (N_174,In_1673,In_1516);
and U175 (N_175,In_6,In_119);
nand U176 (N_176,In_2475,In_823);
or U177 (N_177,In_1992,In_2289);
or U178 (N_178,In_303,In_2805);
or U179 (N_179,In_756,In_1714);
or U180 (N_180,In_983,In_181);
and U181 (N_181,In_1990,In_956);
nand U182 (N_182,In_2903,In_153);
or U183 (N_183,In_2306,In_2428);
and U184 (N_184,In_746,In_2822);
or U185 (N_185,In_350,In_2561);
nor U186 (N_186,In_1964,In_2049);
nor U187 (N_187,In_2218,In_2221);
nand U188 (N_188,In_2397,In_2202);
nor U189 (N_189,In_918,In_2260);
nor U190 (N_190,In_2521,In_329);
and U191 (N_191,In_2217,In_1617);
or U192 (N_192,In_955,In_1152);
nand U193 (N_193,In_1737,In_1936);
and U194 (N_194,In_2847,In_2841);
or U195 (N_195,In_1279,In_1344);
or U196 (N_196,In_899,In_848);
nor U197 (N_197,In_586,In_2179);
xnor U198 (N_198,In_2374,In_2581);
or U199 (N_199,In_2146,In_1222);
xnor U200 (N_200,In_2539,In_1357);
or U201 (N_201,In_1372,In_2379);
nor U202 (N_202,In_257,In_1470);
xor U203 (N_203,In_1649,In_117);
nor U204 (N_204,In_1028,In_990);
nor U205 (N_205,In_205,In_228);
nor U206 (N_206,In_1224,In_2074);
nand U207 (N_207,In_2551,In_1914);
xnor U208 (N_208,In_2943,In_1830);
nand U209 (N_209,In_2764,In_845);
nor U210 (N_210,In_778,In_2099);
or U211 (N_211,In_1386,In_332);
xnor U212 (N_212,In_2896,In_609);
or U213 (N_213,In_703,In_300);
and U214 (N_214,In_1493,In_103);
or U215 (N_215,In_531,In_1614);
and U216 (N_216,In_343,In_351);
and U217 (N_217,In_1987,In_1940);
nor U218 (N_218,In_1103,In_1184);
xor U219 (N_219,In_1101,In_466);
nor U220 (N_220,In_877,In_2535);
nand U221 (N_221,In_1093,In_2301);
or U222 (N_222,In_1744,In_225);
and U223 (N_223,In_809,In_1019);
and U224 (N_224,In_420,In_1728);
and U225 (N_225,In_67,In_64);
nor U226 (N_226,In_1948,In_31);
or U227 (N_227,In_2738,In_1500);
or U228 (N_228,In_2400,In_1007);
or U229 (N_229,In_2436,In_2883);
or U230 (N_230,In_1039,In_344);
nor U231 (N_231,In_1555,In_723);
and U232 (N_232,In_611,In_563);
and U233 (N_233,In_2901,In_590);
or U234 (N_234,In_475,In_794);
nor U235 (N_235,In_1817,In_2464);
nand U236 (N_236,In_1674,In_2781);
xor U237 (N_237,In_2132,In_909);
nand U238 (N_238,In_2015,In_27);
and U239 (N_239,In_2908,In_2586);
or U240 (N_240,In_540,In_1742);
and U241 (N_241,In_1332,In_575);
nor U242 (N_242,In_1813,In_2442);
and U243 (N_243,In_1067,In_852);
and U244 (N_244,In_2715,In_2382);
or U245 (N_245,In_2853,In_1076);
nand U246 (N_246,In_1201,In_1943);
and U247 (N_247,In_2196,In_2754);
nand U248 (N_248,In_2817,In_2994);
or U249 (N_249,In_336,In_2748);
nor U250 (N_250,In_333,In_2498);
nand U251 (N_251,In_1041,In_2704);
or U252 (N_252,In_999,In_926);
nand U253 (N_253,In_2594,In_241);
xor U254 (N_254,In_2560,In_1349);
nand U255 (N_255,In_2640,In_448);
and U256 (N_256,In_2696,In_866);
or U257 (N_257,In_2243,In_263);
nor U258 (N_258,In_33,In_830);
or U259 (N_259,In_2821,In_585);
nor U260 (N_260,In_2341,In_1970);
nand U261 (N_261,In_1654,In_541);
and U262 (N_262,In_974,In_208);
nor U263 (N_263,In_2589,In_2662);
or U264 (N_264,In_1427,In_726);
xor U265 (N_265,In_642,In_2855);
or U266 (N_266,In_951,In_54);
or U267 (N_267,In_1981,In_1884);
or U268 (N_268,In_1198,In_2598);
nor U269 (N_269,In_1281,In_581);
and U270 (N_270,In_1301,In_2088);
and U271 (N_271,In_477,In_1080);
nand U272 (N_272,In_1647,In_1818);
nor U273 (N_273,In_1568,In_2080);
nor U274 (N_274,In_1854,In_412);
and U275 (N_275,In_1492,In_433);
nor U276 (N_276,In_1572,In_769);
xnor U277 (N_277,In_2086,In_693);
and U278 (N_278,In_2172,In_2313);
and U279 (N_279,In_960,In_1034);
or U280 (N_280,In_2330,In_688);
or U281 (N_281,In_2558,In_2750);
and U282 (N_282,In_385,In_2611);
or U283 (N_283,In_1638,In_493);
xnor U284 (N_284,In_2613,In_565);
xnor U285 (N_285,In_422,In_2897);
nor U286 (N_286,In_1829,In_2636);
xor U287 (N_287,In_2700,In_2408);
nor U288 (N_288,In_1123,In_2216);
nand U289 (N_289,In_2145,In_1088);
or U290 (N_290,In_2056,In_2134);
xor U291 (N_291,In_470,In_2045);
or U292 (N_292,In_1874,In_553);
xor U293 (N_293,In_1815,In_178);
xor U294 (N_294,In_1968,In_1428);
nand U295 (N_295,In_799,In_1661);
and U296 (N_296,In_1481,In_1688);
xor U297 (N_297,In_700,In_1474);
nand U298 (N_298,In_979,In_1);
nor U299 (N_299,In_218,In_834);
or U300 (N_300,In_583,In_825);
xor U301 (N_301,In_2810,In_544);
nand U302 (N_302,In_2990,In_2893);
nand U303 (N_303,In_2735,In_147);
xnor U304 (N_304,In_2536,In_784);
xnor U305 (N_305,In_1083,In_2405);
nor U306 (N_306,In_215,In_2222);
or U307 (N_307,In_273,In_1910);
and U308 (N_308,In_1099,In_2880);
nand U309 (N_309,In_1164,In_2999);
and U310 (N_310,In_1741,In_2184);
nor U311 (N_311,In_2830,In_2232);
nand U312 (N_312,In_2466,In_1901);
or U313 (N_313,In_2282,In_184);
xnor U314 (N_314,In_1004,In_408);
or U315 (N_315,In_2197,In_1042);
nor U316 (N_316,In_904,In_1467);
xor U317 (N_317,In_2380,In_859);
and U318 (N_318,In_282,In_671);
xnor U319 (N_319,In_1823,In_719);
and U320 (N_320,In_2017,In_1869);
or U321 (N_321,In_2723,In_1808);
or U322 (N_322,In_1632,In_2854);
xor U323 (N_323,In_1790,In_24);
xnor U324 (N_324,In_2432,In_1194);
nor U325 (N_325,In_2283,In_1746);
and U326 (N_326,In_545,In_2334);
xor U327 (N_327,In_1105,In_790);
nand U328 (N_328,In_389,In_1003);
or U329 (N_329,In_165,In_2641);
or U330 (N_330,In_251,In_1537);
or U331 (N_331,In_255,In_2256);
and U332 (N_332,In_2194,In_2210);
nor U333 (N_333,In_1440,In_808);
or U334 (N_334,In_1701,In_2453);
xnor U335 (N_335,In_1469,In_2769);
or U336 (N_336,In_2010,In_1402);
xnor U337 (N_337,In_646,In_187);
nor U338 (N_338,In_1681,In_2292);
nand U339 (N_339,In_2699,In_1036);
and U340 (N_340,In_1814,In_683);
nor U341 (N_341,In_392,In_1662);
nand U342 (N_342,In_2469,In_1849);
and U343 (N_343,In_2571,In_1952);
nor U344 (N_344,In_1340,In_53);
nor U345 (N_345,In_1407,In_2076);
xor U346 (N_346,In_636,In_1641);
or U347 (N_347,In_1557,In_2568);
nand U348 (N_348,In_806,In_2360);
nor U349 (N_349,In_2538,In_1278);
nand U350 (N_350,In_959,In_1437);
nand U351 (N_351,In_157,In_1838);
xor U352 (N_352,In_2980,In_2310);
nor U353 (N_353,In_1573,In_485);
xor U354 (N_354,In_797,In_1148);
nand U355 (N_355,In_2,In_1447);
or U356 (N_356,In_2574,In_2643);
nor U357 (N_357,In_1436,In_1106);
and U358 (N_358,In_1218,In_1705);
xnor U359 (N_359,In_980,In_2349);
nor U360 (N_360,In_906,In_1636);
and U361 (N_361,In_83,In_68);
and U362 (N_362,In_2299,In_1678);
and U363 (N_363,In_2358,In_2176);
xnor U364 (N_364,In_1043,In_2556);
nand U365 (N_365,In_2348,In_897);
nand U366 (N_366,In_938,In_13);
nand U367 (N_367,In_1454,In_1972);
xnor U368 (N_368,In_1690,In_1431);
and U369 (N_369,In_1348,In_1718);
or U370 (N_370,In_2122,In_1298);
and U371 (N_371,In_1507,In_1091);
and U372 (N_372,In_774,In_1057);
and U373 (N_373,In_1249,In_2458);
nand U374 (N_374,In_2438,In_1424);
and U375 (N_375,In_366,In_2799);
nand U376 (N_376,In_2963,In_1341);
nor U377 (N_377,In_2127,In_2288);
xor U378 (N_378,In_1928,In_620);
and U379 (N_379,In_2147,In_455);
xor U380 (N_380,In_1095,In_342);
and U381 (N_381,In_2333,In_2418);
and U382 (N_382,In_443,In_464);
or U383 (N_383,In_372,In_501);
or U384 (N_384,In_1376,In_1158);
or U385 (N_385,In_2580,In_684);
xnor U386 (N_386,In_2845,In_1685);
nor U387 (N_387,In_534,In_839);
nor U388 (N_388,In_2863,In_2667);
xnor U389 (N_389,In_2430,In_2342);
and U390 (N_390,In_1355,In_765);
or U391 (N_391,In_2311,In_1269);
xor U392 (N_392,In_650,In_1660);
and U393 (N_393,In_1102,In_1518);
xnor U394 (N_394,In_1448,In_1622);
nand U395 (N_395,In_1712,In_142);
or U396 (N_396,In_836,In_840);
nand U397 (N_397,In_410,In_1938);
or U398 (N_398,In_279,In_950);
nor U399 (N_399,In_1986,In_1618);
xnor U400 (N_400,In_2046,In_987);
xor U401 (N_401,In_1965,In_1571);
nor U402 (N_402,In_763,In_2075);
or U403 (N_403,In_2785,In_1022);
nor U404 (N_404,In_1385,In_404);
or U405 (N_405,In_1107,In_2673);
and U406 (N_406,In_1271,In_1761);
nor U407 (N_407,In_2627,In_1593);
and U408 (N_408,In_1717,In_675);
and U409 (N_409,In_1016,In_2261);
xor U410 (N_410,In_1722,In_260);
nand U411 (N_411,In_733,In_2052);
nand U412 (N_412,In_1534,In_2869);
or U413 (N_413,In_2331,In_2368);
xor U414 (N_414,In_1859,In_1822);
nand U415 (N_415,In_2236,In_19);
and U416 (N_416,In_1065,In_821);
xnor U417 (N_417,In_2274,In_2039);
nand U418 (N_418,In_969,In_2730);
and U419 (N_419,In_2717,In_503);
xor U420 (N_420,In_1825,In_2937);
or U421 (N_421,In_681,In_2492);
nor U422 (N_422,In_376,In_917);
xor U423 (N_423,In_2296,In_211);
and U424 (N_424,In_1212,In_547);
nor U425 (N_425,In_931,In_1135);
nor U426 (N_426,In_102,In_1726);
or U427 (N_427,In_214,In_127);
or U428 (N_428,In_633,In_520);
or U429 (N_429,In_2804,In_1170);
nand U430 (N_430,In_724,In_2174);
or U431 (N_431,In_2369,In_1912);
or U432 (N_432,In_601,In_1925);
xnor U433 (N_433,In_1697,In_2634);
xnor U434 (N_434,In_2685,In_1951);
nand U435 (N_435,In_1872,In_1276);
nand U436 (N_436,In_2148,In_2762);
nand U437 (N_437,In_1476,In_2139);
or U438 (N_438,In_1117,In_901);
and U439 (N_439,In_1754,In_1580);
nor U440 (N_440,In_2716,In_2631);
and U441 (N_441,In_915,In_1883);
nand U442 (N_442,In_518,In_120);
nand U443 (N_443,In_2237,In_173);
nand U444 (N_444,In_2135,In_323);
or U445 (N_445,In_2650,In_2276);
or U446 (N_446,In_499,In_2169);
or U447 (N_447,In_472,In_2513);
xor U448 (N_448,In_2593,In_1277);
nand U449 (N_449,In_2945,In_1655);
xnor U450 (N_450,In_2988,In_986);
nor U451 (N_451,In_1337,In_1820);
nor U452 (N_452,In_2064,In_800);
nand U453 (N_453,In_451,In_1085);
and U454 (N_454,In_1700,In_2248);
nor U455 (N_455,In_2991,In_1031);
xor U456 (N_456,In_2029,In_1536);
and U457 (N_457,In_1882,In_1731);
nand U458 (N_458,In_1014,In_320);
nor U459 (N_459,In_43,In_2860);
nand U460 (N_460,In_1664,In_2066);
and U461 (N_461,In_2073,In_1120);
or U462 (N_462,In_1675,In_2363);
nand U463 (N_463,In_994,In_1038);
nand U464 (N_464,In_1183,In_1259);
and U465 (N_465,In_685,In_2193);
xnor U466 (N_466,In_1913,In_1002);
xnor U467 (N_467,In_872,In_2336);
and U468 (N_468,In_729,In_2916);
nand U469 (N_469,In_56,In_364);
nor U470 (N_470,In_548,In_213);
and U471 (N_471,In_232,In_863);
xor U472 (N_472,In_2703,In_1442);
xnor U473 (N_473,In_1368,In_1347);
xor U474 (N_474,In_1953,In_1245);
nor U475 (N_475,In_1543,In_2361);
xnor U476 (N_476,In_1365,In_682);
nand U477 (N_477,In_1311,In_584);
and U478 (N_478,In_643,In_2941);
and U479 (N_479,In_2370,In_648);
or U480 (N_480,In_1564,In_2675);
nor U481 (N_481,In_2280,In_2250);
nor U482 (N_482,In_1186,In_2771);
nor U483 (N_483,In_349,In_2743);
and U484 (N_484,In_8,In_2584);
and U485 (N_485,In_761,In_1356);
nand U486 (N_486,In_1073,In_932);
nand U487 (N_487,In_615,In_2411);
nor U488 (N_488,In_652,In_1591);
and U489 (N_489,In_738,In_1246);
or U490 (N_490,In_9,In_875);
nand U491 (N_491,In_2837,In_660);
xnor U492 (N_492,In_2344,In_869);
and U493 (N_493,In_1127,In_2339);
or U494 (N_494,In_138,In_1497);
nand U495 (N_495,In_2006,In_2016);
nand U496 (N_496,In_2907,In_1515);
nor U497 (N_497,In_1213,In_2262);
nand U498 (N_498,In_2694,In_2376);
and U499 (N_499,In_535,In_912);
xnor U500 (N_500,N_287,In_1628);
nor U501 (N_501,In_1096,In_2653);
and U502 (N_502,In_116,N_463);
nand U503 (N_503,In_2546,In_1561);
nand U504 (N_504,In_2295,In_1907);
and U505 (N_505,In_1539,In_2499);
or U506 (N_506,N_102,N_373);
nor U507 (N_507,In_1202,In_2585);
nand U508 (N_508,In_2032,In_2707);
nor U509 (N_509,In_2372,In_2563);
and U510 (N_510,N_409,In_1509);
nor U511 (N_511,In_2124,N_407);
or U512 (N_512,In_2864,In_2071);
xor U513 (N_513,N_110,In_101);
and U514 (N_514,In_1159,In_110);
xor U515 (N_515,In_2229,In_1300);
nor U516 (N_516,In_459,In_1265);
xnor U517 (N_517,In_629,In_1033);
nand U518 (N_518,In_2482,In_2501);
or U519 (N_519,In_1115,In_1313);
nor U520 (N_520,In_2224,In_2371);
or U521 (N_521,N_90,N_331);
xnor U522 (N_522,In_1582,In_2388);
xnor U523 (N_523,In_1892,In_1141);
and U524 (N_524,N_365,In_2303);
nor U525 (N_525,In_1144,In_390);
xnor U526 (N_526,In_1037,In_1377);
and U527 (N_527,In_833,In_1339);
xnor U528 (N_528,In_2133,In_1495);
xnor U529 (N_529,In_298,In_1001);
or U530 (N_530,In_226,In_1113);
and U531 (N_531,In_949,In_849);
or U532 (N_532,In_2808,In_860);
or U533 (N_533,In_488,In_237);
and U534 (N_534,In_802,In_222);
xnor U535 (N_535,In_662,In_2131);
xor U536 (N_536,In_166,In_2647);
or U537 (N_537,N_495,In_654);
xor U538 (N_538,N_311,In_714);
and U539 (N_539,N_475,In_944);
nand U540 (N_540,In_874,In_1563);
nor U541 (N_541,N_45,In_2981);
or U542 (N_542,In_352,In_2527);
nand U543 (N_543,In_2770,In_2051);
xnor U544 (N_544,In_1934,In_299);
nand U545 (N_545,In_134,In_2975);
or U546 (N_546,N_138,In_957);
nand U547 (N_547,In_460,In_306);
nor U548 (N_548,N_489,In_1226);
and U549 (N_549,In_1153,In_312);
nor U550 (N_550,In_1199,N_298);
and U551 (N_551,N_57,In_707);
or U552 (N_552,In_842,In_1401);
or U553 (N_553,In_1978,In_1157);
xor U554 (N_554,In_229,In_1203);
or U555 (N_555,In_1783,In_1668);
and U556 (N_556,In_2098,In_483);
xor U557 (N_557,N_472,In_1326);
and U558 (N_558,In_1351,In_1219);
nand U559 (N_559,In_691,In_290);
xor U560 (N_560,In_2576,In_2434);
and U561 (N_561,In_695,In_1801);
nand U562 (N_562,In_1615,In_1955);
or U563 (N_563,N_385,In_1327);
nand U564 (N_564,N_265,In_314);
xor U565 (N_565,N_256,N_157);
xnor U566 (N_566,N_51,In_2077);
nor U567 (N_567,N_127,In_307);
and U568 (N_568,In_1262,In_356);
and U569 (N_569,N_307,In_296);
or U570 (N_570,In_2246,In_1071);
nor U571 (N_571,In_1514,N_69);
nand U572 (N_572,N_336,In_1529);
nand U573 (N_573,In_526,In_1650);
nand U574 (N_574,N_56,In_2338);
nor U575 (N_575,In_2270,N_438);
or U576 (N_576,In_2938,N_167);
and U577 (N_577,N_27,In_1139);
or U578 (N_578,In_992,In_186);
nor U579 (N_579,In_1288,In_494);
xor U580 (N_580,In_921,In_238);
and U581 (N_581,In_597,In_1902);
xor U582 (N_582,N_24,In_2141);
and U583 (N_583,In_1263,N_181);
or U584 (N_584,In_783,In_330);
xor U585 (N_585,In_1270,In_1704);
or U586 (N_586,N_126,In_2452);
nand U587 (N_587,In_605,In_831);
and U588 (N_588,In_1331,N_338);
nand U589 (N_589,In_1961,N_481);
nor U590 (N_590,In_1294,In_1011);
nor U591 (N_591,In_887,In_1922);
nor U592 (N_592,In_1137,In_2450);
or U593 (N_593,In_315,In_1715);
and U594 (N_594,In_1252,In_1648);
or U595 (N_595,N_252,In_309);
nand U596 (N_596,In_536,In_554);
nand U597 (N_597,In_1840,In_1378);
xor U598 (N_598,In_246,In_771);
xnor U599 (N_599,In_907,In_1173);
nand U600 (N_600,In_151,In_500);
nand U601 (N_601,In_658,In_2233);
or U602 (N_602,In_2271,In_1072);
xnor U603 (N_603,N_43,In_2541);
and U604 (N_604,In_171,In_439);
xor U605 (N_605,N_372,In_1522);
xnor U606 (N_606,In_2597,In_739);
and U607 (N_607,In_2067,In_998);
xor U608 (N_608,In_2702,In_702);
and U609 (N_609,In_2284,In_432);
xor U610 (N_610,In_25,N_70);
or U611 (N_611,In_1957,In_172);
xnor U612 (N_612,In_855,In_2113);
or U613 (N_613,In_2788,In_2121);
and U614 (N_614,In_1723,In_1525);
and U615 (N_615,In_403,In_244);
nand U616 (N_616,In_621,In_2266);
or U617 (N_617,In_2448,In_1284);
nor U618 (N_618,In_1805,In_233);
nor U619 (N_619,In_130,N_74);
and U620 (N_620,N_299,In_853);
or U621 (N_621,In_745,In_2683);
or U622 (N_622,In_937,In_936);
xor U623 (N_623,In_2933,In_2329);
and U624 (N_624,N_268,In_1484);
xnor U625 (N_625,In_2778,In_491);
xnor U626 (N_626,N_149,In_2413);
and U627 (N_627,In_2462,N_384);
xnor U628 (N_628,In_1635,N_168);
nand U629 (N_629,N_326,In_2228);
nor U630 (N_630,In_640,In_2710);
xnor U631 (N_631,In_1078,In_363);
nor U632 (N_632,N_413,In_2268);
xnor U633 (N_633,In_1185,In_2192);
and U634 (N_634,In_2567,In_2591);
nand U635 (N_635,In_560,In_85);
and U636 (N_636,In_272,In_221);
and U637 (N_637,In_1975,In_1374);
nor U638 (N_638,In_145,In_857);
or U639 (N_639,In_1243,In_430);
and U640 (N_640,In_1904,In_1371);
nand U641 (N_641,In_159,In_2850);
nor U642 (N_642,In_2533,In_487);
and U643 (N_643,N_20,In_2020);
xnor U644 (N_644,In_297,In_1630);
nor U645 (N_645,In_1394,In_2920);
or U646 (N_646,In_2507,In_659);
or U647 (N_647,In_1994,In_427);
or U648 (N_648,In_1542,In_2472);
xnor U649 (N_649,In_2402,In_941);
and U650 (N_650,In_2381,In_1875);
nor U651 (N_651,In_1755,In_2140);
nor U652 (N_652,In_1478,In_935);
xor U653 (N_653,In_1527,In_409);
nand U654 (N_654,In_1063,In_1691);
or U655 (N_655,In_561,N_35);
and U656 (N_656,In_1491,In_2737);
and U657 (N_657,In_1919,N_144);
nor U658 (N_658,In_1121,N_253);
xnor U659 (N_659,In_1982,In_167);
and U660 (N_660,In_2751,In_1128);
or U661 (N_661,In_154,N_408);
nand U662 (N_662,In_1979,In_883);
xor U663 (N_663,In_1005,In_2512);
and U664 (N_664,In_2399,In_248);
nand U665 (N_665,In_2949,In_533);
and U666 (N_666,In_1373,N_211);
nand U667 (N_667,In_1743,In_287);
nand U668 (N_668,N_204,N_14);
or U669 (N_669,In_731,In_49);
or U670 (N_670,In_1482,In_777);
and U671 (N_671,In_162,In_2714);
xor U672 (N_672,In_1472,In_2396);
nand U673 (N_673,In_2162,In_2978);
or U674 (N_674,N_369,In_1779);
nand U675 (N_675,In_2103,In_881);
or U676 (N_676,In_1214,N_223);
or U677 (N_677,N_60,In_1530);
and U678 (N_678,N_275,In_476);
xnor U679 (N_679,In_1379,N_478);
and U680 (N_680,In_437,In_2324);
nand U681 (N_681,In_2726,N_9);
or U682 (N_682,In_889,In_1857);
xor U683 (N_683,In_984,In_1012);
xor U684 (N_684,In_2820,N_62);
nand U685 (N_685,In_313,N_228);
xor U686 (N_686,N_269,In_188);
and U687 (N_687,In_2154,In_1600);
nor U688 (N_688,In_2724,In_1989);
or U689 (N_689,N_75,In_555);
nand U690 (N_690,In_2354,In_2806);
and U691 (N_691,In_811,In_1387);
nand U692 (N_692,N_231,In_1404);
or U693 (N_693,N_163,In_1798);
nor U694 (N_694,In_1066,In_2843);
nand U695 (N_695,In_846,In_1897);
xor U696 (N_696,N_257,In_1466);
xnor U697 (N_697,In_2391,In_413);
nor U698 (N_698,N_278,N_303);
nor U699 (N_699,In_48,In_781);
and U700 (N_700,In_1134,In_1545);
and U701 (N_701,In_1531,In_844);
or U702 (N_702,N_414,In_1196);
or U703 (N_703,In_1000,In_759);
or U704 (N_704,N_366,In_2913);
and U705 (N_705,In_234,N_363);
or U706 (N_706,In_2157,In_2979);
or U707 (N_707,In_1776,N_440);
xor U708 (N_708,In_2649,N_428);
or U709 (N_709,N_476,In_149);
nand U710 (N_710,N_347,N_166);
and U711 (N_711,In_1026,In_1443);
xor U712 (N_712,In_249,In_1504);
and U713 (N_713,In_2620,In_2395);
or U714 (N_714,In_2582,In_884);
xor U715 (N_715,In_2024,In_2158);
xnor U716 (N_716,In_1730,In_1122);
xnor U717 (N_717,In_1353,N_474);
nand U718 (N_718,In_2161,N_54);
nor U719 (N_719,In_2404,In_1993);
and U720 (N_720,In_361,In_2410);
and U721 (N_721,In_2522,N_280);
nor U722 (N_722,In_2904,In_474);
and U723 (N_723,N_4,In_1578);
nand U724 (N_724,In_2691,In_2713);
nand U725 (N_725,In_353,N_189);
and U726 (N_726,In_743,N_66);
nand U727 (N_727,In_2681,In_1318);
and U728 (N_728,In_109,In_1075);
xnor U729 (N_729,In_111,In_712);
nor U730 (N_730,In_2890,In_1605);
xor U731 (N_731,N_258,In_2891);
xor U732 (N_732,N_431,In_59);
xnor U733 (N_733,In_122,In_245);
or U734 (N_734,In_377,In_2287);
and U735 (N_735,In_2198,N_342);
xnor U736 (N_736,N_415,In_1672);
nand U737 (N_737,N_283,In_2630);
nand U738 (N_738,In_2220,N_488);
nand U739 (N_739,N_44,In_2997);
xor U740 (N_740,In_1753,N_281);
nor U741 (N_741,N_421,In_1323);
xor U742 (N_742,In_1886,N_18);
xnor U743 (N_743,N_263,In_1162);
xnor U744 (N_744,In_1160,In_1592);
nor U745 (N_745,In_2661,In_2719);
nor U746 (N_746,In_414,N_249);
nor U747 (N_747,In_2572,In_1295);
nor U748 (N_748,In_2678,In_2431);
nor U749 (N_749,In_176,In_47);
and U750 (N_750,In_880,In_1100);
nand U751 (N_751,N_404,N_175);
nor U752 (N_752,In_2809,In_1533);
xor U753 (N_753,In_1025,In_1802);
xnor U754 (N_754,In_1791,In_1810);
nor U755 (N_755,In_1209,In_2953);
and U756 (N_756,In_2742,In_2866);
or U757 (N_757,In_2414,In_613);
nor U758 (N_758,N_100,In_1689);
xnor U759 (N_759,In_278,In_1052);
nand U760 (N_760,In_1058,In_1995);
or U761 (N_761,N_71,In_1680);
nand U762 (N_762,In_677,In_713);
nor U763 (N_763,In_2496,In_780);
and U764 (N_764,In_2126,In_2666);
nor U765 (N_765,In_2018,In_2831);
nand U766 (N_766,In_1187,In_2429);
or U767 (N_767,In_2959,In_2884);
xnor U768 (N_768,N_47,In_321);
or U769 (N_769,In_1346,In_2107);
xnor U770 (N_770,In_2143,In_2954);
or U771 (N_771,In_1145,In_1398);
and U772 (N_772,In_1788,In_2297);
nand U773 (N_773,N_418,In_2852);
xnor U774 (N_774,N_273,In_2323);
and U775 (N_775,In_2178,In_886);
xor U776 (N_776,In_1208,In_1523);
nor U777 (N_777,In_2326,In_354);
or U778 (N_778,In_1475,In_2902);
nand U779 (N_779,N_241,In_1054);
and U780 (N_780,In_492,In_295);
and U781 (N_781,In_1967,N_350);
nor U782 (N_782,In_2417,In_1866);
nor U783 (N_783,N_430,In_625);
nor U784 (N_784,In_2509,N_316);
nand U785 (N_785,N_272,In_1565);
xnor U786 (N_786,In_2097,N_453);
xnor U787 (N_787,In_426,In_202);
xnor U788 (N_788,In_1577,In_2797);
and U789 (N_789,In_871,In_206);
and U790 (N_790,In_2671,N_88);
and U791 (N_791,In_2939,In_2328);
and U792 (N_792,In_1056,In_1059);
xnor U793 (N_793,In_319,In_23);
xor U794 (N_794,N_445,In_529);
nor U795 (N_795,In_1959,In_1848);
and U796 (N_796,In_1150,In_2269);
and U797 (N_797,N_86,In_568);
nor U798 (N_798,N_254,In_2516);
or U799 (N_799,In_1999,In_2105);
nor U800 (N_800,N_461,In_1881);
nand U801 (N_801,N_295,In_1154);
xnor U802 (N_802,In_2606,In_20);
nand U803 (N_803,In_135,N_262);
or U804 (N_804,N_364,In_2393);
and U805 (N_805,In_2149,In_10);
nor U806 (N_806,In_773,In_280);
or U807 (N_807,In_1188,In_2114);
and U808 (N_808,In_1793,N_134);
nor U809 (N_809,In_728,In_1506);
nand U810 (N_810,In_2007,In_891);
xor U811 (N_811,In_2443,N_349);
nor U812 (N_812,N_215,N_226);
or U813 (N_813,In_1806,N_190);
nand U814 (N_814,N_115,In_1405);
and U815 (N_815,In_2062,In_1268);
nand U816 (N_816,In_895,In_1287);
or U817 (N_817,In_1426,In_155);
nand U818 (N_818,In_2622,In_898);
nor U819 (N_819,In_367,In_634);
xor U820 (N_820,In_1807,In_1477);
nand U821 (N_821,In_447,In_1745);
and U822 (N_822,In_1610,In_35);
nand U823 (N_823,In_514,In_1179);
nand U824 (N_824,In_1833,In_379);
or U825 (N_825,In_1140,In_230);
nand U826 (N_826,In_1369,N_128);
nor U827 (N_827,In_2680,In_311);
nor U828 (N_828,In_2180,In_1596);
nor U829 (N_829,In_199,In_1111);
nor U830 (N_830,In_1670,In_2595);
and U831 (N_831,In_1799,In_1254);
xor U832 (N_832,N_146,In_843);
or U833 (N_833,In_2605,In_696);
or U834 (N_834,In_2824,In_80);
or U835 (N_835,In_2050,In_2621);
xor U836 (N_836,In_2138,In_310);
nor U837 (N_837,In_947,In_2573);
or U838 (N_838,In_1237,In_265);
and U839 (N_839,In_2508,In_90);
and U840 (N_840,In_1891,In_571);
xor U841 (N_841,In_203,In_2037);
and U842 (N_842,In_2078,In_1558);
xor U843 (N_843,In_1710,In_2961);
nor U844 (N_844,N_6,In_1486);
nand U845 (N_845,In_2861,In_2670);
or U846 (N_846,In_1415,N_277);
nor U847 (N_847,In_1393,N_294);
and U848 (N_848,N_68,In_189);
nand U849 (N_849,In_2386,In_1624);
or U850 (N_850,In_793,In_2034);
nand U851 (N_851,In_2842,In_968);
nor U852 (N_852,In_2345,In_1774);
or U853 (N_853,In_2868,In_1831);
nand U854 (N_854,N_87,In_2108);
or U855 (N_855,In_1954,In_1364);
nand U856 (N_856,In_1060,In_175);
xor U857 (N_857,In_65,In_268);
nand U858 (N_858,In_1215,In_2375);
or U859 (N_859,In_1709,N_447);
nor U860 (N_860,In_2259,In_29);
nand U861 (N_861,In_2185,In_2204);
and U862 (N_862,In_291,In_828);
nand U863 (N_863,N_293,In_2766);
nor U864 (N_864,In_274,In_2555);
nor U865 (N_865,In_2247,In_1367);
xnor U866 (N_866,In_753,In_108);
or U867 (N_867,In_1851,In_38);
and U868 (N_868,In_1971,In_104);
nor U869 (N_869,N_1,In_882);
or U870 (N_870,In_870,In_1210);
nand U871 (N_871,N_227,In_1459);
xor U872 (N_872,N_383,In_1366);
or U873 (N_873,In_489,In_465);
and U874 (N_874,In_1465,N_72);
or U875 (N_875,In_1785,In_308);
xnor U876 (N_876,In_1607,In_191);
nor U877 (N_877,N_360,In_1138);
xnor U878 (N_878,N_492,N_98);
nand U879 (N_879,In_1463,In_26);
nand U880 (N_880,In_923,In_1422);
or U881 (N_881,In_1055,In_2800);
or U882 (N_882,In_2065,In_335);
xnor U883 (N_883,In_1334,In_1777);
and U884 (N_884,In_1759,In_2947);
nand U885 (N_885,In_160,In_2190);
nor U886 (N_886,In_1711,In_2364);
xnor U887 (N_887,In_1521,In_2129);
xnor U888 (N_888,In_929,In_398);
nor U889 (N_889,In_428,In_2454);
xor U890 (N_890,In_30,N_242);
and U891 (N_891,In_556,In_2531);
or U892 (N_892,N_483,In_1274);
xor U893 (N_893,In_2109,In_801);
xor U894 (N_894,In_334,In_1230);
nor U895 (N_895,In_185,In_2633);
xor U896 (N_896,In_1816,In_2832);
nand U897 (N_897,In_2275,In_325);
or U898 (N_898,In_2925,In_240);
nand U899 (N_899,In_952,In_125);
xor U900 (N_900,In_2948,N_305);
and U901 (N_901,In_2878,In_1758);
and U902 (N_902,N_313,In_2325);
and U903 (N_903,In_1842,In_219);
nor U904 (N_904,In_1929,In_2340);
or U905 (N_905,N_358,In_2892);
or U906 (N_906,N_5,In_2163);
nand U907 (N_907,In_2263,In_1733);
nor U908 (N_908,In_1077,In_2789);
nand U909 (N_909,In_2780,In_1868);
nor U910 (N_910,In_1253,In_2377);
or U911 (N_911,N_270,In_815);
nand U912 (N_912,In_2116,N_203);
nor U913 (N_913,N_370,In_2231);
and U914 (N_914,In_235,In_598);
nand U915 (N_915,N_21,In_383);
or U916 (N_916,In_741,In_1819);
xor U917 (N_917,In_1703,N_155);
and U918 (N_918,In_2069,In_985);
nor U919 (N_919,In_1266,In_509);
and U920 (N_920,In_1225,In_1414);
or U921 (N_921,N_3,In_1023);
or U922 (N_922,In_1827,In_2815);
xor U923 (N_923,In_1406,In_2188);
xnor U924 (N_924,In_2008,N_210);
xor U925 (N_925,N_426,In_704);
nor U926 (N_926,In_1876,In_207);
or U927 (N_927,In_2698,In_715);
nor U928 (N_928,In_1053,In_1719);
nand U929 (N_929,In_1166,In_2506);
nand U930 (N_930,In_196,N_133);
and U931 (N_931,In_1767,In_76);
nor U932 (N_932,In_1974,In_2905);
nand U933 (N_933,In_2300,In_2213);
and U934 (N_934,In_152,In_749);
xnor U935 (N_935,In_1168,In_158);
xor U936 (N_936,N_135,In_1244);
nand U937 (N_937,In_2663,In_1304);
or U938 (N_938,In_39,In_2565);
and U939 (N_939,N_145,In_209);
or U940 (N_940,In_2373,In_2934);
nor U941 (N_941,In_976,In_981);
or U942 (N_942,In_1296,N_197);
or U943 (N_943,In_2312,In_588);
or U944 (N_944,In_1865,In_973);
nor U945 (N_945,N_398,N_130);
or U946 (N_946,In_522,In_2235);
or U947 (N_947,N_174,In_435);
or U948 (N_948,In_2461,In_1239);
xor U949 (N_949,In_2120,N_132);
nand U950 (N_950,In_721,In_2094);
nor U951 (N_951,In_2827,In_71);
and U952 (N_952,In_2425,N_490);
nand U953 (N_953,N_46,In_1576);
and U954 (N_954,In_2875,N_225);
nand U955 (N_955,In_2935,In_2862);
and U956 (N_956,In_1887,In_328);
nand U957 (N_957,In_2238,In_2592);
nand U958 (N_958,In_2777,In_2041);
or U959 (N_959,In_816,In_1146);
nand U960 (N_960,In_1177,In_2872);
xor U961 (N_961,N_39,N_467);
and U962 (N_962,In_1192,N_33);
nand U963 (N_963,In_711,In_2060);
nand U964 (N_964,In_1286,In_384);
nor U965 (N_965,In_1683,In_506);
and U966 (N_966,In_1490,In_168);
nor U967 (N_967,In_61,In_324);
or U968 (N_968,In_2776,N_381);
xnor U969 (N_969,In_1735,N_341);
xor U970 (N_970,In_1438,In_1667);
nor U971 (N_971,N_217,N_229);
xnor U972 (N_972,N_122,In_551);
or U973 (N_973,In_2343,In_2965);
and U974 (N_974,N_171,In_1642);
xor U975 (N_975,In_2350,In_284);
nor U976 (N_976,In_687,In_2460);
xor U977 (N_977,In_2012,In_1425);
or U978 (N_978,In_1133,In_1413);
and U979 (N_979,In_197,In_2909);
nor U980 (N_980,In_1010,In_1255);
nor U981 (N_981,N_351,In_2969);
and U982 (N_982,In_616,In_1609);
xnor U983 (N_983,N_260,In_2523);
nand U984 (N_984,In_524,In_445);
or U985 (N_985,In_1569,In_2137);
and U986 (N_986,In_2619,In_471);
and U987 (N_987,In_2048,In_381);
nand U988 (N_988,In_1702,In_177);
nand U989 (N_989,N_224,In_1172);
or U990 (N_990,In_1114,In_2615);
nand U991 (N_991,In_1544,N_236);
nand U992 (N_992,In_810,In_2712);
xor U993 (N_993,In_1084,In_16);
or U994 (N_994,In_1092,In_2214);
and U995 (N_995,N_184,N_65);
nor U996 (N_996,In_210,In_86);
nand U997 (N_997,In_2175,In_57);
xor U998 (N_998,In_5,In_2514);
xnor U999 (N_999,In_2774,In_2708);
or U1000 (N_1000,N_220,N_353);
nand U1001 (N_1001,In_896,In_115);
nand U1002 (N_1002,In_2316,N_561);
and U1003 (N_1003,In_717,N_528);
nor U1004 (N_1004,N_137,In_2470);
xor U1005 (N_1005,In_521,In_2922);
nand U1006 (N_1006,In_18,N_820);
nand U1007 (N_1007,In_170,In_1627);
or U1008 (N_1008,N_531,In_2481);
and U1009 (N_1009,In_868,N_560);
nand U1010 (N_1010,In_2441,In_2786);
or U1011 (N_1011,In_789,N_400);
xnor U1012 (N_1012,N_772,In_182);
nand U1013 (N_1013,In_779,In_2455);
nand U1014 (N_1014,N_913,In_1382);
and U1015 (N_1015,In_2859,N_214);
and U1016 (N_1016,N_399,N_330);
xnor U1017 (N_1017,N_963,In_1905);
xnor U1018 (N_1018,In_2063,N_618);
or U1019 (N_1019,N_108,N_15);
and U1020 (N_1020,N_925,N_455);
nor U1021 (N_1021,N_496,N_38);
nor U1022 (N_1022,N_435,N_114);
nor U1023 (N_1023,In_416,In_1236);
or U1024 (N_1024,In_1597,In_1845);
nor U1025 (N_1025,N_866,N_774);
and U1026 (N_1026,N_799,N_705);
nor U1027 (N_1027,N_566,N_835);
and U1028 (N_1028,In_578,In_2803);
and U1029 (N_1029,N_921,In_2677);
nand U1030 (N_1030,In_2833,N_96);
and U1031 (N_1031,N_667,N_991);
and U1032 (N_1032,N_971,In_989);
or U1033 (N_1033,In_752,In_386);
or U1034 (N_1034,In_2917,In_2578);
and U1035 (N_1035,In_2919,In_114);
nor U1036 (N_1036,In_2040,In_1258);
and U1037 (N_1037,In_1408,In_441);
nand U1038 (N_1038,In_1797,In_1496);
nor U1039 (N_1039,N_501,N_199);
nand U1040 (N_1040,In_2682,N_599);
xnor U1041 (N_1041,In_454,In_1824);
or U1042 (N_1042,N_909,N_784);
or U1043 (N_1043,N_967,In_72);
and U1044 (N_1044,In_1679,In_1417);
xor U1045 (N_1045,In_2783,N_781);
nor U1046 (N_1046,In_862,In_1652);
nand U1047 (N_1047,In_2384,In_1812);
or U1048 (N_1048,In_1430,N_535);
or U1049 (N_1049,In_1131,In_1893);
xor U1050 (N_1050,N_99,In_1598);
or U1051 (N_1051,In_2849,In_1923);
or U1052 (N_1052,In_2378,N_738);
nor U1053 (N_1053,In_4,N_194);
xor U1054 (N_1054,N_707,In_2478);
or U1055 (N_1055,In_767,In_2637);
nand U1056 (N_1056,N_195,N_818);
xor U1057 (N_1057,N_150,N_502);
xnor U1058 (N_1058,N_750,N_813);
or U1059 (N_1059,N_454,In_2802);
or U1060 (N_1060,N_810,N_120);
xnor U1061 (N_1061,In_2566,N_302);
nand U1062 (N_1062,In_1180,In_2625);
nand U1063 (N_1063,N_838,In_2881);
nor U1064 (N_1064,In_1885,N_609);
nor U1065 (N_1065,In_2022,N_637);
nor U1066 (N_1066,In_2801,In_2412);
nor U1067 (N_1067,N_582,N_924);
nor U1068 (N_1068,In_243,N_590);
and U1069 (N_1069,N_301,In_1916);
xnor U1070 (N_1070,N_596,In_2674);
nand U1071 (N_1071,In_599,In_680);
nand U1072 (N_1072,In_1308,In_1725);
or U1073 (N_1073,In_1671,N_238);
and U1074 (N_1074,In_1176,N_125);
nor U1075 (N_1075,N_733,In_2973);
or U1076 (N_1076,N_581,In_2639);
nor U1077 (N_1077,In_22,N_629);
or U1078 (N_1078,In_657,In_1554);
nor U1079 (N_1079,In_2357,N_676);
xor U1080 (N_1080,In_2601,In_1360);
and U1081 (N_1081,In_247,In_582);
xnor U1082 (N_1082,N_333,In_2912);
nor U1083 (N_1083,In_446,In_832);
or U1084 (N_1084,In_916,In_2818);
nand U1085 (N_1085,In_2767,In_1178);
or U1086 (N_1086,In_1708,N_863);
nor U1087 (N_1087,In_2676,In_407);
nor U1088 (N_1088,In_720,In_865);
nor U1089 (N_1089,In_98,N_170);
or U1090 (N_1090,In_2984,N_990);
xor U1091 (N_1091,N_465,In_2409);
or U1092 (N_1092,N_169,N_251);
nand U1093 (N_1093,In_1729,N_593);
and U1094 (N_1094,N_981,N_639);
or U1095 (N_1095,In_686,In_2206);
nor U1096 (N_1096,In_2873,N_737);
or U1097 (N_1097,N_335,N_160);
nand U1098 (N_1098,In_100,N_77);
nand U1099 (N_1099,In_1090,In_1299);
nor U1100 (N_1100,In_380,N_624);
xor U1101 (N_1101,N_710,In_434);
and U1102 (N_1102,N_202,N_604);
or U1103 (N_1103,N_811,In_1976);
nand U1104 (N_1104,N_80,In_1416);
nand U1105 (N_1105,In_11,In_1388);
and U1106 (N_1106,In_2446,In_699);
nand U1107 (N_1107,In_2725,N_627);
nor U1108 (N_1108,In_1147,In_1260);
or U1109 (N_1109,N_975,In_345);
nand U1110 (N_1110,In_925,N_569);
or U1111 (N_1111,In_1956,In_1330);
nand U1112 (N_1112,N_427,In_770);
nand U1113 (N_1113,In_1549,N_876);
or U1114 (N_1114,N_577,In_1653);
nand U1115 (N_1115,In_698,N_165);
nor U1116 (N_1116,In_2618,In_1319);
xor U1117 (N_1117,N_958,N_882);
nand U1118 (N_1118,In_1847,N_213);
nor U1119 (N_1119,In_1282,N_429);
and U1120 (N_1120,In_2763,N_446);
and U1121 (N_1121,In_1317,N_230);
and U1122 (N_1122,In_2752,In_894);
xnor U1123 (N_1123,In_183,In_709);
nand U1124 (N_1124,N_486,In_2362);
or U1125 (N_1125,In_2456,In_2932);
nor U1126 (N_1126,In_967,In_1877);
or U1127 (N_1127,N_289,In_734);
nor U1128 (N_1128,N_908,N_906);
nand U1129 (N_1129,In_15,N_576);
nor U1130 (N_1130,In_645,In_970);
or U1131 (N_1131,In_204,N_78);
and U1132 (N_1132,In_2459,In_622);
or U1133 (N_1133,In_2422,In_302);
nor U1134 (N_1134,N_544,In_710);
nand U1135 (N_1135,In_1567,In_1879);
or U1136 (N_1136,N_511,N_960);
and U1137 (N_1137,In_1086,In_1560);
nand U1138 (N_1138,N_359,In_1383);
xnor U1139 (N_1139,In_1030,In_1625);
nand U1140 (N_1140,In_1871,N_416);
and U1141 (N_1141,In_1396,In_1391);
or U1142 (N_1142,N_212,N_555);
and U1143 (N_1143,In_2838,N_97);
nor U1144 (N_1144,In_75,N_25);
nand U1145 (N_1145,In_1909,In_1423);
nor U1146 (N_1146,In_1658,N_665);
and U1147 (N_1147,N_611,N_586);
nor U1148 (N_1148,In_567,N_443);
nor U1149 (N_1149,In_1098,In_2406);
nor U1150 (N_1150,N_509,In_2359);
or U1151 (N_1151,N_942,In_2385);
and U1152 (N_1152,N_436,In_1292);
or U1153 (N_1153,N_780,N_573);
or U1154 (N_1154,In_1410,In_1044);
xor U1155 (N_1155,N_2,N_918);
and U1156 (N_1156,N_638,In_393);
xnor U1157 (N_1157,N_533,N_433);
xor U1158 (N_1158,N_10,In_2829);
and U1159 (N_1159,In_2308,N_140);
nand U1160 (N_1160,N_355,N_206);
nand U1161 (N_1161,In_286,In_1826);
nor U1162 (N_1162,In_1352,In_1677);
or U1163 (N_1163,N_659,N_246);
nand U1164 (N_1164,N_616,N_768);
and U1165 (N_1165,N_221,In_1325);
nand U1166 (N_1166,In_1586,In_2701);
xnor U1167 (N_1167,In_2894,In_2543);
nand U1168 (N_1168,In_1433,In_1399);
xnor U1169 (N_1169,In_1526,N_388);
nand U1170 (N_1170,N_222,In_1585);
or U1171 (N_1171,In_922,In_253);
and U1172 (N_1172,N_143,In_2976);
nor U1173 (N_1173,N_136,In_469);
xnor U1174 (N_1174,In_1045,N_634);
nand U1175 (N_1175,N_41,In_2740);
and U1176 (N_1176,In_2851,In_2684);
or U1177 (N_1177,In_639,In_748);
nor U1178 (N_1178,In_2427,In_1494);
nand U1179 (N_1179,N_371,In_1432);
or U1180 (N_1180,In_2195,In_436);
nor U1181 (N_1181,N_636,In_2100);
xnor U1182 (N_1182,N_758,N_766);
xor U1183 (N_1183,In_517,N_730);
or U1184 (N_1184,In_405,In_892);
or U1185 (N_1185,In_867,N_932);
or U1186 (N_1186,In_511,In_1411);
nand U1187 (N_1187,N_403,N_152);
and U1188 (N_1188,N_600,In_1302);
and U1189 (N_1189,In_1867,N_514);
nor U1190 (N_1190,N_729,N_723);
nor U1191 (N_1191,N_826,N_547);
xor U1192 (N_1192,In_2840,N_491);
nor U1193 (N_1193,In_670,N_988);
xor U1194 (N_1194,N_701,In_930);
and U1195 (N_1195,In_2889,In_269);
nor U1196 (N_1196,N_928,In_1273);
xor U1197 (N_1197,In_1029,In_2319);
or U1198 (N_1198,In_817,In_1540);
and U1199 (N_1199,In_2794,N_324);
nor U1200 (N_1200,In_2123,In_722);
or U1201 (N_1201,N_147,In_1324);
or U1202 (N_1202,N_837,N_93);
nor U1203 (N_1203,In_2915,N_716);
nor U1204 (N_1204,In_1021,In_2502);
xnor U1205 (N_1205,N_621,In_1686);
nand U1206 (N_1206,In_1604,In_668);
nor U1207 (N_1207,In_835,In_666);
and U1208 (N_1208,N_727,In_1458);
or U1209 (N_1209,N_831,In_2962);
nand U1210 (N_1210,In_512,N_420);
nand U1211 (N_1211,N_494,In_2836);
or U1212 (N_1212,In_2950,N_901);
nor U1213 (N_1213,N_538,In_2170);
nor U1214 (N_1214,In_2320,In_754);
nand U1215 (N_1215,In_676,In_576);
and U1216 (N_1216,N_669,In_1595);
nand U1217 (N_1217,In_1035,N_308);
and U1218 (N_1218,In_1081,In_2021);
and U1219 (N_1219,In_914,In_803);
xor U1220 (N_1220,In_2420,N_379);
nand U1221 (N_1221,In_1434,In_1079);
and U1222 (N_1222,In_2104,N_13);
and U1223 (N_1223,N_118,In_46);
nand U1224 (N_1224,In_337,In_2929);
nand U1225 (N_1225,In_2423,In_2255);
nand U1226 (N_1226,In_1241,N_677);
xnor U1227 (N_1227,In_2858,N_944);
nor U1228 (N_1228,In_690,N_759);
and U1229 (N_1229,In_1211,N_864);
xor U1230 (N_1230,In_632,N_304);
and U1231 (N_1231,N_885,In_281);
nor U1232 (N_1232,N_868,N_972);
xor U1233 (N_1233,In_2964,In_2773);
or U1234 (N_1234,In_747,In_2812);
and U1235 (N_1235,In_515,N_207);
or U1236 (N_1236,N_419,In_1285);
nand U1237 (N_1237,In_2439,In_2471);
nand U1238 (N_1238,N_288,In_1116);
nor U1239 (N_1239,N_658,In_2695);
xor U1240 (N_1240,In_1110,In_264);
or U1241 (N_1241,In_1006,N_113);
nand U1242 (N_1242,N_85,N_515);
xnor U1243 (N_1243,In_2811,N_879);
xnor U1244 (N_1244,In_2059,In_2900);
nor U1245 (N_1245,N_89,In_14);
nand U1246 (N_1246,In_1739,N_532);
and U1247 (N_1247,In_2089,N_941);
nor U1248 (N_1248,N_232,In_1880);
xor U1249 (N_1249,In_1165,N_205);
or U1250 (N_1250,N_765,In_338);
xnor U1251 (N_1251,N_675,In_482);
and U1252 (N_1252,In_285,In_1338);
nor U1253 (N_1253,In_148,N_857);
nand U1254 (N_1254,In_635,In_1068);
nor U1255 (N_1255,In_239,In_2383);
xnor U1256 (N_1256,N_601,In_2322);
nor U1257 (N_1257,N_934,In_1047);
xor U1258 (N_1258,In_400,N_622);
and U1259 (N_1259,In_2473,In_1873);
xor U1260 (N_1260,In_2796,In_962);
nor U1261 (N_1261,N_910,In_106);
nor U1262 (N_1262,N_162,N_623);
nand U1263 (N_1263,N_469,N_828);
nand U1264 (N_1264,In_1207,In_440);
and U1265 (N_1265,In_628,N_853);
nand U1266 (N_1266,N_459,N_619);
or U1267 (N_1267,In_2914,In_2447);
xnor U1268 (N_1268,N_394,In_82);
xor U1269 (N_1269,N_683,N_880);
and U1270 (N_1270,In_2230,In_2814);
and U1271 (N_1271,N_898,In_549);
xnor U1272 (N_1272,In_1169,In_1935);
xor U1273 (N_1273,N_323,N_32);
and U1274 (N_1274,In_449,In_174);
xor U1275 (N_1275,N_776,In_2281);
nand U1276 (N_1276,In_965,In_41);
or U1277 (N_1277,N_751,In_1804);
nand U1278 (N_1278,N_954,N_396);
and U1279 (N_1279,N_178,In_124);
or U1280 (N_1280,N_689,In_2026);
and U1281 (N_1281,In_1163,In_2457);
nand U1282 (N_1282,In_2550,N_787);
or U1283 (N_1283,In_1051,N_617);
nand U1284 (N_1284,N_945,In_1303);
nand U1285 (N_1285,In_1316,In_1939);
xor U1286 (N_1286,N_151,In_1669);
nand U1287 (N_1287,In_2057,N_536);
nor U1288 (N_1288,N_712,In_530);
and U1289 (N_1289,In_1275,N_233);
nor U1290 (N_1290,In_2562,N_186);
or U1291 (N_1291,N_565,N_402);
or U1292 (N_1292,In_908,In_1283);
and U1293 (N_1293,N_12,N_55);
or U1294 (N_1294,In_277,N_67);
and U1295 (N_1295,N_139,N_694);
nor U1296 (N_1296,N_891,N_578);
xnor U1297 (N_1297,In_1589,In_2111);
nand U1298 (N_1298,In_317,In_1234);
and U1299 (N_1299,In_2112,In_1206);
xor U1300 (N_1300,In_820,N_728);
xor U1301 (N_1301,In_1862,In_374);
nor U1302 (N_1302,In_2793,In_2416);
xnor U1303 (N_1303,N_931,In_2579);
or U1304 (N_1304,In_276,N_628);
xnor U1305 (N_1305,N_649,In_2687);
nand U1306 (N_1306,N_947,In_1485);
xor U1307 (N_1307,In_2610,In_107);
xnor U1308 (N_1308,In_641,N_375);
or U1309 (N_1309,In_262,N_340);
or U1310 (N_1310,In_2030,In_1850);
xor U1311 (N_1311,In_193,In_2043);
and U1312 (N_1312,N_193,In_732);
or U1313 (N_1313,N_718,N_671);
or U1314 (N_1314,In_2254,In_2318);
or U1315 (N_1315,N_985,In_694);
nand U1316 (N_1316,In_2215,In_2564);
or U1317 (N_1317,In_1864,N_969);
xor U1318 (N_1318,In_2995,In_2587);
nand U1319 (N_1319,N_468,In_259);
xnor U1320 (N_1320,N_339,In_1358);
nand U1321 (N_1321,N_129,In_2337);
nand U1322 (N_1322,In_996,In_1792);
xnor U1323 (N_1323,In_1343,N_786);
and U1324 (N_1324,In_2612,In_1740);
nor U1325 (N_1325,N_473,In_502);
xnor U1326 (N_1326,In_2151,In_1462);
xnor U1327 (N_1327,In_2480,In_2734);
nand U1328 (N_1328,In_1519,In_1264);
xor U1329 (N_1329,N_73,N_953);
nor U1330 (N_1330,In_2517,In_1843);
and U1331 (N_1331,In_1941,In_2118);
nand U1332 (N_1332,N_777,In_1087);
and U1333 (N_1333,In_365,In_2518);
nand U1334 (N_1334,N_49,In_1984);
and U1335 (N_1335,N_959,In_2072);
xor U1336 (N_1336,N_653,N_505);
nor U1337 (N_1337,In_1966,In_550);
xor U1338 (N_1338,In_96,In_2278);
and U1339 (N_1339,In_2286,N_900);
nor U1340 (N_1340,In_528,N_497);
xnor U1341 (N_1341,In_34,In_2164);
and U1342 (N_1342,In_1760,N_652);
or U1343 (N_1343,N_521,N_741);
nor U1344 (N_1344,In_791,In_603);
xnor U1345 (N_1345,In_1483,In_2177);
xor U1346 (N_1346,N_401,N_185);
xor U1347 (N_1347,N_644,N_209);
nor U1348 (N_1348,N_480,In_326);
and U1349 (N_1349,In_2974,In_775);
and U1350 (N_1350,In_2739,N_979);
and U1351 (N_1351,N_153,N_250);
nor U1352 (N_1352,In_322,N_978);
or U1353 (N_1353,N_847,In_1932);
xor U1354 (N_1354,N_588,N_935);
nand U1355 (N_1355,In_851,In_876);
nor U1356 (N_1356,In_223,N_717);
nor U1357 (N_1357,N_841,N_479);
or U1358 (N_1358,N_647,In_716);
xor U1359 (N_1359,In_2291,In_146);
nand U1360 (N_1360,N_116,N_731);
or U1361 (N_1361,N_749,N_279);
and U1362 (N_1362,N_380,In_924);
nor U1363 (N_1363,N_862,N_444);
or U1364 (N_1364,In_357,In_1418);
nor U1365 (N_1365,In_1453,N_607);
xor U1366 (N_1366,N_518,In_1191);
or U1367 (N_1367,In_1333,N_848);
or U1368 (N_1368,In_1696,In_2996);
nor U1369 (N_1369,N_439,N_740);
or U1370 (N_1370,In_201,N_903);
xnor U1371 (N_1371,N_61,N_626);
nor U1372 (N_1372,In_2886,In_252);
nand U1373 (N_1373,N_154,In_2165);
and U1374 (N_1374,N_663,N_949);
nand U1375 (N_1375,In_1409,N_377);
nor U1376 (N_1376,N_761,N_499);
and U1377 (N_1377,N_610,N_161);
nor U1378 (N_1378,In_737,N_922);
nand U1379 (N_1379,N_673,N_656);
or U1380 (N_1380,N_306,In_347);
nand U1381 (N_1381,N_691,In_2686);
xnor U1382 (N_1382,In_2160,N_977);
or U1383 (N_1383,N_702,N_782);
and U1384 (N_1384,N_997,In_1024);
or U1385 (N_1385,N_575,In_217);
nand U1386 (N_1386,N_374,In_220);
nor U1387 (N_1387,N_827,In_2327);
xor U1388 (N_1388,N_754,In_1584);
or U1389 (N_1389,In_1528,N_519);
xnor U1390 (N_1390,In_507,N_452);
xor U1391 (N_1391,N_332,N_354);
or U1392 (N_1392,In_2003,N_121);
and U1393 (N_1393,In_2036,N_48);
xor U1394 (N_1394,N_361,N_393);
nor U1395 (N_1395,N_441,In_1927);
nand U1396 (N_1396,In_873,N_64);
xor U1397 (N_1397,N_955,In_1778);
nor U1398 (N_1398,In_1551,N_82);
and U1399 (N_1399,In_2989,N_996);
and U1400 (N_1400,In_267,N_859);
and U1401 (N_1401,N_836,In_1749);
and U1402 (N_1402,In_2011,In_1736);
nand U1403 (N_1403,N_736,In_1321);
and U1404 (N_1404,In_2660,In_1911);
and U1405 (N_1405,In_1015,In_2009);
nand U1406 (N_1406,In_2130,In_1612);
or U1407 (N_1407,In_1094,In_2693);
nand U1408 (N_1408,N_367,N_989);
and U1409 (N_1409,N_574,N_456);
nor U1410 (N_1410,N_646,N_526);
nor U1411 (N_1411,In_1963,N_783);
and U1412 (N_1412,N_101,In_919);
nand U1413 (N_1413,In_819,In_2199);
or U1414 (N_1414,In_1856,In_40);
xor U1415 (N_1415,In_42,In_519);
and U1416 (N_1416,N_34,In_1380);
nor U1417 (N_1417,N_487,In_2972);
xnor U1418 (N_1418,In_2500,In_2277);
nor U1419 (N_1419,In_627,In_2782);
xor U1420 (N_1420,N_764,In_2772);
nor U1421 (N_1421,N_763,In_2302);
or U1422 (N_1422,In_2435,In_656);
nor U1423 (N_1423,N_587,In_2515);
nand U1424 (N_1424,In_1250,N_968);
nand U1425 (N_1425,In_1429,In_1498);
nand U1426 (N_1426,N_568,In_1297);
nor U1427 (N_1427,N_156,In_966);
and U1428 (N_1428,In_1748,In_3);
or U1429 (N_1429,N_792,In_1734);
xnor U1430 (N_1430,N_123,In_293);
nand U1431 (N_1431,In_508,In_378);
nor U1432 (N_1432,N_318,In_453);
or U1433 (N_1433,N_91,In_2309);
or U1434 (N_1434,In_1855,N_739);
xnor U1435 (N_1435,In_2520,N_541);
xor U1436 (N_1436,N_234,In_612);
xnor U1437 (N_1437,N_584,In_2644);
nand U1438 (N_1438,In_2087,In_1606);
or U1439 (N_1439,In_2093,N_812);
nand U1440 (N_1440,In_516,In_798);
nor U1441 (N_1441,N_894,In_624);
xnor U1442 (N_1442,In_2106,In_1960);
nor U1443 (N_1443,N_883,In_1608);
nor U1444 (N_1444,In_1998,N_734);
nand U1445 (N_1445,In_718,In_2468);
nand U1446 (N_1446,In_1594,In_1707);
or U1447 (N_1447,In_2511,In_1049);
or U1448 (N_1448,In_163,N_557);
xnor U1449 (N_1449,In_1441,N_437);
and U1450 (N_1450,In_837,In_81);
or U1451 (N_1451,N_875,N_788);
nand U1452 (N_1452,In_270,In_2722);
or U1453 (N_1453,In_396,In_2307);
or U1454 (N_1454,N_141,In_1629);
and U1455 (N_1455,N_527,N_594);
xor U1456 (N_1456,N_31,In_1511);
or U1457 (N_1457,N_824,In_1439);
or U1458 (N_1458,N_633,In_995);
xor U1459 (N_1459,In_672,In_1370);
xnor U1460 (N_1460,In_2505,In_2055);
and U1461 (N_1461,In_1074,In_2756);
nand U1462 (N_1462,N_998,In_1389);
nand U1463 (N_1463,In_942,N_974);
or U1464 (N_1464,N_243,N_517);
or U1465 (N_1465,N_105,N_183);
xnor U1466 (N_1466,N_285,In_647);
nand U1467 (N_1467,N_271,In_462);
or U1468 (N_1468,N_595,In_735);
and U1469 (N_1469,In_1395,N_999);
nor U1470 (N_1470,In_2867,In_1947);
nor U1471 (N_1471,In_2524,In_2510);
nand U1472 (N_1472,N_651,N_247);
nand U1473 (N_1473,N_680,In_1766);
nor U1474 (N_1474,In_486,N_679);
nand U1475 (N_1475,N_196,In_1175);
and U1476 (N_1476,In_479,In_1931);
and U1477 (N_1477,In_1832,In_953);
xnor U1478 (N_1478,N_391,N_961);
or U1479 (N_1479,In_250,In_195);
and U1480 (N_1480,In_2697,In_2004);
and U1481 (N_1481,In_573,In_644);
and U1482 (N_1482,In_945,In_1070);
nand U1483 (N_1483,In_664,In_510);
and U1484 (N_1484,N_291,N_321);
nand U1485 (N_1485,In_1261,In_1161);
xnor U1486 (N_1486,In_2096,In_1888);
or U1487 (N_1487,N_640,In_2240);
xor U1488 (N_1488,In_637,In_1384);
or U1489 (N_1489,In_212,In_2635);
nor U1490 (N_1490,N_660,In_1479);
nor U1491 (N_1491,In_1305,In_971);
or U1492 (N_1492,In_2083,In_596);
or U1493 (N_1493,In_473,N_191);
and U1494 (N_1494,N_685,N_951);
nor U1495 (N_1495,In_51,In_782);
nor U1496 (N_1496,In_2451,In_2101);
or U1497 (N_1497,N_926,N_503);
nor U1498 (N_1498,In_762,N_329);
nor U1499 (N_1499,In_1293,In_768);
or U1500 (N_1500,N_1147,N_1472);
and U1501 (N_1501,N_208,N_556);
nand U1502 (N_1502,In_1996,N_1265);
xnor U1503 (N_1503,In_2966,N_579);
nor U1504 (N_1504,In_1616,N_1177);
nand U1505 (N_1505,N_1237,In_2208);
nand U1506 (N_1506,In_2403,N_508);
nor U1507 (N_1507,N_612,N_1126);
nor U1508 (N_1508,In_1772,N_976);
nor U1509 (N_1509,In_401,In_1205);
xnor U1510 (N_1510,In_1643,N_434);
nor U1511 (N_1511,In_1362,In_2911);
nor U1512 (N_1512,N_158,In_1046);
and U1513 (N_1513,N_516,N_829);
xnor U1514 (N_1514,N_52,N_695);
nand U1515 (N_1515,In_2971,In_1763);
and U1516 (N_1516,N_1181,N_1162);
xor U1517 (N_1517,N_1293,In_2044);
nand U1518 (N_1518,In_2257,N_1445);
nor U1519 (N_1519,N_1425,N_589);
nand U1520 (N_1520,In_1601,In_1473);
xnor U1521 (N_1521,In_1918,N_1047);
or U1522 (N_1522,N_1443,N_1042);
or U1523 (N_1523,N_1180,In_32);
nor U1524 (N_1524,In_1973,N_1227);
xnor U1525 (N_1525,In_903,In_1588);
or U1526 (N_1526,In_2807,In_496);
and U1527 (N_1527,N_840,N_1248);
or U1528 (N_1528,N_1383,In_2559);
and U1529 (N_1529,N_1034,N_1277);
nand U1530 (N_1530,N_1362,N_564);
or U1531 (N_1531,N_602,In_692);
and U1532 (N_1532,N_1288,In_818);
or U1533 (N_1533,In_2488,In_143);
and U1534 (N_1534,In_537,N_1153);
and U1535 (N_1535,N_892,In_2874);
nor U1536 (N_1536,In_589,N_543);
nor U1537 (N_1537,In_2775,In_2095);
nand U1538 (N_1538,In_318,N_803);
and U1539 (N_1539,N_530,N_844);
nand U1540 (N_1540,In_574,N_687);
nor U1541 (N_1541,N_28,N_1184);
and U1542 (N_1542,In_948,N_920);
nand U1543 (N_1543,N_613,In_2765);
or U1544 (N_1544,N_1079,N_911);
or U1545 (N_1545,In_1750,N_40);
and U1546 (N_1546,In_564,In_1599);
nor U1547 (N_1547,N_1003,N_1093);
and U1548 (N_1548,N_315,N_1489);
nor U1549 (N_1549,In_373,N_1040);
or U1550 (N_1550,N_1161,In_1765);
or U1551 (N_1551,N_890,N_1340);
and U1552 (N_1552,N_666,In_785);
or U1553 (N_1553,In_431,N_320);
nor U1554 (N_1554,N_1230,In_236);
nor U1555 (N_1555,N_352,In_1566);
and U1556 (N_1556,In_2885,In_1684);
xor U1557 (N_1557,N_550,In_2895);
and U1558 (N_1558,N_1212,In_661);
nand U1559 (N_1559,In_786,In_1713);
nor U1560 (N_1560,N_1104,N_983);
nand U1561 (N_1561,In_1018,In_2525);
and U1562 (N_1562,In_444,N_1440);
and U1563 (N_1563,In_2110,In_2985);
nand U1564 (N_1564,N_591,N_775);
xor U1565 (N_1565,In_2489,In_2616);
or U1566 (N_1566,N_940,N_1236);
nand U1567 (N_1567,N_808,In_2355);
xnor U1568 (N_1568,N_867,N_1057);
xnor U1569 (N_1569,In_674,In_1229);
and U1570 (N_1570,N_1054,N_962);
nand U1571 (N_1571,N_188,N_1364);
nand U1572 (N_1572,N_1239,N_1175);
nand U1573 (N_1573,In_7,N_1399);
or U1574 (N_1574,N_1150,In_1242);
or U1575 (N_1575,N_1048,N_1339);
xnor U1576 (N_1576,In_2672,In_1421);
nand U1577 (N_1577,N_678,In_706);
nor U1578 (N_1578,N_245,N_858);
or U1579 (N_1579,N_927,In_725);
nor U1580 (N_1580,In_2757,N_1455);
xnor U1581 (N_1581,N_30,N_322);
or U1582 (N_1582,N_1458,N_725);
nand U1583 (N_1583,N_1426,In_121);
xnor U1584 (N_1584,N_773,N_1229);
nand U1585 (N_1585,In_1450,N_1046);
and U1586 (N_1586,In_266,In_1721);
xor U1587 (N_1587,N_1470,In_1508);
xor U1588 (N_1588,N_1255,In_1182);
nand U1589 (N_1589,N_1019,In_388);
or U1590 (N_1590,In_1216,N_1446);
nand U1591 (N_1591,N_1356,In_946);
nor U1592 (N_1592,N_1380,N_697);
or U1593 (N_1593,N_917,N_292);
nor U1594 (N_1594,In_346,N_1493);
nand U1595 (N_1595,N_1419,N_1030);
and U1596 (N_1596,In_73,In_1228);
nand U1597 (N_1597,N_1320,In_1361);
nor U1598 (N_1598,N_1039,N_1244);
xnor U1599 (N_1599,In_978,N_1405);
and U1600 (N_1600,In_2727,In_1149);
xnor U1601 (N_1601,N_1077,N_878);
nand U1602 (N_1602,In_2599,In_838);
xnor U1603 (N_1603,In_943,N_1306);
xor U1604 (N_1604,N_1376,N_1112);
or U1605 (N_1605,In_1937,In_1579);
nor U1606 (N_1606,N_1084,In_2992);
nand U1607 (N_1607,In_878,N_1453);
nand U1608 (N_1608,In_1155,N_1452);
and U1609 (N_1609,N_1171,N_1251);
nor U1610 (N_1610,In_92,N_654);
nand U1611 (N_1611,N_950,N_802);
nand U1612 (N_1612,N_744,N_1469);
nand U1613 (N_1613,N_625,N_239);
nand U1614 (N_1614,In_2711,N_392);
or U1615 (N_1615,In_123,N_1270);
or U1616 (N_1616,N_282,N_1250);
xor U1617 (N_1617,N_537,N_0);
nor U1618 (N_1618,N_1013,In_1488);
and U1619 (N_1619,In_1559,In_2483);
nor U1620 (N_1620,In_1322,N_1000);
nand U1621 (N_1621,N_1083,N_1318);
xnor U1622 (N_1622,N_1163,In_136);
xor U1623 (N_1623,In_1471,N_1033);
and U1624 (N_1624,N_1022,N_1105);
and U1625 (N_1625,N_1232,N_1103);
and U1626 (N_1626,In_1125,In_2351);
nand U1627 (N_1627,In_355,N_1085);
or U1628 (N_1628,In_2495,N_1374);
nand U1629 (N_1629,N_1410,In_417);
nor U1630 (N_1630,In_1444,N_1167);
nor U1631 (N_1631,N_559,N_1422);
nor U1632 (N_1632,N_726,In_1232);
and U1633 (N_1633,In_2614,In_927);
nor U1634 (N_1634,N_417,In_2944);
nor U1635 (N_1635,In_2931,N_1435);
and U1636 (N_1636,In_1048,N_1411);
nor U1637 (N_1637,In_2479,N_946);
xnor U1638 (N_1638,N_1494,In_1764);
nor U1639 (N_1639,In_2252,In_2899);
and U1640 (N_1640,N_1051,In_649);
nor U1641 (N_1641,In_94,In_1556);
nand U1642 (N_1642,N_284,In_1720);
and U1643 (N_1643,N_757,In_2791);
nor U1644 (N_1644,N_800,N_684);
nand U1645 (N_1645,In_2437,In_1289);
nand U1646 (N_1646,N_1131,N_111);
and U1647 (N_1647,N_470,N_1151);
or U1648 (N_1648,N_382,N_1207);
or U1649 (N_1649,N_1368,In_1487);
nand U1650 (N_1650,In_2656,N_1461);
nor U1651 (N_1651,N_798,In_1381);
xnor U1652 (N_1652,N_1071,In_2540);
nand U1653 (N_1653,In_1983,N_907);
or U1654 (N_1654,In_617,N_1297);
or U1655 (N_1655,In_1267,In_2476);
xnor U1656 (N_1656,N_938,N_368);
nor U1657 (N_1657,In_2347,N_668);
xor U1658 (N_1658,In_227,N_1415);
nor U1659 (N_1659,N_1140,N_510);
nand U1660 (N_1660,N_957,N_916);
and U1661 (N_1661,In_63,N_1447);
and U1662 (N_1662,N_994,N_187);
xor U1663 (N_1663,In_1390,N_688);
xnor U1664 (N_1664,N_1343,N_395);
nand U1665 (N_1665,N_79,In_62);
xor U1666 (N_1666,N_1402,N_698);
xnor U1667 (N_1667,N_513,N_756);
and U1668 (N_1668,N_424,In_630);
xnor U1669 (N_1669,In_504,In_2534);
and U1670 (N_1670,N_1197,In_331);
xnor U1671 (N_1671,In_1017,N_1498);
nor U1672 (N_1672,In_1811,N_814);
xnor U1673 (N_1673,N_643,N_1097);
nor U1674 (N_1674,N_1393,N_1017);
or U1675 (N_1675,In_2424,In_1220);
nand U1676 (N_1676,N_670,In_2102);
nor U1677 (N_1677,N_839,N_1436);
or U1678 (N_1678,N_300,N_63);
and U1679 (N_1679,N_1286,N_1122);
xnor U1680 (N_1680,N_992,In_2736);
nor U1681 (N_1681,In_2128,N_1347);
xnor U1682 (N_1682,N_631,N_732);
xor U1683 (N_1683,N_423,N_1348);
nand U1684 (N_1684,In_2986,N_793);
xnor U1685 (N_1685,In_2608,N_17);
nand U1686 (N_1686,N_1378,In_2626);
nor U1687 (N_1687,In_2924,In_1858);
nand U1688 (N_1688,N_1325,N_1354);
or U1689 (N_1689,N_1216,In_2150);
nand U1690 (N_1690,N_1262,N_1090);
or U1691 (N_1691,In_2352,N_1370);
xor U1692 (N_1692,N_1166,In_88);
or U1693 (N_1693,In_557,N_1401);
nand U1694 (N_1694,In_256,N_1110);
nand U1695 (N_1695,N_50,N_1224);
and U1696 (N_1696,N_856,In_450);
or U1697 (N_1697,In_1773,N_1333);
nor U1698 (N_1698,N_606,N_1396);
nor U1699 (N_1699,In_394,In_140);
nor U1700 (N_1700,N_797,N_1063);
nor U1701 (N_1701,N_264,N_1011);
nor U1702 (N_1702,In_2227,In_730);
and U1703 (N_1703,N_1468,N_937);
or U1704 (N_1704,N_1064,In_2168);
nand U1705 (N_1705,N_1497,In_2887);
or U1706 (N_1706,N_1138,N_159);
xor U1707 (N_1707,N_442,N_1408);
nand U1708 (N_1708,N_1478,In_231);
xnor U1709 (N_1709,In_1193,N_1012);
and U1710 (N_1710,N_1178,In_1455);
or U1711 (N_1711,N_1466,N_451);
nor U1712 (N_1712,In_1898,N_1205);
nand U1713 (N_1713,N_1298,N_872);
or U1714 (N_1714,In_2090,In_1306);
and U1715 (N_1715,N_785,N_1431);
nor U1716 (N_1716,N_1384,N_603);
and U1717 (N_1717,N_1360,N_1441);
nor U1718 (N_1718,N_893,In_452);
nand U1719 (N_1719,N_109,N_1099);
xnor U1720 (N_1720,N_1133,N_752);
nand U1721 (N_1721,N_484,N_1055);
nand U1722 (N_1722,In_1698,In_1870);
nand U1723 (N_1723,N_1186,N_1459);
and U1724 (N_1724,N_888,In_2921);
and U1725 (N_1725,N_795,In_2187);
xor U1726 (N_1726,In_2664,N_1349);
or U1727 (N_1727,N_148,N_1208);
xor U1728 (N_1728,N_552,N_1142);
or U1729 (N_1729,N_806,N_1463);
xnor U1730 (N_1730,N_1164,N_686);
and U1731 (N_1731,N_970,N_743);
nor U1732 (N_1732,N_173,N_1119);
xnor U1733 (N_1733,N_500,N_58);
nor U1734 (N_1734,N_1066,In_1112);
nand U1735 (N_1735,N_94,In_1985);
nand U1736 (N_1736,In_2119,N_520);
nor U1737 (N_1737,N_762,N_327);
or U1738 (N_1738,N_1242,In_1069);
nand U1739 (N_1739,N_1183,In_2848);
nand U1740 (N_1740,N_572,N_1423);
and U1741 (N_1741,N_558,N_1369);
nor U1742 (N_1742,In_2638,N_362);
or U1743 (N_1743,N_266,In_375);
nor U1744 (N_1744,N_522,In_2449);
and U1745 (N_1745,In_1682,N_929);
nand U1746 (N_1746,N_477,N_312);
and U1747 (N_1747,N_1263,N_1091);
nor U1748 (N_1748,N_172,In_864);
xor U1749 (N_1749,N_1149,In_429);
nor U1750 (N_1750,N_348,N_1135);
xnor U1751 (N_1751,N_540,N_529);
nand U1752 (N_1752,In_1089,N_973);
and U1753 (N_1753,N_1471,N_119);
or U1754 (N_1754,In_97,N_711);
nand U1755 (N_1755,In_2356,In_192);
or U1756 (N_1756,N_1141,In_399);
or U1757 (N_1757,In_2189,N_506);
or U1758 (N_1758,N_1217,N_1258);
nand U1759 (N_1759,N_912,N_1337);
xor U1760 (N_1760,N_1015,N_1328);
or U1761 (N_1761,N_746,N_1361);
nand U1762 (N_1762,In_2023,N_1056);
xor U1763 (N_1763,N_1278,In_1803);
nor U1764 (N_1764,N_1082,N_632);
nand U1765 (N_1765,In_2183,N_1154);
or U1766 (N_1766,N_296,In_758);
nor U1767 (N_1767,In_2665,N_1428);
nor U1768 (N_1768,N_1173,In_1221);
or U1769 (N_1769,N_357,N_1228);
and U1770 (N_1770,In_655,N_735);
xnor U1771 (N_1771,N_846,In_2759);
xor U1772 (N_1772,N_1386,In_1040);
nor U1773 (N_1773,N_767,N_865);
nand U1774 (N_1774,In_1345,In_2226);
nand U1775 (N_1775,N_608,N_842);
or U1776 (N_1776,In_2690,In_751);
or U1777 (N_1777,In_2463,N_1139);
xnor U1778 (N_1778,N_1395,In_879);
or U1779 (N_1779,In_1456,N_770);
xor U1780 (N_1780,N_1213,In_604);
and U1781 (N_1781,N_240,N_645);
and U1782 (N_1782,N_337,N_1220);
and U1783 (N_1783,In_1538,N_1062);
or U1784 (N_1784,N_1276,N_850);
nand U1785 (N_1785,N_693,N_1366);
or U1786 (N_1786,N_1148,N_1215);
xnor U1787 (N_1787,In_44,In_2205);
xnor U1788 (N_1788,In_478,In_2401);
xnor U1789 (N_1789,N_1245,In_2879);
xor U1790 (N_1790,N_1221,N_1407);
and U1791 (N_1791,N_1316,N_1027);
xnor U1792 (N_1792,N_1132,N_498);
xnor U1793 (N_1793,N_1130,In_813);
and U1794 (N_1794,N_1107,In_2834);
nand U1795 (N_1795,In_348,In_546);
or U1796 (N_1796,N_980,In_1693);
nand U1797 (N_1797,In_467,In_1863);
nor U1798 (N_1798,N_1449,N_1143);
nor U1799 (N_1799,N_274,N_1253);
or U1800 (N_1800,N_771,N_852);
or U1801 (N_1801,N_1491,N_42);
xor U1802 (N_1802,In_2629,In_387);
nor U1803 (N_1803,In_481,In_2142);
and U1804 (N_1804,N_630,N_1073);
nand U1805 (N_1805,In_525,In_2602);
or U1806 (N_1806,N_553,N_933);
nand U1807 (N_1807,In_2956,N_899);
or U1808 (N_1808,N_1432,In_1307);
nor U1809 (N_1809,In_1930,N_1365);
xor U1810 (N_1810,N_235,N_23);
nor U1811 (N_1811,N_1256,N_1307);
or U1812 (N_1812,N_1353,N_267);
xnor U1813 (N_1813,N_1192,N_923);
nor U1814 (N_1814,In_2557,In_402);
or U1815 (N_1815,N_1234,In_2857);
nand U1816 (N_1816,N_1314,In_673);
nor U1817 (N_1817,N_471,In_288);
xnor U1818 (N_1818,N_1002,N_112);
xor U1819 (N_1819,In_1132,In_484);
and U1820 (N_1820,N_661,N_319);
nand U1821 (N_1821,N_412,In_2497);
and U1822 (N_1822,In_224,N_834);
nand U1823 (N_1823,In_1784,In_1328);
nand U1824 (N_1824,In_1503,N_1061);
xnor U1825 (N_1825,N_261,N_59);
nor U1826 (N_1826,N_1275,N_1392);
or U1827 (N_1827,N_1301,N_713);
and U1828 (N_1828,N_851,N_201);
nor U1829 (N_1829,N_1488,In_1651);
nand U1830 (N_1830,In_958,In_2705);
and U1831 (N_1831,In_2156,In_665);
and U1832 (N_1832,In_161,In_2967);
xnor U1833 (N_1833,In_1520,In_2918);
or U1834 (N_1834,N_1406,N_177);
nor U1835 (N_1835,In_1280,In_569);
and U1836 (N_1836,In_1770,N_1414);
xnor U1837 (N_1837,In_1665,N_1350);
and U1838 (N_1838,In_1988,In_2609);
or U1839 (N_1839,In_1119,In_1027);
xnor U1840 (N_1840,N_823,In_419);
nor U1841 (N_1841,N_832,In_1062);
xnor U1842 (N_1842,N_982,N_1412);
or U1843 (N_1843,N_948,In_858);
nand U1844 (N_1844,N_1261,In_1656);
nand U1845 (N_1845,N_1257,In_1420);
nand U1846 (N_1846,N_1417,N_8);
and U1847 (N_1847,In_1915,N_378);
nand U1848 (N_1848,In_1846,In_1502);
nand U1849 (N_1849,N_1279,N_1483);
nor U1850 (N_1850,N_1233,In_2732);
nand U1851 (N_1851,N_1450,In_2987);
xor U1852 (N_1852,In_55,N_1117);
and U1853 (N_1853,In_2494,In_316);
or U1854 (N_1854,N_1031,N_1357);
or U1855 (N_1855,N_1273,N_597);
nand U1856 (N_1856,In_2844,N_1254);
xor U1857 (N_1857,In_1227,N_1223);
or U1858 (N_1858,N_1326,N_466);
xor U1859 (N_1859,N_16,N_314);
nor U1860 (N_1860,N_325,N_1351);
nand U1861 (N_1861,N_36,In_2167);
and U1862 (N_1862,N_1067,N_1018);
or U1863 (N_1863,N_179,In_105);
xnor U1864 (N_1864,N_567,In_2542);
nor U1865 (N_1865,N_328,In_2317);
or U1866 (N_1866,N_317,In_2823);
nand U1867 (N_1867,In_1921,N_700);
nand U1868 (N_1868,N_1120,N_1168);
nand U1869 (N_1869,N_1076,N_1487);
and U1870 (N_1870,In_1314,In_1195);
xnor U1871 (N_1871,N_1194,N_1050);
and U1872 (N_1872,N_1137,In_1445);
or U1873 (N_1873,In_1167,N_815);
xnor U1874 (N_1874,N_760,In_275);
nand U1875 (N_1875,In_750,N_703);
or U1876 (N_1876,In_826,In_2440);
xor U1877 (N_1877,In_2526,N_1442);
nor U1878 (N_1878,N_1268,N_995);
nor U1879 (N_1879,N_1264,N_1209);
nor U1880 (N_1880,N_1198,N_825);
nand U1881 (N_1881,N_1144,In_1397);
nand U1882 (N_1882,N_592,N_563);
or U1883 (N_1883,N_1269,N_896);
and U1884 (N_1884,N_81,N_200);
or U1885 (N_1885,N_1280,In_2332);
and U1886 (N_1886,N_1125,N_1211);
nand U1887 (N_1887,In_2529,N_1315);
and U1888 (N_1888,N_791,N_881);
nor U1889 (N_1889,In_66,N_1020);
nor U1890 (N_1890,N_1115,N_1465);
nand U1891 (N_1891,In_2544,N_1032);
or U1892 (N_1892,N_1499,N_248);
or U1893 (N_1893,N_664,N_1113);
xor U1894 (N_1894,N_1202,In_2977);
nand U1895 (N_1895,N_905,N_1310);
or U1896 (N_1896,In_2070,In_283);
and U1897 (N_1897,In_1786,N_598);
and U1898 (N_1898,N_919,In_129);
and U1899 (N_1899,In_2528,N_1165);
and U1900 (N_1900,In_369,N_457);
xnor U1901 (N_1901,N_1334,N_1060);
xnor U1902 (N_1902,In_1272,N_1109);
and U1903 (N_1903,N_966,N_92);
or U1904 (N_1904,In_1621,N_1123);
nor U1905 (N_1905,In_1837,In_1727);
xnor U1906 (N_1906,N_1379,N_1102);
nor U1907 (N_1907,N_142,In_112);
and U1908 (N_1908,N_779,In_2603);
nor U1909 (N_1909,N_1203,In_37);
nand U1910 (N_1910,N_1308,N_1475);
nor U1911 (N_1911,In_1835,N_1421);
and U1912 (N_1912,In_2166,N_164);
nand U1913 (N_1913,In_2826,In_2186);
xor U1914 (N_1914,N_874,N_1456);
nor U1915 (N_1915,N_1158,N_692);
or U1916 (N_1916,In_1174,N_747);
xor U1917 (N_1917,N_724,N_778);
xnor U1918 (N_1918,N_103,N_915);
xnor U1919 (N_1919,N_1344,N_662);
xnor U1920 (N_1920,N_548,N_432);
nor U1921 (N_1921,N_405,In_2504);
nand U1922 (N_1922,N_1400,N_1129);
and U1923 (N_1923,In_358,In_2825);
or U1924 (N_1924,N_1059,In_1375);
xor U1925 (N_1925,In_50,N_1010);
or U1926 (N_1926,N_914,N_1413);
and U1927 (N_1927,In_2537,N_1289);
or U1928 (N_1928,In_2669,N_984);
and U1929 (N_1929,N_605,In_395);
or U1930 (N_1930,In_2728,N_1404);
or U1931 (N_1931,N_708,N_720);
xor U1932 (N_1932,N_830,N_493);
or U1933 (N_1933,N_259,In_2305);
or U1934 (N_1934,N_833,In_1631);
and U1935 (N_1935,N_1200,N_95);
nand U1936 (N_1936,In_614,N_1394);
nand U1937 (N_1937,N_1485,In_1290);
xnor U1938 (N_1938,N_690,N_411);
or U1939 (N_1939,N_1045,N_1290);
xnor U1940 (N_1940,In_2474,N_1156);
and U1941 (N_1941,In_2084,In_795);
nor U1942 (N_1942,In_52,In_1151);
and U1943 (N_1943,In_1603,In_442);
nor U1944 (N_1944,N_198,N_1222);
nor U1945 (N_1945,N_1282,In_2548);
or U1946 (N_1946,N_1021,N_1199);
xnor U1947 (N_1947,In_12,In_543);
or U1948 (N_1948,In_2258,N_1305);
nand U1949 (N_1949,N_176,In_1663);
nor U1950 (N_1950,N_1490,In_1980);
nand U1951 (N_1951,In_2709,In_1109);
or U1952 (N_1952,N_542,N_386);
and U1953 (N_1953,N_722,In_1800);
nor U1954 (N_1954,N_794,In_2888);
and U1955 (N_1955,In_697,N_449);
and U1956 (N_1956,N_1486,In_258);
and U1957 (N_1957,N_1409,In_562);
nor U1958 (N_1958,In_2951,In_2906);
and U1959 (N_1959,N_425,N_1058);
and U1960 (N_1960,N_1182,N_1260);
nand U1961 (N_1961,In_2415,N_1330);
and U1962 (N_1962,N_1038,In_607);
or U1963 (N_1963,N_943,N_1159);
nand U1964 (N_1964,N_1434,N_1096);
nand U1965 (N_1965,N_1391,In_2244);
nand U1966 (N_1966,In_1553,N_1302);
and U1967 (N_1967,N_1295,In_2025);
xor U1968 (N_1968,In_58,N_1127);
or U1969 (N_1969,In_2652,N_1424);
nand U1970 (N_1970,N_1080,In_1009);
nor U1971 (N_1971,In_2314,In_764);
nor U1972 (N_1972,In_137,N_1274);
and U1973 (N_1973,In_2930,N_551);
or U1974 (N_1974,N_524,N_904);
nand U1975 (N_1975,N_1252,N_1352);
or U1976 (N_1976,N_993,N_1291);
or U1977 (N_1977,N_1420,In_406);
nand U1978 (N_1978,N_742,In_2846);
or U1979 (N_1979,N_1128,In_2679);
and U1980 (N_1980,In_2998,N_930);
xor U1981 (N_1981,In_1570,N_1398);
nor U1982 (N_1982,N_571,In_2865);
nor U1983 (N_1983,In_1841,N_583);
nor U1984 (N_1984,N_1016,N_753);
nand U1985 (N_1985,N_1179,N_1101);
and U1986 (N_1986,In_2490,N_297);
nor U1987 (N_1987,In_1933,In_2005);
nand U1988 (N_1988,N_1430,In_663);
xnor U1989 (N_1989,N_344,N_182);
xor U1990 (N_1990,N_539,N_1267);
nand U1991 (N_1991,In_2251,In_1468);
and U1992 (N_1992,N_507,N_1319);
and U1993 (N_1993,N_790,N_1124);
nand U1994 (N_1994,N_389,N_902);
and U1995 (N_1995,N_216,N_546);
nand U1996 (N_1996,N_1448,In_468);
and U1997 (N_1997,N_1444,In_2960);
or U1998 (N_1998,In_2731,In_463);
or U1999 (N_1999,N_965,In_651);
or U2000 (N_2000,N_104,N_1737);
nand U2001 (N_2001,N_719,N_1689);
nand U2002 (N_2002,N_1662,N_1671);
or U2003 (N_2003,In_2790,N_1677);
xnor U2004 (N_2004,N_1788,N_1709);
nor U2005 (N_2005,N_1558,N_1739);
nor U2006 (N_2006,N_1890,N_1926);
or U2007 (N_2007,N_1092,In_708);
nand U2008 (N_2008,In_593,N_1533);
and U2009 (N_2009,N_1007,In_594);
and U2010 (N_2010,N_1427,N_845);
xor U2011 (N_2011,In_179,N_219);
and U2012 (N_2012,N_1931,N_1556);
or U2013 (N_2013,In_2173,N_1539);
and U2014 (N_2014,N_1994,N_1563);
and U2015 (N_2015,N_1882,N_1770);
xnor U2016 (N_2016,N_1800,N_1299);
or U2017 (N_2017,N_674,N_755);
nor U2018 (N_2018,N_1336,N_805);
nand U2019 (N_2019,N_1712,N_1616);
xnor U2020 (N_2020,N_1238,N_180);
xor U2021 (N_2021,In_2648,N_1537);
and U2022 (N_2022,N_1756,N_1721);
nand U2023 (N_2023,N_1824,N_1004);
nand U2024 (N_2024,N_1617,In_1962);
or U2025 (N_2025,N_1598,In_893);
nor U2026 (N_2026,In_1097,N_1385);
xor U2027 (N_2027,N_1474,N_1690);
or U2028 (N_2028,N_460,N_410);
xor U2029 (N_2029,N_1716,N_1789);
xnor U2030 (N_2030,N_1805,N_615);
and U2031 (N_2031,N_1942,In_592);
xnor U2032 (N_2032,N_1975,N_1460);
nand U2033 (N_2033,N_1703,In_2209);
nor U2034 (N_2034,N_1324,N_1542);
and U2035 (N_2035,N_897,N_1724);
and U2036 (N_2036,In_1050,In_824);
nand U2037 (N_2037,N_124,N_1990);
xor U2038 (N_2038,N_1686,N_1196);
and U2039 (N_2039,N_1950,N_1752);
xnor U2040 (N_2040,N_1736,N_1572);
or U2041 (N_2041,N_721,In_888);
nor U2042 (N_2042,N_1645,In_1548);
and U2043 (N_2043,N_1891,In_2910);
and U2044 (N_2044,In_1969,N_1855);
and U2045 (N_2045,N_1874,In_2651);
or U2046 (N_2046,N_1731,N_1190);
nand U2047 (N_2047,N_1861,N_1615);
or U2048 (N_2048,N_1594,In_2144);
xor U2049 (N_2049,N_1226,N_1505);
and U2050 (N_2050,N_1538,N_1652);
or U2051 (N_2051,N_1568,N_1467);
nor U2052 (N_2052,N_1462,N_562);
xor U2053 (N_2053,N_1876,N_1801);
xor U2054 (N_2054,N_1725,N_1624);
xnor U2055 (N_2055,N_1044,N_1372);
xor U2056 (N_2056,N_1697,N_1982);
xor U2057 (N_2057,In_2171,N_1981);
or U2058 (N_2058,N_1292,N_1959);
xnor U2059 (N_2059,N_1642,N_1660);
nand U2060 (N_2060,N_1640,In_1575);
xor U2061 (N_2061,N_406,In_2642);
xnor U2062 (N_2062,N_1160,N_387);
and U2063 (N_2063,N_1699,N_1595);
or U2064 (N_2064,In_1008,N_1917);
nor U2065 (N_2065,N_682,In_1899);
and U2066 (N_2066,N_789,N_1169);
or U2067 (N_2067,N_1849,In_424);
and U2068 (N_2068,N_1549,N_769);
nand U2069 (N_2069,N_1961,N_458);
or U2070 (N_2070,In_2936,N_1718);
or U2071 (N_2071,N_1683,In_1419);
nand U2072 (N_2072,N_1214,N_1311);
xnor U2073 (N_2073,In_2583,In_2353);
xnor U2074 (N_2074,N_570,N_1767);
and U2075 (N_2075,N_1992,N_1188);
nor U2076 (N_2076,N_1860,N_1678);
xnor U2077 (N_2077,N_1812,N_1588);
nor U2078 (N_2078,N_672,N_131);
xnor U2079 (N_2079,N_807,N_1903);
nor U2080 (N_2080,N_1951,In_2068);
xor U2081 (N_2081,N_464,N_1313);
and U2082 (N_2082,In_2445,N_1753);
xor U2083 (N_2083,N_1375,N_1821);
and U2084 (N_2084,N_1185,N_635);
or U2085 (N_2085,N_255,N_1956);
or U2086 (N_2086,In_744,N_1648);
or U2087 (N_2087,In_1583,N_1713);
nor U2088 (N_2088,In_2366,N_1231);
nand U2089 (N_2089,N_1438,N_1464);
nand U2090 (N_2090,N_1074,N_1827);
and U2091 (N_2091,N_1916,N_1934);
and U2092 (N_2092,In_2321,N_1654);
xor U2093 (N_2093,N_1078,N_1807);
nand U2094 (N_2094,N_1358,N_1905);
nor U2095 (N_2095,N_1964,N_869);
nand U2096 (N_2096,N_1772,N_809);
nor U2097 (N_2097,N_1808,N_1977);
and U2098 (N_2098,N_1953,N_1970);
and U2099 (N_2099,N_1546,N_1868);
nand U2100 (N_2100,N_1189,N_1924);
nor U2101 (N_2101,In_2654,N_816);
and U2102 (N_2102,N_1760,N_1680);
xor U2103 (N_2103,N_1439,N_1665);
nor U2104 (N_2104,N_1565,N_26);
or U2105 (N_2105,In_2596,In_2207);
xor U2106 (N_2106,N_1649,N_1936);
nand U2107 (N_2107,N_83,In_2729);
and U2108 (N_2108,N_290,N_1719);
or U2109 (N_2109,N_1390,N_1087);
nand U2110 (N_2110,N_1514,N_1666);
xnor U2111 (N_2111,N_1525,N_1952);
or U2112 (N_2112,N_1495,In_1789);
and U2113 (N_2113,N_1480,N_1941);
or U2114 (N_2114,In_156,N_1973);
and U2115 (N_2115,N_1947,N_1564);
or U2116 (N_2116,N_1647,N_1627);
nor U2117 (N_2117,In_2758,N_1980);
or U2118 (N_2118,In_2153,N_554);
and U2119 (N_2119,N_1433,N_1693);
nand U2120 (N_2120,In_164,In_2733);
xnor U2121 (N_2121,N_237,N_1296);
and U2122 (N_2122,N_1684,In_742);
xor U2123 (N_2123,N_1790,N_1322);
nand U2124 (N_2124,N_1309,In_1787);
and U2125 (N_2125,N_1518,N_1191);
xor U2126 (N_2126,N_1730,In_45);
nand U2127 (N_2127,N_1544,N_1201);
and U2128 (N_2128,N_1509,N_1949);
and U2129 (N_2129,N_1271,In_2870);
xnor U2130 (N_2130,N_1974,In_1320);
and U2131 (N_2131,N_1583,N_650);
xnor U2132 (N_2132,In_532,In_456);
nand U2133 (N_2133,N_1561,N_1553);
and U2134 (N_2134,N_699,N_1816);
nor U2135 (N_2135,N_1701,N_1830);
nand U2136 (N_2136,N_1204,In_669);
or U2137 (N_2137,N_1857,N_1794);
nand U2138 (N_2138,N_1387,In_1633);
xnor U2139 (N_2139,N_1321,N_1235);
and U2140 (N_2140,N_748,N_1714);
nand U2141 (N_2141,In_805,N_1717);
nor U2142 (N_2142,N_1787,N_482);
nand U2143 (N_2143,N_346,N_1041);
nor U2144 (N_2144,N_1667,N_715);
nand U2145 (N_2145,N_704,N_1530);
and U2146 (N_2146,N_821,N_1835);
nor U2147 (N_2147,N_1210,In_2982);
or U2148 (N_2148,N_1779,N_1345);
and U2149 (N_2149,N_1674,N_1089);
nand U2150 (N_2150,In_382,N_1006);
xnor U2151 (N_2151,N_1853,N_1878);
xor U2152 (N_2152,In_271,N_1813);
nor U2153 (N_2153,N_1766,N_1550);
nor U2154 (N_2154,N_1630,N_1866);
nand U2155 (N_2155,In_1949,N_512);
and U2156 (N_2156,N_1176,N_1729);
xnor U2157 (N_2157,N_1075,N_1750);
nor U2158 (N_2158,N_1363,N_1043);
or U2159 (N_2159,In_861,N_1473);
nor U2160 (N_2160,In_911,N_1118);
and U2161 (N_2161,N_1580,N_1521);
nand U2162 (N_2162,N_1519,In_144);
or U2163 (N_2163,N_397,N_1673);
xor U2164 (N_2164,N_1331,In_1695);
or U2165 (N_2165,N_1862,N_106);
or U2166 (N_2166,N_620,N_1833);
and U2167 (N_2167,N_1798,N_1641);
or U2168 (N_2168,N_549,N_1743);
nor U2169 (N_2169,N_1377,In_2493);
and U2170 (N_2170,N_1744,N_1967);
and U2171 (N_2171,N_1969,N_1859);
nor U2172 (N_2172,N_796,N_1700);
nand U2173 (N_2173,N_1873,In_1204);
or U2174 (N_2174,N_1894,N_1838);
nand U2175 (N_2175,N_1935,N_1157);
xnor U2176 (N_2176,N_696,In_95);
nor U2177 (N_2177,N_1740,In_856);
xor U2178 (N_2178,N_1793,N_1851);
xor U2179 (N_2179,N_534,N_1883);
or U2180 (N_2180,N_614,N_1979);
nand U2181 (N_2181,N_1850,In_505);
or U2182 (N_2182,N_1955,N_1836);
or U2183 (N_2183,N_1877,N_1629);
and U2184 (N_2184,N_1479,N_1741);
xnor U2185 (N_2185,N_1571,In_1626);
nand U2186 (N_2186,N_1587,N_1014);
nor U2187 (N_2187,N_1303,N_1763);
and U2188 (N_2188,N_1893,N_1100);
nand U2189 (N_2189,In_2532,N_641);
nand U2190 (N_2190,N_22,N_1944);
nor U2191 (N_2191,N_244,N_986);
nor U2192 (N_2192,N_1477,N_1887);
and U2193 (N_2193,In_755,N_1971);
nor U2194 (N_2194,In_2181,In_78);
nor U2195 (N_2195,N_1778,N_1532);
nand U2196 (N_2196,In_490,N_1567);
and U2197 (N_2197,N_1259,N_1597);
nor U2198 (N_2198,N_817,In_788);
xnor U2199 (N_2199,N_1889,In_1991);
or U2200 (N_2200,N_1611,N_964);
nor U2201 (N_2201,N_1749,N_1581);
and U2202 (N_2202,N_1657,N_1799);
and U2203 (N_2203,N_1886,N_1511);
or U2204 (N_2204,N_1892,N_1599);
nand U2205 (N_2205,N_843,In_804);
or U2206 (N_2206,N_84,N_1715);
nand U2207 (N_2207,N_1895,N_1633);
nor U2208 (N_2208,N_1606,N_1913);
nor U2209 (N_2209,N_1869,N_1728);
nor U2210 (N_2210,N_1094,In_2588);
nand U2211 (N_2211,In_2747,N_1902);
or U2212 (N_2212,N_1884,N_1601);
or U2213 (N_2213,N_1854,N_860);
nor U2214 (N_2214,N_1593,N_1600);
and U2215 (N_2215,N_1656,N_1503);
nor U2216 (N_2216,N_1589,N_1609);
xor U2217 (N_2217,N_1682,N_1653);
and U2218 (N_2218,N_1991,N_1898);
or U2219 (N_2219,N_1508,N_1705);
xnor U2220 (N_2220,N_1081,N_1925);
or U2221 (N_2221,N_1584,N_1679);
nor U2222 (N_2222,In_1590,N_706);
and U2223 (N_2223,N_1136,N_1283);
or U2224 (N_2224,N_1528,N_801);
xor U2225 (N_2225,N_1819,N_1945);
or U2226 (N_2226,In_1460,In_1645);
xor U2227 (N_2227,N_1815,N_1659);
xor U2228 (N_2228,N_1053,In_1781);
or U2229 (N_2229,N_1543,N_485);
nor U2230 (N_2230,In_1926,N_1028);
xnor U2231 (N_2231,In_1032,N_861);
nand U2232 (N_2232,N_504,N_1608);
and U2233 (N_2233,In_619,N_1355);
xnor U2234 (N_2234,N_1134,N_1948);
or U2235 (N_2235,N_1986,In_1480);
nand U2236 (N_2236,N_1909,N_1052);
or U2237 (N_2237,In_423,N_422);
or U2238 (N_2238,N_1603,N_11);
or U2239 (N_2239,N_1848,In_2658);
nor U2240 (N_2240,In_538,In_618);
or U2241 (N_2241,N_1888,N_1285);
and U2242 (N_2242,N_1963,In_1505);
nor U2243 (N_2243,N_1761,N_1243);
xnor U2244 (N_2244,N_1732,N_1579);
nand U2245 (N_2245,In_975,N_1762);
or U2246 (N_2246,N_1317,N_580);
or U2247 (N_2247,N_1901,N_1796);
nand U2248 (N_2248,N_1747,N_1585);
nand U2249 (N_2249,N_1500,N_1586);
nand U2250 (N_2250,N_1636,N_1946);
or U2251 (N_2251,N_1037,N_1416);
or U2252 (N_2252,N_1146,N_1661);
and U2253 (N_2253,N_819,N_1806);
xor U2254 (N_2254,N_1605,N_1622);
xor U2255 (N_2255,N_1669,N_1708);
or U2256 (N_2256,N_376,N_1803);
xnor U2257 (N_2257,In_1512,In_933);
xor U2258 (N_2258,N_1738,N_1823);
nand U2259 (N_2259,N_1998,In_2753);
nor U2260 (N_2260,N_1675,N_1638);
or U2261 (N_2261,N_1938,In_2577);
nor U2262 (N_2262,N_1554,N_1631);
xor U2263 (N_2263,N_1576,N_1943);
or U2264 (N_2264,N_1880,In_261);
and U2265 (N_2265,N_1907,N_1560);
or U2266 (N_2266,N_1769,N_1172);
nor U2267 (N_2267,N_1734,N_804);
nor U2268 (N_2268,N_1958,N_1510);
and U2269 (N_2269,N_1773,In_2392);
nor U2270 (N_2270,N_390,N_1559);
nand U2271 (N_2271,N_1535,N_1707);
nand U2272 (N_2272,N_1828,N_1304);
or U2273 (N_2273,In_1392,N_1195);
nor U2274 (N_2274,N_310,In_2035);
xor U2275 (N_2275,In_1359,N_1482);
xnor U2276 (N_2276,N_1457,N_1987);
or U2277 (N_2277,N_1632,In_1620);
or U2278 (N_2278,N_1818,In_2745);
xnor U2279 (N_2279,In_2926,N_117);
nor U2280 (N_2280,N_1644,In_1780);
nor U2281 (N_2281,N_1098,N_1651);
xnor U2282 (N_2282,N_1775,N_1896);
nor U2283 (N_2283,N_1748,N_334);
xnor U2284 (N_2284,N_1501,N_343);
nand U2285 (N_2285,N_1620,N_895);
nor U2286 (N_2286,N_1751,N_1802);
xnor U2287 (N_2287,N_1484,N_1382);
xor U2288 (N_2288,N_1476,N_1551);
xor U2289 (N_2289,N_1832,N_1036);
nand U2290 (N_2290,In_0,N_956);
xor U2291 (N_2291,N_1937,N_1338);
nand U2292 (N_2292,In_626,N_1668);
nand U2293 (N_2293,N_1663,N_1918);
nand U2294 (N_2294,N_1272,N_1875);
xnor U2295 (N_2295,N_1655,N_1623);
or U2296 (N_2296,N_1695,N_1940);
nand U2297 (N_2297,N_1921,In_566);
xnor U2298 (N_2298,N_107,N_1116);
and U2299 (N_2299,N_1371,In_542);
and U2300 (N_2300,N_1612,N_1246);
nand U2301 (N_2301,N_1626,N_1822);
xnor U2302 (N_2302,N_1768,N_1403);
nand U2303 (N_2303,N_1920,N_855);
xor U2304 (N_2304,N_1915,N_1639);
or U2305 (N_2305,In_766,N_1121);
and U2306 (N_2306,N_1904,N_1531);
and U2307 (N_2307,N_1591,N_37);
nand U2308 (N_2308,N_1170,N_1512);
nor U2309 (N_2309,N_1523,N_1592);
xnor U2310 (N_2310,N_1451,N_1786);
or U2311 (N_2311,In_133,N_1820);
and U2312 (N_2312,N_1389,N_1545);
or U2313 (N_2313,In_438,In_2623);
nand U2314 (N_2314,N_1281,N_1088);
xnor U2315 (N_2315,In_1118,In_2487);
nand U2316 (N_2316,N_714,In_2298);
or U2317 (N_2317,N_1681,N_1694);
nor U2318 (N_2318,N_1993,N_1771);
xnor U2319 (N_2319,N_709,N_1025);
nand U2320 (N_2320,N_1008,N_19);
or U2321 (N_2321,N_545,N_29);
xor U2322 (N_2322,N_1972,N_1764);
xor U2323 (N_2323,N_1831,N_1294);
xor U2324 (N_2324,N_1881,N_1879);
nand U2325 (N_2325,N_1218,N_1804);
nor U2326 (N_2326,N_1702,N_1646);
or U2327 (N_2327,N_1625,N_648);
xnor U2328 (N_2328,N_309,N_1922);
and U2329 (N_2329,N_1997,N_1541);
nor U2330 (N_2330,In_2970,N_1960);
and U2331 (N_2331,N_1247,N_1706);
nand U2332 (N_2332,N_1005,In_595);
or U2333 (N_2333,N_1287,In_812);
and U2334 (N_2334,N_1614,N_936);
and U2335 (N_2335,N_1746,N_854);
or U2336 (N_2336,N_1557,N_877);
or U2337 (N_2337,N_1863,In_1335);
xnor U2338 (N_2338,In_1809,N_1619);
or U2339 (N_2339,N_1792,N_1757);
nor U2340 (N_2340,In_934,N_1381);
nor U2341 (N_2341,N_1284,In_2079);
nand U2342 (N_2342,In_2212,N_356);
nor U2343 (N_2343,N_1754,N_1346);
or U2344 (N_2344,In_580,N_655);
and U2345 (N_2345,N_1507,In_841);
and U2346 (N_2346,N_1578,N_987);
or U2347 (N_2347,N_1540,N_1575);
nand U2348 (N_2348,N_1520,N_1814);
or U2349 (N_2349,N_1841,N_1524);
and U2350 (N_2350,N_1152,In_1524);
xor U2351 (N_2351,N_1929,N_1988);
nand U2352 (N_2352,N_345,In_1256);
xnor U2353 (N_2353,N_448,N_1845);
nor U2354 (N_2354,N_53,N_657);
xor U2355 (N_2355,In_1400,N_1300);
nand U2356 (N_2356,N_1825,N_1711);
nand U2357 (N_2357,N_1726,N_76);
or U2358 (N_2358,N_1574,N_1526);
or U2359 (N_2359,N_1985,N_1784);
xnor U2360 (N_2360,N_1335,In_113);
nand U2361 (N_2361,In_2877,N_1582);
or U2362 (N_2362,N_1009,In_796);
and U2363 (N_2363,N_1536,N_1266);
nor U2364 (N_2364,N_1691,N_1219);
xor U2365 (N_2365,N_1870,In_341);
and U2366 (N_2366,N_1864,N_1954);
or U2367 (N_2367,N_1765,N_1658);
or U2368 (N_2368,N_1502,N_523);
nand U2369 (N_2369,N_1569,N_849);
nor U2370 (N_2370,In_17,N_889);
nand U2371 (N_2371,In_2784,N_1758);
nand U2372 (N_2372,N_1621,N_1897);
nor U2373 (N_2373,N_1872,N_1613);
nand U2374 (N_2374,N_1928,N_1852);
or U2375 (N_2375,N_1847,N_1785);
or U2376 (N_2376,N_1049,In_2001);
and U2377 (N_2377,N_1999,In_1240);
or U2378 (N_2378,N_1596,N_1995);
nor U2379 (N_2379,In_2031,N_1573);
or U2380 (N_2380,N_1932,N_1676);
or U2381 (N_2381,In_631,N_1696);
xnor U2382 (N_2382,N_1885,N_1692);
and U2383 (N_2383,In_940,N_1844);
nand U2384 (N_2384,N_952,In_2390);
and U2385 (N_2385,N_1023,In_2898);
and U2386 (N_2386,N_450,In_2200);
nand U2387 (N_2387,N_1145,N_1914);
nor U2388 (N_2388,N_1174,N_1968);
nand U2389 (N_2389,N_1858,N_1837);
xor U2390 (N_2390,N_1312,N_1397);
nor U2391 (N_2391,N_1225,N_1672);
or U2392 (N_2392,N_1933,N_1341);
and U2393 (N_2393,N_1811,N_1604);
or U2394 (N_2394,N_1437,N_1029);
xnor U2395 (N_2395,N_871,N_1602);
nor U2396 (N_2396,In_2365,N_1240);
and U2397 (N_2397,N_1927,N_1108);
xnor U2398 (N_2398,N_1797,N_1664);
or U2399 (N_2399,N_1249,In_2061);
nor U2400 (N_2400,N_1670,In_84);
nor U2401 (N_2401,In_1611,N_745);
xor U2402 (N_2402,N_1187,N_1068);
nor U2403 (N_2403,N_1782,In_1852);
and U2404 (N_2404,N_1529,N_1418);
nor U2405 (N_2405,N_1906,In_2047);
nand U2406 (N_2406,N_1516,N_1776);
xnor U2407 (N_2407,N_870,N_1504);
and U2408 (N_2408,N_1867,N_1984);
and U2409 (N_2409,N_1562,N_1733);
xnor U2410 (N_2410,N_286,N_1590);
nor U2411 (N_2411,In_2335,N_1856);
nor U2412 (N_2412,N_1791,N_1517);
nor U2413 (N_2413,In_292,In_1329);
xor U2414 (N_2414,In_1844,N_1957);
and U2415 (N_2415,N_1024,N_1026);
xor U2416 (N_2416,N_1577,N_1840);
and U2417 (N_2417,N_1899,N_1635);
and U2418 (N_2418,N_1780,N_1978);
and U2419 (N_2419,In_2549,In_1233);
nor U2420 (N_2420,N_1388,In_1535);
nor U2421 (N_2421,N_1865,N_1742);
and U2422 (N_2422,In_2692,N_1506);
nand U2423 (N_2423,In_1752,N_939);
nor U2424 (N_2424,In_1197,N_1810);
nand U2425 (N_2425,In_2219,In_972);
and U2426 (N_2426,In_1906,N_1329);
xnor U2427 (N_2427,N_1643,N_276);
xor U2428 (N_2428,N_1989,N_1610);
nand U2429 (N_2429,N_1966,In_2755);
xor U2430 (N_2430,N_1688,N_1809);
and U2431 (N_2431,N_1723,N_1547);
xnor U2432 (N_2432,N_1359,In_727);
xnor U2433 (N_2433,N_1035,In_1581);
or U2434 (N_2434,In_1064,In_2444);
nor U2435 (N_2435,N_1839,In_1716);
nor U2436 (N_2436,N_642,In_415);
and U2437 (N_2437,N_1826,N_1795);
nor U2438 (N_2438,N_462,N_1373);
and U2439 (N_2439,N_1983,In_79);
nand U2440 (N_2440,In_760,N_1515);
or U2441 (N_2441,In_2264,N_1111);
or U2442 (N_2442,N_1534,In_776);
nand U2443 (N_2443,N_1072,N_192);
xor U2444 (N_2444,In_458,N_1710);
nand U2445 (N_2445,N_1327,N_1555);
or U2446 (N_2446,N_1939,In_1821);
nand U2447 (N_2447,In_1896,N_1628);
and U2448 (N_2448,N_525,N_1781);
and U2449 (N_2449,N_1552,In_1336);
xor U2450 (N_2450,N_1513,In_1142);
xor U2451 (N_2451,N_1912,In_2688);
or U2452 (N_2452,In_391,N_1996);
or U2453 (N_2453,N_1193,N_1908);
nor U2454 (N_2454,N_1871,N_1001);
xor U2455 (N_2455,In_1895,N_1727);
nand U2456 (N_2456,N_1685,N_1106);
nand U2457 (N_2457,N_1777,N_1069);
and U2458 (N_2458,In_2632,N_585);
and U2459 (N_2459,N_1923,N_1704);
or U2460 (N_2460,N_886,N_1086);
xnor U2461 (N_2461,In_1354,N_1634);
or U2462 (N_2462,N_884,N_1637);
xor U2463 (N_2463,N_1919,N_1755);
nand U2464 (N_2464,N_1698,N_1900);
or U2465 (N_2465,In_2553,N_1548);
nor U2466 (N_2466,N_218,N_1930);
nor U2467 (N_2467,In_2033,N_1687);
and U2468 (N_2468,N_1843,In_93);
xor U2469 (N_2469,In_787,N_1070);
or U2470 (N_2470,N_1155,N_1206);
or U2471 (N_2471,In_2795,N_1842);
nand U2472 (N_2472,N_1522,N_1745);
or U2473 (N_2473,N_1570,N_1323);
nor U2474 (N_2474,N_1735,N_1910);
and U2475 (N_2475,N_1492,N_1429);
xnor U2476 (N_2476,N_1965,N_1454);
xor U2477 (N_2477,N_1846,In_2421);
xor U2478 (N_2478,In_327,N_1114);
nor U2479 (N_2479,N_1911,N_1834);
nor U2480 (N_2480,N_1566,N_822);
and U2481 (N_2481,N_1065,N_1783);
xor U2482 (N_2482,In_1363,In_99);
nor U2483 (N_2483,In_900,N_1241);
xnor U2484 (N_2484,N_1527,N_1496);
xnor U2485 (N_2485,In_2819,N_1720);
xnor U2486 (N_2486,N_1962,N_1618);
or U2487 (N_2487,In_2433,N_873);
and U2488 (N_2488,N_1829,N_1774);
nor U2489 (N_2489,N_681,N_1342);
xnor U2490 (N_2490,In_2225,In_1291);
or U2491 (N_2491,N_1722,In_194);
nand U2492 (N_2492,In_2273,N_1332);
and U2493 (N_2493,N_1095,N_7);
and U2494 (N_2494,N_887,N_1817);
or U2495 (N_2495,In_2389,N_1976);
or U2496 (N_2496,In_1136,N_1607);
and U2497 (N_2497,N_1367,In_964);
nor U2498 (N_2498,N_1759,N_1650);
xnor U2499 (N_2499,N_1481,In_2053);
or U2500 (N_2500,N_2386,N_2446);
nor U2501 (N_2501,N_2192,N_2339);
or U2502 (N_2502,N_2270,N_2186);
nor U2503 (N_2503,N_2040,N_2450);
nor U2504 (N_2504,N_2309,N_2350);
and U2505 (N_2505,N_2373,N_2012);
and U2506 (N_2506,N_2437,N_2301);
or U2507 (N_2507,N_2008,N_2006);
or U2508 (N_2508,N_2380,N_2110);
xor U2509 (N_2509,N_2478,N_2086);
and U2510 (N_2510,N_2062,N_2133);
and U2511 (N_2511,N_2362,N_2410);
xor U2512 (N_2512,N_2498,N_2223);
or U2513 (N_2513,N_2208,N_2112);
nand U2514 (N_2514,N_2003,N_2232);
xnor U2515 (N_2515,N_2409,N_2418);
nor U2516 (N_2516,N_2374,N_2319);
nor U2517 (N_2517,N_2294,N_2162);
xnor U2518 (N_2518,N_2318,N_2233);
and U2519 (N_2519,N_2447,N_2397);
xnor U2520 (N_2520,N_2060,N_2177);
xnor U2521 (N_2521,N_2475,N_2211);
and U2522 (N_2522,N_2368,N_2360);
nor U2523 (N_2523,N_2336,N_2351);
nand U2524 (N_2524,N_2058,N_2050);
nand U2525 (N_2525,N_2170,N_2462);
and U2526 (N_2526,N_2023,N_2343);
nor U2527 (N_2527,N_2458,N_2399);
xnor U2528 (N_2528,N_2004,N_2353);
nor U2529 (N_2529,N_2115,N_2087);
nor U2530 (N_2530,N_2005,N_2098);
nand U2531 (N_2531,N_2202,N_2455);
and U2532 (N_2532,N_2069,N_2246);
xnor U2533 (N_2533,N_2030,N_2381);
and U2534 (N_2534,N_2103,N_2039);
and U2535 (N_2535,N_2032,N_2075);
xor U2536 (N_2536,N_2476,N_2491);
nand U2537 (N_2537,N_2026,N_2416);
xnor U2538 (N_2538,N_2452,N_2434);
or U2539 (N_2539,N_2097,N_2401);
xor U2540 (N_2540,N_2010,N_2147);
nor U2541 (N_2541,N_2481,N_2303);
xor U2542 (N_2542,N_2390,N_2337);
or U2543 (N_2543,N_2290,N_2364);
xor U2544 (N_2544,N_2099,N_2366);
nand U2545 (N_2545,N_2449,N_2304);
and U2546 (N_2546,N_2421,N_2258);
and U2547 (N_2547,N_2033,N_2090);
xor U2548 (N_2548,N_2457,N_2411);
nor U2549 (N_2549,N_2013,N_2260);
or U2550 (N_2550,N_2245,N_2148);
nor U2551 (N_2551,N_2348,N_2046);
or U2552 (N_2552,N_2247,N_2145);
nor U2553 (N_2553,N_2089,N_2044);
and U2554 (N_2554,N_2018,N_2106);
or U2555 (N_2555,N_2150,N_2102);
nor U2556 (N_2556,N_2468,N_2376);
nor U2557 (N_2557,N_2073,N_2173);
nand U2558 (N_2558,N_2315,N_2370);
or U2559 (N_2559,N_2101,N_2430);
xor U2560 (N_2560,N_2190,N_2466);
nand U2561 (N_2561,N_2007,N_2414);
and U2562 (N_2562,N_2083,N_2474);
nor U2563 (N_2563,N_2029,N_2287);
nand U2564 (N_2564,N_2234,N_2194);
nor U2565 (N_2565,N_2307,N_2250);
and U2566 (N_2566,N_2454,N_2469);
nor U2567 (N_2567,N_2059,N_2182);
or U2568 (N_2568,N_2499,N_2436);
xor U2569 (N_2569,N_2000,N_2482);
xnor U2570 (N_2570,N_2225,N_2077);
xnor U2571 (N_2571,N_2117,N_2407);
and U2572 (N_2572,N_2220,N_2057);
or U2573 (N_2573,N_2358,N_2043);
nand U2574 (N_2574,N_2313,N_2453);
and U2575 (N_2575,N_2181,N_2355);
and U2576 (N_2576,N_2009,N_2396);
nor U2577 (N_2577,N_2428,N_2329);
nand U2578 (N_2578,N_2078,N_2398);
or U2579 (N_2579,N_2438,N_2308);
nand U2580 (N_2580,N_2252,N_2174);
or U2581 (N_2581,N_2331,N_2126);
and U2582 (N_2582,N_2152,N_2203);
nand U2583 (N_2583,N_2072,N_2393);
xor U2584 (N_2584,N_2094,N_2274);
and U2585 (N_2585,N_2306,N_2142);
and U2586 (N_2586,N_2022,N_2465);
nor U2587 (N_2587,N_2104,N_2459);
and U2588 (N_2588,N_2317,N_2338);
or U2589 (N_2589,N_2259,N_2066);
or U2590 (N_2590,N_2493,N_2347);
and U2591 (N_2591,N_2253,N_2172);
or U2592 (N_2592,N_2257,N_2034);
xor U2593 (N_2593,N_2121,N_2240);
xor U2594 (N_2594,N_2445,N_2391);
and U2595 (N_2595,N_2357,N_2167);
or U2596 (N_2596,N_2118,N_2199);
nand U2597 (N_2597,N_2156,N_2100);
nand U2598 (N_2598,N_2189,N_2014);
xnor U2599 (N_2599,N_2065,N_2328);
or U2600 (N_2600,N_2201,N_2180);
xnor U2601 (N_2601,N_2345,N_2127);
or U2602 (N_2602,N_2141,N_2042);
xnor U2603 (N_2603,N_2011,N_2496);
nand U2604 (N_2604,N_2241,N_2316);
or U2605 (N_2605,N_2432,N_2282);
and U2606 (N_2606,N_2324,N_2385);
xor U2607 (N_2607,N_2333,N_2206);
xor U2608 (N_2608,N_2144,N_2486);
nor U2609 (N_2609,N_2489,N_2367);
and U2610 (N_2610,N_2064,N_2433);
and U2611 (N_2611,N_2471,N_2213);
nand U2612 (N_2612,N_2425,N_2344);
nor U2613 (N_2613,N_2131,N_2405);
nor U2614 (N_2614,N_2095,N_2485);
and U2615 (N_2615,N_2214,N_2420);
nand U2616 (N_2616,N_2431,N_2284);
nor U2617 (N_2617,N_2487,N_2239);
and U2618 (N_2618,N_2280,N_2265);
xnor U2619 (N_2619,N_2184,N_2268);
nand U2620 (N_2620,N_2341,N_2175);
nand U2621 (N_2621,N_2116,N_2204);
xnor U2622 (N_2622,N_2479,N_2429);
and U2623 (N_2623,N_2249,N_2419);
or U2624 (N_2624,N_2488,N_2224);
nand U2625 (N_2625,N_2404,N_2400);
and U2626 (N_2626,N_2153,N_2051);
and U2627 (N_2627,N_2056,N_2132);
nor U2628 (N_2628,N_2129,N_2084);
xnor U2629 (N_2629,N_2179,N_2076);
nand U2630 (N_2630,N_2169,N_2166);
xor U2631 (N_2631,N_2025,N_2299);
xor U2632 (N_2632,N_2384,N_2114);
nor U2633 (N_2633,N_2359,N_2061);
nand U2634 (N_2634,N_2226,N_2235);
and U2635 (N_2635,N_2130,N_2314);
nand U2636 (N_2636,N_2467,N_2382);
or U2637 (N_2637,N_2251,N_2305);
nor U2638 (N_2638,N_2231,N_2417);
or U2639 (N_2639,N_2352,N_2472);
nor U2640 (N_2640,N_2222,N_2365);
or U2641 (N_2641,N_2266,N_2038);
or U2642 (N_2642,N_2426,N_2293);
and U2643 (N_2643,N_2406,N_2081);
or U2644 (N_2644,N_2016,N_2295);
or U2645 (N_2645,N_2334,N_2326);
and U2646 (N_2646,N_2377,N_2372);
or U2647 (N_2647,N_2219,N_2191);
or U2648 (N_2648,N_2047,N_2238);
nand U2649 (N_2649,N_2197,N_2085);
and U2650 (N_2650,N_2278,N_2441);
xnor U2651 (N_2651,N_2041,N_2490);
and U2652 (N_2652,N_2332,N_2158);
xor U2653 (N_2653,N_2125,N_2248);
xnor U2654 (N_2654,N_2019,N_2124);
nand U2655 (N_2655,N_2160,N_2155);
or U2656 (N_2656,N_2375,N_2298);
xnor U2657 (N_2657,N_2070,N_2193);
nor U2658 (N_2658,N_2477,N_2024);
and U2659 (N_2659,N_2448,N_2164);
nand U2660 (N_2660,N_2207,N_2091);
nor U2661 (N_2661,N_2264,N_2212);
xnor U2662 (N_2662,N_2276,N_2052);
xnor U2663 (N_2663,N_2310,N_2273);
or U2664 (N_2664,N_2335,N_2342);
or U2665 (N_2665,N_2288,N_2187);
or U2666 (N_2666,N_2451,N_2346);
and U2667 (N_2667,N_2463,N_2111);
nand U2668 (N_2668,N_2218,N_2045);
and U2669 (N_2669,N_2484,N_2302);
nand U2670 (N_2670,N_2140,N_2230);
and U2671 (N_2671,N_2296,N_2237);
nand U2672 (N_2672,N_2378,N_2267);
and U2673 (N_2673,N_2210,N_2063);
nor U2674 (N_2674,N_2483,N_2183);
or U2675 (N_2675,N_2443,N_2320);
and U2676 (N_2676,N_2093,N_2027);
xnor U2677 (N_2677,N_2205,N_2105);
and U2678 (N_2678,N_2163,N_2200);
and U2679 (N_2679,N_2456,N_2311);
nor U2680 (N_2680,N_2082,N_2254);
and U2681 (N_2681,N_2263,N_2137);
xnor U2682 (N_2682,N_2439,N_2154);
nand U2683 (N_2683,N_2227,N_2229);
xor U2684 (N_2684,N_2107,N_2113);
xor U2685 (N_2685,N_2242,N_2464);
xor U2686 (N_2686,N_2327,N_2470);
nor U2687 (N_2687,N_2291,N_2143);
and U2688 (N_2688,N_2256,N_2262);
and U2689 (N_2689,N_2289,N_2387);
and U2690 (N_2690,N_2389,N_2074);
and U2691 (N_2691,N_2035,N_2415);
nand U2692 (N_2692,N_2497,N_2427);
xnor U2693 (N_2693,N_2171,N_2067);
and U2694 (N_2694,N_2053,N_2340);
or U2695 (N_2695,N_2403,N_2123);
xor U2696 (N_2696,N_2198,N_2388);
and U2697 (N_2697,N_2321,N_2031);
or U2698 (N_2698,N_2176,N_2136);
or U2699 (N_2699,N_2139,N_2216);
or U2700 (N_2700,N_2215,N_2149);
nor U2701 (N_2701,N_2244,N_2178);
nor U2702 (N_2702,N_2383,N_2300);
nor U2703 (N_2703,N_2394,N_2435);
xor U2704 (N_2704,N_2379,N_2460);
nand U2705 (N_2705,N_2188,N_2422);
nand U2706 (N_2706,N_2236,N_2272);
xnor U2707 (N_2707,N_2195,N_2395);
nor U2708 (N_2708,N_2015,N_2269);
or U2709 (N_2709,N_2279,N_2138);
xor U2710 (N_2710,N_2292,N_2096);
and U2711 (N_2711,N_2330,N_2283);
nor U2712 (N_2712,N_2323,N_2349);
or U2713 (N_2713,N_2440,N_2495);
nor U2714 (N_2714,N_2228,N_2255);
nand U2715 (N_2715,N_2281,N_2088);
xor U2716 (N_2716,N_2261,N_2363);
nor U2717 (N_2717,N_2028,N_2017);
and U2718 (N_2718,N_2120,N_2494);
and U2719 (N_2719,N_2161,N_2135);
nor U2720 (N_2720,N_2275,N_2054);
and U2721 (N_2721,N_2196,N_2165);
and U2722 (N_2722,N_2048,N_2297);
xnor U2723 (N_2723,N_2277,N_2271);
and U2724 (N_2724,N_2356,N_2442);
nor U2725 (N_2725,N_2369,N_2402);
and U2726 (N_2726,N_2217,N_2209);
nand U2727 (N_2727,N_2312,N_2285);
nor U2728 (N_2728,N_2286,N_2021);
and U2729 (N_2729,N_2325,N_2157);
and U2730 (N_2730,N_2080,N_2322);
xor U2731 (N_2731,N_2020,N_2424);
nand U2732 (N_2732,N_2068,N_2159);
nor U2733 (N_2733,N_2146,N_2444);
and U2734 (N_2734,N_2221,N_2109);
and U2735 (N_2735,N_2461,N_2079);
xnor U2736 (N_2736,N_2492,N_2480);
and U2737 (N_2737,N_2108,N_2392);
and U2738 (N_2738,N_2371,N_2122);
or U2739 (N_2739,N_2423,N_2055);
or U2740 (N_2740,N_2168,N_2049);
nor U2741 (N_2741,N_2036,N_2413);
xnor U2742 (N_2742,N_2243,N_2408);
nor U2743 (N_2743,N_2001,N_2361);
nand U2744 (N_2744,N_2354,N_2002);
xnor U2745 (N_2745,N_2092,N_2119);
xor U2746 (N_2746,N_2037,N_2151);
or U2747 (N_2747,N_2134,N_2185);
xor U2748 (N_2748,N_2071,N_2128);
nor U2749 (N_2749,N_2473,N_2412);
nor U2750 (N_2750,N_2319,N_2044);
xor U2751 (N_2751,N_2488,N_2205);
and U2752 (N_2752,N_2126,N_2340);
nor U2753 (N_2753,N_2131,N_2314);
nor U2754 (N_2754,N_2069,N_2237);
xnor U2755 (N_2755,N_2015,N_2194);
nor U2756 (N_2756,N_2317,N_2113);
or U2757 (N_2757,N_2378,N_2250);
xnor U2758 (N_2758,N_2131,N_2079);
nor U2759 (N_2759,N_2157,N_2119);
or U2760 (N_2760,N_2207,N_2120);
and U2761 (N_2761,N_2223,N_2282);
nor U2762 (N_2762,N_2078,N_2282);
nand U2763 (N_2763,N_2206,N_2142);
nor U2764 (N_2764,N_2299,N_2110);
and U2765 (N_2765,N_2453,N_2380);
nand U2766 (N_2766,N_2025,N_2168);
or U2767 (N_2767,N_2486,N_2303);
and U2768 (N_2768,N_2434,N_2345);
nand U2769 (N_2769,N_2479,N_2308);
and U2770 (N_2770,N_2121,N_2096);
and U2771 (N_2771,N_2347,N_2427);
xnor U2772 (N_2772,N_2084,N_2204);
nand U2773 (N_2773,N_2138,N_2055);
and U2774 (N_2774,N_2026,N_2497);
xnor U2775 (N_2775,N_2489,N_2121);
or U2776 (N_2776,N_2469,N_2317);
and U2777 (N_2777,N_2497,N_2169);
nand U2778 (N_2778,N_2128,N_2117);
and U2779 (N_2779,N_2174,N_2363);
or U2780 (N_2780,N_2451,N_2379);
or U2781 (N_2781,N_2173,N_2469);
xnor U2782 (N_2782,N_2188,N_2180);
xnor U2783 (N_2783,N_2137,N_2354);
nor U2784 (N_2784,N_2417,N_2481);
xor U2785 (N_2785,N_2206,N_2017);
nor U2786 (N_2786,N_2214,N_2311);
nor U2787 (N_2787,N_2256,N_2122);
nand U2788 (N_2788,N_2200,N_2197);
nor U2789 (N_2789,N_2036,N_2058);
and U2790 (N_2790,N_2110,N_2302);
or U2791 (N_2791,N_2249,N_2423);
nand U2792 (N_2792,N_2253,N_2109);
nand U2793 (N_2793,N_2406,N_2249);
or U2794 (N_2794,N_2123,N_2165);
nand U2795 (N_2795,N_2192,N_2200);
nand U2796 (N_2796,N_2084,N_2210);
xnor U2797 (N_2797,N_2439,N_2398);
nor U2798 (N_2798,N_2333,N_2039);
and U2799 (N_2799,N_2356,N_2302);
and U2800 (N_2800,N_2033,N_2487);
xor U2801 (N_2801,N_2084,N_2324);
or U2802 (N_2802,N_2036,N_2353);
or U2803 (N_2803,N_2209,N_2263);
nand U2804 (N_2804,N_2217,N_2097);
nand U2805 (N_2805,N_2461,N_2327);
or U2806 (N_2806,N_2320,N_2234);
nor U2807 (N_2807,N_2463,N_2262);
or U2808 (N_2808,N_2275,N_2019);
nor U2809 (N_2809,N_2227,N_2370);
and U2810 (N_2810,N_2112,N_2091);
and U2811 (N_2811,N_2439,N_2301);
xnor U2812 (N_2812,N_2240,N_2462);
or U2813 (N_2813,N_2273,N_2245);
nand U2814 (N_2814,N_2216,N_2225);
nor U2815 (N_2815,N_2398,N_2375);
and U2816 (N_2816,N_2499,N_2453);
xor U2817 (N_2817,N_2121,N_2339);
nand U2818 (N_2818,N_2112,N_2115);
xnor U2819 (N_2819,N_2388,N_2077);
xnor U2820 (N_2820,N_2137,N_2293);
nor U2821 (N_2821,N_2462,N_2192);
nand U2822 (N_2822,N_2461,N_2292);
or U2823 (N_2823,N_2101,N_2367);
xnor U2824 (N_2824,N_2169,N_2225);
xnor U2825 (N_2825,N_2236,N_2477);
or U2826 (N_2826,N_2291,N_2180);
nand U2827 (N_2827,N_2150,N_2423);
nand U2828 (N_2828,N_2172,N_2438);
xor U2829 (N_2829,N_2341,N_2352);
and U2830 (N_2830,N_2063,N_2226);
or U2831 (N_2831,N_2039,N_2092);
and U2832 (N_2832,N_2241,N_2376);
nand U2833 (N_2833,N_2366,N_2442);
nand U2834 (N_2834,N_2077,N_2020);
or U2835 (N_2835,N_2040,N_2106);
xor U2836 (N_2836,N_2271,N_2386);
or U2837 (N_2837,N_2477,N_2288);
and U2838 (N_2838,N_2489,N_2469);
nand U2839 (N_2839,N_2056,N_2486);
nand U2840 (N_2840,N_2352,N_2144);
nand U2841 (N_2841,N_2269,N_2394);
and U2842 (N_2842,N_2496,N_2366);
or U2843 (N_2843,N_2417,N_2449);
or U2844 (N_2844,N_2158,N_2331);
nand U2845 (N_2845,N_2097,N_2199);
or U2846 (N_2846,N_2172,N_2281);
nor U2847 (N_2847,N_2019,N_2120);
or U2848 (N_2848,N_2385,N_2419);
and U2849 (N_2849,N_2113,N_2358);
or U2850 (N_2850,N_2320,N_2017);
and U2851 (N_2851,N_2413,N_2061);
xnor U2852 (N_2852,N_2393,N_2279);
or U2853 (N_2853,N_2010,N_2286);
or U2854 (N_2854,N_2172,N_2399);
xnor U2855 (N_2855,N_2103,N_2078);
nor U2856 (N_2856,N_2134,N_2395);
nand U2857 (N_2857,N_2069,N_2272);
and U2858 (N_2858,N_2348,N_2340);
or U2859 (N_2859,N_2386,N_2382);
nor U2860 (N_2860,N_2478,N_2005);
and U2861 (N_2861,N_2021,N_2424);
nand U2862 (N_2862,N_2477,N_2283);
and U2863 (N_2863,N_2098,N_2069);
or U2864 (N_2864,N_2498,N_2040);
or U2865 (N_2865,N_2249,N_2197);
or U2866 (N_2866,N_2265,N_2222);
nand U2867 (N_2867,N_2140,N_2156);
xnor U2868 (N_2868,N_2261,N_2110);
and U2869 (N_2869,N_2045,N_2217);
xnor U2870 (N_2870,N_2339,N_2223);
nand U2871 (N_2871,N_2434,N_2230);
nand U2872 (N_2872,N_2397,N_2154);
xor U2873 (N_2873,N_2168,N_2322);
nor U2874 (N_2874,N_2300,N_2313);
xnor U2875 (N_2875,N_2389,N_2449);
and U2876 (N_2876,N_2220,N_2399);
and U2877 (N_2877,N_2019,N_2000);
nand U2878 (N_2878,N_2013,N_2278);
nor U2879 (N_2879,N_2175,N_2028);
and U2880 (N_2880,N_2155,N_2013);
nor U2881 (N_2881,N_2000,N_2486);
nor U2882 (N_2882,N_2300,N_2222);
xor U2883 (N_2883,N_2047,N_2494);
or U2884 (N_2884,N_2142,N_2274);
nor U2885 (N_2885,N_2376,N_2004);
and U2886 (N_2886,N_2434,N_2000);
and U2887 (N_2887,N_2068,N_2345);
nor U2888 (N_2888,N_2362,N_2155);
xor U2889 (N_2889,N_2278,N_2473);
nor U2890 (N_2890,N_2300,N_2447);
or U2891 (N_2891,N_2069,N_2261);
and U2892 (N_2892,N_2315,N_2230);
and U2893 (N_2893,N_2012,N_2321);
or U2894 (N_2894,N_2321,N_2210);
nor U2895 (N_2895,N_2456,N_2467);
and U2896 (N_2896,N_2442,N_2003);
or U2897 (N_2897,N_2351,N_2142);
and U2898 (N_2898,N_2480,N_2358);
nor U2899 (N_2899,N_2045,N_2406);
xnor U2900 (N_2900,N_2397,N_2252);
nand U2901 (N_2901,N_2222,N_2479);
and U2902 (N_2902,N_2116,N_2360);
and U2903 (N_2903,N_2353,N_2229);
and U2904 (N_2904,N_2405,N_2116);
or U2905 (N_2905,N_2343,N_2273);
nor U2906 (N_2906,N_2172,N_2258);
and U2907 (N_2907,N_2213,N_2040);
or U2908 (N_2908,N_2115,N_2497);
nand U2909 (N_2909,N_2338,N_2150);
or U2910 (N_2910,N_2182,N_2355);
nand U2911 (N_2911,N_2352,N_2390);
xnor U2912 (N_2912,N_2220,N_2152);
and U2913 (N_2913,N_2435,N_2237);
or U2914 (N_2914,N_2395,N_2152);
xnor U2915 (N_2915,N_2134,N_2372);
nor U2916 (N_2916,N_2257,N_2346);
and U2917 (N_2917,N_2308,N_2329);
xnor U2918 (N_2918,N_2017,N_2346);
xor U2919 (N_2919,N_2284,N_2041);
and U2920 (N_2920,N_2225,N_2337);
or U2921 (N_2921,N_2074,N_2136);
nor U2922 (N_2922,N_2413,N_2307);
nand U2923 (N_2923,N_2097,N_2309);
nand U2924 (N_2924,N_2473,N_2109);
xor U2925 (N_2925,N_2419,N_2087);
and U2926 (N_2926,N_2113,N_2344);
and U2927 (N_2927,N_2059,N_2377);
or U2928 (N_2928,N_2362,N_2416);
and U2929 (N_2929,N_2448,N_2020);
or U2930 (N_2930,N_2462,N_2202);
nor U2931 (N_2931,N_2231,N_2037);
or U2932 (N_2932,N_2452,N_2258);
nor U2933 (N_2933,N_2230,N_2008);
nand U2934 (N_2934,N_2182,N_2016);
xor U2935 (N_2935,N_2372,N_2220);
nand U2936 (N_2936,N_2486,N_2409);
xnor U2937 (N_2937,N_2400,N_2475);
and U2938 (N_2938,N_2428,N_2386);
nand U2939 (N_2939,N_2031,N_2190);
nand U2940 (N_2940,N_2370,N_2039);
or U2941 (N_2941,N_2248,N_2129);
nand U2942 (N_2942,N_2120,N_2237);
or U2943 (N_2943,N_2304,N_2177);
and U2944 (N_2944,N_2184,N_2316);
nand U2945 (N_2945,N_2432,N_2247);
nor U2946 (N_2946,N_2410,N_2268);
nand U2947 (N_2947,N_2444,N_2231);
xor U2948 (N_2948,N_2356,N_2352);
and U2949 (N_2949,N_2000,N_2248);
or U2950 (N_2950,N_2160,N_2470);
or U2951 (N_2951,N_2288,N_2136);
nor U2952 (N_2952,N_2365,N_2236);
and U2953 (N_2953,N_2005,N_2475);
or U2954 (N_2954,N_2250,N_2345);
and U2955 (N_2955,N_2254,N_2376);
xor U2956 (N_2956,N_2341,N_2316);
and U2957 (N_2957,N_2119,N_2343);
nand U2958 (N_2958,N_2202,N_2019);
or U2959 (N_2959,N_2161,N_2413);
nor U2960 (N_2960,N_2202,N_2279);
nand U2961 (N_2961,N_2330,N_2057);
nand U2962 (N_2962,N_2344,N_2284);
nor U2963 (N_2963,N_2485,N_2280);
nor U2964 (N_2964,N_2388,N_2317);
nand U2965 (N_2965,N_2240,N_2012);
and U2966 (N_2966,N_2075,N_2383);
and U2967 (N_2967,N_2422,N_2471);
nor U2968 (N_2968,N_2405,N_2073);
nor U2969 (N_2969,N_2027,N_2439);
nor U2970 (N_2970,N_2058,N_2042);
nor U2971 (N_2971,N_2371,N_2327);
or U2972 (N_2972,N_2240,N_2185);
and U2973 (N_2973,N_2316,N_2081);
xnor U2974 (N_2974,N_2106,N_2332);
and U2975 (N_2975,N_2458,N_2355);
nand U2976 (N_2976,N_2420,N_2241);
and U2977 (N_2977,N_2148,N_2063);
and U2978 (N_2978,N_2237,N_2045);
nor U2979 (N_2979,N_2164,N_2180);
xnor U2980 (N_2980,N_2180,N_2112);
or U2981 (N_2981,N_2004,N_2385);
or U2982 (N_2982,N_2235,N_2180);
xor U2983 (N_2983,N_2364,N_2409);
and U2984 (N_2984,N_2447,N_2045);
xor U2985 (N_2985,N_2084,N_2313);
nand U2986 (N_2986,N_2334,N_2287);
nand U2987 (N_2987,N_2170,N_2329);
nor U2988 (N_2988,N_2028,N_2345);
nor U2989 (N_2989,N_2400,N_2022);
or U2990 (N_2990,N_2396,N_2056);
nand U2991 (N_2991,N_2031,N_2246);
xnor U2992 (N_2992,N_2098,N_2123);
and U2993 (N_2993,N_2148,N_2008);
and U2994 (N_2994,N_2235,N_2074);
and U2995 (N_2995,N_2374,N_2291);
nor U2996 (N_2996,N_2222,N_2418);
or U2997 (N_2997,N_2389,N_2171);
or U2998 (N_2998,N_2139,N_2391);
and U2999 (N_2999,N_2151,N_2252);
or U3000 (N_3000,N_2956,N_2806);
xnor U3001 (N_3001,N_2730,N_2649);
or U3002 (N_3002,N_2713,N_2952);
and U3003 (N_3003,N_2567,N_2736);
xor U3004 (N_3004,N_2845,N_2578);
nand U3005 (N_3005,N_2962,N_2784);
and U3006 (N_3006,N_2528,N_2864);
and U3007 (N_3007,N_2570,N_2771);
nand U3008 (N_3008,N_2708,N_2773);
nand U3009 (N_3009,N_2986,N_2929);
or U3010 (N_3010,N_2810,N_2698);
nor U3011 (N_3011,N_2853,N_2761);
or U3012 (N_3012,N_2823,N_2748);
nor U3013 (N_3013,N_2840,N_2506);
nand U3014 (N_3014,N_2740,N_2620);
and U3015 (N_3015,N_2547,N_2804);
nor U3016 (N_3016,N_2818,N_2747);
xnor U3017 (N_3017,N_2821,N_2731);
nor U3018 (N_3018,N_2874,N_2769);
and U3019 (N_3019,N_2941,N_2777);
xor U3020 (N_3020,N_2607,N_2930);
nor U3021 (N_3021,N_2944,N_2583);
nand U3022 (N_3022,N_2861,N_2873);
and U3023 (N_3023,N_2969,N_2641);
nor U3024 (N_3024,N_2989,N_2838);
and U3025 (N_3025,N_2917,N_2671);
nand U3026 (N_3026,N_2602,N_2545);
nor U3027 (N_3027,N_2667,N_2513);
nor U3028 (N_3028,N_2953,N_2954);
or U3029 (N_3029,N_2554,N_2573);
and U3030 (N_3030,N_2523,N_2887);
nor U3031 (N_3031,N_2681,N_2594);
or U3032 (N_3032,N_2966,N_2694);
nand U3033 (N_3033,N_2750,N_2664);
nor U3034 (N_3034,N_2936,N_2637);
or U3035 (N_3035,N_2520,N_2933);
xor U3036 (N_3036,N_2517,N_2579);
nor U3037 (N_3037,N_2532,N_2587);
and U3038 (N_3038,N_2604,N_2987);
nand U3039 (N_3039,N_2880,N_2580);
xor U3040 (N_3040,N_2510,N_2788);
and U3041 (N_3041,N_2623,N_2854);
xnor U3042 (N_3042,N_2603,N_2836);
nor U3043 (N_3043,N_2676,N_2776);
nand U3044 (N_3044,N_2618,N_2556);
xor U3045 (N_3045,N_2826,N_2514);
xor U3046 (N_3046,N_2527,N_2723);
and U3047 (N_3047,N_2871,N_2862);
nand U3048 (N_3048,N_2765,N_2789);
or U3049 (N_3049,N_2975,N_2687);
and U3050 (N_3050,N_2668,N_2802);
nand U3051 (N_3051,N_2629,N_2877);
nor U3052 (N_3052,N_2856,N_2566);
nor U3053 (N_3053,N_2625,N_2639);
or U3054 (N_3054,N_2548,N_2947);
nand U3055 (N_3055,N_2592,N_2829);
xor U3056 (N_3056,N_2972,N_2820);
xor U3057 (N_3057,N_2522,N_2733);
and U3058 (N_3058,N_2622,N_2725);
nor U3059 (N_3059,N_2882,N_2581);
nand U3060 (N_3060,N_2663,N_2958);
and U3061 (N_3061,N_2648,N_2787);
nand U3062 (N_3062,N_2915,N_2772);
nand U3063 (N_3063,N_2985,N_2586);
and U3064 (N_3064,N_2700,N_2549);
nor U3065 (N_3065,N_2988,N_2857);
nor U3066 (N_3066,N_2844,N_2619);
nand U3067 (N_3067,N_2728,N_2657);
or U3068 (N_3068,N_2998,N_2521);
nand U3069 (N_3069,N_2654,N_2539);
and U3070 (N_3070,N_2881,N_2685);
xnor U3071 (N_3071,N_2828,N_2627);
xnor U3072 (N_3072,N_2632,N_2724);
and U3073 (N_3073,N_2559,N_2614);
nand U3074 (N_3074,N_2875,N_2531);
nor U3075 (N_3075,N_2628,N_2842);
nor U3076 (N_3076,N_2994,N_2591);
xnor U3077 (N_3077,N_2868,N_2735);
or U3078 (N_3078,N_2892,N_2683);
or U3079 (N_3079,N_2851,N_2797);
or U3080 (N_3080,N_2680,N_2919);
and U3081 (N_3081,N_2717,N_2589);
nor U3082 (N_3082,N_2533,N_2764);
xnor U3083 (N_3083,N_2605,N_2889);
nor U3084 (N_3084,N_2912,N_2716);
nor U3085 (N_3085,N_2911,N_2525);
and U3086 (N_3086,N_2643,N_2932);
xnor U3087 (N_3087,N_2707,N_2624);
and U3088 (N_3088,N_2609,N_2600);
and U3089 (N_3089,N_2653,N_2801);
nand U3090 (N_3090,N_2908,N_2902);
or U3091 (N_3091,N_2678,N_2597);
or U3092 (N_3092,N_2760,N_2519);
and U3093 (N_3093,N_2669,N_2568);
xnor U3094 (N_3094,N_2869,N_2688);
or U3095 (N_3095,N_2866,N_2661);
xnor U3096 (N_3096,N_2825,N_2544);
or U3097 (N_3097,N_2710,N_2599);
nor U3098 (N_3098,N_2507,N_2691);
nand U3099 (N_3099,N_2732,N_2951);
nand U3100 (N_3100,N_2768,N_2650);
xor U3101 (N_3101,N_2679,N_2598);
and U3102 (N_3102,N_2860,N_2888);
nand U3103 (N_3103,N_2770,N_2719);
nor U3104 (N_3104,N_2744,N_2867);
or U3105 (N_3105,N_2636,N_2935);
xor U3106 (N_3106,N_2779,N_2885);
or U3107 (N_3107,N_2711,N_2886);
nor U3108 (N_3108,N_2563,N_2968);
nor U3109 (N_3109,N_2626,N_2876);
nand U3110 (N_3110,N_2734,N_2675);
xor U3111 (N_3111,N_2928,N_2982);
or U3112 (N_3112,N_2677,N_2923);
and U3113 (N_3113,N_2572,N_2611);
or U3114 (N_3114,N_2553,N_2909);
nand U3115 (N_3115,N_2645,N_2900);
nor U3116 (N_3116,N_2695,N_2655);
and U3117 (N_3117,N_2756,N_2976);
and U3118 (N_3118,N_2833,N_2658);
xor U3119 (N_3119,N_2799,N_2746);
and U3120 (N_3120,N_2979,N_2530);
nand U3121 (N_3121,N_2963,N_2897);
nand U3122 (N_3122,N_2701,N_2937);
and U3123 (N_3123,N_2714,N_2569);
and U3124 (N_3124,N_2830,N_2615);
nor U3125 (N_3125,N_2722,N_2749);
or U3126 (N_3126,N_2890,N_2762);
and U3127 (N_3127,N_2741,N_2763);
xnor U3128 (N_3128,N_2791,N_2916);
nand U3129 (N_3129,N_2872,N_2684);
nand U3130 (N_3130,N_2500,N_2785);
and U3131 (N_3131,N_2904,N_2546);
nand U3132 (N_3132,N_2766,N_2662);
xor U3133 (N_3133,N_2782,N_2552);
xnor U3134 (N_3134,N_2980,N_2927);
or U3135 (N_3135,N_2959,N_2673);
and U3136 (N_3136,N_2752,N_2925);
xnor U3137 (N_3137,N_2995,N_2848);
nand U3138 (N_3138,N_2803,N_2682);
xor U3139 (N_3139,N_2515,N_2738);
nor U3140 (N_3140,N_2646,N_2905);
xor U3141 (N_3141,N_2751,N_2526);
nor U3142 (N_3142,N_2720,N_2564);
xor U3143 (N_3143,N_2565,N_2990);
or U3144 (N_3144,N_2704,N_2703);
and U3145 (N_3145,N_2942,N_2584);
xnor U3146 (N_3146,N_2938,N_2971);
and U3147 (N_3147,N_2705,N_2635);
and U3148 (N_3148,N_2931,N_2859);
xor U3149 (N_3149,N_2640,N_2835);
xnor U3150 (N_3150,N_2815,N_2977);
and U3151 (N_3151,N_2991,N_2805);
xnor U3152 (N_3152,N_2595,N_2907);
and U3153 (N_3153,N_2666,N_2970);
nor U3154 (N_3154,N_2939,N_2913);
or U3155 (N_3155,N_2950,N_2504);
and U3156 (N_3156,N_2656,N_2898);
nor U3157 (N_3157,N_2692,N_2910);
nand U3158 (N_3158,N_2837,N_2613);
nand U3159 (N_3159,N_2808,N_2754);
nor U3160 (N_3160,N_2807,N_2659);
nand U3161 (N_3161,N_2996,N_2903);
or U3162 (N_3162,N_2999,N_2901);
and U3163 (N_3163,N_2630,N_2914);
xor U3164 (N_3164,N_2538,N_2924);
nor U3165 (N_3165,N_2827,N_2800);
nor U3166 (N_3166,N_2612,N_2955);
or U3167 (N_3167,N_2582,N_2721);
or U3168 (N_3168,N_2518,N_2878);
nand U3169 (N_3169,N_2960,N_2847);
nor U3170 (N_3170,N_2562,N_2729);
nor U3171 (N_3171,N_2855,N_2832);
xnor U3172 (N_3172,N_2967,N_2945);
or U3173 (N_3173,N_2849,N_2974);
nand U3174 (N_3174,N_2540,N_2588);
nor U3175 (N_3175,N_2718,N_2879);
nand U3176 (N_3176,N_2537,N_2561);
or U3177 (N_3177,N_2896,N_2555);
or U3178 (N_3178,N_2621,N_2920);
and U3179 (N_3179,N_2696,N_2993);
and U3180 (N_3180,N_2774,N_2505);
xor U3181 (N_3181,N_2686,N_2786);
and U3182 (N_3182,N_2557,N_2997);
nor U3183 (N_3183,N_2783,N_2781);
nor U3184 (N_3184,N_2961,N_2727);
xor U3185 (N_3185,N_2922,N_2906);
xnor U3186 (N_3186,N_2652,N_2690);
nand U3187 (N_3187,N_2894,N_2992);
nor U3188 (N_3188,N_2948,N_2775);
nand U3189 (N_3189,N_2865,N_2610);
or U3190 (N_3190,N_2697,N_2558);
nand U3191 (N_3191,N_2753,N_2755);
nand U3192 (N_3192,N_2593,N_2817);
nand U3193 (N_3193,N_2590,N_2709);
nand U3194 (N_3194,N_2536,N_2585);
nor U3195 (N_3195,N_2651,N_2819);
nand U3196 (N_3196,N_2811,N_2790);
or U3197 (N_3197,N_2693,N_2502);
nor U3198 (N_3198,N_2631,N_2633);
xnor U3199 (N_3199,N_2535,N_2895);
xnor U3200 (N_3200,N_2576,N_2793);
nor U3201 (N_3201,N_2918,N_2780);
nor U3202 (N_3202,N_2670,N_2813);
and U3203 (N_3203,N_2891,N_2617);
or U3204 (N_3204,N_2699,N_2616);
nand U3205 (N_3205,N_2560,N_2665);
or U3206 (N_3206,N_2795,N_2973);
nand U3207 (N_3207,N_2926,N_2822);
xnor U3208 (N_3208,N_2949,N_2863);
or U3209 (N_3209,N_2824,N_2672);
nand U3210 (N_3210,N_2745,N_2759);
and U3211 (N_3211,N_2839,N_2647);
nor U3212 (N_3212,N_2883,N_2606);
nand U3213 (N_3213,N_2934,N_2737);
or U3214 (N_3214,N_2812,N_2981);
nor U3215 (N_3215,N_2984,N_2816);
and U3216 (N_3216,N_2541,N_2706);
nor U3217 (N_3217,N_2534,N_2767);
nand U3218 (N_3218,N_2644,N_2608);
and U3219 (N_3219,N_2712,N_2757);
and U3220 (N_3220,N_2965,N_2846);
nand U3221 (N_3221,N_2571,N_2512);
or U3222 (N_3222,N_2943,N_2634);
nand U3223 (N_3223,N_2834,N_2794);
and U3224 (N_3224,N_2638,N_2550);
nand U3225 (N_3225,N_2858,N_2809);
or U3226 (N_3226,N_2742,N_2524);
xor U3227 (N_3227,N_2574,N_2508);
or U3228 (N_3228,N_2978,N_2739);
nand U3229 (N_3229,N_2940,N_2577);
and U3230 (N_3230,N_2726,N_2743);
nor U3231 (N_3231,N_2509,N_2792);
nor U3232 (N_3232,N_2884,N_2921);
xor U3233 (N_3233,N_2642,N_2983);
xnor U3234 (N_3234,N_2852,N_2596);
nand U3235 (N_3235,N_2796,N_2841);
nand U3236 (N_3236,N_2542,N_2511);
or U3237 (N_3237,N_2964,N_2843);
xnor U3238 (N_3238,N_2516,N_2957);
nor U3239 (N_3239,N_2893,N_2758);
and U3240 (N_3240,N_2850,N_2601);
and U3241 (N_3241,N_2870,N_2798);
and U3242 (N_3242,N_2660,N_2831);
and U3243 (N_3243,N_2814,N_2529);
xor U3244 (N_3244,N_2946,N_2501);
and U3245 (N_3245,N_2702,N_2689);
nor U3246 (N_3246,N_2543,N_2899);
nor U3247 (N_3247,N_2575,N_2674);
xor U3248 (N_3248,N_2778,N_2551);
nand U3249 (N_3249,N_2715,N_2503);
or U3250 (N_3250,N_2700,N_2824);
nor U3251 (N_3251,N_2696,N_2681);
and U3252 (N_3252,N_2930,N_2868);
xnor U3253 (N_3253,N_2596,N_2861);
or U3254 (N_3254,N_2710,N_2950);
or U3255 (N_3255,N_2895,N_2945);
and U3256 (N_3256,N_2676,N_2597);
and U3257 (N_3257,N_2701,N_2517);
nor U3258 (N_3258,N_2907,N_2847);
and U3259 (N_3259,N_2666,N_2776);
or U3260 (N_3260,N_2659,N_2907);
or U3261 (N_3261,N_2691,N_2944);
nand U3262 (N_3262,N_2591,N_2858);
nor U3263 (N_3263,N_2810,N_2598);
and U3264 (N_3264,N_2743,N_2909);
and U3265 (N_3265,N_2662,N_2776);
and U3266 (N_3266,N_2547,N_2989);
xor U3267 (N_3267,N_2684,N_2894);
or U3268 (N_3268,N_2658,N_2775);
and U3269 (N_3269,N_2533,N_2983);
or U3270 (N_3270,N_2763,N_2888);
or U3271 (N_3271,N_2895,N_2741);
xor U3272 (N_3272,N_2649,N_2626);
xor U3273 (N_3273,N_2965,N_2532);
and U3274 (N_3274,N_2604,N_2920);
nor U3275 (N_3275,N_2704,N_2891);
nand U3276 (N_3276,N_2771,N_2833);
or U3277 (N_3277,N_2670,N_2845);
xor U3278 (N_3278,N_2559,N_2612);
or U3279 (N_3279,N_2915,N_2545);
nor U3280 (N_3280,N_2577,N_2808);
nor U3281 (N_3281,N_2863,N_2690);
and U3282 (N_3282,N_2881,N_2709);
and U3283 (N_3283,N_2623,N_2566);
xnor U3284 (N_3284,N_2680,N_2938);
and U3285 (N_3285,N_2927,N_2843);
xnor U3286 (N_3286,N_2939,N_2917);
xnor U3287 (N_3287,N_2539,N_2556);
nor U3288 (N_3288,N_2691,N_2532);
nand U3289 (N_3289,N_2800,N_2644);
nand U3290 (N_3290,N_2646,N_2691);
and U3291 (N_3291,N_2751,N_2534);
and U3292 (N_3292,N_2900,N_2898);
and U3293 (N_3293,N_2869,N_2739);
nand U3294 (N_3294,N_2833,N_2633);
and U3295 (N_3295,N_2784,N_2939);
or U3296 (N_3296,N_2661,N_2942);
and U3297 (N_3297,N_2561,N_2686);
nand U3298 (N_3298,N_2750,N_2660);
and U3299 (N_3299,N_2871,N_2553);
xnor U3300 (N_3300,N_2953,N_2651);
or U3301 (N_3301,N_2719,N_2883);
nor U3302 (N_3302,N_2735,N_2593);
nand U3303 (N_3303,N_2527,N_2894);
and U3304 (N_3304,N_2567,N_2885);
and U3305 (N_3305,N_2503,N_2603);
nor U3306 (N_3306,N_2519,N_2769);
xor U3307 (N_3307,N_2993,N_2799);
nand U3308 (N_3308,N_2525,N_2631);
and U3309 (N_3309,N_2524,N_2623);
xor U3310 (N_3310,N_2943,N_2783);
and U3311 (N_3311,N_2840,N_2740);
xnor U3312 (N_3312,N_2921,N_2889);
xnor U3313 (N_3313,N_2733,N_2600);
xnor U3314 (N_3314,N_2846,N_2906);
xnor U3315 (N_3315,N_2807,N_2702);
nor U3316 (N_3316,N_2544,N_2943);
nor U3317 (N_3317,N_2821,N_2684);
nor U3318 (N_3318,N_2506,N_2939);
nor U3319 (N_3319,N_2820,N_2709);
nand U3320 (N_3320,N_2763,N_2553);
xnor U3321 (N_3321,N_2523,N_2918);
or U3322 (N_3322,N_2641,N_2539);
and U3323 (N_3323,N_2521,N_2979);
and U3324 (N_3324,N_2524,N_2688);
nand U3325 (N_3325,N_2648,N_2506);
and U3326 (N_3326,N_2502,N_2781);
or U3327 (N_3327,N_2979,N_2572);
or U3328 (N_3328,N_2682,N_2977);
xor U3329 (N_3329,N_2684,N_2739);
xnor U3330 (N_3330,N_2896,N_2980);
or U3331 (N_3331,N_2513,N_2891);
xnor U3332 (N_3332,N_2991,N_2855);
nand U3333 (N_3333,N_2729,N_2655);
xor U3334 (N_3334,N_2716,N_2521);
or U3335 (N_3335,N_2683,N_2904);
nand U3336 (N_3336,N_2591,N_2545);
nand U3337 (N_3337,N_2960,N_2826);
nor U3338 (N_3338,N_2966,N_2742);
nor U3339 (N_3339,N_2952,N_2537);
nand U3340 (N_3340,N_2532,N_2958);
and U3341 (N_3341,N_2724,N_2700);
or U3342 (N_3342,N_2798,N_2911);
nand U3343 (N_3343,N_2560,N_2674);
nor U3344 (N_3344,N_2646,N_2864);
xor U3345 (N_3345,N_2845,N_2544);
nand U3346 (N_3346,N_2810,N_2739);
nor U3347 (N_3347,N_2551,N_2992);
and U3348 (N_3348,N_2725,N_2841);
or U3349 (N_3349,N_2979,N_2595);
nor U3350 (N_3350,N_2810,N_2641);
nand U3351 (N_3351,N_2788,N_2500);
nor U3352 (N_3352,N_2978,N_2929);
xnor U3353 (N_3353,N_2975,N_2656);
and U3354 (N_3354,N_2592,N_2645);
nor U3355 (N_3355,N_2779,N_2975);
xnor U3356 (N_3356,N_2561,N_2522);
xnor U3357 (N_3357,N_2541,N_2657);
and U3358 (N_3358,N_2548,N_2788);
and U3359 (N_3359,N_2715,N_2531);
xor U3360 (N_3360,N_2892,N_2617);
or U3361 (N_3361,N_2614,N_2721);
nor U3362 (N_3362,N_2553,N_2560);
xnor U3363 (N_3363,N_2787,N_2586);
nand U3364 (N_3364,N_2835,N_2850);
xor U3365 (N_3365,N_2749,N_2550);
and U3366 (N_3366,N_2551,N_2518);
and U3367 (N_3367,N_2611,N_2786);
and U3368 (N_3368,N_2758,N_2525);
xnor U3369 (N_3369,N_2729,N_2541);
or U3370 (N_3370,N_2568,N_2828);
xnor U3371 (N_3371,N_2534,N_2963);
and U3372 (N_3372,N_2808,N_2832);
and U3373 (N_3373,N_2841,N_2537);
or U3374 (N_3374,N_2771,N_2870);
nor U3375 (N_3375,N_2526,N_2969);
nand U3376 (N_3376,N_2912,N_2931);
nor U3377 (N_3377,N_2720,N_2732);
nand U3378 (N_3378,N_2643,N_2866);
xnor U3379 (N_3379,N_2527,N_2923);
xnor U3380 (N_3380,N_2682,N_2743);
or U3381 (N_3381,N_2719,N_2766);
nor U3382 (N_3382,N_2859,N_2735);
nand U3383 (N_3383,N_2698,N_2572);
nor U3384 (N_3384,N_2999,N_2528);
nor U3385 (N_3385,N_2734,N_2810);
xnor U3386 (N_3386,N_2908,N_2939);
nand U3387 (N_3387,N_2937,N_2939);
nand U3388 (N_3388,N_2689,N_2857);
nor U3389 (N_3389,N_2838,N_2688);
xor U3390 (N_3390,N_2927,N_2502);
xnor U3391 (N_3391,N_2579,N_2823);
nor U3392 (N_3392,N_2584,N_2865);
and U3393 (N_3393,N_2796,N_2925);
xor U3394 (N_3394,N_2518,N_2963);
xor U3395 (N_3395,N_2528,N_2773);
nand U3396 (N_3396,N_2718,N_2830);
and U3397 (N_3397,N_2581,N_2660);
and U3398 (N_3398,N_2953,N_2607);
nand U3399 (N_3399,N_2648,N_2716);
or U3400 (N_3400,N_2984,N_2638);
nand U3401 (N_3401,N_2861,N_2964);
nor U3402 (N_3402,N_2510,N_2938);
and U3403 (N_3403,N_2821,N_2505);
xor U3404 (N_3404,N_2880,N_2609);
or U3405 (N_3405,N_2683,N_2862);
or U3406 (N_3406,N_2963,N_2543);
xnor U3407 (N_3407,N_2723,N_2684);
xnor U3408 (N_3408,N_2797,N_2639);
nand U3409 (N_3409,N_2622,N_2803);
nand U3410 (N_3410,N_2972,N_2529);
and U3411 (N_3411,N_2659,N_2986);
or U3412 (N_3412,N_2904,N_2717);
nand U3413 (N_3413,N_2811,N_2896);
and U3414 (N_3414,N_2622,N_2934);
or U3415 (N_3415,N_2884,N_2827);
xnor U3416 (N_3416,N_2523,N_2592);
nand U3417 (N_3417,N_2747,N_2542);
nand U3418 (N_3418,N_2629,N_2687);
xor U3419 (N_3419,N_2670,N_2962);
nor U3420 (N_3420,N_2506,N_2822);
nand U3421 (N_3421,N_2993,N_2992);
or U3422 (N_3422,N_2823,N_2897);
nor U3423 (N_3423,N_2708,N_2567);
or U3424 (N_3424,N_2739,N_2881);
and U3425 (N_3425,N_2889,N_2538);
nand U3426 (N_3426,N_2913,N_2558);
nor U3427 (N_3427,N_2800,N_2989);
nand U3428 (N_3428,N_2787,N_2568);
xor U3429 (N_3429,N_2805,N_2583);
xnor U3430 (N_3430,N_2514,N_2550);
nand U3431 (N_3431,N_2705,N_2918);
nand U3432 (N_3432,N_2623,N_2659);
xor U3433 (N_3433,N_2622,N_2802);
and U3434 (N_3434,N_2989,N_2825);
nand U3435 (N_3435,N_2743,N_2731);
nor U3436 (N_3436,N_2624,N_2572);
xnor U3437 (N_3437,N_2896,N_2822);
nand U3438 (N_3438,N_2504,N_2773);
and U3439 (N_3439,N_2624,N_2884);
xnor U3440 (N_3440,N_2911,N_2757);
nor U3441 (N_3441,N_2897,N_2625);
nand U3442 (N_3442,N_2808,N_2731);
xor U3443 (N_3443,N_2596,N_2954);
nand U3444 (N_3444,N_2699,N_2565);
and U3445 (N_3445,N_2684,N_2649);
or U3446 (N_3446,N_2501,N_2671);
xnor U3447 (N_3447,N_2881,N_2889);
or U3448 (N_3448,N_2880,N_2753);
nand U3449 (N_3449,N_2793,N_2724);
and U3450 (N_3450,N_2998,N_2511);
xor U3451 (N_3451,N_2679,N_2860);
or U3452 (N_3452,N_2883,N_2859);
nor U3453 (N_3453,N_2817,N_2730);
xor U3454 (N_3454,N_2673,N_2875);
nor U3455 (N_3455,N_2888,N_2962);
nand U3456 (N_3456,N_2689,N_2900);
nor U3457 (N_3457,N_2561,N_2707);
nor U3458 (N_3458,N_2985,N_2506);
xnor U3459 (N_3459,N_2965,N_2646);
nor U3460 (N_3460,N_2885,N_2630);
or U3461 (N_3461,N_2976,N_2828);
and U3462 (N_3462,N_2898,N_2865);
nor U3463 (N_3463,N_2764,N_2921);
nor U3464 (N_3464,N_2591,N_2729);
nand U3465 (N_3465,N_2897,N_2567);
and U3466 (N_3466,N_2655,N_2573);
nor U3467 (N_3467,N_2744,N_2933);
xnor U3468 (N_3468,N_2819,N_2950);
or U3469 (N_3469,N_2533,N_2798);
nor U3470 (N_3470,N_2967,N_2917);
or U3471 (N_3471,N_2509,N_2520);
nand U3472 (N_3472,N_2850,N_2985);
nor U3473 (N_3473,N_2617,N_2850);
or U3474 (N_3474,N_2882,N_2655);
nand U3475 (N_3475,N_2844,N_2705);
or U3476 (N_3476,N_2534,N_2929);
nor U3477 (N_3477,N_2949,N_2648);
nor U3478 (N_3478,N_2905,N_2870);
and U3479 (N_3479,N_2985,N_2519);
xor U3480 (N_3480,N_2519,N_2674);
nand U3481 (N_3481,N_2944,N_2733);
or U3482 (N_3482,N_2654,N_2842);
and U3483 (N_3483,N_2554,N_2546);
and U3484 (N_3484,N_2506,N_2854);
xor U3485 (N_3485,N_2532,N_2898);
nor U3486 (N_3486,N_2775,N_2793);
nand U3487 (N_3487,N_2924,N_2998);
nand U3488 (N_3488,N_2639,N_2887);
nor U3489 (N_3489,N_2565,N_2679);
or U3490 (N_3490,N_2963,N_2736);
or U3491 (N_3491,N_2880,N_2786);
nor U3492 (N_3492,N_2828,N_2842);
and U3493 (N_3493,N_2762,N_2522);
or U3494 (N_3494,N_2986,N_2901);
and U3495 (N_3495,N_2772,N_2943);
or U3496 (N_3496,N_2782,N_2509);
or U3497 (N_3497,N_2700,N_2727);
nand U3498 (N_3498,N_2895,N_2753);
nand U3499 (N_3499,N_2771,N_2737);
or U3500 (N_3500,N_3110,N_3095);
and U3501 (N_3501,N_3055,N_3128);
xnor U3502 (N_3502,N_3438,N_3333);
nor U3503 (N_3503,N_3354,N_3083);
or U3504 (N_3504,N_3497,N_3000);
and U3505 (N_3505,N_3455,N_3239);
or U3506 (N_3506,N_3261,N_3327);
nor U3507 (N_3507,N_3335,N_3402);
and U3508 (N_3508,N_3213,N_3278);
nor U3509 (N_3509,N_3043,N_3324);
and U3510 (N_3510,N_3027,N_3207);
nand U3511 (N_3511,N_3134,N_3181);
xor U3512 (N_3512,N_3193,N_3107);
nand U3513 (N_3513,N_3016,N_3168);
or U3514 (N_3514,N_3205,N_3295);
nand U3515 (N_3515,N_3386,N_3224);
nand U3516 (N_3516,N_3070,N_3190);
or U3517 (N_3517,N_3155,N_3432);
nor U3518 (N_3518,N_3123,N_3150);
nand U3519 (N_3519,N_3434,N_3476);
nand U3520 (N_3520,N_3373,N_3477);
and U3521 (N_3521,N_3360,N_3267);
nor U3522 (N_3522,N_3462,N_3313);
or U3523 (N_3523,N_3217,N_3316);
nor U3524 (N_3524,N_3252,N_3045);
or U3525 (N_3525,N_3347,N_3145);
nand U3526 (N_3526,N_3189,N_3035);
nand U3527 (N_3527,N_3307,N_3254);
xor U3528 (N_3528,N_3240,N_3486);
nand U3529 (N_3529,N_3187,N_3305);
xor U3530 (N_3530,N_3162,N_3409);
nand U3531 (N_3531,N_3484,N_3265);
nor U3532 (N_3532,N_3222,N_3433);
xnor U3533 (N_3533,N_3303,N_3285);
nor U3534 (N_3534,N_3269,N_3118);
or U3535 (N_3535,N_3298,N_3198);
or U3536 (N_3536,N_3358,N_3283);
or U3537 (N_3537,N_3447,N_3268);
and U3538 (N_3538,N_3258,N_3166);
or U3539 (N_3539,N_3159,N_3342);
nor U3540 (N_3540,N_3341,N_3381);
nor U3541 (N_3541,N_3499,N_3359);
xor U3542 (N_3542,N_3385,N_3280);
xnor U3543 (N_3543,N_3022,N_3453);
nand U3544 (N_3544,N_3312,N_3364);
or U3545 (N_3545,N_3304,N_3158);
and U3546 (N_3546,N_3318,N_3214);
nor U3547 (N_3547,N_3445,N_3257);
nor U3548 (N_3548,N_3369,N_3441);
or U3549 (N_3549,N_3101,N_3117);
or U3550 (N_3550,N_3173,N_3363);
or U3551 (N_3551,N_3452,N_3064);
xor U3552 (N_3552,N_3401,N_3093);
or U3553 (N_3553,N_3211,N_3379);
nand U3554 (N_3554,N_3010,N_3351);
or U3555 (N_3555,N_3326,N_3036);
or U3556 (N_3556,N_3308,N_3290);
nor U3557 (N_3557,N_3418,N_3439);
or U3558 (N_3558,N_3137,N_3249);
xor U3559 (N_3559,N_3081,N_3130);
nor U3560 (N_3560,N_3311,N_3400);
nor U3561 (N_3561,N_3136,N_3459);
or U3562 (N_3562,N_3389,N_3460);
and U3563 (N_3563,N_3355,N_3245);
xnor U3564 (N_3564,N_3057,N_3349);
xnor U3565 (N_3565,N_3466,N_3023);
or U3566 (N_3566,N_3328,N_3446);
or U3567 (N_3567,N_3058,N_3156);
or U3568 (N_3568,N_3376,N_3241);
and U3569 (N_3569,N_3197,N_3132);
and U3570 (N_3570,N_3171,N_3006);
or U3571 (N_3571,N_3378,N_3431);
nor U3572 (N_3572,N_3297,N_3282);
nand U3573 (N_3573,N_3203,N_3073);
nor U3574 (N_3574,N_3230,N_3106);
nor U3575 (N_3575,N_3273,N_3002);
nor U3576 (N_3576,N_3019,N_3076);
or U3577 (N_3577,N_3048,N_3480);
nand U3578 (N_3578,N_3122,N_3017);
nand U3579 (N_3579,N_3039,N_3040);
xnor U3580 (N_3580,N_3125,N_3191);
and U3581 (N_3581,N_3068,N_3437);
or U3582 (N_3582,N_3321,N_3296);
or U3583 (N_3583,N_3127,N_3228);
or U3584 (N_3584,N_3302,N_3416);
and U3585 (N_3585,N_3208,N_3247);
and U3586 (N_3586,N_3094,N_3129);
or U3587 (N_3587,N_3229,N_3148);
nand U3588 (N_3588,N_3102,N_3395);
nand U3589 (N_3589,N_3263,N_3215);
nand U3590 (N_3590,N_3352,N_3427);
nand U3591 (N_3591,N_3422,N_3080);
nand U3592 (N_3592,N_3377,N_3075);
or U3593 (N_3593,N_3424,N_3274);
xor U3594 (N_3594,N_3090,N_3147);
xnor U3595 (N_3595,N_3406,N_3233);
nor U3596 (N_3596,N_3049,N_3196);
nand U3597 (N_3597,N_3264,N_3182);
and U3598 (N_3598,N_3192,N_3420);
nand U3599 (N_3599,N_3115,N_3275);
and U3600 (N_3600,N_3103,N_3315);
nor U3601 (N_3601,N_3028,N_3470);
and U3602 (N_3602,N_3001,N_3344);
xor U3603 (N_3603,N_3210,N_3003);
and U3604 (N_3604,N_3170,N_3236);
xnor U3605 (N_3605,N_3113,N_3216);
nand U3606 (N_3606,N_3338,N_3025);
and U3607 (N_3607,N_3448,N_3253);
and U3608 (N_3608,N_3151,N_3119);
and U3609 (N_3609,N_3059,N_3133);
or U3610 (N_3610,N_3111,N_3060);
nand U3611 (N_3611,N_3415,N_3085);
nand U3612 (N_3612,N_3331,N_3371);
nor U3613 (N_3613,N_3412,N_3323);
or U3614 (N_3614,N_3082,N_3436);
or U3615 (N_3615,N_3238,N_3367);
or U3616 (N_3616,N_3219,N_3317);
nor U3617 (N_3617,N_3291,N_3054);
and U3618 (N_3618,N_3366,N_3015);
nand U3619 (N_3619,N_3343,N_3260);
or U3620 (N_3620,N_3186,N_3078);
nor U3621 (N_3621,N_3272,N_3161);
nand U3622 (N_3622,N_3177,N_3287);
nor U3623 (N_3623,N_3013,N_3374);
nand U3624 (N_3624,N_3180,N_3139);
and U3625 (N_3625,N_3276,N_3114);
nand U3626 (N_3626,N_3485,N_3362);
nor U3627 (N_3627,N_3361,N_3306);
nand U3628 (N_3628,N_3489,N_3146);
and U3629 (N_3629,N_3310,N_3353);
nand U3630 (N_3630,N_3467,N_3046);
nor U3631 (N_3631,N_3126,N_3227);
xor U3632 (N_3632,N_3277,N_3174);
or U3633 (N_3633,N_3011,N_3121);
and U3634 (N_3634,N_3077,N_3281);
nor U3635 (N_3635,N_3108,N_3246);
xnor U3636 (N_3636,N_3383,N_3469);
and U3637 (N_3637,N_3243,N_3340);
nor U3638 (N_3638,N_3405,N_3206);
or U3639 (N_3639,N_3397,N_3152);
nor U3640 (N_3640,N_3050,N_3138);
nand U3641 (N_3641,N_3120,N_3100);
nor U3642 (N_3642,N_3200,N_3012);
nor U3643 (N_3643,N_3483,N_3270);
xnor U3644 (N_3644,N_3443,N_3149);
or U3645 (N_3645,N_3185,N_3334);
and U3646 (N_3646,N_3345,N_3284);
or U3647 (N_3647,N_3124,N_3092);
and U3648 (N_3648,N_3346,N_3047);
and U3649 (N_3649,N_3250,N_3116);
and U3650 (N_3650,N_3201,N_3212);
nand U3651 (N_3651,N_3232,N_3348);
nor U3652 (N_3652,N_3375,N_3319);
nand U3653 (N_3653,N_3498,N_3248);
and U3654 (N_3654,N_3104,N_3098);
nand U3655 (N_3655,N_3289,N_3465);
xnor U3656 (N_3656,N_3256,N_3163);
or U3657 (N_3657,N_3225,N_3131);
nor U3658 (N_3658,N_3018,N_3444);
and U3659 (N_3659,N_3069,N_3194);
nand U3660 (N_3660,N_3286,N_3429);
xnor U3661 (N_3661,N_3329,N_3112);
or U3662 (N_3662,N_3365,N_3183);
or U3663 (N_3663,N_3410,N_3195);
and U3664 (N_3664,N_3488,N_3479);
or U3665 (N_3665,N_3178,N_3288);
or U3666 (N_3666,N_3266,N_3086);
xnor U3667 (N_3667,N_3299,N_3255);
xnor U3668 (N_3668,N_3105,N_3387);
or U3669 (N_3669,N_3020,N_3021);
nor U3670 (N_3670,N_3392,N_3079);
xor U3671 (N_3671,N_3417,N_3160);
nand U3672 (N_3672,N_3008,N_3393);
xor U3673 (N_3673,N_3141,N_3388);
and U3674 (N_3674,N_3394,N_3458);
xnor U3675 (N_3675,N_3271,N_3144);
nor U3676 (N_3676,N_3457,N_3014);
or U3677 (N_3677,N_3164,N_3034);
and U3678 (N_3678,N_3165,N_3033);
or U3679 (N_3679,N_3005,N_3099);
nor U3680 (N_3680,N_3423,N_3184);
and U3681 (N_3681,N_3172,N_3450);
or U3682 (N_3682,N_3259,N_3398);
nand U3683 (N_3683,N_3157,N_3053);
nand U3684 (N_3684,N_3314,N_3024);
xnor U3685 (N_3685,N_3067,N_3234);
nor U3686 (N_3686,N_3370,N_3066);
or U3687 (N_3687,N_3380,N_3482);
nor U3688 (N_3688,N_3411,N_3390);
and U3689 (N_3689,N_3451,N_3474);
nand U3690 (N_3690,N_3044,N_3071);
xnor U3691 (N_3691,N_3204,N_3065);
or U3692 (N_3692,N_3494,N_3218);
or U3693 (N_3693,N_3478,N_3062);
xnor U3694 (N_3694,N_3292,N_3475);
xor U3695 (N_3695,N_3235,N_3339);
and U3696 (N_3696,N_3325,N_3421);
nand U3697 (N_3697,N_3169,N_3029);
nor U3698 (N_3698,N_3142,N_3337);
xnor U3699 (N_3699,N_3493,N_3300);
or U3700 (N_3700,N_3336,N_3413);
xnor U3701 (N_3701,N_3089,N_3087);
or U3702 (N_3702,N_3440,N_3179);
nor U3703 (N_3703,N_3220,N_3430);
or U3704 (N_3704,N_3221,N_3188);
nand U3705 (N_3705,N_3384,N_3030);
or U3706 (N_3706,N_3391,N_3251);
nand U3707 (N_3707,N_3135,N_3332);
or U3708 (N_3708,N_3403,N_3056);
xnor U3709 (N_3709,N_3231,N_3419);
and U3710 (N_3710,N_3209,N_3320);
nand U3711 (N_3711,N_3396,N_3454);
nor U3712 (N_3712,N_3140,N_3496);
and U3713 (N_3713,N_3242,N_3154);
xor U3714 (N_3714,N_3244,N_3202);
xnor U3715 (N_3715,N_3472,N_3226);
nand U3716 (N_3716,N_3051,N_3372);
xor U3717 (N_3717,N_3279,N_3031);
or U3718 (N_3718,N_3097,N_3153);
nand U3719 (N_3719,N_3009,N_3426);
nand U3720 (N_3720,N_3032,N_3425);
and U3721 (N_3721,N_3461,N_3088);
xnor U3722 (N_3722,N_3143,N_3492);
xnor U3723 (N_3723,N_3301,N_3468);
xor U3724 (N_3724,N_3495,N_3223);
and U3725 (N_3725,N_3042,N_3463);
xnor U3726 (N_3726,N_3061,N_3330);
or U3727 (N_3727,N_3491,N_3490);
or U3728 (N_3728,N_3435,N_3038);
or U3729 (N_3729,N_3404,N_3072);
nor U3730 (N_3730,N_3473,N_3464);
or U3731 (N_3731,N_3176,N_3408);
nor U3732 (N_3732,N_3442,N_3399);
and U3733 (N_3733,N_3471,N_3026);
nand U3734 (N_3734,N_3294,N_3041);
or U3735 (N_3735,N_3199,N_3428);
nand U3736 (N_3736,N_3109,N_3091);
nor U3737 (N_3737,N_3167,N_3357);
nand U3738 (N_3738,N_3481,N_3368);
xnor U3739 (N_3739,N_3309,N_3074);
or U3740 (N_3740,N_3293,N_3414);
nor U3741 (N_3741,N_3356,N_3007);
nor U3742 (N_3742,N_3262,N_3487);
or U3743 (N_3743,N_3456,N_3237);
and U3744 (N_3744,N_3382,N_3052);
nand U3745 (N_3745,N_3449,N_3084);
nor U3746 (N_3746,N_3037,N_3004);
nor U3747 (N_3747,N_3096,N_3175);
xor U3748 (N_3748,N_3407,N_3350);
nor U3749 (N_3749,N_3322,N_3063);
nand U3750 (N_3750,N_3424,N_3448);
and U3751 (N_3751,N_3246,N_3380);
nor U3752 (N_3752,N_3401,N_3363);
nor U3753 (N_3753,N_3035,N_3407);
xor U3754 (N_3754,N_3124,N_3326);
or U3755 (N_3755,N_3471,N_3432);
xor U3756 (N_3756,N_3432,N_3182);
nand U3757 (N_3757,N_3141,N_3344);
xnor U3758 (N_3758,N_3481,N_3371);
nand U3759 (N_3759,N_3018,N_3100);
xor U3760 (N_3760,N_3370,N_3362);
nor U3761 (N_3761,N_3456,N_3169);
or U3762 (N_3762,N_3274,N_3209);
and U3763 (N_3763,N_3350,N_3075);
and U3764 (N_3764,N_3253,N_3005);
xnor U3765 (N_3765,N_3135,N_3403);
xnor U3766 (N_3766,N_3014,N_3003);
nor U3767 (N_3767,N_3483,N_3420);
nor U3768 (N_3768,N_3260,N_3436);
or U3769 (N_3769,N_3180,N_3319);
xor U3770 (N_3770,N_3312,N_3151);
xnor U3771 (N_3771,N_3211,N_3261);
xor U3772 (N_3772,N_3335,N_3417);
and U3773 (N_3773,N_3083,N_3473);
xnor U3774 (N_3774,N_3163,N_3343);
and U3775 (N_3775,N_3232,N_3188);
nand U3776 (N_3776,N_3356,N_3467);
and U3777 (N_3777,N_3449,N_3310);
and U3778 (N_3778,N_3004,N_3132);
xnor U3779 (N_3779,N_3030,N_3258);
xor U3780 (N_3780,N_3037,N_3343);
or U3781 (N_3781,N_3290,N_3080);
xor U3782 (N_3782,N_3174,N_3168);
nand U3783 (N_3783,N_3306,N_3468);
nor U3784 (N_3784,N_3316,N_3337);
or U3785 (N_3785,N_3256,N_3399);
xnor U3786 (N_3786,N_3233,N_3439);
xnor U3787 (N_3787,N_3055,N_3019);
or U3788 (N_3788,N_3392,N_3223);
and U3789 (N_3789,N_3384,N_3150);
nand U3790 (N_3790,N_3186,N_3264);
nor U3791 (N_3791,N_3129,N_3309);
and U3792 (N_3792,N_3005,N_3495);
xor U3793 (N_3793,N_3178,N_3113);
nand U3794 (N_3794,N_3056,N_3043);
or U3795 (N_3795,N_3048,N_3025);
and U3796 (N_3796,N_3327,N_3392);
or U3797 (N_3797,N_3297,N_3215);
and U3798 (N_3798,N_3119,N_3115);
or U3799 (N_3799,N_3378,N_3413);
and U3800 (N_3800,N_3053,N_3236);
and U3801 (N_3801,N_3493,N_3374);
and U3802 (N_3802,N_3447,N_3454);
nand U3803 (N_3803,N_3046,N_3383);
or U3804 (N_3804,N_3036,N_3432);
nor U3805 (N_3805,N_3266,N_3322);
or U3806 (N_3806,N_3025,N_3090);
or U3807 (N_3807,N_3296,N_3315);
xor U3808 (N_3808,N_3272,N_3189);
xor U3809 (N_3809,N_3405,N_3435);
nor U3810 (N_3810,N_3342,N_3219);
and U3811 (N_3811,N_3489,N_3132);
nand U3812 (N_3812,N_3216,N_3394);
or U3813 (N_3813,N_3488,N_3126);
or U3814 (N_3814,N_3280,N_3347);
nor U3815 (N_3815,N_3122,N_3407);
or U3816 (N_3816,N_3386,N_3080);
nor U3817 (N_3817,N_3028,N_3359);
and U3818 (N_3818,N_3413,N_3174);
xor U3819 (N_3819,N_3212,N_3451);
and U3820 (N_3820,N_3479,N_3328);
nand U3821 (N_3821,N_3061,N_3354);
and U3822 (N_3822,N_3075,N_3161);
or U3823 (N_3823,N_3465,N_3121);
nand U3824 (N_3824,N_3443,N_3132);
nand U3825 (N_3825,N_3099,N_3439);
nand U3826 (N_3826,N_3191,N_3105);
xnor U3827 (N_3827,N_3279,N_3222);
or U3828 (N_3828,N_3258,N_3403);
nand U3829 (N_3829,N_3365,N_3405);
or U3830 (N_3830,N_3488,N_3296);
nor U3831 (N_3831,N_3167,N_3052);
nor U3832 (N_3832,N_3380,N_3403);
nand U3833 (N_3833,N_3044,N_3025);
or U3834 (N_3834,N_3390,N_3285);
or U3835 (N_3835,N_3455,N_3225);
and U3836 (N_3836,N_3195,N_3015);
or U3837 (N_3837,N_3319,N_3403);
or U3838 (N_3838,N_3321,N_3127);
nor U3839 (N_3839,N_3493,N_3157);
nand U3840 (N_3840,N_3043,N_3090);
nor U3841 (N_3841,N_3040,N_3131);
and U3842 (N_3842,N_3201,N_3461);
nand U3843 (N_3843,N_3314,N_3393);
and U3844 (N_3844,N_3364,N_3321);
and U3845 (N_3845,N_3385,N_3491);
and U3846 (N_3846,N_3034,N_3301);
xnor U3847 (N_3847,N_3090,N_3470);
nor U3848 (N_3848,N_3251,N_3029);
nor U3849 (N_3849,N_3187,N_3061);
xnor U3850 (N_3850,N_3083,N_3058);
or U3851 (N_3851,N_3181,N_3313);
and U3852 (N_3852,N_3177,N_3144);
xnor U3853 (N_3853,N_3173,N_3401);
or U3854 (N_3854,N_3319,N_3006);
and U3855 (N_3855,N_3078,N_3165);
and U3856 (N_3856,N_3471,N_3376);
nand U3857 (N_3857,N_3221,N_3019);
xor U3858 (N_3858,N_3328,N_3167);
and U3859 (N_3859,N_3457,N_3187);
nand U3860 (N_3860,N_3388,N_3313);
xor U3861 (N_3861,N_3211,N_3127);
xnor U3862 (N_3862,N_3468,N_3081);
xnor U3863 (N_3863,N_3003,N_3218);
nor U3864 (N_3864,N_3384,N_3052);
nor U3865 (N_3865,N_3256,N_3288);
nor U3866 (N_3866,N_3269,N_3492);
nand U3867 (N_3867,N_3040,N_3228);
nor U3868 (N_3868,N_3302,N_3448);
nor U3869 (N_3869,N_3171,N_3323);
and U3870 (N_3870,N_3081,N_3209);
xor U3871 (N_3871,N_3347,N_3217);
and U3872 (N_3872,N_3477,N_3491);
nand U3873 (N_3873,N_3058,N_3179);
nand U3874 (N_3874,N_3059,N_3496);
and U3875 (N_3875,N_3281,N_3434);
and U3876 (N_3876,N_3030,N_3461);
xnor U3877 (N_3877,N_3304,N_3430);
or U3878 (N_3878,N_3289,N_3257);
xor U3879 (N_3879,N_3300,N_3077);
nor U3880 (N_3880,N_3136,N_3313);
nand U3881 (N_3881,N_3360,N_3497);
or U3882 (N_3882,N_3075,N_3276);
xor U3883 (N_3883,N_3071,N_3256);
nand U3884 (N_3884,N_3113,N_3339);
and U3885 (N_3885,N_3444,N_3187);
nor U3886 (N_3886,N_3382,N_3325);
and U3887 (N_3887,N_3478,N_3101);
nand U3888 (N_3888,N_3307,N_3455);
and U3889 (N_3889,N_3411,N_3493);
xnor U3890 (N_3890,N_3408,N_3247);
nand U3891 (N_3891,N_3068,N_3177);
xnor U3892 (N_3892,N_3295,N_3196);
nor U3893 (N_3893,N_3317,N_3257);
nor U3894 (N_3894,N_3014,N_3440);
nor U3895 (N_3895,N_3430,N_3104);
or U3896 (N_3896,N_3428,N_3406);
nand U3897 (N_3897,N_3116,N_3308);
and U3898 (N_3898,N_3096,N_3282);
xor U3899 (N_3899,N_3269,N_3027);
nand U3900 (N_3900,N_3046,N_3010);
xor U3901 (N_3901,N_3218,N_3236);
or U3902 (N_3902,N_3218,N_3495);
nor U3903 (N_3903,N_3150,N_3430);
or U3904 (N_3904,N_3104,N_3067);
and U3905 (N_3905,N_3084,N_3448);
nand U3906 (N_3906,N_3348,N_3337);
nor U3907 (N_3907,N_3232,N_3000);
and U3908 (N_3908,N_3131,N_3401);
and U3909 (N_3909,N_3441,N_3077);
nand U3910 (N_3910,N_3291,N_3131);
and U3911 (N_3911,N_3064,N_3031);
nand U3912 (N_3912,N_3306,N_3144);
nor U3913 (N_3913,N_3177,N_3002);
nor U3914 (N_3914,N_3035,N_3140);
and U3915 (N_3915,N_3008,N_3321);
or U3916 (N_3916,N_3061,N_3480);
and U3917 (N_3917,N_3289,N_3040);
or U3918 (N_3918,N_3285,N_3154);
xnor U3919 (N_3919,N_3166,N_3172);
nand U3920 (N_3920,N_3039,N_3181);
xor U3921 (N_3921,N_3460,N_3258);
and U3922 (N_3922,N_3173,N_3043);
or U3923 (N_3923,N_3163,N_3038);
and U3924 (N_3924,N_3392,N_3250);
nor U3925 (N_3925,N_3217,N_3324);
xor U3926 (N_3926,N_3091,N_3182);
xor U3927 (N_3927,N_3283,N_3016);
xnor U3928 (N_3928,N_3315,N_3194);
nor U3929 (N_3929,N_3012,N_3216);
or U3930 (N_3930,N_3200,N_3250);
nand U3931 (N_3931,N_3449,N_3482);
nand U3932 (N_3932,N_3001,N_3483);
and U3933 (N_3933,N_3295,N_3280);
nand U3934 (N_3934,N_3191,N_3453);
nor U3935 (N_3935,N_3337,N_3242);
and U3936 (N_3936,N_3267,N_3078);
nor U3937 (N_3937,N_3450,N_3373);
and U3938 (N_3938,N_3256,N_3459);
xnor U3939 (N_3939,N_3140,N_3442);
nand U3940 (N_3940,N_3407,N_3255);
xnor U3941 (N_3941,N_3421,N_3007);
nor U3942 (N_3942,N_3173,N_3309);
nand U3943 (N_3943,N_3225,N_3083);
nand U3944 (N_3944,N_3026,N_3029);
nand U3945 (N_3945,N_3413,N_3326);
xor U3946 (N_3946,N_3053,N_3188);
xor U3947 (N_3947,N_3097,N_3499);
xor U3948 (N_3948,N_3319,N_3135);
or U3949 (N_3949,N_3105,N_3383);
nand U3950 (N_3950,N_3318,N_3390);
nand U3951 (N_3951,N_3312,N_3249);
nand U3952 (N_3952,N_3117,N_3222);
nor U3953 (N_3953,N_3052,N_3415);
or U3954 (N_3954,N_3164,N_3454);
xor U3955 (N_3955,N_3137,N_3100);
or U3956 (N_3956,N_3429,N_3049);
or U3957 (N_3957,N_3144,N_3278);
xnor U3958 (N_3958,N_3104,N_3020);
xnor U3959 (N_3959,N_3054,N_3470);
or U3960 (N_3960,N_3423,N_3471);
nor U3961 (N_3961,N_3034,N_3190);
nor U3962 (N_3962,N_3300,N_3388);
xnor U3963 (N_3963,N_3496,N_3145);
and U3964 (N_3964,N_3445,N_3047);
nand U3965 (N_3965,N_3239,N_3304);
or U3966 (N_3966,N_3159,N_3141);
or U3967 (N_3967,N_3047,N_3419);
and U3968 (N_3968,N_3496,N_3309);
nand U3969 (N_3969,N_3304,N_3485);
xor U3970 (N_3970,N_3314,N_3427);
or U3971 (N_3971,N_3264,N_3283);
or U3972 (N_3972,N_3265,N_3146);
or U3973 (N_3973,N_3029,N_3128);
nor U3974 (N_3974,N_3302,N_3420);
nor U3975 (N_3975,N_3459,N_3458);
nor U3976 (N_3976,N_3317,N_3292);
nand U3977 (N_3977,N_3436,N_3496);
nor U3978 (N_3978,N_3374,N_3154);
nor U3979 (N_3979,N_3238,N_3437);
or U3980 (N_3980,N_3317,N_3223);
nor U3981 (N_3981,N_3257,N_3488);
nor U3982 (N_3982,N_3274,N_3004);
nand U3983 (N_3983,N_3374,N_3036);
xnor U3984 (N_3984,N_3472,N_3320);
nor U3985 (N_3985,N_3327,N_3088);
nor U3986 (N_3986,N_3028,N_3291);
xnor U3987 (N_3987,N_3435,N_3385);
nor U3988 (N_3988,N_3318,N_3014);
and U3989 (N_3989,N_3160,N_3297);
or U3990 (N_3990,N_3080,N_3423);
or U3991 (N_3991,N_3296,N_3308);
nand U3992 (N_3992,N_3292,N_3375);
or U3993 (N_3993,N_3407,N_3271);
and U3994 (N_3994,N_3117,N_3160);
nor U3995 (N_3995,N_3280,N_3351);
xnor U3996 (N_3996,N_3172,N_3384);
xor U3997 (N_3997,N_3062,N_3488);
and U3998 (N_3998,N_3115,N_3194);
or U3999 (N_3999,N_3371,N_3394);
or U4000 (N_4000,N_3570,N_3531);
nand U4001 (N_4001,N_3734,N_3840);
xor U4002 (N_4002,N_3832,N_3998);
and U4003 (N_4003,N_3640,N_3748);
or U4004 (N_4004,N_3954,N_3710);
and U4005 (N_4005,N_3899,N_3881);
nor U4006 (N_4006,N_3850,N_3908);
and U4007 (N_4007,N_3993,N_3631);
nor U4008 (N_4008,N_3842,N_3544);
nor U4009 (N_4009,N_3501,N_3791);
and U4010 (N_4010,N_3648,N_3591);
xor U4011 (N_4011,N_3976,N_3938);
nor U4012 (N_4012,N_3510,N_3575);
xor U4013 (N_4013,N_3893,N_3636);
nor U4014 (N_4014,N_3922,N_3981);
and U4015 (N_4015,N_3848,N_3685);
nand U4016 (N_4016,N_3637,N_3997);
nor U4017 (N_4017,N_3694,N_3578);
or U4018 (N_4018,N_3798,N_3617);
or U4019 (N_4019,N_3776,N_3619);
and U4020 (N_4020,N_3825,N_3777);
and U4021 (N_4021,N_3602,N_3500);
nand U4022 (N_4022,N_3901,N_3810);
nand U4023 (N_4023,N_3876,N_3698);
xor U4024 (N_4024,N_3562,N_3768);
or U4025 (N_4025,N_3638,N_3749);
nor U4026 (N_4026,N_3868,N_3610);
nor U4027 (N_4027,N_3650,N_3763);
and U4028 (N_4028,N_3944,N_3984);
xor U4029 (N_4029,N_3590,N_3793);
xor U4030 (N_4030,N_3764,N_3985);
xor U4031 (N_4031,N_3601,N_3503);
nand U4032 (N_4032,N_3577,N_3589);
and U4033 (N_4033,N_3582,N_3936);
or U4034 (N_4034,N_3773,N_3704);
xor U4035 (N_4035,N_3753,N_3872);
nor U4036 (N_4036,N_3940,N_3626);
or U4037 (N_4037,N_3526,N_3863);
nand U4038 (N_4038,N_3635,N_3731);
nor U4039 (N_4039,N_3913,N_3581);
nand U4040 (N_4040,N_3599,N_3992);
xnor U4041 (N_4041,N_3966,N_3683);
or U4042 (N_4042,N_3870,N_3645);
xnor U4043 (N_4043,N_3717,N_3835);
or U4044 (N_4044,N_3625,N_3929);
nand U4045 (N_4045,N_3928,N_3541);
nor U4046 (N_4046,N_3950,N_3979);
and U4047 (N_4047,N_3968,N_3829);
or U4048 (N_4048,N_3911,N_3546);
or U4049 (N_4049,N_3925,N_3812);
nand U4050 (N_4050,N_3836,N_3527);
xor U4051 (N_4051,N_3666,N_3797);
and U4052 (N_4052,N_3540,N_3779);
and U4053 (N_4053,N_3695,N_3831);
xor U4054 (N_4054,N_3909,N_3604);
xor U4055 (N_4055,N_3709,N_3658);
and U4056 (N_4056,N_3708,N_3897);
nand U4057 (N_4057,N_3550,N_3691);
xnor U4058 (N_4058,N_3719,N_3743);
and U4059 (N_4059,N_3644,N_3706);
xnor U4060 (N_4060,N_3888,N_3623);
xor U4061 (N_4061,N_3711,N_3547);
nor U4062 (N_4062,N_3978,N_3530);
xor U4063 (N_4063,N_3697,N_3517);
and U4064 (N_4064,N_3600,N_3630);
nor U4065 (N_4065,N_3785,N_3947);
or U4066 (N_4066,N_3543,N_3745);
and U4067 (N_4067,N_3766,N_3952);
and U4068 (N_4068,N_3960,N_3827);
xnor U4069 (N_4069,N_3584,N_3632);
xor U4070 (N_4070,N_3548,N_3505);
xnor U4071 (N_4071,N_3539,N_3613);
nand U4072 (N_4072,N_3535,N_3524);
nor U4073 (N_4073,N_3620,N_3756);
nand U4074 (N_4074,N_3730,N_3882);
nand U4075 (N_4075,N_3678,N_3885);
xor U4076 (N_4076,N_3627,N_3890);
or U4077 (N_4077,N_3747,N_3813);
and U4078 (N_4078,N_3659,N_3877);
xor U4079 (N_4079,N_3516,N_3560);
nand U4080 (N_4080,N_3639,N_3845);
xor U4081 (N_4081,N_3927,N_3563);
nand U4082 (N_4082,N_3667,N_3671);
or U4083 (N_4083,N_3824,N_3867);
or U4084 (N_4084,N_3515,N_3712);
and U4085 (N_4085,N_3843,N_3826);
or U4086 (N_4086,N_3880,N_3705);
nor U4087 (N_4087,N_3849,N_3995);
xnor U4088 (N_4088,N_3693,N_3977);
nor U4089 (N_4089,N_3994,N_3741);
nor U4090 (N_4090,N_3969,N_3643);
nor U4091 (N_4091,N_3742,N_3512);
or U4092 (N_4092,N_3957,N_3651);
nor U4093 (N_4093,N_3844,N_3528);
or U4094 (N_4094,N_3941,N_3989);
or U4095 (N_4095,N_3809,N_3507);
xor U4096 (N_4096,N_3884,N_3751);
and U4097 (N_4097,N_3733,N_3783);
or U4098 (N_4098,N_3805,N_3525);
xor U4099 (N_4099,N_3815,N_3769);
and U4100 (N_4100,N_3830,N_3687);
and U4101 (N_4101,N_3971,N_3921);
nand U4102 (N_4102,N_3724,N_3784);
or U4103 (N_4103,N_3789,N_3757);
nand U4104 (N_4104,N_3714,N_3518);
and U4105 (N_4105,N_3738,N_3537);
nor U4106 (N_4106,N_3961,N_3934);
nand U4107 (N_4107,N_3973,N_3910);
and U4108 (N_4108,N_3556,N_3871);
and U4109 (N_4109,N_3838,N_3655);
xnor U4110 (N_4110,N_3847,N_3780);
nor U4111 (N_4111,N_3545,N_3522);
xor U4112 (N_4112,N_3588,N_3737);
or U4113 (N_4113,N_3608,N_3624);
and U4114 (N_4114,N_3752,N_3728);
and U4115 (N_4115,N_3772,N_3834);
nand U4116 (N_4116,N_3787,N_3502);
nand U4117 (N_4117,N_3820,N_3605);
or U4118 (N_4118,N_3725,N_3907);
nor U4119 (N_4119,N_3926,N_3726);
xor U4120 (N_4120,N_3949,N_3837);
or U4121 (N_4121,N_3958,N_3696);
xor U4122 (N_4122,N_3965,N_3740);
nand U4123 (N_4123,N_3767,N_3814);
xor U4124 (N_4124,N_3661,N_3504);
xnor U4125 (N_4125,N_3657,N_3816);
and U4126 (N_4126,N_3664,N_3951);
or U4127 (N_4127,N_3953,N_3569);
nor U4128 (N_4128,N_3754,N_3675);
xnor U4129 (N_4129,N_3758,N_3692);
xnor U4130 (N_4130,N_3795,N_3796);
or U4131 (N_4131,N_3653,N_3823);
or U4132 (N_4132,N_3746,N_3663);
and U4133 (N_4133,N_3778,N_3962);
xor U4134 (N_4134,N_3920,N_3860);
nor U4135 (N_4135,N_3916,N_3794);
nor U4136 (N_4136,N_3828,N_3851);
nor U4137 (N_4137,N_3946,N_3833);
nor U4138 (N_4138,N_3647,N_3665);
xor U4139 (N_4139,N_3856,N_3558);
or U4140 (N_4140,N_3662,N_3593);
xnor U4141 (N_4141,N_3883,N_3603);
nor U4142 (N_4142,N_3686,N_3846);
nand U4143 (N_4143,N_3607,N_3732);
or U4144 (N_4144,N_3554,N_3821);
or U4145 (N_4145,N_3807,N_3853);
or U4146 (N_4146,N_3879,N_3980);
xnor U4147 (N_4147,N_3576,N_3932);
nor U4148 (N_4148,N_3990,N_3839);
nor U4149 (N_4149,N_3739,N_3891);
or U4150 (N_4150,N_3878,N_3781);
and U4151 (N_4151,N_3771,N_3786);
and U4152 (N_4152,N_3873,N_3761);
nor U4153 (N_4153,N_3895,N_3713);
xor U4154 (N_4154,N_3621,N_3765);
nand U4155 (N_4155,N_3750,N_3649);
or U4156 (N_4156,N_3963,N_3534);
xnor U4157 (N_4157,N_3629,N_3808);
and U4158 (N_4158,N_3520,N_3991);
xnor U4159 (N_4159,N_3536,N_3803);
and U4160 (N_4160,N_3887,N_3633);
nor U4161 (N_4161,N_3718,N_3673);
and U4162 (N_4162,N_3583,N_3755);
and U4163 (N_4163,N_3677,N_3970);
nand U4164 (N_4164,N_3668,N_3646);
xor U4165 (N_4165,N_3587,N_3854);
xnor U4166 (N_4166,N_3679,N_3506);
nor U4167 (N_4167,N_3735,N_3565);
nor U4168 (N_4168,N_3948,N_3799);
and U4169 (N_4169,N_3945,N_3841);
xor U4170 (N_4170,N_3906,N_3521);
xnor U4171 (N_4171,N_3792,N_3919);
xnor U4172 (N_4172,N_3615,N_3902);
nor U4173 (N_4173,N_3669,N_3811);
nand U4174 (N_4174,N_3744,N_3964);
nand U4175 (N_4175,N_3672,N_3555);
xnor U4176 (N_4176,N_3802,N_3759);
nor U4177 (N_4177,N_3788,N_3579);
nor U4178 (N_4178,N_3592,N_3903);
nor U4179 (N_4179,N_3727,N_3523);
nand U4180 (N_4180,N_3701,N_3889);
xnor U4181 (N_4181,N_3762,N_3806);
and U4182 (N_4182,N_3865,N_3596);
or U4183 (N_4183,N_3652,N_3818);
and U4184 (N_4184,N_3720,N_3931);
nor U4185 (N_4185,N_3999,N_3801);
xor U4186 (N_4186,N_3656,N_3559);
or U4187 (N_4187,N_3959,N_3574);
nand U4188 (N_4188,N_3972,N_3606);
nand U4189 (N_4189,N_3939,N_3680);
nand U4190 (N_4190,N_3896,N_3866);
xnor U4191 (N_4191,N_3716,N_3861);
nor U4192 (N_4192,N_3551,N_3622);
or U4193 (N_4193,N_3508,N_3612);
nor U4194 (N_4194,N_3942,N_3943);
nand U4195 (N_4195,N_3690,N_3611);
and U4196 (N_4196,N_3996,N_3855);
xnor U4197 (N_4197,N_3519,N_3886);
xnor U4198 (N_4198,N_3987,N_3923);
nand U4199 (N_4199,N_3864,N_3595);
xnor U4200 (N_4200,N_3736,N_3513);
nor U4201 (N_4201,N_3819,N_3975);
nand U4202 (N_4202,N_3924,N_3580);
xor U4203 (N_4203,N_3557,N_3509);
and U4204 (N_4204,N_3723,N_3874);
nor U4205 (N_4205,N_3988,N_3585);
and U4206 (N_4206,N_3641,N_3770);
nor U4207 (N_4207,N_3715,N_3986);
nand U4208 (N_4208,N_3782,N_3571);
nor U4209 (N_4209,N_3628,N_3682);
nand U4210 (N_4210,N_3933,N_3775);
and U4211 (N_4211,N_3642,N_3822);
or U4212 (N_4212,N_3894,N_3654);
nor U4213 (N_4213,N_3956,N_3618);
nor U4214 (N_4214,N_3549,N_3586);
nand U4215 (N_4215,N_3597,N_3561);
and U4216 (N_4216,N_3905,N_3538);
nand U4217 (N_4217,N_3688,N_3699);
and U4218 (N_4218,N_3915,N_3983);
xor U4219 (N_4219,N_3703,N_3729);
nor U4220 (N_4220,N_3898,N_3598);
xnor U4221 (N_4221,N_3670,N_3935);
nor U4222 (N_4222,N_3532,N_3674);
nand U4223 (N_4223,N_3566,N_3676);
nor U4224 (N_4224,N_3760,N_3702);
and U4225 (N_4225,N_3552,N_3616);
nand U4226 (N_4226,N_3721,N_3857);
xnor U4227 (N_4227,N_3914,N_3930);
nand U4228 (N_4228,N_3858,N_3573);
nor U4229 (N_4229,N_3790,N_3917);
and U4230 (N_4230,N_3681,N_3817);
or U4231 (N_4231,N_3904,N_3700);
xor U4232 (N_4232,N_3852,N_3774);
xnor U4233 (N_4233,N_3609,N_3511);
nand U4234 (N_4234,N_3660,N_3564);
xnor U4235 (N_4235,N_3875,N_3862);
nand U4236 (N_4236,N_3684,N_3614);
or U4237 (N_4237,N_3568,N_3937);
xor U4238 (N_4238,N_3974,N_3955);
xnor U4239 (N_4239,N_3967,N_3918);
nand U4240 (N_4240,N_3634,N_3567);
nand U4241 (N_4241,N_3514,N_3707);
nor U4242 (N_4242,N_3804,N_3594);
and U4243 (N_4243,N_3800,N_3553);
and U4244 (N_4244,N_3912,N_3722);
and U4245 (N_4245,N_3859,N_3572);
nand U4246 (N_4246,N_3689,N_3900);
and U4247 (N_4247,N_3982,N_3869);
nand U4248 (N_4248,N_3892,N_3529);
nor U4249 (N_4249,N_3533,N_3542);
nor U4250 (N_4250,N_3818,N_3837);
nor U4251 (N_4251,N_3767,N_3857);
and U4252 (N_4252,N_3704,N_3517);
and U4253 (N_4253,N_3500,N_3568);
or U4254 (N_4254,N_3752,N_3566);
nand U4255 (N_4255,N_3722,N_3595);
nand U4256 (N_4256,N_3532,N_3852);
and U4257 (N_4257,N_3644,N_3586);
nand U4258 (N_4258,N_3951,N_3793);
or U4259 (N_4259,N_3913,N_3853);
nor U4260 (N_4260,N_3994,N_3963);
or U4261 (N_4261,N_3656,N_3899);
or U4262 (N_4262,N_3968,N_3999);
nand U4263 (N_4263,N_3909,N_3513);
nand U4264 (N_4264,N_3529,N_3800);
or U4265 (N_4265,N_3687,N_3986);
and U4266 (N_4266,N_3641,N_3831);
xnor U4267 (N_4267,N_3765,N_3900);
xnor U4268 (N_4268,N_3833,N_3935);
xnor U4269 (N_4269,N_3823,N_3758);
xor U4270 (N_4270,N_3823,N_3660);
and U4271 (N_4271,N_3770,N_3795);
nand U4272 (N_4272,N_3696,N_3540);
nand U4273 (N_4273,N_3989,N_3708);
nand U4274 (N_4274,N_3779,N_3865);
or U4275 (N_4275,N_3918,N_3715);
xor U4276 (N_4276,N_3540,N_3888);
or U4277 (N_4277,N_3616,N_3579);
nor U4278 (N_4278,N_3704,N_3600);
nor U4279 (N_4279,N_3631,N_3511);
xnor U4280 (N_4280,N_3900,N_3729);
or U4281 (N_4281,N_3695,N_3552);
or U4282 (N_4282,N_3854,N_3668);
nand U4283 (N_4283,N_3682,N_3942);
and U4284 (N_4284,N_3509,N_3870);
xor U4285 (N_4285,N_3756,N_3568);
nand U4286 (N_4286,N_3910,N_3853);
nand U4287 (N_4287,N_3736,N_3514);
nand U4288 (N_4288,N_3565,N_3971);
xor U4289 (N_4289,N_3703,N_3957);
and U4290 (N_4290,N_3655,N_3618);
or U4291 (N_4291,N_3597,N_3769);
nand U4292 (N_4292,N_3742,N_3859);
xnor U4293 (N_4293,N_3530,N_3917);
nor U4294 (N_4294,N_3951,N_3848);
nand U4295 (N_4295,N_3549,N_3676);
nand U4296 (N_4296,N_3793,N_3613);
or U4297 (N_4297,N_3701,N_3590);
nand U4298 (N_4298,N_3936,N_3827);
nand U4299 (N_4299,N_3947,N_3994);
and U4300 (N_4300,N_3949,N_3595);
or U4301 (N_4301,N_3798,N_3631);
xnor U4302 (N_4302,N_3847,N_3874);
nand U4303 (N_4303,N_3619,N_3680);
nand U4304 (N_4304,N_3684,N_3721);
or U4305 (N_4305,N_3737,N_3630);
or U4306 (N_4306,N_3819,N_3917);
and U4307 (N_4307,N_3942,N_3771);
and U4308 (N_4308,N_3571,N_3554);
and U4309 (N_4309,N_3867,N_3862);
nor U4310 (N_4310,N_3839,N_3529);
nor U4311 (N_4311,N_3676,N_3820);
and U4312 (N_4312,N_3705,N_3967);
and U4313 (N_4313,N_3786,N_3950);
or U4314 (N_4314,N_3952,N_3521);
or U4315 (N_4315,N_3876,N_3941);
and U4316 (N_4316,N_3517,N_3789);
nor U4317 (N_4317,N_3898,N_3893);
nand U4318 (N_4318,N_3519,N_3938);
and U4319 (N_4319,N_3713,N_3723);
or U4320 (N_4320,N_3736,N_3732);
nand U4321 (N_4321,N_3594,N_3921);
xor U4322 (N_4322,N_3529,N_3625);
xnor U4323 (N_4323,N_3513,N_3835);
nor U4324 (N_4324,N_3868,N_3639);
nor U4325 (N_4325,N_3766,N_3665);
nand U4326 (N_4326,N_3721,N_3995);
or U4327 (N_4327,N_3912,N_3986);
and U4328 (N_4328,N_3761,N_3809);
nor U4329 (N_4329,N_3718,N_3764);
and U4330 (N_4330,N_3706,N_3757);
or U4331 (N_4331,N_3782,N_3502);
and U4332 (N_4332,N_3764,N_3820);
or U4333 (N_4333,N_3880,N_3582);
xnor U4334 (N_4334,N_3991,N_3764);
and U4335 (N_4335,N_3970,N_3797);
nor U4336 (N_4336,N_3902,N_3974);
nand U4337 (N_4337,N_3675,N_3945);
or U4338 (N_4338,N_3982,N_3956);
xor U4339 (N_4339,N_3648,N_3927);
xnor U4340 (N_4340,N_3717,N_3760);
and U4341 (N_4341,N_3975,N_3786);
or U4342 (N_4342,N_3946,N_3725);
and U4343 (N_4343,N_3844,N_3501);
xor U4344 (N_4344,N_3931,N_3773);
or U4345 (N_4345,N_3629,N_3621);
xor U4346 (N_4346,N_3979,N_3772);
nand U4347 (N_4347,N_3743,N_3730);
nand U4348 (N_4348,N_3524,N_3818);
and U4349 (N_4349,N_3763,N_3574);
and U4350 (N_4350,N_3938,N_3884);
nand U4351 (N_4351,N_3983,N_3746);
xor U4352 (N_4352,N_3734,N_3750);
or U4353 (N_4353,N_3957,N_3881);
nand U4354 (N_4354,N_3681,N_3932);
nor U4355 (N_4355,N_3776,N_3955);
nor U4356 (N_4356,N_3628,N_3945);
xnor U4357 (N_4357,N_3989,N_3604);
and U4358 (N_4358,N_3843,N_3922);
or U4359 (N_4359,N_3727,N_3671);
and U4360 (N_4360,N_3820,N_3973);
nand U4361 (N_4361,N_3848,N_3564);
nand U4362 (N_4362,N_3581,N_3967);
xor U4363 (N_4363,N_3776,N_3675);
nand U4364 (N_4364,N_3750,N_3678);
or U4365 (N_4365,N_3926,N_3911);
nand U4366 (N_4366,N_3825,N_3634);
nor U4367 (N_4367,N_3933,N_3910);
nand U4368 (N_4368,N_3719,N_3562);
or U4369 (N_4369,N_3706,N_3530);
nand U4370 (N_4370,N_3901,N_3719);
nand U4371 (N_4371,N_3717,N_3620);
nand U4372 (N_4372,N_3918,N_3716);
or U4373 (N_4373,N_3880,N_3825);
xor U4374 (N_4374,N_3704,N_3950);
xor U4375 (N_4375,N_3783,N_3697);
nand U4376 (N_4376,N_3919,N_3529);
and U4377 (N_4377,N_3913,N_3631);
or U4378 (N_4378,N_3535,N_3842);
nand U4379 (N_4379,N_3604,N_3534);
nand U4380 (N_4380,N_3707,N_3732);
xor U4381 (N_4381,N_3530,N_3862);
nor U4382 (N_4382,N_3901,N_3825);
or U4383 (N_4383,N_3723,N_3831);
nor U4384 (N_4384,N_3866,N_3961);
xnor U4385 (N_4385,N_3713,N_3868);
xor U4386 (N_4386,N_3688,N_3509);
and U4387 (N_4387,N_3885,N_3650);
nand U4388 (N_4388,N_3959,N_3606);
or U4389 (N_4389,N_3858,N_3961);
nor U4390 (N_4390,N_3923,N_3772);
and U4391 (N_4391,N_3703,N_3641);
xor U4392 (N_4392,N_3519,N_3524);
nor U4393 (N_4393,N_3577,N_3546);
xnor U4394 (N_4394,N_3953,N_3783);
xnor U4395 (N_4395,N_3814,N_3501);
nand U4396 (N_4396,N_3620,N_3918);
and U4397 (N_4397,N_3669,N_3731);
or U4398 (N_4398,N_3635,N_3845);
nand U4399 (N_4399,N_3515,N_3705);
and U4400 (N_4400,N_3774,N_3753);
or U4401 (N_4401,N_3565,N_3684);
xor U4402 (N_4402,N_3752,N_3968);
xnor U4403 (N_4403,N_3908,N_3899);
and U4404 (N_4404,N_3910,N_3506);
or U4405 (N_4405,N_3647,N_3503);
or U4406 (N_4406,N_3888,N_3993);
and U4407 (N_4407,N_3606,N_3820);
or U4408 (N_4408,N_3591,N_3546);
nor U4409 (N_4409,N_3660,N_3815);
nor U4410 (N_4410,N_3726,N_3579);
and U4411 (N_4411,N_3818,N_3874);
or U4412 (N_4412,N_3539,N_3684);
nand U4413 (N_4413,N_3979,N_3591);
xor U4414 (N_4414,N_3859,N_3916);
nor U4415 (N_4415,N_3805,N_3721);
nand U4416 (N_4416,N_3766,N_3595);
nand U4417 (N_4417,N_3960,N_3796);
or U4418 (N_4418,N_3629,N_3617);
xnor U4419 (N_4419,N_3720,N_3758);
or U4420 (N_4420,N_3963,N_3914);
or U4421 (N_4421,N_3846,N_3974);
xor U4422 (N_4422,N_3571,N_3757);
and U4423 (N_4423,N_3507,N_3563);
nor U4424 (N_4424,N_3941,N_3690);
nand U4425 (N_4425,N_3676,N_3712);
nand U4426 (N_4426,N_3807,N_3582);
xnor U4427 (N_4427,N_3647,N_3756);
or U4428 (N_4428,N_3708,N_3820);
nand U4429 (N_4429,N_3926,N_3758);
nand U4430 (N_4430,N_3703,N_3880);
nor U4431 (N_4431,N_3726,N_3752);
nand U4432 (N_4432,N_3738,N_3611);
nand U4433 (N_4433,N_3624,N_3750);
nand U4434 (N_4434,N_3972,N_3938);
nand U4435 (N_4435,N_3973,N_3983);
nand U4436 (N_4436,N_3765,N_3738);
nand U4437 (N_4437,N_3721,N_3772);
nand U4438 (N_4438,N_3658,N_3754);
and U4439 (N_4439,N_3949,N_3555);
nor U4440 (N_4440,N_3508,N_3507);
xor U4441 (N_4441,N_3750,N_3721);
and U4442 (N_4442,N_3631,N_3639);
and U4443 (N_4443,N_3630,N_3611);
or U4444 (N_4444,N_3707,N_3931);
nand U4445 (N_4445,N_3788,N_3705);
or U4446 (N_4446,N_3754,N_3719);
nor U4447 (N_4447,N_3559,N_3622);
nor U4448 (N_4448,N_3981,N_3816);
and U4449 (N_4449,N_3945,N_3714);
or U4450 (N_4450,N_3684,N_3958);
nand U4451 (N_4451,N_3855,N_3682);
nor U4452 (N_4452,N_3531,N_3961);
nand U4453 (N_4453,N_3592,N_3774);
nand U4454 (N_4454,N_3771,N_3814);
nor U4455 (N_4455,N_3978,N_3567);
and U4456 (N_4456,N_3557,N_3730);
or U4457 (N_4457,N_3758,N_3680);
and U4458 (N_4458,N_3657,N_3585);
or U4459 (N_4459,N_3605,N_3789);
and U4460 (N_4460,N_3845,N_3784);
nor U4461 (N_4461,N_3741,N_3530);
and U4462 (N_4462,N_3841,N_3666);
or U4463 (N_4463,N_3756,N_3738);
and U4464 (N_4464,N_3658,N_3645);
or U4465 (N_4465,N_3527,N_3858);
xor U4466 (N_4466,N_3672,N_3650);
xor U4467 (N_4467,N_3534,N_3561);
nand U4468 (N_4468,N_3586,N_3778);
and U4469 (N_4469,N_3883,N_3646);
nand U4470 (N_4470,N_3656,N_3962);
nand U4471 (N_4471,N_3979,N_3574);
xor U4472 (N_4472,N_3879,N_3627);
nor U4473 (N_4473,N_3836,N_3607);
xor U4474 (N_4474,N_3705,N_3810);
nand U4475 (N_4475,N_3696,N_3914);
nand U4476 (N_4476,N_3594,N_3798);
or U4477 (N_4477,N_3502,N_3664);
nor U4478 (N_4478,N_3506,N_3523);
nor U4479 (N_4479,N_3684,N_3696);
xor U4480 (N_4480,N_3864,N_3948);
xor U4481 (N_4481,N_3829,N_3606);
nor U4482 (N_4482,N_3625,N_3731);
or U4483 (N_4483,N_3660,N_3726);
nor U4484 (N_4484,N_3526,N_3643);
nor U4485 (N_4485,N_3712,N_3897);
nand U4486 (N_4486,N_3542,N_3552);
nor U4487 (N_4487,N_3768,N_3743);
or U4488 (N_4488,N_3937,N_3671);
nand U4489 (N_4489,N_3958,N_3649);
nand U4490 (N_4490,N_3508,N_3547);
nand U4491 (N_4491,N_3985,N_3905);
nor U4492 (N_4492,N_3501,N_3669);
nor U4493 (N_4493,N_3972,N_3648);
and U4494 (N_4494,N_3760,N_3712);
nand U4495 (N_4495,N_3695,N_3856);
xor U4496 (N_4496,N_3775,N_3772);
and U4497 (N_4497,N_3962,N_3800);
and U4498 (N_4498,N_3860,N_3675);
and U4499 (N_4499,N_3563,N_3989);
xnor U4500 (N_4500,N_4229,N_4198);
nand U4501 (N_4501,N_4097,N_4443);
nand U4502 (N_4502,N_4210,N_4247);
or U4503 (N_4503,N_4024,N_4311);
and U4504 (N_4504,N_4479,N_4172);
xor U4505 (N_4505,N_4269,N_4287);
or U4506 (N_4506,N_4262,N_4019);
and U4507 (N_4507,N_4179,N_4098);
and U4508 (N_4508,N_4038,N_4093);
or U4509 (N_4509,N_4017,N_4104);
nand U4510 (N_4510,N_4480,N_4185);
nor U4511 (N_4511,N_4232,N_4349);
and U4512 (N_4512,N_4228,N_4113);
and U4513 (N_4513,N_4096,N_4066);
and U4514 (N_4514,N_4486,N_4469);
and U4515 (N_4515,N_4495,N_4295);
or U4516 (N_4516,N_4300,N_4277);
nand U4517 (N_4517,N_4355,N_4122);
xnor U4518 (N_4518,N_4099,N_4014);
or U4519 (N_4519,N_4147,N_4164);
nand U4520 (N_4520,N_4379,N_4466);
nand U4521 (N_4521,N_4196,N_4163);
xor U4522 (N_4522,N_4442,N_4430);
nor U4523 (N_4523,N_4450,N_4491);
nor U4524 (N_4524,N_4174,N_4129);
or U4525 (N_4525,N_4286,N_4380);
and U4526 (N_4526,N_4411,N_4091);
and U4527 (N_4527,N_4125,N_4114);
xnor U4528 (N_4528,N_4165,N_4485);
nor U4529 (N_4529,N_4244,N_4094);
xnor U4530 (N_4530,N_4472,N_4463);
nand U4531 (N_4531,N_4135,N_4307);
or U4532 (N_4532,N_4461,N_4141);
nor U4533 (N_4533,N_4157,N_4256);
nor U4534 (N_4534,N_4366,N_4407);
nand U4535 (N_4535,N_4376,N_4102);
nor U4536 (N_4536,N_4271,N_4230);
xor U4537 (N_4537,N_4358,N_4332);
or U4538 (N_4538,N_4206,N_4464);
nand U4539 (N_4539,N_4248,N_4103);
nand U4540 (N_4540,N_4352,N_4363);
or U4541 (N_4541,N_4436,N_4148);
nand U4542 (N_4542,N_4426,N_4109);
nor U4543 (N_4543,N_4181,N_4496);
nor U4544 (N_4544,N_4408,N_4108);
and U4545 (N_4545,N_4333,N_4153);
xnor U4546 (N_4546,N_4137,N_4123);
or U4547 (N_4547,N_4126,N_4204);
or U4548 (N_4548,N_4007,N_4351);
or U4549 (N_4549,N_4004,N_4214);
nand U4550 (N_4550,N_4315,N_4342);
nand U4551 (N_4551,N_4487,N_4133);
or U4552 (N_4552,N_4305,N_4199);
and U4553 (N_4553,N_4494,N_4360);
xnor U4554 (N_4554,N_4321,N_4111);
or U4555 (N_4555,N_4330,N_4193);
and U4556 (N_4556,N_4130,N_4465);
nor U4557 (N_4557,N_4418,N_4377);
nor U4558 (N_4558,N_4023,N_4467);
or U4559 (N_4559,N_4219,N_4057);
xor U4560 (N_4560,N_4266,N_4370);
nor U4561 (N_4561,N_4394,N_4453);
xnor U4562 (N_4562,N_4470,N_4446);
xnor U4563 (N_4563,N_4184,N_4150);
nand U4564 (N_4564,N_4209,N_4237);
xnor U4565 (N_4565,N_4183,N_4278);
nor U4566 (N_4566,N_4420,N_4445);
nor U4567 (N_4567,N_4387,N_4346);
nand U4568 (N_4568,N_4146,N_4044);
xnor U4569 (N_4569,N_4344,N_4251);
or U4570 (N_4570,N_4434,N_4216);
or U4571 (N_4571,N_4390,N_4213);
xor U4572 (N_4572,N_4492,N_4238);
and U4573 (N_4573,N_4144,N_4364);
nor U4574 (N_4574,N_4036,N_4059);
or U4575 (N_4575,N_4325,N_4161);
nor U4576 (N_4576,N_4458,N_4138);
nor U4577 (N_4577,N_4200,N_4233);
or U4578 (N_4578,N_4421,N_4030);
and U4579 (N_4579,N_4134,N_4497);
or U4580 (N_4580,N_4312,N_4025);
nand U4581 (N_4581,N_4428,N_4357);
xor U4582 (N_4582,N_4293,N_4063);
nor U4583 (N_4583,N_4289,N_4035);
nor U4584 (N_4584,N_4031,N_4086);
xnor U4585 (N_4585,N_4477,N_4338);
or U4586 (N_4586,N_4462,N_4431);
nor U4587 (N_4587,N_4043,N_4404);
or U4588 (N_4588,N_4132,N_4076);
nor U4589 (N_4589,N_4118,N_4062);
and U4590 (N_4590,N_4074,N_4382);
and U4591 (N_4591,N_4476,N_4362);
nand U4592 (N_4592,N_4499,N_4197);
xor U4593 (N_4593,N_4245,N_4011);
nand U4594 (N_4594,N_4003,N_4396);
or U4595 (N_4595,N_4010,N_4265);
xnor U4596 (N_4596,N_4455,N_4367);
nand U4597 (N_4597,N_4393,N_4322);
or U4598 (N_4598,N_4084,N_4303);
nand U4599 (N_4599,N_4423,N_4166);
nand U4600 (N_4600,N_4405,N_4128);
and U4601 (N_4601,N_4309,N_4227);
and U4602 (N_4602,N_4397,N_4054);
or U4603 (N_4603,N_4107,N_4241);
or U4604 (N_4604,N_4015,N_4211);
and U4605 (N_4605,N_4456,N_4273);
nand U4606 (N_4606,N_4173,N_4026);
nand U4607 (N_4607,N_4222,N_4317);
xnor U4608 (N_4608,N_4383,N_4432);
nor U4609 (N_4609,N_4270,N_4037);
xnor U4610 (N_4610,N_4186,N_4374);
nand U4611 (N_4611,N_4116,N_4279);
and U4612 (N_4612,N_4369,N_4047);
nand U4613 (N_4613,N_4473,N_4437);
or U4614 (N_4614,N_4429,N_4189);
or U4615 (N_4615,N_4159,N_4140);
nand U4616 (N_4616,N_4253,N_4373);
nand U4617 (N_4617,N_4051,N_4168);
xnor U4618 (N_4618,N_4061,N_4410);
or U4619 (N_4619,N_4398,N_4482);
nor U4620 (N_4620,N_4090,N_4267);
nor U4621 (N_4621,N_4117,N_4053);
and U4622 (N_4622,N_4281,N_4202);
and U4623 (N_4623,N_4016,N_4291);
or U4624 (N_4624,N_4389,N_4208);
or U4625 (N_4625,N_4155,N_4112);
xnor U4626 (N_4626,N_4257,N_4177);
xnor U4627 (N_4627,N_4060,N_4223);
nor U4628 (N_4628,N_4039,N_4475);
or U4629 (N_4629,N_4288,N_4478);
or U4630 (N_4630,N_4081,N_4386);
xnor U4631 (N_4631,N_4250,N_4336);
xor U4632 (N_4632,N_4064,N_4029);
xor U4633 (N_4633,N_4018,N_4127);
nor U4634 (N_4634,N_4215,N_4483);
and U4635 (N_4635,N_4335,N_4220);
nand U4636 (N_4636,N_4041,N_4368);
and U4637 (N_4637,N_4079,N_4145);
or U4638 (N_4638,N_4224,N_4070);
nand U4639 (N_4639,N_4028,N_4372);
xnor U4640 (N_4640,N_4182,N_4371);
xnor U4641 (N_4641,N_4195,N_4488);
xor U4642 (N_4642,N_4381,N_4378);
nand U4643 (N_4643,N_4484,N_4457);
and U4644 (N_4644,N_4318,N_4105);
nor U4645 (N_4645,N_4136,N_4027);
nor U4646 (N_4646,N_4474,N_4399);
and U4647 (N_4647,N_4106,N_4152);
nand U4648 (N_4648,N_4424,N_4190);
nor U4649 (N_4649,N_4260,N_4331);
nand U4650 (N_4650,N_4348,N_4042);
or U4651 (N_4651,N_4416,N_4412);
nand U4652 (N_4652,N_4313,N_4045);
and U4653 (N_4653,N_4236,N_4121);
nor U4654 (N_4654,N_4217,N_4449);
and U4655 (N_4655,N_4441,N_4391);
or U4656 (N_4656,N_4304,N_4100);
xor U4657 (N_4657,N_4069,N_4032);
xor U4658 (N_4658,N_4264,N_4320);
nor U4659 (N_4659,N_4268,N_4323);
nor U4660 (N_4660,N_4192,N_4249);
xnor U4661 (N_4661,N_4154,N_4075);
nor U4662 (N_4662,N_4340,N_4298);
or U4663 (N_4663,N_4329,N_4403);
xor U4664 (N_4664,N_4252,N_4427);
and U4665 (N_4665,N_4359,N_4046);
or U4666 (N_4666,N_4156,N_4115);
and U4667 (N_4667,N_4422,N_4120);
or U4668 (N_4668,N_4083,N_4337);
nor U4669 (N_4669,N_4440,N_4413);
nand U4670 (N_4670,N_4008,N_4065);
nand U4671 (N_4671,N_4048,N_4071);
xnor U4672 (N_4672,N_4176,N_4400);
nor U4673 (N_4673,N_4297,N_4301);
xnor U4674 (N_4674,N_4385,N_4218);
or U4675 (N_4675,N_4272,N_4077);
or U4676 (N_4676,N_4101,N_4392);
and U4677 (N_4677,N_4080,N_4341);
or U4678 (N_4678,N_4388,N_4055);
or U4679 (N_4679,N_4406,N_4020);
and U4680 (N_4680,N_4231,N_4384);
or U4681 (N_4681,N_4324,N_4021);
and U4682 (N_4682,N_4149,N_4275);
nor U4683 (N_4683,N_4205,N_4243);
nor U4684 (N_4684,N_4082,N_4263);
nor U4685 (N_4685,N_4292,N_4162);
nand U4686 (N_4686,N_4188,N_4092);
and U4687 (N_4687,N_4191,N_4415);
xnor U4688 (N_4688,N_4451,N_4012);
xor U4689 (N_4689,N_4178,N_4239);
nand U4690 (N_4690,N_4435,N_4087);
xor U4691 (N_4691,N_4258,N_4274);
and U4692 (N_4692,N_4319,N_4171);
xnor U4693 (N_4693,N_4068,N_4327);
nor U4694 (N_4694,N_4498,N_4361);
and U4695 (N_4695,N_4234,N_4095);
nor U4696 (N_4696,N_4306,N_4414);
and U4697 (N_4697,N_4447,N_4124);
nand U4698 (N_4698,N_4481,N_4471);
or U4699 (N_4699,N_4169,N_4294);
or U4700 (N_4700,N_4131,N_4139);
nand U4701 (N_4701,N_4085,N_4459);
nand U4702 (N_4702,N_4240,N_4034);
and U4703 (N_4703,N_4354,N_4246);
nand U4704 (N_4704,N_4290,N_4006);
or U4705 (N_4705,N_4401,N_4326);
and U4706 (N_4706,N_4187,N_4242);
nor U4707 (N_4707,N_4142,N_4143);
nand U4708 (N_4708,N_4347,N_4050);
nor U4709 (N_4709,N_4439,N_4402);
or U4710 (N_4710,N_4261,N_4067);
nor U4711 (N_4711,N_4282,N_4203);
nand U4712 (N_4712,N_4078,N_4255);
nand U4713 (N_4713,N_4259,N_4343);
and U4714 (N_4714,N_4073,N_4180);
and U4715 (N_4715,N_4058,N_4052);
nand U4716 (N_4716,N_4119,N_4170);
nand U4717 (N_4717,N_4089,N_4158);
xnor U4718 (N_4718,N_4225,N_4284);
xnor U4719 (N_4719,N_4444,N_4452);
or U4720 (N_4720,N_4285,N_4493);
and U4721 (N_4721,N_4490,N_4151);
xor U4722 (N_4722,N_4448,N_4207);
or U4723 (N_4723,N_4002,N_4302);
xnor U4724 (N_4724,N_4001,N_4088);
or U4725 (N_4725,N_4460,N_4235);
nand U4726 (N_4726,N_4356,N_4334);
nor U4727 (N_4727,N_4438,N_4417);
xnor U4728 (N_4728,N_4345,N_4419);
nor U4729 (N_4729,N_4254,N_4296);
or U4730 (N_4730,N_4425,N_4072);
and U4731 (N_4731,N_4299,N_4350);
or U4732 (N_4732,N_4310,N_4033);
and U4733 (N_4733,N_4489,N_4283);
xnor U4734 (N_4734,N_4276,N_4221);
nand U4735 (N_4735,N_4468,N_4175);
and U4736 (N_4736,N_4040,N_4013);
xnor U4737 (N_4737,N_4194,N_4316);
or U4738 (N_4738,N_4022,N_4353);
nor U4739 (N_4739,N_4314,N_4308);
xnor U4740 (N_4740,N_4056,N_4005);
nor U4741 (N_4741,N_4433,N_4454);
or U4742 (N_4742,N_4365,N_4375);
nand U4743 (N_4743,N_4167,N_4110);
nand U4744 (N_4744,N_4339,N_4201);
nor U4745 (N_4745,N_4212,N_4049);
and U4746 (N_4746,N_4009,N_4226);
xnor U4747 (N_4747,N_4280,N_4160);
nand U4748 (N_4748,N_4328,N_4395);
nand U4749 (N_4749,N_4000,N_4409);
or U4750 (N_4750,N_4024,N_4373);
xnor U4751 (N_4751,N_4248,N_4434);
nand U4752 (N_4752,N_4480,N_4355);
or U4753 (N_4753,N_4296,N_4147);
nor U4754 (N_4754,N_4203,N_4453);
nor U4755 (N_4755,N_4396,N_4023);
nor U4756 (N_4756,N_4464,N_4180);
and U4757 (N_4757,N_4271,N_4272);
xnor U4758 (N_4758,N_4194,N_4276);
and U4759 (N_4759,N_4178,N_4273);
xor U4760 (N_4760,N_4170,N_4415);
nor U4761 (N_4761,N_4236,N_4487);
and U4762 (N_4762,N_4326,N_4264);
xnor U4763 (N_4763,N_4410,N_4030);
xor U4764 (N_4764,N_4064,N_4384);
and U4765 (N_4765,N_4356,N_4111);
xor U4766 (N_4766,N_4071,N_4049);
or U4767 (N_4767,N_4420,N_4085);
xor U4768 (N_4768,N_4252,N_4275);
and U4769 (N_4769,N_4073,N_4431);
nand U4770 (N_4770,N_4051,N_4077);
nand U4771 (N_4771,N_4245,N_4259);
xnor U4772 (N_4772,N_4290,N_4478);
or U4773 (N_4773,N_4131,N_4489);
nor U4774 (N_4774,N_4486,N_4412);
or U4775 (N_4775,N_4202,N_4437);
nand U4776 (N_4776,N_4482,N_4063);
xnor U4777 (N_4777,N_4105,N_4054);
or U4778 (N_4778,N_4023,N_4191);
nor U4779 (N_4779,N_4442,N_4326);
or U4780 (N_4780,N_4321,N_4330);
nor U4781 (N_4781,N_4240,N_4118);
nor U4782 (N_4782,N_4130,N_4074);
and U4783 (N_4783,N_4470,N_4380);
or U4784 (N_4784,N_4413,N_4368);
nand U4785 (N_4785,N_4312,N_4089);
xnor U4786 (N_4786,N_4114,N_4018);
nand U4787 (N_4787,N_4477,N_4480);
xnor U4788 (N_4788,N_4085,N_4049);
or U4789 (N_4789,N_4481,N_4240);
nor U4790 (N_4790,N_4130,N_4327);
nor U4791 (N_4791,N_4368,N_4180);
and U4792 (N_4792,N_4015,N_4370);
and U4793 (N_4793,N_4408,N_4430);
nor U4794 (N_4794,N_4142,N_4416);
nor U4795 (N_4795,N_4291,N_4195);
or U4796 (N_4796,N_4183,N_4405);
nand U4797 (N_4797,N_4360,N_4465);
or U4798 (N_4798,N_4266,N_4094);
or U4799 (N_4799,N_4146,N_4388);
nor U4800 (N_4800,N_4074,N_4028);
nor U4801 (N_4801,N_4209,N_4436);
nand U4802 (N_4802,N_4151,N_4378);
and U4803 (N_4803,N_4042,N_4237);
xnor U4804 (N_4804,N_4296,N_4333);
or U4805 (N_4805,N_4342,N_4007);
or U4806 (N_4806,N_4095,N_4437);
and U4807 (N_4807,N_4076,N_4488);
nor U4808 (N_4808,N_4473,N_4250);
xor U4809 (N_4809,N_4136,N_4081);
nor U4810 (N_4810,N_4340,N_4168);
nand U4811 (N_4811,N_4232,N_4324);
nand U4812 (N_4812,N_4216,N_4189);
and U4813 (N_4813,N_4431,N_4448);
nand U4814 (N_4814,N_4235,N_4397);
nor U4815 (N_4815,N_4097,N_4031);
and U4816 (N_4816,N_4058,N_4121);
and U4817 (N_4817,N_4174,N_4096);
xnor U4818 (N_4818,N_4350,N_4091);
xnor U4819 (N_4819,N_4191,N_4478);
nor U4820 (N_4820,N_4454,N_4046);
and U4821 (N_4821,N_4223,N_4266);
xnor U4822 (N_4822,N_4268,N_4369);
or U4823 (N_4823,N_4440,N_4019);
and U4824 (N_4824,N_4113,N_4087);
and U4825 (N_4825,N_4373,N_4219);
nand U4826 (N_4826,N_4447,N_4186);
or U4827 (N_4827,N_4173,N_4051);
nor U4828 (N_4828,N_4019,N_4352);
nor U4829 (N_4829,N_4449,N_4404);
nor U4830 (N_4830,N_4123,N_4129);
nand U4831 (N_4831,N_4401,N_4462);
nand U4832 (N_4832,N_4369,N_4498);
xor U4833 (N_4833,N_4350,N_4237);
or U4834 (N_4834,N_4488,N_4015);
nor U4835 (N_4835,N_4292,N_4073);
nor U4836 (N_4836,N_4357,N_4447);
xnor U4837 (N_4837,N_4351,N_4367);
xor U4838 (N_4838,N_4310,N_4009);
or U4839 (N_4839,N_4306,N_4312);
xnor U4840 (N_4840,N_4288,N_4078);
xor U4841 (N_4841,N_4152,N_4095);
and U4842 (N_4842,N_4272,N_4031);
nand U4843 (N_4843,N_4215,N_4212);
nor U4844 (N_4844,N_4476,N_4132);
or U4845 (N_4845,N_4052,N_4175);
nor U4846 (N_4846,N_4402,N_4382);
xor U4847 (N_4847,N_4461,N_4142);
xnor U4848 (N_4848,N_4154,N_4298);
xor U4849 (N_4849,N_4246,N_4350);
nor U4850 (N_4850,N_4003,N_4168);
nand U4851 (N_4851,N_4121,N_4131);
xor U4852 (N_4852,N_4164,N_4247);
xor U4853 (N_4853,N_4482,N_4024);
nor U4854 (N_4854,N_4344,N_4018);
nand U4855 (N_4855,N_4008,N_4044);
xor U4856 (N_4856,N_4422,N_4334);
nand U4857 (N_4857,N_4253,N_4139);
and U4858 (N_4858,N_4386,N_4379);
or U4859 (N_4859,N_4430,N_4267);
or U4860 (N_4860,N_4179,N_4338);
or U4861 (N_4861,N_4109,N_4312);
or U4862 (N_4862,N_4128,N_4150);
nand U4863 (N_4863,N_4209,N_4352);
and U4864 (N_4864,N_4350,N_4168);
xor U4865 (N_4865,N_4245,N_4167);
xor U4866 (N_4866,N_4006,N_4481);
nand U4867 (N_4867,N_4199,N_4361);
and U4868 (N_4868,N_4059,N_4386);
and U4869 (N_4869,N_4362,N_4110);
and U4870 (N_4870,N_4309,N_4045);
nand U4871 (N_4871,N_4257,N_4079);
nand U4872 (N_4872,N_4393,N_4297);
and U4873 (N_4873,N_4440,N_4013);
xor U4874 (N_4874,N_4178,N_4426);
nand U4875 (N_4875,N_4427,N_4265);
or U4876 (N_4876,N_4337,N_4393);
or U4877 (N_4877,N_4238,N_4162);
or U4878 (N_4878,N_4132,N_4109);
xnor U4879 (N_4879,N_4371,N_4205);
nand U4880 (N_4880,N_4183,N_4450);
nor U4881 (N_4881,N_4256,N_4426);
nor U4882 (N_4882,N_4368,N_4406);
and U4883 (N_4883,N_4446,N_4283);
nand U4884 (N_4884,N_4365,N_4381);
and U4885 (N_4885,N_4494,N_4396);
xor U4886 (N_4886,N_4319,N_4429);
or U4887 (N_4887,N_4279,N_4401);
nor U4888 (N_4888,N_4158,N_4041);
xnor U4889 (N_4889,N_4421,N_4189);
and U4890 (N_4890,N_4371,N_4251);
xnor U4891 (N_4891,N_4156,N_4314);
nand U4892 (N_4892,N_4396,N_4168);
nand U4893 (N_4893,N_4417,N_4254);
xnor U4894 (N_4894,N_4321,N_4469);
nor U4895 (N_4895,N_4002,N_4109);
and U4896 (N_4896,N_4238,N_4260);
xor U4897 (N_4897,N_4238,N_4490);
xnor U4898 (N_4898,N_4265,N_4378);
xor U4899 (N_4899,N_4432,N_4366);
xnor U4900 (N_4900,N_4288,N_4302);
or U4901 (N_4901,N_4369,N_4089);
or U4902 (N_4902,N_4483,N_4024);
nor U4903 (N_4903,N_4132,N_4357);
xor U4904 (N_4904,N_4396,N_4443);
nand U4905 (N_4905,N_4146,N_4252);
and U4906 (N_4906,N_4244,N_4235);
nand U4907 (N_4907,N_4432,N_4357);
xor U4908 (N_4908,N_4040,N_4324);
and U4909 (N_4909,N_4414,N_4089);
xnor U4910 (N_4910,N_4248,N_4057);
nor U4911 (N_4911,N_4260,N_4056);
nand U4912 (N_4912,N_4255,N_4280);
nor U4913 (N_4913,N_4231,N_4138);
nand U4914 (N_4914,N_4123,N_4162);
nand U4915 (N_4915,N_4211,N_4292);
xnor U4916 (N_4916,N_4059,N_4335);
and U4917 (N_4917,N_4082,N_4141);
nand U4918 (N_4918,N_4065,N_4197);
xor U4919 (N_4919,N_4428,N_4124);
nor U4920 (N_4920,N_4187,N_4465);
xnor U4921 (N_4921,N_4423,N_4111);
nor U4922 (N_4922,N_4445,N_4457);
xor U4923 (N_4923,N_4391,N_4263);
and U4924 (N_4924,N_4127,N_4200);
xnor U4925 (N_4925,N_4092,N_4229);
xnor U4926 (N_4926,N_4217,N_4097);
nor U4927 (N_4927,N_4266,N_4165);
nand U4928 (N_4928,N_4382,N_4090);
and U4929 (N_4929,N_4379,N_4245);
nor U4930 (N_4930,N_4297,N_4302);
and U4931 (N_4931,N_4030,N_4166);
nand U4932 (N_4932,N_4275,N_4122);
nand U4933 (N_4933,N_4461,N_4052);
or U4934 (N_4934,N_4399,N_4202);
xor U4935 (N_4935,N_4375,N_4015);
and U4936 (N_4936,N_4263,N_4160);
nand U4937 (N_4937,N_4278,N_4292);
nor U4938 (N_4938,N_4288,N_4111);
nand U4939 (N_4939,N_4426,N_4375);
or U4940 (N_4940,N_4239,N_4317);
nand U4941 (N_4941,N_4186,N_4203);
and U4942 (N_4942,N_4117,N_4178);
xnor U4943 (N_4943,N_4000,N_4120);
and U4944 (N_4944,N_4414,N_4052);
xnor U4945 (N_4945,N_4288,N_4475);
or U4946 (N_4946,N_4384,N_4077);
nand U4947 (N_4947,N_4041,N_4206);
xor U4948 (N_4948,N_4062,N_4223);
and U4949 (N_4949,N_4049,N_4360);
and U4950 (N_4950,N_4254,N_4159);
xor U4951 (N_4951,N_4200,N_4298);
or U4952 (N_4952,N_4482,N_4466);
nand U4953 (N_4953,N_4280,N_4032);
and U4954 (N_4954,N_4187,N_4179);
nor U4955 (N_4955,N_4109,N_4247);
or U4956 (N_4956,N_4336,N_4194);
or U4957 (N_4957,N_4352,N_4050);
nor U4958 (N_4958,N_4384,N_4460);
and U4959 (N_4959,N_4364,N_4029);
nand U4960 (N_4960,N_4287,N_4315);
nand U4961 (N_4961,N_4200,N_4225);
xnor U4962 (N_4962,N_4417,N_4293);
xor U4963 (N_4963,N_4106,N_4079);
nand U4964 (N_4964,N_4169,N_4130);
nor U4965 (N_4965,N_4279,N_4308);
and U4966 (N_4966,N_4274,N_4304);
nand U4967 (N_4967,N_4303,N_4473);
or U4968 (N_4968,N_4473,N_4018);
nor U4969 (N_4969,N_4045,N_4065);
xnor U4970 (N_4970,N_4423,N_4173);
and U4971 (N_4971,N_4304,N_4073);
and U4972 (N_4972,N_4115,N_4360);
nand U4973 (N_4973,N_4425,N_4312);
xor U4974 (N_4974,N_4024,N_4276);
or U4975 (N_4975,N_4053,N_4445);
xor U4976 (N_4976,N_4053,N_4061);
or U4977 (N_4977,N_4411,N_4247);
and U4978 (N_4978,N_4157,N_4209);
xor U4979 (N_4979,N_4073,N_4106);
nor U4980 (N_4980,N_4423,N_4219);
and U4981 (N_4981,N_4451,N_4430);
xor U4982 (N_4982,N_4289,N_4108);
nor U4983 (N_4983,N_4136,N_4230);
or U4984 (N_4984,N_4113,N_4384);
nor U4985 (N_4985,N_4122,N_4099);
nor U4986 (N_4986,N_4196,N_4259);
and U4987 (N_4987,N_4123,N_4259);
nor U4988 (N_4988,N_4286,N_4155);
nand U4989 (N_4989,N_4201,N_4100);
nand U4990 (N_4990,N_4081,N_4153);
nor U4991 (N_4991,N_4152,N_4434);
nor U4992 (N_4992,N_4080,N_4163);
nand U4993 (N_4993,N_4459,N_4106);
or U4994 (N_4994,N_4155,N_4311);
and U4995 (N_4995,N_4284,N_4241);
or U4996 (N_4996,N_4361,N_4195);
and U4997 (N_4997,N_4316,N_4058);
and U4998 (N_4998,N_4104,N_4158);
or U4999 (N_4999,N_4017,N_4037);
or U5000 (N_5000,N_4724,N_4966);
and U5001 (N_5001,N_4763,N_4872);
and U5002 (N_5002,N_4714,N_4535);
nor U5003 (N_5003,N_4762,N_4732);
and U5004 (N_5004,N_4868,N_4682);
xor U5005 (N_5005,N_4978,N_4559);
nand U5006 (N_5006,N_4787,N_4963);
nor U5007 (N_5007,N_4620,N_4687);
or U5008 (N_5008,N_4920,N_4610);
and U5009 (N_5009,N_4623,N_4648);
xor U5010 (N_5010,N_4696,N_4771);
nand U5011 (N_5011,N_4749,N_4924);
xnor U5012 (N_5012,N_4841,N_4901);
nand U5013 (N_5013,N_4852,N_4800);
and U5014 (N_5014,N_4776,N_4955);
or U5015 (N_5015,N_4946,N_4662);
nand U5016 (N_5016,N_4899,N_4839);
nand U5017 (N_5017,N_4542,N_4884);
nor U5018 (N_5018,N_4793,N_4590);
and U5019 (N_5019,N_4902,N_4900);
nor U5020 (N_5020,N_4862,N_4953);
nor U5021 (N_5021,N_4529,N_4616);
or U5022 (N_5022,N_4710,N_4971);
xor U5023 (N_5023,N_4723,N_4758);
nand U5024 (N_5024,N_4661,N_4842);
or U5025 (N_5025,N_4601,N_4995);
nand U5026 (N_5026,N_4861,N_4830);
nand U5027 (N_5027,N_4980,N_4999);
or U5028 (N_5028,N_4608,N_4572);
nor U5029 (N_5029,N_4904,N_4893);
xor U5030 (N_5030,N_4782,N_4936);
nand U5031 (N_5031,N_4961,N_4650);
nand U5032 (N_5032,N_4919,N_4840);
and U5033 (N_5033,N_4870,N_4792);
xor U5034 (N_5034,N_4905,N_4511);
or U5035 (N_5035,N_4979,N_4939);
nand U5036 (N_5036,N_4821,N_4533);
nor U5037 (N_5037,N_4863,N_4796);
nor U5038 (N_5038,N_4672,N_4715);
xor U5039 (N_5039,N_4618,N_4867);
xnor U5040 (N_5040,N_4640,N_4848);
xor U5041 (N_5041,N_4945,N_4778);
xnor U5042 (N_5042,N_4630,N_4673);
nor U5043 (N_5043,N_4909,N_4998);
or U5044 (N_5044,N_4865,N_4777);
nor U5045 (N_5045,N_4784,N_4697);
nand U5046 (N_5046,N_4949,N_4745);
nor U5047 (N_5047,N_4947,N_4752);
and U5048 (N_5048,N_4894,N_4910);
nand U5049 (N_5049,N_4578,N_4730);
or U5050 (N_5050,N_4587,N_4864);
or U5051 (N_5051,N_4605,N_4526);
nor U5052 (N_5052,N_4755,N_4689);
or U5053 (N_5053,N_4622,N_4935);
and U5054 (N_5054,N_4674,N_4825);
nand U5055 (N_5055,N_4850,N_4520);
xnor U5056 (N_5056,N_4898,N_4659);
or U5057 (N_5057,N_4907,N_4754);
or U5058 (N_5058,N_4964,N_4957);
and U5059 (N_5059,N_4958,N_4703);
and U5060 (N_5060,N_4582,N_4985);
nand U5061 (N_5061,N_4765,N_4568);
and U5062 (N_5062,N_4678,N_4942);
xor U5063 (N_5063,N_4744,N_4836);
and U5064 (N_5064,N_4604,N_4545);
nor U5065 (N_5065,N_4691,N_4737);
xnor U5066 (N_5066,N_4917,N_4888);
and U5067 (N_5067,N_4515,N_4562);
or U5068 (N_5068,N_4538,N_4834);
nand U5069 (N_5069,N_4510,N_4976);
nor U5070 (N_5070,N_4973,N_4873);
or U5071 (N_5071,N_4594,N_4619);
xnor U5072 (N_5072,N_4517,N_4783);
nand U5073 (N_5073,N_4932,N_4660);
nor U5074 (N_5074,N_4588,N_4531);
or U5075 (N_5075,N_4606,N_4555);
xnor U5076 (N_5076,N_4788,N_4600);
nand U5077 (N_5077,N_4720,N_4812);
or U5078 (N_5078,N_4719,N_4558);
and U5079 (N_5079,N_4746,N_4688);
nand U5080 (N_5080,N_4892,N_4532);
nand U5081 (N_5081,N_4882,N_4977);
xor U5082 (N_5082,N_4665,N_4641);
nand U5083 (N_5083,N_4943,N_4718);
nor U5084 (N_5084,N_4518,N_4785);
xnor U5085 (N_5085,N_4769,N_4704);
xor U5086 (N_5086,N_4611,N_4997);
nand U5087 (N_5087,N_4602,N_4599);
nor U5088 (N_5088,N_4613,N_4818);
nand U5089 (N_5089,N_4504,N_4926);
or U5090 (N_5090,N_4815,N_4759);
xor U5091 (N_5091,N_4933,N_4685);
nor U5092 (N_5092,N_4938,N_4743);
and U5093 (N_5093,N_4982,N_4856);
nor U5094 (N_5094,N_4584,N_4760);
xnor U5095 (N_5095,N_4657,N_4679);
nand U5096 (N_5096,N_4536,N_4524);
nand U5097 (N_5097,N_4652,N_4780);
and U5098 (N_5098,N_4645,N_4881);
and U5099 (N_5099,N_4811,N_4621);
nor U5100 (N_5100,N_4866,N_4670);
and U5101 (N_5101,N_4695,N_4607);
nand U5102 (N_5102,N_4734,N_4625);
and U5103 (N_5103,N_4740,N_4786);
nand U5104 (N_5104,N_4806,N_4757);
and U5105 (N_5105,N_4651,N_4557);
nor U5106 (N_5106,N_4553,N_4564);
nand U5107 (N_5107,N_4647,N_4684);
xnor U5108 (N_5108,N_4658,N_4772);
nand U5109 (N_5109,N_4883,N_4521);
nor U5110 (N_5110,N_4539,N_4874);
and U5111 (N_5111,N_4925,N_4628);
xor U5112 (N_5112,N_4992,N_4916);
nor U5113 (N_5113,N_4827,N_4911);
nor U5114 (N_5114,N_4574,N_4726);
nor U5115 (N_5115,N_4931,N_4950);
nand U5116 (N_5116,N_4844,N_4741);
and U5117 (N_5117,N_4692,N_4843);
nand U5118 (N_5118,N_4736,N_4956);
nor U5119 (N_5119,N_4716,N_4871);
and U5120 (N_5120,N_4891,N_4686);
and U5121 (N_5121,N_4879,N_4951);
and U5122 (N_5122,N_4937,N_4722);
or U5123 (N_5123,N_4617,N_4566);
nand U5124 (N_5124,N_4592,N_4857);
or U5125 (N_5125,N_4699,N_4913);
or U5126 (N_5126,N_4683,N_4975);
xor U5127 (N_5127,N_4808,N_4767);
nor U5128 (N_5128,N_4805,N_4912);
xnor U5129 (N_5129,N_4996,N_4634);
or U5130 (N_5130,N_4819,N_4537);
xnor U5131 (N_5131,N_4693,N_4575);
nand U5132 (N_5132,N_4751,N_4706);
nand U5133 (N_5133,N_4506,N_4642);
nor U5134 (N_5134,N_4802,N_4663);
nor U5135 (N_5135,N_4709,N_4753);
xor U5136 (N_5136,N_4838,N_4795);
nor U5137 (N_5137,N_4666,N_4550);
and U5138 (N_5138,N_4549,N_4577);
nand U5139 (N_5139,N_4847,N_4581);
nand U5140 (N_5140,N_4858,N_4569);
xor U5141 (N_5141,N_4514,N_4738);
nand U5142 (N_5142,N_4895,N_4986);
xnor U5143 (N_5143,N_4877,N_4707);
nand U5144 (N_5144,N_4712,N_4708);
xor U5145 (N_5145,N_4988,N_4598);
nand U5146 (N_5146,N_4629,N_4766);
nor U5147 (N_5147,N_4887,N_4944);
xor U5148 (N_5148,N_4530,N_4576);
nor U5149 (N_5149,N_4906,N_4505);
xnor U5150 (N_5150,N_4713,N_4929);
xnor U5151 (N_5151,N_4972,N_4993);
or U5152 (N_5152,N_4756,N_4897);
or U5153 (N_5153,N_4561,N_4789);
or U5154 (N_5154,N_4711,N_4624);
or U5155 (N_5155,N_4702,N_4967);
nor U5156 (N_5156,N_4656,N_4954);
nor U5157 (N_5157,N_4774,N_4813);
nor U5158 (N_5158,N_4579,N_4921);
or U5159 (N_5159,N_4959,N_4728);
or U5160 (N_5160,N_4934,N_4750);
nand U5161 (N_5161,N_4890,N_4855);
nand U5162 (N_5162,N_4994,N_4653);
nor U5163 (N_5163,N_4508,N_4705);
or U5164 (N_5164,N_4570,N_4835);
nor U5165 (N_5165,N_4962,N_4914);
and U5166 (N_5166,N_4540,N_4637);
xnor U5167 (N_5167,N_4770,N_4922);
nor U5168 (N_5168,N_4991,N_4960);
nor U5169 (N_5169,N_4927,N_4987);
or U5170 (N_5170,N_4814,N_4826);
nand U5171 (N_5171,N_4876,N_4729);
nor U5172 (N_5172,N_4853,N_4968);
or U5173 (N_5173,N_4773,N_4593);
or U5174 (N_5174,N_4727,N_4655);
xnor U5175 (N_5175,N_4546,N_4747);
nand U5176 (N_5176,N_4970,N_4580);
and U5177 (N_5177,N_4822,N_4829);
and U5178 (N_5178,N_4644,N_4528);
xnor U5179 (N_5179,N_4984,N_4591);
nor U5180 (N_5180,N_4596,N_4854);
nor U5181 (N_5181,N_4810,N_4664);
nand U5182 (N_5182,N_4627,N_4516);
xor U5183 (N_5183,N_4507,N_4519);
and U5184 (N_5184,N_4768,N_4824);
and U5185 (N_5185,N_4573,N_4928);
and U5186 (N_5186,N_4845,N_4809);
nand U5187 (N_5187,N_4509,N_4556);
nor U5188 (N_5188,N_4614,N_4551);
and U5189 (N_5189,N_4626,N_4885);
and U5190 (N_5190,N_4681,N_4930);
nor U5191 (N_5191,N_4502,N_4731);
nand U5192 (N_5192,N_4525,N_4503);
xor U5193 (N_5193,N_4837,N_4941);
or U5194 (N_5194,N_4552,N_4595);
or U5195 (N_5195,N_4677,N_4761);
nand U5196 (N_5196,N_4615,N_4875);
xnor U5197 (N_5197,N_4764,N_4804);
and U5198 (N_5198,N_4880,N_4903);
xor U5199 (N_5199,N_4981,N_4725);
xor U5200 (N_5200,N_4869,N_4832);
and U5201 (N_5201,N_4820,N_4523);
and U5202 (N_5202,N_4527,N_4721);
and U5203 (N_5203,N_4700,N_4965);
nand U5204 (N_5204,N_4649,N_4923);
or U5205 (N_5205,N_4638,N_4636);
or U5206 (N_5206,N_4586,N_4541);
xor U5207 (N_5207,N_4989,N_4676);
and U5208 (N_5208,N_4646,N_4823);
nor U5209 (N_5209,N_4612,N_4548);
nand U5210 (N_5210,N_4969,N_4775);
xor U5211 (N_5211,N_4990,N_4816);
or U5212 (N_5212,N_4735,N_4654);
nand U5213 (N_5213,N_4799,N_4781);
xor U5214 (N_5214,N_4896,N_4831);
or U5215 (N_5215,N_4639,N_4733);
and U5216 (N_5216,N_4739,N_4797);
nand U5217 (N_5217,N_4940,N_4918);
or U5218 (N_5218,N_4803,N_4878);
nand U5219 (N_5219,N_4585,N_4886);
nor U5220 (N_5220,N_4798,N_4974);
and U5221 (N_5221,N_4597,N_4522);
or U5222 (N_5222,N_4675,N_4690);
nand U5223 (N_5223,N_4513,N_4668);
nor U5224 (N_5224,N_4632,N_4849);
or U5225 (N_5225,N_4748,N_4952);
nor U5226 (N_5226,N_4512,N_4833);
and U5227 (N_5227,N_4609,N_4851);
or U5228 (N_5228,N_4948,N_4667);
xor U5229 (N_5229,N_4500,N_4571);
nor U5230 (N_5230,N_4791,N_4554);
nand U5231 (N_5231,N_4671,N_4543);
nand U5232 (N_5232,N_4983,N_4828);
nand U5233 (N_5233,N_4633,N_4889);
nand U5234 (N_5234,N_4565,N_4790);
or U5235 (N_5235,N_4846,N_4742);
nand U5236 (N_5236,N_4908,N_4603);
nor U5237 (N_5237,N_4779,N_4860);
and U5238 (N_5238,N_4698,N_4859);
nor U5239 (N_5239,N_4669,N_4801);
nor U5240 (N_5240,N_4643,N_4701);
xor U5241 (N_5241,N_4635,N_4807);
or U5242 (N_5242,N_4694,N_4544);
nand U5243 (N_5243,N_4817,N_4680);
xnor U5244 (N_5244,N_4501,N_4915);
nand U5245 (N_5245,N_4717,N_4794);
nand U5246 (N_5246,N_4547,N_4583);
xor U5247 (N_5247,N_4560,N_4589);
xor U5248 (N_5248,N_4631,N_4567);
nor U5249 (N_5249,N_4534,N_4563);
nand U5250 (N_5250,N_4814,N_4760);
or U5251 (N_5251,N_4895,N_4930);
nand U5252 (N_5252,N_4959,N_4622);
xor U5253 (N_5253,N_4507,N_4973);
nand U5254 (N_5254,N_4749,N_4622);
or U5255 (N_5255,N_4508,N_4971);
and U5256 (N_5256,N_4673,N_4515);
nor U5257 (N_5257,N_4593,N_4684);
xor U5258 (N_5258,N_4832,N_4911);
xnor U5259 (N_5259,N_4655,N_4654);
and U5260 (N_5260,N_4760,N_4995);
nor U5261 (N_5261,N_4968,N_4922);
and U5262 (N_5262,N_4751,N_4959);
nand U5263 (N_5263,N_4961,N_4759);
xnor U5264 (N_5264,N_4566,N_4765);
and U5265 (N_5265,N_4738,N_4753);
nand U5266 (N_5266,N_4720,N_4997);
and U5267 (N_5267,N_4591,N_4710);
and U5268 (N_5268,N_4599,N_4983);
or U5269 (N_5269,N_4639,N_4918);
nor U5270 (N_5270,N_4956,N_4780);
or U5271 (N_5271,N_4749,N_4799);
or U5272 (N_5272,N_4598,N_4597);
and U5273 (N_5273,N_4896,N_4910);
and U5274 (N_5274,N_4642,N_4609);
xor U5275 (N_5275,N_4587,N_4613);
and U5276 (N_5276,N_4611,N_4604);
or U5277 (N_5277,N_4763,N_4805);
nor U5278 (N_5278,N_4815,N_4899);
nor U5279 (N_5279,N_4961,N_4897);
and U5280 (N_5280,N_4581,N_4621);
nor U5281 (N_5281,N_4747,N_4870);
or U5282 (N_5282,N_4717,N_4964);
and U5283 (N_5283,N_4515,N_4670);
nand U5284 (N_5284,N_4663,N_4705);
xor U5285 (N_5285,N_4790,N_4795);
nor U5286 (N_5286,N_4569,N_4718);
nor U5287 (N_5287,N_4615,N_4669);
or U5288 (N_5288,N_4584,N_4780);
xnor U5289 (N_5289,N_4555,N_4559);
nand U5290 (N_5290,N_4687,N_4588);
and U5291 (N_5291,N_4845,N_4908);
or U5292 (N_5292,N_4817,N_4634);
nor U5293 (N_5293,N_4888,N_4645);
or U5294 (N_5294,N_4772,N_4815);
nor U5295 (N_5295,N_4876,N_4867);
or U5296 (N_5296,N_4630,N_4621);
xnor U5297 (N_5297,N_4665,N_4983);
nor U5298 (N_5298,N_4581,N_4901);
xor U5299 (N_5299,N_4812,N_4602);
nand U5300 (N_5300,N_4656,N_4817);
xnor U5301 (N_5301,N_4765,N_4769);
and U5302 (N_5302,N_4799,N_4816);
or U5303 (N_5303,N_4672,N_4872);
or U5304 (N_5304,N_4826,N_4528);
or U5305 (N_5305,N_4961,N_4842);
or U5306 (N_5306,N_4901,N_4856);
or U5307 (N_5307,N_4970,N_4588);
xnor U5308 (N_5308,N_4798,N_4582);
or U5309 (N_5309,N_4721,N_4800);
nand U5310 (N_5310,N_4941,N_4659);
and U5311 (N_5311,N_4595,N_4624);
nor U5312 (N_5312,N_4945,N_4543);
xnor U5313 (N_5313,N_4688,N_4791);
or U5314 (N_5314,N_4945,N_4856);
xor U5315 (N_5315,N_4772,N_4794);
or U5316 (N_5316,N_4854,N_4590);
and U5317 (N_5317,N_4736,N_4745);
nand U5318 (N_5318,N_4745,N_4766);
and U5319 (N_5319,N_4882,N_4756);
and U5320 (N_5320,N_4748,N_4997);
or U5321 (N_5321,N_4766,N_4566);
and U5322 (N_5322,N_4967,N_4857);
xor U5323 (N_5323,N_4979,N_4833);
nor U5324 (N_5324,N_4527,N_4995);
and U5325 (N_5325,N_4646,N_4589);
nor U5326 (N_5326,N_4674,N_4554);
xnor U5327 (N_5327,N_4838,N_4616);
or U5328 (N_5328,N_4679,N_4991);
and U5329 (N_5329,N_4961,N_4559);
xor U5330 (N_5330,N_4597,N_4574);
or U5331 (N_5331,N_4872,N_4893);
nor U5332 (N_5332,N_4502,N_4956);
nor U5333 (N_5333,N_4795,N_4837);
nor U5334 (N_5334,N_4962,N_4880);
xor U5335 (N_5335,N_4792,N_4750);
nor U5336 (N_5336,N_4699,N_4750);
and U5337 (N_5337,N_4656,N_4843);
and U5338 (N_5338,N_4735,N_4661);
nor U5339 (N_5339,N_4796,N_4833);
nor U5340 (N_5340,N_4842,N_4713);
or U5341 (N_5341,N_4880,N_4542);
and U5342 (N_5342,N_4645,N_4552);
and U5343 (N_5343,N_4811,N_4645);
xnor U5344 (N_5344,N_4661,N_4520);
or U5345 (N_5345,N_4874,N_4819);
xnor U5346 (N_5346,N_4796,N_4676);
xnor U5347 (N_5347,N_4876,N_4511);
nor U5348 (N_5348,N_4928,N_4980);
or U5349 (N_5349,N_4552,N_4548);
nor U5350 (N_5350,N_4776,N_4875);
nor U5351 (N_5351,N_4653,N_4593);
nand U5352 (N_5352,N_4930,N_4661);
xnor U5353 (N_5353,N_4909,N_4685);
or U5354 (N_5354,N_4739,N_4705);
xor U5355 (N_5355,N_4510,N_4889);
nor U5356 (N_5356,N_4901,N_4826);
nor U5357 (N_5357,N_4640,N_4961);
nand U5358 (N_5358,N_4744,N_4994);
nor U5359 (N_5359,N_4862,N_4825);
and U5360 (N_5360,N_4510,N_4681);
and U5361 (N_5361,N_4652,N_4875);
or U5362 (N_5362,N_4639,N_4824);
nor U5363 (N_5363,N_4909,N_4590);
xnor U5364 (N_5364,N_4846,N_4822);
xnor U5365 (N_5365,N_4659,N_4868);
nand U5366 (N_5366,N_4696,N_4629);
nand U5367 (N_5367,N_4641,N_4711);
nor U5368 (N_5368,N_4822,N_4852);
nand U5369 (N_5369,N_4995,N_4708);
nor U5370 (N_5370,N_4913,N_4892);
nor U5371 (N_5371,N_4725,N_4845);
and U5372 (N_5372,N_4582,N_4699);
nor U5373 (N_5373,N_4608,N_4681);
or U5374 (N_5374,N_4921,N_4818);
xnor U5375 (N_5375,N_4675,N_4599);
and U5376 (N_5376,N_4833,N_4867);
or U5377 (N_5377,N_4562,N_4589);
nor U5378 (N_5378,N_4539,N_4500);
nand U5379 (N_5379,N_4737,N_4940);
nand U5380 (N_5380,N_4972,N_4896);
or U5381 (N_5381,N_4553,N_4603);
and U5382 (N_5382,N_4968,N_4838);
or U5383 (N_5383,N_4534,N_4837);
and U5384 (N_5384,N_4554,N_4625);
and U5385 (N_5385,N_4993,N_4549);
or U5386 (N_5386,N_4612,N_4811);
or U5387 (N_5387,N_4964,N_4572);
nor U5388 (N_5388,N_4779,N_4839);
nand U5389 (N_5389,N_4628,N_4904);
nand U5390 (N_5390,N_4875,N_4893);
xnor U5391 (N_5391,N_4543,N_4617);
xor U5392 (N_5392,N_4805,N_4760);
nor U5393 (N_5393,N_4868,N_4858);
xor U5394 (N_5394,N_4742,N_4567);
xnor U5395 (N_5395,N_4852,N_4905);
and U5396 (N_5396,N_4659,N_4662);
and U5397 (N_5397,N_4673,N_4935);
xnor U5398 (N_5398,N_4901,N_4618);
xnor U5399 (N_5399,N_4899,N_4542);
nor U5400 (N_5400,N_4963,N_4679);
nand U5401 (N_5401,N_4586,N_4805);
and U5402 (N_5402,N_4867,N_4812);
or U5403 (N_5403,N_4911,N_4879);
nand U5404 (N_5404,N_4677,N_4869);
xnor U5405 (N_5405,N_4860,N_4512);
nor U5406 (N_5406,N_4677,N_4908);
xor U5407 (N_5407,N_4997,N_4765);
nor U5408 (N_5408,N_4990,N_4874);
and U5409 (N_5409,N_4523,N_4705);
or U5410 (N_5410,N_4803,N_4523);
and U5411 (N_5411,N_4624,N_4659);
nor U5412 (N_5412,N_4907,N_4585);
and U5413 (N_5413,N_4744,N_4503);
nand U5414 (N_5414,N_4781,N_4546);
or U5415 (N_5415,N_4524,N_4976);
nor U5416 (N_5416,N_4960,N_4674);
and U5417 (N_5417,N_4937,N_4510);
and U5418 (N_5418,N_4920,N_4696);
or U5419 (N_5419,N_4634,N_4626);
nor U5420 (N_5420,N_4972,N_4601);
nand U5421 (N_5421,N_4772,N_4952);
nand U5422 (N_5422,N_4838,N_4703);
xor U5423 (N_5423,N_4546,N_4671);
or U5424 (N_5424,N_4590,N_4690);
nor U5425 (N_5425,N_4759,N_4565);
or U5426 (N_5426,N_4858,N_4594);
or U5427 (N_5427,N_4846,N_4804);
and U5428 (N_5428,N_4852,N_4783);
and U5429 (N_5429,N_4522,N_4508);
nor U5430 (N_5430,N_4711,N_4650);
or U5431 (N_5431,N_4752,N_4713);
xor U5432 (N_5432,N_4649,N_4580);
and U5433 (N_5433,N_4572,N_4573);
xnor U5434 (N_5434,N_4816,N_4971);
or U5435 (N_5435,N_4563,N_4639);
and U5436 (N_5436,N_4795,N_4701);
or U5437 (N_5437,N_4867,N_4903);
nand U5438 (N_5438,N_4673,N_4788);
or U5439 (N_5439,N_4615,N_4811);
and U5440 (N_5440,N_4948,N_4577);
nor U5441 (N_5441,N_4748,N_4941);
and U5442 (N_5442,N_4529,N_4840);
nor U5443 (N_5443,N_4525,N_4545);
nor U5444 (N_5444,N_4693,N_4624);
nor U5445 (N_5445,N_4559,N_4861);
nor U5446 (N_5446,N_4574,N_4562);
nand U5447 (N_5447,N_4644,N_4537);
nand U5448 (N_5448,N_4625,N_4521);
or U5449 (N_5449,N_4861,N_4572);
xnor U5450 (N_5450,N_4663,N_4785);
xor U5451 (N_5451,N_4942,N_4944);
nor U5452 (N_5452,N_4679,N_4744);
and U5453 (N_5453,N_4555,N_4738);
or U5454 (N_5454,N_4941,N_4946);
and U5455 (N_5455,N_4779,N_4926);
and U5456 (N_5456,N_4993,N_4562);
xnor U5457 (N_5457,N_4725,N_4963);
xnor U5458 (N_5458,N_4709,N_4813);
xnor U5459 (N_5459,N_4614,N_4998);
and U5460 (N_5460,N_4565,N_4947);
or U5461 (N_5461,N_4547,N_4798);
and U5462 (N_5462,N_4980,N_4968);
nand U5463 (N_5463,N_4829,N_4972);
and U5464 (N_5464,N_4658,N_4560);
and U5465 (N_5465,N_4932,N_4697);
nand U5466 (N_5466,N_4581,N_4778);
or U5467 (N_5467,N_4844,N_4815);
xnor U5468 (N_5468,N_4889,N_4896);
nand U5469 (N_5469,N_4727,N_4915);
or U5470 (N_5470,N_4823,N_4508);
and U5471 (N_5471,N_4749,N_4659);
or U5472 (N_5472,N_4634,N_4527);
nand U5473 (N_5473,N_4598,N_4767);
and U5474 (N_5474,N_4627,N_4729);
xor U5475 (N_5475,N_4767,N_4634);
or U5476 (N_5476,N_4600,N_4928);
and U5477 (N_5477,N_4730,N_4786);
nor U5478 (N_5478,N_4542,N_4593);
or U5479 (N_5479,N_4887,N_4737);
or U5480 (N_5480,N_4698,N_4533);
nor U5481 (N_5481,N_4628,N_4754);
nand U5482 (N_5482,N_4831,N_4595);
and U5483 (N_5483,N_4844,N_4761);
or U5484 (N_5484,N_4526,N_4788);
and U5485 (N_5485,N_4687,N_4579);
and U5486 (N_5486,N_4713,N_4534);
nor U5487 (N_5487,N_4539,N_4824);
nor U5488 (N_5488,N_4634,N_4974);
or U5489 (N_5489,N_4766,N_4637);
nand U5490 (N_5490,N_4689,N_4654);
nand U5491 (N_5491,N_4833,N_4572);
or U5492 (N_5492,N_4604,N_4567);
and U5493 (N_5493,N_4999,N_4709);
or U5494 (N_5494,N_4665,N_4885);
or U5495 (N_5495,N_4807,N_4778);
nor U5496 (N_5496,N_4702,N_4782);
nand U5497 (N_5497,N_4935,N_4942);
and U5498 (N_5498,N_4671,N_4816);
and U5499 (N_5499,N_4772,N_4887);
xnor U5500 (N_5500,N_5130,N_5468);
or U5501 (N_5501,N_5185,N_5294);
and U5502 (N_5502,N_5056,N_5104);
xnor U5503 (N_5503,N_5298,N_5050);
or U5504 (N_5504,N_5193,N_5313);
or U5505 (N_5505,N_5043,N_5096);
xor U5506 (N_5506,N_5387,N_5004);
and U5507 (N_5507,N_5240,N_5138);
nand U5508 (N_5508,N_5071,N_5220);
xnor U5509 (N_5509,N_5396,N_5171);
nand U5510 (N_5510,N_5151,N_5196);
nor U5511 (N_5511,N_5353,N_5486);
xnor U5512 (N_5512,N_5101,N_5016);
nand U5513 (N_5513,N_5251,N_5238);
nand U5514 (N_5514,N_5014,N_5037);
and U5515 (N_5515,N_5273,N_5178);
and U5516 (N_5516,N_5122,N_5257);
nand U5517 (N_5517,N_5027,N_5350);
xor U5518 (N_5518,N_5323,N_5364);
xor U5519 (N_5519,N_5428,N_5328);
or U5520 (N_5520,N_5392,N_5301);
nor U5521 (N_5521,N_5186,N_5034);
nand U5522 (N_5522,N_5290,N_5357);
nand U5523 (N_5523,N_5054,N_5343);
xnor U5524 (N_5524,N_5095,N_5459);
and U5525 (N_5525,N_5379,N_5431);
xnor U5526 (N_5526,N_5441,N_5053);
or U5527 (N_5527,N_5136,N_5391);
and U5528 (N_5528,N_5417,N_5451);
xnor U5529 (N_5529,N_5013,N_5117);
or U5530 (N_5530,N_5134,N_5242);
xor U5531 (N_5531,N_5079,N_5354);
and U5532 (N_5532,N_5211,N_5411);
nor U5533 (N_5533,N_5112,N_5369);
or U5534 (N_5534,N_5331,N_5169);
and U5535 (N_5535,N_5320,N_5030);
xnor U5536 (N_5536,N_5135,N_5231);
and U5537 (N_5537,N_5336,N_5157);
xor U5538 (N_5538,N_5064,N_5176);
nand U5539 (N_5539,N_5165,N_5312);
nand U5540 (N_5540,N_5006,N_5254);
or U5541 (N_5541,N_5308,N_5052);
and U5542 (N_5542,N_5275,N_5339);
xor U5543 (N_5543,N_5198,N_5069);
or U5544 (N_5544,N_5348,N_5478);
or U5545 (N_5545,N_5229,N_5470);
and U5546 (N_5546,N_5084,N_5010);
xnor U5547 (N_5547,N_5103,N_5460);
and U5548 (N_5548,N_5111,N_5453);
and U5549 (N_5549,N_5435,N_5091);
nand U5550 (N_5550,N_5160,N_5397);
nor U5551 (N_5551,N_5184,N_5114);
nand U5552 (N_5552,N_5144,N_5373);
and U5553 (N_5553,N_5481,N_5132);
nand U5554 (N_5554,N_5370,N_5154);
xnor U5555 (N_5555,N_5085,N_5330);
or U5556 (N_5556,N_5081,N_5093);
and U5557 (N_5557,N_5035,N_5281);
nor U5558 (N_5558,N_5018,N_5306);
nor U5559 (N_5559,N_5271,N_5058);
or U5560 (N_5560,N_5378,N_5433);
nand U5561 (N_5561,N_5142,N_5246);
and U5562 (N_5562,N_5147,N_5244);
nand U5563 (N_5563,N_5127,N_5083);
and U5564 (N_5564,N_5248,N_5456);
or U5565 (N_5565,N_5405,N_5119);
nor U5566 (N_5566,N_5082,N_5066);
xnor U5567 (N_5567,N_5349,N_5159);
or U5568 (N_5568,N_5197,N_5466);
or U5569 (N_5569,N_5036,N_5444);
nand U5570 (N_5570,N_5356,N_5292);
nand U5571 (N_5571,N_5247,N_5001);
or U5572 (N_5572,N_5123,N_5252);
nand U5573 (N_5573,N_5048,N_5042);
or U5574 (N_5574,N_5299,N_5263);
or U5575 (N_5575,N_5146,N_5163);
nor U5576 (N_5576,N_5170,N_5126);
xor U5577 (N_5577,N_5094,N_5346);
or U5578 (N_5578,N_5311,N_5216);
nand U5579 (N_5579,N_5177,N_5166);
nand U5580 (N_5580,N_5497,N_5297);
or U5581 (N_5581,N_5187,N_5332);
xnor U5582 (N_5582,N_5499,N_5285);
or U5583 (N_5583,N_5394,N_5181);
xnor U5584 (N_5584,N_5333,N_5141);
nand U5585 (N_5585,N_5498,N_5194);
or U5586 (N_5586,N_5173,N_5237);
or U5587 (N_5587,N_5318,N_5334);
and U5588 (N_5588,N_5259,N_5145);
and U5589 (N_5589,N_5201,N_5125);
nand U5590 (N_5590,N_5372,N_5189);
xor U5591 (N_5591,N_5070,N_5152);
and U5592 (N_5592,N_5469,N_5310);
xnor U5593 (N_5593,N_5404,N_5492);
or U5594 (N_5594,N_5162,N_5324);
or U5595 (N_5595,N_5287,N_5218);
xor U5596 (N_5596,N_5366,N_5129);
xor U5597 (N_5597,N_5408,N_5009);
and U5598 (N_5598,N_5258,N_5245);
nand U5599 (N_5599,N_5026,N_5304);
and U5600 (N_5600,N_5222,N_5174);
xor U5601 (N_5601,N_5403,N_5462);
or U5602 (N_5602,N_5335,N_5401);
and U5603 (N_5603,N_5434,N_5179);
xor U5604 (N_5604,N_5046,N_5190);
nand U5605 (N_5605,N_5291,N_5494);
xor U5606 (N_5606,N_5293,N_5075);
and U5607 (N_5607,N_5137,N_5424);
or U5608 (N_5608,N_5063,N_5191);
and U5609 (N_5609,N_5284,N_5395);
xnor U5610 (N_5610,N_5358,N_5315);
xor U5611 (N_5611,N_5002,N_5041);
and U5612 (N_5612,N_5448,N_5068);
nor U5613 (N_5613,N_5383,N_5439);
nand U5614 (N_5614,N_5471,N_5180);
nand U5615 (N_5615,N_5051,N_5380);
and U5616 (N_5616,N_5419,N_5228);
and U5617 (N_5617,N_5376,N_5011);
nand U5618 (N_5618,N_5235,N_5020);
nor U5619 (N_5619,N_5450,N_5413);
nand U5620 (N_5620,N_5362,N_5164);
and U5621 (N_5621,N_5402,N_5426);
nand U5622 (N_5622,N_5022,N_5430);
and U5623 (N_5623,N_5115,N_5195);
or U5624 (N_5624,N_5361,N_5175);
nor U5625 (N_5625,N_5300,N_5233);
or U5626 (N_5626,N_5480,N_5414);
or U5627 (N_5627,N_5044,N_5032);
nor U5628 (N_5628,N_5266,N_5337);
nor U5629 (N_5629,N_5224,N_5283);
nor U5630 (N_5630,N_5386,N_5326);
xnor U5631 (N_5631,N_5289,N_5472);
and U5632 (N_5632,N_5409,N_5088);
and U5633 (N_5633,N_5024,N_5213);
or U5634 (N_5634,N_5340,N_5092);
or U5635 (N_5635,N_5208,N_5250);
or U5636 (N_5636,N_5427,N_5133);
nand U5637 (N_5637,N_5078,N_5467);
nand U5638 (N_5638,N_5317,N_5377);
nor U5639 (N_5639,N_5074,N_5038);
and U5640 (N_5640,N_5400,N_5031);
nor U5641 (N_5641,N_5168,N_5345);
or U5642 (N_5642,N_5440,N_5442);
or U5643 (N_5643,N_5230,N_5412);
and U5644 (N_5644,N_5342,N_5033);
nand U5645 (N_5645,N_5012,N_5329);
and U5646 (N_5646,N_5473,N_5067);
xor U5647 (N_5647,N_5295,N_5347);
nand U5648 (N_5648,N_5015,N_5118);
nand U5649 (N_5649,N_5143,N_5206);
nand U5650 (N_5650,N_5087,N_5028);
or U5651 (N_5651,N_5495,N_5445);
nand U5652 (N_5652,N_5458,N_5205);
and U5653 (N_5653,N_5019,N_5363);
xor U5654 (N_5654,N_5000,N_5124);
and U5655 (N_5655,N_5368,N_5319);
nor U5656 (N_5656,N_5393,N_5496);
nand U5657 (N_5657,N_5029,N_5105);
nor U5658 (N_5658,N_5107,N_5351);
and U5659 (N_5659,N_5077,N_5097);
or U5660 (N_5660,N_5385,N_5327);
nor U5661 (N_5661,N_5270,N_5243);
nand U5662 (N_5662,N_5389,N_5390);
or U5663 (N_5663,N_5479,N_5061);
nor U5664 (N_5664,N_5484,N_5371);
nor U5665 (N_5665,N_5374,N_5367);
and U5666 (N_5666,N_5416,N_5199);
xor U5667 (N_5667,N_5429,N_5399);
or U5668 (N_5668,N_5321,N_5073);
nor U5669 (N_5669,N_5260,N_5447);
nor U5670 (N_5670,N_5485,N_5446);
or U5671 (N_5671,N_5388,N_5454);
xnor U5672 (N_5672,N_5025,N_5214);
xnor U5673 (N_5673,N_5482,N_5307);
nand U5674 (N_5674,N_5491,N_5221);
xnor U5675 (N_5675,N_5155,N_5261);
or U5676 (N_5676,N_5161,N_5226);
nor U5677 (N_5677,N_5204,N_5352);
xor U5678 (N_5678,N_5065,N_5277);
nor U5679 (N_5679,N_5282,N_5463);
xor U5680 (N_5680,N_5080,N_5200);
nand U5681 (N_5681,N_5443,N_5128);
or U5682 (N_5682,N_5272,N_5420);
xnor U5683 (N_5683,N_5382,N_5172);
and U5684 (N_5684,N_5149,N_5457);
nor U5685 (N_5685,N_5375,N_5212);
nor U5686 (N_5686,N_5089,N_5415);
nor U5687 (N_5687,N_5007,N_5288);
nand U5688 (N_5688,N_5269,N_5278);
nand U5689 (N_5689,N_5274,N_5265);
and U5690 (N_5690,N_5359,N_5120);
nand U5691 (N_5691,N_5072,N_5102);
or U5692 (N_5692,N_5234,N_5236);
xnor U5693 (N_5693,N_5483,N_5465);
xor U5694 (N_5694,N_5438,N_5316);
xnor U5695 (N_5695,N_5188,N_5182);
xnor U5696 (N_5696,N_5215,N_5207);
nor U5697 (N_5697,N_5150,N_5076);
xnor U5698 (N_5698,N_5021,N_5422);
nor U5699 (N_5699,N_5309,N_5202);
nand U5700 (N_5700,N_5280,N_5449);
and U5701 (N_5701,N_5057,N_5455);
or U5702 (N_5702,N_5437,N_5488);
xor U5703 (N_5703,N_5086,N_5108);
nand U5704 (N_5704,N_5062,N_5060);
xor U5705 (N_5705,N_5003,N_5217);
or U5706 (N_5706,N_5140,N_5410);
nor U5707 (N_5707,N_5249,N_5055);
nand U5708 (N_5708,N_5475,N_5477);
or U5709 (N_5709,N_5338,N_5279);
or U5710 (N_5710,N_5156,N_5148);
nand U5711 (N_5711,N_5039,N_5268);
xnor U5712 (N_5712,N_5232,N_5109);
and U5713 (N_5713,N_5464,N_5227);
nand U5714 (N_5714,N_5253,N_5131);
and U5715 (N_5715,N_5017,N_5203);
or U5716 (N_5716,N_5099,N_5487);
xor U5717 (N_5717,N_5365,N_5040);
or U5718 (N_5718,N_5407,N_5239);
nand U5719 (N_5719,N_5059,N_5423);
and U5720 (N_5720,N_5241,N_5425);
xnor U5721 (N_5721,N_5139,N_5286);
xnor U5722 (N_5722,N_5406,N_5432);
nor U5723 (N_5723,N_5106,N_5113);
xnor U5724 (N_5724,N_5267,N_5045);
xnor U5725 (N_5725,N_5489,N_5047);
xnor U5726 (N_5726,N_5322,N_5219);
nor U5727 (N_5727,N_5305,N_5116);
xnor U5728 (N_5728,N_5476,N_5344);
or U5729 (N_5729,N_5223,N_5005);
nand U5730 (N_5730,N_5167,N_5262);
or U5731 (N_5731,N_5303,N_5153);
xor U5732 (N_5732,N_5210,N_5255);
nor U5733 (N_5733,N_5452,N_5341);
nand U5734 (N_5734,N_5121,N_5023);
xor U5735 (N_5735,N_5225,N_5256);
and U5736 (N_5736,N_5314,N_5110);
nor U5737 (N_5737,N_5381,N_5355);
or U5738 (N_5738,N_5325,N_5100);
nand U5739 (N_5739,N_5192,N_5209);
xnor U5740 (N_5740,N_5008,N_5302);
and U5741 (N_5741,N_5360,N_5474);
or U5742 (N_5742,N_5098,N_5398);
nor U5743 (N_5743,N_5436,N_5296);
nand U5744 (N_5744,N_5461,N_5384);
and U5745 (N_5745,N_5493,N_5418);
nor U5746 (N_5746,N_5090,N_5158);
or U5747 (N_5747,N_5276,N_5490);
and U5748 (N_5748,N_5264,N_5049);
xnor U5749 (N_5749,N_5421,N_5183);
or U5750 (N_5750,N_5313,N_5278);
nor U5751 (N_5751,N_5068,N_5006);
nand U5752 (N_5752,N_5207,N_5088);
nor U5753 (N_5753,N_5402,N_5112);
and U5754 (N_5754,N_5292,N_5249);
xor U5755 (N_5755,N_5167,N_5486);
nor U5756 (N_5756,N_5474,N_5198);
or U5757 (N_5757,N_5161,N_5337);
nor U5758 (N_5758,N_5110,N_5366);
or U5759 (N_5759,N_5171,N_5051);
nor U5760 (N_5760,N_5011,N_5488);
nand U5761 (N_5761,N_5295,N_5076);
nor U5762 (N_5762,N_5180,N_5108);
or U5763 (N_5763,N_5341,N_5162);
or U5764 (N_5764,N_5377,N_5174);
xor U5765 (N_5765,N_5010,N_5093);
and U5766 (N_5766,N_5216,N_5385);
nand U5767 (N_5767,N_5310,N_5163);
or U5768 (N_5768,N_5249,N_5032);
nor U5769 (N_5769,N_5198,N_5353);
xor U5770 (N_5770,N_5272,N_5496);
xnor U5771 (N_5771,N_5266,N_5411);
and U5772 (N_5772,N_5069,N_5420);
nand U5773 (N_5773,N_5400,N_5425);
or U5774 (N_5774,N_5305,N_5209);
nor U5775 (N_5775,N_5051,N_5033);
nor U5776 (N_5776,N_5118,N_5177);
nor U5777 (N_5777,N_5008,N_5499);
and U5778 (N_5778,N_5335,N_5348);
or U5779 (N_5779,N_5496,N_5498);
or U5780 (N_5780,N_5340,N_5095);
nor U5781 (N_5781,N_5441,N_5133);
or U5782 (N_5782,N_5172,N_5063);
nor U5783 (N_5783,N_5481,N_5393);
nand U5784 (N_5784,N_5201,N_5207);
nor U5785 (N_5785,N_5142,N_5054);
xor U5786 (N_5786,N_5049,N_5461);
and U5787 (N_5787,N_5032,N_5390);
or U5788 (N_5788,N_5128,N_5221);
nor U5789 (N_5789,N_5105,N_5301);
or U5790 (N_5790,N_5451,N_5022);
nor U5791 (N_5791,N_5195,N_5107);
nand U5792 (N_5792,N_5119,N_5394);
xor U5793 (N_5793,N_5118,N_5492);
and U5794 (N_5794,N_5295,N_5226);
and U5795 (N_5795,N_5435,N_5170);
nand U5796 (N_5796,N_5205,N_5388);
xnor U5797 (N_5797,N_5475,N_5014);
and U5798 (N_5798,N_5006,N_5420);
and U5799 (N_5799,N_5495,N_5033);
xor U5800 (N_5800,N_5251,N_5282);
or U5801 (N_5801,N_5060,N_5493);
xor U5802 (N_5802,N_5124,N_5244);
xor U5803 (N_5803,N_5124,N_5370);
xor U5804 (N_5804,N_5140,N_5034);
and U5805 (N_5805,N_5272,N_5491);
and U5806 (N_5806,N_5269,N_5190);
or U5807 (N_5807,N_5220,N_5078);
nor U5808 (N_5808,N_5377,N_5473);
or U5809 (N_5809,N_5306,N_5285);
nand U5810 (N_5810,N_5171,N_5473);
and U5811 (N_5811,N_5286,N_5199);
nand U5812 (N_5812,N_5348,N_5129);
nand U5813 (N_5813,N_5230,N_5241);
or U5814 (N_5814,N_5015,N_5386);
nor U5815 (N_5815,N_5433,N_5207);
or U5816 (N_5816,N_5272,N_5220);
nor U5817 (N_5817,N_5015,N_5194);
xor U5818 (N_5818,N_5211,N_5298);
and U5819 (N_5819,N_5133,N_5067);
xor U5820 (N_5820,N_5015,N_5321);
xor U5821 (N_5821,N_5207,N_5365);
xnor U5822 (N_5822,N_5387,N_5051);
xnor U5823 (N_5823,N_5100,N_5146);
nor U5824 (N_5824,N_5376,N_5196);
nand U5825 (N_5825,N_5350,N_5176);
xor U5826 (N_5826,N_5348,N_5117);
and U5827 (N_5827,N_5009,N_5487);
nand U5828 (N_5828,N_5013,N_5159);
and U5829 (N_5829,N_5486,N_5118);
or U5830 (N_5830,N_5402,N_5147);
and U5831 (N_5831,N_5119,N_5092);
nor U5832 (N_5832,N_5053,N_5083);
and U5833 (N_5833,N_5053,N_5188);
nand U5834 (N_5834,N_5462,N_5133);
or U5835 (N_5835,N_5484,N_5006);
or U5836 (N_5836,N_5435,N_5128);
nand U5837 (N_5837,N_5397,N_5132);
nor U5838 (N_5838,N_5009,N_5363);
or U5839 (N_5839,N_5490,N_5314);
nand U5840 (N_5840,N_5031,N_5387);
or U5841 (N_5841,N_5290,N_5141);
and U5842 (N_5842,N_5353,N_5418);
and U5843 (N_5843,N_5350,N_5144);
and U5844 (N_5844,N_5268,N_5163);
nand U5845 (N_5845,N_5211,N_5451);
or U5846 (N_5846,N_5410,N_5083);
and U5847 (N_5847,N_5325,N_5228);
xnor U5848 (N_5848,N_5050,N_5278);
or U5849 (N_5849,N_5093,N_5275);
or U5850 (N_5850,N_5368,N_5119);
xnor U5851 (N_5851,N_5487,N_5485);
and U5852 (N_5852,N_5440,N_5378);
xnor U5853 (N_5853,N_5032,N_5472);
nand U5854 (N_5854,N_5302,N_5373);
nor U5855 (N_5855,N_5250,N_5004);
or U5856 (N_5856,N_5233,N_5262);
or U5857 (N_5857,N_5154,N_5009);
xnor U5858 (N_5858,N_5321,N_5183);
nor U5859 (N_5859,N_5037,N_5296);
nor U5860 (N_5860,N_5372,N_5176);
xor U5861 (N_5861,N_5024,N_5460);
nand U5862 (N_5862,N_5209,N_5299);
nor U5863 (N_5863,N_5364,N_5199);
nor U5864 (N_5864,N_5268,N_5145);
or U5865 (N_5865,N_5407,N_5203);
xor U5866 (N_5866,N_5493,N_5323);
nand U5867 (N_5867,N_5156,N_5093);
xor U5868 (N_5868,N_5000,N_5476);
xnor U5869 (N_5869,N_5033,N_5446);
xnor U5870 (N_5870,N_5073,N_5178);
nand U5871 (N_5871,N_5357,N_5064);
nand U5872 (N_5872,N_5239,N_5364);
nand U5873 (N_5873,N_5028,N_5287);
and U5874 (N_5874,N_5453,N_5465);
nand U5875 (N_5875,N_5117,N_5293);
or U5876 (N_5876,N_5023,N_5210);
and U5877 (N_5877,N_5010,N_5194);
nor U5878 (N_5878,N_5125,N_5164);
xor U5879 (N_5879,N_5011,N_5205);
and U5880 (N_5880,N_5393,N_5273);
xnor U5881 (N_5881,N_5115,N_5231);
and U5882 (N_5882,N_5121,N_5353);
or U5883 (N_5883,N_5436,N_5161);
xnor U5884 (N_5884,N_5254,N_5180);
xnor U5885 (N_5885,N_5126,N_5365);
xor U5886 (N_5886,N_5079,N_5271);
or U5887 (N_5887,N_5226,N_5165);
nand U5888 (N_5888,N_5168,N_5330);
or U5889 (N_5889,N_5285,N_5391);
nand U5890 (N_5890,N_5094,N_5224);
or U5891 (N_5891,N_5473,N_5092);
or U5892 (N_5892,N_5348,N_5033);
and U5893 (N_5893,N_5424,N_5491);
xnor U5894 (N_5894,N_5323,N_5467);
or U5895 (N_5895,N_5440,N_5062);
xor U5896 (N_5896,N_5146,N_5433);
nand U5897 (N_5897,N_5146,N_5446);
and U5898 (N_5898,N_5115,N_5142);
nand U5899 (N_5899,N_5466,N_5078);
and U5900 (N_5900,N_5298,N_5046);
or U5901 (N_5901,N_5289,N_5115);
or U5902 (N_5902,N_5352,N_5018);
nand U5903 (N_5903,N_5487,N_5391);
nand U5904 (N_5904,N_5062,N_5068);
nor U5905 (N_5905,N_5393,N_5317);
or U5906 (N_5906,N_5064,N_5277);
nor U5907 (N_5907,N_5215,N_5415);
or U5908 (N_5908,N_5192,N_5305);
and U5909 (N_5909,N_5404,N_5222);
and U5910 (N_5910,N_5150,N_5027);
or U5911 (N_5911,N_5401,N_5083);
and U5912 (N_5912,N_5381,N_5275);
nand U5913 (N_5913,N_5138,N_5200);
nor U5914 (N_5914,N_5065,N_5221);
nor U5915 (N_5915,N_5360,N_5045);
and U5916 (N_5916,N_5288,N_5185);
nand U5917 (N_5917,N_5440,N_5476);
or U5918 (N_5918,N_5435,N_5341);
xnor U5919 (N_5919,N_5459,N_5398);
nand U5920 (N_5920,N_5456,N_5075);
and U5921 (N_5921,N_5415,N_5220);
xnor U5922 (N_5922,N_5090,N_5199);
and U5923 (N_5923,N_5337,N_5273);
xnor U5924 (N_5924,N_5454,N_5475);
or U5925 (N_5925,N_5449,N_5001);
nand U5926 (N_5926,N_5290,N_5356);
nor U5927 (N_5927,N_5154,N_5016);
nor U5928 (N_5928,N_5212,N_5410);
and U5929 (N_5929,N_5389,N_5125);
xnor U5930 (N_5930,N_5249,N_5366);
or U5931 (N_5931,N_5208,N_5066);
nor U5932 (N_5932,N_5291,N_5480);
nor U5933 (N_5933,N_5063,N_5468);
or U5934 (N_5934,N_5149,N_5285);
nor U5935 (N_5935,N_5164,N_5291);
and U5936 (N_5936,N_5098,N_5478);
xnor U5937 (N_5937,N_5339,N_5350);
nand U5938 (N_5938,N_5148,N_5022);
nor U5939 (N_5939,N_5494,N_5194);
nor U5940 (N_5940,N_5332,N_5390);
or U5941 (N_5941,N_5408,N_5065);
nand U5942 (N_5942,N_5158,N_5157);
nor U5943 (N_5943,N_5006,N_5424);
nor U5944 (N_5944,N_5105,N_5434);
nor U5945 (N_5945,N_5130,N_5049);
nor U5946 (N_5946,N_5455,N_5287);
nand U5947 (N_5947,N_5172,N_5441);
and U5948 (N_5948,N_5042,N_5019);
xnor U5949 (N_5949,N_5117,N_5447);
or U5950 (N_5950,N_5440,N_5219);
xor U5951 (N_5951,N_5092,N_5126);
and U5952 (N_5952,N_5285,N_5400);
xnor U5953 (N_5953,N_5284,N_5477);
and U5954 (N_5954,N_5410,N_5077);
nor U5955 (N_5955,N_5308,N_5009);
nor U5956 (N_5956,N_5104,N_5377);
nand U5957 (N_5957,N_5325,N_5448);
and U5958 (N_5958,N_5332,N_5475);
nor U5959 (N_5959,N_5335,N_5442);
and U5960 (N_5960,N_5015,N_5008);
nand U5961 (N_5961,N_5166,N_5120);
and U5962 (N_5962,N_5149,N_5121);
xnor U5963 (N_5963,N_5285,N_5398);
nand U5964 (N_5964,N_5423,N_5078);
and U5965 (N_5965,N_5273,N_5216);
nand U5966 (N_5966,N_5073,N_5302);
nor U5967 (N_5967,N_5190,N_5002);
xnor U5968 (N_5968,N_5320,N_5280);
and U5969 (N_5969,N_5210,N_5357);
xor U5970 (N_5970,N_5146,N_5357);
or U5971 (N_5971,N_5037,N_5196);
nor U5972 (N_5972,N_5045,N_5320);
or U5973 (N_5973,N_5485,N_5080);
and U5974 (N_5974,N_5439,N_5278);
nor U5975 (N_5975,N_5452,N_5474);
or U5976 (N_5976,N_5049,N_5141);
nor U5977 (N_5977,N_5365,N_5255);
xnor U5978 (N_5978,N_5304,N_5456);
nor U5979 (N_5979,N_5315,N_5294);
xnor U5980 (N_5980,N_5410,N_5390);
nor U5981 (N_5981,N_5142,N_5336);
nand U5982 (N_5982,N_5308,N_5344);
xnor U5983 (N_5983,N_5175,N_5258);
nand U5984 (N_5984,N_5345,N_5084);
and U5985 (N_5985,N_5414,N_5470);
or U5986 (N_5986,N_5080,N_5015);
and U5987 (N_5987,N_5025,N_5063);
and U5988 (N_5988,N_5307,N_5479);
and U5989 (N_5989,N_5156,N_5291);
xor U5990 (N_5990,N_5381,N_5298);
nor U5991 (N_5991,N_5271,N_5484);
and U5992 (N_5992,N_5156,N_5281);
nor U5993 (N_5993,N_5084,N_5382);
nor U5994 (N_5994,N_5342,N_5233);
nor U5995 (N_5995,N_5201,N_5457);
xnor U5996 (N_5996,N_5325,N_5279);
nor U5997 (N_5997,N_5302,N_5415);
nand U5998 (N_5998,N_5113,N_5303);
nand U5999 (N_5999,N_5447,N_5456);
xnor U6000 (N_6000,N_5996,N_5902);
nor U6001 (N_6001,N_5565,N_5643);
nand U6002 (N_6002,N_5557,N_5761);
nor U6003 (N_6003,N_5857,N_5630);
or U6004 (N_6004,N_5701,N_5707);
nand U6005 (N_6005,N_5552,N_5845);
nand U6006 (N_6006,N_5659,N_5534);
or U6007 (N_6007,N_5673,N_5698);
xnor U6008 (N_6008,N_5619,N_5992);
xor U6009 (N_6009,N_5684,N_5522);
or U6010 (N_6010,N_5878,N_5514);
or U6011 (N_6011,N_5589,N_5638);
nand U6012 (N_6012,N_5733,N_5752);
and U6013 (N_6013,N_5766,N_5590);
nor U6014 (N_6014,N_5769,N_5743);
nand U6015 (N_6015,N_5583,N_5646);
and U6016 (N_6016,N_5689,N_5692);
and U6017 (N_6017,N_5874,N_5645);
and U6018 (N_6018,N_5838,N_5687);
xnor U6019 (N_6019,N_5528,N_5779);
nor U6020 (N_6020,N_5603,N_5559);
nor U6021 (N_6021,N_5828,N_5988);
xnor U6022 (N_6022,N_5745,N_5994);
or U6023 (N_6023,N_5516,N_5520);
nor U6024 (N_6024,N_5765,N_5946);
nor U6025 (N_6025,N_5637,N_5688);
xnor U6026 (N_6026,N_5958,N_5921);
or U6027 (N_6027,N_5605,N_5502);
or U6028 (N_6028,N_5535,N_5933);
xor U6029 (N_6029,N_5968,N_5756);
xor U6030 (N_6030,N_5817,N_5686);
nand U6031 (N_6031,N_5714,N_5571);
nand U6032 (N_6032,N_5651,N_5883);
nor U6033 (N_6033,N_5711,N_5639);
nand U6034 (N_6034,N_5831,N_5539);
or U6035 (N_6035,N_5863,N_5697);
or U6036 (N_6036,N_5950,N_5771);
xnor U6037 (N_6037,N_5533,N_5772);
and U6038 (N_6038,N_5678,N_5650);
and U6039 (N_6039,N_5691,N_5724);
nand U6040 (N_6040,N_5912,N_5781);
xor U6041 (N_6041,N_5987,N_5696);
and U6042 (N_6042,N_5908,N_5703);
nand U6043 (N_6043,N_5901,N_5844);
nor U6044 (N_6044,N_5961,N_5775);
nand U6045 (N_6045,N_5903,N_5825);
nor U6046 (N_6046,N_5575,N_5892);
or U6047 (N_6047,N_5753,N_5602);
xor U6048 (N_6048,N_5975,N_5983);
xnor U6049 (N_6049,N_5521,N_5974);
nand U6050 (N_6050,N_5882,N_5768);
and U6051 (N_6051,N_5633,N_5869);
and U6052 (N_6052,N_5661,N_5670);
or U6053 (N_6053,N_5674,N_5702);
nand U6054 (N_6054,N_5508,N_5699);
nand U6055 (N_6055,N_5834,N_5896);
nor U6056 (N_6056,N_5525,N_5647);
nand U6057 (N_6057,N_5764,N_5635);
xor U6058 (N_6058,N_5770,N_5550);
nor U6059 (N_6059,N_5695,N_5666);
nor U6060 (N_6060,N_5739,N_5510);
xor U6061 (N_6061,N_5564,N_5949);
nand U6062 (N_6062,N_5814,N_5986);
xnor U6063 (N_6063,N_5862,N_5569);
xor U6064 (N_6064,N_5748,N_5945);
nor U6065 (N_6065,N_5805,N_5801);
and U6066 (N_6066,N_5601,N_5663);
xor U6067 (N_6067,N_5894,N_5504);
xor U6068 (N_6068,N_5736,N_5860);
xor U6069 (N_6069,N_5581,N_5540);
xnor U6070 (N_6070,N_5624,N_5578);
nand U6071 (N_6071,N_5920,N_5759);
nor U6072 (N_6072,N_5959,N_5623);
and U6073 (N_6073,N_5917,N_5873);
nor U6074 (N_6074,N_5893,N_5880);
nor U6075 (N_6075,N_5820,N_5685);
and U6076 (N_6076,N_5962,N_5890);
or U6077 (N_6077,N_5997,N_5829);
and U6078 (N_6078,N_5762,N_5792);
and U6079 (N_6079,N_5970,N_5784);
nor U6080 (N_6080,N_5807,N_5795);
nand U6081 (N_6081,N_5816,N_5984);
nand U6082 (N_6082,N_5856,N_5990);
nor U6083 (N_6083,N_5708,N_5927);
and U6084 (N_6084,N_5910,N_5727);
nand U6085 (N_6085,N_5938,N_5562);
or U6086 (N_6086,N_5730,N_5806);
nand U6087 (N_6087,N_5723,N_5568);
nand U6088 (N_6088,N_5563,N_5715);
nor U6089 (N_6089,N_5636,N_5821);
xnor U6090 (N_6090,N_5813,N_5802);
xnor U6091 (N_6091,N_5812,N_5907);
xnor U6092 (N_6092,N_5751,N_5660);
xor U6093 (N_6093,N_5536,N_5631);
or U6094 (N_6094,N_5529,N_5725);
xnor U6095 (N_6095,N_5717,N_5995);
xor U6096 (N_6096,N_5587,N_5704);
or U6097 (N_6097,N_5613,N_5665);
or U6098 (N_6098,N_5930,N_5774);
or U6099 (N_6099,N_5669,N_5788);
nor U6100 (N_6100,N_5610,N_5577);
and U6101 (N_6101,N_5981,N_5541);
and U6102 (N_6102,N_5729,N_5767);
xnor U6103 (N_6103,N_5754,N_5848);
or U6104 (N_6104,N_5738,N_5554);
nand U6105 (N_6105,N_5763,N_5957);
or U6106 (N_6106,N_5586,N_5721);
or U6107 (N_6107,N_5573,N_5998);
or U6108 (N_6108,N_5544,N_5747);
xor U6109 (N_6109,N_5681,N_5700);
and U6110 (N_6110,N_5888,N_5582);
xnor U6111 (N_6111,N_5800,N_5822);
nor U6112 (N_6112,N_5913,N_5694);
or U6113 (N_6113,N_5966,N_5566);
nor U6114 (N_6114,N_5750,N_5895);
nand U6115 (N_6115,N_5668,N_5855);
or U6116 (N_6116,N_5606,N_5597);
and U6117 (N_6117,N_5979,N_5936);
nand U6118 (N_6118,N_5524,N_5911);
nand U6119 (N_6119,N_5517,N_5918);
or U6120 (N_6120,N_5940,N_5942);
xor U6121 (N_6121,N_5627,N_5909);
or U6122 (N_6122,N_5955,N_5532);
and U6123 (N_6123,N_5899,N_5889);
or U6124 (N_6124,N_5654,N_5712);
nor U6125 (N_6125,N_5853,N_5652);
xor U6126 (N_6126,N_5755,N_5876);
nand U6127 (N_6127,N_5783,N_5680);
nand U6128 (N_6128,N_5791,N_5655);
xnor U6129 (N_6129,N_5512,N_5594);
nor U6130 (N_6130,N_5985,N_5591);
nor U6131 (N_6131,N_5953,N_5891);
and U6132 (N_6132,N_5870,N_5518);
xor U6133 (N_6133,N_5972,N_5809);
nor U6134 (N_6134,N_5549,N_5648);
nor U6135 (N_6135,N_5509,N_5746);
nor U6136 (N_6136,N_5600,N_5794);
xor U6137 (N_6137,N_5886,N_5667);
nand U6138 (N_6138,N_5914,N_5790);
nand U6139 (N_6139,N_5599,N_5991);
and U6140 (N_6140,N_5542,N_5948);
nand U6141 (N_6141,N_5861,N_5887);
nor U6142 (N_6142,N_5789,N_5851);
or U6143 (N_6143,N_5963,N_5506);
or U6144 (N_6144,N_5737,N_5951);
and U6145 (N_6145,N_5758,N_5622);
xnor U6146 (N_6146,N_5875,N_5999);
nor U6147 (N_6147,N_5644,N_5931);
nor U6148 (N_6148,N_5634,N_5713);
and U6149 (N_6149,N_5798,N_5682);
xor U6150 (N_6150,N_5881,N_5960);
xnor U6151 (N_6151,N_5584,N_5993);
and U6152 (N_6152,N_5925,N_5824);
xnor U6153 (N_6153,N_5941,N_5973);
or U6154 (N_6154,N_5935,N_5572);
or U6155 (N_6155,N_5830,N_5937);
or U6156 (N_6156,N_5980,N_5850);
or U6157 (N_6157,N_5579,N_5731);
or U6158 (N_6158,N_5604,N_5641);
nand U6159 (N_6159,N_5977,N_5726);
and U6160 (N_6160,N_5864,N_5629);
and U6161 (N_6161,N_5580,N_5773);
or U6162 (N_6162,N_5932,N_5956);
nor U6163 (N_6163,N_5511,N_5916);
and U6164 (N_6164,N_5978,N_5501);
and U6165 (N_6165,N_5574,N_5615);
nand U6166 (N_6166,N_5849,N_5675);
xor U6167 (N_6167,N_5939,N_5560);
nor U6168 (N_6168,N_5526,N_5679);
and U6169 (N_6169,N_5545,N_5934);
and U6170 (N_6170,N_5546,N_5519);
or U6171 (N_6171,N_5561,N_5760);
or U6172 (N_6172,N_5553,N_5804);
nor U6173 (N_6173,N_5785,N_5811);
nor U6174 (N_6174,N_5926,N_5662);
nand U6175 (N_6175,N_5922,N_5558);
nor U6176 (N_6176,N_5915,N_5796);
nand U6177 (N_6177,N_5867,N_5719);
xnor U6178 (N_6178,N_5858,N_5841);
xor U6179 (N_6179,N_5866,N_5823);
or U6180 (N_6180,N_5551,N_5879);
nor U6181 (N_6181,N_5943,N_5744);
nor U6182 (N_6182,N_5632,N_5954);
and U6183 (N_6183,N_5884,N_5705);
xnor U6184 (N_6184,N_5843,N_5778);
nor U6185 (N_6185,N_5819,N_5657);
or U6186 (N_6186,N_5854,N_5500);
and U6187 (N_6187,N_5810,N_5836);
nor U6188 (N_6188,N_5906,N_5904);
or U6189 (N_6189,N_5923,N_5971);
xnor U6190 (N_6190,N_5982,N_5722);
xor U6191 (N_6191,N_5608,N_5897);
or U6192 (N_6192,N_5656,N_5965);
and U6193 (N_6193,N_5618,N_5515);
or U6194 (N_6194,N_5852,N_5538);
nor U6195 (N_6195,N_5842,N_5596);
nand U6196 (N_6196,N_5693,N_5642);
xor U6197 (N_6197,N_5531,N_5826);
or U6198 (N_6198,N_5924,N_5543);
nor U6199 (N_6199,N_5640,N_5588);
nor U6200 (N_6200,N_5537,N_5570);
or U6201 (N_6201,N_5846,N_5944);
or U6202 (N_6202,N_5720,N_5782);
nor U6203 (N_6203,N_5793,N_5740);
or U6204 (N_6204,N_5620,N_5612);
xnor U6205 (N_6205,N_5840,N_5947);
or U6206 (N_6206,N_5653,N_5555);
nor U6207 (N_6207,N_5609,N_5626);
or U6208 (N_6208,N_5732,N_5690);
and U6209 (N_6209,N_5595,N_5611);
nand U6210 (N_6210,N_5742,N_5585);
or U6211 (N_6211,N_5776,N_5616);
nand U6212 (N_6212,N_5503,N_5929);
and U6213 (N_6213,N_5706,N_5787);
nor U6214 (N_6214,N_5989,N_5530);
nor U6215 (N_6215,N_5523,N_5847);
nand U6216 (N_6216,N_5777,N_5741);
xnor U6217 (N_6217,N_5839,N_5658);
nor U6218 (N_6218,N_5928,N_5718);
and U6219 (N_6219,N_5786,N_5919);
and U6220 (N_6220,N_5803,N_5877);
nand U6221 (N_6221,N_5598,N_5976);
and U6222 (N_6222,N_5513,N_5709);
nand U6223 (N_6223,N_5734,N_5617);
xnor U6224 (N_6224,N_5799,N_5757);
nand U6225 (N_6225,N_5507,N_5818);
xnor U6226 (N_6226,N_5556,N_5676);
nor U6227 (N_6227,N_5710,N_5749);
or U6228 (N_6228,N_5835,N_5865);
xor U6229 (N_6229,N_5905,N_5716);
and U6230 (N_6230,N_5872,N_5885);
nand U6231 (N_6231,N_5859,N_5898);
nand U6232 (N_6232,N_5621,N_5683);
nand U6233 (N_6233,N_5628,N_5548);
xnor U6234 (N_6234,N_5728,N_5827);
nand U6235 (N_6235,N_5625,N_5567);
nor U6236 (N_6236,N_5505,N_5833);
nand U6237 (N_6237,N_5607,N_5547);
nor U6238 (N_6238,N_5592,N_5969);
xnor U6239 (N_6239,N_5780,N_5964);
or U6240 (N_6240,N_5815,N_5871);
nor U6241 (N_6241,N_5593,N_5868);
or U6242 (N_6242,N_5576,N_5677);
xor U6243 (N_6243,N_5952,N_5664);
nand U6244 (N_6244,N_5672,N_5671);
xnor U6245 (N_6245,N_5797,N_5527);
nor U6246 (N_6246,N_5735,N_5614);
or U6247 (N_6247,N_5967,N_5808);
nand U6248 (N_6248,N_5837,N_5832);
nand U6249 (N_6249,N_5649,N_5900);
xnor U6250 (N_6250,N_5989,N_5529);
or U6251 (N_6251,N_5606,N_5594);
or U6252 (N_6252,N_5640,N_5530);
nand U6253 (N_6253,N_5979,N_5704);
xor U6254 (N_6254,N_5787,N_5990);
nand U6255 (N_6255,N_5519,N_5677);
nor U6256 (N_6256,N_5648,N_5948);
xor U6257 (N_6257,N_5720,N_5998);
or U6258 (N_6258,N_5804,N_5584);
or U6259 (N_6259,N_5850,N_5753);
and U6260 (N_6260,N_5753,N_5616);
nand U6261 (N_6261,N_5625,N_5658);
xor U6262 (N_6262,N_5684,N_5922);
nand U6263 (N_6263,N_5933,N_5807);
nand U6264 (N_6264,N_5975,N_5724);
or U6265 (N_6265,N_5581,N_5827);
xnor U6266 (N_6266,N_5823,N_5945);
and U6267 (N_6267,N_5945,N_5862);
nor U6268 (N_6268,N_5964,N_5538);
nand U6269 (N_6269,N_5698,N_5980);
nand U6270 (N_6270,N_5665,N_5648);
xnor U6271 (N_6271,N_5727,N_5868);
xnor U6272 (N_6272,N_5907,N_5916);
xor U6273 (N_6273,N_5997,N_5616);
nor U6274 (N_6274,N_5880,N_5667);
xor U6275 (N_6275,N_5528,N_5808);
nand U6276 (N_6276,N_5840,N_5601);
or U6277 (N_6277,N_5757,N_5948);
and U6278 (N_6278,N_5687,N_5575);
or U6279 (N_6279,N_5806,N_5996);
xor U6280 (N_6280,N_5741,N_5855);
nor U6281 (N_6281,N_5811,N_5843);
nand U6282 (N_6282,N_5761,N_5831);
nand U6283 (N_6283,N_5651,N_5540);
nand U6284 (N_6284,N_5541,N_5630);
or U6285 (N_6285,N_5657,N_5954);
xor U6286 (N_6286,N_5998,N_5722);
nor U6287 (N_6287,N_5529,N_5690);
and U6288 (N_6288,N_5924,N_5516);
nand U6289 (N_6289,N_5547,N_5972);
and U6290 (N_6290,N_5855,N_5963);
xor U6291 (N_6291,N_5563,N_5728);
nor U6292 (N_6292,N_5892,N_5792);
or U6293 (N_6293,N_5910,N_5609);
or U6294 (N_6294,N_5887,N_5562);
and U6295 (N_6295,N_5688,N_5588);
and U6296 (N_6296,N_5929,N_5758);
or U6297 (N_6297,N_5839,N_5699);
and U6298 (N_6298,N_5884,N_5678);
nor U6299 (N_6299,N_5846,N_5586);
nor U6300 (N_6300,N_5678,N_5848);
nand U6301 (N_6301,N_5506,N_5773);
nor U6302 (N_6302,N_5710,N_5843);
nand U6303 (N_6303,N_5728,N_5603);
or U6304 (N_6304,N_5667,N_5751);
or U6305 (N_6305,N_5637,N_5514);
xnor U6306 (N_6306,N_5837,N_5993);
nand U6307 (N_6307,N_5977,N_5943);
xor U6308 (N_6308,N_5613,N_5891);
or U6309 (N_6309,N_5568,N_5724);
or U6310 (N_6310,N_5993,N_5746);
nor U6311 (N_6311,N_5847,N_5574);
nor U6312 (N_6312,N_5658,N_5638);
and U6313 (N_6313,N_5826,N_5808);
nand U6314 (N_6314,N_5945,N_5603);
and U6315 (N_6315,N_5655,N_5926);
nand U6316 (N_6316,N_5607,N_5859);
nor U6317 (N_6317,N_5818,N_5751);
nand U6318 (N_6318,N_5883,N_5525);
xor U6319 (N_6319,N_5608,N_5500);
nor U6320 (N_6320,N_5626,N_5820);
or U6321 (N_6321,N_5738,N_5673);
xnor U6322 (N_6322,N_5585,N_5650);
and U6323 (N_6323,N_5838,N_5820);
nand U6324 (N_6324,N_5904,N_5919);
nor U6325 (N_6325,N_5755,N_5762);
nor U6326 (N_6326,N_5756,N_5922);
nor U6327 (N_6327,N_5553,N_5883);
nand U6328 (N_6328,N_5728,N_5839);
or U6329 (N_6329,N_5635,N_5570);
or U6330 (N_6330,N_5738,N_5684);
or U6331 (N_6331,N_5619,N_5834);
and U6332 (N_6332,N_5914,N_5811);
nor U6333 (N_6333,N_5918,N_5815);
xor U6334 (N_6334,N_5948,N_5773);
nor U6335 (N_6335,N_5503,N_5533);
or U6336 (N_6336,N_5848,N_5639);
xor U6337 (N_6337,N_5627,N_5584);
or U6338 (N_6338,N_5711,N_5653);
nand U6339 (N_6339,N_5546,N_5516);
nor U6340 (N_6340,N_5656,N_5667);
nand U6341 (N_6341,N_5788,N_5654);
nor U6342 (N_6342,N_5511,N_5786);
or U6343 (N_6343,N_5684,N_5776);
nor U6344 (N_6344,N_5930,N_5525);
nor U6345 (N_6345,N_5928,N_5820);
xnor U6346 (N_6346,N_5899,N_5644);
nand U6347 (N_6347,N_5689,N_5632);
nor U6348 (N_6348,N_5705,N_5532);
or U6349 (N_6349,N_5683,N_5612);
and U6350 (N_6350,N_5808,N_5745);
or U6351 (N_6351,N_5858,N_5998);
or U6352 (N_6352,N_5651,N_5948);
nor U6353 (N_6353,N_5727,N_5822);
or U6354 (N_6354,N_5883,N_5988);
nor U6355 (N_6355,N_5659,N_5543);
or U6356 (N_6356,N_5714,N_5547);
nor U6357 (N_6357,N_5601,N_5589);
or U6358 (N_6358,N_5555,N_5779);
and U6359 (N_6359,N_5964,N_5877);
xor U6360 (N_6360,N_5864,N_5767);
nand U6361 (N_6361,N_5732,N_5864);
or U6362 (N_6362,N_5824,N_5525);
xor U6363 (N_6363,N_5676,N_5501);
nand U6364 (N_6364,N_5640,N_5677);
nand U6365 (N_6365,N_5827,N_5697);
nor U6366 (N_6366,N_5831,N_5521);
or U6367 (N_6367,N_5918,N_5828);
and U6368 (N_6368,N_5742,N_5699);
nand U6369 (N_6369,N_5691,N_5986);
xor U6370 (N_6370,N_5679,N_5901);
and U6371 (N_6371,N_5642,N_5760);
xnor U6372 (N_6372,N_5885,N_5807);
xnor U6373 (N_6373,N_5808,N_5661);
or U6374 (N_6374,N_5550,N_5870);
nor U6375 (N_6375,N_5729,N_5762);
xnor U6376 (N_6376,N_5817,N_5890);
or U6377 (N_6377,N_5820,N_5592);
nor U6378 (N_6378,N_5959,N_5681);
xor U6379 (N_6379,N_5994,N_5798);
xor U6380 (N_6380,N_5524,N_5965);
nand U6381 (N_6381,N_5909,N_5511);
or U6382 (N_6382,N_5720,N_5795);
or U6383 (N_6383,N_5690,N_5815);
xnor U6384 (N_6384,N_5924,N_5697);
or U6385 (N_6385,N_5575,N_5546);
or U6386 (N_6386,N_5752,N_5853);
nor U6387 (N_6387,N_5584,N_5863);
or U6388 (N_6388,N_5830,N_5958);
nor U6389 (N_6389,N_5678,N_5725);
nand U6390 (N_6390,N_5712,N_5592);
nor U6391 (N_6391,N_5720,N_5963);
and U6392 (N_6392,N_5526,N_5616);
nand U6393 (N_6393,N_5500,N_5818);
nor U6394 (N_6394,N_5607,N_5994);
nor U6395 (N_6395,N_5515,N_5581);
xnor U6396 (N_6396,N_5555,N_5820);
xor U6397 (N_6397,N_5621,N_5818);
xnor U6398 (N_6398,N_5810,N_5882);
or U6399 (N_6399,N_5912,N_5798);
nand U6400 (N_6400,N_5995,N_5654);
nand U6401 (N_6401,N_5871,N_5731);
xnor U6402 (N_6402,N_5994,N_5788);
and U6403 (N_6403,N_5609,N_5722);
or U6404 (N_6404,N_5672,N_5946);
or U6405 (N_6405,N_5742,N_5836);
or U6406 (N_6406,N_5961,N_5551);
nand U6407 (N_6407,N_5905,N_5922);
xnor U6408 (N_6408,N_5762,N_5731);
or U6409 (N_6409,N_5844,N_5630);
nand U6410 (N_6410,N_5932,N_5822);
xnor U6411 (N_6411,N_5918,N_5814);
nor U6412 (N_6412,N_5845,N_5570);
nor U6413 (N_6413,N_5966,N_5517);
or U6414 (N_6414,N_5899,N_5995);
nor U6415 (N_6415,N_5500,N_5507);
nand U6416 (N_6416,N_5938,N_5838);
or U6417 (N_6417,N_5700,N_5830);
nor U6418 (N_6418,N_5500,N_5674);
xor U6419 (N_6419,N_5901,N_5814);
or U6420 (N_6420,N_5612,N_5913);
and U6421 (N_6421,N_5823,N_5979);
nor U6422 (N_6422,N_5785,N_5917);
xor U6423 (N_6423,N_5949,N_5511);
nand U6424 (N_6424,N_5901,N_5591);
nand U6425 (N_6425,N_5772,N_5520);
xnor U6426 (N_6426,N_5942,N_5910);
nand U6427 (N_6427,N_5522,N_5785);
nor U6428 (N_6428,N_5592,N_5602);
or U6429 (N_6429,N_5994,N_5981);
nand U6430 (N_6430,N_5937,N_5908);
xor U6431 (N_6431,N_5732,N_5529);
nor U6432 (N_6432,N_5527,N_5511);
nand U6433 (N_6433,N_5938,N_5654);
or U6434 (N_6434,N_5974,N_5554);
and U6435 (N_6435,N_5748,N_5572);
or U6436 (N_6436,N_5878,N_5542);
xnor U6437 (N_6437,N_5877,N_5993);
nor U6438 (N_6438,N_5874,N_5637);
and U6439 (N_6439,N_5593,N_5858);
or U6440 (N_6440,N_5769,N_5678);
nand U6441 (N_6441,N_5930,N_5809);
xor U6442 (N_6442,N_5571,N_5878);
nand U6443 (N_6443,N_5827,N_5563);
or U6444 (N_6444,N_5595,N_5888);
or U6445 (N_6445,N_5942,N_5860);
nor U6446 (N_6446,N_5752,N_5868);
or U6447 (N_6447,N_5510,N_5695);
or U6448 (N_6448,N_5867,N_5895);
nor U6449 (N_6449,N_5516,N_5531);
nor U6450 (N_6450,N_5791,N_5746);
and U6451 (N_6451,N_5747,N_5775);
nor U6452 (N_6452,N_5716,N_5691);
xor U6453 (N_6453,N_5716,N_5755);
and U6454 (N_6454,N_5923,N_5697);
xnor U6455 (N_6455,N_5594,N_5980);
nand U6456 (N_6456,N_5601,N_5943);
nand U6457 (N_6457,N_5944,N_5940);
or U6458 (N_6458,N_5545,N_5550);
xor U6459 (N_6459,N_5510,N_5524);
and U6460 (N_6460,N_5971,N_5974);
xnor U6461 (N_6461,N_5656,N_5953);
xnor U6462 (N_6462,N_5910,N_5821);
or U6463 (N_6463,N_5731,N_5583);
nor U6464 (N_6464,N_5984,N_5566);
nor U6465 (N_6465,N_5753,N_5515);
or U6466 (N_6466,N_5836,N_5887);
nor U6467 (N_6467,N_5989,N_5870);
and U6468 (N_6468,N_5967,N_5600);
nor U6469 (N_6469,N_5594,N_5969);
nor U6470 (N_6470,N_5926,N_5802);
nor U6471 (N_6471,N_5681,N_5804);
and U6472 (N_6472,N_5582,N_5682);
and U6473 (N_6473,N_5832,N_5537);
nor U6474 (N_6474,N_5550,N_5579);
or U6475 (N_6475,N_5894,N_5926);
xnor U6476 (N_6476,N_5955,N_5937);
and U6477 (N_6477,N_5844,N_5764);
nand U6478 (N_6478,N_5873,N_5797);
or U6479 (N_6479,N_5524,N_5815);
and U6480 (N_6480,N_5998,N_5523);
nor U6481 (N_6481,N_5604,N_5683);
and U6482 (N_6482,N_5794,N_5550);
nand U6483 (N_6483,N_5729,N_5739);
nand U6484 (N_6484,N_5870,N_5722);
and U6485 (N_6485,N_5535,N_5550);
or U6486 (N_6486,N_5684,N_5859);
xnor U6487 (N_6487,N_5626,N_5947);
nor U6488 (N_6488,N_5571,N_5860);
and U6489 (N_6489,N_5779,N_5524);
or U6490 (N_6490,N_5529,N_5703);
nor U6491 (N_6491,N_5761,N_5673);
xnor U6492 (N_6492,N_5870,N_5752);
nor U6493 (N_6493,N_5775,N_5748);
xor U6494 (N_6494,N_5648,N_5537);
nand U6495 (N_6495,N_5694,N_5646);
nand U6496 (N_6496,N_5728,N_5577);
xor U6497 (N_6497,N_5565,N_5662);
nor U6498 (N_6498,N_5979,N_5675);
xnor U6499 (N_6499,N_5515,N_5533);
xnor U6500 (N_6500,N_6478,N_6465);
xnor U6501 (N_6501,N_6157,N_6317);
or U6502 (N_6502,N_6011,N_6102);
nand U6503 (N_6503,N_6467,N_6235);
and U6504 (N_6504,N_6329,N_6381);
and U6505 (N_6505,N_6370,N_6158);
nand U6506 (N_6506,N_6496,N_6197);
or U6507 (N_6507,N_6130,N_6208);
or U6508 (N_6508,N_6117,N_6286);
or U6509 (N_6509,N_6249,N_6207);
or U6510 (N_6510,N_6195,N_6283);
xor U6511 (N_6511,N_6120,N_6420);
and U6512 (N_6512,N_6499,N_6042);
or U6513 (N_6513,N_6231,N_6243);
xnor U6514 (N_6514,N_6343,N_6264);
nand U6515 (N_6515,N_6245,N_6081);
nor U6516 (N_6516,N_6144,N_6429);
or U6517 (N_6517,N_6362,N_6482);
and U6518 (N_6518,N_6058,N_6006);
and U6519 (N_6519,N_6206,N_6457);
or U6520 (N_6520,N_6497,N_6349);
nand U6521 (N_6521,N_6475,N_6167);
and U6522 (N_6522,N_6080,N_6209);
nor U6523 (N_6523,N_6131,N_6160);
xor U6524 (N_6524,N_6422,N_6280);
or U6525 (N_6525,N_6187,N_6313);
nor U6526 (N_6526,N_6380,N_6299);
xor U6527 (N_6527,N_6139,N_6005);
and U6528 (N_6528,N_6142,N_6214);
and U6529 (N_6529,N_6059,N_6481);
or U6530 (N_6530,N_6169,N_6382);
and U6531 (N_6531,N_6010,N_6109);
and U6532 (N_6532,N_6057,N_6495);
and U6533 (N_6533,N_6066,N_6052);
xor U6534 (N_6534,N_6087,N_6035);
nand U6535 (N_6535,N_6076,N_6145);
xnor U6536 (N_6536,N_6082,N_6347);
nor U6537 (N_6537,N_6443,N_6425);
and U6538 (N_6538,N_6350,N_6150);
or U6539 (N_6539,N_6267,N_6315);
and U6540 (N_6540,N_6152,N_6348);
nor U6541 (N_6541,N_6427,N_6200);
and U6542 (N_6542,N_6259,N_6466);
nor U6543 (N_6543,N_6319,N_6141);
or U6544 (N_6544,N_6106,N_6376);
xnor U6545 (N_6545,N_6405,N_6357);
or U6546 (N_6546,N_6312,N_6045);
nand U6547 (N_6547,N_6198,N_6426);
nor U6548 (N_6548,N_6128,N_6203);
nand U6549 (N_6549,N_6251,N_6262);
nand U6550 (N_6550,N_6124,N_6322);
nand U6551 (N_6551,N_6114,N_6016);
xnor U6552 (N_6552,N_6476,N_6110);
nand U6553 (N_6553,N_6374,N_6234);
or U6554 (N_6554,N_6335,N_6159);
nand U6555 (N_6555,N_6423,N_6233);
xnor U6556 (N_6556,N_6301,N_6040);
nor U6557 (N_6557,N_6250,N_6260);
xnor U6558 (N_6558,N_6441,N_6053);
nand U6559 (N_6559,N_6397,N_6171);
or U6560 (N_6560,N_6229,N_6015);
xor U6561 (N_6561,N_6153,N_6133);
or U6562 (N_6562,N_6306,N_6196);
xnor U6563 (N_6563,N_6135,N_6077);
xor U6564 (N_6564,N_6492,N_6271);
nand U6565 (N_6565,N_6324,N_6212);
or U6566 (N_6566,N_6433,N_6377);
or U6567 (N_6567,N_6225,N_6177);
nor U6568 (N_6568,N_6173,N_6417);
or U6569 (N_6569,N_6136,N_6162);
and U6570 (N_6570,N_6257,N_6182);
xnor U6571 (N_6571,N_6291,N_6351);
nand U6572 (N_6572,N_6273,N_6289);
nor U6573 (N_6573,N_6092,N_6089);
nand U6574 (N_6574,N_6134,N_6193);
xnor U6575 (N_6575,N_6412,N_6118);
or U6576 (N_6576,N_6444,N_6383);
nor U6577 (N_6577,N_6388,N_6330);
xnor U6578 (N_6578,N_6334,N_6305);
nor U6579 (N_6579,N_6339,N_6392);
nand U6580 (N_6580,N_6189,N_6237);
or U6581 (N_6581,N_6013,N_6358);
and U6582 (N_6582,N_6075,N_6228);
nor U6583 (N_6583,N_6068,N_6007);
nand U6584 (N_6584,N_6211,N_6147);
xor U6585 (N_6585,N_6464,N_6097);
or U6586 (N_6586,N_6384,N_6111);
xnor U6587 (N_6587,N_6137,N_6026);
or U6588 (N_6588,N_6373,N_6226);
nand U6589 (N_6589,N_6093,N_6085);
nand U6590 (N_6590,N_6004,N_6454);
xor U6591 (N_6591,N_6101,N_6017);
nor U6592 (N_6592,N_6385,N_6029);
xor U6593 (N_6593,N_6073,N_6183);
nor U6594 (N_6594,N_6435,N_6000);
or U6595 (N_6595,N_6399,N_6166);
xnor U6596 (N_6596,N_6178,N_6254);
or U6597 (N_6597,N_6161,N_6459);
or U6598 (N_6598,N_6261,N_6105);
nor U6599 (N_6599,N_6170,N_6400);
nor U6600 (N_6600,N_6368,N_6325);
nand U6601 (N_6601,N_6001,N_6044);
and U6602 (N_6602,N_6323,N_6436);
nand U6603 (N_6603,N_6474,N_6176);
nor U6604 (N_6604,N_6471,N_6409);
xor U6605 (N_6605,N_6164,N_6486);
xor U6606 (N_6606,N_6270,N_6483);
or U6607 (N_6607,N_6210,N_6281);
and U6608 (N_6608,N_6452,N_6022);
nand U6609 (N_6609,N_6084,N_6356);
xnor U6610 (N_6610,N_6309,N_6043);
and U6611 (N_6611,N_6055,N_6300);
nor U6612 (N_6612,N_6445,N_6020);
or U6613 (N_6613,N_6121,N_6463);
nor U6614 (N_6614,N_6078,N_6242);
nand U6615 (N_6615,N_6155,N_6326);
xor U6616 (N_6616,N_6314,N_6132);
xor U6617 (N_6617,N_6151,N_6218);
nor U6618 (N_6618,N_6367,N_6244);
nand U6619 (N_6619,N_6424,N_6100);
xor U6620 (N_6620,N_6091,N_6072);
nor U6621 (N_6621,N_6494,N_6294);
nor U6622 (N_6622,N_6031,N_6061);
nand U6623 (N_6623,N_6217,N_6473);
and U6624 (N_6624,N_6258,N_6490);
nand U6625 (N_6625,N_6023,N_6440);
and U6626 (N_6626,N_6402,N_6297);
nor U6627 (N_6627,N_6449,N_6416);
nor U6628 (N_6628,N_6069,N_6143);
and U6629 (N_6629,N_6174,N_6192);
nor U6630 (N_6630,N_6282,N_6307);
nor U6631 (N_6631,N_6185,N_6221);
xor U6632 (N_6632,N_6468,N_6122);
xnor U6633 (N_6633,N_6034,N_6298);
nand U6634 (N_6634,N_6012,N_6239);
or U6635 (N_6635,N_6332,N_6126);
or U6636 (N_6636,N_6071,N_6403);
and U6637 (N_6637,N_6352,N_6363);
nor U6638 (N_6638,N_6172,N_6320);
xnor U6639 (N_6639,N_6096,N_6140);
nor U6640 (N_6640,N_6246,N_6318);
or U6641 (N_6641,N_6024,N_6149);
nor U6642 (N_6642,N_6014,N_6008);
nor U6643 (N_6643,N_6255,N_6458);
xnor U6644 (N_6644,N_6461,N_6252);
or U6645 (N_6645,N_6387,N_6491);
xnor U6646 (N_6646,N_6048,N_6009);
and U6647 (N_6647,N_6472,N_6265);
nand U6648 (N_6648,N_6179,N_6268);
nor U6649 (N_6649,N_6067,N_6365);
xor U6650 (N_6650,N_6107,N_6213);
xnor U6651 (N_6651,N_6359,N_6263);
nand U6652 (N_6652,N_6095,N_6060);
nand U6653 (N_6653,N_6431,N_6275);
nand U6654 (N_6654,N_6484,N_6498);
and U6655 (N_6655,N_6308,N_6401);
xnor U6656 (N_6656,N_6099,N_6232);
or U6657 (N_6657,N_6127,N_6311);
or U6658 (N_6658,N_6108,N_6278);
nand U6659 (N_6659,N_6393,N_6202);
and U6660 (N_6660,N_6079,N_6274);
nor U6661 (N_6661,N_6364,N_6293);
nor U6662 (N_6662,N_6333,N_6337);
nor U6663 (N_6663,N_6404,N_6215);
xor U6664 (N_6664,N_6340,N_6038);
xnor U6665 (N_6665,N_6050,N_6037);
xor U6666 (N_6666,N_6236,N_6375);
and U6667 (N_6667,N_6063,N_6480);
nand U6668 (N_6668,N_6406,N_6303);
xnor U6669 (N_6669,N_6002,N_6386);
nor U6670 (N_6670,N_6361,N_6338);
and U6671 (N_6671,N_6489,N_6088);
or U6672 (N_6672,N_6446,N_6408);
or U6673 (N_6673,N_6223,N_6154);
and U6674 (N_6674,N_6181,N_6028);
xor U6675 (N_6675,N_6276,N_6342);
and U6676 (N_6676,N_6451,N_6290);
nor U6677 (N_6677,N_6391,N_6240);
or U6678 (N_6678,N_6470,N_6190);
xnor U6679 (N_6679,N_6287,N_6410);
xor U6680 (N_6680,N_6025,N_6455);
and U6681 (N_6681,N_6032,N_6201);
nand U6682 (N_6682,N_6477,N_6241);
nand U6683 (N_6683,N_6113,N_6186);
and U6684 (N_6684,N_6411,N_6456);
nand U6685 (N_6685,N_6021,N_6033);
nand U6686 (N_6686,N_6331,N_6414);
and U6687 (N_6687,N_6062,N_6086);
and U6688 (N_6688,N_6041,N_6430);
and U6689 (N_6689,N_6194,N_6205);
or U6690 (N_6690,N_6366,N_6390);
nand U6691 (N_6691,N_6328,N_6418);
nor U6692 (N_6692,N_6094,N_6238);
and U6693 (N_6693,N_6056,N_6064);
and U6694 (N_6694,N_6074,N_6285);
and U6695 (N_6695,N_6460,N_6396);
or U6696 (N_6696,N_6219,N_6098);
xor U6697 (N_6697,N_6310,N_6054);
and U6698 (N_6698,N_6493,N_6046);
nand U6699 (N_6699,N_6447,N_6407);
nand U6700 (N_6700,N_6116,N_6138);
or U6701 (N_6701,N_6369,N_6360);
nor U6702 (N_6702,N_6372,N_6394);
nor U6703 (N_6703,N_6292,N_6302);
nor U6704 (N_6704,N_6353,N_6413);
nand U6705 (N_6705,N_6419,N_6327);
nor U6706 (N_6706,N_6277,N_6119);
nand U6707 (N_6707,N_6123,N_6224);
nand U6708 (N_6708,N_6272,N_6304);
or U6709 (N_6709,N_6487,N_6036);
and U6710 (N_6710,N_6230,N_6103);
or U6711 (N_6711,N_6165,N_6288);
nand U6712 (N_6712,N_6180,N_6438);
xnor U6713 (N_6713,N_6469,N_6432);
or U6714 (N_6714,N_6415,N_6039);
xor U6715 (N_6715,N_6070,N_6247);
or U6716 (N_6716,N_6453,N_6354);
nor U6717 (N_6717,N_6090,N_6346);
or U6718 (N_6718,N_6345,N_6148);
or U6719 (N_6719,N_6027,N_6175);
and U6720 (N_6720,N_6341,N_6485);
and U6721 (N_6721,N_6437,N_6191);
nand U6722 (N_6722,N_6065,N_6316);
or U6723 (N_6723,N_6129,N_6389);
nand U6724 (N_6724,N_6216,N_6163);
or U6725 (N_6725,N_6336,N_6488);
or U6726 (N_6726,N_6434,N_6115);
nand U6727 (N_6727,N_6321,N_6284);
and U6728 (N_6728,N_6083,N_6104);
and U6729 (N_6729,N_6256,N_6395);
nand U6730 (N_6730,N_6156,N_6248);
xor U6731 (N_6731,N_6030,N_6448);
or U6732 (N_6732,N_6371,N_6125);
nor U6733 (N_6733,N_6220,N_6378);
nand U6734 (N_6734,N_6344,N_6479);
and U6735 (N_6735,N_6222,N_6146);
nor U6736 (N_6736,N_6398,N_6266);
and U6737 (N_6737,N_6355,N_6450);
and U6738 (N_6738,N_6253,N_6188);
nand U6739 (N_6739,N_6049,N_6442);
nor U6740 (N_6740,N_6428,N_6204);
or U6741 (N_6741,N_6051,N_6019);
and U6742 (N_6742,N_6295,N_6279);
and U6743 (N_6743,N_6379,N_6047);
and U6744 (N_6744,N_6184,N_6003);
or U6745 (N_6745,N_6227,N_6112);
nor U6746 (N_6746,N_6296,N_6421);
nand U6747 (N_6747,N_6462,N_6439);
nor U6748 (N_6748,N_6269,N_6168);
nand U6749 (N_6749,N_6199,N_6018);
nor U6750 (N_6750,N_6110,N_6184);
nor U6751 (N_6751,N_6105,N_6204);
xnor U6752 (N_6752,N_6485,N_6244);
and U6753 (N_6753,N_6313,N_6030);
xor U6754 (N_6754,N_6151,N_6326);
nor U6755 (N_6755,N_6432,N_6204);
or U6756 (N_6756,N_6066,N_6233);
xor U6757 (N_6757,N_6041,N_6221);
and U6758 (N_6758,N_6128,N_6325);
nand U6759 (N_6759,N_6321,N_6015);
nor U6760 (N_6760,N_6355,N_6249);
or U6761 (N_6761,N_6212,N_6351);
nand U6762 (N_6762,N_6426,N_6197);
and U6763 (N_6763,N_6325,N_6073);
xor U6764 (N_6764,N_6425,N_6197);
nand U6765 (N_6765,N_6125,N_6267);
and U6766 (N_6766,N_6300,N_6470);
or U6767 (N_6767,N_6339,N_6499);
or U6768 (N_6768,N_6476,N_6033);
nand U6769 (N_6769,N_6178,N_6223);
or U6770 (N_6770,N_6315,N_6240);
nand U6771 (N_6771,N_6429,N_6284);
xor U6772 (N_6772,N_6496,N_6017);
xnor U6773 (N_6773,N_6329,N_6325);
or U6774 (N_6774,N_6320,N_6178);
and U6775 (N_6775,N_6074,N_6280);
nor U6776 (N_6776,N_6086,N_6373);
and U6777 (N_6777,N_6289,N_6124);
or U6778 (N_6778,N_6480,N_6175);
nor U6779 (N_6779,N_6142,N_6323);
or U6780 (N_6780,N_6163,N_6449);
nand U6781 (N_6781,N_6403,N_6074);
or U6782 (N_6782,N_6069,N_6395);
nand U6783 (N_6783,N_6336,N_6152);
nor U6784 (N_6784,N_6196,N_6286);
or U6785 (N_6785,N_6261,N_6455);
xor U6786 (N_6786,N_6030,N_6362);
and U6787 (N_6787,N_6044,N_6474);
nor U6788 (N_6788,N_6304,N_6493);
xor U6789 (N_6789,N_6229,N_6160);
xor U6790 (N_6790,N_6207,N_6219);
or U6791 (N_6791,N_6016,N_6499);
xor U6792 (N_6792,N_6147,N_6187);
xor U6793 (N_6793,N_6246,N_6169);
and U6794 (N_6794,N_6140,N_6249);
or U6795 (N_6795,N_6099,N_6285);
and U6796 (N_6796,N_6467,N_6200);
and U6797 (N_6797,N_6150,N_6013);
nand U6798 (N_6798,N_6111,N_6375);
or U6799 (N_6799,N_6155,N_6231);
and U6800 (N_6800,N_6414,N_6406);
nor U6801 (N_6801,N_6214,N_6315);
or U6802 (N_6802,N_6253,N_6123);
nand U6803 (N_6803,N_6335,N_6420);
and U6804 (N_6804,N_6438,N_6198);
and U6805 (N_6805,N_6030,N_6006);
nor U6806 (N_6806,N_6151,N_6123);
nor U6807 (N_6807,N_6302,N_6332);
xnor U6808 (N_6808,N_6331,N_6406);
or U6809 (N_6809,N_6071,N_6315);
or U6810 (N_6810,N_6471,N_6376);
xnor U6811 (N_6811,N_6130,N_6307);
nand U6812 (N_6812,N_6041,N_6128);
nor U6813 (N_6813,N_6433,N_6337);
xor U6814 (N_6814,N_6159,N_6281);
xor U6815 (N_6815,N_6454,N_6195);
or U6816 (N_6816,N_6458,N_6302);
and U6817 (N_6817,N_6079,N_6425);
xnor U6818 (N_6818,N_6474,N_6379);
or U6819 (N_6819,N_6390,N_6029);
or U6820 (N_6820,N_6497,N_6033);
nand U6821 (N_6821,N_6133,N_6349);
xor U6822 (N_6822,N_6440,N_6073);
xor U6823 (N_6823,N_6353,N_6358);
xnor U6824 (N_6824,N_6050,N_6489);
nor U6825 (N_6825,N_6082,N_6091);
nand U6826 (N_6826,N_6091,N_6272);
or U6827 (N_6827,N_6496,N_6485);
nand U6828 (N_6828,N_6050,N_6140);
nand U6829 (N_6829,N_6079,N_6234);
nand U6830 (N_6830,N_6308,N_6112);
xor U6831 (N_6831,N_6451,N_6177);
nand U6832 (N_6832,N_6311,N_6001);
nand U6833 (N_6833,N_6087,N_6392);
and U6834 (N_6834,N_6383,N_6220);
xnor U6835 (N_6835,N_6479,N_6101);
xor U6836 (N_6836,N_6188,N_6260);
xor U6837 (N_6837,N_6126,N_6261);
and U6838 (N_6838,N_6072,N_6436);
or U6839 (N_6839,N_6174,N_6215);
xnor U6840 (N_6840,N_6344,N_6127);
or U6841 (N_6841,N_6297,N_6370);
nand U6842 (N_6842,N_6274,N_6080);
nor U6843 (N_6843,N_6479,N_6473);
nand U6844 (N_6844,N_6499,N_6185);
xor U6845 (N_6845,N_6467,N_6400);
nand U6846 (N_6846,N_6492,N_6375);
or U6847 (N_6847,N_6300,N_6363);
xnor U6848 (N_6848,N_6243,N_6352);
xor U6849 (N_6849,N_6166,N_6285);
nor U6850 (N_6850,N_6364,N_6203);
nand U6851 (N_6851,N_6236,N_6309);
xor U6852 (N_6852,N_6449,N_6490);
nand U6853 (N_6853,N_6100,N_6416);
xor U6854 (N_6854,N_6235,N_6034);
nand U6855 (N_6855,N_6394,N_6353);
nor U6856 (N_6856,N_6271,N_6493);
nor U6857 (N_6857,N_6419,N_6317);
nor U6858 (N_6858,N_6063,N_6368);
and U6859 (N_6859,N_6054,N_6084);
and U6860 (N_6860,N_6470,N_6311);
or U6861 (N_6861,N_6182,N_6461);
and U6862 (N_6862,N_6398,N_6229);
nand U6863 (N_6863,N_6193,N_6070);
and U6864 (N_6864,N_6342,N_6192);
or U6865 (N_6865,N_6248,N_6041);
nor U6866 (N_6866,N_6412,N_6185);
nor U6867 (N_6867,N_6406,N_6338);
and U6868 (N_6868,N_6117,N_6137);
nand U6869 (N_6869,N_6166,N_6290);
nor U6870 (N_6870,N_6411,N_6497);
xor U6871 (N_6871,N_6347,N_6456);
or U6872 (N_6872,N_6476,N_6480);
nor U6873 (N_6873,N_6384,N_6311);
or U6874 (N_6874,N_6015,N_6177);
or U6875 (N_6875,N_6403,N_6275);
nor U6876 (N_6876,N_6373,N_6212);
xor U6877 (N_6877,N_6369,N_6478);
nand U6878 (N_6878,N_6462,N_6236);
xnor U6879 (N_6879,N_6070,N_6305);
nand U6880 (N_6880,N_6108,N_6305);
and U6881 (N_6881,N_6125,N_6470);
and U6882 (N_6882,N_6212,N_6238);
xnor U6883 (N_6883,N_6124,N_6115);
nand U6884 (N_6884,N_6047,N_6423);
xnor U6885 (N_6885,N_6446,N_6499);
or U6886 (N_6886,N_6163,N_6404);
and U6887 (N_6887,N_6106,N_6311);
nand U6888 (N_6888,N_6194,N_6421);
nand U6889 (N_6889,N_6269,N_6499);
xor U6890 (N_6890,N_6304,N_6186);
and U6891 (N_6891,N_6453,N_6176);
nand U6892 (N_6892,N_6489,N_6173);
and U6893 (N_6893,N_6363,N_6223);
xnor U6894 (N_6894,N_6175,N_6293);
nand U6895 (N_6895,N_6343,N_6348);
nor U6896 (N_6896,N_6453,N_6369);
nor U6897 (N_6897,N_6455,N_6224);
xnor U6898 (N_6898,N_6490,N_6118);
and U6899 (N_6899,N_6055,N_6398);
nor U6900 (N_6900,N_6058,N_6196);
and U6901 (N_6901,N_6186,N_6409);
nor U6902 (N_6902,N_6270,N_6124);
or U6903 (N_6903,N_6220,N_6237);
nand U6904 (N_6904,N_6338,N_6295);
nand U6905 (N_6905,N_6426,N_6136);
nand U6906 (N_6906,N_6274,N_6431);
xor U6907 (N_6907,N_6440,N_6436);
or U6908 (N_6908,N_6425,N_6471);
nor U6909 (N_6909,N_6381,N_6295);
or U6910 (N_6910,N_6189,N_6049);
nor U6911 (N_6911,N_6101,N_6176);
nor U6912 (N_6912,N_6497,N_6160);
nand U6913 (N_6913,N_6189,N_6361);
or U6914 (N_6914,N_6139,N_6125);
nor U6915 (N_6915,N_6190,N_6068);
nor U6916 (N_6916,N_6047,N_6365);
nand U6917 (N_6917,N_6388,N_6109);
xor U6918 (N_6918,N_6169,N_6015);
or U6919 (N_6919,N_6040,N_6419);
or U6920 (N_6920,N_6207,N_6206);
xor U6921 (N_6921,N_6024,N_6296);
xnor U6922 (N_6922,N_6099,N_6427);
or U6923 (N_6923,N_6327,N_6258);
nand U6924 (N_6924,N_6104,N_6241);
nor U6925 (N_6925,N_6314,N_6018);
xnor U6926 (N_6926,N_6204,N_6332);
nor U6927 (N_6927,N_6239,N_6458);
xor U6928 (N_6928,N_6302,N_6047);
nor U6929 (N_6929,N_6222,N_6010);
nor U6930 (N_6930,N_6426,N_6274);
xor U6931 (N_6931,N_6468,N_6113);
xnor U6932 (N_6932,N_6203,N_6485);
nand U6933 (N_6933,N_6270,N_6187);
and U6934 (N_6934,N_6172,N_6095);
nor U6935 (N_6935,N_6422,N_6232);
nor U6936 (N_6936,N_6225,N_6239);
nand U6937 (N_6937,N_6224,N_6097);
nor U6938 (N_6938,N_6159,N_6186);
nand U6939 (N_6939,N_6062,N_6037);
and U6940 (N_6940,N_6205,N_6228);
nor U6941 (N_6941,N_6179,N_6091);
or U6942 (N_6942,N_6102,N_6192);
and U6943 (N_6943,N_6015,N_6157);
nand U6944 (N_6944,N_6237,N_6400);
nand U6945 (N_6945,N_6048,N_6163);
and U6946 (N_6946,N_6121,N_6024);
xnor U6947 (N_6947,N_6000,N_6204);
and U6948 (N_6948,N_6350,N_6443);
nand U6949 (N_6949,N_6409,N_6166);
nor U6950 (N_6950,N_6186,N_6442);
xor U6951 (N_6951,N_6464,N_6100);
and U6952 (N_6952,N_6025,N_6173);
or U6953 (N_6953,N_6016,N_6134);
or U6954 (N_6954,N_6161,N_6442);
nand U6955 (N_6955,N_6137,N_6410);
nor U6956 (N_6956,N_6116,N_6253);
and U6957 (N_6957,N_6256,N_6043);
xnor U6958 (N_6958,N_6022,N_6479);
or U6959 (N_6959,N_6177,N_6046);
nand U6960 (N_6960,N_6493,N_6316);
and U6961 (N_6961,N_6171,N_6255);
nand U6962 (N_6962,N_6146,N_6071);
or U6963 (N_6963,N_6169,N_6453);
or U6964 (N_6964,N_6410,N_6007);
xor U6965 (N_6965,N_6040,N_6376);
xnor U6966 (N_6966,N_6483,N_6232);
xor U6967 (N_6967,N_6380,N_6454);
and U6968 (N_6968,N_6215,N_6049);
xor U6969 (N_6969,N_6385,N_6290);
and U6970 (N_6970,N_6218,N_6429);
or U6971 (N_6971,N_6250,N_6351);
nand U6972 (N_6972,N_6062,N_6491);
nand U6973 (N_6973,N_6455,N_6189);
nand U6974 (N_6974,N_6437,N_6484);
or U6975 (N_6975,N_6055,N_6492);
xnor U6976 (N_6976,N_6280,N_6088);
xor U6977 (N_6977,N_6420,N_6185);
xor U6978 (N_6978,N_6048,N_6438);
and U6979 (N_6979,N_6311,N_6193);
and U6980 (N_6980,N_6111,N_6151);
xnor U6981 (N_6981,N_6244,N_6361);
nor U6982 (N_6982,N_6161,N_6380);
nor U6983 (N_6983,N_6421,N_6048);
nor U6984 (N_6984,N_6300,N_6060);
and U6985 (N_6985,N_6033,N_6131);
xor U6986 (N_6986,N_6340,N_6468);
nor U6987 (N_6987,N_6389,N_6027);
xor U6988 (N_6988,N_6395,N_6085);
and U6989 (N_6989,N_6024,N_6497);
nor U6990 (N_6990,N_6265,N_6219);
or U6991 (N_6991,N_6192,N_6120);
xnor U6992 (N_6992,N_6162,N_6428);
nand U6993 (N_6993,N_6109,N_6401);
and U6994 (N_6994,N_6138,N_6256);
or U6995 (N_6995,N_6490,N_6369);
nor U6996 (N_6996,N_6174,N_6237);
nor U6997 (N_6997,N_6006,N_6170);
nor U6998 (N_6998,N_6138,N_6456);
xnor U6999 (N_6999,N_6476,N_6344);
or U7000 (N_7000,N_6847,N_6877);
and U7001 (N_7001,N_6541,N_6763);
or U7002 (N_7002,N_6741,N_6955);
and U7003 (N_7003,N_6635,N_6904);
or U7004 (N_7004,N_6890,N_6585);
and U7005 (N_7005,N_6582,N_6559);
nand U7006 (N_7006,N_6719,N_6994);
nand U7007 (N_7007,N_6803,N_6907);
nand U7008 (N_7008,N_6882,N_6522);
and U7009 (N_7009,N_6927,N_6628);
and U7010 (N_7010,N_6985,N_6968);
xor U7011 (N_7011,N_6864,N_6814);
nor U7012 (N_7012,N_6571,N_6948);
or U7013 (N_7013,N_6788,N_6731);
and U7014 (N_7014,N_6641,N_6746);
or U7015 (N_7015,N_6798,N_6695);
xnor U7016 (N_7016,N_6850,N_6956);
nand U7017 (N_7017,N_6880,N_6509);
nor U7018 (N_7018,N_6970,N_6644);
or U7019 (N_7019,N_6657,N_6769);
and U7020 (N_7020,N_6820,N_6512);
xnor U7021 (N_7021,N_6526,N_6900);
nand U7022 (N_7022,N_6716,N_6781);
and U7023 (N_7023,N_6954,N_6605);
and U7024 (N_7024,N_6910,N_6825);
nand U7025 (N_7025,N_6940,N_6666);
and U7026 (N_7026,N_6663,N_6711);
xnor U7027 (N_7027,N_6751,N_6578);
xor U7028 (N_7028,N_6561,N_6755);
or U7029 (N_7029,N_6744,N_6545);
nor U7030 (N_7030,N_6809,N_6501);
xnor U7031 (N_7031,N_6996,N_6566);
nand U7032 (N_7032,N_6713,N_6967);
and U7033 (N_7033,N_6849,N_6584);
xnor U7034 (N_7034,N_6911,N_6888);
and U7035 (N_7035,N_6873,N_6599);
nor U7036 (N_7036,N_6913,N_6560);
and U7037 (N_7037,N_6852,N_6548);
xnor U7038 (N_7038,N_6879,N_6859);
nor U7039 (N_7039,N_6619,N_6683);
or U7040 (N_7040,N_6924,N_6909);
or U7041 (N_7041,N_6588,N_6524);
nand U7042 (N_7042,N_6801,N_6887);
or U7043 (N_7043,N_6530,N_6831);
nor U7044 (N_7044,N_6700,N_6777);
or U7045 (N_7045,N_6670,N_6997);
or U7046 (N_7046,N_6813,N_6511);
nand U7047 (N_7047,N_6822,N_6577);
xor U7048 (N_7048,N_6868,N_6923);
nor U7049 (N_7049,N_6527,N_6608);
or U7050 (N_7050,N_6915,N_6826);
and U7051 (N_7051,N_6782,N_6840);
xnor U7052 (N_7052,N_6963,N_6538);
and U7053 (N_7053,N_6710,N_6544);
or U7054 (N_7054,N_6691,N_6689);
xnor U7055 (N_7055,N_6676,N_6866);
and U7056 (N_7056,N_6837,N_6944);
and U7057 (N_7057,N_6978,N_6598);
xnor U7058 (N_7058,N_6858,N_6523);
nand U7059 (N_7059,N_6917,N_6974);
and U7060 (N_7060,N_6836,N_6933);
and U7061 (N_7061,N_6543,N_6694);
nand U7062 (N_7062,N_6747,N_6816);
or U7063 (N_7063,N_6611,N_6602);
or U7064 (N_7064,N_6701,N_6680);
nand U7065 (N_7065,N_6965,N_6827);
and U7066 (N_7066,N_6568,N_6705);
nor U7067 (N_7067,N_6515,N_6895);
or U7068 (N_7068,N_6762,N_6966);
and U7069 (N_7069,N_6946,N_6606);
nor U7070 (N_7070,N_6627,N_6596);
and U7071 (N_7071,N_6648,N_6776);
nor U7072 (N_7072,N_6665,N_6554);
or U7073 (N_7073,N_6844,N_6754);
nor U7074 (N_7074,N_6703,N_6579);
nand U7075 (N_7075,N_6592,N_6929);
or U7076 (N_7076,N_6613,N_6991);
nor U7077 (N_7077,N_6727,N_6979);
or U7078 (N_7078,N_6576,N_6764);
and U7079 (N_7079,N_6516,N_6630);
and U7080 (N_7080,N_6500,N_6674);
nor U7081 (N_7081,N_6614,N_6875);
nand U7082 (N_7082,N_6563,N_6797);
xnor U7083 (N_7083,N_6787,N_6988);
or U7084 (N_7084,N_6658,N_6999);
nor U7085 (N_7085,N_6779,N_6730);
nor U7086 (N_7086,N_6867,N_6672);
xor U7087 (N_7087,N_6681,N_6745);
or U7088 (N_7088,N_6795,N_6589);
nor U7089 (N_7089,N_6704,N_6732);
or U7090 (N_7090,N_6505,N_6819);
nor U7091 (N_7091,N_6686,N_6564);
nor U7092 (N_7092,N_6637,N_6977);
nand U7093 (N_7093,N_6855,N_6671);
xnor U7094 (N_7094,N_6862,N_6918);
or U7095 (N_7095,N_6941,N_6542);
nor U7096 (N_7096,N_6600,N_6891);
or U7097 (N_7097,N_6869,N_6612);
nor U7098 (N_7098,N_6934,N_6659);
nor U7099 (N_7099,N_6921,N_6793);
nand U7100 (N_7100,N_6894,N_6765);
nand U7101 (N_7101,N_6930,N_6513);
nor U7102 (N_7102,N_6536,N_6987);
xor U7103 (N_7103,N_6848,N_6767);
xnor U7104 (N_7104,N_6992,N_6722);
nand U7105 (N_7105,N_6631,N_6636);
nor U7106 (N_7106,N_6706,N_6652);
and U7107 (N_7107,N_6539,N_6950);
nor U7108 (N_7108,N_6558,N_6519);
nand U7109 (N_7109,N_6724,N_6983);
nor U7110 (N_7110,N_6982,N_6808);
nand U7111 (N_7111,N_6789,N_6839);
and U7112 (N_7112,N_6651,N_6533);
and U7113 (N_7113,N_6573,N_6502);
and U7114 (N_7114,N_6698,N_6734);
nand U7115 (N_7115,N_6699,N_6726);
and U7116 (N_7116,N_6626,N_6766);
and U7117 (N_7117,N_6667,N_6936);
xor U7118 (N_7118,N_6898,N_6802);
and U7119 (N_7119,N_6846,N_6521);
nand U7120 (N_7120,N_6785,N_6647);
nor U7121 (N_7121,N_6622,N_6957);
xor U7122 (N_7122,N_6749,N_6534);
or U7123 (N_7123,N_6832,N_6897);
and U7124 (N_7124,N_6908,N_6640);
nor U7125 (N_7125,N_6770,N_6572);
nor U7126 (N_7126,N_6595,N_6684);
or U7127 (N_7127,N_6815,N_6581);
xnor U7128 (N_7128,N_6899,N_6871);
nand U7129 (N_7129,N_6893,N_6980);
or U7130 (N_7130,N_6790,N_6857);
nand U7131 (N_7131,N_6853,N_6823);
nand U7132 (N_7132,N_6675,N_6620);
or U7133 (N_7133,N_6773,N_6737);
and U7134 (N_7134,N_6903,N_6661);
or U7135 (N_7135,N_6817,N_6778);
nand U7136 (N_7136,N_6796,N_6646);
and U7137 (N_7137,N_6972,N_6553);
and U7138 (N_7138,N_6607,N_6926);
nand U7139 (N_7139,N_6811,N_6570);
or U7140 (N_7140,N_6738,N_6678);
nand U7141 (N_7141,N_6506,N_6531);
and U7142 (N_7142,N_6914,N_6717);
nand U7143 (N_7143,N_6696,N_6679);
nand U7144 (N_7144,N_6725,N_6551);
nand U7145 (N_7145,N_6775,N_6842);
and U7146 (N_7146,N_6884,N_6721);
nor U7147 (N_7147,N_6960,N_6750);
xor U7148 (N_7148,N_6885,N_6510);
nand U7149 (N_7149,N_6922,N_6669);
and U7150 (N_7150,N_6593,N_6949);
xnor U7151 (N_7151,N_6952,N_6958);
and U7152 (N_7152,N_6739,N_6756);
xor U7153 (N_7153,N_6951,N_6935);
or U7154 (N_7154,N_6520,N_6580);
and U7155 (N_7155,N_6990,N_6919);
or U7156 (N_7156,N_6861,N_6625);
xnor U7157 (N_7157,N_6537,N_6673);
xnor U7158 (N_7158,N_6708,N_6591);
and U7159 (N_7159,N_6702,N_6889);
or U7160 (N_7160,N_6805,N_6780);
nor U7161 (N_7161,N_6791,N_6690);
xor U7162 (N_7162,N_6757,N_6604);
and U7163 (N_7163,N_6616,N_6540);
or U7164 (N_7164,N_6851,N_6892);
nand U7165 (N_7165,N_6712,N_6902);
and U7166 (N_7166,N_6733,N_6574);
nand U7167 (N_7167,N_6752,N_6761);
and U7168 (N_7168,N_6723,N_6655);
or U7169 (N_7169,N_6845,N_6740);
nor U7170 (N_7170,N_6772,N_6828);
or U7171 (N_7171,N_6975,N_6925);
xor U7172 (N_7172,N_6800,N_6742);
xnor U7173 (N_7173,N_6938,N_6807);
nand U7174 (N_7174,N_6718,N_6986);
nand U7175 (N_7175,N_6664,N_6901);
xnor U7176 (N_7176,N_6623,N_6586);
and U7177 (N_7177,N_6629,N_6618);
and U7178 (N_7178,N_6682,N_6896);
and U7179 (N_7179,N_6945,N_6624);
nor U7180 (N_7180,N_6714,N_6784);
xnor U7181 (N_7181,N_6841,N_6514);
nand U7182 (N_7182,N_6931,N_6878);
nor U7183 (N_7183,N_6621,N_6818);
xnor U7184 (N_7184,N_6947,N_6617);
nand U7185 (N_7185,N_6920,N_6662);
nor U7186 (N_7186,N_6874,N_6964);
nand U7187 (N_7187,N_6928,N_6653);
nor U7188 (N_7188,N_6830,N_6633);
and U7189 (N_7189,N_6565,N_6771);
xnor U7190 (N_7190,N_6833,N_6870);
xor U7191 (N_7191,N_6504,N_6609);
and U7192 (N_7192,N_6525,N_6863);
nor U7193 (N_7193,N_6507,N_6768);
nand U7194 (N_7194,N_6720,N_6692);
and U7195 (N_7195,N_6760,N_6656);
xor U7196 (N_7196,N_6989,N_6654);
and U7197 (N_7197,N_6856,N_6995);
xnor U7198 (N_7198,N_6806,N_6562);
or U7199 (N_7199,N_6594,N_6804);
nor U7200 (N_7200,N_6835,N_6953);
nor U7201 (N_7201,N_6906,N_6555);
nor U7202 (N_7202,N_6829,N_6687);
nor U7203 (N_7203,N_6984,N_6993);
nor U7204 (N_7204,N_6677,N_6615);
nor U7205 (N_7205,N_6552,N_6834);
xnor U7206 (N_7206,N_6697,N_6735);
xnor U7207 (N_7207,N_6883,N_6729);
xor U7208 (N_7208,N_6799,N_6583);
and U7209 (N_7209,N_6812,N_6645);
nand U7210 (N_7210,N_6550,N_6529);
and U7211 (N_7211,N_6753,N_6961);
xnor U7212 (N_7212,N_6707,N_6971);
and U7213 (N_7213,N_6546,N_6532);
and U7214 (N_7214,N_6556,N_6969);
and U7215 (N_7215,N_6643,N_6557);
or U7216 (N_7216,N_6998,N_6547);
xor U7217 (N_7217,N_6528,N_6569);
nand U7218 (N_7218,N_6603,N_6792);
nor U7219 (N_7219,N_6508,N_6821);
or U7220 (N_7220,N_6728,N_6709);
nand U7221 (N_7221,N_6549,N_6786);
and U7222 (N_7222,N_6597,N_6876);
nor U7223 (N_7223,N_6905,N_6824);
nor U7224 (N_7224,N_6976,N_6872);
or U7225 (N_7225,N_6517,N_6937);
nor U7226 (N_7226,N_6575,N_6783);
or U7227 (N_7227,N_6590,N_6774);
nor U7228 (N_7228,N_6838,N_6518);
or U7229 (N_7229,N_6794,N_6962);
nand U7230 (N_7230,N_6668,N_6973);
or U7231 (N_7231,N_6881,N_6810);
nor U7232 (N_7232,N_6634,N_6649);
or U7233 (N_7233,N_6610,N_6685);
or U7234 (N_7234,N_6642,N_6693);
xor U7235 (N_7235,N_6959,N_6865);
or U7236 (N_7236,N_6736,N_6759);
nor U7237 (N_7237,N_6860,N_6503);
nor U7238 (N_7238,N_6932,N_6639);
nor U7239 (N_7239,N_6743,N_6942);
and U7240 (N_7240,N_6715,N_6660);
nand U7241 (N_7241,N_6758,N_6567);
nor U7242 (N_7242,N_6638,N_6939);
xnor U7243 (N_7243,N_6688,N_6632);
nand U7244 (N_7244,N_6843,N_6535);
xnor U7245 (N_7245,N_6943,N_6981);
or U7246 (N_7246,N_6587,N_6601);
xnor U7247 (N_7247,N_6886,N_6650);
nand U7248 (N_7248,N_6854,N_6916);
or U7249 (N_7249,N_6912,N_6748);
or U7250 (N_7250,N_6528,N_6596);
nand U7251 (N_7251,N_6736,N_6866);
nor U7252 (N_7252,N_6703,N_6938);
and U7253 (N_7253,N_6819,N_6665);
nor U7254 (N_7254,N_6563,N_6936);
or U7255 (N_7255,N_6999,N_6789);
nand U7256 (N_7256,N_6692,N_6711);
nand U7257 (N_7257,N_6648,N_6689);
nand U7258 (N_7258,N_6547,N_6696);
nor U7259 (N_7259,N_6841,N_6845);
nand U7260 (N_7260,N_6880,N_6518);
and U7261 (N_7261,N_6558,N_6916);
and U7262 (N_7262,N_6595,N_6809);
nor U7263 (N_7263,N_6718,N_6543);
nand U7264 (N_7264,N_6829,N_6694);
xnor U7265 (N_7265,N_6690,N_6623);
nor U7266 (N_7266,N_6965,N_6792);
xor U7267 (N_7267,N_6612,N_6574);
and U7268 (N_7268,N_6798,N_6919);
nand U7269 (N_7269,N_6963,N_6598);
or U7270 (N_7270,N_6909,N_6806);
nand U7271 (N_7271,N_6965,N_6503);
nand U7272 (N_7272,N_6850,N_6573);
nor U7273 (N_7273,N_6603,N_6503);
or U7274 (N_7274,N_6857,N_6733);
nor U7275 (N_7275,N_6929,N_6988);
nand U7276 (N_7276,N_6944,N_6565);
nand U7277 (N_7277,N_6719,N_6856);
or U7278 (N_7278,N_6710,N_6679);
xnor U7279 (N_7279,N_6553,N_6869);
xor U7280 (N_7280,N_6593,N_6697);
nor U7281 (N_7281,N_6522,N_6951);
nor U7282 (N_7282,N_6526,N_6853);
xnor U7283 (N_7283,N_6751,N_6733);
xor U7284 (N_7284,N_6601,N_6733);
xnor U7285 (N_7285,N_6785,N_6681);
nor U7286 (N_7286,N_6693,N_6592);
nor U7287 (N_7287,N_6733,N_6692);
xnor U7288 (N_7288,N_6687,N_6606);
xor U7289 (N_7289,N_6599,N_6945);
and U7290 (N_7290,N_6998,N_6946);
and U7291 (N_7291,N_6585,N_6619);
xnor U7292 (N_7292,N_6773,N_6711);
xnor U7293 (N_7293,N_6655,N_6740);
or U7294 (N_7294,N_6689,N_6517);
or U7295 (N_7295,N_6941,N_6573);
or U7296 (N_7296,N_6936,N_6969);
or U7297 (N_7297,N_6746,N_6749);
nor U7298 (N_7298,N_6860,N_6517);
xor U7299 (N_7299,N_6646,N_6818);
or U7300 (N_7300,N_6556,N_6936);
nor U7301 (N_7301,N_6694,N_6600);
nand U7302 (N_7302,N_6970,N_6851);
nor U7303 (N_7303,N_6878,N_6927);
nand U7304 (N_7304,N_6924,N_6875);
xor U7305 (N_7305,N_6690,N_6983);
or U7306 (N_7306,N_6752,N_6662);
nand U7307 (N_7307,N_6820,N_6901);
nand U7308 (N_7308,N_6722,N_6965);
nand U7309 (N_7309,N_6748,N_6905);
or U7310 (N_7310,N_6908,N_6975);
or U7311 (N_7311,N_6847,N_6934);
or U7312 (N_7312,N_6610,N_6717);
xor U7313 (N_7313,N_6779,N_6587);
and U7314 (N_7314,N_6733,N_6713);
nor U7315 (N_7315,N_6622,N_6760);
or U7316 (N_7316,N_6942,N_6627);
nor U7317 (N_7317,N_6706,N_6685);
xor U7318 (N_7318,N_6889,N_6563);
nand U7319 (N_7319,N_6603,N_6627);
nand U7320 (N_7320,N_6532,N_6517);
nand U7321 (N_7321,N_6670,N_6941);
nand U7322 (N_7322,N_6994,N_6580);
nor U7323 (N_7323,N_6884,N_6646);
and U7324 (N_7324,N_6731,N_6881);
xnor U7325 (N_7325,N_6939,N_6911);
nor U7326 (N_7326,N_6705,N_6662);
or U7327 (N_7327,N_6516,N_6664);
and U7328 (N_7328,N_6685,N_6861);
xnor U7329 (N_7329,N_6948,N_6787);
and U7330 (N_7330,N_6948,N_6610);
nand U7331 (N_7331,N_6980,N_6957);
or U7332 (N_7332,N_6504,N_6584);
nor U7333 (N_7333,N_6545,N_6740);
or U7334 (N_7334,N_6695,N_6687);
xor U7335 (N_7335,N_6853,N_6661);
xnor U7336 (N_7336,N_6973,N_6705);
nor U7337 (N_7337,N_6961,N_6772);
and U7338 (N_7338,N_6898,N_6658);
and U7339 (N_7339,N_6617,N_6702);
nand U7340 (N_7340,N_6703,N_6572);
or U7341 (N_7341,N_6932,N_6501);
or U7342 (N_7342,N_6728,N_6914);
xor U7343 (N_7343,N_6849,N_6958);
nor U7344 (N_7344,N_6586,N_6860);
nand U7345 (N_7345,N_6819,N_6606);
xnor U7346 (N_7346,N_6763,N_6658);
xor U7347 (N_7347,N_6576,N_6651);
xnor U7348 (N_7348,N_6906,N_6718);
and U7349 (N_7349,N_6865,N_6784);
and U7350 (N_7350,N_6860,N_6533);
and U7351 (N_7351,N_6985,N_6764);
nor U7352 (N_7352,N_6515,N_6839);
nor U7353 (N_7353,N_6815,N_6504);
or U7354 (N_7354,N_6995,N_6514);
nand U7355 (N_7355,N_6825,N_6628);
nand U7356 (N_7356,N_6739,N_6974);
or U7357 (N_7357,N_6866,N_6886);
or U7358 (N_7358,N_6804,N_6671);
xor U7359 (N_7359,N_6656,N_6738);
nor U7360 (N_7360,N_6519,N_6690);
nor U7361 (N_7361,N_6935,N_6706);
xor U7362 (N_7362,N_6848,N_6503);
nor U7363 (N_7363,N_6792,N_6674);
nor U7364 (N_7364,N_6806,N_6645);
and U7365 (N_7365,N_6591,N_6627);
and U7366 (N_7366,N_6682,N_6932);
nand U7367 (N_7367,N_6693,N_6580);
nand U7368 (N_7368,N_6677,N_6880);
nand U7369 (N_7369,N_6609,N_6818);
nor U7370 (N_7370,N_6695,N_6944);
nor U7371 (N_7371,N_6952,N_6902);
nand U7372 (N_7372,N_6924,N_6502);
and U7373 (N_7373,N_6969,N_6903);
nor U7374 (N_7374,N_6788,N_6768);
nor U7375 (N_7375,N_6864,N_6800);
nor U7376 (N_7376,N_6690,N_6748);
nand U7377 (N_7377,N_6551,N_6517);
or U7378 (N_7378,N_6550,N_6912);
nand U7379 (N_7379,N_6796,N_6585);
xor U7380 (N_7380,N_6790,N_6568);
or U7381 (N_7381,N_6845,N_6923);
nor U7382 (N_7382,N_6655,N_6813);
xnor U7383 (N_7383,N_6540,N_6719);
xnor U7384 (N_7384,N_6767,N_6954);
xor U7385 (N_7385,N_6614,N_6743);
or U7386 (N_7386,N_6789,N_6709);
nor U7387 (N_7387,N_6774,N_6979);
and U7388 (N_7388,N_6987,N_6889);
xor U7389 (N_7389,N_6592,N_6850);
or U7390 (N_7390,N_6797,N_6959);
or U7391 (N_7391,N_6705,N_6796);
xor U7392 (N_7392,N_6664,N_6948);
nand U7393 (N_7393,N_6723,N_6553);
or U7394 (N_7394,N_6619,N_6862);
and U7395 (N_7395,N_6802,N_6974);
nor U7396 (N_7396,N_6686,N_6837);
xnor U7397 (N_7397,N_6818,N_6740);
or U7398 (N_7398,N_6969,N_6916);
or U7399 (N_7399,N_6591,N_6940);
xor U7400 (N_7400,N_6823,N_6558);
or U7401 (N_7401,N_6560,N_6793);
nor U7402 (N_7402,N_6973,N_6600);
and U7403 (N_7403,N_6994,N_6675);
nand U7404 (N_7404,N_6877,N_6916);
or U7405 (N_7405,N_6966,N_6548);
xnor U7406 (N_7406,N_6671,N_6824);
and U7407 (N_7407,N_6573,N_6548);
or U7408 (N_7408,N_6848,N_6909);
nor U7409 (N_7409,N_6803,N_6842);
and U7410 (N_7410,N_6640,N_6539);
xor U7411 (N_7411,N_6703,N_6567);
and U7412 (N_7412,N_6939,N_6887);
or U7413 (N_7413,N_6561,N_6662);
and U7414 (N_7414,N_6513,N_6712);
and U7415 (N_7415,N_6999,N_6802);
and U7416 (N_7416,N_6545,N_6716);
and U7417 (N_7417,N_6813,N_6776);
nor U7418 (N_7418,N_6762,N_6976);
or U7419 (N_7419,N_6945,N_6556);
xor U7420 (N_7420,N_6629,N_6909);
and U7421 (N_7421,N_6685,N_6680);
nand U7422 (N_7422,N_6755,N_6749);
xor U7423 (N_7423,N_6519,N_6790);
and U7424 (N_7424,N_6603,N_6577);
xnor U7425 (N_7425,N_6753,N_6996);
and U7426 (N_7426,N_6883,N_6994);
and U7427 (N_7427,N_6863,N_6538);
nor U7428 (N_7428,N_6713,N_6613);
nor U7429 (N_7429,N_6546,N_6681);
or U7430 (N_7430,N_6588,N_6584);
and U7431 (N_7431,N_6834,N_6653);
xnor U7432 (N_7432,N_6969,N_6878);
xor U7433 (N_7433,N_6739,N_6791);
nor U7434 (N_7434,N_6529,N_6617);
xor U7435 (N_7435,N_6861,N_6891);
and U7436 (N_7436,N_6949,N_6760);
and U7437 (N_7437,N_6975,N_6863);
xor U7438 (N_7438,N_6862,N_6638);
nand U7439 (N_7439,N_6644,N_6503);
and U7440 (N_7440,N_6659,N_6843);
nand U7441 (N_7441,N_6846,N_6664);
xor U7442 (N_7442,N_6950,N_6966);
nor U7443 (N_7443,N_6623,N_6536);
and U7444 (N_7444,N_6873,N_6688);
xnor U7445 (N_7445,N_6599,N_6819);
nand U7446 (N_7446,N_6711,N_6937);
nand U7447 (N_7447,N_6900,N_6561);
or U7448 (N_7448,N_6703,N_6791);
xnor U7449 (N_7449,N_6694,N_6729);
or U7450 (N_7450,N_6838,N_6697);
xnor U7451 (N_7451,N_6852,N_6848);
nand U7452 (N_7452,N_6615,N_6907);
and U7453 (N_7453,N_6506,N_6988);
or U7454 (N_7454,N_6925,N_6585);
and U7455 (N_7455,N_6778,N_6710);
nand U7456 (N_7456,N_6843,N_6984);
xor U7457 (N_7457,N_6690,N_6546);
nor U7458 (N_7458,N_6867,N_6907);
xor U7459 (N_7459,N_6570,N_6675);
nor U7460 (N_7460,N_6908,N_6549);
nor U7461 (N_7461,N_6719,N_6882);
nand U7462 (N_7462,N_6598,N_6752);
xnor U7463 (N_7463,N_6726,N_6832);
or U7464 (N_7464,N_6668,N_6889);
nand U7465 (N_7465,N_6751,N_6547);
or U7466 (N_7466,N_6742,N_6608);
and U7467 (N_7467,N_6959,N_6925);
nor U7468 (N_7468,N_6956,N_6619);
nor U7469 (N_7469,N_6962,N_6762);
nor U7470 (N_7470,N_6641,N_6515);
nand U7471 (N_7471,N_6672,N_6919);
xor U7472 (N_7472,N_6541,N_6602);
xor U7473 (N_7473,N_6851,N_6518);
nand U7474 (N_7474,N_6776,N_6517);
or U7475 (N_7475,N_6750,N_6666);
nor U7476 (N_7476,N_6737,N_6558);
xnor U7477 (N_7477,N_6766,N_6922);
and U7478 (N_7478,N_6921,N_6576);
xnor U7479 (N_7479,N_6779,N_6834);
xor U7480 (N_7480,N_6858,N_6585);
xnor U7481 (N_7481,N_6817,N_6862);
and U7482 (N_7482,N_6563,N_6827);
nand U7483 (N_7483,N_6989,N_6745);
and U7484 (N_7484,N_6838,N_6893);
xor U7485 (N_7485,N_6828,N_6549);
or U7486 (N_7486,N_6536,N_6828);
nor U7487 (N_7487,N_6835,N_6649);
xnor U7488 (N_7488,N_6753,N_6932);
or U7489 (N_7489,N_6941,N_6771);
nor U7490 (N_7490,N_6878,N_6535);
nand U7491 (N_7491,N_6767,N_6599);
and U7492 (N_7492,N_6738,N_6829);
nand U7493 (N_7493,N_6543,N_6937);
or U7494 (N_7494,N_6736,N_6919);
or U7495 (N_7495,N_6881,N_6666);
xor U7496 (N_7496,N_6893,N_6954);
and U7497 (N_7497,N_6826,N_6997);
nand U7498 (N_7498,N_6981,N_6725);
nand U7499 (N_7499,N_6728,N_6575);
nand U7500 (N_7500,N_7105,N_7282);
nor U7501 (N_7501,N_7014,N_7439);
and U7502 (N_7502,N_7336,N_7353);
and U7503 (N_7503,N_7308,N_7498);
nand U7504 (N_7504,N_7421,N_7157);
or U7505 (N_7505,N_7447,N_7395);
xor U7506 (N_7506,N_7436,N_7495);
nor U7507 (N_7507,N_7010,N_7485);
or U7508 (N_7508,N_7231,N_7237);
nand U7509 (N_7509,N_7446,N_7479);
nand U7510 (N_7510,N_7420,N_7211);
nor U7511 (N_7511,N_7210,N_7468);
nor U7512 (N_7512,N_7108,N_7112);
or U7513 (N_7513,N_7104,N_7304);
xnor U7514 (N_7514,N_7118,N_7367);
nand U7515 (N_7515,N_7122,N_7141);
or U7516 (N_7516,N_7114,N_7250);
xnor U7517 (N_7517,N_7131,N_7084);
or U7518 (N_7518,N_7195,N_7351);
or U7519 (N_7519,N_7204,N_7324);
nor U7520 (N_7520,N_7275,N_7064);
or U7521 (N_7521,N_7368,N_7085);
nor U7522 (N_7522,N_7340,N_7228);
and U7523 (N_7523,N_7291,N_7068);
and U7524 (N_7524,N_7441,N_7080);
xor U7525 (N_7525,N_7355,N_7247);
xnor U7526 (N_7526,N_7425,N_7328);
nor U7527 (N_7527,N_7102,N_7057);
nor U7528 (N_7528,N_7238,N_7123);
xnor U7529 (N_7529,N_7369,N_7430);
nor U7530 (N_7530,N_7256,N_7482);
xnor U7531 (N_7531,N_7045,N_7161);
or U7532 (N_7532,N_7315,N_7071);
nand U7533 (N_7533,N_7026,N_7394);
nor U7534 (N_7534,N_7097,N_7410);
nor U7535 (N_7535,N_7134,N_7082);
and U7536 (N_7536,N_7263,N_7153);
nor U7537 (N_7537,N_7448,N_7246);
and U7538 (N_7538,N_7453,N_7329);
xnor U7539 (N_7539,N_7213,N_7138);
nand U7540 (N_7540,N_7005,N_7463);
nor U7541 (N_7541,N_7478,N_7489);
xor U7542 (N_7542,N_7345,N_7396);
or U7543 (N_7543,N_7036,N_7350);
or U7544 (N_7544,N_7307,N_7376);
nor U7545 (N_7545,N_7063,N_7229);
or U7546 (N_7546,N_7127,N_7059);
nor U7547 (N_7547,N_7265,N_7168);
nand U7548 (N_7548,N_7040,N_7389);
nor U7549 (N_7549,N_7381,N_7046);
nand U7550 (N_7550,N_7431,N_7303);
xnor U7551 (N_7551,N_7072,N_7144);
or U7552 (N_7552,N_7243,N_7332);
nand U7553 (N_7553,N_7067,N_7322);
nor U7554 (N_7554,N_7337,N_7320);
and U7555 (N_7555,N_7158,N_7013);
and U7556 (N_7556,N_7496,N_7470);
nor U7557 (N_7557,N_7272,N_7270);
nand U7558 (N_7558,N_7205,N_7370);
and U7559 (N_7559,N_7424,N_7075);
nand U7560 (N_7560,N_7401,N_7339);
nand U7561 (N_7561,N_7358,N_7499);
or U7562 (N_7562,N_7461,N_7148);
xor U7563 (N_7563,N_7186,N_7066);
or U7564 (N_7564,N_7288,N_7090);
and U7565 (N_7565,N_7312,N_7459);
xnor U7566 (N_7566,N_7306,N_7305);
or U7567 (N_7567,N_7255,N_7054);
nor U7568 (N_7568,N_7009,N_7083);
nand U7569 (N_7569,N_7091,N_7024);
nand U7570 (N_7570,N_7442,N_7217);
nor U7571 (N_7571,N_7294,N_7295);
and U7572 (N_7572,N_7034,N_7433);
nand U7573 (N_7573,N_7357,N_7239);
and U7574 (N_7574,N_7412,N_7208);
or U7575 (N_7575,N_7119,N_7454);
xor U7576 (N_7576,N_7146,N_7175);
and U7577 (N_7577,N_7223,N_7077);
and U7578 (N_7578,N_7343,N_7450);
nor U7579 (N_7579,N_7363,N_7260);
nand U7580 (N_7580,N_7487,N_7182);
nand U7581 (N_7581,N_7342,N_7098);
nand U7582 (N_7582,N_7230,N_7011);
nor U7583 (N_7583,N_7032,N_7474);
nand U7584 (N_7584,N_7361,N_7140);
xnor U7585 (N_7585,N_7379,N_7143);
nand U7586 (N_7586,N_7225,N_7375);
xnor U7587 (N_7587,N_7111,N_7006);
nor U7588 (N_7588,N_7429,N_7462);
and U7589 (N_7589,N_7422,N_7214);
nand U7590 (N_7590,N_7173,N_7188);
and U7591 (N_7591,N_7364,N_7299);
xor U7592 (N_7592,N_7321,N_7314);
xor U7593 (N_7593,N_7331,N_7047);
or U7594 (N_7594,N_7194,N_7289);
nand U7595 (N_7595,N_7458,N_7028);
and U7596 (N_7596,N_7497,N_7349);
nand U7597 (N_7597,N_7055,N_7050);
xor U7598 (N_7598,N_7016,N_7117);
and U7599 (N_7599,N_7488,N_7087);
nor U7600 (N_7600,N_7169,N_7440);
and U7601 (N_7601,N_7027,N_7100);
xnor U7602 (N_7602,N_7233,N_7124);
or U7603 (N_7603,N_7444,N_7346);
nor U7604 (N_7604,N_7391,N_7212);
nor U7605 (N_7605,N_7130,N_7192);
nand U7606 (N_7606,N_7224,N_7457);
nor U7607 (N_7607,N_7001,N_7177);
nand U7608 (N_7608,N_7409,N_7107);
or U7609 (N_7609,N_7252,N_7285);
xnor U7610 (N_7610,N_7387,N_7022);
or U7611 (N_7611,N_7044,N_7435);
and U7612 (N_7612,N_7018,N_7283);
and U7613 (N_7613,N_7008,N_7456);
or U7614 (N_7614,N_7003,N_7347);
nand U7615 (N_7615,N_7360,N_7215);
nor U7616 (N_7616,N_7033,N_7164);
or U7617 (N_7617,N_7202,N_7413);
and U7618 (N_7618,N_7133,N_7234);
or U7619 (N_7619,N_7327,N_7472);
xnor U7620 (N_7620,N_7354,N_7253);
and U7621 (N_7621,N_7103,N_7120);
or U7622 (N_7622,N_7019,N_7390);
nand U7623 (N_7623,N_7335,N_7060);
xnor U7624 (N_7624,N_7415,N_7382);
and U7625 (N_7625,N_7070,N_7172);
and U7626 (N_7626,N_7051,N_7196);
nand U7627 (N_7627,N_7065,N_7159);
xnor U7628 (N_7628,N_7061,N_7317);
and U7629 (N_7629,N_7235,N_7484);
nor U7630 (N_7630,N_7372,N_7128);
xor U7631 (N_7631,N_7414,N_7269);
and U7632 (N_7632,N_7388,N_7197);
and U7633 (N_7633,N_7284,N_7185);
xor U7634 (N_7634,N_7190,N_7418);
nor U7635 (N_7635,N_7226,N_7330);
nor U7636 (N_7636,N_7262,N_7281);
or U7637 (N_7637,N_7445,N_7416);
or U7638 (N_7638,N_7493,N_7467);
xor U7639 (N_7639,N_7030,N_7166);
or U7640 (N_7640,N_7203,N_7280);
xor U7641 (N_7641,N_7249,N_7222);
nand U7642 (N_7642,N_7469,N_7240);
nand U7643 (N_7643,N_7475,N_7135);
or U7644 (N_7644,N_7277,N_7058);
nand U7645 (N_7645,N_7121,N_7259);
and U7646 (N_7646,N_7311,N_7297);
nor U7647 (N_7647,N_7216,N_7298);
nor U7648 (N_7648,N_7261,N_7296);
nor U7649 (N_7649,N_7139,N_7145);
xnor U7650 (N_7650,N_7007,N_7244);
and U7651 (N_7651,N_7325,N_7359);
xor U7652 (N_7652,N_7113,N_7266);
or U7653 (N_7653,N_7397,N_7333);
and U7654 (N_7654,N_7126,N_7483);
nand U7655 (N_7655,N_7073,N_7428);
nor U7656 (N_7656,N_7000,N_7081);
nand U7657 (N_7657,N_7076,N_7242);
nand U7658 (N_7658,N_7257,N_7180);
nor U7659 (N_7659,N_7227,N_7417);
nand U7660 (N_7660,N_7356,N_7096);
or U7661 (N_7661,N_7344,N_7089);
xor U7662 (N_7662,N_7200,N_7116);
nand U7663 (N_7663,N_7452,N_7432);
nor U7664 (N_7664,N_7163,N_7110);
or U7665 (N_7665,N_7207,N_7268);
xor U7666 (N_7666,N_7136,N_7362);
nand U7667 (N_7667,N_7017,N_7221);
or U7668 (N_7668,N_7206,N_7151);
nor U7669 (N_7669,N_7443,N_7251);
nand U7670 (N_7670,N_7167,N_7012);
and U7671 (N_7671,N_7301,N_7209);
xor U7672 (N_7672,N_7385,N_7147);
or U7673 (N_7673,N_7095,N_7399);
nor U7674 (N_7674,N_7309,N_7160);
or U7675 (N_7675,N_7092,N_7101);
and U7676 (N_7676,N_7155,N_7366);
nand U7677 (N_7677,N_7002,N_7174);
nor U7678 (N_7678,N_7189,N_7201);
nor U7679 (N_7679,N_7302,N_7142);
xnor U7680 (N_7680,N_7094,N_7115);
nor U7681 (N_7681,N_7481,N_7198);
nor U7682 (N_7682,N_7464,N_7193);
and U7683 (N_7683,N_7220,N_7150);
nand U7684 (N_7684,N_7245,N_7403);
or U7685 (N_7685,N_7029,N_7477);
nor U7686 (N_7686,N_7181,N_7035);
nand U7687 (N_7687,N_7020,N_7053);
and U7688 (N_7688,N_7373,N_7025);
and U7689 (N_7689,N_7313,N_7348);
nand U7690 (N_7690,N_7406,N_7393);
xnor U7691 (N_7691,N_7377,N_7079);
and U7692 (N_7692,N_7264,N_7310);
or U7693 (N_7693,N_7438,N_7316);
nand U7694 (N_7694,N_7038,N_7405);
or U7695 (N_7695,N_7383,N_7183);
nor U7696 (N_7696,N_7088,N_7292);
nand U7697 (N_7697,N_7179,N_7187);
nand U7698 (N_7698,N_7279,N_7274);
xnor U7699 (N_7699,N_7241,N_7232);
or U7700 (N_7700,N_7052,N_7041);
and U7701 (N_7701,N_7062,N_7476);
and U7702 (N_7702,N_7300,N_7352);
nor U7703 (N_7703,N_7437,N_7184);
and U7704 (N_7704,N_7293,N_7248);
nand U7705 (N_7705,N_7460,N_7392);
or U7706 (N_7706,N_7049,N_7434);
or U7707 (N_7707,N_7219,N_7465);
xor U7708 (N_7708,N_7491,N_7191);
xnor U7709 (N_7709,N_7466,N_7323);
nor U7710 (N_7710,N_7176,N_7093);
or U7711 (N_7711,N_7318,N_7109);
or U7712 (N_7712,N_7154,N_7426);
or U7713 (N_7713,N_7099,N_7170);
nor U7714 (N_7714,N_7402,N_7129);
nand U7715 (N_7715,N_7199,N_7037);
nand U7716 (N_7716,N_7334,N_7031);
or U7717 (N_7717,N_7069,N_7152);
xnor U7718 (N_7718,N_7236,N_7449);
nand U7719 (N_7719,N_7162,N_7384);
nor U7720 (N_7720,N_7286,N_7451);
or U7721 (N_7721,N_7125,N_7290);
nor U7722 (N_7722,N_7149,N_7043);
and U7723 (N_7723,N_7380,N_7423);
and U7724 (N_7724,N_7374,N_7386);
nor U7725 (N_7725,N_7106,N_7015);
xnor U7726 (N_7726,N_7048,N_7039);
nor U7727 (N_7727,N_7455,N_7056);
or U7728 (N_7728,N_7004,N_7378);
xnor U7729 (N_7729,N_7074,N_7398);
nor U7730 (N_7730,N_7419,N_7427);
or U7731 (N_7731,N_7400,N_7341);
nand U7732 (N_7732,N_7254,N_7165);
xor U7733 (N_7733,N_7480,N_7486);
xnor U7734 (N_7734,N_7276,N_7492);
nand U7735 (N_7735,N_7326,N_7023);
and U7736 (N_7736,N_7267,N_7258);
nand U7737 (N_7737,N_7365,N_7086);
or U7738 (N_7738,N_7137,N_7042);
or U7739 (N_7739,N_7319,N_7021);
and U7740 (N_7740,N_7411,N_7407);
xnor U7741 (N_7741,N_7171,N_7132);
nand U7742 (N_7742,N_7408,N_7338);
xnor U7743 (N_7743,N_7473,N_7371);
nand U7744 (N_7744,N_7218,N_7178);
nor U7745 (N_7745,N_7471,N_7078);
xor U7746 (N_7746,N_7404,N_7490);
nand U7747 (N_7747,N_7278,N_7287);
nand U7748 (N_7748,N_7273,N_7271);
nand U7749 (N_7749,N_7156,N_7494);
and U7750 (N_7750,N_7144,N_7289);
nor U7751 (N_7751,N_7234,N_7460);
and U7752 (N_7752,N_7369,N_7240);
nor U7753 (N_7753,N_7103,N_7404);
xor U7754 (N_7754,N_7331,N_7119);
and U7755 (N_7755,N_7257,N_7156);
xor U7756 (N_7756,N_7300,N_7046);
or U7757 (N_7757,N_7131,N_7499);
or U7758 (N_7758,N_7088,N_7068);
nand U7759 (N_7759,N_7498,N_7005);
xnor U7760 (N_7760,N_7258,N_7147);
and U7761 (N_7761,N_7115,N_7065);
or U7762 (N_7762,N_7003,N_7302);
and U7763 (N_7763,N_7015,N_7084);
nand U7764 (N_7764,N_7499,N_7493);
xor U7765 (N_7765,N_7430,N_7417);
nor U7766 (N_7766,N_7194,N_7033);
nand U7767 (N_7767,N_7454,N_7010);
xor U7768 (N_7768,N_7035,N_7028);
or U7769 (N_7769,N_7130,N_7258);
nand U7770 (N_7770,N_7190,N_7117);
nor U7771 (N_7771,N_7312,N_7352);
and U7772 (N_7772,N_7433,N_7434);
nand U7773 (N_7773,N_7063,N_7064);
xor U7774 (N_7774,N_7400,N_7468);
and U7775 (N_7775,N_7320,N_7336);
and U7776 (N_7776,N_7417,N_7344);
nor U7777 (N_7777,N_7356,N_7316);
or U7778 (N_7778,N_7410,N_7308);
xor U7779 (N_7779,N_7011,N_7199);
or U7780 (N_7780,N_7147,N_7397);
nand U7781 (N_7781,N_7453,N_7377);
and U7782 (N_7782,N_7220,N_7273);
xnor U7783 (N_7783,N_7350,N_7268);
nor U7784 (N_7784,N_7031,N_7317);
nor U7785 (N_7785,N_7412,N_7359);
and U7786 (N_7786,N_7290,N_7133);
xnor U7787 (N_7787,N_7026,N_7457);
nand U7788 (N_7788,N_7327,N_7499);
and U7789 (N_7789,N_7037,N_7315);
xnor U7790 (N_7790,N_7181,N_7280);
nor U7791 (N_7791,N_7114,N_7408);
or U7792 (N_7792,N_7221,N_7215);
nor U7793 (N_7793,N_7378,N_7122);
and U7794 (N_7794,N_7062,N_7447);
nand U7795 (N_7795,N_7075,N_7338);
xnor U7796 (N_7796,N_7480,N_7024);
nor U7797 (N_7797,N_7147,N_7474);
or U7798 (N_7798,N_7417,N_7483);
nand U7799 (N_7799,N_7001,N_7348);
xnor U7800 (N_7800,N_7145,N_7488);
and U7801 (N_7801,N_7375,N_7164);
and U7802 (N_7802,N_7090,N_7433);
and U7803 (N_7803,N_7444,N_7082);
nor U7804 (N_7804,N_7307,N_7140);
or U7805 (N_7805,N_7215,N_7419);
xor U7806 (N_7806,N_7153,N_7018);
or U7807 (N_7807,N_7159,N_7272);
xnor U7808 (N_7808,N_7453,N_7472);
nor U7809 (N_7809,N_7310,N_7250);
or U7810 (N_7810,N_7304,N_7382);
xor U7811 (N_7811,N_7260,N_7383);
xnor U7812 (N_7812,N_7101,N_7399);
and U7813 (N_7813,N_7240,N_7178);
nand U7814 (N_7814,N_7240,N_7288);
or U7815 (N_7815,N_7090,N_7151);
and U7816 (N_7816,N_7434,N_7289);
and U7817 (N_7817,N_7485,N_7025);
or U7818 (N_7818,N_7306,N_7244);
xor U7819 (N_7819,N_7294,N_7429);
nand U7820 (N_7820,N_7151,N_7493);
nor U7821 (N_7821,N_7381,N_7009);
xnor U7822 (N_7822,N_7128,N_7065);
xor U7823 (N_7823,N_7037,N_7253);
nor U7824 (N_7824,N_7220,N_7328);
xnor U7825 (N_7825,N_7172,N_7440);
nand U7826 (N_7826,N_7110,N_7469);
nand U7827 (N_7827,N_7269,N_7218);
nand U7828 (N_7828,N_7499,N_7289);
and U7829 (N_7829,N_7433,N_7304);
and U7830 (N_7830,N_7173,N_7217);
and U7831 (N_7831,N_7056,N_7298);
nand U7832 (N_7832,N_7013,N_7182);
and U7833 (N_7833,N_7095,N_7051);
nor U7834 (N_7834,N_7062,N_7418);
or U7835 (N_7835,N_7402,N_7421);
xor U7836 (N_7836,N_7493,N_7047);
or U7837 (N_7837,N_7127,N_7254);
or U7838 (N_7838,N_7489,N_7365);
nor U7839 (N_7839,N_7252,N_7383);
xnor U7840 (N_7840,N_7312,N_7292);
and U7841 (N_7841,N_7272,N_7256);
and U7842 (N_7842,N_7435,N_7318);
and U7843 (N_7843,N_7399,N_7076);
nand U7844 (N_7844,N_7032,N_7210);
or U7845 (N_7845,N_7142,N_7393);
xnor U7846 (N_7846,N_7011,N_7137);
nand U7847 (N_7847,N_7041,N_7263);
and U7848 (N_7848,N_7190,N_7385);
xnor U7849 (N_7849,N_7398,N_7019);
or U7850 (N_7850,N_7447,N_7263);
nand U7851 (N_7851,N_7142,N_7263);
xnor U7852 (N_7852,N_7186,N_7052);
nor U7853 (N_7853,N_7464,N_7023);
nor U7854 (N_7854,N_7346,N_7316);
or U7855 (N_7855,N_7022,N_7458);
xnor U7856 (N_7856,N_7272,N_7171);
and U7857 (N_7857,N_7412,N_7211);
xor U7858 (N_7858,N_7350,N_7389);
nor U7859 (N_7859,N_7077,N_7238);
xor U7860 (N_7860,N_7387,N_7196);
nor U7861 (N_7861,N_7125,N_7491);
nand U7862 (N_7862,N_7307,N_7207);
and U7863 (N_7863,N_7011,N_7271);
and U7864 (N_7864,N_7185,N_7404);
nor U7865 (N_7865,N_7294,N_7109);
nor U7866 (N_7866,N_7461,N_7330);
nor U7867 (N_7867,N_7163,N_7492);
or U7868 (N_7868,N_7031,N_7439);
xor U7869 (N_7869,N_7041,N_7476);
and U7870 (N_7870,N_7071,N_7482);
or U7871 (N_7871,N_7413,N_7016);
or U7872 (N_7872,N_7411,N_7104);
nor U7873 (N_7873,N_7053,N_7493);
nand U7874 (N_7874,N_7088,N_7017);
and U7875 (N_7875,N_7437,N_7118);
nand U7876 (N_7876,N_7153,N_7231);
and U7877 (N_7877,N_7046,N_7404);
nor U7878 (N_7878,N_7104,N_7313);
nor U7879 (N_7879,N_7236,N_7092);
nor U7880 (N_7880,N_7191,N_7207);
or U7881 (N_7881,N_7298,N_7459);
and U7882 (N_7882,N_7281,N_7265);
nor U7883 (N_7883,N_7118,N_7349);
xnor U7884 (N_7884,N_7285,N_7374);
xnor U7885 (N_7885,N_7474,N_7343);
nor U7886 (N_7886,N_7080,N_7410);
nor U7887 (N_7887,N_7161,N_7496);
nor U7888 (N_7888,N_7086,N_7482);
xnor U7889 (N_7889,N_7261,N_7382);
nand U7890 (N_7890,N_7223,N_7382);
nand U7891 (N_7891,N_7474,N_7244);
nor U7892 (N_7892,N_7251,N_7417);
nand U7893 (N_7893,N_7283,N_7417);
or U7894 (N_7894,N_7361,N_7292);
nor U7895 (N_7895,N_7467,N_7040);
nand U7896 (N_7896,N_7193,N_7194);
xor U7897 (N_7897,N_7383,N_7466);
nor U7898 (N_7898,N_7065,N_7147);
xor U7899 (N_7899,N_7202,N_7240);
xor U7900 (N_7900,N_7347,N_7183);
and U7901 (N_7901,N_7164,N_7396);
xnor U7902 (N_7902,N_7333,N_7206);
nor U7903 (N_7903,N_7184,N_7343);
nor U7904 (N_7904,N_7441,N_7195);
and U7905 (N_7905,N_7029,N_7411);
and U7906 (N_7906,N_7057,N_7159);
and U7907 (N_7907,N_7134,N_7307);
nor U7908 (N_7908,N_7403,N_7213);
nor U7909 (N_7909,N_7200,N_7294);
xnor U7910 (N_7910,N_7269,N_7261);
and U7911 (N_7911,N_7182,N_7169);
xnor U7912 (N_7912,N_7345,N_7182);
and U7913 (N_7913,N_7085,N_7425);
or U7914 (N_7914,N_7273,N_7345);
xor U7915 (N_7915,N_7029,N_7233);
or U7916 (N_7916,N_7466,N_7441);
xnor U7917 (N_7917,N_7071,N_7393);
nor U7918 (N_7918,N_7358,N_7223);
nor U7919 (N_7919,N_7457,N_7267);
xnor U7920 (N_7920,N_7065,N_7006);
nor U7921 (N_7921,N_7198,N_7050);
xor U7922 (N_7922,N_7086,N_7019);
or U7923 (N_7923,N_7170,N_7127);
or U7924 (N_7924,N_7257,N_7301);
and U7925 (N_7925,N_7367,N_7374);
nand U7926 (N_7926,N_7102,N_7167);
and U7927 (N_7927,N_7070,N_7314);
nand U7928 (N_7928,N_7325,N_7431);
or U7929 (N_7929,N_7403,N_7393);
or U7930 (N_7930,N_7464,N_7440);
and U7931 (N_7931,N_7126,N_7352);
xnor U7932 (N_7932,N_7089,N_7021);
xor U7933 (N_7933,N_7203,N_7417);
and U7934 (N_7934,N_7119,N_7304);
or U7935 (N_7935,N_7487,N_7448);
nor U7936 (N_7936,N_7047,N_7319);
nor U7937 (N_7937,N_7053,N_7478);
nand U7938 (N_7938,N_7346,N_7020);
or U7939 (N_7939,N_7215,N_7090);
nand U7940 (N_7940,N_7328,N_7350);
xor U7941 (N_7941,N_7016,N_7069);
and U7942 (N_7942,N_7457,N_7023);
nor U7943 (N_7943,N_7476,N_7036);
and U7944 (N_7944,N_7196,N_7140);
xnor U7945 (N_7945,N_7451,N_7426);
xor U7946 (N_7946,N_7397,N_7269);
nand U7947 (N_7947,N_7086,N_7493);
xnor U7948 (N_7948,N_7482,N_7026);
nor U7949 (N_7949,N_7015,N_7097);
or U7950 (N_7950,N_7253,N_7441);
nor U7951 (N_7951,N_7316,N_7385);
xor U7952 (N_7952,N_7194,N_7024);
nand U7953 (N_7953,N_7207,N_7122);
nor U7954 (N_7954,N_7234,N_7421);
or U7955 (N_7955,N_7234,N_7409);
nand U7956 (N_7956,N_7018,N_7013);
nor U7957 (N_7957,N_7494,N_7142);
nor U7958 (N_7958,N_7137,N_7417);
xor U7959 (N_7959,N_7088,N_7066);
xor U7960 (N_7960,N_7160,N_7433);
xnor U7961 (N_7961,N_7414,N_7423);
or U7962 (N_7962,N_7184,N_7120);
and U7963 (N_7963,N_7233,N_7178);
or U7964 (N_7964,N_7127,N_7140);
xor U7965 (N_7965,N_7171,N_7308);
nor U7966 (N_7966,N_7351,N_7180);
nor U7967 (N_7967,N_7347,N_7329);
and U7968 (N_7968,N_7431,N_7052);
nand U7969 (N_7969,N_7159,N_7137);
xor U7970 (N_7970,N_7252,N_7262);
or U7971 (N_7971,N_7359,N_7482);
xnor U7972 (N_7972,N_7378,N_7351);
xor U7973 (N_7973,N_7366,N_7282);
or U7974 (N_7974,N_7389,N_7050);
nand U7975 (N_7975,N_7247,N_7457);
nor U7976 (N_7976,N_7077,N_7131);
nand U7977 (N_7977,N_7268,N_7449);
nand U7978 (N_7978,N_7429,N_7377);
or U7979 (N_7979,N_7436,N_7017);
or U7980 (N_7980,N_7340,N_7078);
xnor U7981 (N_7981,N_7191,N_7230);
nand U7982 (N_7982,N_7412,N_7461);
and U7983 (N_7983,N_7109,N_7381);
nand U7984 (N_7984,N_7091,N_7447);
nand U7985 (N_7985,N_7208,N_7291);
or U7986 (N_7986,N_7476,N_7104);
or U7987 (N_7987,N_7466,N_7186);
nand U7988 (N_7988,N_7298,N_7136);
nor U7989 (N_7989,N_7116,N_7142);
or U7990 (N_7990,N_7021,N_7022);
and U7991 (N_7991,N_7445,N_7028);
nand U7992 (N_7992,N_7423,N_7112);
or U7993 (N_7993,N_7203,N_7100);
or U7994 (N_7994,N_7150,N_7425);
and U7995 (N_7995,N_7047,N_7221);
nand U7996 (N_7996,N_7304,N_7373);
and U7997 (N_7997,N_7384,N_7250);
or U7998 (N_7998,N_7460,N_7048);
xnor U7999 (N_7999,N_7175,N_7027);
or U8000 (N_8000,N_7575,N_7977);
nand U8001 (N_8001,N_7634,N_7723);
and U8002 (N_8002,N_7798,N_7815);
xnor U8003 (N_8003,N_7651,N_7691);
nand U8004 (N_8004,N_7900,N_7533);
or U8005 (N_8005,N_7629,N_7732);
xor U8006 (N_8006,N_7992,N_7585);
xor U8007 (N_8007,N_7853,N_7554);
nor U8008 (N_8008,N_7694,N_7521);
or U8009 (N_8009,N_7983,N_7705);
and U8010 (N_8010,N_7539,N_7903);
nand U8011 (N_8011,N_7702,N_7614);
and U8012 (N_8012,N_7590,N_7657);
and U8013 (N_8013,N_7734,N_7846);
nor U8014 (N_8014,N_7699,N_7701);
xnor U8015 (N_8015,N_7787,N_7932);
xor U8016 (N_8016,N_7564,N_7746);
or U8017 (N_8017,N_7872,N_7592);
and U8018 (N_8018,N_7529,N_7631);
and U8019 (N_8019,N_7973,N_7678);
xor U8020 (N_8020,N_7580,N_7781);
or U8021 (N_8021,N_7530,N_7740);
nor U8022 (N_8022,N_7837,N_7537);
or U8023 (N_8023,N_7961,N_7532);
and U8024 (N_8024,N_7658,N_7712);
or U8025 (N_8025,N_7984,N_7777);
xor U8026 (N_8026,N_7510,N_7996);
nor U8027 (N_8027,N_7736,N_7639);
or U8028 (N_8028,N_7671,N_7560);
or U8029 (N_8029,N_7820,N_7758);
or U8030 (N_8030,N_7790,N_7550);
or U8031 (N_8031,N_7951,N_7504);
or U8032 (N_8032,N_7928,N_7827);
nand U8033 (N_8033,N_7733,N_7954);
nor U8034 (N_8034,N_7659,N_7735);
xor U8035 (N_8035,N_7764,N_7591);
nor U8036 (N_8036,N_7674,N_7909);
and U8037 (N_8037,N_7782,N_7826);
and U8038 (N_8038,N_7524,N_7690);
xnor U8039 (N_8039,N_7942,N_7599);
nor U8040 (N_8040,N_7601,N_7650);
xnor U8041 (N_8041,N_7817,N_7958);
and U8042 (N_8042,N_7507,N_7776);
nor U8043 (N_8043,N_7930,N_7627);
and U8044 (N_8044,N_7636,N_7774);
nand U8045 (N_8045,N_7654,N_7881);
nor U8046 (N_8046,N_7664,N_7514);
nor U8047 (N_8047,N_7578,N_7802);
nor U8048 (N_8048,N_7948,N_7588);
or U8049 (N_8049,N_7834,N_7784);
or U8050 (N_8050,N_7613,N_7512);
nand U8051 (N_8051,N_7933,N_7797);
xor U8052 (N_8052,N_7552,N_7811);
and U8053 (N_8053,N_7675,N_7718);
or U8054 (N_8054,N_7878,N_7898);
or U8055 (N_8055,N_7786,N_7936);
nand U8056 (N_8056,N_7813,N_7663);
nand U8057 (N_8057,N_7891,N_7848);
or U8058 (N_8058,N_7941,N_7644);
nor U8059 (N_8059,N_7757,N_7828);
nand U8060 (N_8060,N_7637,N_7794);
or U8061 (N_8061,N_7950,N_7756);
nor U8062 (N_8062,N_7804,N_7576);
nor U8063 (N_8063,N_7994,N_7693);
and U8064 (N_8064,N_7688,N_7840);
nand U8065 (N_8065,N_7628,N_7752);
or U8066 (N_8066,N_7921,N_7750);
xor U8067 (N_8067,N_7621,N_7880);
nor U8068 (N_8068,N_7569,N_7582);
or U8069 (N_8069,N_7581,N_7511);
and U8070 (N_8070,N_7976,N_7742);
or U8071 (N_8071,N_7667,N_7715);
or U8072 (N_8072,N_7971,N_7847);
xnor U8073 (N_8073,N_7687,N_7632);
and U8074 (N_8074,N_7801,N_7761);
nand U8075 (N_8075,N_7868,N_7620);
and U8076 (N_8076,N_7913,N_7985);
xor U8077 (N_8077,N_7818,N_7656);
and U8078 (N_8078,N_7616,N_7940);
and U8079 (N_8079,N_7653,N_7907);
and U8080 (N_8080,N_7630,N_7871);
nand U8081 (N_8081,N_7624,N_7584);
nand U8082 (N_8082,N_7684,N_7540);
and U8083 (N_8083,N_7517,N_7759);
nand U8084 (N_8084,N_7548,N_7743);
and U8085 (N_8085,N_7589,N_7819);
or U8086 (N_8086,N_7549,N_7830);
and U8087 (N_8087,N_7566,N_7643);
and U8088 (N_8088,N_7987,N_7775);
and U8089 (N_8089,N_7768,N_7875);
or U8090 (N_8090,N_7547,N_7997);
and U8091 (N_8091,N_7905,N_7860);
or U8092 (N_8092,N_7763,N_7812);
or U8093 (N_8093,N_7720,N_7660);
xor U8094 (N_8094,N_7896,N_7852);
nor U8095 (N_8095,N_7672,N_7755);
xnor U8096 (N_8096,N_7882,N_7574);
xnor U8097 (N_8097,N_7648,N_7666);
nand U8098 (N_8098,N_7854,N_7642);
and U8099 (N_8099,N_7841,N_7518);
or U8100 (N_8100,N_7908,N_7717);
or U8101 (N_8101,N_7760,N_7595);
nor U8102 (N_8102,N_7865,N_7778);
nor U8103 (N_8103,N_7914,N_7683);
xor U8104 (N_8104,N_7978,N_7993);
nor U8105 (N_8105,N_7970,N_7986);
and U8106 (N_8106,N_7710,N_7615);
nand U8107 (N_8107,N_7806,N_7894);
and U8108 (N_8108,N_7551,N_7893);
nand U8109 (N_8109,N_7945,N_7528);
nor U8110 (N_8110,N_7682,N_7968);
nor U8111 (N_8111,N_7886,N_7836);
nor U8112 (N_8112,N_7638,N_7522);
and U8113 (N_8113,N_7623,N_7887);
or U8114 (N_8114,N_7889,N_7707);
xnor U8115 (N_8115,N_7570,N_7737);
and U8116 (N_8116,N_7857,N_7824);
or U8117 (N_8117,N_7649,N_7525);
nor U8118 (N_8118,N_7662,N_7708);
xnor U8119 (N_8119,N_7618,N_7668);
nand U8120 (N_8120,N_7888,N_7706);
or U8121 (N_8121,N_7747,N_7519);
and U8122 (N_8122,N_7803,N_7696);
or U8123 (N_8123,N_7527,N_7714);
or U8124 (N_8124,N_7845,N_7739);
nor U8125 (N_8125,N_7625,N_7929);
nand U8126 (N_8126,N_7679,N_7609);
nor U8127 (N_8127,N_7677,N_7729);
and U8128 (N_8128,N_7711,N_7766);
and U8129 (N_8129,N_7633,N_7937);
and U8130 (N_8130,N_7995,N_7593);
xnor U8131 (N_8131,N_7587,N_7922);
xnor U8132 (N_8132,N_7859,N_7622);
nor U8133 (N_8133,N_7738,N_7920);
and U8134 (N_8134,N_7681,N_7829);
or U8135 (N_8135,N_7831,N_7918);
nand U8136 (N_8136,N_7669,N_7698);
and U8137 (N_8137,N_7953,N_7655);
nand U8138 (N_8138,N_7923,N_7748);
xor U8139 (N_8139,N_7981,N_7538);
and U8140 (N_8140,N_7769,N_7912);
and U8141 (N_8141,N_7573,N_7509);
nand U8142 (N_8142,N_7611,N_7899);
and U8143 (N_8143,N_7725,N_7884);
xnor U8144 (N_8144,N_7716,N_7562);
nor U8145 (N_8145,N_7925,N_7862);
and U8146 (N_8146,N_7814,N_7979);
xnor U8147 (N_8147,N_7988,N_7944);
nand U8148 (N_8148,N_7980,N_7572);
nor U8149 (N_8149,N_7544,N_7788);
or U8150 (N_8150,N_7500,N_7861);
nor U8151 (N_8151,N_7858,N_7741);
nor U8152 (N_8152,N_7646,N_7640);
and U8153 (N_8153,N_7598,N_7885);
or U8154 (N_8154,N_7559,N_7565);
or U8155 (N_8155,N_7919,N_7515);
and U8156 (N_8156,N_7608,N_7523);
or U8157 (N_8157,N_7876,N_7526);
or U8158 (N_8158,N_7771,N_7571);
or U8159 (N_8159,N_7943,N_7603);
and U8160 (N_8160,N_7703,N_7610);
xnor U8161 (N_8161,N_7753,N_7892);
nor U8162 (N_8162,N_7809,N_7821);
xor U8163 (N_8163,N_7982,N_7520);
or U8164 (N_8164,N_7835,N_7805);
nand U8165 (N_8165,N_7879,N_7931);
xnor U8166 (N_8166,N_7842,N_7935);
xnor U8167 (N_8167,N_7939,N_7780);
or U8168 (N_8168,N_7967,N_7901);
and U8169 (N_8169,N_7851,N_7779);
or U8170 (N_8170,N_7721,N_7567);
nand U8171 (N_8171,N_7745,N_7545);
xnor U8172 (N_8172,N_7989,N_7904);
and U8173 (N_8173,N_7676,N_7765);
nor U8174 (N_8174,N_7700,N_7906);
xor U8175 (N_8175,N_7536,N_7555);
nor U8176 (N_8176,N_7999,N_7917);
nor U8177 (N_8177,N_7762,N_7534);
nor U8178 (N_8178,N_7863,N_7955);
xor U8179 (N_8179,N_7607,N_7849);
xnor U8180 (N_8180,N_7516,N_7531);
nand U8181 (N_8181,N_7974,N_7619);
xor U8182 (N_8182,N_7969,N_7855);
xor U8183 (N_8183,N_7927,N_7506);
xnor U8184 (N_8184,N_7807,N_7785);
xnor U8185 (N_8185,N_7513,N_7946);
and U8186 (N_8186,N_7661,N_7800);
and U8187 (N_8187,N_7825,N_7724);
or U8188 (N_8188,N_7645,N_7652);
xnor U8189 (N_8189,N_7924,N_7586);
xor U8190 (N_8190,N_7895,N_7641);
nor U8191 (N_8191,N_7543,N_7966);
nor U8192 (N_8192,N_7686,N_7874);
or U8193 (N_8193,N_7568,N_7556);
or U8194 (N_8194,N_7727,N_7704);
nor U8195 (N_8195,N_7685,N_7956);
and U8196 (N_8196,N_7563,N_7843);
xor U8197 (N_8197,N_7990,N_7728);
nor U8198 (N_8198,N_7867,N_7998);
and U8199 (N_8199,N_7810,N_7902);
or U8200 (N_8200,N_7502,N_7557);
and U8201 (N_8201,N_7934,N_7952);
and U8202 (N_8202,N_7938,N_7612);
xnor U8203 (N_8203,N_7647,N_7635);
xnor U8204 (N_8204,N_7796,N_7719);
nand U8205 (N_8205,N_7960,N_7561);
nand U8206 (N_8206,N_7816,N_7697);
and U8207 (N_8207,N_7542,N_7577);
and U8208 (N_8208,N_7808,N_7505);
nor U8209 (N_8209,N_7709,N_7838);
and U8210 (N_8210,N_7503,N_7910);
nand U8211 (N_8211,N_7673,N_7689);
xnor U8212 (N_8212,N_7926,N_7770);
or U8213 (N_8213,N_7680,N_7692);
xnor U8214 (N_8214,N_7916,N_7864);
and U8215 (N_8215,N_7832,N_7964);
nand U8216 (N_8216,N_7963,N_7959);
nand U8217 (N_8217,N_7722,N_7626);
and U8218 (N_8218,N_7597,N_7546);
nor U8219 (N_8219,N_7911,N_7957);
nand U8220 (N_8220,N_7594,N_7749);
nand U8221 (N_8221,N_7877,N_7866);
nand U8222 (N_8222,N_7744,N_7856);
nor U8223 (N_8223,N_7870,N_7604);
or U8224 (N_8224,N_7713,N_7869);
nand U8225 (N_8225,N_7823,N_7972);
nor U8226 (N_8226,N_7795,N_7890);
and U8227 (N_8227,N_7670,N_7949);
nor U8228 (N_8228,N_7541,N_7789);
xor U8229 (N_8229,N_7839,N_7754);
or U8230 (N_8230,N_7773,N_7726);
and U8231 (N_8231,N_7844,N_7600);
and U8232 (N_8232,N_7799,N_7731);
nand U8233 (N_8233,N_7772,N_7553);
nor U8234 (N_8234,N_7617,N_7915);
nor U8235 (N_8235,N_7730,N_7579);
and U8236 (N_8236,N_7947,N_7873);
nor U8237 (N_8237,N_7558,N_7962);
or U8238 (N_8238,N_7822,N_7606);
or U8239 (N_8239,N_7783,N_7695);
or U8240 (N_8240,N_7897,N_7991);
xnor U8241 (N_8241,N_7792,N_7751);
xnor U8242 (N_8242,N_7975,N_7965);
xor U8243 (N_8243,N_7605,N_7791);
or U8244 (N_8244,N_7583,N_7501);
nand U8245 (N_8245,N_7883,N_7767);
nor U8246 (N_8246,N_7535,N_7850);
and U8247 (N_8247,N_7665,N_7602);
nand U8248 (N_8248,N_7833,N_7596);
and U8249 (N_8249,N_7793,N_7508);
or U8250 (N_8250,N_7610,N_7572);
nand U8251 (N_8251,N_7538,N_7576);
nand U8252 (N_8252,N_7945,N_7626);
or U8253 (N_8253,N_7904,N_7523);
nand U8254 (N_8254,N_7521,N_7555);
nand U8255 (N_8255,N_7802,N_7852);
xnor U8256 (N_8256,N_7688,N_7884);
and U8257 (N_8257,N_7725,N_7760);
nand U8258 (N_8258,N_7789,N_7559);
nor U8259 (N_8259,N_7692,N_7534);
nand U8260 (N_8260,N_7507,N_7616);
xnor U8261 (N_8261,N_7991,N_7639);
nor U8262 (N_8262,N_7650,N_7945);
xnor U8263 (N_8263,N_7747,N_7848);
and U8264 (N_8264,N_7525,N_7726);
xor U8265 (N_8265,N_7821,N_7624);
and U8266 (N_8266,N_7862,N_7743);
xor U8267 (N_8267,N_7996,N_7799);
and U8268 (N_8268,N_7593,N_7936);
xor U8269 (N_8269,N_7851,N_7875);
or U8270 (N_8270,N_7807,N_7990);
and U8271 (N_8271,N_7645,N_7700);
nor U8272 (N_8272,N_7508,N_7951);
and U8273 (N_8273,N_7831,N_7742);
nand U8274 (N_8274,N_7870,N_7653);
and U8275 (N_8275,N_7696,N_7911);
and U8276 (N_8276,N_7749,N_7741);
xnor U8277 (N_8277,N_7620,N_7723);
nand U8278 (N_8278,N_7538,N_7531);
nand U8279 (N_8279,N_7931,N_7921);
nand U8280 (N_8280,N_7922,N_7996);
or U8281 (N_8281,N_7923,N_7659);
nand U8282 (N_8282,N_7876,N_7758);
nand U8283 (N_8283,N_7687,N_7766);
and U8284 (N_8284,N_7837,N_7636);
and U8285 (N_8285,N_7579,N_7510);
and U8286 (N_8286,N_7547,N_7808);
xor U8287 (N_8287,N_7730,N_7914);
or U8288 (N_8288,N_7995,N_7976);
nand U8289 (N_8289,N_7595,N_7822);
nand U8290 (N_8290,N_7645,N_7511);
and U8291 (N_8291,N_7981,N_7529);
xnor U8292 (N_8292,N_7721,N_7510);
nand U8293 (N_8293,N_7543,N_7625);
nor U8294 (N_8294,N_7831,N_7605);
and U8295 (N_8295,N_7567,N_7859);
and U8296 (N_8296,N_7643,N_7572);
xor U8297 (N_8297,N_7628,N_7787);
and U8298 (N_8298,N_7965,N_7681);
or U8299 (N_8299,N_7900,N_7876);
nor U8300 (N_8300,N_7902,N_7527);
or U8301 (N_8301,N_7778,N_7940);
nand U8302 (N_8302,N_7802,N_7572);
nand U8303 (N_8303,N_7846,N_7909);
xor U8304 (N_8304,N_7811,N_7874);
nor U8305 (N_8305,N_7527,N_7694);
or U8306 (N_8306,N_7510,N_7979);
and U8307 (N_8307,N_7641,N_7947);
or U8308 (N_8308,N_7709,N_7743);
and U8309 (N_8309,N_7956,N_7737);
nand U8310 (N_8310,N_7960,N_7891);
nand U8311 (N_8311,N_7797,N_7771);
nand U8312 (N_8312,N_7594,N_7797);
nand U8313 (N_8313,N_7923,N_7707);
nand U8314 (N_8314,N_7653,N_7595);
xnor U8315 (N_8315,N_7750,N_7511);
nand U8316 (N_8316,N_7722,N_7650);
nor U8317 (N_8317,N_7976,N_7792);
and U8318 (N_8318,N_7668,N_7995);
nor U8319 (N_8319,N_7736,N_7712);
or U8320 (N_8320,N_7751,N_7513);
nor U8321 (N_8321,N_7570,N_7909);
nor U8322 (N_8322,N_7729,N_7823);
or U8323 (N_8323,N_7609,N_7795);
nor U8324 (N_8324,N_7571,N_7971);
xor U8325 (N_8325,N_7521,N_7949);
xnor U8326 (N_8326,N_7764,N_7740);
and U8327 (N_8327,N_7955,N_7609);
xnor U8328 (N_8328,N_7993,N_7620);
and U8329 (N_8329,N_7510,N_7665);
or U8330 (N_8330,N_7928,N_7962);
xnor U8331 (N_8331,N_7934,N_7625);
nor U8332 (N_8332,N_7986,N_7993);
nand U8333 (N_8333,N_7895,N_7583);
nor U8334 (N_8334,N_7535,N_7790);
nand U8335 (N_8335,N_7613,N_7636);
nor U8336 (N_8336,N_7851,N_7987);
nor U8337 (N_8337,N_7957,N_7853);
xnor U8338 (N_8338,N_7894,N_7587);
and U8339 (N_8339,N_7869,N_7972);
nand U8340 (N_8340,N_7768,N_7939);
or U8341 (N_8341,N_7922,N_7915);
or U8342 (N_8342,N_7707,N_7622);
xor U8343 (N_8343,N_7847,N_7780);
nand U8344 (N_8344,N_7968,N_7970);
nor U8345 (N_8345,N_7936,N_7887);
xnor U8346 (N_8346,N_7802,N_7544);
xor U8347 (N_8347,N_7853,N_7623);
or U8348 (N_8348,N_7726,N_7511);
nor U8349 (N_8349,N_7580,N_7691);
nand U8350 (N_8350,N_7799,N_7771);
or U8351 (N_8351,N_7971,N_7863);
nor U8352 (N_8352,N_7761,N_7967);
nor U8353 (N_8353,N_7608,N_7996);
nor U8354 (N_8354,N_7797,N_7553);
or U8355 (N_8355,N_7827,N_7829);
or U8356 (N_8356,N_7735,N_7905);
nor U8357 (N_8357,N_7562,N_7680);
and U8358 (N_8358,N_7940,N_7999);
xor U8359 (N_8359,N_7985,N_7684);
or U8360 (N_8360,N_7849,N_7566);
or U8361 (N_8361,N_7586,N_7816);
nor U8362 (N_8362,N_7605,N_7565);
and U8363 (N_8363,N_7956,N_7946);
nor U8364 (N_8364,N_7833,N_7618);
nand U8365 (N_8365,N_7707,N_7739);
nand U8366 (N_8366,N_7542,N_7893);
xor U8367 (N_8367,N_7921,N_7609);
or U8368 (N_8368,N_7669,N_7667);
and U8369 (N_8369,N_7928,N_7721);
or U8370 (N_8370,N_7837,N_7992);
or U8371 (N_8371,N_7592,N_7689);
nand U8372 (N_8372,N_7677,N_7680);
nand U8373 (N_8373,N_7919,N_7595);
xnor U8374 (N_8374,N_7637,N_7723);
and U8375 (N_8375,N_7856,N_7504);
xor U8376 (N_8376,N_7765,N_7598);
nand U8377 (N_8377,N_7540,N_7724);
or U8378 (N_8378,N_7514,N_7710);
nand U8379 (N_8379,N_7903,N_7968);
or U8380 (N_8380,N_7901,N_7889);
xnor U8381 (N_8381,N_7794,N_7763);
xnor U8382 (N_8382,N_7658,N_7982);
nor U8383 (N_8383,N_7620,N_7903);
nor U8384 (N_8384,N_7785,N_7690);
and U8385 (N_8385,N_7826,N_7979);
xnor U8386 (N_8386,N_7686,N_7981);
and U8387 (N_8387,N_7973,N_7559);
nor U8388 (N_8388,N_7876,N_7639);
nand U8389 (N_8389,N_7583,N_7676);
xor U8390 (N_8390,N_7996,N_7758);
or U8391 (N_8391,N_7956,N_7926);
nand U8392 (N_8392,N_7523,N_7846);
or U8393 (N_8393,N_7618,N_7545);
nor U8394 (N_8394,N_7629,N_7708);
nand U8395 (N_8395,N_7886,N_7969);
or U8396 (N_8396,N_7913,N_7578);
or U8397 (N_8397,N_7700,N_7920);
nand U8398 (N_8398,N_7874,N_7526);
or U8399 (N_8399,N_7815,N_7708);
nand U8400 (N_8400,N_7854,N_7850);
nand U8401 (N_8401,N_7546,N_7772);
and U8402 (N_8402,N_7845,N_7745);
nand U8403 (N_8403,N_7878,N_7946);
nand U8404 (N_8404,N_7911,N_7701);
nand U8405 (N_8405,N_7844,N_7869);
nand U8406 (N_8406,N_7710,N_7848);
xor U8407 (N_8407,N_7506,N_7756);
or U8408 (N_8408,N_7693,N_7727);
or U8409 (N_8409,N_7851,N_7955);
nand U8410 (N_8410,N_7754,N_7888);
nor U8411 (N_8411,N_7585,N_7874);
nand U8412 (N_8412,N_7635,N_7591);
nor U8413 (N_8413,N_7911,N_7606);
nor U8414 (N_8414,N_7931,N_7961);
nand U8415 (N_8415,N_7651,N_7632);
nand U8416 (N_8416,N_7554,N_7735);
or U8417 (N_8417,N_7949,N_7688);
xnor U8418 (N_8418,N_7514,N_7915);
xor U8419 (N_8419,N_7613,N_7803);
or U8420 (N_8420,N_7976,N_7818);
xor U8421 (N_8421,N_7742,N_7759);
and U8422 (N_8422,N_7912,N_7836);
xnor U8423 (N_8423,N_7959,N_7544);
nor U8424 (N_8424,N_7663,N_7735);
nand U8425 (N_8425,N_7848,N_7541);
nand U8426 (N_8426,N_7900,N_7886);
nand U8427 (N_8427,N_7727,N_7510);
and U8428 (N_8428,N_7697,N_7520);
nor U8429 (N_8429,N_7879,N_7665);
nor U8430 (N_8430,N_7999,N_7862);
nand U8431 (N_8431,N_7989,N_7844);
or U8432 (N_8432,N_7889,N_7514);
nand U8433 (N_8433,N_7683,N_7994);
nor U8434 (N_8434,N_7570,N_7835);
and U8435 (N_8435,N_7923,N_7901);
nor U8436 (N_8436,N_7984,N_7511);
xor U8437 (N_8437,N_7956,N_7759);
or U8438 (N_8438,N_7705,N_7852);
and U8439 (N_8439,N_7604,N_7714);
xor U8440 (N_8440,N_7863,N_7705);
nand U8441 (N_8441,N_7520,N_7503);
xnor U8442 (N_8442,N_7690,N_7712);
nand U8443 (N_8443,N_7695,N_7711);
nor U8444 (N_8444,N_7876,N_7510);
and U8445 (N_8445,N_7879,N_7913);
nand U8446 (N_8446,N_7562,N_7794);
and U8447 (N_8447,N_7716,N_7919);
or U8448 (N_8448,N_7933,N_7614);
nor U8449 (N_8449,N_7778,N_7643);
and U8450 (N_8450,N_7719,N_7875);
and U8451 (N_8451,N_7727,N_7908);
xor U8452 (N_8452,N_7994,N_7520);
nor U8453 (N_8453,N_7854,N_7915);
nand U8454 (N_8454,N_7771,N_7870);
nand U8455 (N_8455,N_7712,N_7816);
nand U8456 (N_8456,N_7943,N_7673);
or U8457 (N_8457,N_7806,N_7540);
xor U8458 (N_8458,N_7538,N_7577);
or U8459 (N_8459,N_7892,N_7809);
nand U8460 (N_8460,N_7963,N_7844);
nand U8461 (N_8461,N_7823,N_7944);
and U8462 (N_8462,N_7864,N_7663);
or U8463 (N_8463,N_7759,N_7911);
xor U8464 (N_8464,N_7550,N_7548);
and U8465 (N_8465,N_7617,N_7644);
nor U8466 (N_8466,N_7714,N_7958);
and U8467 (N_8467,N_7877,N_7926);
xnor U8468 (N_8468,N_7661,N_7897);
xnor U8469 (N_8469,N_7783,N_7676);
nor U8470 (N_8470,N_7789,N_7612);
nand U8471 (N_8471,N_7579,N_7898);
nor U8472 (N_8472,N_7881,N_7684);
or U8473 (N_8473,N_7879,N_7854);
and U8474 (N_8474,N_7720,N_7951);
nor U8475 (N_8475,N_7689,N_7712);
nor U8476 (N_8476,N_7884,N_7848);
and U8477 (N_8477,N_7565,N_7739);
nand U8478 (N_8478,N_7510,N_7582);
xor U8479 (N_8479,N_7548,N_7789);
nor U8480 (N_8480,N_7539,N_7752);
nand U8481 (N_8481,N_7989,N_7940);
nand U8482 (N_8482,N_7502,N_7611);
or U8483 (N_8483,N_7915,N_7931);
and U8484 (N_8484,N_7761,N_7841);
nand U8485 (N_8485,N_7810,N_7922);
or U8486 (N_8486,N_7549,N_7862);
nor U8487 (N_8487,N_7677,N_7895);
nand U8488 (N_8488,N_7935,N_7530);
xor U8489 (N_8489,N_7542,N_7848);
and U8490 (N_8490,N_7765,N_7604);
nand U8491 (N_8491,N_7831,N_7538);
nor U8492 (N_8492,N_7912,N_7626);
or U8493 (N_8493,N_7875,N_7665);
nand U8494 (N_8494,N_7927,N_7576);
xor U8495 (N_8495,N_7905,N_7733);
or U8496 (N_8496,N_7876,N_7614);
and U8497 (N_8497,N_7772,N_7840);
and U8498 (N_8498,N_7647,N_7701);
nand U8499 (N_8499,N_7864,N_7726);
xor U8500 (N_8500,N_8015,N_8356);
nor U8501 (N_8501,N_8277,N_8234);
xor U8502 (N_8502,N_8261,N_8117);
or U8503 (N_8503,N_8096,N_8390);
nand U8504 (N_8504,N_8355,N_8030);
xor U8505 (N_8505,N_8276,N_8058);
or U8506 (N_8506,N_8463,N_8149);
or U8507 (N_8507,N_8422,N_8293);
nand U8508 (N_8508,N_8286,N_8453);
nand U8509 (N_8509,N_8391,N_8244);
and U8510 (N_8510,N_8387,N_8256);
nand U8511 (N_8511,N_8367,N_8037);
xor U8512 (N_8512,N_8473,N_8112);
and U8513 (N_8513,N_8179,N_8181);
nand U8514 (N_8514,N_8359,N_8205);
or U8515 (N_8515,N_8141,N_8364);
or U8516 (N_8516,N_8492,N_8378);
or U8517 (N_8517,N_8070,N_8371);
or U8518 (N_8518,N_8447,N_8430);
nand U8519 (N_8519,N_8002,N_8101);
or U8520 (N_8520,N_8079,N_8300);
nor U8521 (N_8521,N_8084,N_8050);
nand U8522 (N_8522,N_8423,N_8115);
nand U8523 (N_8523,N_8382,N_8097);
or U8524 (N_8524,N_8196,N_8026);
or U8525 (N_8525,N_8369,N_8021);
or U8526 (N_8526,N_8241,N_8311);
and U8527 (N_8527,N_8278,N_8043);
nand U8528 (N_8528,N_8366,N_8162);
or U8529 (N_8529,N_8439,N_8333);
or U8530 (N_8530,N_8236,N_8006);
nand U8531 (N_8531,N_8136,N_8290);
nand U8532 (N_8532,N_8393,N_8239);
xnor U8533 (N_8533,N_8232,N_8274);
nor U8534 (N_8534,N_8312,N_8123);
xor U8535 (N_8535,N_8100,N_8034);
xnor U8536 (N_8536,N_8316,N_8103);
or U8537 (N_8537,N_8342,N_8251);
or U8538 (N_8538,N_8013,N_8442);
and U8539 (N_8539,N_8040,N_8271);
or U8540 (N_8540,N_8477,N_8011);
or U8541 (N_8541,N_8093,N_8479);
or U8542 (N_8542,N_8491,N_8405);
xnor U8543 (N_8543,N_8113,N_8332);
xor U8544 (N_8544,N_8116,N_8017);
or U8545 (N_8545,N_8353,N_8090);
or U8546 (N_8546,N_8475,N_8468);
nand U8547 (N_8547,N_8207,N_8417);
nor U8548 (N_8548,N_8171,N_8133);
xnor U8549 (N_8549,N_8395,N_8338);
xnor U8550 (N_8550,N_8357,N_8461);
nand U8551 (N_8551,N_8374,N_8047);
nand U8552 (N_8552,N_8018,N_8172);
xor U8553 (N_8553,N_8418,N_8296);
or U8554 (N_8554,N_8137,N_8464);
xnor U8555 (N_8555,N_8210,N_8309);
xor U8556 (N_8556,N_8295,N_8036);
or U8557 (N_8557,N_8019,N_8023);
xnor U8558 (N_8558,N_8028,N_8089);
and U8559 (N_8559,N_8465,N_8164);
xnor U8560 (N_8560,N_8283,N_8246);
and U8561 (N_8561,N_8159,N_8305);
nor U8562 (N_8562,N_8257,N_8206);
and U8563 (N_8563,N_8303,N_8494);
nor U8564 (N_8564,N_8456,N_8401);
nor U8565 (N_8565,N_8068,N_8376);
nand U8566 (N_8566,N_8291,N_8451);
nand U8567 (N_8567,N_8433,N_8269);
and U8568 (N_8568,N_8202,N_8027);
nor U8569 (N_8569,N_8302,N_8424);
or U8570 (N_8570,N_8022,N_8299);
and U8571 (N_8571,N_8310,N_8488);
xor U8572 (N_8572,N_8098,N_8126);
or U8573 (N_8573,N_8386,N_8052);
nand U8574 (N_8574,N_8368,N_8016);
nor U8575 (N_8575,N_8069,N_8443);
or U8576 (N_8576,N_8223,N_8199);
or U8577 (N_8577,N_8320,N_8258);
nor U8578 (N_8578,N_8224,N_8243);
or U8579 (N_8579,N_8020,N_8249);
nor U8580 (N_8580,N_8389,N_8358);
and U8581 (N_8581,N_8003,N_8194);
or U8582 (N_8582,N_8111,N_8265);
and U8583 (N_8583,N_8125,N_8445);
nand U8584 (N_8584,N_8412,N_8087);
nor U8585 (N_8585,N_8250,N_8345);
xor U8586 (N_8586,N_8263,N_8252);
nand U8587 (N_8587,N_8275,N_8260);
nand U8588 (N_8588,N_8381,N_8336);
xnor U8589 (N_8589,N_8402,N_8304);
nand U8590 (N_8590,N_8388,N_8215);
or U8591 (N_8591,N_8347,N_8362);
nor U8592 (N_8592,N_8048,N_8165);
nand U8593 (N_8593,N_8313,N_8054);
nor U8594 (N_8594,N_8499,N_8483);
and U8595 (N_8595,N_8247,N_8448);
or U8596 (N_8596,N_8348,N_8327);
or U8597 (N_8597,N_8352,N_8325);
and U8598 (N_8598,N_8081,N_8363);
nor U8599 (N_8599,N_8268,N_8490);
and U8600 (N_8600,N_8014,N_8486);
or U8601 (N_8601,N_8351,N_8346);
xnor U8602 (N_8602,N_8025,N_8072);
xor U8603 (N_8603,N_8163,N_8044);
and U8604 (N_8604,N_8114,N_8001);
xor U8605 (N_8605,N_8394,N_8091);
nand U8606 (N_8606,N_8365,N_8071);
and U8607 (N_8607,N_8287,N_8480);
or U8608 (N_8608,N_8398,N_8130);
nand U8609 (N_8609,N_8000,N_8339);
and U8610 (N_8610,N_8235,N_8143);
nand U8611 (N_8611,N_8200,N_8487);
or U8612 (N_8612,N_8231,N_8450);
and U8613 (N_8613,N_8142,N_8214);
or U8614 (N_8614,N_8331,N_8484);
or U8615 (N_8615,N_8148,N_8057);
nand U8616 (N_8616,N_8184,N_8078);
nor U8617 (N_8617,N_8183,N_8471);
nor U8618 (N_8618,N_8322,N_8272);
xor U8619 (N_8619,N_8004,N_8399);
and U8620 (N_8620,N_8055,N_8462);
nand U8621 (N_8621,N_8161,N_8110);
nor U8622 (N_8622,N_8493,N_8062);
xor U8623 (N_8623,N_8012,N_8420);
nand U8624 (N_8624,N_8074,N_8452);
xor U8625 (N_8625,N_8242,N_8255);
xnor U8626 (N_8626,N_8178,N_8308);
nand U8627 (N_8627,N_8222,N_8167);
nand U8628 (N_8628,N_8419,N_8086);
or U8629 (N_8629,N_8253,N_8458);
nor U8630 (N_8630,N_8160,N_8416);
nand U8631 (N_8631,N_8318,N_8248);
and U8632 (N_8632,N_8099,N_8129);
nor U8633 (N_8633,N_8193,N_8176);
or U8634 (N_8634,N_8280,N_8496);
or U8635 (N_8635,N_8228,N_8024);
or U8636 (N_8636,N_8383,N_8120);
and U8637 (N_8637,N_8005,N_8436);
or U8638 (N_8638,N_8220,N_8227);
or U8639 (N_8639,N_8121,N_8059);
nor U8640 (N_8640,N_8427,N_8122);
nand U8641 (N_8641,N_8226,N_8370);
or U8642 (N_8642,N_8188,N_8341);
nor U8643 (N_8643,N_8254,N_8454);
or U8644 (N_8644,N_8108,N_8481);
or U8645 (N_8645,N_8307,N_8482);
and U8646 (N_8646,N_8440,N_8426);
nand U8647 (N_8647,N_8413,N_8127);
nor U8648 (N_8648,N_8498,N_8198);
or U8649 (N_8649,N_8185,N_8191);
and U8650 (N_8650,N_8384,N_8407);
xnor U8651 (N_8651,N_8095,N_8186);
and U8652 (N_8652,N_8134,N_8170);
and U8653 (N_8653,N_8400,N_8315);
or U8654 (N_8654,N_8404,N_8201);
xor U8655 (N_8655,N_8282,N_8033);
xnor U8656 (N_8656,N_8211,N_8213);
xnor U8657 (N_8657,N_8195,N_8009);
xor U8658 (N_8658,N_8372,N_8306);
xor U8659 (N_8659,N_8415,N_8489);
nand U8660 (N_8660,N_8008,N_8466);
and U8661 (N_8661,N_8007,N_8139);
and U8662 (N_8662,N_8182,N_8107);
nor U8663 (N_8663,N_8067,N_8219);
and U8664 (N_8664,N_8153,N_8173);
xnor U8665 (N_8665,N_8301,N_8428);
nor U8666 (N_8666,N_8403,N_8075);
xor U8667 (N_8667,N_8289,N_8083);
and U8668 (N_8668,N_8324,N_8180);
nand U8669 (N_8669,N_8425,N_8495);
xor U8670 (N_8670,N_8344,N_8411);
and U8671 (N_8671,N_8349,N_8140);
nand U8672 (N_8672,N_8414,N_8203);
nor U8673 (N_8673,N_8077,N_8334);
nand U8674 (N_8674,N_8124,N_8192);
or U8675 (N_8675,N_8266,N_8061);
nand U8676 (N_8676,N_8225,N_8157);
or U8677 (N_8677,N_8259,N_8063);
or U8678 (N_8678,N_8467,N_8102);
nand U8679 (N_8679,N_8264,N_8262);
nor U8680 (N_8680,N_8175,N_8190);
or U8681 (N_8681,N_8189,N_8237);
nand U8682 (N_8682,N_8267,N_8229);
nor U8683 (N_8683,N_8314,N_8435);
xnor U8684 (N_8684,N_8429,N_8151);
or U8685 (N_8685,N_8065,N_8146);
and U8686 (N_8686,N_8329,N_8457);
nand U8687 (N_8687,N_8377,N_8088);
and U8688 (N_8688,N_8379,N_8460);
xnor U8689 (N_8689,N_8446,N_8292);
xnor U8690 (N_8690,N_8217,N_8340);
and U8691 (N_8691,N_8221,N_8177);
nor U8692 (N_8692,N_8455,N_8029);
or U8693 (N_8693,N_8397,N_8233);
or U8694 (N_8694,N_8469,N_8056);
xnor U8695 (N_8695,N_8106,N_8270);
nand U8696 (N_8696,N_8046,N_8441);
xor U8697 (N_8697,N_8330,N_8049);
and U8698 (N_8698,N_8238,N_8144);
nor U8699 (N_8699,N_8152,N_8444);
nor U8700 (N_8700,N_8150,N_8031);
nor U8701 (N_8701,N_8474,N_8373);
nand U8702 (N_8702,N_8038,N_8204);
nand U8703 (N_8703,N_8156,N_8392);
or U8704 (N_8704,N_8361,N_8218);
and U8705 (N_8705,N_8459,N_8209);
nor U8706 (N_8706,N_8166,N_8051);
xnor U8707 (N_8707,N_8297,N_8279);
nand U8708 (N_8708,N_8406,N_8119);
or U8709 (N_8709,N_8135,N_8409);
xnor U8710 (N_8710,N_8449,N_8076);
nor U8711 (N_8711,N_8288,N_8039);
xor U8712 (N_8712,N_8350,N_8138);
nand U8713 (N_8713,N_8131,N_8158);
xor U8714 (N_8714,N_8208,N_8434);
nand U8715 (N_8715,N_8317,N_8216);
and U8716 (N_8716,N_8410,N_8328);
or U8717 (N_8717,N_8094,N_8169);
nor U8718 (N_8718,N_8060,N_8155);
nor U8719 (N_8719,N_8294,N_8174);
xor U8720 (N_8720,N_8092,N_8323);
xnor U8721 (N_8721,N_8375,N_8082);
xor U8722 (N_8722,N_8335,N_8360);
or U8723 (N_8723,N_8497,N_8041);
nor U8724 (N_8724,N_8042,N_8281);
nor U8725 (N_8725,N_8478,N_8154);
xnor U8726 (N_8726,N_8032,N_8431);
or U8727 (N_8727,N_8128,N_8326);
xnor U8728 (N_8728,N_8168,N_8354);
nor U8729 (N_8729,N_8470,N_8298);
and U8730 (N_8730,N_8421,N_8145);
nand U8731 (N_8731,N_8476,N_8285);
nor U8732 (N_8732,N_8337,N_8045);
xnor U8733 (N_8733,N_8104,N_8385);
or U8734 (N_8734,N_8380,N_8066);
nor U8735 (N_8735,N_8118,N_8053);
or U8736 (N_8736,N_8432,N_8105);
or U8737 (N_8737,N_8109,N_8073);
xor U8738 (N_8738,N_8197,N_8132);
nor U8739 (N_8739,N_8472,N_8230);
nand U8740 (N_8740,N_8147,N_8212);
or U8741 (N_8741,N_8273,N_8187);
nand U8742 (N_8742,N_8319,N_8245);
or U8743 (N_8743,N_8080,N_8064);
and U8744 (N_8744,N_8437,N_8343);
nor U8745 (N_8745,N_8485,N_8240);
nand U8746 (N_8746,N_8408,N_8085);
and U8747 (N_8747,N_8035,N_8396);
and U8748 (N_8748,N_8438,N_8321);
or U8749 (N_8749,N_8284,N_8010);
nand U8750 (N_8750,N_8212,N_8206);
nor U8751 (N_8751,N_8499,N_8012);
nand U8752 (N_8752,N_8100,N_8136);
nor U8753 (N_8753,N_8211,N_8286);
xor U8754 (N_8754,N_8342,N_8227);
or U8755 (N_8755,N_8118,N_8256);
or U8756 (N_8756,N_8091,N_8081);
nor U8757 (N_8757,N_8035,N_8101);
nor U8758 (N_8758,N_8453,N_8207);
nand U8759 (N_8759,N_8239,N_8463);
or U8760 (N_8760,N_8098,N_8143);
or U8761 (N_8761,N_8126,N_8384);
or U8762 (N_8762,N_8077,N_8198);
and U8763 (N_8763,N_8451,N_8401);
nand U8764 (N_8764,N_8028,N_8469);
nand U8765 (N_8765,N_8373,N_8336);
and U8766 (N_8766,N_8157,N_8428);
nand U8767 (N_8767,N_8422,N_8380);
xnor U8768 (N_8768,N_8313,N_8291);
or U8769 (N_8769,N_8167,N_8138);
nand U8770 (N_8770,N_8231,N_8000);
or U8771 (N_8771,N_8027,N_8459);
or U8772 (N_8772,N_8154,N_8230);
xnor U8773 (N_8773,N_8291,N_8193);
xnor U8774 (N_8774,N_8336,N_8158);
nand U8775 (N_8775,N_8191,N_8427);
or U8776 (N_8776,N_8124,N_8140);
xnor U8777 (N_8777,N_8430,N_8392);
and U8778 (N_8778,N_8323,N_8355);
xor U8779 (N_8779,N_8224,N_8027);
nor U8780 (N_8780,N_8203,N_8216);
xnor U8781 (N_8781,N_8053,N_8241);
nor U8782 (N_8782,N_8243,N_8027);
xor U8783 (N_8783,N_8455,N_8354);
nand U8784 (N_8784,N_8453,N_8442);
xnor U8785 (N_8785,N_8065,N_8170);
nor U8786 (N_8786,N_8319,N_8220);
nand U8787 (N_8787,N_8382,N_8303);
or U8788 (N_8788,N_8360,N_8236);
or U8789 (N_8789,N_8260,N_8242);
and U8790 (N_8790,N_8297,N_8119);
and U8791 (N_8791,N_8109,N_8279);
xor U8792 (N_8792,N_8067,N_8073);
or U8793 (N_8793,N_8012,N_8307);
nand U8794 (N_8794,N_8439,N_8070);
or U8795 (N_8795,N_8235,N_8142);
and U8796 (N_8796,N_8025,N_8470);
xnor U8797 (N_8797,N_8386,N_8474);
nor U8798 (N_8798,N_8172,N_8337);
and U8799 (N_8799,N_8404,N_8443);
nor U8800 (N_8800,N_8414,N_8250);
nor U8801 (N_8801,N_8074,N_8415);
nand U8802 (N_8802,N_8434,N_8268);
and U8803 (N_8803,N_8071,N_8212);
nor U8804 (N_8804,N_8294,N_8175);
or U8805 (N_8805,N_8484,N_8173);
and U8806 (N_8806,N_8154,N_8473);
and U8807 (N_8807,N_8046,N_8058);
and U8808 (N_8808,N_8398,N_8430);
xnor U8809 (N_8809,N_8469,N_8024);
nor U8810 (N_8810,N_8085,N_8223);
nand U8811 (N_8811,N_8268,N_8088);
nor U8812 (N_8812,N_8414,N_8375);
nor U8813 (N_8813,N_8135,N_8119);
or U8814 (N_8814,N_8343,N_8006);
or U8815 (N_8815,N_8425,N_8175);
or U8816 (N_8816,N_8163,N_8361);
or U8817 (N_8817,N_8338,N_8305);
nand U8818 (N_8818,N_8249,N_8277);
nor U8819 (N_8819,N_8258,N_8197);
nand U8820 (N_8820,N_8269,N_8353);
xor U8821 (N_8821,N_8059,N_8024);
nand U8822 (N_8822,N_8495,N_8019);
nor U8823 (N_8823,N_8207,N_8142);
xor U8824 (N_8824,N_8332,N_8383);
xnor U8825 (N_8825,N_8129,N_8327);
or U8826 (N_8826,N_8476,N_8265);
or U8827 (N_8827,N_8370,N_8011);
and U8828 (N_8828,N_8198,N_8114);
nand U8829 (N_8829,N_8200,N_8410);
nor U8830 (N_8830,N_8167,N_8285);
and U8831 (N_8831,N_8339,N_8334);
or U8832 (N_8832,N_8194,N_8425);
or U8833 (N_8833,N_8028,N_8002);
nor U8834 (N_8834,N_8207,N_8483);
nand U8835 (N_8835,N_8413,N_8438);
xor U8836 (N_8836,N_8340,N_8324);
and U8837 (N_8837,N_8192,N_8087);
xnor U8838 (N_8838,N_8232,N_8483);
and U8839 (N_8839,N_8442,N_8110);
nand U8840 (N_8840,N_8427,N_8417);
nor U8841 (N_8841,N_8082,N_8147);
nor U8842 (N_8842,N_8011,N_8037);
and U8843 (N_8843,N_8049,N_8297);
xnor U8844 (N_8844,N_8489,N_8140);
nand U8845 (N_8845,N_8285,N_8429);
nor U8846 (N_8846,N_8070,N_8370);
and U8847 (N_8847,N_8374,N_8043);
nand U8848 (N_8848,N_8300,N_8260);
nand U8849 (N_8849,N_8154,N_8125);
nand U8850 (N_8850,N_8171,N_8402);
or U8851 (N_8851,N_8275,N_8216);
and U8852 (N_8852,N_8093,N_8426);
nand U8853 (N_8853,N_8144,N_8233);
nor U8854 (N_8854,N_8286,N_8138);
and U8855 (N_8855,N_8357,N_8001);
and U8856 (N_8856,N_8223,N_8046);
and U8857 (N_8857,N_8298,N_8402);
and U8858 (N_8858,N_8124,N_8240);
nand U8859 (N_8859,N_8421,N_8132);
xnor U8860 (N_8860,N_8313,N_8159);
nor U8861 (N_8861,N_8109,N_8016);
xor U8862 (N_8862,N_8102,N_8335);
nand U8863 (N_8863,N_8418,N_8330);
xor U8864 (N_8864,N_8148,N_8053);
xor U8865 (N_8865,N_8247,N_8202);
xor U8866 (N_8866,N_8214,N_8286);
nor U8867 (N_8867,N_8229,N_8118);
nand U8868 (N_8868,N_8376,N_8157);
and U8869 (N_8869,N_8336,N_8228);
nor U8870 (N_8870,N_8284,N_8495);
xnor U8871 (N_8871,N_8315,N_8496);
xnor U8872 (N_8872,N_8492,N_8145);
and U8873 (N_8873,N_8286,N_8091);
nand U8874 (N_8874,N_8092,N_8349);
nor U8875 (N_8875,N_8428,N_8437);
nand U8876 (N_8876,N_8439,N_8345);
xnor U8877 (N_8877,N_8452,N_8470);
nand U8878 (N_8878,N_8383,N_8026);
or U8879 (N_8879,N_8072,N_8391);
nor U8880 (N_8880,N_8444,N_8383);
nor U8881 (N_8881,N_8383,N_8485);
or U8882 (N_8882,N_8180,N_8125);
and U8883 (N_8883,N_8235,N_8463);
nor U8884 (N_8884,N_8095,N_8079);
nor U8885 (N_8885,N_8306,N_8096);
or U8886 (N_8886,N_8453,N_8305);
and U8887 (N_8887,N_8397,N_8051);
xor U8888 (N_8888,N_8235,N_8440);
nor U8889 (N_8889,N_8357,N_8149);
or U8890 (N_8890,N_8447,N_8483);
and U8891 (N_8891,N_8441,N_8471);
nand U8892 (N_8892,N_8236,N_8471);
and U8893 (N_8893,N_8040,N_8078);
or U8894 (N_8894,N_8491,N_8452);
nor U8895 (N_8895,N_8110,N_8176);
nor U8896 (N_8896,N_8294,N_8154);
xnor U8897 (N_8897,N_8479,N_8250);
or U8898 (N_8898,N_8297,N_8378);
nor U8899 (N_8899,N_8388,N_8477);
or U8900 (N_8900,N_8042,N_8308);
nand U8901 (N_8901,N_8458,N_8109);
or U8902 (N_8902,N_8225,N_8044);
nor U8903 (N_8903,N_8220,N_8428);
and U8904 (N_8904,N_8011,N_8184);
nor U8905 (N_8905,N_8042,N_8360);
nand U8906 (N_8906,N_8158,N_8481);
or U8907 (N_8907,N_8121,N_8310);
nand U8908 (N_8908,N_8456,N_8151);
nand U8909 (N_8909,N_8365,N_8229);
and U8910 (N_8910,N_8496,N_8035);
xor U8911 (N_8911,N_8041,N_8489);
or U8912 (N_8912,N_8243,N_8136);
nand U8913 (N_8913,N_8041,N_8190);
xnor U8914 (N_8914,N_8233,N_8213);
nand U8915 (N_8915,N_8056,N_8493);
nand U8916 (N_8916,N_8469,N_8198);
nor U8917 (N_8917,N_8010,N_8051);
nor U8918 (N_8918,N_8191,N_8321);
nand U8919 (N_8919,N_8133,N_8379);
and U8920 (N_8920,N_8066,N_8334);
nand U8921 (N_8921,N_8129,N_8370);
or U8922 (N_8922,N_8401,N_8316);
nor U8923 (N_8923,N_8472,N_8207);
xor U8924 (N_8924,N_8005,N_8492);
xor U8925 (N_8925,N_8490,N_8485);
nor U8926 (N_8926,N_8043,N_8459);
nand U8927 (N_8927,N_8080,N_8245);
or U8928 (N_8928,N_8219,N_8332);
and U8929 (N_8929,N_8007,N_8384);
nor U8930 (N_8930,N_8055,N_8301);
or U8931 (N_8931,N_8218,N_8395);
and U8932 (N_8932,N_8048,N_8443);
and U8933 (N_8933,N_8142,N_8051);
xnor U8934 (N_8934,N_8270,N_8105);
nor U8935 (N_8935,N_8386,N_8077);
xnor U8936 (N_8936,N_8157,N_8426);
or U8937 (N_8937,N_8415,N_8181);
nand U8938 (N_8938,N_8082,N_8193);
nor U8939 (N_8939,N_8170,N_8184);
or U8940 (N_8940,N_8084,N_8078);
nor U8941 (N_8941,N_8242,N_8283);
xnor U8942 (N_8942,N_8090,N_8275);
or U8943 (N_8943,N_8026,N_8015);
or U8944 (N_8944,N_8219,N_8329);
nor U8945 (N_8945,N_8253,N_8453);
xnor U8946 (N_8946,N_8390,N_8114);
or U8947 (N_8947,N_8459,N_8228);
or U8948 (N_8948,N_8477,N_8079);
and U8949 (N_8949,N_8441,N_8143);
nor U8950 (N_8950,N_8011,N_8399);
xor U8951 (N_8951,N_8405,N_8117);
nor U8952 (N_8952,N_8449,N_8447);
xor U8953 (N_8953,N_8341,N_8026);
nand U8954 (N_8954,N_8207,N_8136);
and U8955 (N_8955,N_8099,N_8421);
xor U8956 (N_8956,N_8228,N_8480);
or U8957 (N_8957,N_8024,N_8044);
and U8958 (N_8958,N_8018,N_8249);
and U8959 (N_8959,N_8394,N_8103);
and U8960 (N_8960,N_8026,N_8295);
or U8961 (N_8961,N_8326,N_8394);
or U8962 (N_8962,N_8025,N_8344);
nor U8963 (N_8963,N_8417,N_8160);
nand U8964 (N_8964,N_8162,N_8312);
xor U8965 (N_8965,N_8054,N_8342);
nand U8966 (N_8966,N_8118,N_8253);
nor U8967 (N_8967,N_8393,N_8255);
nand U8968 (N_8968,N_8004,N_8269);
xor U8969 (N_8969,N_8297,N_8490);
or U8970 (N_8970,N_8133,N_8184);
and U8971 (N_8971,N_8126,N_8016);
xor U8972 (N_8972,N_8335,N_8402);
nand U8973 (N_8973,N_8111,N_8026);
or U8974 (N_8974,N_8245,N_8047);
xor U8975 (N_8975,N_8147,N_8478);
or U8976 (N_8976,N_8300,N_8310);
xor U8977 (N_8977,N_8428,N_8307);
or U8978 (N_8978,N_8161,N_8216);
nor U8979 (N_8979,N_8189,N_8254);
or U8980 (N_8980,N_8293,N_8455);
xor U8981 (N_8981,N_8410,N_8119);
and U8982 (N_8982,N_8141,N_8393);
nand U8983 (N_8983,N_8116,N_8246);
xor U8984 (N_8984,N_8476,N_8450);
and U8985 (N_8985,N_8211,N_8326);
nand U8986 (N_8986,N_8184,N_8294);
or U8987 (N_8987,N_8317,N_8406);
and U8988 (N_8988,N_8312,N_8387);
nand U8989 (N_8989,N_8437,N_8223);
nand U8990 (N_8990,N_8327,N_8491);
and U8991 (N_8991,N_8454,N_8460);
nor U8992 (N_8992,N_8323,N_8473);
nand U8993 (N_8993,N_8159,N_8194);
nand U8994 (N_8994,N_8352,N_8365);
or U8995 (N_8995,N_8249,N_8408);
xnor U8996 (N_8996,N_8397,N_8132);
and U8997 (N_8997,N_8418,N_8139);
xnor U8998 (N_8998,N_8278,N_8123);
nand U8999 (N_8999,N_8071,N_8045);
nand U9000 (N_9000,N_8815,N_8744);
and U9001 (N_9001,N_8674,N_8836);
nor U9002 (N_9002,N_8641,N_8905);
and U9003 (N_9003,N_8998,N_8933);
or U9004 (N_9004,N_8520,N_8653);
and U9005 (N_9005,N_8665,N_8545);
nor U9006 (N_9006,N_8870,N_8848);
nand U9007 (N_9007,N_8553,N_8658);
nand U9008 (N_9008,N_8805,N_8590);
nor U9009 (N_9009,N_8881,N_8779);
xor U9010 (N_9010,N_8627,N_8776);
or U9011 (N_9011,N_8622,N_8742);
and U9012 (N_9012,N_8885,N_8555);
xnor U9013 (N_9013,N_8646,N_8681);
or U9014 (N_9014,N_8542,N_8584);
xnor U9015 (N_9015,N_8867,N_8823);
and U9016 (N_9016,N_8526,N_8951);
and U9017 (N_9017,N_8800,N_8821);
nor U9018 (N_9018,N_8513,N_8615);
or U9019 (N_9019,N_8792,N_8928);
and U9020 (N_9020,N_8771,N_8747);
and U9021 (N_9021,N_8927,N_8803);
nor U9022 (N_9022,N_8826,N_8856);
and U9023 (N_9023,N_8983,N_8900);
nand U9024 (N_9024,N_8739,N_8713);
and U9025 (N_9025,N_8997,N_8620);
nand U9026 (N_9026,N_8539,N_8849);
nand U9027 (N_9027,N_8810,N_8637);
nand U9028 (N_9028,N_8970,N_8669);
xor U9029 (N_9029,N_8813,N_8563);
nor U9030 (N_9030,N_8929,N_8524);
xor U9031 (N_9031,N_8847,N_8985);
xnor U9032 (N_9032,N_8668,N_8572);
and U9033 (N_9033,N_8599,N_8683);
xor U9034 (N_9034,N_8897,N_8649);
and U9035 (N_9035,N_8611,N_8760);
nand U9036 (N_9036,N_8922,N_8509);
xor U9037 (N_9037,N_8945,N_8861);
and U9038 (N_9038,N_8872,N_8921);
nand U9039 (N_9039,N_8934,N_8659);
nor U9040 (N_9040,N_8876,N_8636);
xor U9041 (N_9041,N_8950,N_8574);
or U9042 (N_9042,N_8576,N_8698);
nor U9043 (N_9043,N_8548,N_8505);
nand U9044 (N_9044,N_8736,N_8535);
or U9045 (N_9045,N_8979,N_8875);
xor U9046 (N_9046,N_8651,N_8871);
and U9047 (N_9047,N_8931,N_8525);
and U9048 (N_9048,N_8634,N_8925);
and U9049 (N_9049,N_8581,N_8775);
and U9050 (N_9050,N_8570,N_8814);
and U9051 (N_9051,N_8840,N_8903);
and U9052 (N_9052,N_8600,N_8781);
xor U9053 (N_9053,N_8948,N_8991);
nand U9054 (N_9054,N_8886,N_8918);
or U9055 (N_9055,N_8729,N_8660);
or U9056 (N_9056,N_8715,N_8710);
and U9057 (N_9057,N_8566,N_8911);
nand U9058 (N_9058,N_8994,N_8967);
and U9059 (N_9059,N_8961,N_8853);
and U9060 (N_9060,N_8989,N_8841);
nor U9061 (N_9061,N_8583,N_8746);
nand U9062 (N_9062,N_8694,N_8935);
nor U9063 (N_9063,N_8774,N_8626);
nor U9064 (N_9064,N_8788,N_8569);
xor U9065 (N_9065,N_8733,N_8724);
xor U9066 (N_9066,N_8944,N_8974);
nand U9067 (N_9067,N_8832,N_8968);
nand U9068 (N_9068,N_8690,N_8888);
nor U9069 (N_9069,N_8824,N_8633);
xnor U9070 (N_9070,N_8995,N_8768);
xor U9071 (N_9071,N_8816,N_8504);
nand U9072 (N_9072,N_8552,N_8707);
xor U9073 (N_9073,N_8812,N_8829);
nand U9074 (N_9074,N_8625,N_8947);
or U9075 (N_9075,N_8766,N_8703);
or U9076 (N_9076,N_8869,N_8663);
xor U9077 (N_9077,N_8891,N_8882);
nor U9078 (N_9078,N_8577,N_8786);
and U9079 (N_9079,N_8868,N_8657);
nor U9080 (N_9080,N_8941,N_8664);
nor U9081 (N_9081,N_8873,N_8680);
xor U9082 (N_9082,N_8516,N_8671);
and U9083 (N_9083,N_8817,N_8688);
nor U9084 (N_9084,N_8589,N_8579);
nand U9085 (N_9085,N_8758,N_8936);
or U9086 (N_9086,N_8644,N_8978);
or U9087 (N_9087,N_8559,N_8784);
and U9088 (N_9088,N_8924,N_8613);
nand U9089 (N_9089,N_8981,N_8679);
xnor U9090 (N_9090,N_8798,N_8656);
and U9091 (N_9091,N_8631,N_8783);
and U9092 (N_9092,N_8670,N_8635);
and U9093 (N_9093,N_8842,N_8986);
nor U9094 (N_9094,N_8558,N_8820);
nor U9095 (N_9095,N_8639,N_8791);
xnor U9096 (N_9096,N_8585,N_8692);
and U9097 (N_9097,N_8597,N_8643);
and U9098 (N_9098,N_8699,N_8790);
and U9099 (N_9099,N_8762,N_8735);
or U9100 (N_9100,N_8866,N_8773);
xor U9101 (N_9101,N_8892,N_8789);
nand U9102 (N_9102,N_8508,N_8580);
xnor U9103 (N_9103,N_8538,N_8568);
and U9104 (N_9104,N_8958,N_8706);
xor U9105 (N_9105,N_8887,N_8598);
and U9106 (N_9106,N_8737,N_8624);
or U9107 (N_9107,N_8603,N_8547);
xnor U9108 (N_9108,N_8962,N_8727);
and U9109 (N_9109,N_8592,N_8720);
nand U9110 (N_9110,N_8953,N_8952);
nand U9111 (N_9111,N_8554,N_8537);
nand U9112 (N_9112,N_8731,N_8647);
nand U9113 (N_9113,N_8667,N_8761);
or U9114 (N_9114,N_8898,N_8763);
nand U9115 (N_9115,N_8769,N_8977);
or U9116 (N_9116,N_8987,N_8595);
xor U9117 (N_9117,N_8531,N_8591);
or U9118 (N_9118,N_8618,N_8894);
and U9119 (N_9119,N_8793,N_8772);
or U9120 (N_9120,N_8807,N_8878);
or U9121 (N_9121,N_8770,N_8621);
or U9122 (N_9122,N_8920,N_8966);
xor U9123 (N_9123,N_8850,N_8880);
nor U9124 (N_9124,N_8993,N_8719);
nand U9125 (N_9125,N_8732,N_8556);
nand U9126 (N_9126,N_8912,N_8972);
nor U9127 (N_9127,N_8907,N_8695);
nor U9128 (N_9128,N_8976,N_8623);
and U9129 (N_9129,N_8743,N_8540);
nand U9130 (N_9130,N_8839,N_8677);
nor U9131 (N_9131,N_8612,N_8844);
xnor U9132 (N_9132,N_8596,N_8687);
and U9133 (N_9133,N_8652,N_8514);
xor U9134 (N_9134,N_8711,N_8702);
nand U9135 (N_9135,N_8716,N_8831);
nand U9136 (N_9136,N_8586,N_8883);
nor U9137 (N_9137,N_8956,N_8607);
nor U9138 (N_9138,N_8648,N_8796);
or U9139 (N_9139,N_8517,N_8666);
xnor U9140 (N_9140,N_8534,N_8500);
nand U9141 (N_9141,N_8879,N_8999);
or U9142 (N_9142,N_8510,N_8661);
and U9143 (N_9143,N_8971,N_8594);
xnor U9144 (N_9144,N_8960,N_8593);
xnor U9145 (N_9145,N_8862,N_8910);
and U9146 (N_9146,N_8723,N_8859);
or U9147 (N_9147,N_8946,N_8700);
or U9148 (N_9148,N_8527,N_8588);
nand U9149 (N_9149,N_8632,N_8765);
xor U9150 (N_9150,N_8754,N_8899);
nand U9151 (N_9151,N_8794,N_8806);
nand U9152 (N_9152,N_8819,N_8511);
and U9153 (N_9153,N_8601,N_8686);
xnor U9154 (N_9154,N_8908,N_8565);
nor U9155 (N_9155,N_8830,N_8799);
or U9156 (N_9156,N_8914,N_8619);
or U9157 (N_9157,N_8777,N_8884);
nor U9158 (N_9158,N_8551,N_8521);
xnor U9159 (N_9159,N_8696,N_8506);
or U9160 (N_9160,N_8895,N_8852);
and U9161 (N_9161,N_8738,N_8795);
xor U9162 (N_9162,N_8544,N_8782);
xnor U9163 (N_9163,N_8536,N_8837);
nand U9164 (N_9164,N_8955,N_8709);
nand U9165 (N_9165,N_8726,N_8797);
nand U9166 (N_9166,N_8606,N_8825);
xnor U9167 (N_9167,N_8750,N_8909);
nor U9168 (N_9168,N_8751,N_8529);
xnor U9169 (N_9169,N_8969,N_8678);
and U9170 (N_9170,N_8838,N_8860);
or U9171 (N_9171,N_8843,N_8512);
nand U9172 (N_9172,N_8864,N_8756);
nor U9173 (N_9173,N_8917,N_8578);
or U9174 (N_9174,N_8515,N_8858);
or U9175 (N_9175,N_8693,N_8827);
and U9176 (N_9176,N_8673,N_8642);
xor U9177 (N_9177,N_8902,N_8582);
xor U9178 (N_9178,N_8501,N_8571);
and U9179 (N_9179,N_8801,N_8630);
nand U9180 (N_9180,N_8503,N_8802);
xor U9181 (N_9181,N_8865,N_8889);
nand U9182 (N_9182,N_8655,N_8752);
xnor U9183 (N_9183,N_8780,N_8759);
nand U9184 (N_9184,N_8753,N_8982);
and U9185 (N_9185,N_8609,N_8988);
or U9186 (N_9186,N_8682,N_8638);
nor U9187 (N_9187,N_8672,N_8822);
or U9188 (N_9188,N_8573,N_8764);
nor U9189 (N_9189,N_8640,N_8877);
xnor U9190 (N_9190,N_8519,N_8629);
xnor U9191 (N_9191,N_8662,N_8518);
xor U9192 (N_9192,N_8930,N_8602);
nand U9193 (N_9193,N_8973,N_8533);
xor U9194 (N_9194,N_8835,N_8734);
nor U9195 (N_9195,N_8992,N_8705);
or U9196 (N_9196,N_8916,N_8704);
and U9197 (N_9197,N_8650,N_8575);
and U9198 (N_9198,N_8728,N_8560);
nand U9199 (N_9199,N_8616,N_8749);
nand U9200 (N_9200,N_8778,N_8507);
or U9201 (N_9201,N_8804,N_8740);
xnor U9202 (N_9202,N_8522,N_8854);
and U9203 (N_9203,N_8628,N_8846);
and U9204 (N_9204,N_8562,N_8863);
or U9205 (N_9205,N_8939,N_8890);
nand U9206 (N_9206,N_8697,N_8959);
nor U9207 (N_9207,N_8787,N_8901);
or U9208 (N_9208,N_8975,N_8675);
and U9209 (N_9209,N_8818,N_8604);
nand U9210 (N_9210,N_8845,N_8617);
and U9211 (N_9211,N_8550,N_8923);
nor U9212 (N_9212,N_8708,N_8567);
xor U9213 (N_9213,N_8718,N_8717);
xor U9214 (N_9214,N_8587,N_8714);
nor U9215 (N_9215,N_8964,N_8684);
xor U9216 (N_9216,N_8828,N_8757);
nor U9217 (N_9217,N_8712,N_8857);
nor U9218 (N_9218,N_8532,N_8808);
nor U9219 (N_9219,N_8748,N_8676);
nor U9220 (N_9220,N_8701,N_8906);
and U9221 (N_9221,N_8874,N_8541);
xnor U9222 (N_9222,N_8564,N_8926);
and U9223 (N_9223,N_8689,N_8990);
nand U9224 (N_9224,N_8502,N_8963);
xnor U9225 (N_9225,N_8546,N_8893);
xor U9226 (N_9226,N_8608,N_8855);
xnor U9227 (N_9227,N_8645,N_8943);
or U9228 (N_9228,N_8722,N_8557);
nor U9229 (N_9229,N_8932,N_8543);
nand U9230 (N_9230,N_8745,N_8913);
nand U9231 (N_9231,N_8957,N_8730);
and U9232 (N_9232,N_8523,N_8833);
or U9233 (N_9233,N_8965,N_8549);
nor U9234 (N_9234,N_8785,N_8851);
or U9235 (N_9235,N_8755,N_8530);
and U9236 (N_9236,N_8721,N_8937);
nand U9237 (N_9237,N_8811,N_8741);
xnor U9238 (N_9238,N_8919,N_8996);
nand U9239 (N_9239,N_8984,N_8980);
xnor U9240 (N_9240,N_8915,N_8949);
or U9241 (N_9241,N_8685,N_8940);
or U9242 (N_9242,N_8528,N_8896);
xnor U9243 (N_9243,N_8904,N_8691);
and U9244 (N_9244,N_8834,N_8767);
nor U9245 (N_9245,N_8938,N_8954);
or U9246 (N_9246,N_8614,N_8654);
xor U9247 (N_9247,N_8725,N_8942);
nor U9248 (N_9248,N_8605,N_8561);
nor U9249 (N_9249,N_8809,N_8610);
and U9250 (N_9250,N_8865,N_8504);
or U9251 (N_9251,N_8698,N_8536);
and U9252 (N_9252,N_8813,N_8671);
and U9253 (N_9253,N_8790,N_8913);
or U9254 (N_9254,N_8559,N_8895);
and U9255 (N_9255,N_8668,N_8694);
nand U9256 (N_9256,N_8725,N_8878);
nand U9257 (N_9257,N_8979,N_8556);
nand U9258 (N_9258,N_8646,N_8629);
or U9259 (N_9259,N_8997,N_8696);
nor U9260 (N_9260,N_8632,N_8996);
or U9261 (N_9261,N_8765,N_8926);
and U9262 (N_9262,N_8916,N_8881);
or U9263 (N_9263,N_8890,N_8731);
and U9264 (N_9264,N_8920,N_8944);
xor U9265 (N_9265,N_8739,N_8762);
or U9266 (N_9266,N_8938,N_8800);
nor U9267 (N_9267,N_8638,N_8952);
and U9268 (N_9268,N_8857,N_8942);
or U9269 (N_9269,N_8749,N_8754);
or U9270 (N_9270,N_8576,N_8757);
nand U9271 (N_9271,N_8581,N_8589);
and U9272 (N_9272,N_8759,N_8778);
and U9273 (N_9273,N_8625,N_8796);
nand U9274 (N_9274,N_8729,N_8622);
nor U9275 (N_9275,N_8938,N_8631);
nor U9276 (N_9276,N_8505,N_8815);
and U9277 (N_9277,N_8865,N_8886);
nand U9278 (N_9278,N_8550,N_8692);
nor U9279 (N_9279,N_8760,N_8736);
nor U9280 (N_9280,N_8882,N_8655);
xnor U9281 (N_9281,N_8806,N_8739);
and U9282 (N_9282,N_8743,N_8901);
nor U9283 (N_9283,N_8838,N_8670);
and U9284 (N_9284,N_8891,N_8602);
xnor U9285 (N_9285,N_8932,N_8536);
nor U9286 (N_9286,N_8907,N_8960);
xor U9287 (N_9287,N_8540,N_8822);
nand U9288 (N_9288,N_8587,N_8823);
or U9289 (N_9289,N_8904,N_8750);
nand U9290 (N_9290,N_8737,N_8931);
or U9291 (N_9291,N_8695,N_8827);
or U9292 (N_9292,N_8730,N_8639);
nand U9293 (N_9293,N_8894,N_8530);
or U9294 (N_9294,N_8797,N_8608);
xnor U9295 (N_9295,N_8942,N_8513);
xnor U9296 (N_9296,N_8941,N_8655);
xnor U9297 (N_9297,N_8861,N_8508);
or U9298 (N_9298,N_8781,N_8940);
xnor U9299 (N_9299,N_8548,N_8954);
nor U9300 (N_9300,N_8923,N_8647);
nor U9301 (N_9301,N_8915,N_8726);
nor U9302 (N_9302,N_8939,N_8610);
xnor U9303 (N_9303,N_8611,N_8968);
nand U9304 (N_9304,N_8594,N_8643);
nand U9305 (N_9305,N_8671,N_8993);
nand U9306 (N_9306,N_8932,N_8669);
or U9307 (N_9307,N_8629,N_8883);
nand U9308 (N_9308,N_8925,N_8943);
nor U9309 (N_9309,N_8606,N_8918);
nor U9310 (N_9310,N_8614,N_8727);
nand U9311 (N_9311,N_8737,N_8848);
nor U9312 (N_9312,N_8752,N_8914);
xor U9313 (N_9313,N_8815,N_8724);
xor U9314 (N_9314,N_8996,N_8585);
nand U9315 (N_9315,N_8588,N_8987);
nor U9316 (N_9316,N_8965,N_8571);
nand U9317 (N_9317,N_8997,N_8985);
nand U9318 (N_9318,N_8820,N_8915);
or U9319 (N_9319,N_8866,N_8774);
and U9320 (N_9320,N_8574,N_8912);
or U9321 (N_9321,N_8999,N_8803);
xnor U9322 (N_9322,N_8690,N_8741);
xnor U9323 (N_9323,N_8585,N_8988);
nor U9324 (N_9324,N_8835,N_8948);
nor U9325 (N_9325,N_8618,N_8594);
and U9326 (N_9326,N_8777,N_8981);
xnor U9327 (N_9327,N_8801,N_8907);
nor U9328 (N_9328,N_8739,N_8683);
or U9329 (N_9329,N_8835,N_8796);
nand U9330 (N_9330,N_8762,N_8585);
and U9331 (N_9331,N_8808,N_8669);
or U9332 (N_9332,N_8727,N_8636);
nand U9333 (N_9333,N_8527,N_8517);
nor U9334 (N_9334,N_8927,N_8896);
nor U9335 (N_9335,N_8823,N_8778);
nor U9336 (N_9336,N_8763,N_8902);
nand U9337 (N_9337,N_8738,N_8881);
or U9338 (N_9338,N_8918,N_8632);
xnor U9339 (N_9339,N_8663,N_8851);
nor U9340 (N_9340,N_8874,N_8964);
xnor U9341 (N_9341,N_8726,N_8840);
and U9342 (N_9342,N_8803,N_8721);
or U9343 (N_9343,N_8977,N_8875);
and U9344 (N_9344,N_8691,N_8932);
xnor U9345 (N_9345,N_8829,N_8900);
xnor U9346 (N_9346,N_8652,N_8856);
or U9347 (N_9347,N_8749,N_8692);
nor U9348 (N_9348,N_8777,N_8775);
or U9349 (N_9349,N_8742,N_8891);
xnor U9350 (N_9350,N_8567,N_8563);
and U9351 (N_9351,N_8595,N_8752);
and U9352 (N_9352,N_8748,N_8953);
and U9353 (N_9353,N_8719,N_8899);
xnor U9354 (N_9354,N_8983,N_8721);
and U9355 (N_9355,N_8543,N_8974);
xor U9356 (N_9356,N_8719,N_8724);
and U9357 (N_9357,N_8551,N_8810);
and U9358 (N_9358,N_8841,N_8518);
nor U9359 (N_9359,N_8738,N_8639);
nand U9360 (N_9360,N_8605,N_8513);
xnor U9361 (N_9361,N_8569,N_8675);
xnor U9362 (N_9362,N_8875,N_8553);
and U9363 (N_9363,N_8604,N_8912);
xnor U9364 (N_9364,N_8920,N_8546);
nand U9365 (N_9365,N_8747,N_8942);
nand U9366 (N_9366,N_8788,N_8594);
or U9367 (N_9367,N_8729,N_8929);
xnor U9368 (N_9368,N_8920,N_8589);
nand U9369 (N_9369,N_8860,N_8982);
and U9370 (N_9370,N_8554,N_8684);
or U9371 (N_9371,N_8829,N_8820);
xnor U9372 (N_9372,N_8607,N_8663);
nand U9373 (N_9373,N_8857,N_8759);
nand U9374 (N_9374,N_8982,N_8989);
xor U9375 (N_9375,N_8804,N_8681);
xnor U9376 (N_9376,N_8666,N_8923);
and U9377 (N_9377,N_8812,N_8854);
and U9378 (N_9378,N_8988,N_8925);
nor U9379 (N_9379,N_8626,N_8693);
nor U9380 (N_9380,N_8881,N_8692);
xor U9381 (N_9381,N_8697,N_8585);
and U9382 (N_9382,N_8755,N_8585);
or U9383 (N_9383,N_8826,N_8726);
xnor U9384 (N_9384,N_8877,N_8965);
nand U9385 (N_9385,N_8873,N_8752);
xor U9386 (N_9386,N_8791,N_8691);
and U9387 (N_9387,N_8703,N_8742);
or U9388 (N_9388,N_8558,N_8715);
nand U9389 (N_9389,N_8930,N_8677);
nor U9390 (N_9390,N_8843,N_8918);
xor U9391 (N_9391,N_8951,N_8889);
and U9392 (N_9392,N_8622,N_8792);
xnor U9393 (N_9393,N_8667,N_8521);
nor U9394 (N_9394,N_8881,N_8689);
nand U9395 (N_9395,N_8868,N_8917);
xor U9396 (N_9396,N_8629,N_8837);
nor U9397 (N_9397,N_8682,N_8838);
and U9398 (N_9398,N_8785,N_8791);
nor U9399 (N_9399,N_8989,N_8729);
nand U9400 (N_9400,N_8719,N_8706);
or U9401 (N_9401,N_8952,N_8988);
nand U9402 (N_9402,N_8713,N_8899);
nand U9403 (N_9403,N_8756,N_8637);
and U9404 (N_9404,N_8734,N_8550);
or U9405 (N_9405,N_8848,N_8581);
nand U9406 (N_9406,N_8968,N_8980);
nand U9407 (N_9407,N_8933,N_8925);
or U9408 (N_9408,N_8910,N_8554);
nand U9409 (N_9409,N_8818,N_8552);
nor U9410 (N_9410,N_8586,N_8724);
nor U9411 (N_9411,N_8954,N_8673);
and U9412 (N_9412,N_8730,N_8831);
nor U9413 (N_9413,N_8950,N_8676);
or U9414 (N_9414,N_8653,N_8676);
and U9415 (N_9415,N_8806,N_8816);
or U9416 (N_9416,N_8803,N_8598);
or U9417 (N_9417,N_8733,N_8699);
and U9418 (N_9418,N_8808,N_8751);
or U9419 (N_9419,N_8515,N_8695);
or U9420 (N_9420,N_8593,N_8917);
or U9421 (N_9421,N_8764,N_8593);
nor U9422 (N_9422,N_8956,N_8513);
or U9423 (N_9423,N_8719,N_8866);
xnor U9424 (N_9424,N_8994,N_8761);
xnor U9425 (N_9425,N_8910,N_8898);
nor U9426 (N_9426,N_8592,N_8502);
or U9427 (N_9427,N_8911,N_8637);
or U9428 (N_9428,N_8727,N_8992);
nand U9429 (N_9429,N_8757,N_8859);
nand U9430 (N_9430,N_8875,N_8958);
nand U9431 (N_9431,N_8572,N_8698);
nand U9432 (N_9432,N_8506,N_8887);
and U9433 (N_9433,N_8691,N_8770);
nor U9434 (N_9434,N_8541,N_8905);
and U9435 (N_9435,N_8527,N_8821);
and U9436 (N_9436,N_8770,N_8633);
nand U9437 (N_9437,N_8566,N_8822);
or U9438 (N_9438,N_8522,N_8608);
xor U9439 (N_9439,N_8753,N_8510);
nand U9440 (N_9440,N_8976,N_8739);
and U9441 (N_9441,N_8977,N_8964);
nor U9442 (N_9442,N_8633,N_8524);
nand U9443 (N_9443,N_8575,N_8845);
nor U9444 (N_9444,N_8772,N_8586);
or U9445 (N_9445,N_8701,N_8889);
xor U9446 (N_9446,N_8656,N_8873);
or U9447 (N_9447,N_8991,N_8885);
nor U9448 (N_9448,N_8966,N_8640);
nor U9449 (N_9449,N_8774,N_8829);
nand U9450 (N_9450,N_8574,N_8725);
nand U9451 (N_9451,N_8798,N_8752);
nand U9452 (N_9452,N_8543,N_8652);
nand U9453 (N_9453,N_8664,N_8624);
or U9454 (N_9454,N_8690,N_8769);
xnor U9455 (N_9455,N_8623,N_8534);
nand U9456 (N_9456,N_8743,N_8742);
xnor U9457 (N_9457,N_8954,N_8952);
xnor U9458 (N_9458,N_8812,N_8897);
and U9459 (N_9459,N_8831,N_8579);
nor U9460 (N_9460,N_8971,N_8576);
nor U9461 (N_9461,N_8619,N_8930);
xor U9462 (N_9462,N_8940,N_8996);
or U9463 (N_9463,N_8981,N_8568);
xnor U9464 (N_9464,N_8650,N_8845);
nor U9465 (N_9465,N_8718,N_8845);
nand U9466 (N_9466,N_8959,N_8857);
or U9467 (N_9467,N_8859,N_8634);
and U9468 (N_9468,N_8866,N_8971);
xor U9469 (N_9469,N_8879,N_8762);
and U9470 (N_9470,N_8774,N_8523);
and U9471 (N_9471,N_8966,N_8836);
nor U9472 (N_9472,N_8519,N_8951);
and U9473 (N_9473,N_8507,N_8858);
or U9474 (N_9474,N_8634,N_8799);
and U9475 (N_9475,N_8668,N_8777);
nor U9476 (N_9476,N_8794,N_8892);
xor U9477 (N_9477,N_8867,N_8658);
or U9478 (N_9478,N_8817,N_8720);
or U9479 (N_9479,N_8711,N_8570);
xor U9480 (N_9480,N_8859,N_8914);
xnor U9481 (N_9481,N_8702,N_8843);
and U9482 (N_9482,N_8903,N_8930);
xnor U9483 (N_9483,N_8659,N_8549);
nor U9484 (N_9484,N_8662,N_8837);
nor U9485 (N_9485,N_8747,N_8643);
nor U9486 (N_9486,N_8537,N_8752);
nand U9487 (N_9487,N_8965,N_8794);
nand U9488 (N_9488,N_8634,N_8926);
xnor U9489 (N_9489,N_8787,N_8960);
and U9490 (N_9490,N_8684,N_8517);
or U9491 (N_9491,N_8909,N_8572);
nor U9492 (N_9492,N_8625,N_8633);
and U9493 (N_9493,N_8858,N_8660);
or U9494 (N_9494,N_8965,N_8633);
xor U9495 (N_9495,N_8716,N_8945);
nand U9496 (N_9496,N_8743,N_8534);
nor U9497 (N_9497,N_8716,N_8563);
nand U9498 (N_9498,N_8643,N_8793);
nor U9499 (N_9499,N_8660,N_8608);
and U9500 (N_9500,N_9219,N_9495);
xnor U9501 (N_9501,N_9178,N_9408);
nor U9502 (N_9502,N_9275,N_9488);
and U9503 (N_9503,N_9431,N_9459);
nand U9504 (N_9504,N_9252,N_9198);
nor U9505 (N_9505,N_9155,N_9071);
nand U9506 (N_9506,N_9236,N_9205);
xnor U9507 (N_9507,N_9381,N_9383);
and U9508 (N_9508,N_9203,N_9407);
or U9509 (N_9509,N_9005,N_9070);
nor U9510 (N_9510,N_9182,N_9377);
and U9511 (N_9511,N_9111,N_9413);
nand U9512 (N_9512,N_9346,N_9397);
and U9513 (N_9513,N_9253,N_9196);
nor U9514 (N_9514,N_9031,N_9278);
xor U9515 (N_9515,N_9138,N_9026);
xor U9516 (N_9516,N_9463,N_9127);
or U9517 (N_9517,N_9404,N_9243);
nand U9518 (N_9518,N_9467,N_9051);
nand U9519 (N_9519,N_9064,N_9422);
nor U9520 (N_9520,N_9200,N_9106);
or U9521 (N_9521,N_9021,N_9487);
nor U9522 (N_9522,N_9328,N_9464);
xor U9523 (N_9523,N_9359,N_9398);
nor U9524 (N_9524,N_9014,N_9365);
and U9525 (N_9525,N_9101,N_9184);
or U9526 (N_9526,N_9323,N_9391);
xor U9527 (N_9527,N_9033,N_9396);
nor U9528 (N_9528,N_9117,N_9376);
and U9529 (N_9529,N_9284,N_9137);
or U9530 (N_9530,N_9439,N_9457);
or U9531 (N_9531,N_9177,N_9499);
xnor U9532 (N_9532,N_9250,N_9139);
or U9533 (N_9533,N_9379,N_9313);
and U9534 (N_9534,N_9481,N_9388);
nor U9535 (N_9535,N_9267,N_9287);
xnor U9536 (N_9536,N_9126,N_9295);
nor U9537 (N_9537,N_9226,N_9047);
nor U9538 (N_9538,N_9272,N_9086);
nor U9539 (N_9539,N_9339,N_9333);
or U9540 (N_9540,N_9228,N_9460);
nand U9541 (N_9541,N_9306,N_9124);
nand U9542 (N_9542,N_9445,N_9330);
nand U9543 (N_9543,N_9251,N_9092);
and U9544 (N_9544,N_9472,N_9027);
or U9545 (N_9545,N_9428,N_9085);
or U9546 (N_9546,N_9289,N_9151);
and U9547 (N_9547,N_9188,N_9357);
nand U9548 (N_9548,N_9290,N_9262);
nor U9549 (N_9549,N_9220,N_9077);
nor U9550 (N_9550,N_9208,N_9104);
or U9551 (N_9551,N_9406,N_9225);
nor U9552 (N_9552,N_9187,N_9288);
xor U9553 (N_9553,N_9038,N_9058);
xnor U9554 (N_9554,N_9024,N_9018);
and U9555 (N_9555,N_9122,N_9436);
nor U9556 (N_9556,N_9240,N_9114);
nand U9557 (N_9557,N_9174,N_9405);
and U9558 (N_9558,N_9373,N_9239);
nand U9559 (N_9559,N_9040,N_9202);
nand U9560 (N_9560,N_9341,N_9103);
or U9561 (N_9561,N_9008,N_9229);
nand U9562 (N_9562,N_9019,N_9455);
nor U9563 (N_9563,N_9003,N_9474);
and U9564 (N_9564,N_9172,N_9055);
and U9565 (N_9565,N_9012,N_9490);
nand U9566 (N_9566,N_9110,N_9331);
and U9567 (N_9567,N_9180,N_9334);
nor U9568 (N_9568,N_9209,N_9217);
nor U9569 (N_9569,N_9448,N_9157);
nand U9570 (N_9570,N_9468,N_9056);
nand U9571 (N_9571,N_9044,N_9268);
and U9572 (N_9572,N_9492,N_9001);
nand U9573 (N_9573,N_9062,N_9261);
and U9574 (N_9574,N_9446,N_9199);
nand U9575 (N_9575,N_9310,N_9393);
nand U9576 (N_9576,N_9338,N_9016);
xnor U9577 (N_9577,N_9241,N_9344);
and U9578 (N_9578,N_9382,N_9255);
and U9579 (N_9579,N_9152,N_9471);
xor U9580 (N_9580,N_9115,N_9311);
xor U9581 (N_9581,N_9447,N_9080);
nand U9582 (N_9582,N_9285,N_9011);
xor U9583 (N_9583,N_9109,N_9061);
and U9584 (N_9584,N_9482,N_9166);
and U9585 (N_9585,N_9073,N_9129);
nand U9586 (N_9586,N_9034,N_9132);
nor U9587 (N_9587,N_9093,N_9102);
xor U9588 (N_9588,N_9247,N_9060);
nand U9589 (N_9589,N_9269,N_9475);
nand U9590 (N_9590,N_9192,N_9023);
and U9591 (N_9591,N_9270,N_9171);
and U9592 (N_9592,N_9312,N_9150);
nand U9593 (N_9593,N_9299,N_9082);
nor U9594 (N_9594,N_9458,N_9135);
or U9595 (N_9595,N_9244,N_9319);
or U9596 (N_9596,N_9211,N_9466);
xnor U9597 (N_9597,N_9195,N_9036);
and U9598 (N_9598,N_9302,N_9399);
nor U9599 (N_9599,N_9079,N_9469);
nor U9600 (N_9600,N_9444,N_9232);
and U9601 (N_9601,N_9291,N_9176);
and U9602 (N_9602,N_9321,N_9175);
or U9603 (N_9603,N_9286,N_9017);
and U9604 (N_9604,N_9013,N_9162);
and U9605 (N_9605,N_9361,N_9304);
or U9606 (N_9606,N_9142,N_9048);
and U9607 (N_9607,N_9378,N_9462);
nor U9608 (N_9608,N_9052,N_9189);
or U9609 (N_9609,N_9190,N_9230);
xnor U9610 (N_9610,N_9158,N_9427);
and U9611 (N_9611,N_9207,N_9078);
nand U9612 (N_9612,N_9185,N_9496);
or U9613 (N_9613,N_9238,N_9410);
nand U9614 (N_9614,N_9067,N_9303);
or U9615 (N_9615,N_9298,N_9032);
xor U9616 (N_9616,N_9053,N_9213);
nor U9617 (N_9617,N_9029,N_9293);
nor U9618 (N_9618,N_9392,N_9435);
and U9619 (N_9619,N_9325,N_9348);
nand U9620 (N_9620,N_9368,N_9258);
nor U9621 (N_9621,N_9300,N_9315);
xor U9622 (N_9622,N_9453,N_9497);
or U9623 (N_9623,N_9116,N_9374);
or U9624 (N_9624,N_9429,N_9146);
or U9625 (N_9625,N_9354,N_9485);
and U9626 (N_9626,N_9133,N_9327);
xor U9627 (N_9627,N_9028,N_9409);
and U9628 (N_9628,N_9163,N_9169);
or U9629 (N_9629,N_9130,N_9441);
nor U9630 (N_9630,N_9181,N_9096);
xnor U9631 (N_9631,N_9273,N_9477);
and U9632 (N_9632,N_9476,N_9186);
nor U9633 (N_9633,N_9025,N_9423);
nor U9634 (N_9634,N_9486,N_9194);
and U9635 (N_9635,N_9483,N_9349);
or U9636 (N_9636,N_9254,N_9165);
nor U9637 (N_9637,N_9307,N_9193);
nand U9638 (N_9638,N_9366,N_9353);
and U9639 (N_9639,N_9314,N_9416);
nor U9640 (N_9640,N_9227,N_9414);
xor U9641 (N_9641,N_9385,N_9156);
or U9642 (N_9642,N_9161,N_9400);
xor U9643 (N_9643,N_9280,N_9363);
or U9644 (N_9644,N_9223,N_9305);
xnor U9645 (N_9645,N_9168,N_9437);
nor U9646 (N_9646,N_9113,N_9432);
nor U9647 (N_9647,N_9141,N_9440);
xnor U9648 (N_9648,N_9235,N_9206);
nand U9649 (N_9649,N_9332,N_9351);
and U9650 (N_9650,N_9420,N_9371);
and U9651 (N_9651,N_9418,N_9030);
nor U9652 (N_9652,N_9043,N_9140);
xor U9653 (N_9653,N_9277,N_9380);
xnor U9654 (N_9654,N_9345,N_9342);
nand U9655 (N_9655,N_9249,N_9045);
nor U9656 (N_9656,N_9010,N_9069);
and U9657 (N_9657,N_9072,N_9257);
nand U9658 (N_9658,N_9362,N_9179);
nand U9659 (N_9659,N_9395,N_9105);
xor U9660 (N_9660,N_9478,N_9294);
xnor U9661 (N_9661,N_9450,N_9279);
nand U9662 (N_9662,N_9022,N_9148);
xor U9663 (N_9663,N_9042,N_9340);
xor U9664 (N_9664,N_9170,N_9136);
xnor U9665 (N_9665,N_9498,N_9390);
or U9666 (N_9666,N_9087,N_9066);
nand U9667 (N_9667,N_9411,N_9107);
nand U9668 (N_9668,N_9083,N_9095);
nor U9669 (N_9669,N_9118,N_9320);
and U9670 (N_9670,N_9183,N_9276);
nand U9671 (N_9671,N_9317,N_9143);
nand U9672 (N_9672,N_9245,N_9167);
nor U9673 (N_9673,N_9329,N_9074);
xnor U9674 (N_9674,N_9356,N_9394);
xnor U9675 (N_9675,N_9004,N_9246);
or U9676 (N_9676,N_9387,N_9063);
and U9677 (N_9677,N_9059,N_9352);
and U9678 (N_9678,N_9049,N_9210);
and U9679 (N_9679,N_9197,N_9046);
and U9680 (N_9680,N_9057,N_9484);
nand U9681 (N_9681,N_9369,N_9318);
and U9682 (N_9682,N_9283,N_9403);
xor U9683 (N_9683,N_9098,N_9430);
nor U9684 (N_9684,N_9084,N_9364);
nand U9685 (N_9685,N_9054,N_9360);
nor U9686 (N_9686,N_9326,N_9037);
and U9687 (N_9687,N_9234,N_9120);
nand U9688 (N_9688,N_9343,N_9191);
nand U9689 (N_9689,N_9454,N_9144);
nor U9690 (N_9690,N_9009,N_9216);
xnor U9691 (N_9691,N_9108,N_9480);
nand U9692 (N_9692,N_9370,N_9433);
nor U9693 (N_9693,N_9421,N_9389);
xnor U9694 (N_9694,N_9489,N_9296);
and U9695 (N_9695,N_9274,N_9164);
and U9696 (N_9696,N_9375,N_9099);
and U9697 (N_9697,N_9424,N_9000);
and U9698 (N_9698,N_9425,N_9050);
and U9699 (N_9699,N_9218,N_9035);
nor U9700 (N_9700,N_9263,N_9076);
or U9701 (N_9701,N_9426,N_9266);
or U9702 (N_9702,N_9449,N_9149);
xor U9703 (N_9703,N_9123,N_9125);
nand U9704 (N_9704,N_9041,N_9452);
or U9705 (N_9705,N_9015,N_9401);
xor U9706 (N_9706,N_9282,N_9419);
xnor U9707 (N_9707,N_9367,N_9100);
nor U9708 (N_9708,N_9324,N_9204);
xnor U9709 (N_9709,N_9159,N_9336);
or U9710 (N_9710,N_9248,N_9214);
nand U9711 (N_9711,N_9089,N_9119);
or U9712 (N_9712,N_9358,N_9402);
and U9713 (N_9713,N_9039,N_9075);
xnor U9714 (N_9714,N_9081,N_9442);
nand U9715 (N_9715,N_9128,N_9097);
xnor U9716 (N_9716,N_9301,N_9221);
nand U9717 (N_9717,N_9006,N_9091);
and U9718 (N_9718,N_9237,N_9242);
nor U9719 (N_9719,N_9002,N_9337);
xor U9720 (N_9720,N_9201,N_9020);
and U9721 (N_9721,N_9335,N_9465);
nor U9722 (N_9722,N_9309,N_9347);
and U9723 (N_9723,N_9145,N_9131);
or U9724 (N_9724,N_9065,N_9265);
xnor U9725 (N_9725,N_9260,N_9350);
nor U9726 (N_9726,N_9160,N_9153);
xor U9727 (N_9727,N_9438,N_9493);
or U9728 (N_9728,N_9112,N_9007);
and U9729 (N_9729,N_9147,N_9308);
nand U9730 (N_9730,N_9443,N_9479);
nor U9731 (N_9731,N_9212,N_9281);
and U9732 (N_9732,N_9271,N_9224);
nor U9733 (N_9733,N_9384,N_9386);
xnor U9734 (N_9734,N_9256,N_9292);
and U9735 (N_9735,N_9233,N_9494);
nor U9736 (N_9736,N_9264,N_9316);
nor U9737 (N_9737,N_9297,N_9094);
xor U9738 (N_9738,N_9259,N_9231);
and U9739 (N_9739,N_9068,N_9154);
nor U9740 (N_9740,N_9322,N_9473);
and U9741 (N_9741,N_9173,N_9451);
or U9742 (N_9742,N_9434,N_9355);
or U9743 (N_9743,N_9461,N_9470);
nor U9744 (N_9744,N_9090,N_9088);
nand U9745 (N_9745,N_9417,N_9415);
or U9746 (N_9746,N_9491,N_9215);
or U9747 (N_9747,N_9134,N_9222);
xnor U9748 (N_9748,N_9412,N_9372);
nor U9749 (N_9749,N_9456,N_9121);
or U9750 (N_9750,N_9308,N_9234);
or U9751 (N_9751,N_9305,N_9231);
and U9752 (N_9752,N_9200,N_9261);
nand U9753 (N_9753,N_9142,N_9379);
nand U9754 (N_9754,N_9053,N_9331);
or U9755 (N_9755,N_9025,N_9054);
nand U9756 (N_9756,N_9281,N_9365);
nand U9757 (N_9757,N_9343,N_9018);
nand U9758 (N_9758,N_9484,N_9225);
or U9759 (N_9759,N_9491,N_9197);
and U9760 (N_9760,N_9263,N_9426);
nand U9761 (N_9761,N_9365,N_9096);
and U9762 (N_9762,N_9067,N_9120);
and U9763 (N_9763,N_9407,N_9127);
nor U9764 (N_9764,N_9043,N_9242);
and U9765 (N_9765,N_9225,N_9420);
and U9766 (N_9766,N_9004,N_9044);
nor U9767 (N_9767,N_9031,N_9046);
and U9768 (N_9768,N_9152,N_9223);
nor U9769 (N_9769,N_9224,N_9373);
or U9770 (N_9770,N_9106,N_9224);
and U9771 (N_9771,N_9413,N_9410);
and U9772 (N_9772,N_9421,N_9202);
nand U9773 (N_9773,N_9166,N_9084);
or U9774 (N_9774,N_9318,N_9340);
and U9775 (N_9775,N_9484,N_9195);
or U9776 (N_9776,N_9161,N_9120);
or U9777 (N_9777,N_9080,N_9292);
and U9778 (N_9778,N_9095,N_9263);
or U9779 (N_9779,N_9100,N_9190);
and U9780 (N_9780,N_9378,N_9149);
nand U9781 (N_9781,N_9377,N_9137);
and U9782 (N_9782,N_9362,N_9130);
xnor U9783 (N_9783,N_9294,N_9418);
nand U9784 (N_9784,N_9438,N_9362);
xnor U9785 (N_9785,N_9475,N_9315);
nor U9786 (N_9786,N_9211,N_9230);
nor U9787 (N_9787,N_9137,N_9465);
and U9788 (N_9788,N_9429,N_9172);
xnor U9789 (N_9789,N_9015,N_9460);
nor U9790 (N_9790,N_9098,N_9383);
and U9791 (N_9791,N_9180,N_9052);
nand U9792 (N_9792,N_9083,N_9351);
nand U9793 (N_9793,N_9342,N_9036);
xnor U9794 (N_9794,N_9043,N_9149);
nor U9795 (N_9795,N_9435,N_9036);
nand U9796 (N_9796,N_9059,N_9213);
xor U9797 (N_9797,N_9283,N_9221);
nand U9798 (N_9798,N_9463,N_9263);
nand U9799 (N_9799,N_9472,N_9178);
or U9800 (N_9800,N_9334,N_9125);
and U9801 (N_9801,N_9144,N_9311);
or U9802 (N_9802,N_9077,N_9249);
nand U9803 (N_9803,N_9389,N_9447);
nor U9804 (N_9804,N_9497,N_9226);
or U9805 (N_9805,N_9356,N_9218);
nor U9806 (N_9806,N_9468,N_9159);
xor U9807 (N_9807,N_9242,N_9317);
xor U9808 (N_9808,N_9395,N_9019);
xnor U9809 (N_9809,N_9494,N_9474);
and U9810 (N_9810,N_9476,N_9185);
nor U9811 (N_9811,N_9319,N_9251);
xnor U9812 (N_9812,N_9335,N_9251);
or U9813 (N_9813,N_9239,N_9096);
and U9814 (N_9814,N_9161,N_9265);
xor U9815 (N_9815,N_9080,N_9307);
nor U9816 (N_9816,N_9336,N_9434);
xor U9817 (N_9817,N_9023,N_9467);
nor U9818 (N_9818,N_9457,N_9432);
or U9819 (N_9819,N_9265,N_9295);
xor U9820 (N_9820,N_9138,N_9386);
nor U9821 (N_9821,N_9087,N_9421);
or U9822 (N_9822,N_9062,N_9250);
xnor U9823 (N_9823,N_9498,N_9275);
xor U9824 (N_9824,N_9485,N_9326);
nand U9825 (N_9825,N_9445,N_9499);
and U9826 (N_9826,N_9471,N_9332);
or U9827 (N_9827,N_9052,N_9295);
and U9828 (N_9828,N_9067,N_9394);
nand U9829 (N_9829,N_9017,N_9031);
and U9830 (N_9830,N_9249,N_9288);
or U9831 (N_9831,N_9101,N_9104);
xnor U9832 (N_9832,N_9329,N_9090);
nand U9833 (N_9833,N_9367,N_9252);
nand U9834 (N_9834,N_9287,N_9015);
nand U9835 (N_9835,N_9333,N_9377);
or U9836 (N_9836,N_9400,N_9435);
nor U9837 (N_9837,N_9290,N_9494);
or U9838 (N_9838,N_9242,N_9011);
nand U9839 (N_9839,N_9184,N_9070);
nor U9840 (N_9840,N_9129,N_9057);
and U9841 (N_9841,N_9402,N_9080);
and U9842 (N_9842,N_9291,N_9385);
xor U9843 (N_9843,N_9142,N_9244);
nand U9844 (N_9844,N_9431,N_9151);
nor U9845 (N_9845,N_9196,N_9247);
xor U9846 (N_9846,N_9495,N_9498);
and U9847 (N_9847,N_9438,N_9005);
or U9848 (N_9848,N_9387,N_9404);
nand U9849 (N_9849,N_9166,N_9316);
or U9850 (N_9850,N_9246,N_9060);
and U9851 (N_9851,N_9154,N_9161);
and U9852 (N_9852,N_9211,N_9052);
or U9853 (N_9853,N_9431,N_9271);
and U9854 (N_9854,N_9373,N_9031);
nor U9855 (N_9855,N_9108,N_9341);
and U9856 (N_9856,N_9264,N_9391);
and U9857 (N_9857,N_9469,N_9140);
nand U9858 (N_9858,N_9211,N_9336);
and U9859 (N_9859,N_9307,N_9402);
or U9860 (N_9860,N_9377,N_9194);
nand U9861 (N_9861,N_9299,N_9237);
nand U9862 (N_9862,N_9293,N_9365);
nand U9863 (N_9863,N_9417,N_9004);
nand U9864 (N_9864,N_9469,N_9151);
nand U9865 (N_9865,N_9474,N_9026);
and U9866 (N_9866,N_9023,N_9319);
xor U9867 (N_9867,N_9260,N_9160);
and U9868 (N_9868,N_9328,N_9483);
and U9869 (N_9869,N_9040,N_9439);
nand U9870 (N_9870,N_9302,N_9362);
xor U9871 (N_9871,N_9407,N_9346);
and U9872 (N_9872,N_9081,N_9162);
nand U9873 (N_9873,N_9472,N_9403);
xnor U9874 (N_9874,N_9145,N_9478);
nor U9875 (N_9875,N_9257,N_9461);
or U9876 (N_9876,N_9016,N_9004);
xor U9877 (N_9877,N_9226,N_9066);
or U9878 (N_9878,N_9332,N_9110);
xor U9879 (N_9879,N_9311,N_9482);
nor U9880 (N_9880,N_9059,N_9438);
and U9881 (N_9881,N_9030,N_9186);
nand U9882 (N_9882,N_9490,N_9242);
and U9883 (N_9883,N_9382,N_9268);
or U9884 (N_9884,N_9302,N_9157);
or U9885 (N_9885,N_9162,N_9230);
nor U9886 (N_9886,N_9485,N_9215);
or U9887 (N_9887,N_9368,N_9456);
nor U9888 (N_9888,N_9359,N_9219);
nor U9889 (N_9889,N_9076,N_9355);
xor U9890 (N_9890,N_9241,N_9016);
xor U9891 (N_9891,N_9007,N_9364);
or U9892 (N_9892,N_9109,N_9277);
or U9893 (N_9893,N_9196,N_9322);
xor U9894 (N_9894,N_9095,N_9092);
nand U9895 (N_9895,N_9012,N_9170);
and U9896 (N_9896,N_9276,N_9291);
and U9897 (N_9897,N_9039,N_9069);
or U9898 (N_9898,N_9317,N_9046);
and U9899 (N_9899,N_9307,N_9105);
xnor U9900 (N_9900,N_9467,N_9395);
and U9901 (N_9901,N_9092,N_9493);
and U9902 (N_9902,N_9226,N_9164);
or U9903 (N_9903,N_9097,N_9227);
nand U9904 (N_9904,N_9370,N_9235);
nand U9905 (N_9905,N_9126,N_9150);
nand U9906 (N_9906,N_9347,N_9315);
nand U9907 (N_9907,N_9360,N_9105);
or U9908 (N_9908,N_9445,N_9494);
nand U9909 (N_9909,N_9361,N_9171);
nand U9910 (N_9910,N_9330,N_9468);
xnor U9911 (N_9911,N_9293,N_9323);
nand U9912 (N_9912,N_9168,N_9267);
or U9913 (N_9913,N_9369,N_9310);
nor U9914 (N_9914,N_9475,N_9390);
and U9915 (N_9915,N_9339,N_9247);
nand U9916 (N_9916,N_9205,N_9413);
nand U9917 (N_9917,N_9260,N_9110);
nor U9918 (N_9918,N_9197,N_9069);
and U9919 (N_9919,N_9050,N_9104);
xnor U9920 (N_9920,N_9234,N_9294);
nand U9921 (N_9921,N_9452,N_9154);
and U9922 (N_9922,N_9069,N_9311);
nand U9923 (N_9923,N_9394,N_9075);
or U9924 (N_9924,N_9100,N_9091);
or U9925 (N_9925,N_9076,N_9472);
xor U9926 (N_9926,N_9345,N_9035);
nor U9927 (N_9927,N_9003,N_9002);
xor U9928 (N_9928,N_9366,N_9395);
nand U9929 (N_9929,N_9433,N_9441);
and U9930 (N_9930,N_9106,N_9228);
and U9931 (N_9931,N_9229,N_9477);
xnor U9932 (N_9932,N_9215,N_9174);
and U9933 (N_9933,N_9193,N_9185);
or U9934 (N_9934,N_9473,N_9349);
xor U9935 (N_9935,N_9431,N_9452);
and U9936 (N_9936,N_9209,N_9311);
nand U9937 (N_9937,N_9240,N_9260);
and U9938 (N_9938,N_9482,N_9325);
nor U9939 (N_9939,N_9217,N_9488);
nand U9940 (N_9940,N_9203,N_9389);
nor U9941 (N_9941,N_9097,N_9463);
nor U9942 (N_9942,N_9130,N_9160);
nor U9943 (N_9943,N_9020,N_9279);
and U9944 (N_9944,N_9422,N_9306);
nor U9945 (N_9945,N_9338,N_9313);
nor U9946 (N_9946,N_9027,N_9495);
and U9947 (N_9947,N_9165,N_9006);
and U9948 (N_9948,N_9398,N_9022);
and U9949 (N_9949,N_9007,N_9477);
and U9950 (N_9950,N_9134,N_9329);
xnor U9951 (N_9951,N_9353,N_9058);
or U9952 (N_9952,N_9347,N_9363);
nand U9953 (N_9953,N_9497,N_9242);
or U9954 (N_9954,N_9062,N_9337);
and U9955 (N_9955,N_9374,N_9465);
or U9956 (N_9956,N_9177,N_9328);
nor U9957 (N_9957,N_9272,N_9160);
nor U9958 (N_9958,N_9228,N_9323);
nor U9959 (N_9959,N_9014,N_9088);
nand U9960 (N_9960,N_9359,N_9174);
or U9961 (N_9961,N_9380,N_9032);
or U9962 (N_9962,N_9448,N_9268);
nor U9963 (N_9963,N_9473,N_9433);
xor U9964 (N_9964,N_9482,N_9180);
xnor U9965 (N_9965,N_9018,N_9304);
nor U9966 (N_9966,N_9331,N_9026);
or U9967 (N_9967,N_9191,N_9288);
and U9968 (N_9968,N_9003,N_9360);
nand U9969 (N_9969,N_9150,N_9071);
xor U9970 (N_9970,N_9127,N_9380);
and U9971 (N_9971,N_9211,N_9158);
xor U9972 (N_9972,N_9047,N_9325);
nand U9973 (N_9973,N_9098,N_9091);
nor U9974 (N_9974,N_9128,N_9298);
nor U9975 (N_9975,N_9032,N_9163);
and U9976 (N_9976,N_9242,N_9472);
and U9977 (N_9977,N_9347,N_9210);
nand U9978 (N_9978,N_9430,N_9034);
and U9979 (N_9979,N_9142,N_9320);
xnor U9980 (N_9980,N_9138,N_9339);
xnor U9981 (N_9981,N_9265,N_9312);
or U9982 (N_9982,N_9129,N_9314);
nand U9983 (N_9983,N_9491,N_9270);
and U9984 (N_9984,N_9154,N_9268);
or U9985 (N_9985,N_9090,N_9150);
xnor U9986 (N_9986,N_9088,N_9290);
and U9987 (N_9987,N_9268,N_9443);
nand U9988 (N_9988,N_9378,N_9148);
or U9989 (N_9989,N_9238,N_9344);
or U9990 (N_9990,N_9256,N_9479);
nand U9991 (N_9991,N_9454,N_9447);
nor U9992 (N_9992,N_9288,N_9009);
and U9993 (N_9993,N_9223,N_9145);
xnor U9994 (N_9994,N_9358,N_9278);
nand U9995 (N_9995,N_9458,N_9107);
xnor U9996 (N_9996,N_9325,N_9294);
nand U9997 (N_9997,N_9319,N_9125);
xnor U9998 (N_9998,N_9280,N_9442);
xor U9999 (N_9999,N_9151,N_9272);
nand U10000 (N_10000,N_9542,N_9749);
or U10001 (N_10001,N_9680,N_9660);
or U10002 (N_10002,N_9616,N_9653);
xnor U10003 (N_10003,N_9772,N_9933);
and U10004 (N_10004,N_9605,N_9964);
nand U10005 (N_10005,N_9826,N_9587);
xor U10006 (N_10006,N_9619,N_9506);
nor U10007 (N_10007,N_9716,N_9531);
and U10008 (N_10008,N_9567,N_9645);
nand U10009 (N_10009,N_9612,N_9811);
and U10010 (N_10010,N_9953,N_9800);
nand U10011 (N_10011,N_9941,N_9902);
nand U10012 (N_10012,N_9701,N_9508);
and U10013 (N_10013,N_9685,N_9980);
or U10014 (N_10014,N_9971,N_9954);
and U10015 (N_10015,N_9895,N_9924);
nor U10016 (N_10016,N_9695,N_9607);
nor U10017 (N_10017,N_9593,N_9982);
or U10018 (N_10018,N_9650,N_9577);
and U10019 (N_10019,N_9925,N_9763);
or U10020 (N_10020,N_9875,N_9665);
nor U10021 (N_10021,N_9663,N_9718);
nor U10022 (N_10022,N_9684,N_9598);
xnor U10023 (N_10023,N_9503,N_9519);
nand U10024 (N_10024,N_9602,N_9702);
nor U10025 (N_10025,N_9706,N_9719);
nand U10026 (N_10026,N_9740,N_9891);
or U10027 (N_10027,N_9956,N_9700);
nand U10028 (N_10028,N_9734,N_9876);
or U10029 (N_10029,N_9563,N_9546);
and U10030 (N_10030,N_9738,N_9972);
xnor U10031 (N_10031,N_9750,N_9929);
or U10032 (N_10032,N_9640,N_9917);
or U10033 (N_10033,N_9785,N_9830);
and U10034 (N_10034,N_9769,N_9987);
nor U10035 (N_10035,N_9687,N_9812);
or U10036 (N_10036,N_9720,N_9921);
xnor U10037 (N_10037,N_9864,N_9568);
or U10038 (N_10038,N_9910,N_9846);
and U10039 (N_10039,N_9938,N_9809);
nor U10040 (N_10040,N_9784,N_9990);
or U10041 (N_10041,N_9621,N_9748);
nor U10042 (N_10042,N_9544,N_9714);
xor U10043 (N_10043,N_9948,N_9996);
nand U10044 (N_10044,N_9855,N_9658);
nor U10045 (N_10045,N_9713,N_9761);
nand U10046 (N_10046,N_9558,N_9777);
nand U10047 (N_10047,N_9952,N_9881);
and U10048 (N_10048,N_9535,N_9973);
xnor U10049 (N_10049,N_9967,N_9501);
nor U10050 (N_10050,N_9538,N_9798);
and U10051 (N_10051,N_9717,N_9509);
and U10052 (N_10052,N_9984,N_9868);
and U10053 (N_10053,N_9715,N_9553);
nor U10054 (N_10054,N_9835,N_9795);
or U10055 (N_10055,N_9975,N_9656);
or U10056 (N_10056,N_9574,N_9634);
or U10057 (N_10057,N_9570,N_9675);
nor U10058 (N_10058,N_9859,N_9500);
or U10059 (N_10059,N_9539,N_9974);
xnor U10060 (N_10060,N_9869,N_9609);
and U10061 (N_10061,N_9960,N_9521);
nand U10062 (N_10062,N_9721,N_9683);
nor U10063 (N_10063,N_9594,N_9635);
or U10064 (N_10064,N_9845,N_9833);
nand U10065 (N_10065,N_9927,N_9779);
nor U10066 (N_10066,N_9930,N_9743);
and U10067 (N_10067,N_9644,N_9912);
nand U10068 (N_10068,N_9918,N_9831);
xnor U10069 (N_10069,N_9828,N_9551);
and U10070 (N_10070,N_9857,N_9856);
nand U10071 (N_10071,N_9937,N_9591);
or U10072 (N_10072,N_9518,N_9822);
xnor U10073 (N_10073,N_9988,N_9842);
and U10074 (N_10074,N_9911,N_9699);
and U10075 (N_10075,N_9914,N_9642);
nand U10076 (N_10076,N_9969,N_9810);
xnor U10077 (N_10077,N_9849,N_9801);
and U10078 (N_10078,N_9628,N_9999);
and U10079 (N_10079,N_9746,N_9620);
nand U10080 (N_10080,N_9780,N_9540);
nor U10081 (N_10081,N_9981,N_9840);
xor U10082 (N_10082,N_9808,N_9708);
xnor U10083 (N_10083,N_9890,N_9992);
or U10084 (N_10084,N_9589,N_9916);
nor U10085 (N_10085,N_9732,N_9892);
nor U10086 (N_10086,N_9580,N_9958);
nand U10087 (N_10087,N_9636,N_9806);
nor U10088 (N_10088,N_9727,N_9774);
xor U10089 (N_10089,N_9843,N_9555);
xnor U10090 (N_10090,N_9829,N_9860);
nor U10091 (N_10091,N_9782,N_9586);
nor U10092 (N_10092,N_9511,N_9571);
and U10093 (N_10093,N_9565,N_9704);
and U10094 (N_10094,N_9652,N_9976);
nor U10095 (N_10095,N_9893,N_9961);
or U10096 (N_10096,N_9900,N_9994);
or U10097 (N_10097,N_9936,N_9686);
nor U10098 (N_10098,N_9677,N_9670);
nand U10099 (N_10099,N_9804,N_9525);
xor U10100 (N_10100,N_9932,N_9703);
or U10101 (N_10101,N_9898,N_9608);
nor U10102 (N_10102,N_9659,N_9903);
nor U10103 (N_10103,N_9541,N_9852);
nand U10104 (N_10104,N_9696,N_9611);
nand U10105 (N_10105,N_9585,N_9579);
or U10106 (N_10106,N_9604,N_9943);
xor U10107 (N_10107,N_9643,N_9873);
or U10108 (N_10108,N_9775,N_9639);
nand U10109 (N_10109,N_9764,N_9671);
nor U10110 (N_10110,N_9882,N_9783);
nand U10111 (N_10111,N_9631,N_9790);
xnor U10112 (N_10112,N_9979,N_9517);
xor U10113 (N_10113,N_9633,N_9865);
nor U10114 (N_10114,N_9733,N_9588);
nand U10115 (N_10115,N_9818,N_9934);
and U10116 (N_10116,N_9600,N_9747);
or U10117 (N_10117,N_9854,N_9786);
or U10118 (N_10118,N_9926,N_9705);
and U10119 (N_10119,N_9897,N_9931);
or U10120 (N_10120,N_9877,N_9759);
or U10121 (N_10121,N_9836,N_9504);
nand U10122 (N_10122,N_9762,N_9618);
nor U10123 (N_10123,N_9613,N_9879);
or U10124 (N_10124,N_9978,N_9906);
xnor U10125 (N_10125,N_9824,N_9723);
xnor U10126 (N_10126,N_9625,N_9657);
or U10127 (N_10127,N_9524,N_9851);
or U10128 (N_10128,N_9788,N_9655);
or U10129 (N_10129,N_9742,N_9622);
or U10130 (N_10130,N_9681,N_9942);
nand U10131 (N_10131,N_9512,N_9582);
xor U10132 (N_10132,N_9710,N_9729);
xnor U10133 (N_10133,N_9691,N_9887);
or U10134 (N_10134,N_9737,N_9970);
nor U10135 (N_10135,N_9726,N_9615);
and U10136 (N_10136,N_9692,N_9949);
or U10137 (N_10137,N_9673,N_9610);
nor U10138 (N_10138,N_9522,N_9755);
xor U10139 (N_10139,N_9977,N_9799);
nor U10140 (N_10140,N_9915,N_9819);
nand U10141 (N_10141,N_9662,N_9814);
and U10142 (N_10142,N_9690,N_9728);
nand U10143 (N_10143,N_9821,N_9638);
or U10144 (N_10144,N_9813,N_9792);
and U10145 (N_10145,N_9739,N_9534);
xnor U10146 (N_10146,N_9666,N_9678);
nand U10147 (N_10147,N_9507,N_9794);
xnor U10148 (N_10148,N_9510,N_9989);
and U10149 (N_10149,N_9965,N_9664);
nand U10150 (N_10150,N_9709,N_9844);
or U10151 (N_10151,N_9584,N_9575);
or U10152 (N_10152,N_9871,N_9781);
and U10153 (N_10153,N_9847,N_9793);
xnor U10154 (N_10154,N_9791,N_9532);
nand U10155 (N_10155,N_9564,N_9880);
nor U10156 (N_10156,N_9955,N_9923);
nor U10157 (N_10157,N_9735,N_9578);
nand U10158 (N_10158,N_9773,N_9878);
and U10159 (N_10159,N_9654,N_9566);
or U10160 (N_10160,N_9672,N_9862);
nand U10161 (N_10161,N_9533,N_9630);
nand U10162 (N_10162,N_9968,N_9632);
nor U10163 (N_10163,N_9523,N_9668);
nor U10164 (N_10164,N_9629,N_9946);
nand U10165 (N_10165,N_9527,N_9957);
nor U10166 (N_10166,N_9920,N_9827);
nand U10167 (N_10167,N_9816,N_9516);
nor U10168 (N_10168,N_9647,N_9866);
and U10169 (N_10169,N_9861,N_9805);
or U10170 (N_10170,N_9627,N_9557);
and U10171 (N_10171,N_9637,N_9985);
nor U10172 (N_10172,N_9530,N_9757);
and U10173 (N_10173,N_9597,N_9939);
and U10174 (N_10174,N_9590,N_9682);
and U10175 (N_10175,N_9765,N_9803);
xor U10176 (N_10176,N_9698,N_9730);
nand U10177 (N_10177,N_9641,N_9919);
or U10178 (N_10178,N_9559,N_9562);
nand U10179 (N_10179,N_9513,N_9909);
or U10180 (N_10180,N_9863,N_9603);
xor U10181 (N_10181,N_9888,N_9502);
or U10182 (N_10182,N_9679,N_9547);
nand U10183 (N_10183,N_9731,N_9736);
xnor U10184 (N_10184,N_9561,N_9697);
or U10185 (N_10185,N_9741,N_9991);
nand U10186 (N_10186,N_9537,N_9676);
nand U10187 (N_10187,N_9935,N_9928);
or U10188 (N_10188,N_9617,N_9867);
or U10189 (N_10189,N_9694,N_9669);
or U10190 (N_10190,N_9581,N_9778);
or U10191 (N_10191,N_9550,N_9688);
or U10192 (N_10192,N_9962,N_9986);
nor U10193 (N_10193,N_9945,N_9908);
and U10194 (N_10194,N_9767,N_9549);
or U10195 (N_10195,N_9815,N_9725);
nand U10196 (N_10196,N_9649,N_9707);
xnor U10197 (N_10197,N_9545,N_9886);
nor U10198 (N_10198,N_9853,N_9839);
or U10199 (N_10199,N_9883,N_9983);
xor U10200 (N_10200,N_9997,N_9848);
nand U10201 (N_10201,N_9722,N_9768);
xor U10202 (N_10202,N_9560,N_9998);
xnor U10203 (N_10203,N_9623,N_9907);
nand U10204 (N_10204,N_9536,N_9624);
and U10205 (N_10205,N_9940,N_9807);
xnor U10206 (N_10206,N_9751,N_9899);
nand U10207 (N_10207,N_9858,N_9894);
nand U10208 (N_10208,N_9959,N_9651);
xor U10209 (N_10209,N_9950,N_9874);
xor U10210 (N_10210,N_9554,N_9797);
or U10211 (N_10211,N_9556,N_9760);
xor U10212 (N_10212,N_9825,N_9648);
nor U10213 (N_10213,N_9817,N_9756);
nand U10214 (N_10214,N_9552,N_9922);
nand U10215 (N_10215,N_9599,N_9766);
and U10216 (N_10216,N_9572,N_9904);
nor U10217 (N_10217,N_9592,N_9884);
xor U10218 (N_10218,N_9947,N_9711);
and U10219 (N_10219,N_9896,N_9712);
xnor U10220 (N_10220,N_9838,N_9520);
nand U10221 (N_10221,N_9913,N_9758);
xnor U10222 (N_10222,N_9951,N_9872);
nand U10223 (N_10223,N_9601,N_9505);
or U10224 (N_10224,N_9529,N_9820);
and U10225 (N_10225,N_9626,N_9514);
or U10226 (N_10226,N_9595,N_9771);
nor U10227 (N_10227,N_9693,N_9841);
nand U10228 (N_10228,N_9832,N_9889);
xor U10229 (N_10229,N_9744,N_9966);
xnor U10230 (N_10230,N_9548,N_9993);
nor U10231 (N_10231,N_9667,N_9543);
or U10232 (N_10232,N_9674,N_9837);
nor U10233 (N_10233,N_9944,N_9569);
xnor U10234 (N_10234,N_9870,N_9796);
or U10235 (N_10235,N_9661,N_9583);
xor U10236 (N_10236,N_9646,N_9526);
nand U10237 (N_10237,N_9905,N_9745);
xor U10238 (N_10238,N_9752,N_9724);
nand U10239 (N_10239,N_9515,N_9528);
nand U10240 (N_10240,N_9787,N_9753);
and U10241 (N_10241,N_9963,N_9850);
and U10242 (N_10242,N_9614,N_9596);
or U10243 (N_10243,N_9770,N_9823);
nor U10244 (N_10244,N_9776,N_9834);
xor U10245 (N_10245,N_9995,N_9789);
or U10246 (N_10246,N_9606,N_9901);
nor U10247 (N_10247,N_9802,N_9573);
xnor U10248 (N_10248,N_9576,N_9689);
nand U10249 (N_10249,N_9754,N_9885);
or U10250 (N_10250,N_9578,N_9880);
nor U10251 (N_10251,N_9689,N_9652);
nor U10252 (N_10252,N_9747,N_9748);
or U10253 (N_10253,N_9825,N_9791);
nor U10254 (N_10254,N_9692,N_9858);
nand U10255 (N_10255,N_9644,N_9516);
or U10256 (N_10256,N_9503,N_9975);
nand U10257 (N_10257,N_9644,N_9997);
nor U10258 (N_10258,N_9937,N_9845);
nor U10259 (N_10259,N_9537,N_9553);
or U10260 (N_10260,N_9532,N_9752);
nor U10261 (N_10261,N_9769,N_9841);
and U10262 (N_10262,N_9612,N_9856);
and U10263 (N_10263,N_9750,N_9680);
and U10264 (N_10264,N_9730,N_9847);
nor U10265 (N_10265,N_9952,N_9705);
and U10266 (N_10266,N_9947,N_9978);
and U10267 (N_10267,N_9653,N_9603);
and U10268 (N_10268,N_9992,N_9981);
nand U10269 (N_10269,N_9715,N_9617);
nand U10270 (N_10270,N_9606,N_9915);
xor U10271 (N_10271,N_9689,N_9797);
xor U10272 (N_10272,N_9853,N_9595);
nor U10273 (N_10273,N_9869,N_9871);
or U10274 (N_10274,N_9753,N_9662);
nor U10275 (N_10275,N_9564,N_9763);
xnor U10276 (N_10276,N_9997,N_9944);
nand U10277 (N_10277,N_9903,N_9683);
or U10278 (N_10278,N_9972,N_9838);
nand U10279 (N_10279,N_9506,N_9873);
and U10280 (N_10280,N_9987,N_9748);
or U10281 (N_10281,N_9877,N_9962);
or U10282 (N_10282,N_9538,N_9996);
and U10283 (N_10283,N_9512,N_9819);
or U10284 (N_10284,N_9708,N_9834);
nand U10285 (N_10285,N_9595,N_9509);
nor U10286 (N_10286,N_9681,N_9917);
nand U10287 (N_10287,N_9589,N_9930);
xnor U10288 (N_10288,N_9987,N_9954);
and U10289 (N_10289,N_9766,N_9821);
nand U10290 (N_10290,N_9723,N_9675);
xnor U10291 (N_10291,N_9825,N_9935);
or U10292 (N_10292,N_9580,N_9535);
xor U10293 (N_10293,N_9913,N_9804);
xor U10294 (N_10294,N_9678,N_9855);
nand U10295 (N_10295,N_9810,N_9872);
or U10296 (N_10296,N_9851,N_9933);
nand U10297 (N_10297,N_9798,N_9905);
nand U10298 (N_10298,N_9649,N_9608);
nor U10299 (N_10299,N_9694,N_9994);
nand U10300 (N_10300,N_9877,N_9996);
nand U10301 (N_10301,N_9989,N_9649);
nor U10302 (N_10302,N_9641,N_9806);
or U10303 (N_10303,N_9776,N_9573);
and U10304 (N_10304,N_9668,N_9913);
and U10305 (N_10305,N_9504,N_9740);
nand U10306 (N_10306,N_9928,N_9584);
or U10307 (N_10307,N_9881,N_9879);
nand U10308 (N_10308,N_9711,N_9551);
xnor U10309 (N_10309,N_9847,N_9691);
or U10310 (N_10310,N_9929,N_9923);
nand U10311 (N_10311,N_9947,N_9721);
or U10312 (N_10312,N_9718,N_9511);
and U10313 (N_10313,N_9645,N_9941);
nand U10314 (N_10314,N_9747,N_9778);
nand U10315 (N_10315,N_9650,N_9786);
xor U10316 (N_10316,N_9939,N_9714);
nor U10317 (N_10317,N_9561,N_9905);
xnor U10318 (N_10318,N_9628,N_9831);
nand U10319 (N_10319,N_9643,N_9800);
nor U10320 (N_10320,N_9870,N_9886);
or U10321 (N_10321,N_9708,N_9860);
nand U10322 (N_10322,N_9982,N_9741);
nor U10323 (N_10323,N_9881,N_9630);
and U10324 (N_10324,N_9888,N_9981);
and U10325 (N_10325,N_9720,N_9767);
nand U10326 (N_10326,N_9778,N_9786);
nand U10327 (N_10327,N_9608,N_9538);
nand U10328 (N_10328,N_9856,N_9761);
nor U10329 (N_10329,N_9621,N_9703);
or U10330 (N_10330,N_9901,N_9664);
nor U10331 (N_10331,N_9785,N_9589);
nand U10332 (N_10332,N_9937,N_9967);
and U10333 (N_10333,N_9800,N_9592);
nand U10334 (N_10334,N_9956,N_9941);
or U10335 (N_10335,N_9620,N_9717);
and U10336 (N_10336,N_9868,N_9672);
or U10337 (N_10337,N_9922,N_9878);
nor U10338 (N_10338,N_9629,N_9993);
or U10339 (N_10339,N_9838,N_9598);
and U10340 (N_10340,N_9901,N_9869);
nand U10341 (N_10341,N_9967,N_9976);
or U10342 (N_10342,N_9842,N_9900);
nand U10343 (N_10343,N_9648,N_9577);
nor U10344 (N_10344,N_9743,N_9991);
xnor U10345 (N_10345,N_9723,N_9851);
nor U10346 (N_10346,N_9971,N_9560);
or U10347 (N_10347,N_9564,N_9895);
xnor U10348 (N_10348,N_9990,N_9925);
and U10349 (N_10349,N_9923,N_9686);
nand U10350 (N_10350,N_9723,N_9706);
nor U10351 (N_10351,N_9510,N_9994);
nor U10352 (N_10352,N_9770,N_9827);
and U10353 (N_10353,N_9770,N_9877);
nand U10354 (N_10354,N_9774,N_9962);
or U10355 (N_10355,N_9858,N_9610);
and U10356 (N_10356,N_9876,N_9689);
or U10357 (N_10357,N_9828,N_9877);
nor U10358 (N_10358,N_9898,N_9800);
and U10359 (N_10359,N_9833,N_9783);
nand U10360 (N_10360,N_9887,N_9895);
and U10361 (N_10361,N_9865,N_9983);
nand U10362 (N_10362,N_9910,N_9647);
or U10363 (N_10363,N_9805,N_9783);
or U10364 (N_10364,N_9962,N_9752);
and U10365 (N_10365,N_9974,N_9661);
nor U10366 (N_10366,N_9669,N_9550);
or U10367 (N_10367,N_9624,N_9817);
nand U10368 (N_10368,N_9635,N_9810);
or U10369 (N_10369,N_9988,N_9849);
nor U10370 (N_10370,N_9958,N_9904);
nor U10371 (N_10371,N_9886,N_9593);
nor U10372 (N_10372,N_9789,N_9709);
and U10373 (N_10373,N_9852,N_9725);
or U10374 (N_10374,N_9727,N_9723);
xnor U10375 (N_10375,N_9532,N_9595);
and U10376 (N_10376,N_9634,N_9936);
nand U10377 (N_10377,N_9815,N_9921);
nor U10378 (N_10378,N_9654,N_9561);
nand U10379 (N_10379,N_9790,N_9923);
and U10380 (N_10380,N_9950,N_9525);
xor U10381 (N_10381,N_9602,N_9628);
xor U10382 (N_10382,N_9795,N_9511);
or U10383 (N_10383,N_9540,N_9604);
nor U10384 (N_10384,N_9574,N_9914);
nand U10385 (N_10385,N_9924,N_9929);
xnor U10386 (N_10386,N_9561,N_9651);
or U10387 (N_10387,N_9835,N_9611);
nor U10388 (N_10388,N_9702,N_9724);
and U10389 (N_10389,N_9768,N_9874);
nand U10390 (N_10390,N_9761,N_9649);
and U10391 (N_10391,N_9896,N_9698);
and U10392 (N_10392,N_9700,N_9655);
and U10393 (N_10393,N_9918,N_9898);
and U10394 (N_10394,N_9968,N_9888);
and U10395 (N_10395,N_9759,N_9545);
nor U10396 (N_10396,N_9513,N_9505);
xnor U10397 (N_10397,N_9698,N_9783);
xor U10398 (N_10398,N_9736,N_9718);
xor U10399 (N_10399,N_9697,N_9851);
xnor U10400 (N_10400,N_9675,N_9690);
or U10401 (N_10401,N_9900,N_9911);
nand U10402 (N_10402,N_9727,N_9981);
xor U10403 (N_10403,N_9584,N_9912);
xnor U10404 (N_10404,N_9893,N_9665);
nand U10405 (N_10405,N_9522,N_9630);
xnor U10406 (N_10406,N_9519,N_9705);
nand U10407 (N_10407,N_9531,N_9891);
xor U10408 (N_10408,N_9770,N_9800);
and U10409 (N_10409,N_9690,N_9759);
xnor U10410 (N_10410,N_9821,N_9784);
nor U10411 (N_10411,N_9733,N_9789);
xnor U10412 (N_10412,N_9539,N_9572);
nand U10413 (N_10413,N_9622,N_9970);
and U10414 (N_10414,N_9600,N_9855);
nor U10415 (N_10415,N_9891,N_9592);
and U10416 (N_10416,N_9786,N_9841);
xnor U10417 (N_10417,N_9524,N_9621);
or U10418 (N_10418,N_9679,N_9506);
xor U10419 (N_10419,N_9958,N_9988);
or U10420 (N_10420,N_9787,N_9590);
and U10421 (N_10421,N_9957,N_9882);
nor U10422 (N_10422,N_9878,N_9630);
or U10423 (N_10423,N_9889,N_9794);
nand U10424 (N_10424,N_9819,N_9563);
and U10425 (N_10425,N_9554,N_9636);
xor U10426 (N_10426,N_9790,N_9504);
and U10427 (N_10427,N_9792,N_9542);
xor U10428 (N_10428,N_9938,N_9793);
nor U10429 (N_10429,N_9826,N_9837);
xor U10430 (N_10430,N_9811,N_9728);
xnor U10431 (N_10431,N_9607,N_9512);
xor U10432 (N_10432,N_9949,N_9907);
or U10433 (N_10433,N_9697,N_9641);
and U10434 (N_10434,N_9753,N_9872);
or U10435 (N_10435,N_9979,N_9835);
nor U10436 (N_10436,N_9684,N_9681);
nor U10437 (N_10437,N_9607,N_9501);
xnor U10438 (N_10438,N_9794,N_9792);
and U10439 (N_10439,N_9870,N_9613);
and U10440 (N_10440,N_9610,N_9978);
or U10441 (N_10441,N_9753,N_9640);
nor U10442 (N_10442,N_9771,N_9819);
nor U10443 (N_10443,N_9950,N_9640);
xor U10444 (N_10444,N_9823,N_9503);
nand U10445 (N_10445,N_9828,N_9902);
and U10446 (N_10446,N_9834,N_9622);
nand U10447 (N_10447,N_9952,N_9930);
xnor U10448 (N_10448,N_9535,N_9527);
xnor U10449 (N_10449,N_9501,N_9880);
nor U10450 (N_10450,N_9845,N_9985);
or U10451 (N_10451,N_9528,N_9539);
nor U10452 (N_10452,N_9949,N_9759);
nor U10453 (N_10453,N_9905,N_9945);
xnor U10454 (N_10454,N_9736,N_9765);
xor U10455 (N_10455,N_9927,N_9880);
nor U10456 (N_10456,N_9670,N_9516);
nor U10457 (N_10457,N_9620,N_9915);
xor U10458 (N_10458,N_9520,N_9989);
nand U10459 (N_10459,N_9680,N_9543);
xnor U10460 (N_10460,N_9762,N_9672);
or U10461 (N_10461,N_9786,N_9717);
and U10462 (N_10462,N_9982,N_9510);
or U10463 (N_10463,N_9992,N_9563);
or U10464 (N_10464,N_9617,N_9813);
and U10465 (N_10465,N_9799,N_9734);
or U10466 (N_10466,N_9839,N_9789);
and U10467 (N_10467,N_9825,N_9543);
and U10468 (N_10468,N_9832,N_9781);
or U10469 (N_10469,N_9734,N_9720);
xnor U10470 (N_10470,N_9535,N_9665);
nor U10471 (N_10471,N_9573,N_9900);
nor U10472 (N_10472,N_9932,N_9503);
xor U10473 (N_10473,N_9555,N_9868);
or U10474 (N_10474,N_9784,N_9834);
nor U10475 (N_10475,N_9981,N_9917);
or U10476 (N_10476,N_9815,N_9841);
nand U10477 (N_10477,N_9860,N_9838);
nand U10478 (N_10478,N_9563,N_9981);
nor U10479 (N_10479,N_9880,N_9566);
xnor U10480 (N_10480,N_9911,N_9781);
nor U10481 (N_10481,N_9742,N_9836);
nor U10482 (N_10482,N_9517,N_9625);
nor U10483 (N_10483,N_9507,N_9762);
xor U10484 (N_10484,N_9769,N_9745);
nor U10485 (N_10485,N_9529,N_9861);
or U10486 (N_10486,N_9500,N_9869);
nand U10487 (N_10487,N_9825,N_9562);
xor U10488 (N_10488,N_9805,N_9741);
or U10489 (N_10489,N_9720,N_9850);
nor U10490 (N_10490,N_9536,N_9905);
nor U10491 (N_10491,N_9990,N_9844);
nor U10492 (N_10492,N_9853,N_9782);
xor U10493 (N_10493,N_9990,N_9711);
nand U10494 (N_10494,N_9796,N_9682);
xor U10495 (N_10495,N_9831,N_9538);
nand U10496 (N_10496,N_9542,N_9783);
nand U10497 (N_10497,N_9553,N_9818);
nor U10498 (N_10498,N_9582,N_9678);
nor U10499 (N_10499,N_9882,N_9832);
nand U10500 (N_10500,N_10213,N_10167);
or U10501 (N_10501,N_10077,N_10411);
nand U10502 (N_10502,N_10138,N_10107);
or U10503 (N_10503,N_10399,N_10208);
nor U10504 (N_10504,N_10016,N_10192);
nor U10505 (N_10505,N_10229,N_10253);
nand U10506 (N_10506,N_10326,N_10439);
or U10507 (N_10507,N_10378,N_10033);
nand U10508 (N_10508,N_10484,N_10174);
xor U10509 (N_10509,N_10460,N_10139);
nand U10510 (N_10510,N_10130,N_10136);
nor U10511 (N_10511,N_10282,N_10267);
nor U10512 (N_10512,N_10092,N_10088);
nand U10513 (N_10513,N_10274,N_10242);
xor U10514 (N_10514,N_10142,N_10472);
nor U10515 (N_10515,N_10100,N_10252);
nand U10516 (N_10516,N_10473,N_10395);
and U10517 (N_10517,N_10367,N_10416);
and U10518 (N_10518,N_10007,N_10161);
or U10519 (N_10519,N_10042,N_10302);
or U10520 (N_10520,N_10384,N_10349);
nor U10521 (N_10521,N_10261,N_10243);
and U10522 (N_10522,N_10178,N_10443);
nor U10523 (N_10523,N_10148,N_10177);
nand U10524 (N_10524,N_10386,N_10227);
nand U10525 (N_10525,N_10280,N_10388);
and U10526 (N_10526,N_10464,N_10097);
nor U10527 (N_10527,N_10478,N_10342);
or U10528 (N_10528,N_10311,N_10036);
nand U10529 (N_10529,N_10245,N_10365);
or U10530 (N_10530,N_10061,N_10423);
nor U10531 (N_10531,N_10249,N_10413);
nor U10532 (N_10532,N_10380,N_10090);
nor U10533 (N_10533,N_10398,N_10043);
or U10534 (N_10534,N_10364,N_10166);
nor U10535 (N_10535,N_10372,N_10465);
xor U10536 (N_10536,N_10412,N_10264);
nand U10537 (N_10537,N_10442,N_10429);
nand U10538 (N_10538,N_10225,N_10308);
or U10539 (N_10539,N_10011,N_10094);
nor U10540 (N_10540,N_10057,N_10405);
and U10541 (N_10541,N_10153,N_10341);
and U10542 (N_10542,N_10029,N_10389);
nor U10543 (N_10543,N_10487,N_10024);
or U10544 (N_10544,N_10068,N_10417);
xnor U10545 (N_10545,N_10294,N_10497);
nor U10546 (N_10546,N_10015,N_10322);
or U10547 (N_10547,N_10231,N_10445);
nand U10548 (N_10548,N_10441,N_10432);
nor U10549 (N_10549,N_10123,N_10209);
xor U10550 (N_10550,N_10408,N_10105);
xnor U10551 (N_10551,N_10397,N_10014);
or U10552 (N_10552,N_10390,N_10205);
or U10553 (N_10553,N_10108,N_10137);
or U10554 (N_10554,N_10430,N_10184);
nand U10555 (N_10555,N_10290,N_10330);
and U10556 (N_10556,N_10495,N_10112);
nor U10557 (N_10557,N_10147,N_10312);
and U10558 (N_10558,N_10296,N_10003);
xor U10559 (N_10559,N_10146,N_10196);
and U10560 (N_10560,N_10496,N_10054);
nand U10561 (N_10561,N_10086,N_10075);
and U10562 (N_10562,N_10391,N_10375);
or U10563 (N_10563,N_10027,N_10292);
xnor U10564 (N_10564,N_10317,N_10045);
or U10565 (N_10565,N_10435,N_10396);
or U10566 (N_10566,N_10345,N_10303);
xor U10567 (N_10567,N_10127,N_10175);
nand U10568 (N_10568,N_10169,N_10255);
nor U10569 (N_10569,N_10216,N_10499);
xor U10570 (N_10570,N_10431,N_10101);
xor U10571 (N_10571,N_10286,N_10369);
nor U10572 (N_10572,N_10293,N_10082);
nand U10573 (N_10573,N_10403,N_10055);
or U10574 (N_10574,N_10450,N_10032);
nand U10575 (N_10575,N_10247,N_10026);
or U10576 (N_10576,N_10006,N_10018);
xor U10577 (N_10577,N_10114,N_10052);
nand U10578 (N_10578,N_10193,N_10474);
or U10579 (N_10579,N_10037,N_10250);
or U10580 (N_10580,N_10228,N_10222);
nand U10581 (N_10581,N_10324,N_10427);
nor U10582 (N_10582,N_10258,N_10093);
nor U10583 (N_10583,N_10218,N_10336);
nor U10584 (N_10584,N_10475,N_10051);
nand U10585 (N_10585,N_10103,N_10220);
nand U10586 (N_10586,N_10272,N_10156);
nand U10587 (N_10587,N_10344,N_10482);
nor U10588 (N_10588,N_10154,N_10201);
and U10589 (N_10589,N_10410,N_10304);
nor U10590 (N_10590,N_10230,N_10362);
xnor U10591 (N_10591,N_10351,N_10115);
and U10592 (N_10592,N_10168,N_10125);
xnor U10593 (N_10593,N_10207,N_10120);
nor U10594 (N_10594,N_10301,N_10260);
xnor U10595 (N_10595,N_10124,N_10102);
nand U10596 (N_10596,N_10279,N_10488);
nor U10597 (N_10597,N_10001,N_10060);
nor U10598 (N_10598,N_10116,N_10238);
xnor U10599 (N_10599,N_10486,N_10240);
or U10600 (N_10600,N_10471,N_10083);
or U10601 (N_10601,N_10234,N_10226);
nor U10602 (N_10602,N_10009,N_10492);
nand U10603 (N_10603,N_10309,N_10407);
or U10604 (N_10604,N_10490,N_10025);
xor U10605 (N_10605,N_10203,N_10109);
nor U10606 (N_10606,N_10098,N_10266);
xor U10607 (N_10607,N_10058,N_10313);
nand U10608 (N_10608,N_10096,N_10182);
nor U10609 (N_10609,N_10382,N_10121);
or U10610 (N_10610,N_10048,N_10299);
nand U10611 (N_10611,N_10318,N_10180);
nor U10612 (N_10612,N_10087,N_10110);
and U10613 (N_10613,N_10067,N_10377);
nand U10614 (N_10614,N_10401,N_10469);
or U10615 (N_10615,N_10359,N_10288);
xnor U10616 (N_10616,N_10425,N_10062);
xnor U10617 (N_10617,N_10409,N_10072);
or U10618 (N_10618,N_10353,N_10485);
nand U10619 (N_10619,N_10119,N_10295);
xor U10620 (N_10620,N_10447,N_10046);
and U10621 (N_10621,N_10004,N_10172);
xor U10622 (N_10622,N_10211,N_10152);
nor U10623 (N_10623,N_10244,N_10204);
or U10624 (N_10624,N_10269,N_10298);
xor U10625 (N_10625,N_10257,N_10337);
nor U10626 (N_10626,N_10106,N_10145);
xnor U10627 (N_10627,N_10481,N_10468);
or U10628 (N_10628,N_10248,N_10104);
xnor U10629 (N_10629,N_10433,N_10289);
or U10630 (N_10630,N_10185,N_10078);
and U10631 (N_10631,N_10348,N_10246);
and U10632 (N_10632,N_10195,N_10002);
and U10633 (N_10633,N_10080,N_10183);
xor U10634 (N_10634,N_10023,N_10385);
or U10635 (N_10635,N_10459,N_10005);
xor U10636 (N_10636,N_10162,N_10189);
and U10637 (N_10637,N_10237,N_10111);
nand U10638 (N_10638,N_10419,N_10360);
xnor U10639 (N_10639,N_10470,N_10436);
and U10640 (N_10640,N_10323,N_10340);
nand U10641 (N_10641,N_10163,N_10448);
and U10642 (N_10642,N_10186,N_10164);
nor U10643 (N_10643,N_10181,N_10347);
nand U10644 (N_10644,N_10035,N_10132);
and U10645 (N_10645,N_10031,N_10453);
nor U10646 (N_10646,N_10066,N_10073);
xor U10647 (N_10647,N_10376,N_10074);
and U10648 (N_10648,N_10297,N_10306);
nor U10649 (N_10649,N_10452,N_10170);
nor U10650 (N_10650,N_10259,N_10118);
xnor U10651 (N_10651,N_10331,N_10489);
nor U10652 (N_10652,N_10328,N_10140);
nand U10653 (N_10653,N_10095,N_10199);
and U10654 (N_10654,N_10329,N_10020);
nor U10655 (N_10655,N_10270,N_10291);
nor U10656 (N_10656,N_10383,N_10327);
xor U10657 (N_10657,N_10333,N_10085);
nor U10658 (N_10658,N_10373,N_10129);
or U10659 (N_10659,N_10179,N_10421);
nor U10660 (N_10660,N_10063,N_10210);
and U10661 (N_10661,N_10305,N_10091);
nand U10662 (N_10662,N_10415,N_10158);
or U10663 (N_10663,N_10477,N_10420);
nor U10664 (N_10664,N_10437,N_10366);
nand U10665 (N_10665,N_10017,N_10314);
and U10666 (N_10666,N_10038,N_10350);
xnor U10667 (N_10667,N_10155,N_10206);
nor U10668 (N_10668,N_10099,N_10198);
and U10669 (N_10669,N_10346,N_10379);
and U10670 (N_10670,N_10173,N_10150);
nor U10671 (N_10671,N_10339,N_10008);
and U10672 (N_10672,N_10165,N_10480);
nand U10673 (N_10673,N_10493,N_10363);
nand U10674 (N_10674,N_10334,N_10357);
and U10675 (N_10675,N_10461,N_10273);
nor U10676 (N_10676,N_10149,N_10019);
nor U10677 (N_10677,N_10265,N_10133);
and U10678 (N_10678,N_10466,N_10422);
nor U10679 (N_10679,N_10194,N_10176);
nand U10680 (N_10680,N_10268,N_10089);
and U10681 (N_10681,N_10444,N_10232);
and U10682 (N_10682,N_10219,N_10426);
and U10683 (N_10683,N_10053,N_10440);
xnor U10684 (N_10684,N_10144,N_10354);
nor U10685 (N_10685,N_10224,N_10113);
or U10686 (N_10686,N_10000,N_10361);
nand U10687 (N_10687,N_10159,N_10457);
nand U10688 (N_10688,N_10332,N_10316);
and U10689 (N_10689,N_10212,N_10498);
xnor U10690 (N_10690,N_10307,N_10315);
and U10691 (N_10691,N_10300,N_10040);
xnor U10692 (N_10692,N_10277,N_10451);
xor U10693 (N_10693,N_10117,N_10462);
nand U10694 (N_10694,N_10276,N_10134);
nor U10695 (N_10695,N_10251,N_10059);
and U10696 (N_10696,N_10319,N_10171);
or U10697 (N_10697,N_10418,N_10013);
nand U10698 (N_10698,N_10187,N_10064);
and U10699 (N_10699,N_10143,N_10233);
nor U10700 (N_10700,N_10325,N_10065);
and U10701 (N_10701,N_10283,N_10200);
and U10702 (N_10702,N_10079,N_10160);
or U10703 (N_10703,N_10284,N_10263);
and U10704 (N_10704,N_10402,N_10494);
xnor U10705 (N_10705,N_10278,N_10394);
nor U10706 (N_10706,N_10356,N_10456);
nor U10707 (N_10707,N_10320,N_10022);
and U10708 (N_10708,N_10197,N_10393);
and U10709 (N_10709,N_10381,N_10049);
nand U10710 (N_10710,N_10076,N_10338);
nor U10711 (N_10711,N_10491,N_10215);
and U10712 (N_10712,N_10281,N_10028);
and U10713 (N_10713,N_10454,N_10157);
nor U10714 (N_10714,N_10030,N_10188);
or U10715 (N_10715,N_10400,N_10126);
and U10716 (N_10716,N_10371,N_10071);
and U10717 (N_10717,N_10217,N_10335);
xnor U10718 (N_10718,N_10056,N_10476);
or U10719 (N_10719,N_10368,N_10483);
xor U10720 (N_10720,N_10202,N_10039);
or U10721 (N_10721,N_10455,N_10241);
nor U10722 (N_10722,N_10438,N_10012);
nor U10723 (N_10723,N_10010,N_10034);
nor U10724 (N_10724,N_10223,N_10190);
nand U10725 (N_10725,N_10463,N_10084);
and U10726 (N_10726,N_10271,N_10310);
nand U10727 (N_10727,N_10358,N_10047);
nor U10728 (N_10728,N_10414,N_10221);
nand U10729 (N_10729,N_10321,N_10070);
nand U10730 (N_10730,N_10287,N_10131);
or U10731 (N_10731,N_10050,N_10479);
and U10732 (N_10732,N_10262,N_10352);
nand U10733 (N_10733,N_10122,N_10467);
and U10734 (N_10734,N_10392,N_10021);
and U10735 (N_10735,N_10191,N_10406);
nor U10736 (N_10736,N_10343,N_10135);
nor U10737 (N_10737,N_10214,N_10275);
nor U10738 (N_10738,N_10141,N_10458);
and U10739 (N_10739,N_10151,N_10128);
nor U10740 (N_10740,N_10041,N_10387);
nor U10741 (N_10741,N_10424,N_10374);
or U10742 (N_10742,N_10355,N_10449);
or U10743 (N_10743,N_10254,N_10256);
nand U10744 (N_10744,N_10434,N_10236);
xnor U10745 (N_10745,N_10235,N_10370);
or U10746 (N_10746,N_10239,N_10428);
nand U10747 (N_10747,N_10081,N_10044);
nor U10748 (N_10748,N_10404,N_10446);
xor U10749 (N_10749,N_10069,N_10285);
nor U10750 (N_10750,N_10454,N_10434);
nor U10751 (N_10751,N_10400,N_10060);
or U10752 (N_10752,N_10171,N_10333);
and U10753 (N_10753,N_10049,N_10244);
and U10754 (N_10754,N_10418,N_10278);
and U10755 (N_10755,N_10122,N_10199);
xnor U10756 (N_10756,N_10406,N_10281);
xnor U10757 (N_10757,N_10316,N_10037);
nor U10758 (N_10758,N_10013,N_10193);
nor U10759 (N_10759,N_10479,N_10029);
or U10760 (N_10760,N_10419,N_10178);
or U10761 (N_10761,N_10429,N_10107);
or U10762 (N_10762,N_10081,N_10380);
or U10763 (N_10763,N_10285,N_10041);
and U10764 (N_10764,N_10423,N_10067);
nand U10765 (N_10765,N_10485,N_10179);
nor U10766 (N_10766,N_10009,N_10378);
or U10767 (N_10767,N_10368,N_10409);
xor U10768 (N_10768,N_10020,N_10118);
nand U10769 (N_10769,N_10472,N_10295);
and U10770 (N_10770,N_10141,N_10194);
xnor U10771 (N_10771,N_10370,N_10455);
or U10772 (N_10772,N_10486,N_10412);
nand U10773 (N_10773,N_10268,N_10032);
and U10774 (N_10774,N_10273,N_10413);
or U10775 (N_10775,N_10016,N_10216);
xor U10776 (N_10776,N_10245,N_10437);
or U10777 (N_10777,N_10236,N_10383);
nand U10778 (N_10778,N_10318,N_10428);
nor U10779 (N_10779,N_10151,N_10390);
nand U10780 (N_10780,N_10491,N_10307);
xnor U10781 (N_10781,N_10418,N_10094);
xor U10782 (N_10782,N_10483,N_10442);
or U10783 (N_10783,N_10161,N_10095);
or U10784 (N_10784,N_10314,N_10312);
and U10785 (N_10785,N_10345,N_10299);
or U10786 (N_10786,N_10064,N_10456);
xnor U10787 (N_10787,N_10490,N_10317);
nand U10788 (N_10788,N_10056,N_10294);
nand U10789 (N_10789,N_10094,N_10270);
and U10790 (N_10790,N_10384,N_10312);
nand U10791 (N_10791,N_10410,N_10185);
nand U10792 (N_10792,N_10497,N_10371);
or U10793 (N_10793,N_10419,N_10456);
xor U10794 (N_10794,N_10303,N_10118);
nor U10795 (N_10795,N_10478,N_10422);
and U10796 (N_10796,N_10213,N_10067);
or U10797 (N_10797,N_10284,N_10094);
or U10798 (N_10798,N_10027,N_10092);
nand U10799 (N_10799,N_10412,N_10127);
or U10800 (N_10800,N_10499,N_10088);
or U10801 (N_10801,N_10310,N_10355);
xor U10802 (N_10802,N_10067,N_10138);
nor U10803 (N_10803,N_10488,N_10243);
nor U10804 (N_10804,N_10032,N_10128);
nand U10805 (N_10805,N_10499,N_10315);
xor U10806 (N_10806,N_10216,N_10005);
or U10807 (N_10807,N_10088,N_10435);
and U10808 (N_10808,N_10188,N_10089);
nor U10809 (N_10809,N_10227,N_10207);
nand U10810 (N_10810,N_10425,N_10140);
nand U10811 (N_10811,N_10483,N_10303);
or U10812 (N_10812,N_10242,N_10140);
and U10813 (N_10813,N_10118,N_10010);
nor U10814 (N_10814,N_10191,N_10376);
nand U10815 (N_10815,N_10107,N_10351);
xor U10816 (N_10816,N_10486,N_10308);
nor U10817 (N_10817,N_10411,N_10188);
or U10818 (N_10818,N_10395,N_10038);
xor U10819 (N_10819,N_10469,N_10373);
nor U10820 (N_10820,N_10334,N_10201);
or U10821 (N_10821,N_10201,N_10439);
nand U10822 (N_10822,N_10264,N_10052);
xor U10823 (N_10823,N_10369,N_10362);
nor U10824 (N_10824,N_10252,N_10074);
nand U10825 (N_10825,N_10202,N_10265);
xor U10826 (N_10826,N_10092,N_10204);
nand U10827 (N_10827,N_10434,N_10440);
and U10828 (N_10828,N_10374,N_10375);
nor U10829 (N_10829,N_10173,N_10437);
and U10830 (N_10830,N_10179,N_10288);
or U10831 (N_10831,N_10075,N_10182);
and U10832 (N_10832,N_10283,N_10241);
or U10833 (N_10833,N_10355,N_10314);
xor U10834 (N_10834,N_10398,N_10121);
and U10835 (N_10835,N_10421,N_10057);
nor U10836 (N_10836,N_10460,N_10360);
nor U10837 (N_10837,N_10117,N_10380);
xnor U10838 (N_10838,N_10311,N_10135);
xor U10839 (N_10839,N_10381,N_10418);
xor U10840 (N_10840,N_10367,N_10192);
nand U10841 (N_10841,N_10315,N_10327);
nor U10842 (N_10842,N_10219,N_10441);
xor U10843 (N_10843,N_10287,N_10314);
and U10844 (N_10844,N_10123,N_10045);
and U10845 (N_10845,N_10331,N_10376);
xor U10846 (N_10846,N_10065,N_10390);
or U10847 (N_10847,N_10173,N_10460);
and U10848 (N_10848,N_10042,N_10313);
nor U10849 (N_10849,N_10070,N_10368);
nor U10850 (N_10850,N_10352,N_10141);
xnor U10851 (N_10851,N_10198,N_10473);
and U10852 (N_10852,N_10152,N_10018);
nor U10853 (N_10853,N_10206,N_10340);
nor U10854 (N_10854,N_10038,N_10329);
nand U10855 (N_10855,N_10240,N_10158);
nor U10856 (N_10856,N_10151,N_10073);
and U10857 (N_10857,N_10026,N_10016);
nand U10858 (N_10858,N_10203,N_10317);
nand U10859 (N_10859,N_10213,N_10412);
xor U10860 (N_10860,N_10091,N_10419);
nand U10861 (N_10861,N_10398,N_10271);
xnor U10862 (N_10862,N_10399,N_10291);
nor U10863 (N_10863,N_10425,N_10002);
nor U10864 (N_10864,N_10145,N_10167);
or U10865 (N_10865,N_10139,N_10272);
or U10866 (N_10866,N_10370,N_10296);
or U10867 (N_10867,N_10419,N_10475);
nor U10868 (N_10868,N_10035,N_10415);
xor U10869 (N_10869,N_10315,N_10127);
or U10870 (N_10870,N_10281,N_10183);
xor U10871 (N_10871,N_10162,N_10116);
xnor U10872 (N_10872,N_10427,N_10206);
xnor U10873 (N_10873,N_10362,N_10119);
nor U10874 (N_10874,N_10467,N_10293);
nor U10875 (N_10875,N_10192,N_10150);
and U10876 (N_10876,N_10423,N_10058);
nand U10877 (N_10877,N_10169,N_10477);
nand U10878 (N_10878,N_10367,N_10351);
nand U10879 (N_10879,N_10436,N_10172);
or U10880 (N_10880,N_10430,N_10270);
nand U10881 (N_10881,N_10031,N_10187);
nor U10882 (N_10882,N_10392,N_10068);
and U10883 (N_10883,N_10094,N_10476);
or U10884 (N_10884,N_10139,N_10079);
xor U10885 (N_10885,N_10068,N_10293);
or U10886 (N_10886,N_10496,N_10229);
and U10887 (N_10887,N_10402,N_10225);
nor U10888 (N_10888,N_10014,N_10358);
nand U10889 (N_10889,N_10022,N_10251);
xnor U10890 (N_10890,N_10206,N_10381);
and U10891 (N_10891,N_10431,N_10320);
nor U10892 (N_10892,N_10327,N_10158);
and U10893 (N_10893,N_10265,N_10413);
or U10894 (N_10894,N_10214,N_10189);
or U10895 (N_10895,N_10478,N_10187);
or U10896 (N_10896,N_10246,N_10302);
nand U10897 (N_10897,N_10056,N_10038);
xnor U10898 (N_10898,N_10187,N_10355);
and U10899 (N_10899,N_10328,N_10095);
and U10900 (N_10900,N_10041,N_10010);
and U10901 (N_10901,N_10147,N_10205);
nand U10902 (N_10902,N_10388,N_10386);
or U10903 (N_10903,N_10257,N_10031);
or U10904 (N_10904,N_10232,N_10474);
xnor U10905 (N_10905,N_10367,N_10108);
nor U10906 (N_10906,N_10442,N_10282);
and U10907 (N_10907,N_10085,N_10266);
or U10908 (N_10908,N_10196,N_10441);
nor U10909 (N_10909,N_10136,N_10109);
nor U10910 (N_10910,N_10378,N_10011);
and U10911 (N_10911,N_10464,N_10236);
or U10912 (N_10912,N_10170,N_10242);
xor U10913 (N_10913,N_10426,N_10061);
or U10914 (N_10914,N_10074,N_10329);
and U10915 (N_10915,N_10439,N_10031);
xnor U10916 (N_10916,N_10323,N_10270);
and U10917 (N_10917,N_10368,N_10125);
or U10918 (N_10918,N_10361,N_10231);
nand U10919 (N_10919,N_10068,N_10248);
and U10920 (N_10920,N_10135,N_10410);
and U10921 (N_10921,N_10087,N_10398);
xor U10922 (N_10922,N_10054,N_10293);
or U10923 (N_10923,N_10292,N_10367);
and U10924 (N_10924,N_10152,N_10188);
nor U10925 (N_10925,N_10172,N_10077);
xor U10926 (N_10926,N_10346,N_10308);
nor U10927 (N_10927,N_10477,N_10342);
xnor U10928 (N_10928,N_10220,N_10147);
xor U10929 (N_10929,N_10245,N_10119);
nand U10930 (N_10930,N_10121,N_10412);
xor U10931 (N_10931,N_10089,N_10198);
and U10932 (N_10932,N_10318,N_10271);
nand U10933 (N_10933,N_10152,N_10106);
nor U10934 (N_10934,N_10134,N_10497);
or U10935 (N_10935,N_10220,N_10444);
nor U10936 (N_10936,N_10304,N_10056);
nand U10937 (N_10937,N_10323,N_10355);
xnor U10938 (N_10938,N_10484,N_10442);
nor U10939 (N_10939,N_10089,N_10018);
and U10940 (N_10940,N_10311,N_10260);
xnor U10941 (N_10941,N_10397,N_10079);
or U10942 (N_10942,N_10054,N_10133);
or U10943 (N_10943,N_10222,N_10411);
and U10944 (N_10944,N_10179,N_10359);
xor U10945 (N_10945,N_10341,N_10226);
nor U10946 (N_10946,N_10056,N_10420);
nand U10947 (N_10947,N_10448,N_10116);
nand U10948 (N_10948,N_10305,N_10403);
xor U10949 (N_10949,N_10157,N_10287);
and U10950 (N_10950,N_10442,N_10108);
and U10951 (N_10951,N_10205,N_10117);
xor U10952 (N_10952,N_10231,N_10285);
xnor U10953 (N_10953,N_10396,N_10293);
nand U10954 (N_10954,N_10054,N_10083);
and U10955 (N_10955,N_10236,N_10473);
nand U10956 (N_10956,N_10300,N_10270);
xor U10957 (N_10957,N_10322,N_10337);
xnor U10958 (N_10958,N_10031,N_10120);
nand U10959 (N_10959,N_10349,N_10157);
xor U10960 (N_10960,N_10177,N_10365);
xor U10961 (N_10961,N_10118,N_10170);
nand U10962 (N_10962,N_10479,N_10301);
and U10963 (N_10963,N_10372,N_10087);
or U10964 (N_10964,N_10047,N_10148);
nand U10965 (N_10965,N_10192,N_10418);
and U10966 (N_10966,N_10275,N_10391);
and U10967 (N_10967,N_10121,N_10180);
or U10968 (N_10968,N_10292,N_10161);
or U10969 (N_10969,N_10090,N_10394);
nand U10970 (N_10970,N_10113,N_10269);
nor U10971 (N_10971,N_10073,N_10009);
nand U10972 (N_10972,N_10005,N_10178);
xor U10973 (N_10973,N_10465,N_10255);
and U10974 (N_10974,N_10489,N_10205);
nand U10975 (N_10975,N_10414,N_10251);
nand U10976 (N_10976,N_10102,N_10237);
nor U10977 (N_10977,N_10276,N_10260);
or U10978 (N_10978,N_10219,N_10130);
nor U10979 (N_10979,N_10166,N_10375);
and U10980 (N_10980,N_10460,N_10209);
and U10981 (N_10981,N_10206,N_10459);
and U10982 (N_10982,N_10470,N_10384);
xor U10983 (N_10983,N_10096,N_10323);
nor U10984 (N_10984,N_10257,N_10018);
nor U10985 (N_10985,N_10369,N_10406);
nand U10986 (N_10986,N_10137,N_10240);
xnor U10987 (N_10987,N_10360,N_10275);
nand U10988 (N_10988,N_10147,N_10104);
or U10989 (N_10989,N_10142,N_10207);
nand U10990 (N_10990,N_10045,N_10420);
nand U10991 (N_10991,N_10416,N_10117);
nor U10992 (N_10992,N_10061,N_10487);
and U10993 (N_10993,N_10063,N_10389);
or U10994 (N_10994,N_10373,N_10481);
nand U10995 (N_10995,N_10085,N_10141);
xor U10996 (N_10996,N_10415,N_10383);
and U10997 (N_10997,N_10488,N_10233);
and U10998 (N_10998,N_10097,N_10204);
and U10999 (N_10999,N_10138,N_10203);
or U11000 (N_11000,N_10613,N_10631);
or U11001 (N_11001,N_10707,N_10832);
xnor U11002 (N_11002,N_10863,N_10811);
nand U11003 (N_11003,N_10929,N_10992);
xor U11004 (N_11004,N_10847,N_10702);
or U11005 (N_11005,N_10500,N_10727);
and U11006 (N_11006,N_10800,N_10924);
and U11007 (N_11007,N_10955,N_10751);
nand U11008 (N_11008,N_10828,N_10681);
nor U11009 (N_11009,N_10700,N_10773);
xnor U11010 (N_11010,N_10553,N_10522);
nand U11011 (N_11011,N_10972,N_10777);
or U11012 (N_11012,N_10634,N_10752);
or U11013 (N_11013,N_10802,N_10982);
xor U11014 (N_11014,N_10525,N_10557);
nor U11015 (N_11015,N_10670,N_10621);
and U11016 (N_11016,N_10644,N_10560);
xnor U11017 (N_11017,N_10510,N_10834);
nand U11018 (N_11018,N_10555,N_10552);
nor U11019 (N_11019,N_10551,N_10550);
nand U11020 (N_11020,N_10537,N_10583);
xor U11021 (N_11021,N_10960,N_10520);
nor U11022 (N_11022,N_10829,N_10657);
and U11023 (N_11023,N_10755,N_10893);
nand U11024 (N_11024,N_10630,N_10650);
and U11025 (N_11025,N_10734,N_10705);
nor U11026 (N_11026,N_10845,N_10598);
xnor U11027 (N_11027,N_10660,N_10771);
nor U11028 (N_11028,N_10596,N_10742);
and U11029 (N_11029,N_10533,N_10712);
xor U11030 (N_11030,N_10874,N_10656);
or U11031 (N_11031,N_10838,N_10590);
or U11032 (N_11032,N_10808,N_10766);
nor U11033 (N_11033,N_10900,N_10840);
and U11034 (N_11034,N_10781,N_10703);
and U11035 (N_11035,N_10692,N_10579);
nand U11036 (N_11036,N_10722,N_10977);
xnor U11037 (N_11037,N_10693,N_10930);
xor U11038 (N_11038,N_10503,N_10654);
or U11039 (N_11039,N_10882,N_10589);
nor U11040 (N_11040,N_10797,N_10895);
xor U11041 (N_11041,N_10758,N_10878);
and U11042 (N_11042,N_10715,N_10852);
and U11043 (N_11043,N_10810,N_10736);
xor U11044 (N_11044,N_10666,N_10535);
and U11045 (N_11045,N_10603,N_10678);
xnor U11046 (N_11046,N_10515,N_10890);
or U11047 (N_11047,N_10668,N_10954);
nor U11048 (N_11048,N_10606,N_10881);
nor U11049 (N_11049,N_10908,N_10566);
nor U11050 (N_11050,N_10577,N_10661);
nor U11051 (N_11051,N_10764,N_10719);
or U11052 (N_11052,N_10573,N_10540);
nand U11053 (N_11053,N_10897,N_10701);
and U11054 (N_11054,N_10854,N_10993);
nand U11055 (N_11055,N_10633,N_10990);
nor U11056 (N_11056,N_10676,N_10793);
xnor U11057 (N_11057,N_10568,N_10902);
nor U11058 (N_11058,N_10501,N_10912);
nor U11059 (N_11059,N_10718,N_10920);
or U11060 (N_11060,N_10870,N_10695);
or U11061 (N_11061,N_10575,N_10664);
and U11062 (N_11062,N_10985,N_10667);
and U11063 (N_11063,N_10710,N_10507);
or U11064 (N_11064,N_10943,N_10933);
nand U11065 (N_11065,N_10542,N_10697);
nand U11066 (N_11066,N_10625,N_10856);
nand U11067 (N_11067,N_10523,N_10822);
nand U11068 (N_11068,N_10794,N_10949);
nand U11069 (N_11069,N_10947,N_10782);
or U11070 (N_11070,N_10941,N_10818);
xor U11071 (N_11071,N_10658,N_10620);
xnor U11072 (N_11072,N_10546,N_10669);
xor U11073 (N_11073,N_10858,N_10789);
or U11074 (N_11074,N_10763,N_10745);
and U11075 (N_11075,N_10584,N_10823);
or U11076 (N_11076,N_10593,N_10968);
and U11077 (N_11077,N_10820,N_10735);
or U11078 (N_11078,N_10898,N_10617);
nor U11079 (N_11079,N_10975,N_10663);
nand U11080 (N_11080,N_10910,N_10772);
xnor U11081 (N_11081,N_10792,N_10647);
and U11082 (N_11082,N_10964,N_10967);
nor U11083 (N_11083,N_10877,N_10855);
and U11084 (N_11084,N_10601,N_10865);
xor U11085 (N_11085,N_10738,N_10916);
or U11086 (N_11086,N_10925,N_10754);
xor U11087 (N_11087,N_10588,N_10850);
xnor U11088 (N_11088,N_10641,N_10795);
nand U11089 (N_11089,N_10514,N_10830);
nand U11090 (N_11090,N_10979,N_10944);
and U11091 (N_11091,N_10974,N_10932);
nand U11092 (N_11092,N_10645,N_10775);
nor U11093 (N_11093,N_10605,N_10909);
or U11094 (N_11094,N_10814,N_10713);
xor U11095 (N_11095,N_10765,N_10779);
and U11096 (N_11096,N_10659,N_10996);
or U11097 (N_11097,N_10788,N_10649);
nor U11098 (N_11098,N_10615,N_10917);
xnor U11099 (N_11099,N_10841,N_10937);
and U11100 (N_11100,N_10831,N_10687);
nor U11101 (N_11101,N_10871,N_10739);
nor U11102 (N_11102,N_10971,N_10757);
nand U11103 (N_11103,N_10688,N_10939);
or U11104 (N_11104,N_10652,N_10685);
and U11105 (N_11105,N_10572,N_10873);
and U11106 (N_11106,N_10699,N_10511);
nand U11107 (N_11107,N_10776,N_10635);
nor U11108 (N_11108,N_10582,N_10839);
or U11109 (N_11109,N_10686,N_10906);
xnor U11110 (N_11110,N_10524,N_10885);
and U11111 (N_11111,N_10821,N_10867);
and U11112 (N_11112,N_10962,N_10804);
xnor U11113 (N_11113,N_10945,N_10998);
nand U11114 (N_11114,N_10724,N_10516);
nor U11115 (N_11115,N_10767,N_10696);
or U11116 (N_11116,N_10622,N_10760);
xnor U11117 (N_11117,N_10959,N_10869);
and U11118 (N_11118,N_10716,N_10543);
nor U11119 (N_11119,N_10581,N_10903);
and U11120 (N_11120,N_10899,N_10623);
nor U11121 (N_11121,N_10927,N_10809);
nor U11122 (N_11122,N_10883,N_10534);
nand U11123 (N_11123,N_10539,N_10892);
xor U11124 (N_11124,N_10733,N_10536);
nand U11125 (N_11125,N_10558,N_10774);
nor U11126 (N_11126,N_10571,N_10853);
and U11127 (N_11127,N_10879,N_10729);
and U11128 (N_11128,N_10966,N_10901);
and U11129 (N_11129,N_10561,N_10548);
nand U11130 (N_11130,N_10642,N_10679);
and U11131 (N_11131,N_10691,N_10973);
xor U11132 (N_11132,N_10704,N_10835);
and U11133 (N_11133,N_10612,N_10628);
and U11134 (N_11134,N_10837,N_10690);
nor U11135 (N_11135,N_10915,N_10559);
xnor U11136 (N_11136,N_10565,N_10787);
and U11137 (N_11137,N_10848,N_10948);
nor U11138 (N_11138,N_10585,N_10896);
and U11139 (N_11139,N_10940,N_10639);
or U11140 (N_11140,N_10721,N_10849);
and U11141 (N_11141,N_10769,N_10725);
xnor U11142 (N_11142,N_10988,N_10714);
nor U11143 (N_11143,N_10815,N_10907);
and U11144 (N_11144,N_10604,N_10609);
and U11145 (N_11145,N_10783,N_10616);
and U11146 (N_11146,N_10860,N_10756);
nor U11147 (N_11147,N_10567,N_10816);
or U11148 (N_11148,N_10506,N_10935);
nand U11149 (N_11149,N_10651,N_10862);
xnor U11150 (N_11150,N_10570,N_10994);
xor U11151 (N_11151,N_10737,N_10806);
nand U11152 (N_11152,N_10951,N_10614);
nor U11153 (N_11153,N_10646,N_10961);
nand U11154 (N_11154,N_10619,N_10526);
nand U11155 (N_11155,N_10600,N_10938);
nand U11156 (N_11156,N_10711,N_10889);
nand U11157 (N_11157,N_10905,N_10698);
or U11158 (N_11158,N_10842,N_10790);
nand U11159 (N_11159,N_10513,N_10741);
and U11160 (N_11160,N_10564,N_10866);
nand U11161 (N_11161,N_10872,N_10743);
or U11162 (N_11162,N_10762,N_10984);
and U11163 (N_11163,N_10965,N_10638);
nor U11164 (N_11164,N_10934,N_10827);
and U11165 (N_11165,N_10529,N_10655);
nand U11166 (N_11166,N_10544,N_10978);
nor U11167 (N_11167,N_10851,N_10904);
and U11168 (N_11168,N_10740,N_10509);
and U11169 (N_11169,N_10749,N_10610);
nor U11170 (N_11170,N_10956,N_10894);
and U11171 (N_11171,N_10844,N_10530);
or U11172 (N_11172,N_10708,N_10611);
nor U11173 (N_11173,N_10886,N_10674);
and U11174 (N_11174,N_10958,N_10914);
nor U11175 (N_11175,N_10911,N_10928);
xnor U11176 (N_11176,N_10723,N_10980);
or U11177 (N_11177,N_10648,N_10784);
nor U11178 (N_11178,N_10876,N_10868);
nand U11179 (N_11179,N_10887,N_10683);
or U11180 (N_11180,N_10950,N_10813);
nand U11181 (N_11181,N_10921,N_10595);
or U11182 (N_11182,N_10919,N_10549);
and U11183 (N_11183,N_10786,N_10987);
nand U11184 (N_11184,N_10983,N_10618);
or U11185 (N_11185,N_10976,N_10836);
nor U11186 (N_11186,N_10521,N_10969);
nor U11187 (N_11187,N_10778,N_10799);
and U11188 (N_11188,N_10770,N_10519);
xnor U11189 (N_11189,N_10750,N_10833);
and U11190 (N_11190,N_10594,N_10576);
nor U11191 (N_11191,N_10953,N_10592);
and U11192 (N_11192,N_10512,N_10671);
or U11193 (N_11193,N_10597,N_10759);
xor U11194 (N_11194,N_10824,N_10846);
nor U11195 (N_11195,N_10732,N_10677);
or U11196 (N_11196,N_10508,N_10607);
and U11197 (N_11197,N_10785,N_10817);
xnor U11198 (N_11198,N_10665,N_10826);
nor U11199 (N_11199,N_10747,N_10636);
and U11200 (N_11200,N_10569,N_10918);
xnor U11201 (N_11201,N_10626,N_10689);
nand U11202 (N_11202,N_10819,N_10629);
or U11203 (N_11203,N_10528,N_10580);
and U11204 (N_11204,N_10502,N_10706);
nand U11205 (N_11205,N_10922,N_10527);
nor U11206 (N_11206,N_10717,N_10643);
nand U11207 (N_11207,N_10554,N_10875);
xor U11208 (N_11208,N_10673,N_10518);
and U11209 (N_11209,N_10672,N_10591);
nor U11210 (N_11210,N_10861,N_10926);
and U11211 (N_11211,N_10562,N_10627);
xnor U11212 (N_11212,N_10709,N_10768);
xor U11213 (N_11213,N_10728,N_10680);
or U11214 (N_11214,N_10505,N_10517);
nor U11215 (N_11215,N_10744,N_10963);
nor U11216 (N_11216,N_10888,N_10946);
and U11217 (N_11217,N_10857,N_10602);
and U11218 (N_11218,N_10803,N_10545);
xor U11219 (N_11219,N_10730,N_10624);
or U11220 (N_11220,N_10748,N_10913);
nor U11221 (N_11221,N_10942,N_10504);
nand U11222 (N_11222,N_10931,N_10952);
nand U11223 (N_11223,N_10989,N_10599);
and U11224 (N_11224,N_10694,N_10957);
nand U11225 (N_11225,N_10981,N_10586);
and U11226 (N_11226,N_10807,N_10997);
nor U11227 (N_11227,N_10801,N_10991);
nand U11228 (N_11228,N_10798,N_10936);
nand U11229 (N_11229,N_10556,N_10812);
nand U11230 (N_11230,N_10753,N_10578);
or U11231 (N_11231,N_10970,N_10531);
xor U11232 (N_11232,N_10761,N_10682);
or U11233 (N_11233,N_10780,N_10796);
xnor U11234 (N_11234,N_10843,N_10640);
nor U11235 (N_11235,N_10805,N_10662);
nor U11236 (N_11236,N_10541,N_10532);
or U11237 (N_11237,N_10986,N_10684);
nand U11238 (N_11238,N_10538,N_10864);
nor U11239 (N_11239,N_10563,N_10880);
nor U11240 (N_11240,N_10547,N_10653);
nor U11241 (N_11241,N_10746,N_10608);
xnor U11242 (N_11242,N_10632,N_10859);
or U11243 (N_11243,N_10923,N_10720);
xor U11244 (N_11244,N_10731,N_10999);
nand U11245 (N_11245,N_10675,N_10574);
or U11246 (N_11246,N_10587,N_10726);
or U11247 (N_11247,N_10791,N_10995);
or U11248 (N_11248,N_10884,N_10825);
nand U11249 (N_11249,N_10891,N_10637);
nand U11250 (N_11250,N_10803,N_10630);
nor U11251 (N_11251,N_10972,N_10652);
or U11252 (N_11252,N_10906,N_10612);
nand U11253 (N_11253,N_10901,N_10786);
nor U11254 (N_11254,N_10760,N_10660);
or U11255 (N_11255,N_10883,N_10526);
xnor U11256 (N_11256,N_10686,N_10729);
xnor U11257 (N_11257,N_10863,N_10542);
nand U11258 (N_11258,N_10652,N_10665);
nand U11259 (N_11259,N_10651,N_10604);
nor U11260 (N_11260,N_10631,N_10623);
nor U11261 (N_11261,N_10998,N_10986);
and U11262 (N_11262,N_10828,N_10955);
nand U11263 (N_11263,N_10803,N_10897);
and U11264 (N_11264,N_10975,N_10792);
and U11265 (N_11265,N_10670,N_10972);
or U11266 (N_11266,N_10972,N_10981);
xnor U11267 (N_11267,N_10640,N_10575);
and U11268 (N_11268,N_10674,N_10681);
and U11269 (N_11269,N_10892,N_10831);
nand U11270 (N_11270,N_10906,N_10564);
or U11271 (N_11271,N_10691,N_10730);
nand U11272 (N_11272,N_10933,N_10681);
nor U11273 (N_11273,N_10793,N_10938);
and U11274 (N_11274,N_10837,N_10872);
nor U11275 (N_11275,N_10815,N_10677);
or U11276 (N_11276,N_10953,N_10967);
xnor U11277 (N_11277,N_10635,N_10712);
or U11278 (N_11278,N_10789,N_10737);
or U11279 (N_11279,N_10994,N_10531);
and U11280 (N_11280,N_10882,N_10540);
nand U11281 (N_11281,N_10749,N_10870);
and U11282 (N_11282,N_10845,N_10631);
nor U11283 (N_11283,N_10703,N_10889);
or U11284 (N_11284,N_10916,N_10754);
nor U11285 (N_11285,N_10544,N_10849);
xor U11286 (N_11286,N_10922,N_10537);
xor U11287 (N_11287,N_10616,N_10765);
nand U11288 (N_11288,N_10626,N_10680);
nor U11289 (N_11289,N_10502,N_10730);
and U11290 (N_11290,N_10851,N_10560);
and U11291 (N_11291,N_10798,N_10861);
nand U11292 (N_11292,N_10991,N_10516);
nand U11293 (N_11293,N_10904,N_10650);
or U11294 (N_11294,N_10626,N_10757);
and U11295 (N_11295,N_10586,N_10922);
and U11296 (N_11296,N_10959,N_10742);
nor U11297 (N_11297,N_10563,N_10760);
xnor U11298 (N_11298,N_10846,N_10537);
nand U11299 (N_11299,N_10972,N_10802);
or U11300 (N_11300,N_10529,N_10745);
nor U11301 (N_11301,N_10950,N_10850);
xor U11302 (N_11302,N_10864,N_10559);
nand U11303 (N_11303,N_10786,N_10742);
nand U11304 (N_11304,N_10588,N_10513);
nor U11305 (N_11305,N_10621,N_10958);
nor U11306 (N_11306,N_10760,N_10520);
nand U11307 (N_11307,N_10932,N_10898);
and U11308 (N_11308,N_10728,N_10633);
nor U11309 (N_11309,N_10778,N_10800);
nand U11310 (N_11310,N_10862,N_10506);
nor U11311 (N_11311,N_10888,N_10940);
nand U11312 (N_11312,N_10678,N_10909);
xnor U11313 (N_11313,N_10801,N_10550);
and U11314 (N_11314,N_10620,N_10728);
nand U11315 (N_11315,N_10777,N_10928);
nor U11316 (N_11316,N_10727,N_10718);
and U11317 (N_11317,N_10834,N_10618);
nand U11318 (N_11318,N_10565,N_10640);
nand U11319 (N_11319,N_10846,N_10692);
nand U11320 (N_11320,N_10721,N_10916);
xnor U11321 (N_11321,N_10671,N_10517);
and U11322 (N_11322,N_10667,N_10997);
nor U11323 (N_11323,N_10847,N_10972);
nor U11324 (N_11324,N_10949,N_10554);
or U11325 (N_11325,N_10694,N_10655);
nor U11326 (N_11326,N_10526,N_10817);
and U11327 (N_11327,N_10880,N_10555);
and U11328 (N_11328,N_10739,N_10901);
or U11329 (N_11329,N_10902,N_10813);
and U11330 (N_11330,N_10825,N_10722);
and U11331 (N_11331,N_10739,N_10830);
xnor U11332 (N_11332,N_10950,N_10508);
xor U11333 (N_11333,N_10579,N_10546);
or U11334 (N_11334,N_10718,N_10935);
nand U11335 (N_11335,N_10797,N_10639);
and U11336 (N_11336,N_10979,N_10738);
or U11337 (N_11337,N_10901,N_10893);
and U11338 (N_11338,N_10541,N_10512);
nand U11339 (N_11339,N_10755,N_10838);
nor U11340 (N_11340,N_10986,N_10508);
nor U11341 (N_11341,N_10661,N_10808);
nand U11342 (N_11342,N_10513,N_10693);
and U11343 (N_11343,N_10548,N_10801);
and U11344 (N_11344,N_10503,N_10799);
and U11345 (N_11345,N_10713,N_10828);
and U11346 (N_11346,N_10946,N_10940);
xnor U11347 (N_11347,N_10919,N_10844);
xor U11348 (N_11348,N_10762,N_10929);
and U11349 (N_11349,N_10724,N_10920);
nor U11350 (N_11350,N_10770,N_10628);
xor U11351 (N_11351,N_10531,N_10791);
nand U11352 (N_11352,N_10918,N_10772);
or U11353 (N_11353,N_10540,N_10621);
xor U11354 (N_11354,N_10734,N_10836);
or U11355 (N_11355,N_10887,N_10726);
or U11356 (N_11356,N_10796,N_10992);
and U11357 (N_11357,N_10774,N_10733);
and U11358 (N_11358,N_10788,N_10567);
or U11359 (N_11359,N_10775,N_10686);
nor U11360 (N_11360,N_10593,N_10642);
nor U11361 (N_11361,N_10912,N_10980);
nor U11362 (N_11362,N_10722,N_10983);
or U11363 (N_11363,N_10729,N_10904);
xor U11364 (N_11364,N_10670,N_10649);
and U11365 (N_11365,N_10853,N_10871);
or U11366 (N_11366,N_10502,N_10766);
nor U11367 (N_11367,N_10747,N_10864);
or U11368 (N_11368,N_10912,N_10667);
or U11369 (N_11369,N_10830,N_10696);
nor U11370 (N_11370,N_10510,N_10755);
nand U11371 (N_11371,N_10958,N_10818);
or U11372 (N_11372,N_10667,N_10918);
xor U11373 (N_11373,N_10689,N_10882);
nor U11374 (N_11374,N_10609,N_10904);
nor U11375 (N_11375,N_10828,N_10701);
xnor U11376 (N_11376,N_10887,N_10532);
nor U11377 (N_11377,N_10921,N_10703);
xnor U11378 (N_11378,N_10981,N_10706);
nor U11379 (N_11379,N_10509,N_10685);
nand U11380 (N_11380,N_10904,N_10726);
and U11381 (N_11381,N_10504,N_10685);
and U11382 (N_11382,N_10557,N_10874);
nand U11383 (N_11383,N_10586,N_10543);
xor U11384 (N_11384,N_10500,N_10983);
or U11385 (N_11385,N_10920,N_10884);
nor U11386 (N_11386,N_10685,N_10687);
and U11387 (N_11387,N_10761,N_10624);
nor U11388 (N_11388,N_10571,N_10521);
nand U11389 (N_11389,N_10984,N_10834);
or U11390 (N_11390,N_10690,N_10518);
nor U11391 (N_11391,N_10657,N_10963);
nor U11392 (N_11392,N_10925,N_10842);
xnor U11393 (N_11393,N_10735,N_10598);
nor U11394 (N_11394,N_10933,N_10999);
nand U11395 (N_11395,N_10702,N_10539);
and U11396 (N_11396,N_10737,N_10982);
nand U11397 (N_11397,N_10763,N_10753);
nand U11398 (N_11398,N_10643,N_10612);
nand U11399 (N_11399,N_10787,N_10764);
or U11400 (N_11400,N_10728,N_10936);
or U11401 (N_11401,N_10789,N_10702);
nand U11402 (N_11402,N_10532,N_10827);
nor U11403 (N_11403,N_10988,N_10504);
nand U11404 (N_11404,N_10714,N_10797);
xnor U11405 (N_11405,N_10931,N_10627);
nor U11406 (N_11406,N_10749,N_10821);
xor U11407 (N_11407,N_10908,N_10787);
nor U11408 (N_11408,N_10557,N_10776);
or U11409 (N_11409,N_10534,N_10750);
and U11410 (N_11410,N_10813,N_10688);
nor U11411 (N_11411,N_10812,N_10972);
nor U11412 (N_11412,N_10821,N_10933);
or U11413 (N_11413,N_10573,N_10666);
nand U11414 (N_11414,N_10795,N_10734);
nor U11415 (N_11415,N_10888,N_10957);
nor U11416 (N_11416,N_10687,N_10765);
nor U11417 (N_11417,N_10744,N_10966);
nor U11418 (N_11418,N_10504,N_10587);
or U11419 (N_11419,N_10946,N_10831);
or U11420 (N_11420,N_10855,N_10665);
and U11421 (N_11421,N_10873,N_10725);
nand U11422 (N_11422,N_10893,N_10859);
or U11423 (N_11423,N_10931,N_10675);
or U11424 (N_11424,N_10687,N_10645);
or U11425 (N_11425,N_10563,N_10551);
or U11426 (N_11426,N_10682,N_10566);
or U11427 (N_11427,N_10572,N_10840);
and U11428 (N_11428,N_10634,N_10869);
nor U11429 (N_11429,N_10880,N_10539);
or U11430 (N_11430,N_10789,N_10621);
nand U11431 (N_11431,N_10627,N_10519);
and U11432 (N_11432,N_10554,N_10784);
nor U11433 (N_11433,N_10622,N_10682);
and U11434 (N_11434,N_10600,N_10674);
xnor U11435 (N_11435,N_10510,N_10718);
nand U11436 (N_11436,N_10610,N_10732);
nor U11437 (N_11437,N_10554,N_10776);
nor U11438 (N_11438,N_10782,N_10892);
or U11439 (N_11439,N_10732,N_10830);
nor U11440 (N_11440,N_10873,N_10539);
and U11441 (N_11441,N_10852,N_10720);
nand U11442 (N_11442,N_10901,N_10804);
xnor U11443 (N_11443,N_10528,N_10805);
nand U11444 (N_11444,N_10965,N_10885);
xor U11445 (N_11445,N_10665,N_10891);
xnor U11446 (N_11446,N_10615,N_10856);
or U11447 (N_11447,N_10660,N_10986);
and U11448 (N_11448,N_10718,N_10612);
nand U11449 (N_11449,N_10738,N_10545);
and U11450 (N_11450,N_10956,N_10995);
or U11451 (N_11451,N_10679,N_10762);
nor U11452 (N_11452,N_10836,N_10921);
and U11453 (N_11453,N_10501,N_10814);
xnor U11454 (N_11454,N_10694,N_10921);
nand U11455 (N_11455,N_10734,N_10851);
nor U11456 (N_11456,N_10617,N_10894);
nor U11457 (N_11457,N_10762,N_10864);
xor U11458 (N_11458,N_10581,N_10695);
and U11459 (N_11459,N_10974,N_10855);
nand U11460 (N_11460,N_10648,N_10623);
xor U11461 (N_11461,N_10776,N_10654);
and U11462 (N_11462,N_10962,N_10771);
and U11463 (N_11463,N_10778,N_10586);
nor U11464 (N_11464,N_10790,N_10882);
nand U11465 (N_11465,N_10608,N_10974);
nand U11466 (N_11466,N_10996,N_10843);
nor U11467 (N_11467,N_10886,N_10809);
xor U11468 (N_11468,N_10626,N_10911);
or U11469 (N_11469,N_10554,N_10790);
and U11470 (N_11470,N_10725,N_10956);
xor U11471 (N_11471,N_10748,N_10765);
xor U11472 (N_11472,N_10734,N_10579);
nor U11473 (N_11473,N_10995,N_10934);
nand U11474 (N_11474,N_10711,N_10835);
nand U11475 (N_11475,N_10677,N_10702);
nor U11476 (N_11476,N_10727,N_10768);
xnor U11477 (N_11477,N_10682,N_10999);
and U11478 (N_11478,N_10951,N_10743);
nand U11479 (N_11479,N_10871,N_10626);
and U11480 (N_11480,N_10968,N_10956);
and U11481 (N_11481,N_10502,N_10782);
xnor U11482 (N_11482,N_10945,N_10737);
or U11483 (N_11483,N_10640,N_10899);
xnor U11484 (N_11484,N_10630,N_10749);
xnor U11485 (N_11485,N_10580,N_10819);
xnor U11486 (N_11486,N_10684,N_10530);
xor U11487 (N_11487,N_10992,N_10993);
nand U11488 (N_11488,N_10552,N_10835);
nor U11489 (N_11489,N_10945,N_10722);
nand U11490 (N_11490,N_10859,N_10880);
xnor U11491 (N_11491,N_10670,N_10603);
nor U11492 (N_11492,N_10779,N_10839);
and U11493 (N_11493,N_10866,N_10787);
and U11494 (N_11494,N_10580,N_10988);
and U11495 (N_11495,N_10544,N_10952);
and U11496 (N_11496,N_10885,N_10818);
or U11497 (N_11497,N_10675,N_10695);
and U11498 (N_11498,N_10524,N_10786);
nand U11499 (N_11499,N_10748,N_10744);
nor U11500 (N_11500,N_11297,N_11330);
or U11501 (N_11501,N_11464,N_11028);
and U11502 (N_11502,N_11125,N_11012);
or U11503 (N_11503,N_11335,N_11339);
xor U11504 (N_11504,N_11134,N_11313);
nor U11505 (N_11505,N_11244,N_11346);
xor U11506 (N_11506,N_11331,N_11496);
and U11507 (N_11507,N_11337,N_11165);
xor U11508 (N_11508,N_11401,N_11392);
and U11509 (N_11509,N_11135,N_11215);
xnor U11510 (N_11510,N_11426,N_11262);
or U11511 (N_11511,N_11365,N_11196);
xor U11512 (N_11512,N_11322,N_11203);
xnor U11513 (N_11513,N_11433,N_11066);
xnor U11514 (N_11514,N_11311,N_11382);
xnor U11515 (N_11515,N_11372,N_11105);
or U11516 (N_11516,N_11047,N_11438);
or U11517 (N_11517,N_11217,N_11497);
nor U11518 (N_11518,N_11082,N_11178);
xnor U11519 (N_11519,N_11170,N_11027);
and U11520 (N_11520,N_11257,N_11294);
and U11521 (N_11521,N_11317,N_11273);
nor U11522 (N_11522,N_11298,N_11256);
nor U11523 (N_11523,N_11046,N_11344);
xor U11524 (N_11524,N_11149,N_11428);
xnor U11525 (N_11525,N_11449,N_11320);
nand U11526 (N_11526,N_11448,N_11143);
or U11527 (N_11527,N_11173,N_11126);
nand U11528 (N_11528,N_11148,N_11390);
and U11529 (N_11529,N_11356,N_11423);
or U11530 (N_11530,N_11160,N_11247);
or U11531 (N_11531,N_11106,N_11415);
and U11532 (N_11532,N_11179,N_11471);
nor U11533 (N_11533,N_11068,N_11245);
nand U11534 (N_11534,N_11169,N_11272);
or U11535 (N_11535,N_11358,N_11013);
xor U11536 (N_11536,N_11296,N_11034);
nor U11537 (N_11537,N_11109,N_11067);
and U11538 (N_11538,N_11050,N_11209);
and U11539 (N_11539,N_11024,N_11376);
or U11540 (N_11540,N_11118,N_11277);
xnor U11541 (N_11541,N_11220,N_11212);
or U11542 (N_11542,N_11491,N_11015);
and U11543 (N_11543,N_11480,N_11379);
nor U11544 (N_11544,N_11299,N_11091);
nor U11545 (N_11545,N_11072,N_11281);
nor U11546 (N_11546,N_11111,N_11351);
nor U11547 (N_11547,N_11269,N_11253);
or U11548 (N_11548,N_11435,N_11210);
nor U11549 (N_11549,N_11267,N_11248);
xor U11550 (N_11550,N_11176,N_11123);
and U11551 (N_11551,N_11167,N_11040);
and U11552 (N_11552,N_11338,N_11218);
xnor U11553 (N_11553,N_11285,N_11062);
xor U11554 (N_11554,N_11033,N_11293);
xor U11555 (N_11555,N_11226,N_11292);
or U11556 (N_11556,N_11171,N_11432);
nor U11557 (N_11557,N_11429,N_11185);
nand U11558 (N_11558,N_11343,N_11271);
xnor U11559 (N_11559,N_11348,N_11147);
nand U11560 (N_11560,N_11200,N_11043);
and U11561 (N_11561,N_11159,N_11307);
xnor U11562 (N_11562,N_11407,N_11085);
or U11563 (N_11563,N_11460,N_11194);
and U11564 (N_11564,N_11304,N_11058);
xor U11565 (N_11565,N_11439,N_11396);
and U11566 (N_11566,N_11265,N_11350);
nor U11567 (N_11567,N_11150,N_11009);
nand U11568 (N_11568,N_11347,N_11456);
or U11569 (N_11569,N_11475,N_11057);
xor U11570 (N_11570,N_11008,N_11342);
nor U11571 (N_11571,N_11071,N_11386);
and U11572 (N_11572,N_11395,N_11295);
xnor U11573 (N_11573,N_11375,N_11142);
nor U11574 (N_11574,N_11486,N_11286);
nand U11575 (N_11575,N_11039,N_11184);
nand U11576 (N_11576,N_11181,N_11090);
or U11577 (N_11577,N_11198,N_11060);
nor U11578 (N_11578,N_11369,N_11122);
or U11579 (N_11579,N_11233,N_11325);
nand U11580 (N_11580,N_11484,N_11107);
nand U11581 (N_11581,N_11055,N_11195);
nand U11582 (N_11582,N_11202,N_11110);
nor U11583 (N_11583,N_11468,N_11373);
xnor U11584 (N_11584,N_11444,N_11461);
nor U11585 (N_11585,N_11450,N_11153);
nor U11586 (N_11586,N_11139,N_11476);
or U11587 (N_11587,N_11264,N_11467);
or U11588 (N_11588,N_11228,N_11070);
or U11589 (N_11589,N_11000,N_11494);
xor U11590 (N_11590,N_11029,N_11145);
and U11591 (N_11591,N_11154,N_11499);
nor U11592 (N_11592,N_11458,N_11457);
and U11593 (N_11593,N_11427,N_11364);
and U11594 (N_11594,N_11214,N_11132);
xor U11595 (N_11595,N_11182,N_11394);
or U11596 (N_11596,N_11414,N_11199);
or U11597 (N_11597,N_11026,N_11133);
xor U11598 (N_11598,N_11278,N_11225);
xnor U11599 (N_11599,N_11341,N_11319);
nand U11600 (N_11600,N_11451,N_11190);
or U11601 (N_11601,N_11310,N_11096);
xnor U11602 (N_11602,N_11422,N_11436);
or U11603 (N_11603,N_11406,N_11137);
nand U11604 (N_11604,N_11124,N_11121);
and U11605 (N_11605,N_11250,N_11288);
or U11606 (N_11606,N_11321,N_11352);
or U11607 (N_11607,N_11227,N_11175);
nor U11608 (N_11608,N_11318,N_11400);
and U11609 (N_11609,N_11483,N_11038);
nor U11610 (N_11610,N_11465,N_11023);
nor U11611 (N_11611,N_11128,N_11187);
or U11612 (N_11612,N_11254,N_11037);
and U11613 (N_11613,N_11355,N_11088);
nand U11614 (N_11614,N_11064,N_11136);
nand U11615 (N_11615,N_11489,N_11002);
nand U11616 (N_11616,N_11092,N_11409);
or U11617 (N_11617,N_11157,N_11316);
nor U11618 (N_11618,N_11001,N_11353);
nand U11619 (N_11619,N_11418,N_11324);
and U11620 (N_11620,N_11059,N_11018);
and U11621 (N_11621,N_11016,N_11385);
nand U11622 (N_11622,N_11381,N_11208);
or U11623 (N_11623,N_11243,N_11114);
xor U11624 (N_11624,N_11455,N_11201);
nand U11625 (N_11625,N_11222,N_11367);
nor U11626 (N_11626,N_11030,N_11240);
nand U11627 (N_11627,N_11302,N_11162);
nor U11628 (N_11628,N_11417,N_11261);
xnor U11629 (N_11629,N_11477,N_11259);
and U11630 (N_11630,N_11100,N_11025);
or U11631 (N_11631,N_11260,N_11393);
nand U11632 (N_11632,N_11340,N_11473);
nor U11633 (N_11633,N_11357,N_11099);
and U11634 (N_11634,N_11279,N_11239);
or U11635 (N_11635,N_11230,N_11014);
xor U11636 (N_11636,N_11236,N_11021);
nand U11637 (N_11637,N_11301,N_11005);
and U11638 (N_11638,N_11087,N_11127);
nand U11639 (N_11639,N_11078,N_11398);
xor U11640 (N_11640,N_11183,N_11174);
or U11641 (N_11641,N_11280,N_11421);
nor U11642 (N_11642,N_11152,N_11470);
and U11643 (N_11643,N_11097,N_11413);
nand U11644 (N_11644,N_11361,N_11481);
or U11645 (N_11645,N_11130,N_11052);
and U11646 (N_11646,N_11479,N_11300);
nand U11647 (N_11647,N_11388,N_11075);
nand U11648 (N_11648,N_11430,N_11424);
nor U11649 (N_11649,N_11419,N_11258);
nor U11650 (N_11650,N_11094,N_11079);
and U11651 (N_11651,N_11263,N_11158);
or U11652 (N_11652,N_11336,N_11354);
nor U11653 (N_11653,N_11086,N_11129);
and U11654 (N_11654,N_11490,N_11384);
or U11655 (N_11655,N_11076,N_11303);
and U11656 (N_11656,N_11144,N_11207);
nor U11657 (N_11657,N_11411,N_11268);
nor U11658 (N_11658,N_11309,N_11054);
xnor U11659 (N_11659,N_11363,N_11266);
or U11660 (N_11660,N_11161,N_11425);
nor U11661 (N_11661,N_11290,N_11443);
nand U11662 (N_11662,N_11377,N_11042);
or U11663 (N_11663,N_11420,N_11334);
xnor U11664 (N_11664,N_11482,N_11234);
and U11665 (N_11665,N_11332,N_11103);
or U11666 (N_11666,N_11083,N_11387);
xnor U11667 (N_11667,N_11229,N_11431);
nor U11668 (N_11668,N_11498,N_11305);
or U11669 (N_11669,N_11360,N_11485);
and U11670 (N_11670,N_11323,N_11437);
xor U11671 (N_11671,N_11252,N_11463);
xor U11672 (N_11672,N_11069,N_11020);
xnor U11673 (N_11673,N_11368,N_11146);
nand U11674 (N_11674,N_11495,N_11093);
nor U11675 (N_11675,N_11061,N_11188);
nor U11676 (N_11676,N_11180,N_11131);
nor U11677 (N_11677,N_11073,N_11041);
or U11678 (N_11678,N_11410,N_11232);
or U11679 (N_11679,N_11216,N_11077);
nor U11680 (N_11680,N_11312,N_11004);
nand U11681 (N_11681,N_11080,N_11459);
xor U11682 (N_11682,N_11466,N_11276);
or U11683 (N_11683,N_11151,N_11095);
and U11684 (N_11684,N_11446,N_11397);
nor U11685 (N_11685,N_11287,N_11156);
and U11686 (N_11686,N_11275,N_11308);
nand U11687 (N_11687,N_11333,N_11035);
nand U11688 (N_11688,N_11447,N_11140);
nor U11689 (N_11689,N_11172,N_11006);
xnor U11690 (N_11690,N_11440,N_11063);
xnor U11691 (N_11691,N_11102,N_11168);
nor U11692 (N_11692,N_11474,N_11166);
xor U11693 (N_11693,N_11488,N_11327);
xnor U11694 (N_11694,N_11402,N_11326);
xor U11695 (N_11695,N_11469,N_11044);
nor U11696 (N_11696,N_11383,N_11119);
and U11697 (N_11697,N_11003,N_11138);
xor U11698 (N_11698,N_11283,N_11163);
nor U11699 (N_11699,N_11362,N_11370);
nand U11700 (N_11700,N_11115,N_11051);
nor U11701 (N_11701,N_11315,N_11291);
nor U11702 (N_11702,N_11306,N_11206);
nor U11703 (N_11703,N_11434,N_11492);
xor U11704 (N_11704,N_11022,N_11270);
and U11705 (N_11705,N_11445,N_11186);
and U11706 (N_11706,N_11045,N_11011);
nor U11707 (N_11707,N_11412,N_11191);
and U11708 (N_11708,N_11274,N_11284);
or U11709 (N_11709,N_11017,N_11231);
or U11710 (N_11710,N_11141,N_11189);
xor U11711 (N_11711,N_11249,N_11242);
nand U11712 (N_11712,N_11112,N_11241);
or U11713 (N_11713,N_11053,N_11329);
nand U11714 (N_11714,N_11224,N_11098);
or U11715 (N_11715,N_11223,N_11031);
xor U11716 (N_11716,N_11391,N_11197);
nand U11717 (N_11717,N_11049,N_11113);
and U11718 (N_11718,N_11048,N_11032);
and U11719 (N_11719,N_11116,N_11378);
or U11720 (N_11720,N_11416,N_11453);
nor U11721 (N_11721,N_11193,N_11246);
and U11722 (N_11722,N_11380,N_11487);
xnor U11723 (N_11723,N_11371,N_11235);
and U11724 (N_11724,N_11036,N_11404);
xor U11725 (N_11725,N_11019,N_11205);
xnor U11726 (N_11726,N_11462,N_11211);
xor U11727 (N_11727,N_11084,N_11101);
and U11728 (N_11728,N_11255,N_11056);
xnor U11729 (N_11729,N_11408,N_11289);
nor U11730 (N_11730,N_11221,N_11007);
or U11731 (N_11731,N_11164,N_11010);
or U11732 (N_11732,N_11441,N_11345);
xor U11733 (N_11733,N_11081,N_11374);
xnor U11734 (N_11734,N_11219,N_11366);
and U11735 (N_11735,N_11359,N_11454);
nor U11736 (N_11736,N_11204,N_11238);
xor U11737 (N_11737,N_11314,N_11120);
nand U11738 (N_11738,N_11403,N_11237);
nand U11739 (N_11739,N_11213,N_11472);
nand U11740 (N_11740,N_11328,N_11177);
and U11741 (N_11741,N_11065,N_11405);
nor U11742 (N_11742,N_11089,N_11452);
xor U11743 (N_11743,N_11399,N_11155);
xnor U11744 (N_11744,N_11389,N_11478);
nor U11745 (N_11745,N_11349,N_11493);
and U11746 (N_11746,N_11117,N_11251);
nand U11747 (N_11747,N_11192,N_11282);
or U11748 (N_11748,N_11104,N_11442);
or U11749 (N_11749,N_11108,N_11074);
or U11750 (N_11750,N_11235,N_11164);
nor U11751 (N_11751,N_11413,N_11179);
or U11752 (N_11752,N_11138,N_11086);
xor U11753 (N_11753,N_11462,N_11092);
or U11754 (N_11754,N_11185,N_11034);
and U11755 (N_11755,N_11395,N_11044);
nand U11756 (N_11756,N_11103,N_11274);
nor U11757 (N_11757,N_11117,N_11437);
and U11758 (N_11758,N_11479,N_11206);
nand U11759 (N_11759,N_11028,N_11363);
nor U11760 (N_11760,N_11281,N_11419);
and U11761 (N_11761,N_11004,N_11317);
xor U11762 (N_11762,N_11055,N_11438);
xnor U11763 (N_11763,N_11244,N_11258);
nand U11764 (N_11764,N_11175,N_11256);
nand U11765 (N_11765,N_11249,N_11357);
or U11766 (N_11766,N_11201,N_11369);
nand U11767 (N_11767,N_11358,N_11123);
xnor U11768 (N_11768,N_11142,N_11166);
xnor U11769 (N_11769,N_11130,N_11223);
xor U11770 (N_11770,N_11447,N_11473);
and U11771 (N_11771,N_11074,N_11118);
nor U11772 (N_11772,N_11379,N_11142);
nor U11773 (N_11773,N_11437,N_11227);
or U11774 (N_11774,N_11097,N_11298);
and U11775 (N_11775,N_11145,N_11062);
and U11776 (N_11776,N_11000,N_11449);
nand U11777 (N_11777,N_11168,N_11234);
nor U11778 (N_11778,N_11297,N_11004);
nor U11779 (N_11779,N_11254,N_11195);
and U11780 (N_11780,N_11045,N_11130);
nor U11781 (N_11781,N_11395,N_11043);
xnor U11782 (N_11782,N_11113,N_11466);
and U11783 (N_11783,N_11211,N_11464);
or U11784 (N_11784,N_11184,N_11059);
or U11785 (N_11785,N_11107,N_11200);
nor U11786 (N_11786,N_11477,N_11434);
nand U11787 (N_11787,N_11356,N_11087);
nor U11788 (N_11788,N_11065,N_11176);
nor U11789 (N_11789,N_11383,N_11312);
nor U11790 (N_11790,N_11105,N_11271);
xnor U11791 (N_11791,N_11199,N_11311);
or U11792 (N_11792,N_11373,N_11383);
or U11793 (N_11793,N_11183,N_11104);
and U11794 (N_11794,N_11126,N_11295);
or U11795 (N_11795,N_11470,N_11086);
xor U11796 (N_11796,N_11263,N_11424);
or U11797 (N_11797,N_11343,N_11045);
nor U11798 (N_11798,N_11180,N_11127);
and U11799 (N_11799,N_11425,N_11330);
nand U11800 (N_11800,N_11000,N_11279);
nor U11801 (N_11801,N_11288,N_11338);
nor U11802 (N_11802,N_11378,N_11055);
nor U11803 (N_11803,N_11002,N_11460);
xor U11804 (N_11804,N_11318,N_11342);
nand U11805 (N_11805,N_11241,N_11273);
or U11806 (N_11806,N_11376,N_11377);
nand U11807 (N_11807,N_11232,N_11185);
xnor U11808 (N_11808,N_11318,N_11445);
nor U11809 (N_11809,N_11267,N_11156);
nor U11810 (N_11810,N_11098,N_11142);
nor U11811 (N_11811,N_11368,N_11003);
or U11812 (N_11812,N_11169,N_11495);
or U11813 (N_11813,N_11425,N_11024);
xor U11814 (N_11814,N_11373,N_11200);
and U11815 (N_11815,N_11309,N_11430);
or U11816 (N_11816,N_11021,N_11096);
nor U11817 (N_11817,N_11462,N_11016);
xor U11818 (N_11818,N_11404,N_11442);
nor U11819 (N_11819,N_11141,N_11305);
and U11820 (N_11820,N_11338,N_11428);
nand U11821 (N_11821,N_11150,N_11219);
xnor U11822 (N_11822,N_11416,N_11066);
and U11823 (N_11823,N_11384,N_11485);
nor U11824 (N_11824,N_11262,N_11197);
xnor U11825 (N_11825,N_11054,N_11220);
or U11826 (N_11826,N_11251,N_11293);
or U11827 (N_11827,N_11472,N_11421);
nor U11828 (N_11828,N_11258,N_11087);
nor U11829 (N_11829,N_11231,N_11093);
nor U11830 (N_11830,N_11044,N_11465);
xor U11831 (N_11831,N_11130,N_11461);
nor U11832 (N_11832,N_11424,N_11207);
nand U11833 (N_11833,N_11328,N_11141);
xnor U11834 (N_11834,N_11142,N_11489);
nor U11835 (N_11835,N_11284,N_11207);
or U11836 (N_11836,N_11285,N_11315);
nor U11837 (N_11837,N_11436,N_11259);
and U11838 (N_11838,N_11416,N_11282);
and U11839 (N_11839,N_11470,N_11281);
or U11840 (N_11840,N_11424,N_11419);
xnor U11841 (N_11841,N_11262,N_11356);
and U11842 (N_11842,N_11260,N_11315);
nor U11843 (N_11843,N_11039,N_11180);
or U11844 (N_11844,N_11171,N_11020);
nor U11845 (N_11845,N_11395,N_11472);
nor U11846 (N_11846,N_11258,N_11261);
or U11847 (N_11847,N_11420,N_11469);
and U11848 (N_11848,N_11025,N_11454);
or U11849 (N_11849,N_11015,N_11419);
xnor U11850 (N_11850,N_11339,N_11341);
or U11851 (N_11851,N_11455,N_11499);
and U11852 (N_11852,N_11200,N_11097);
xnor U11853 (N_11853,N_11480,N_11478);
nand U11854 (N_11854,N_11012,N_11455);
nand U11855 (N_11855,N_11048,N_11290);
or U11856 (N_11856,N_11277,N_11369);
and U11857 (N_11857,N_11349,N_11281);
nor U11858 (N_11858,N_11457,N_11046);
and U11859 (N_11859,N_11427,N_11441);
and U11860 (N_11860,N_11072,N_11446);
nor U11861 (N_11861,N_11456,N_11389);
and U11862 (N_11862,N_11493,N_11085);
or U11863 (N_11863,N_11180,N_11034);
xor U11864 (N_11864,N_11090,N_11495);
xnor U11865 (N_11865,N_11319,N_11113);
nor U11866 (N_11866,N_11089,N_11196);
and U11867 (N_11867,N_11175,N_11390);
and U11868 (N_11868,N_11362,N_11036);
nand U11869 (N_11869,N_11303,N_11048);
and U11870 (N_11870,N_11323,N_11198);
and U11871 (N_11871,N_11025,N_11096);
or U11872 (N_11872,N_11157,N_11422);
nor U11873 (N_11873,N_11043,N_11478);
xnor U11874 (N_11874,N_11276,N_11025);
or U11875 (N_11875,N_11055,N_11340);
nor U11876 (N_11876,N_11417,N_11361);
nor U11877 (N_11877,N_11237,N_11140);
and U11878 (N_11878,N_11033,N_11322);
xnor U11879 (N_11879,N_11097,N_11082);
and U11880 (N_11880,N_11383,N_11344);
and U11881 (N_11881,N_11034,N_11434);
and U11882 (N_11882,N_11039,N_11086);
nor U11883 (N_11883,N_11381,N_11336);
nor U11884 (N_11884,N_11104,N_11496);
nor U11885 (N_11885,N_11233,N_11156);
nand U11886 (N_11886,N_11102,N_11176);
or U11887 (N_11887,N_11496,N_11335);
and U11888 (N_11888,N_11196,N_11451);
xnor U11889 (N_11889,N_11467,N_11091);
nand U11890 (N_11890,N_11381,N_11176);
and U11891 (N_11891,N_11054,N_11033);
and U11892 (N_11892,N_11254,N_11097);
nand U11893 (N_11893,N_11460,N_11405);
nand U11894 (N_11894,N_11098,N_11182);
nand U11895 (N_11895,N_11261,N_11177);
and U11896 (N_11896,N_11015,N_11308);
xnor U11897 (N_11897,N_11476,N_11029);
or U11898 (N_11898,N_11043,N_11029);
xnor U11899 (N_11899,N_11281,N_11110);
nor U11900 (N_11900,N_11126,N_11460);
or U11901 (N_11901,N_11381,N_11165);
nor U11902 (N_11902,N_11182,N_11360);
and U11903 (N_11903,N_11373,N_11242);
nor U11904 (N_11904,N_11293,N_11236);
xor U11905 (N_11905,N_11485,N_11317);
and U11906 (N_11906,N_11426,N_11261);
xor U11907 (N_11907,N_11273,N_11169);
nor U11908 (N_11908,N_11415,N_11057);
and U11909 (N_11909,N_11381,N_11207);
or U11910 (N_11910,N_11453,N_11396);
or U11911 (N_11911,N_11277,N_11117);
or U11912 (N_11912,N_11278,N_11415);
xor U11913 (N_11913,N_11349,N_11325);
xnor U11914 (N_11914,N_11212,N_11094);
xnor U11915 (N_11915,N_11139,N_11050);
and U11916 (N_11916,N_11092,N_11033);
nor U11917 (N_11917,N_11271,N_11053);
or U11918 (N_11918,N_11302,N_11422);
nor U11919 (N_11919,N_11334,N_11192);
or U11920 (N_11920,N_11036,N_11296);
nor U11921 (N_11921,N_11474,N_11312);
or U11922 (N_11922,N_11089,N_11305);
xnor U11923 (N_11923,N_11024,N_11401);
nand U11924 (N_11924,N_11218,N_11475);
and U11925 (N_11925,N_11006,N_11058);
xor U11926 (N_11926,N_11237,N_11135);
and U11927 (N_11927,N_11144,N_11137);
nor U11928 (N_11928,N_11480,N_11472);
nor U11929 (N_11929,N_11252,N_11234);
or U11930 (N_11930,N_11060,N_11223);
nor U11931 (N_11931,N_11338,N_11062);
or U11932 (N_11932,N_11120,N_11195);
nand U11933 (N_11933,N_11044,N_11277);
nor U11934 (N_11934,N_11318,N_11114);
nor U11935 (N_11935,N_11373,N_11226);
and U11936 (N_11936,N_11176,N_11036);
nor U11937 (N_11937,N_11346,N_11058);
xor U11938 (N_11938,N_11122,N_11104);
xnor U11939 (N_11939,N_11215,N_11226);
or U11940 (N_11940,N_11273,N_11314);
and U11941 (N_11941,N_11444,N_11278);
xnor U11942 (N_11942,N_11225,N_11306);
or U11943 (N_11943,N_11464,N_11466);
and U11944 (N_11944,N_11366,N_11250);
nand U11945 (N_11945,N_11109,N_11253);
nand U11946 (N_11946,N_11077,N_11049);
and U11947 (N_11947,N_11185,N_11395);
or U11948 (N_11948,N_11004,N_11056);
or U11949 (N_11949,N_11462,N_11192);
or U11950 (N_11950,N_11326,N_11170);
nor U11951 (N_11951,N_11122,N_11038);
or U11952 (N_11952,N_11066,N_11041);
nor U11953 (N_11953,N_11192,N_11052);
nor U11954 (N_11954,N_11248,N_11306);
nand U11955 (N_11955,N_11234,N_11492);
xor U11956 (N_11956,N_11236,N_11229);
nand U11957 (N_11957,N_11348,N_11397);
or U11958 (N_11958,N_11403,N_11417);
and U11959 (N_11959,N_11483,N_11062);
and U11960 (N_11960,N_11359,N_11119);
nand U11961 (N_11961,N_11423,N_11088);
and U11962 (N_11962,N_11184,N_11323);
and U11963 (N_11963,N_11253,N_11291);
xor U11964 (N_11964,N_11362,N_11450);
xnor U11965 (N_11965,N_11097,N_11366);
nand U11966 (N_11966,N_11206,N_11063);
nor U11967 (N_11967,N_11009,N_11454);
xor U11968 (N_11968,N_11454,N_11213);
nand U11969 (N_11969,N_11268,N_11279);
or U11970 (N_11970,N_11405,N_11085);
xnor U11971 (N_11971,N_11002,N_11046);
nand U11972 (N_11972,N_11218,N_11137);
and U11973 (N_11973,N_11085,N_11424);
nand U11974 (N_11974,N_11380,N_11095);
xor U11975 (N_11975,N_11106,N_11215);
or U11976 (N_11976,N_11056,N_11138);
nor U11977 (N_11977,N_11470,N_11061);
and U11978 (N_11978,N_11030,N_11057);
and U11979 (N_11979,N_11201,N_11159);
and U11980 (N_11980,N_11024,N_11375);
or U11981 (N_11981,N_11460,N_11073);
or U11982 (N_11982,N_11349,N_11122);
or U11983 (N_11983,N_11488,N_11060);
nand U11984 (N_11984,N_11279,N_11299);
nand U11985 (N_11985,N_11369,N_11375);
nand U11986 (N_11986,N_11246,N_11303);
or U11987 (N_11987,N_11074,N_11166);
and U11988 (N_11988,N_11036,N_11446);
or U11989 (N_11989,N_11132,N_11247);
and U11990 (N_11990,N_11371,N_11229);
and U11991 (N_11991,N_11168,N_11262);
xnor U11992 (N_11992,N_11317,N_11145);
and U11993 (N_11993,N_11486,N_11013);
or U11994 (N_11994,N_11336,N_11180);
xor U11995 (N_11995,N_11238,N_11255);
nor U11996 (N_11996,N_11327,N_11497);
nand U11997 (N_11997,N_11495,N_11183);
xnor U11998 (N_11998,N_11267,N_11216);
xor U11999 (N_11999,N_11472,N_11173);
nor U12000 (N_12000,N_11848,N_11851);
nand U12001 (N_12001,N_11897,N_11528);
xor U12002 (N_12002,N_11920,N_11932);
nor U12003 (N_12003,N_11909,N_11625);
xnor U12004 (N_12004,N_11512,N_11551);
and U12005 (N_12005,N_11902,N_11925);
and U12006 (N_12006,N_11756,N_11919);
xor U12007 (N_12007,N_11542,N_11559);
nor U12008 (N_12008,N_11639,N_11739);
xnor U12009 (N_12009,N_11588,N_11899);
and U12010 (N_12010,N_11573,N_11650);
xnor U12011 (N_12011,N_11572,N_11627);
nand U12012 (N_12012,N_11679,N_11574);
nor U12013 (N_12013,N_11613,N_11640);
nor U12014 (N_12014,N_11963,N_11652);
nand U12015 (N_12015,N_11847,N_11991);
nand U12016 (N_12016,N_11808,N_11835);
nor U12017 (N_12017,N_11675,N_11669);
nand U12018 (N_12018,N_11630,N_11868);
and U12019 (N_12019,N_11700,N_11540);
or U12020 (N_12020,N_11961,N_11693);
nand U12021 (N_12021,N_11730,N_11837);
nand U12022 (N_12022,N_11803,N_11695);
nor U12023 (N_12023,N_11834,N_11629);
nand U12024 (N_12024,N_11880,N_11800);
or U12025 (N_12025,N_11710,N_11951);
xor U12026 (N_12026,N_11780,N_11998);
or U12027 (N_12027,N_11947,N_11738);
or U12028 (N_12028,N_11860,N_11624);
and U12029 (N_12029,N_11841,N_11724);
and U12030 (N_12030,N_11802,N_11770);
nor U12031 (N_12031,N_11832,N_11545);
or U12032 (N_12032,N_11744,N_11691);
nand U12033 (N_12033,N_11687,N_11760);
and U12034 (N_12034,N_11535,N_11748);
nor U12035 (N_12035,N_11642,N_11976);
nand U12036 (N_12036,N_11987,N_11591);
nor U12037 (N_12037,N_11912,N_11906);
xnor U12038 (N_12038,N_11798,N_11615);
xnor U12039 (N_12039,N_11531,N_11946);
and U12040 (N_12040,N_11578,N_11816);
nor U12041 (N_12041,N_11978,N_11933);
nand U12042 (N_12042,N_11564,N_11633);
nor U12043 (N_12043,N_11929,N_11890);
and U12044 (N_12044,N_11818,N_11930);
nand U12045 (N_12045,N_11656,N_11701);
xor U12046 (N_12046,N_11555,N_11715);
xor U12047 (N_12047,N_11955,N_11966);
nand U12048 (N_12048,N_11924,N_11733);
nand U12049 (N_12049,N_11567,N_11839);
nor U12050 (N_12050,N_11773,N_11943);
and U12051 (N_12051,N_11510,N_11603);
nand U12052 (N_12052,N_11529,N_11979);
nor U12053 (N_12053,N_11647,N_11741);
and U12054 (N_12054,N_11788,N_11637);
nor U12055 (N_12055,N_11654,N_11792);
or U12056 (N_12056,N_11942,N_11882);
xor U12057 (N_12057,N_11742,N_11774);
nor U12058 (N_12058,N_11984,N_11621);
nand U12059 (N_12059,N_11757,N_11673);
xor U12060 (N_12060,N_11922,N_11521);
nand U12061 (N_12061,N_11692,N_11634);
or U12062 (N_12062,N_11655,N_11846);
nor U12063 (N_12063,N_11905,N_11986);
or U12064 (N_12064,N_11599,N_11525);
xnor U12065 (N_12065,N_11826,N_11879);
or U12066 (N_12066,N_11505,N_11660);
and U12067 (N_12067,N_11815,N_11716);
nor U12068 (N_12068,N_11838,N_11936);
nand U12069 (N_12069,N_11901,N_11580);
and U12070 (N_12070,N_11791,N_11990);
and U12071 (N_12071,N_11611,N_11758);
xnor U12072 (N_12072,N_11607,N_11606);
and U12073 (N_12073,N_11950,N_11831);
xnor U12074 (N_12074,N_11889,N_11518);
or U12075 (N_12075,N_11814,N_11558);
and U12076 (N_12076,N_11549,N_11817);
nand U12077 (N_12077,N_11556,N_11843);
nor U12078 (N_12078,N_11534,N_11977);
nand U12079 (N_12079,N_11553,N_11938);
nor U12080 (N_12080,N_11579,N_11811);
xor U12081 (N_12081,N_11727,N_11997);
or U12082 (N_12082,N_11777,N_11644);
nand U12083 (N_12083,N_11728,N_11753);
or U12084 (N_12084,N_11543,N_11921);
or U12085 (N_12085,N_11911,N_11563);
nand U12086 (N_12086,N_11871,N_11520);
xnor U12087 (N_12087,N_11861,N_11807);
nor U12088 (N_12088,N_11891,N_11632);
nor U12089 (N_12089,N_11845,N_11853);
xor U12090 (N_12090,N_11796,N_11604);
or U12091 (N_12091,N_11527,N_11949);
or U12092 (N_12092,N_11994,N_11532);
nand U12093 (N_12093,N_11821,N_11928);
nor U12094 (N_12094,N_11988,N_11885);
or U12095 (N_12095,N_11504,N_11867);
nor U12096 (N_12096,N_11752,N_11643);
xnor U12097 (N_12097,N_11694,N_11702);
nor U12098 (N_12098,N_11734,N_11721);
nor U12099 (N_12099,N_11598,N_11971);
nor U12100 (N_12100,N_11849,N_11562);
xnor U12101 (N_12101,N_11590,N_11722);
or U12102 (N_12102,N_11648,N_11676);
or U12103 (N_12103,N_11863,N_11503);
nor U12104 (N_12104,N_11541,N_11893);
nand U12105 (N_12105,N_11511,N_11548);
or U12106 (N_12106,N_11517,N_11641);
or U12107 (N_12107,N_11959,N_11805);
nor U12108 (N_12108,N_11884,N_11539);
or U12109 (N_12109,N_11931,N_11554);
or U12110 (N_12110,N_11595,N_11664);
and U12111 (N_12111,N_11516,N_11619);
or U12112 (N_12112,N_11717,N_11769);
and U12113 (N_12113,N_11646,N_11618);
nand U12114 (N_12114,N_11689,N_11898);
nor U12115 (N_12115,N_11612,N_11530);
xor U12116 (N_12116,N_11859,N_11869);
xor U12117 (N_12117,N_11957,N_11965);
or U12118 (N_12118,N_11996,N_11718);
nand U12119 (N_12119,N_11740,N_11836);
xor U12120 (N_12120,N_11969,N_11833);
xor U12121 (N_12121,N_11690,N_11712);
and U12122 (N_12122,N_11824,N_11610);
nand U12123 (N_12123,N_11866,N_11508);
nand U12124 (N_12124,N_11678,N_11743);
and U12125 (N_12125,N_11674,N_11775);
nand U12126 (N_12126,N_11609,N_11887);
nor U12127 (N_12127,N_11751,N_11784);
and U12128 (N_12128,N_11729,N_11662);
nand U12129 (N_12129,N_11940,N_11723);
and U12130 (N_12130,N_11948,N_11763);
and U12131 (N_12131,N_11522,N_11623);
xor U12132 (N_12132,N_11820,N_11713);
xnor U12133 (N_12133,N_11571,N_11683);
or U12134 (N_12134,N_11636,N_11903);
nor U12135 (N_12135,N_11651,N_11585);
xnor U12136 (N_12136,N_11711,N_11794);
nand U12137 (N_12137,N_11680,N_11810);
nor U12138 (N_12138,N_11941,N_11628);
and U12139 (N_12139,N_11745,N_11536);
nor U12140 (N_12140,N_11685,N_11755);
nor U12141 (N_12141,N_11750,N_11876);
nand U12142 (N_12142,N_11703,N_11993);
or U12143 (N_12143,N_11953,N_11746);
nor U12144 (N_12144,N_11705,N_11915);
nand U12145 (N_12145,N_11557,N_11658);
xnor U12146 (N_12146,N_11981,N_11666);
nand U12147 (N_12147,N_11601,N_11875);
nand U12148 (N_12148,N_11787,N_11631);
or U12149 (N_12149,N_11954,N_11989);
nor U12150 (N_12150,N_11779,N_11561);
or U12151 (N_12151,N_11801,N_11550);
and U12152 (N_12152,N_11972,N_11560);
and U12153 (N_12153,N_11697,N_11668);
nand U12154 (N_12154,N_11638,N_11892);
nor U12155 (N_12155,N_11790,N_11914);
or U12156 (N_12156,N_11614,N_11747);
and U12157 (N_12157,N_11813,N_11663);
and U12158 (N_12158,N_11827,N_11570);
xnor U12159 (N_12159,N_11956,N_11513);
nor U12160 (N_12160,N_11622,N_11519);
nand U12161 (N_12161,N_11907,N_11895);
nand U12162 (N_12162,N_11985,N_11719);
nand U12163 (N_12163,N_11913,N_11785);
xnor U12164 (N_12164,N_11501,N_11576);
nand U12165 (N_12165,N_11605,N_11967);
or U12166 (N_12166,N_11962,N_11799);
nand U12167 (N_12167,N_11939,N_11789);
and U12168 (N_12168,N_11584,N_11533);
nor U12169 (N_12169,N_11686,N_11823);
or U12170 (N_12170,N_11857,N_11698);
nand U12171 (N_12171,N_11995,N_11569);
xnor U12172 (N_12172,N_11649,N_11538);
or U12173 (N_12173,N_11586,N_11749);
or U12174 (N_12174,N_11626,N_11776);
xor U12175 (N_12175,N_11688,N_11782);
nand U12176 (N_12176,N_11877,N_11594);
xor U12177 (N_12177,N_11781,N_11864);
nor U12178 (N_12178,N_11577,N_11944);
nand U12179 (N_12179,N_11926,N_11617);
and U12180 (N_12180,N_11506,N_11886);
and U12181 (N_12181,N_11980,N_11582);
and U12182 (N_12182,N_11523,N_11597);
nand U12183 (N_12183,N_11720,N_11795);
or U12184 (N_12184,N_11900,N_11865);
nand U12185 (N_12185,N_11968,N_11916);
or U12186 (N_12186,N_11767,N_11587);
and U12187 (N_12187,N_11819,N_11592);
or U12188 (N_12188,N_11754,N_11888);
nor U12189 (N_12189,N_11565,N_11896);
or U12190 (N_12190,N_11667,N_11546);
nand U12191 (N_12191,N_11927,N_11677);
and U12192 (N_12192,N_11681,N_11672);
or U12193 (N_12193,N_11575,N_11507);
xor U12194 (N_12194,N_11862,N_11772);
nand U12195 (N_12195,N_11706,N_11960);
nor U12196 (N_12196,N_11699,N_11937);
nand U12197 (N_12197,N_11502,N_11858);
and U12198 (N_12198,N_11958,N_11602);
nor U12199 (N_12199,N_11657,N_11684);
or U12200 (N_12200,N_11830,N_11975);
nand U12201 (N_12201,N_11894,N_11825);
and U12202 (N_12202,N_11544,N_11616);
nor U12203 (N_12203,N_11704,N_11771);
nand U12204 (N_12204,N_11589,N_11881);
and U12205 (N_12205,N_11515,N_11822);
or U12206 (N_12206,N_11970,N_11537);
nor U12207 (N_12207,N_11661,N_11804);
nor U12208 (N_12208,N_11854,N_11806);
nand U12209 (N_12209,N_11840,N_11952);
nand U12210 (N_12210,N_11793,N_11682);
nor U12211 (N_12211,N_11762,N_11736);
and U12212 (N_12212,N_11870,N_11620);
nor U12213 (N_12213,N_11500,N_11809);
or U12214 (N_12214,N_11526,N_11708);
xor U12215 (N_12215,N_11908,N_11765);
xnor U12216 (N_12216,N_11973,N_11737);
xnor U12217 (N_12217,N_11645,N_11910);
xnor U12218 (N_12218,N_11593,N_11874);
nand U12219 (N_12219,N_11778,N_11923);
and U12220 (N_12220,N_11581,N_11797);
and U12221 (N_12221,N_11917,N_11583);
xor U12222 (N_12222,N_11566,N_11735);
xnor U12223 (N_12223,N_11608,N_11709);
or U12224 (N_12224,N_11596,N_11935);
or U12225 (N_12225,N_11726,N_11600);
xor U12226 (N_12226,N_11828,N_11509);
xor U12227 (N_12227,N_11524,N_11872);
xor U12228 (N_12228,N_11635,N_11904);
or U12229 (N_12229,N_11918,N_11759);
or U12230 (N_12230,N_11761,N_11964);
and U12231 (N_12231,N_11732,N_11934);
nand U12232 (N_12232,N_11768,N_11552);
and U12233 (N_12233,N_11670,N_11992);
or U12234 (N_12234,N_11653,N_11983);
nor U12235 (N_12235,N_11878,N_11786);
nor U12236 (N_12236,N_11852,N_11665);
nand U12237 (N_12237,N_11783,N_11547);
xor U12238 (N_12238,N_11514,N_11568);
or U12239 (N_12239,N_11856,N_11842);
nand U12240 (N_12240,N_11659,N_11850);
or U12241 (N_12241,N_11982,N_11974);
or U12242 (N_12242,N_11873,N_11764);
xnor U12243 (N_12243,N_11829,N_11999);
nor U12244 (N_12244,N_11855,N_11731);
or U12245 (N_12245,N_11707,N_11812);
nand U12246 (N_12246,N_11766,N_11714);
nor U12247 (N_12247,N_11725,N_11883);
nand U12248 (N_12248,N_11671,N_11696);
nand U12249 (N_12249,N_11844,N_11945);
or U12250 (N_12250,N_11696,N_11617);
nand U12251 (N_12251,N_11817,N_11883);
or U12252 (N_12252,N_11907,N_11597);
nand U12253 (N_12253,N_11872,N_11822);
xnor U12254 (N_12254,N_11887,N_11831);
or U12255 (N_12255,N_11676,N_11894);
and U12256 (N_12256,N_11623,N_11607);
nor U12257 (N_12257,N_11593,N_11770);
and U12258 (N_12258,N_11606,N_11892);
nand U12259 (N_12259,N_11894,N_11801);
xor U12260 (N_12260,N_11870,N_11915);
nand U12261 (N_12261,N_11921,N_11804);
xor U12262 (N_12262,N_11720,N_11916);
xnor U12263 (N_12263,N_11819,N_11733);
or U12264 (N_12264,N_11745,N_11884);
nand U12265 (N_12265,N_11648,N_11982);
or U12266 (N_12266,N_11685,N_11976);
nor U12267 (N_12267,N_11766,N_11719);
xnor U12268 (N_12268,N_11890,N_11628);
and U12269 (N_12269,N_11891,N_11620);
and U12270 (N_12270,N_11719,N_11763);
xnor U12271 (N_12271,N_11644,N_11887);
or U12272 (N_12272,N_11965,N_11587);
xor U12273 (N_12273,N_11958,N_11695);
nor U12274 (N_12274,N_11550,N_11856);
nand U12275 (N_12275,N_11642,N_11568);
and U12276 (N_12276,N_11882,N_11508);
and U12277 (N_12277,N_11836,N_11771);
and U12278 (N_12278,N_11651,N_11905);
or U12279 (N_12279,N_11905,N_11785);
nor U12280 (N_12280,N_11951,N_11846);
or U12281 (N_12281,N_11760,N_11647);
xnor U12282 (N_12282,N_11584,N_11798);
nor U12283 (N_12283,N_11648,N_11774);
or U12284 (N_12284,N_11541,N_11708);
xnor U12285 (N_12285,N_11587,N_11853);
or U12286 (N_12286,N_11769,N_11624);
nand U12287 (N_12287,N_11832,N_11899);
nand U12288 (N_12288,N_11804,N_11674);
nor U12289 (N_12289,N_11871,N_11867);
or U12290 (N_12290,N_11540,N_11513);
or U12291 (N_12291,N_11617,N_11758);
nand U12292 (N_12292,N_11730,N_11500);
or U12293 (N_12293,N_11903,N_11877);
or U12294 (N_12294,N_11868,N_11761);
xnor U12295 (N_12295,N_11706,N_11894);
nand U12296 (N_12296,N_11698,N_11644);
nor U12297 (N_12297,N_11766,N_11755);
nand U12298 (N_12298,N_11617,N_11795);
or U12299 (N_12299,N_11744,N_11554);
or U12300 (N_12300,N_11845,N_11937);
nor U12301 (N_12301,N_11636,N_11732);
and U12302 (N_12302,N_11679,N_11855);
or U12303 (N_12303,N_11793,N_11907);
nor U12304 (N_12304,N_11969,N_11595);
and U12305 (N_12305,N_11793,N_11835);
or U12306 (N_12306,N_11724,N_11776);
or U12307 (N_12307,N_11903,N_11835);
nand U12308 (N_12308,N_11680,N_11503);
xor U12309 (N_12309,N_11788,N_11869);
or U12310 (N_12310,N_11695,N_11621);
xor U12311 (N_12311,N_11868,N_11582);
nor U12312 (N_12312,N_11948,N_11951);
xor U12313 (N_12313,N_11514,N_11936);
or U12314 (N_12314,N_11644,N_11561);
nor U12315 (N_12315,N_11997,N_11814);
xor U12316 (N_12316,N_11849,N_11824);
and U12317 (N_12317,N_11777,N_11525);
or U12318 (N_12318,N_11750,N_11591);
or U12319 (N_12319,N_11723,N_11830);
and U12320 (N_12320,N_11741,N_11868);
nor U12321 (N_12321,N_11611,N_11504);
nand U12322 (N_12322,N_11789,N_11852);
and U12323 (N_12323,N_11885,N_11995);
or U12324 (N_12324,N_11576,N_11694);
nor U12325 (N_12325,N_11660,N_11616);
nor U12326 (N_12326,N_11642,N_11940);
nor U12327 (N_12327,N_11665,N_11945);
or U12328 (N_12328,N_11716,N_11694);
and U12329 (N_12329,N_11986,N_11633);
nor U12330 (N_12330,N_11741,N_11593);
xnor U12331 (N_12331,N_11726,N_11807);
nor U12332 (N_12332,N_11960,N_11844);
nor U12333 (N_12333,N_11543,N_11787);
and U12334 (N_12334,N_11722,N_11671);
or U12335 (N_12335,N_11513,N_11658);
nor U12336 (N_12336,N_11900,N_11846);
and U12337 (N_12337,N_11882,N_11939);
nor U12338 (N_12338,N_11786,N_11851);
nor U12339 (N_12339,N_11509,N_11521);
and U12340 (N_12340,N_11964,N_11907);
and U12341 (N_12341,N_11969,N_11816);
nor U12342 (N_12342,N_11783,N_11788);
nand U12343 (N_12343,N_11810,N_11907);
or U12344 (N_12344,N_11727,N_11971);
or U12345 (N_12345,N_11770,N_11908);
nand U12346 (N_12346,N_11649,N_11586);
nor U12347 (N_12347,N_11719,N_11614);
or U12348 (N_12348,N_11682,N_11605);
xnor U12349 (N_12349,N_11573,N_11956);
nor U12350 (N_12350,N_11614,N_11900);
nor U12351 (N_12351,N_11870,N_11747);
nor U12352 (N_12352,N_11797,N_11800);
xor U12353 (N_12353,N_11593,N_11968);
nand U12354 (N_12354,N_11638,N_11659);
nand U12355 (N_12355,N_11933,N_11599);
nor U12356 (N_12356,N_11972,N_11890);
nand U12357 (N_12357,N_11933,N_11739);
or U12358 (N_12358,N_11762,N_11601);
and U12359 (N_12359,N_11842,N_11816);
and U12360 (N_12360,N_11772,N_11580);
nand U12361 (N_12361,N_11892,N_11791);
nand U12362 (N_12362,N_11598,N_11831);
and U12363 (N_12363,N_11637,N_11596);
nand U12364 (N_12364,N_11832,N_11537);
and U12365 (N_12365,N_11521,N_11654);
or U12366 (N_12366,N_11746,N_11956);
nor U12367 (N_12367,N_11649,N_11606);
nand U12368 (N_12368,N_11727,N_11634);
xnor U12369 (N_12369,N_11764,N_11723);
nor U12370 (N_12370,N_11613,N_11872);
or U12371 (N_12371,N_11834,N_11939);
or U12372 (N_12372,N_11696,N_11602);
nor U12373 (N_12373,N_11788,N_11560);
nand U12374 (N_12374,N_11894,N_11507);
nor U12375 (N_12375,N_11901,N_11727);
nor U12376 (N_12376,N_11631,N_11942);
or U12377 (N_12377,N_11566,N_11959);
nor U12378 (N_12378,N_11855,N_11532);
xor U12379 (N_12379,N_11684,N_11949);
or U12380 (N_12380,N_11642,N_11775);
nand U12381 (N_12381,N_11855,N_11854);
xnor U12382 (N_12382,N_11972,N_11940);
nand U12383 (N_12383,N_11640,N_11538);
nor U12384 (N_12384,N_11679,N_11504);
xnor U12385 (N_12385,N_11629,N_11811);
nand U12386 (N_12386,N_11746,N_11629);
xor U12387 (N_12387,N_11782,N_11676);
and U12388 (N_12388,N_11589,N_11991);
and U12389 (N_12389,N_11511,N_11718);
nand U12390 (N_12390,N_11873,N_11519);
or U12391 (N_12391,N_11629,N_11832);
nor U12392 (N_12392,N_11638,N_11662);
or U12393 (N_12393,N_11588,N_11982);
and U12394 (N_12394,N_11809,N_11841);
nor U12395 (N_12395,N_11680,N_11940);
nand U12396 (N_12396,N_11607,N_11952);
nand U12397 (N_12397,N_11685,N_11851);
and U12398 (N_12398,N_11718,N_11968);
and U12399 (N_12399,N_11823,N_11904);
or U12400 (N_12400,N_11981,N_11959);
xor U12401 (N_12401,N_11526,N_11975);
and U12402 (N_12402,N_11887,N_11819);
nor U12403 (N_12403,N_11707,N_11926);
nand U12404 (N_12404,N_11642,N_11986);
nand U12405 (N_12405,N_11749,N_11990);
and U12406 (N_12406,N_11728,N_11805);
xor U12407 (N_12407,N_11501,N_11515);
xnor U12408 (N_12408,N_11820,N_11714);
and U12409 (N_12409,N_11790,N_11588);
and U12410 (N_12410,N_11690,N_11762);
nor U12411 (N_12411,N_11878,N_11880);
or U12412 (N_12412,N_11539,N_11774);
or U12413 (N_12413,N_11843,N_11585);
or U12414 (N_12414,N_11997,N_11755);
nor U12415 (N_12415,N_11793,N_11573);
nand U12416 (N_12416,N_11575,N_11878);
nor U12417 (N_12417,N_11647,N_11855);
nand U12418 (N_12418,N_11592,N_11793);
nor U12419 (N_12419,N_11957,N_11568);
and U12420 (N_12420,N_11840,N_11936);
xnor U12421 (N_12421,N_11946,N_11738);
and U12422 (N_12422,N_11818,N_11978);
xnor U12423 (N_12423,N_11944,N_11889);
nor U12424 (N_12424,N_11675,N_11606);
and U12425 (N_12425,N_11610,N_11774);
or U12426 (N_12426,N_11580,N_11731);
or U12427 (N_12427,N_11676,N_11710);
or U12428 (N_12428,N_11815,N_11537);
xor U12429 (N_12429,N_11726,N_11776);
nor U12430 (N_12430,N_11701,N_11786);
xor U12431 (N_12431,N_11733,N_11935);
or U12432 (N_12432,N_11745,N_11665);
xor U12433 (N_12433,N_11619,N_11840);
nand U12434 (N_12434,N_11585,N_11753);
xor U12435 (N_12435,N_11745,N_11593);
or U12436 (N_12436,N_11848,N_11767);
and U12437 (N_12437,N_11657,N_11816);
nor U12438 (N_12438,N_11847,N_11532);
xor U12439 (N_12439,N_11880,N_11782);
nor U12440 (N_12440,N_11936,N_11571);
and U12441 (N_12441,N_11908,N_11976);
and U12442 (N_12442,N_11705,N_11675);
nor U12443 (N_12443,N_11730,N_11644);
or U12444 (N_12444,N_11809,N_11865);
or U12445 (N_12445,N_11814,N_11584);
xor U12446 (N_12446,N_11643,N_11591);
and U12447 (N_12447,N_11592,N_11849);
or U12448 (N_12448,N_11537,N_11779);
nand U12449 (N_12449,N_11950,N_11980);
nand U12450 (N_12450,N_11572,N_11901);
xnor U12451 (N_12451,N_11829,N_11897);
nor U12452 (N_12452,N_11793,N_11633);
and U12453 (N_12453,N_11727,N_11798);
and U12454 (N_12454,N_11951,N_11764);
or U12455 (N_12455,N_11517,N_11902);
or U12456 (N_12456,N_11661,N_11959);
and U12457 (N_12457,N_11680,N_11654);
nor U12458 (N_12458,N_11672,N_11546);
and U12459 (N_12459,N_11625,N_11864);
nand U12460 (N_12460,N_11734,N_11951);
xor U12461 (N_12461,N_11779,N_11501);
and U12462 (N_12462,N_11732,N_11796);
nand U12463 (N_12463,N_11685,N_11528);
xnor U12464 (N_12464,N_11737,N_11839);
nor U12465 (N_12465,N_11958,N_11764);
or U12466 (N_12466,N_11956,N_11589);
xnor U12467 (N_12467,N_11619,N_11954);
nor U12468 (N_12468,N_11624,N_11670);
or U12469 (N_12469,N_11628,N_11892);
and U12470 (N_12470,N_11945,N_11662);
nand U12471 (N_12471,N_11725,N_11926);
nor U12472 (N_12472,N_11782,N_11761);
nor U12473 (N_12473,N_11574,N_11806);
xor U12474 (N_12474,N_11603,N_11600);
or U12475 (N_12475,N_11824,N_11873);
nand U12476 (N_12476,N_11919,N_11640);
xor U12477 (N_12477,N_11704,N_11764);
and U12478 (N_12478,N_11860,N_11838);
nand U12479 (N_12479,N_11755,N_11877);
nor U12480 (N_12480,N_11914,N_11913);
nor U12481 (N_12481,N_11693,N_11778);
xnor U12482 (N_12482,N_11961,N_11925);
or U12483 (N_12483,N_11750,N_11942);
xor U12484 (N_12484,N_11503,N_11619);
or U12485 (N_12485,N_11842,N_11991);
and U12486 (N_12486,N_11598,N_11507);
or U12487 (N_12487,N_11552,N_11837);
and U12488 (N_12488,N_11631,N_11567);
nand U12489 (N_12489,N_11799,N_11674);
or U12490 (N_12490,N_11717,N_11875);
or U12491 (N_12491,N_11826,N_11913);
or U12492 (N_12492,N_11870,N_11503);
nor U12493 (N_12493,N_11717,N_11888);
or U12494 (N_12494,N_11526,N_11984);
xor U12495 (N_12495,N_11547,N_11698);
or U12496 (N_12496,N_11510,N_11873);
or U12497 (N_12497,N_11611,N_11737);
or U12498 (N_12498,N_11882,N_11908);
nand U12499 (N_12499,N_11562,N_11710);
nor U12500 (N_12500,N_12401,N_12046);
or U12501 (N_12501,N_12071,N_12354);
or U12502 (N_12502,N_12229,N_12481);
nand U12503 (N_12503,N_12063,N_12365);
nand U12504 (N_12504,N_12259,N_12136);
and U12505 (N_12505,N_12329,N_12215);
nand U12506 (N_12506,N_12435,N_12403);
nor U12507 (N_12507,N_12393,N_12429);
xor U12508 (N_12508,N_12366,N_12019);
nor U12509 (N_12509,N_12073,N_12317);
and U12510 (N_12510,N_12166,N_12474);
and U12511 (N_12511,N_12367,N_12271);
xnor U12512 (N_12512,N_12458,N_12344);
xor U12513 (N_12513,N_12488,N_12133);
xor U12514 (N_12514,N_12285,N_12316);
nand U12515 (N_12515,N_12235,N_12418);
nor U12516 (N_12516,N_12269,N_12041);
or U12517 (N_12517,N_12203,N_12146);
and U12518 (N_12518,N_12086,N_12011);
nand U12519 (N_12519,N_12070,N_12113);
nand U12520 (N_12520,N_12274,N_12424);
or U12521 (N_12521,N_12022,N_12192);
nand U12522 (N_12522,N_12137,N_12441);
nor U12523 (N_12523,N_12395,N_12094);
nor U12524 (N_12524,N_12260,N_12195);
and U12525 (N_12525,N_12152,N_12191);
nand U12526 (N_12526,N_12079,N_12357);
and U12527 (N_12527,N_12258,N_12278);
and U12528 (N_12528,N_12287,N_12108);
nor U12529 (N_12529,N_12382,N_12480);
nand U12530 (N_12530,N_12331,N_12369);
and U12531 (N_12531,N_12005,N_12358);
nor U12532 (N_12532,N_12110,N_12225);
and U12533 (N_12533,N_12330,N_12179);
nor U12534 (N_12534,N_12163,N_12302);
xor U12535 (N_12535,N_12037,N_12123);
nor U12536 (N_12536,N_12056,N_12135);
xnor U12537 (N_12537,N_12157,N_12456);
nor U12538 (N_12538,N_12476,N_12010);
and U12539 (N_12539,N_12262,N_12144);
and U12540 (N_12540,N_12104,N_12340);
nor U12541 (N_12541,N_12018,N_12082);
and U12542 (N_12542,N_12003,N_12077);
nor U12543 (N_12543,N_12143,N_12318);
nand U12544 (N_12544,N_12402,N_12155);
nor U12545 (N_12545,N_12413,N_12031);
nand U12546 (N_12546,N_12176,N_12292);
nor U12547 (N_12547,N_12351,N_12112);
xor U12548 (N_12548,N_12220,N_12058);
nand U12549 (N_12549,N_12178,N_12069);
or U12550 (N_12550,N_12015,N_12106);
nand U12551 (N_12551,N_12439,N_12045);
xnor U12552 (N_12552,N_12012,N_12428);
and U12553 (N_12553,N_12291,N_12383);
xor U12554 (N_12554,N_12423,N_12490);
or U12555 (N_12555,N_12475,N_12341);
nor U12556 (N_12556,N_12328,N_12371);
and U12557 (N_12557,N_12335,N_12312);
nor U12558 (N_12558,N_12414,N_12283);
nand U12559 (N_12559,N_12160,N_12391);
and U12560 (N_12560,N_12360,N_12432);
nand U12561 (N_12561,N_12333,N_12057);
nor U12562 (N_12562,N_12245,N_12405);
xor U12563 (N_12563,N_12232,N_12088);
or U12564 (N_12564,N_12009,N_12489);
and U12565 (N_12565,N_12452,N_12187);
or U12566 (N_12566,N_12255,N_12281);
nand U12567 (N_12567,N_12483,N_12089);
xnor U12568 (N_12568,N_12052,N_12267);
and U12569 (N_12569,N_12184,N_12059);
xnor U12570 (N_12570,N_12427,N_12487);
and U12571 (N_12571,N_12068,N_12445);
nor U12572 (N_12572,N_12120,N_12398);
nor U12573 (N_12573,N_12219,N_12381);
nand U12574 (N_12574,N_12349,N_12313);
nor U12575 (N_12575,N_12115,N_12242);
and U12576 (N_12576,N_12356,N_12327);
and U12577 (N_12577,N_12226,N_12223);
or U12578 (N_12578,N_12126,N_12270);
nand U12579 (N_12579,N_12492,N_12170);
xnor U12580 (N_12580,N_12433,N_12197);
nor U12581 (N_12581,N_12091,N_12023);
xor U12582 (N_12582,N_12156,N_12017);
or U12583 (N_12583,N_12127,N_12224);
xnor U12584 (N_12584,N_12114,N_12420);
nand U12585 (N_12585,N_12043,N_12185);
nand U12586 (N_12586,N_12380,N_12392);
nand U12587 (N_12587,N_12048,N_12298);
and U12588 (N_12588,N_12499,N_12305);
and U12589 (N_12589,N_12442,N_12062);
or U12590 (N_12590,N_12254,N_12199);
and U12591 (N_12591,N_12096,N_12284);
and U12592 (N_12592,N_12040,N_12250);
nand U12593 (N_12593,N_12465,N_12026);
nand U12594 (N_12594,N_12411,N_12213);
xnor U12595 (N_12595,N_12308,N_12081);
nand U12596 (N_12596,N_12374,N_12246);
and U12597 (N_12597,N_12373,N_12189);
and U12598 (N_12598,N_12454,N_12438);
or U12599 (N_12599,N_12347,N_12422);
nand U12600 (N_12600,N_12378,N_12322);
and U12601 (N_12601,N_12303,N_12129);
nor U12602 (N_12602,N_12496,N_12072);
or U12603 (N_12603,N_12007,N_12247);
xnor U12604 (N_12604,N_12440,N_12416);
xor U12605 (N_12605,N_12389,N_12482);
and U12606 (N_12606,N_12093,N_12447);
xnor U12607 (N_12607,N_12065,N_12066);
xnor U12608 (N_12608,N_12034,N_12362);
nor U12609 (N_12609,N_12139,N_12148);
or U12610 (N_12610,N_12460,N_12338);
and U12611 (N_12611,N_12122,N_12206);
nand U12612 (N_12612,N_12299,N_12241);
and U12613 (N_12613,N_12103,N_12307);
and U12614 (N_12614,N_12154,N_12297);
and U12615 (N_12615,N_12293,N_12196);
and U12616 (N_12616,N_12234,N_12060);
nor U12617 (N_12617,N_12061,N_12171);
nand U12618 (N_12618,N_12159,N_12484);
xor U12619 (N_12619,N_12263,N_12463);
nand U12620 (N_12620,N_12013,N_12055);
nand U12621 (N_12621,N_12032,N_12147);
xor U12622 (N_12622,N_12453,N_12355);
or U12623 (N_12623,N_12397,N_12211);
or U12624 (N_12624,N_12231,N_12486);
nand U12625 (N_12625,N_12468,N_12001);
nand U12626 (N_12626,N_12132,N_12352);
and U12627 (N_12627,N_12109,N_12205);
and U12628 (N_12628,N_12124,N_12310);
nor U12629 (N_12629,N_12078,N_12400);
nand U12630 (N_12630,N_12105,N_12167);
or U12631 (N_12631,N_12377,N_12087);
xor U12632 (N_12632,N_12473,N_12212);
and U12633 (N_12633,N_12464,N_12044);
or U12634 (N_12634,N_12183,N_12346);
nand U12635 (N_12635,N_12150,N_12296);
nor U12636 (N_12636,N_12158,N_12200);
xnor U12637 (N_12637,N_12051,N_12099);
nand U12638 (N_12638,N_12387,N_12319);
nand U12639 (N_12639,N_12384,N_12497);
xor U12640 (N_12640,N_12261,N_12240);
or U12641 (N_12641,N_12425,N_12020);
or U12642 (N_12642,N_12151,N_12016);
or U12643 (N_12643,N_12207,N_12042);
or U12644 (N_12644,N_12233,N_12201);
or U12645 (N_12645,N_12165,N_12290);
nor U12646 (N_12646,N_12326,N_12478);
nand U12647 (N_12647,N_12006,N_12116);
nand U12648 (N_12648,N_12268,N_12372);
nand U12649 (N_12649,N_12090,N_12021);
nand U12650 (N_12650,N_12238,N_12498);
xnor U12651 (N_12651,N_12080,N_12332);
xnor U12652 (N_12652,N_12054,N_12415);
and U12653 (N_12653,N_12208,N_12406);
and U12654 (N_12654,N_12138,N_12162);
nand U12655 (N_12655,N_12265,N_12444);
xor U12656 (N_12656,N_12097,N_12353);
nor U12657 (N_12657,N_12153,N_12202);
or U12658 (N_12658,N_12095,N_12248);
nor U12659 (N_12659,N_12495,N_12198);
and U12660 (N_12660,N_12450,N_12469);
nand U12661 (N_12661,N_12479,N_12188);
nor U12662 (N_12662,N_12455,N_12204);
nand U12663 (N_12663,N_12494,N_12027);
and U12664 (N_12664,N_12343,N_12304);
nor U12665 (N_12665,N_12277,N_12128);
or U12666 (N_12666,N_12074,N_12471);
and U12667 (N_12667,N_12323,N_12396);
nor U12668 (N_12668,N_12222,N_12436);
xnor U12669 (N_12669,N_12337,N_12430);
nor U12670 (N_12670,N_12002,N_12085);
nor U12671 (N_12671,N_12361,N_12239);
and U12672 (N_12672,N_12190,N_12272);
xnor U12673 (N_12673,N_12121,N_12325);
xor U12674 (N_12674,N_12467,N_12100);
and U12675 (N_12675,N_12014,N_12379);
or U12676 (N_12676,N_12294,N_12142);
or U12677 (N_12677,N_12098,N_12092);
nor U12678 (N_12678,N_12030,N_12174);
or U12679 (N_12679,N_12491,N_12049);
nand U12680 (N_12680,N_12459,N_12193);
nand U12681 (N_12681,N_12407,N_12446);
xor U12682 (N_12682,N_12408,N_12388);
or U12683 (N_12683,N_12359,N_12449);
or U12684 (N_12684,N_12172,N_12145);
and U12685 (N_12685,N_12161,N_12177);
or U12686 (N_12686,N_12461,N_12107);
and U12687 (N_12687,N_12493,N_12025);
xnor U12688 (N_12688,N_12364,N_12466);
xnor U12689 (N_12689,N_12300,N_12140);
and U12690 (N_12690,N_12306,N_12035);
nand U12691 (N_12691,N_12181,N_12472);
and U12692 (N_12692,N_12209,N_12409);
or U12693 (N_12693,N_12311,N_12173);
nand U12694 (N_12694,N_12214,N_12053);
or U12695 (N_12695,N_12036,N_12218);
nor U12696 (N_12696,N_12350,N_12175);
and U12697 (N_12697,N_12180,N_12102);
or U12698 (N_12698,N_12434,N_12288);
xor U12699 (N_12699,N_12426,N_12394);
or U12700 (N_12700,N_12216,N_12348);
and U12701 (N_12701,N_12280,N_12370);
or U12702 (N_12702,N_12169,N_12399);
or U12703 (N_12703,N_12038,N_12485);
xor U12704 (N_12704,N_12470,N_12314);
nand U12705 (N_12705,N_12342,N_12028);
or U12706 (N_12706,N_12264,N_12324);
nand U12707 (N_12707,N_12320,N_12033);
and U12708 (N_12708,N_12286,N_12462);
xor U12709 (N_12709,N_12279,N_12321);
and U12710 (N_12710,N_12168,N_12273);
xnor U12711 (N_12711,N_12363,N_12421);
nor U12712 (N_12712,N_12282,N_12275);
xnor U12713 (N_12713,N_12039,N_12024);
xnor U12714 (N_12714,N_12130,N_12417);
and U12715 (N_12715,N_12230,N_12276);
xor U12716 (N_12716,N_12210,N_12228);
or U12717 (N_12717,N_12131,N_12125);
xor U12718 (N_12718,N_12050,N_12243);
xor U12719 (N_12719,N_12194,N_12118);
and U12720 (N_12720,N_12345,N_12227);
or U12721 (N_12721,N_12075,N_12149);
nand U12722 (N_12722,N_12004,N_12237);
and U12723 (N_12723,N_12252,N_12376);
xor U12724 (N_12724,N_12217,N_12000);
nor U12725 (N_12725,N_12244,N_12111);
or U12726 (N_12726,N_12477,N_12257);
or U12727 (N_12727,N_12315,N_12412);
or U12728 (N_12728,N_12141,N_12084);
nand U12729 (N_12729,N_12134,N_12431);
nor U12730 (N_12730,N_12386,N_12119);
nor U12731 (N_12731,N_12251,N_12375);
and U12732 (N_12732,N_12253,N_12256);
nand U12733 (N_12733,N_12164,N_12064);
nand U12734 (N_12734,N_12443,N_12008);
and U12735 (N_12735,N_12368,N_12457);
or U12736 (N_12736,N_12047,N_12117);
and U12737 (N_12737,N_12083,N_12410);
nor U12738 (N_12738,N_12404,N_12289);
or U12739 (N_12739,N_12067,N_12295);
nor U12740 (N_12740,N_12236,N_12221);
nor U12741 (N_12741,N_12266,N_12182);
nand U12742 (N_12742,N_12186,N_12419);
and U12743 (N_12743,N_12437,N_12451);
nor U12744 (N_12744,N_12339,N_12336);
and U12745 (N_12745,N_12101,N_12249);
and U12746 (N_12746,N_12029,N_12390);
and U12747 (N_12747,N_12301,N_12385);
nor U12748 (N_12748,N_12309,N_12334);
or U12749 (N_12749,N_12448,N_12076);
nor U12750 (N_12750,N_12396,N_12449);
nor U12751 (N_12751,N_12019,N_12048);
nor U12752 (N_12752,N_12023,N_12293);
xnor U12753 (N_12753,N_12309,N_12316);
xor U12754 (N_12754,N_12119,N_12398);
xor U12755 (N_12755,N_12177,N_12214);
and U12756 (N_12756,N_12101,N_12325);
xnor U12757 (N_12757,N_12468,N_12103);
or U12758 (N_12758,N_12345,N_12268);
nor U12759 (N_12759,N_12138,N_12386);
xnor U12760 (N_12760,N_12465,N_12440);
xnor U12761 (N_12761,N_12068,N_12117);
and U12762 (N_12762,N_12340,N_12074);
and U12763 (N_12763,N_12492,N_12276);
nand U12764 (N_12764,N_12373,N_12447);
or U12765 (N_12765,N_12447,N_12217);
nor U12766 (N_12766,N_12269,N_12292);
or U12767 (N_12767,N_12128,N_12043);
nor U12768 (N_12768,N_12401,N_12057);
xor U12769 (N_12769,N_12366,N_12154);
or U12770 (N_12770,N_12293,N_12331);
or U12771 (N_12771,N_12364,N_12473);
nand U12772 (N_12772,N_12337,N_12194);
xnor U12773 (N_12773,N_12177,N_12287);
nand U12774 (N_12774,N_12038,N_12117);
xor U12775 (N_12775,N_12394,N_12487);
nor U12776 (N_12776,N_12222,N_12021);
xor U12777 (N_12777,N_12109,N_12215);
and U12778 (N_12778,N_12396,N_12499);
or U12779 (N_12779,N_12356,N_12313);
and U12780 (N_12780,N_12056,N_12235);
and U12781 (N_12781,N_12029,N_12005);
and U12782 (N_12782,N_12028,N_12366);
or U12783 (N_12783,N_12056,N_12349);
nand U12784 (N_12784,N_12351,N_12341);
and U12785 (N_12785,N_12144,N_12034);
nand U12786 (N_12786,N_12047,N_12245);
nor U12787 (N_12787,N_12331,N_12377);
xor U12788 (N_12788,N_12334,N_12350);
xnor U12789 (N_12789,N_12470,N_12334);
nor U12790 (N_12790,N_12398,N_12295);
or U12791 (N_12791,N_12309,N_12157);
nand U12792 (N_12792,N_12378,N_12174);
and U12793 (N_12793,N_12495,N_12267);
and U12794 (N_12794,N_12204,N_12309);
nor U12795 (N_12795,N_12100,N_12320);
xor U12796 (N_12796,N_12343,N_12483);
nor U12797 (N_12797,N_12392,N_12494);
or U12798 (N_12798,N_12449,N_12312);
xor U12799 (N_12799,N_12004,N_12363);
xor U12800 (N_12800,N_12058,N_12172);
or U12801 (N_12801,N_12008,N_12230);
or U12802 (N_12802,N_12153,N_12015);
nand U12803 (N_12803,N_12190,N_12092);
and U12804 (N_12804,N_12195,N_12363);
and U12805 (N_12805,N_12447,N_12395);
xnor U12806 (N_12806,N_12342,N_12324);
nand U12807 (N_12807,N_12102,N_12455);
nor U12808 (N_12808,N_12401,N_12072);
or U12809 (N_12809,N_12003,N_12112);
nand U12810 (N_12810,N_12292,N_12227);
nor U12811 (N_12811,N_12141,N_12274);
and U12812 (N_12812,N_12087,N_12213);
or U12813 (N_12813,N_12118,N_12161);
xnor U12814 (N_12814,N_12039,N_12206);
xor U12815 (N_12815,N_12185,N_12181);
xor U12816 (N_12816,N_12161,N_12349);
nand U12817 (N_12817,N_12047,N_12310);
and U12818 (N_12818,N_12265,N_12179);
or U12819 (N_12819,N_12163,N_12006);
nor U12820 (N_12820,N_12429,N_12084);
nand U12821 (N_12821,N_12192,N_12237);
and U12822 (N_12822,N_12265,N_12115);
and U12823 (N_12823,N_12363,N_12424);
xnor U12824 (N_12824,N_12119,N_12091);
nor U12825 (N_12825,N_12331,N_12312);
and U12826 (N_12826,N_12193,N_12177);
or U12827 (N_12827,N_12369,N_12484);
nor U12828 (N_12828,N_12015,N_12462);
and U12829 (N_12829,N_12238,N_12198);
nand U12830 (N_12830,N_12031,N_12132);
and U12831 (N_12831,N_12402,N_12078);
nor U12832 (N_12832,N_12163,N_12066);
nand U12833 (N_12833,N_12188,N_12308);
and U12834 (N_12834,N_12295,N_12346);
nand U12835 (N_12835,N_12459,N_12291);
nand U12836 (N_12836,N_12232,N_12205);
nor U12837 (N_12837,N_12133,N_12409);
and U12838 (N_12838,N_12355,N_12147);
nand U12839 (N_12839,N_12148,N_12021);
nor U12840 (N_12840,N_12430,N_12227);
nand U12841 (N_12841,N_12387,N_12431);
nand U12842 (N_12842,N_12348,N_12214);
nor U12843 (N_12843,N_12207,N_12407);
or U12844 (N_12844,N_12006,N_12033);
and U12845 (N_12845,N_12351,N_12155);
nor U12846 (N_12846,N_12356,N_12442);
and U12847 (N_12847,N_12353,N_12134);
xor U12848 (N_12848,N_12377,N_12328);
xnor U12849 (N_12849,N_12351,N_12357);
xnor U12850 (N_12850,N_12499,N_12121);
nand U12851 (N_12851,N_12294,N_12009);
nand U12852 (N_12852,N_12400,N_12383);
or U12853 (N_12853,N_12362,N_12116);
or U12854 (N_12854,N_12213,N_12028);
or U12855 (N_12855,N_12377,N_12060);
nor U12856 (N_12856,N_12433,N_12403);
and U12857 (N_12857,N_12230,N_12192);
and U12858 (N_12858,N_12070,N_12276);
nor U12859 (N_12859,N_12331,N_12223);
and U12860 (N_12860,N_12481,N_12352);
nand U12861 (N_12861,N_12180,N_12382);
xnor U12862 (N_12862,N_12180,N_12030);
nor U12863 (N_12863,N_12265,N_12499);
and U12864 (N_12864,N_12345,N_12262);
and U12865 (N_12865,N_12056,N_12261);
xnor U12866 (N_12866,N_12218,N_12448);
or U12867 (N_12867,N_12100,N_12494);
and U12868 (N_12868,N_12474,N_12015);
and U12869 (N_12869,N_12389,N_12445);
or U12870 (N_12870,N_12008,N_12471);
or U12871 (N_12871,N_12158,N_12028);
xor U12872 (N_12872,N_12119,N_12420);
or U12873 (N_12873,N_12071,N_12462);
nand U12874 (N_12874,N_12108,N_12064);
and U12875 (N_12875,N_12303,N_12405);
nand U12876 (N_12876,N_12083,N_12104);
nor U12877 (N_12877,N_12422,N_12343);
nand U12878 (N_12878,N_12007,N_12458);
and U12879 (N_12879,N_12323,N_12039);
or U12880 (N_12880,N_12032,N_12376);
or U12881 (N_12881,N_12241,N_12490);
xor U12882 (N_12882,N_12323,N_12220);
nand U12883 (N_12883,N_12130,N_12238);
xor U12884 (N_12884,N_12467,N_12021);
nor U12885 (N_12885,N_12434,N_12174);
xnor U12886 (N_12886,N_12268,N_12092);
nand U12887 (N_12887,N_12034,N_12175);
nand U12888 (N_12888,N_12267,N_12240);
nand U12889 (N_12889,N_12161,N_12180);
nand U12890 (N_12890,N_12150,N_12178);
nor U12891 (N_12891,N_12265,N_12496);
and U12892 (N_12892,N_12300,N_12131);
xnor U12893 (N_12893,N_12338,N_12020);
nor U12894 (N_12894,N_12488,N_12234);
xnor U12895 (N_12895,N_12216,N_12424);
and U12896 (N_12896,N_12193,N_12329);
nand U12897 (N_12897,N_12218,N_12064);
and U12898 (N_12898,N_12267,N_12152);
or U12899 (N_12899,N_12038,N_12291);
nor U12900 (N_12900,N_12380,N_12017);
nand U12901 (N_12901,N_12369,N_12435);
and U12902 (N_12902,N_12255,N_12286);
nor U12903 (N_12903,N_12290,N_12144);
nor U12904 (N_12904,N_12213,N_12497);
and U12905 (N_12905,N_12111,N_12245);
or U12906 (N_12906,N_12050,N_12375);
or U12907 (N_12907,N_12425,N_12334);
or U12908 (N_12908,N_12232,N_12228);
or U12909 (N_12909,N_12135,N_12066);
or U12910 (N_12910,N_12136,N_12223);
nand U12911 (N_12911,N_12293,N_12221);
nor U12912 (N_12912,N_12066,N_12355);
xnor U12913 (N_12913,N_12357,N_12326);
xor U12914 (N_12914,N_12283,N_12011);
or U12915 (N_12915,N_12452,N_12482);
or U12916 (N_12916,N_12012,N_12130);
and U12917 (N_12917,N_12202,N_12035);
nor U12918 (N_12918,N_12268,N_12216);
or U12919 (N_12919,N_12451,N_12068);
or U12920 (N_12920,N_12205,N_12400);
xor U12921 (N_12921,N_12291,N_12323);
nor U12922 (N_12922,N_12362,N_12463);
and U12923 (N_12923,N_12411,N_12201);
nor U12924 (N_12924,N_12368,N_12261);
xnor U12925 (N_12925,N_12419,N_12331);
or U12926 (N_12926,N_12156,N_12323);
or U12927 (N_12927,N_12193,N_12246);
xnor U12928 (N_12928,N_12268,N_12094);
xor U12929 (N_12929,N_12046,N_12041);
and U12930 (N_12930,N_12446,N_12161);
xor U12931 (N_12931,N_12179,N_12247);
or U12932 (N_12932,N_12202,N_12414);
nand U12933 (N_12933,N_12260,N_12376);
nand U12934 (N_12934,N_12008,N_12013);
and U12935 (N_12935,N_12401,N_12023);
xor U12936 (N_12936,N_12167,N_12473);
xnor U12937 (N_12937,N_12190,N_12192);
xnor U12938 (N_12938,N_12069,N_12430);
nand U12939 (N_12939,N_12444,N_12092);
and U12940 (N_12940,N_12494,N_12316);
nand U12941 (N_12941,N_12348,N_12356);
xor U12942 (N_12942,N_12023,N_12274);
xnor U12943 (N_12943,N_12044,N_12147);
xor U12944 (N_12944,N_12423,N_12246);
or U12945 (N_12945,N_12491,N_12259);
xnor U12946 (N_12946,N_12434,N_12201);
nand U12947 (N_12947,N_12091,N_12149);
nor U12948 (N_12948,N_12422,N_12008);
and U12949 (N_12949,N_12023,N_12219);
nor U12950 (N_12950,N_12218,N_12484);
xnor U12951 (N_12951,N_12038,N_12343);
nand U12952 (N_12952,N_12293,N_12253);
and U12953 (N_12953,N_12266,N_12201);
xor U12954 (N_12954,N_12329,N_12370);
xnor U12955 (N_12955,N_12047,N_12053);
nor U12956 (N_12956,N_12370,N_12461);
nand U12957 (N_12957,N_12153,N_12091);
xor U12958 (N_12958,N_12015,N_12324);
or U12959 (N_12959,N_12307,N_12121);
or U12960 (N_12960,N_12426,N_12465);
xor U12961 (N_12961,N_12150,N_12181);
nand U12962 (N_12962,N_12232,N_12191);
nand U12963 (N_12963,N_12388,N_12475);
xor U12964 (N_12964,N_12105,N_12386);
nand U12965 (N_12965,N_12483,N_12222);
nor U12966 (N_12966,N_12462,N_12474);
or U12967 (N_12967,N_12225,N_12487);
xnor U12968 (N_12968,N_12251,N_12491);
xnor U12969 (N_12969,N_12078,N_12357);
or U12970 (N_12970,N_12267,N_12029);
or U12971 (N_12971,N_12477,N_12227);
nand U12972 (N_12972,N_12002,N_12161);
nand U12973 (N_12973,N_12004,N_12464);
or U12974 (N_12974,N_12190,N_12208);
nand U12975 (N_12975,N_12221,N_12217);
or U12976 (N_12976,N_12099,N_12341);
nor U12977 (N_12977,N_12179,N_12454);
nor U12978 (N_12978,N_12237,N_12137);
xnor U12979 (N_12979,N_12233,N_12090);
and U12980 (N_12980,N_12450,N_12096);
xor U12981 (N_12981,N_12190,N_12194);
nand U12982 (N_12982,N_12058,N_12075);
and U12983 (N_12983,N_12294,N_12217);
and U12984 (N_12984,N_12082,N_12452);
xor U12985 (N_12985,N_12479,N_12000);
and U12986 (N_12986,N_12008,N_12419);
or U12987 (N_12987,N_12191,N_12157);
xnor U12988 (N_12988,N_12000,N_12465);
nand U12989 (N_12989,N_12489,N_12343);
nor U12990 (N_12990,N_12106,N_12208);
or U12991 (N_12991,N_12341,N_12452);
or U12992 (N_12992,N_12024,N_12074);
nor U12993 (N_12993,N_12412,N_12336);
and U12994 (N_12994,N_12476,N_12236);
and U12995 (N_12995,N_12406,N_12091);
nor U12996 (N_12996,N_12100,N_12390);
or U12997 (N_12997,N_12194,N_12207);
or U12998 (N_12998,N_12376,N_12190);
xor U12999 (N_12999,N_12014,N_12163);
or U13000 (N_13000,N_12854,N_12727);
and U13001 (N_13001,N_12524,N_12826);
and U13002 (N_13002,N_12614,N_12970);
and U13003 (N_13003,N_12540,N_12682);
and U13004 (N_13004,N_12937,N_12581);
nand U13005 (N_13005,N_12534,N_12747);
nand U13006 (N_13006,N_12945,N_12926);
nand U13007 (N_13007,N_12652,N_12579);
and U13008 (N_13008,N_12716,N_12967);
nor U13009 (N_13009,N_12944,N_12882);
or U13010 (N_13010,N_12809,N_12609);
and U13011 (N_13011,N_12521,N_12756);
or U13012 (N_13012,N_12653,N_12822);
or U13013 (N_13013,N_12684,N_12541);
or U13014 (N_13014,N_12845,N_12896);
nand U13015 (N_13015,N_12743,N_12794);
or U13016 (N_13016,N_12879,N_12580);
or U13017 (N_13017,N_12648,N_12764);
and U13018 (N_13018,N_12948,N_12694);
nor U13019 (N_13019,N_12889,N_12615);
nor U13020 (N_13020,N_12739,N_12770);
and U13021 (N_13021,N_12563,N_12760);
or U13022 (N_13022,N_12925,N_12874);
nand U13023 (N_13023,N_12998,N_12832);
nand U13024 (N_13024,N_12724,N_12641);
nand U13025 (N_13025,N_12976,N_12938);
xor U13026 (N_13026,N_12550,N_12960);
nand U13027 (N_13027,N_12836,N_12806);
nand U13028 (N_13028,N_12628,N_12509);
nor U13029 (N_13029,N_12588,N_12936);
xor U13030 (N_13030,N_12557,N_12574);
or U13031 (N_13031,N_12840,N_12767);
nand U13032 (N_13032,N_12920,N_12860);
nand U13033 (N_13033,N_12867,N_12545);
xor U13034 (N_13034,N_12754,N_12971);
nor U13035 (N_13035,N_12635,N_12798);
or U13036 (N_13036,N_12714,N_12984);
nand U13037 (N_13037,N_12622,N_12911);
xnor U13038 (N_13038,N_12607,N_12780);
xor U13039 (N_13039,N_12923,N_12632);
or U13040 (N_13040,N_12807,N_12931);
xnor U13041 (N_13041,N_12691,N_12616);
and U13042 (N_13042,N_12802,N_12745);
and U13043 (N_13043,N_12858,N_12873);
nand U13044 (N_13044,N_12603,N_12582);
or U13045 (N_13045,N_12748,N_12916);
nor U13046 (N_13046,N_12728,N_12823);
nand U13047 (N_13047,N_12990,N_12543);
or U13048 (N_13048,N_12980,N_12850);
and U13049 (N_13049,N_12642,N_12585);
or U13050 (N_13050,N_12940,N_12846);
and U13051 (N_13051,N_12902,N_12988);
and U13052 (N_13052,N_12819,N_12611);
nand U13053 (N_13053,N_12932,N_12561);
xor U13054 (N_13054,N_12839,N_12878);
or U13055 (N_13055,N_12578,N_12784);
or U13056 (N_13056,N_12966,N_12590);
nand U13057 (N_13057,N_12949,N_12863);
nor U13058 (N_13058,N_12700,N_12710);
and U13059 (N_13059,N_12569,N_12892);
or U13060 (N_13060,N_12505,N_12522);
or U13061 (N_13061,N_12801,N_12978);
xnor U13062 (N_13062,N_12644,N_12538);
nor U13063 (N_13063,N_12888,N_12929);
and U13064 (N_13064,N_12816,N_12564);
nand U13065 (N_13065,N_12856,N_12908);
nand U13066 (N_13066,N_12898,N_12752);
xnor U13067 (N_13067,N_12958,N_12987);
and U13068 (N_13068,N_12847,N_12577);
nand U13069 (N_13069,N_12876,N_12708);
and U13070 (N_13070,N_12733,N_12812);
and U13071 (N_13071,N_12514,N_12587);
or U13072 (N_13072,N_12963,N_12969);
xnor U13073 (N_13073,N_12877,N_12654);
or U13074 (N_13074,N_12986,N_12893);
and U13075 (N_13075,N_12713,N_12705);
nor U13076 (N_13076,N_12551,N_12595);
xor U13077 (N_13077,N_12928,N_12720);
nor U13078 (N_13078,N_12885,N_12501);
or U13079 (N_13079,N_12518,N_12679);
xor U13080 (N_13080,N_12975,N_12701);
nor U13081 (N_13081,N_12688,N_12608);
and U13082 (N_13082,N_12934,N_12573);
nor U13083 (N_13083,N_12983,N_12895);
nor U13084 (N_13084,N_12690,N_12755);
and U13085 (N_13085,N_12567,N_12526);
nor U13086 (N_13086,N_12849,N_12951);
nor U13087 (N_13087,N_12829,N_12516);
or U13088 (N_13088,N_12736,N_12602);
nor U13089 (N_13089,N_12670,N_12558);
nand U13090 (N_13090,N_12537,N_12974);
xnor U13091 (N_13091,N_12552,N_12500);
or U13092 (N_13092,N_12848,N_12715);
nor U13093 (N_13093,N_12637,N_12775);
nor U13094 (N_13094,N_12942,N_12852);
or U13095 (N_13095,N_12766,N_12671);
nor U13096 (N_13096,N_12726,N_12999);
and U13097 (N_13097,N_12553,N_12589);
nand U13098 (N_13098,N_12805,N_12697);
or U13099 (N_13099,N_12681,N_12592);
nand U13100 (N_13100,N_12687,N_12881);
nor U13101 (N_13101,N_12827,N_12719);
and U13102 (N_13102,N_12831,N_12717);
nor U13103 (N_13103,N_12952,N_12953);
xor U13104 (N_13104,N_12572,N_12771);
and U13105 (N_13105,N_12869,N_12957);
xnor U13106 (N_13106,N_12907,N_12744);
nor U13107 (N_13107,N_12870,N_12525);
or U13108 (N_13108,N_12502,N_12663);
nand U13109 (N_13109,N_12964,N_12790);
or U13110 (N_13110,N_12946,N_12555);
nand U13111 (N_13111,N_12650,N_12512);
xor U13112 (N_13112,N_12620,N_12955);
and U13113 (N_13113,N_12818,N_12520);
xnor U13114 (N_13114,N_12596,N_12666);
or U13115 (N_13115,N_12735,N_12627);
xor U13116 (N_13116,N_12712,N_12914);
and U13117 (N_13117,N_12789,N_12785);
or U13118 (N_13118,N_12751,N_12664);
xor U13119 (N_13119,N_12662,N_12732);
nor U13120 (N_13120,N_12842,N_12997);
nand U13121 (N_13121,N_12773,N_12610);
nor U13122 (N_13122,N_12597,N_12950);
nor U13123 (N_13123,N_12549,N_12750);
nor U13124 (N_13124,N_12741,N_12706);
nor U13125 (N_13125,N_12880,N_12927);
nand U13126 (N_13126,N_12939,N_12919);
and U13127 (N_13127,N_12542,N_12638);
or U13128 (N_13128,N_12841,N_12566);
nor U13129 (N_13129,N_12527,N_12834);
xnor U13130 (N_13130,N_12676,N_12556);
or U13131 (N_13131,N_12782,N_12612);
xnor U13132 (N_13132,N_12899,N_12658);
or U13133 (N_13133,N_12996,N_12593);
or U13134 (N_13134,N_12859,N_12630);
xor U13135 (N_13135,N_12804,N_12740);
and U13136 (N_13136,N_12776,N_12544);
nand U13137 (N_13137,N_12995,N_12718);
xnor U13138 (N_13138,N_12890,N_12699);
and U13139 (N_13139,N_12901,N_12667);
nor U13140 (N_13140,N_12972,N_12956);
nand U13141 (N_13141,N_12821,N_12924);
nor U13142 (N_13142,N_12973,N_12698);
xor U13143 (N_13143,N_12598,N_12977);
and U13144 (N_13144,N_12692,N_12979);
or U13145 (N_13145,N_12617,N_12606);
and U13146 (N_13146,N_12918,N_12904);
and U13147 (N_13147,N_12721,N_12817);
and U13148 (N_13148,N_12626,N_12959);
xnor U13149 (N_13149,N_12825,N_12601);
nand U13150 (N_13150,N_12772,N_12643);
or U13151 (N_13151,N_12591,N_12695);
or U13152 (N_13152,N_12729,N_12922);
xor U13153 (N_13153,N_12660,N_12930);
nand U13154 (N_13154,N_12562,N_12613);
or U13155 (N_13155,N_12962,N_12799);
or U13156 (N_13156,N_12680,N_12599);
nand U13157 (N_13157,N_12504,N_12909);
and U13158 (N_13158,N_12851,N_12730);
or U13159 (N_13159,N_12709,N_12533);
xor U13160 (N_13160,N_12765,N_12968);
nand U13161 (N_13161,N_12810,N_12529);
or U13162 (N_13162,N_12689,N_12570);
xnor U13163 (N_13163,N_12887,N_12649);
or U13164 (N_13164,N_12894,N_12864);
nand U13165 (N_13165,N_12528,N_12758);
xor U13166 (N_13166,N_12665,N_12795);
and U13167 (N_13167,N_12933,N_12546);
and U13168 (N_13168,N_12875,N_12655);
and U13169 (N_13169,N_12943,N_12631);
nor U13170 (N_13170,N_12742,N_12903);
or U13171 (N_13171,N_12530,N_12539);
xor U13172 (N_13172,N_12668,N_12575);
xnor U13173 (N_13173,N_12624,N_12868);
xnor U13174 (N_13174,N_12523,N_12757);
xnor U13175 (N_13175,N_12947,N_12559);
nand U13176 (N_13176,N_12814,N_12835);
nand U13177 (N_13177,N_12781,N_12915);
nand U13178 (N_13178,N_12905,N_12672);
and U13179 (N_13179,N_12731,N_12656);
nor U13180 (N_13180,N_12503,N_12853);
nor U13181 (N_13181,N_12838,N_12866);
xor U13182 (N_13182,N_12686,N_12833);
or U13183 (N_13183,N_12511,N_12723);
nand U13184 (N_13184,N_12912,N_12640);
nand U13185 (N_13185,N_12633,N_12808);
or U13186 (N_13186,N_12862,N_12722);
and U13187 (N_13187,N_12634,N_12800);
nand U13188 (N_13188,N_12855,N_12657);
or U13189 (N_13189,N_12636,N_12759);
nor U13190 (N_13190,N_12793,N_12677);
nor U13191 (N_13191,N_12571,N_12796);
and U13192 (N_13192,N_12777,N_12820);
or U13193 (N_13193,N_12913,N_12897);
xnor U13194 (N_13194,N_12583,N_12508);
or U13195 (N_13195,N_12917,N_12515);
xnor U13196 (N_13196,N_12576,N_12813);
xnor U13197 (N_13197,N_12623,N_12992);
and U13198 (N_13198,N_12778,N_12749);
nor U13199 (N_13199,N_12910,N_12683);
and U13200 (N_13200,N_12769,N_12678);
xor U13201 (N_13201,N_12815,N_12661);
xor U13202 (N_13202,N_12872,N_12535);
nor U13203 (N_13203,N_12941,N_12738);
nor U13204 (N_13204,N_12803,N_12685);
nor U13205 (N_13205,N_12547,N_12675);
or U13206 (N_13206,N_12843,N_12991);
nor U13207 (N_13207,N_12761,N_12961);
and U13208 (N_13208,N_12993,N_12981);
and U13209 (N_13209,N_12768,N_12763);
nor U13210 (N_13210,N_12548,N_12513);
and U13211 (N_13211,N_12792,N_12629);
xnor U13212 (N_13212,N_12506,N_12703);
xnor U13213 (N_13213,N_12600,N_12619);
and U13214 (N_13214,N_12965,N_12783);
xor U13215 (N_13215,N_12532,N_12791);
xnor U13216 (N_13216,N_12921,N_12737);
xor U13217 (N_13217,N_12646,N_12647);
and U13218 (N_13218,N_12510,N_12886);
and U13219 (N_13219,N_12669,N_12568);
xnor U13220 (N_13220,N_12797,N_12884);
xor U13221 (N_13221,N_12746,N_12985);
xor U13222 (N_13222,N_12954,N_12711);
or U13223 (N_13223,N_12519,N_12674);
nand U13224 (N_13224,N_12762,N_12734);
nor U13225 (N_13225,N_12517,N_12645);
xnor U13226 (N_13226,N_12865,N_12704);
nand U13227 (N_13227,N_12693,N_12618);
xor U13228 (N_13228,N_12786,N_12621);
and U13229 (N_13229,N_12586,N_12707);
nand U13230 (N_13230,N_12702,N_12560);
or U13231 (N_13231,N_12625,N_12774);
or U13232 (N_13232,N_12696,N_12753);
xor U13233 (N_13233,N_12659,N_12788);
or U13234 (N_13234,N_12906,N_12565);
nor U13235 (N_13235,N_12507,N_12935);
xor U13236 (N_13236,N_12830,N_12651);
xor U13237 (N_13237,N_12787,N_12824);
xnor U13238 (N_13238,N_12994,N_12837);
or U13239 (N_13239,N_12871,N_12594);
xnor U13240 (N_13240,N_12861,N_12844);
nor U13241 (N_13241,N_12900,N_12605);
xnor U13242 (N_13242,N_12531,N_12828);
nor U13243 (N_13243,N_12982,N_12725);
nor U13244 (N_13244,N_12604,N_12554);
nand U13245 (N_13245,N_12584,N_12989);
or U13246 (N_13246,N_12891,N_12536);
nand U13247 (N_13247,N_12883,N_12779);
xnor U13248 (N_13248,N_12673,N_12811);
and U13249 (N_13249,N_12857,N_12639);
or U13250 (N_13250,N_12505,N_12650);
or U13251 (N_13251,N_12931,N_12969);
or U13252 (N_13252,N_12711,N_12615);
nand U13253 (N_13253,N_12602,N_12915);
xnor U13254 (N_13254,N_12825,N_12609);
nand U13255 (N_13255,N_12553,N_12786);
or U13256 (N_13256,N_12939,N_12531);
nand U13257 (N_13257,N_12997,N_12858);
or U13258 (N_13258,N_12986,N_12575);
or U13259 (N_13259,N_12984,N_12816);
nor U13260 (N_13260,N_12526,N_12644);
nor U13261 (N_13261,N_12935,N_12983);
or U13262 (N_13262,N_12631,N_12930);
and U13263 (N_13263,N_12732,N_12538);
and U13264 (N_13264,N_12779,N_12830);
nand U13265 (N_13265,N_12595,N_12524);
xor U13266 (N_13266,N_12982,N_12621);
nand U13267 (N_13267,N_12641,N_12757);
nand U13268 (N_13268,N_12858,N_12952);
nand U13269 (N_13269,N_12864,N_12821);
nand U13270 (N_13270,N_12933,N_12841);
nor U13271 (N_13271,N_12554,N_12898);
nand U13272 (N_13272,N_12695,N_12810);
nand U13273 (N_13273,N_12710,N_12598);
and U13274 (N_13274,N_12653,N_12901);
or U13275 (N_13275,N_12726,N_12793);
xnor U13276 (N_13276,N_12763,N_12847);
and U13277 (N_13277,N_12770,N_12930);
and U13278 (N_13278,N_12649,N_12805);
nor U13279 (N_13279,N_12903,N_12635);
nor U13280 (N_13280,N_12531,N_12566);
xnor U13281 (N_13281,N_12952,N_12722);
or U13282 (N_13282,N_12523,N_12931);
nand U13283 (N_13283,N_12620,N_12877);
or U13284 (N_13284,N_12941,N_12749);
or U13285 (N_13285,N_12522,N_12882);
or U13286 (N_13286,N_12725,N_12744);
nand U13287 (N_13287,N_12569,N_12869);
nor U13288 (N_13288,N_12629,N_12590);
nor U13289 (N_13289,N_12923,N_12866);
nor U13290 (N_13290,N_12931,N_12923);
nor U13291 (N_13291,N_12563,N_12898);
nor U13292 (N_13292,N_12552,N_12890);
and U13293 (N_13293,N_12817,N_12685);
nand U13294 (N_13294,N_12656,N_12923);
nand U13295 (N_13295,N_12517,N_12582);
xnor U13296 (N_13296,N_12682,N_12725);
nand U13297 (N_13297,N_12554,N_12546);
or U13298 (N_13298,N_12685,N_12717);
xor U13299 (N_13299,N_12938,N_12994);
xnor U13300 (N_13300,N_12670,N_12933);
or U13301 (N_13301,N_12578,N_12601);
nand U13302 (N_13302,N_12881,N_12565);
and U13303 (N_13303,N_12653,N_12613);
nor U13304 (N_13304,N_12512,N_12542);
xor U13305 (N_13305,N_12726,N_12734);
nor U13306 (N_13306,N_12514,N_12848);
nand U13307 (N_13307,N_12909,N_12741);
and U13308 (N_13308,N_12921,N_12519);
or U13309 (N_13309,N_12669,N_12644);
or U13310 (N_13310,N_12959,N_12995);
or U13311 (N_13311,N_12603,N_12867);
and U13312 (N_13312,N_12730,N_12829);
and U13313 (N_13313,N_12510,N_12621);
nor U13314 (N_13314,N_12835,N_12821);
xor U13315 (N_13315,N_12745,N_12894);
or U13316 (N_13316,N_12815,N_12615);
nor U13317 (N_13317,N_12767,N_12633);
nand U13318 (N_13318,N_12551,N_12519);
xor U13319 (N_13319,N_12897,N_12579);
and U13320 (N_13320,N_12930,N_12678);
nor U13321 (N_13321,N_12969,N_12986);
nor U13322 (N_13322,N_12635,N_12568);
nand U13323 (N_13323,N_12919,N_12582);
and U13324 (N_13324,N_12945,N_12573);
xor U13325 (N_13325,N_12998,N_12592);
nand U13326 (N_13326,N_12665,N_12906);
nor U13327 (N_13327,N_12567,N_12663);
and U13328 (N_13328,N_12502,N_12795);
or U13329 (N_13329,N_12633,N_12895);
or U13330 (N_13330,N_12727,N_12969);
or U13331 (N_13331,N_12567,N_12806);
xor U13332 (N_13332,N_12540,N_12987);
and U13333 (N_13333,N_12798,N_12762);
nand U13334 (N_13334,N_12819,N_12636);
xnor U13335 (N_13335,N_12555,N_12687);
or U13336 (N_13336,N_12521,N_12727);
nand U13337 (N_13337,N_12868,N_12880);
and U13338 (N_13338,N_12631,N_12528);
xor U13339 (N_13339,N_12538,N_12930);
nand U13340 (N_13340,N_12617,N_12584);
nor U13341 (N_13341,N_12992,N_12641);
xnor U13342 (N_13342,N_12770,N_12702);
or U13343 (N_13343,N_12548,N_12514);
nand U13344 (N_13344,N_12688,N_12894);
or U13345 (N_13345,N_12975,N_12753);
nor U13346 (N_13346,N_12705,N_12807);
nand U13347 (N_13347,N_12774,N_12699);
and U13348 (N_13348,N_12567,N_12659);
nor U13349 (N_13349,N_12516,N_12982);
and U13350 (N_13350,N_12576,N_12957);
nand U13351 (N_13351,N_12982,N_12672);
nand U13352 (N_13352,N_12765,N_12976);
nor U13353 (N_13353,N_12868,N_12954);
and U13354 (N_13354,N_12906,N_12957);
nor U13355 (N_13355,N_12694,N_12906);
xor U13356 (N_13356,N_12995,N_12763);
and U13357 (N_13357,N_12874,N_12632);
nor U13358 (N_13358,N_12948,N_12902);
nand U13359 (N_13359,N_12824,N_12997);
and U13360 (N_13360,N_12614,N_12620);
xnor U13361 (N_13361,N_12773,N_12890);
or U13362 (N_13362,N_12686,N_12632);
or U13363 (N_13363,N_12632,N_12671);
and U13364 (N_13364,N_12865,N_12738);
nor U13365 (N_13365,N_12904,N_12552);
xor U13366 (N_13366,N_12509,N_12711);
and U13367 (N_13367,N_12714,N_12772);
and U13368 (N_13368,N_12923,N_12949);
or U13369 (N_13369,N_12996,N_12814);
nor U13370 (N_13370,N_12755,N_12597);
nand U13371 (N_13371,N_12944,N_12789);
or U13372 (N_13372,N_12930,N_12995);
nand U13373 (N_13373,N_12940,N_12946);
and U13374 (N_13374,N_12711,N_12769);
xor U13375 (N_13375,N_12577,N_12567);
nor U13376 (N_13376,N_12556,N_12542);
xnor U13377 (N_13377,N_12529,N_12725);
nor U13378 (N_13378,N_12542,N_12912);
and U13379 (N_13379,N_12652,N_12609);
or U13380 (N_13380,N_12624,N_12974);
and U13381 (N_13381,N_12881,N_12798);
nor U13382 (N_13382,N_12800,N_12783);
or U13383 (N_13383,N_12946,N_12682);
xor U13384 (N_13384,N_12890,N_12918);
xnor U13385 (N_13385,N_12513,N_12881);
or U13386 (N_13386,N_12631,N_12850);
xor U13387 (N_13387,N_12930,N_12519);
and U13388 (N_13388,N_12976,N_12742);
nor U13389 (N_13389,N_12757,N_12976);
nor U13390 (N_13390,N_12603,N_12829);
nor U13391 (N_13391,N_12974,N_12881);
and U13392 (N_13392,N_12947,N_12906);
nor U13393 (N_13393,N_12533,N_12811);
nand U13394 (N_13394,N_12513,N_12912);
nor U13395 (N_13395,N_12744,N_12568);
nand U13396 (N_13396,N_12933,N_12818);
xnor U13397 (N_13397,N_12643,N_12979);
xor U13398 (N_13398,N_12840,N_12950);
and U13399 (N_13399,N_12982,N_12786);
or U13400 (N_13400,N_12810,N_12593);
or U13401 (N_13401,N_12958,N_12719);
and U13402 (N_13402,N_12763,N_12738);
nor U13403 (N_13403,N_12614,N_12980);
xor U13404 (N_13404,N_12622,N_12941);
or U13405 (N_13405,N_12879,N_12824);
nor U13406 (N_13406,N_12909,N_12652);
or U13407 (N_13407,N_12507,N_12603);
nor U13408 (N_13408,N_12798,N_12550);
or U13409 (N_13409,N_12582,N_12839);
and U13410 (N_13410,N_12686,N_12758);
and U13411 (N_13411,N_12992,N_12511);
or U13412 (N_13412,N_12597,N_12622);
or U13413 (N_13413,N_12586,N_12549);
or U13414 (N_13414,N_12619,N_12593);
and U13415 (N_13415,N_12943,N_12993);
and U13416 (N_13416,N_12726,N_12914);
xnor U13417 (N_13417,N_12911,N_12726);
nor U13418 (N_13418,N_12652,N_12713);
nand U13419 (N_13419,N_12579,N_12603);
xnor U13420 (N_13420,N_12968,N_12735);
nand U13421 (N_13421,N_12829,N_12681);
nor U13422 (N_13422,N_12881,N_12699);
and U13423 (N_13423,N_12698,N_12934);
xnor U13424 (N_13424,N_12964,N_12624);
xnor U13425 (N_13425,N_12837,N_12757);
nor U13426 (N_13426,N_12597,N_12523);
xor U13427 (N_13427,N_12831,N_12926);
xnor U13428 (N_13428,N_12686,N_12780);
nor U13429 (N_13429,N_12838,N_12929);
xor U13430 (N_13430,N_12865,N_12871);
or U13431 (N_13431,N_12544,N_12997);
xor U13432 (N_13432,N_12701,N_12507);
nand U13433 (N_13433,N_12784,N_12529);
xor U13434 (N_13434,N_12642,N_12768);
xor U13435 (N_13435,N_12929,N_12526);
nor U13436 (N_13436,N_12779,N_12600);
nor U13437 (N_13437,N_12728,N_12500);
xor U13438 (N_13438,N_12702,N_12548);
or U13439 (N_13439,N_12916,N_12719);
xnor U13440 (N_13440,N_12801,N_12673);
and U13441 (N_13441,N_12666,N_12880);
xor U13442 (N_13442,N_12788,N_12745);
and U13443 (N_13443,N_12876,N_12994);
nand U13444 (N_13444,N_12772,N_12771);
nand U13445 (N_13445,N_12507,N_12964);
nor U13446 (N_13446,N_12642,N_12865);
nand U13447 (N_13447,N_12611,N_12650);
and U13448 (N_13448,N_12894,N_12785);
nand U13449 (N_13449,N_12675,N_12596);
xor U13450 (N_13450,N_12742,N_12996);
or U13451 (N_13451,N_12679,N_12984);
and U13452 (N_13452,N_12844,N_12583);
nor U13453 (N_13453,N_12925,N_12653);
nor U13454 (N_13454,N_12872,N_12726);
nor U13455 (N_13455,N_12860,N_12854);
nand U13456 (N_13456,N_12893,N_12846);
and U13457 (N_13457,N_12539,N_12802);
xnor U13458 (N_13458,N_12643,N_12621);
and U13459 (N_13459,N_12571,N_12504);
or U13460 (N_13460,N_12804,N_12986);
nand U13461 (N_13461,N_12988,N_12810);
xor U13462 (N_13462,N_12725,N_12955);
and U13463 (N_13463,N_12872,N_12837);
and U13464 (N_13464,N_12974,N_12566);
nand U13465 (N_13465,N_12507,N_12669);
nor U13466 (N_13466,N_12795,N_12746);
xor U13467 (N_13467,N_12968,N_12884);
and U13468 (N_13468,N_12611,N_12784);
nor U13469 (N_13469,N_12650,N_12977);
nand U13470 (N_13470,N_12704,N_12681);
xnor U13471 (N_13471,N_12839,N_12835);
xnor U13472 (N_13472,N_12725,N_12690);
nand U13473 (N_13473,N_12866,N_12517);
and U13474 (N_13474,N_12794,N_12845);
or U13475 (N_13475,N_12887,N_12844);
or U13476 (N_13476,N_12635,N_12865);
or U13477 (N_13477,N_12851,N_12983);
nor U13478 (N_13478,N_12996,N_12610);
nand U13479 (N_13479,N_12756,N_12984);
or U13480 (N_13480,N_12539,N_12833);
nand U13481 (N_13481,N_12709,N_12664);
nor U13482 (N_13482,N_12641,N_12668);
nor U13483 (N_13483,N_12773,N_12782);
xor U13484 (N_13484,N_12885,N_12814);
xnor U13485 (N_13485,N_12570,N_12900);
and U13486 (N_13486,N_12512,N_12649);
and U13487 (N_13487,N_12821,N_12609);
or U13488 (N_13488,N_12677,N_12532);
nor U13489 (N_13489,N_12924,N_12647);
nand U13490 (N_13490,N_12678,N_12952);
or U13491 (N_13491,N_12684,N_12534);
nor U13492 (N_13492,N_12709,N_12565);
xnor U13493 (N_13493,N_12518,N_12620);
nor U13494 (N_13494,N_12588,N_12539);
nor U13495 (N_13495,N_12592,N_12590);
nor U13496 (N_13496,N_12699,N_12613);
and U13497 (N_13497,N_12998,N_12974);
or U13498 (N_13498,N_12713,N_12775);
or U13499 (N_13499,N_12530,N_12560);
and U13500 (N_13500,N_13180,N_13206);
xnor U13501 (N_13501,N_13380,N_13412);
and U13502 (N_13502,N_13210,N_13216);
xor U13503 (N_13503,N_13125,N_13014);
nand U13504 (N_13504,N_13346,N_13266);
or U13505 (N_13505,N_13110,N_13005);
nor U13506 (N_13506,N_13384,N_13421);
or U13507 (N_13507,N_13133,N_13079);
nand U13508 (N_13508,N_13259,N_13068);
xor U13509 (N_13509,N_13186,N_13177);
nor U13510 (N_13510,N_13343,N_13003);
or U13511 (N_13511,N_13132,N_13127);
nor U13512 (N_13512,N_13417,N_13371);
nand U13513 (N_13513,N_13398,N_13195);
nand U13514 (N_13514,N_13016,N_13205);
or U13515 (N_13515,N_13162,N_13355);
nor U13516 (N_13516,N_13023,N_13336);
and U13517 (N_13517,N_13374,N_13252);
and U13518 (N_13518,N_13303,N_13238);
and U13519 (N_13519,N_13328,N_13473);
and U13520 (N_13520,N_13159,N_13296);
nor U13521 (N_13521,N_13078,N_13393);
xor U13522 (N_13522,N_13489,N_13203);
or U13523 (N_13523,N_13100,N_13348);
xnor U13524 (N_13524,N_13308,N_13474);
nor U13525 (N_13525,N_13418,N_13283);
or U13526 (N_13526,N_13265,N_13332);
nor U13527 (N_13527,N_13490,N_13425);
or U13528 (N_13528,N_13179,N_13157);
nand U13529 (N_13529,N_13229,N_13001);
nand U13530 (N_13530,N_13315,N_13470);
or U13531 (N_13531,N_13258,N_13431);
xnor U13532 (N_13532,N_13277,N_13046);
and U13533 (N_13533,N_13423,N_13092);
xor U13534 (N_13534,N_13300,N_13434);
xor U13535 (N_13535,N_13217,N_13399);
and U13536 (N_13536,N_13268,N_13056);
xor U13537 (N_13537,N_13144,N_13072);
nand U13538 (N_13538,N_13174,N_13230);
nand U13539 (N_13539,N_13040,N_13207);
or U13540 (N_13540,N_13166,N_13290);
nor U13541 (N_13541,N_13089,N_13349);
xnor U13542 (N_13542,N_13242,N_13435);
or U13543 (N_13543,N_13262,N_13221);
nand U13544 (N_13544,N_13376,N_13225);
nand U13545 (N_13545,N_13416,N_13467);
or U13546 (N_13546,N_13015,N_13134);
and U13547 (N_13547,N_13481,N_13136);
or U13548 (N_13548,N_13447,N_13152);
and U13549 (N_13549,N_13008,N_13156);
nand U13550 (N_13550,N_13382,N_13451);
and U13551 (N_13551,N_13345,N_13298);
or U13552 (N_13552,N_13269,N_13281);
xnor U13553 (N_13553,N_13459,N_13471);
nor U13554 (N_13554,N_13226,N_13139);
or U13555 (N_13555,N_13084,N_13487);
xor U13556 (N_13556,N_13063,N_13352);
xnor U13557 (N_13557,N_13436,N_13301);
nand U13558 (N_13558,N_13129,N_13083);
nand U13559 (N_13559,N_13131,N_13038);
and U13560 (N_13560,N_13227,N_13271);
nand U13561 (N_13561,N_13429,N_13354);
nand U13562 (N_13562,N_13275,N_13458);
or U13563 (N_13563,N_13051,N_13394);
nand U13564 (N_13564,N_13383,N_13415);
nor U13565 (N_13565,N_13342,N_13304);
and U13566 (N_13566,N_13197,N_13094);
xor U13567 (N_13567,N_13276,N_13433);
and U13568 (N_13568,N_13414,N_13239);
or U13569 (N_13569,N_13189,N_13147);
nand U13570 (N_13570,N_13082,N_13396);
and U13571 (N_13571,N_13172,N_13466);
or U13572 (N_13572,N_13282,N_13309);
or U13573 (N_13573,N_13360,N_13462);
xnor U13574 (N_13574,N_13333,N_13143);
xnor U13575 (N_13575,N_13187,N_13020);
nor U13576 (N_13576,N_13455,N_13220);
nor U13577 (N_13577,N_13101,N_13438);
and U13578 (N_13578,N_13019,N_13310);
xnor U13579 (N_13579,N_13256,N_13363);
nor U13580 (N_13580,N_13108,N_13233);
and U13581 (N_13581,N_13488,N_13379);
nand U13582 (N_13582,N_13006,N_13437);
xnor U13583 (N_13583,N_13316,N_13090);
and U13584 (N_13584,N_13158,N_13322);
nand U13585 (N_13585,N_13375,N_13218);
or U13586 (N_13586,N_13299,N_13391);
nor U13587 (N_13587,N_13495,N_13204);
or U13588 (N_13588,N_13492,N_13284);
or U13589 (N_13589,N_13424,N_13340);
xor U13590 (N_13590,N_13171,N_13366);
or U13591 (N_13591,N_13215,N_13306);
nand U13592 (N_13592,N_13460,N_13130);
nand U13593 (N_13593,N_13052,N_13167);
xnor U13594 (N_13594,N_13024,N_13194);
nand U13595 (N_13595,N_13011,N_13445);
nor U13596 (N_13596,N_13286,N_13041);
and U13597 (N_13597,N_13295,N_13141);
or U13598 (N_13598,N_13037,N_13021);
and U13599 (N_13599,N_13175,N_13137);
or U13600 (N_13600,N_13381,N_13270);
and U13601 (N_13601,N_13185,N_13369);
or U13602 (N_13602,N_13211,N_13080);
or U13603 (N_13603,N_13420,N_13116);
xnor U13604 (N_13604,N_13331,N_13066);
and U13605 (N_13605,N_13472,N_13287);
xnor U13606 (N_13606,N_13311,N_13285);
nor U13607 (N_13607,N_13188,N_13231);
and U13608 (N_13608,N_13441,N_13043);
and U13609 (N_13609,N_13073,N_13182);
or U13610 (N_13610,N_13449,N_13390);
or U13611 (N_13611,N_13497,N_13294);
nor U13612 (N_13612,N_13480,N_13029);
and U13613 (N_13613,N_13479,N_13465);
xnor U13614 (N_13614,N_13446,N_13104);
and U13615 (N_13615,N_13368,N_13067);
xnor U13616 (N_13616,N_13193,N_13170);
nor U13617 (N_13617,N_13361,N_13148);
and U13618 (N_13618,N_13060,N_13452);
and U13619 (N_13619,N_13358,N_13126);
nand U13620 (N_13620,N_13181,N_13138);
xor U13621 (N_13621,N_13404,N_13121);
nor U13622 (N_13622,N_13337,N_13103);
nand U13623 (N_13623,N_13491,N_13260);
xnor U13624 (N_13624,N_13150,N_13261);
or U13625 (N_13625,N_13199,N_13419);
and U13626 (N_13626,N_13411,N_13440);
nor U13627 (N_13627,N_13044,N_13432);
nand U13628 (N_13628,N_13042,N_13442);
xor U13629 (N_13629,N_13324,N_13002);
and U13630 (N_13630,N_13200,N_13191);
nand U13631 (N_13631,N_13255,N_13085);
or U13632 (N_13632,N_13054,N_13022);
xnor U13633 (N_13633,N_13025,N_13061);
or U13634 (N_13634,N_13228,N_13192);
and U13635 (N_13635,N_13293,N_13034);
or U13636 (N_13636,N_13109,N_13305);
xor U13637 (N_13637,N_13367,N_13102);
and U13638 (N_13638,N_13064,N_13169);
and U13639 (N_13639,N_13407,N_13254);
nand U13640 (N_13640,N_13307,N_13069);
nor U13641 (N_13641,N_13273,N_13235);
xnor U13642 (N_13642,N_13246,N_13013);
nor U13643 (N_13643,N_13461,N_13074);
and U13644 (N_13644,N_13476,N_13028);
nor U13645 (N_13645,N_13055,N_13482);
or U13646 (N_13646,N_13049,N_13081);
xor U13647 (N_13647,N_13119,N_13009);
and U13648 (N_13648,N_13389,N_13243);
and U13649 (N_13649,N_13164,N_13244);
nor U13650 (N_13650,N_13344,N_13234);
and U13651 (N_13651,N_13257,N_13422);
or U13652 (N_13652,N_13091,N_13012);
or U13653 (N_13653,N_13184,N_13124);
or U13654 (N_13654,N_13334,N_13359);
nor U13655 (N_13655,N_13302,N_13160);
xnor U13656 (N_13656,N_13312,N_13475);
and U13657 (N_13657,N_13032,N_13253);
nor U13658 (N_13658,N_13178,N_13356);
nor U13659 (N_13659,N_13112,N_13107);
nand U13660 (N_13660,N_13325,N_13088);
and U13661 (N_13661,N_13053,N_13223);
and U13662 (N_13662,N_13071,N_13105);
xnor U13663 (N_13663,N_13122,N_13250);
nor U13664 (N_13664,N_13386,N_13026);
nor U13665 (N_13665,N_13161,N_13149);
nand U13666 (N_13666,N_13267,N_13209);
xor U13667 (N_13667,N_13494,N_13483);
nor U13668 (N_13668,N_13196,N_13403);
nand U13669 (N_13669,N_13426,N_13400);
or U13670 (N_13670,N_13117,N_13120);
or U13671 (N_13671,N_13245,N_13496);
nand U13672 (N_13672,N_13030,N_13077);
nand U13673 (N_13673,N_13314,N_13444);
nand U13674 (N_13674,N_13154,N_13151);
and U13675 (N_13675,N_13280,N_13168);
xor U13676 (N_13676,N_13454,N_13163);
xor U13677 (N_13677,N_13341,N_13027);
nand U13678 (N_13678,N_13288,N_13405);
xnor U13679 (N_13679,N_13330,N_13321);
nand U13680 (N_13680,N_13153,N_13232);
or U13681 (N_13681,N_13428,N_13443);
nor U13682 (N_13682,N_13395,N_13362);
and U13683 (N_13683,N_13183,N_13329);
or U13684 (N_13684,N_13372,N_13058);
or U13685 (N_13685,N_13050,N_13377);
and U13686 (N_13686,N_13448,N_13469);
and U13687 (N_13687,N_13145,N_13075);
nor U13688 (N_13688,N_13350,N_13247);
nand U13689 (N_13689,N_13097,N_13408);
and U13690 (N_13690,N_13010,N_13439);
nor U13691 (N_13691,N_13427,N_13140);
and U13692 (N_13692,N_13039,N_13409);
and U13693 (N_13693,N_13387,N_13219);
xor U13694 (N_13694,N_13320,N_13018);
or U13695 (N_13695,N_13498,N_13224);
or U13696 (N_13696,N_13087,N_13031);
or U13697 (N_13697,N_13353,N_13142);
nand U13698 (N_13698,N_13033,N_13456);
nor U13699 (N_13699,N_13155,N_13463);
xnor U13700 (N_13700,N_13236,N_13222);
or U13701 (N_13701,N_13251,N_13297);
nor U13702 (N_13702,N_13327,N_13323);
or U13703 (N_13703,N_13004,N_13086);
nand U13704 (N_13704,N_13453,N_13098);
nand U13705 (N_13705,N_13478,N_13289);
nor U13706 (N_13706,N_13198,N_13347);
nand U13707 (N_13707,N_13272,N_13485);
xnor U13708 (N_13708,N_13201,N_13190);
nand U13709 (N_13709,N_13278,N_13240);
nor U13710 (N_13710,N_13113,N_13406);
nor U13711 (N_13711,N_13385,N_13292);
and U13712 (N_13712,N_13319,N_13176);
nor U13713 (N_13713,N_13000,N_13413);
nor U13714 (N_13714,N_13450,N_13202);
xnor U13715 (N_13715,N_13326,N_13095);
or U13716 (N_13716,N_13128,N_13263);
nor U13717 (N_13717,N_13173,N_13378);
and U13718 (N_13718,N_13313,N_13388);
and U13719 (N_13719,N_13123,N_13096);
nand U13720 (N_13720,N_13036,N_13468);
nor U13721 (N_13721,N_13070,N_13062);
or U13722 (N_13722,N_13241,N_13017);
xnor U13723 (N_13723,N_13111,N_13370);
xnor U13724 (N_13724,N_13339,N_13047);
xor U13725 (N_13725,N_13402,N_13397);
nor U13726 (N_13726,N_13045,N_13248);
xor U13727 (N_13727,N_13237,N_13165);
and U13728 (N_13728,N_13457,N_13410);
xor U13729 (N_13729,N_13351,N_13114);
and U13730 (N_13730,N_13059,N_13065);
nor U13731 (N_13731,N_13099,N_13493);
and U13732 (N_13732,N_13213,N_13373);
or U13733 (N_13733,N_13279,N_13106);
or U13734 (N_13734,N_13093,N_13274);
and U13735 (N_13735,N_13484,N_13076);
nand U13736 (N_13736,N_13499,N_13057);
or U13737 (N_13737,N_13338,N_13035);
nand U13738 (N_13738,N_13146,N_13135);
xnor U13739 (N_13739,N_13118,N_13048);
or U13740 (N_13740,N_13264,N_13318);
nand U13741 (N_13741,N_13212,N_13317);
and U13742 (N_13742,N_13364,N_13214);
nor U13743 (N_13743,N_13430,N_13357);
nand U13744 (N_13744,N_13401,N_13007);
nand U13745 (N_13745,N_13392,N_13464);
nor U13746 (N_13746,N_13335,N_13477);
and U13747 (N_13747,N_13249,N_13365);
nand U13748 (N_13748,N_13486,N_13208);
nand U13749 (N_13749,N_13115,N_13291);
nor U13750 (N_13750,N_13009,N_13392);
nor U13751 (N_13751,N_13097,N_13269);
or U13752 (N_13752,N_13003,N_13186);
nor U13753 (N_13753,N_13248,N_13282);
or U13754 (N_13754,N_13102,N_13394);
nand U13755 (N_13755,N_13366,N_13215);
xor U13756 (N_13756,N_13365,N_13008);
nor U13757 (N_13757,N_13319,N_13022);
and U13758 (N_13758,N_13240,N_13321);
or U13759 (N_13759,N_13444,N_13294);
xor U13760 (N_13760,N_13029,N_13416);
xnor U13761 (N_13761,N_13336,N_13163);
xnor U13762 (N_13762,N_13131,N_13097);
or U13763 (N_13763,N_13432,N_13374);
nor U13764 (N_13764,N_13239,N_13406);
or U13765 (N_13765,N_13071,N_13142);
nor U13766 (N_13766,N_13322,N_13120);
and U13767 (N_13767,N_13233,N_13176);
nand U13768 (N_13768,N_13334,N_13125);
nor U13769 (N_13769,N_13290,N_13262);
xor U13770 (N_13770,N_13464,N_13461);
nor U13771 (N_13771,N_13112,N_13079);
or U13772 (N_13772,N_13403,N_13127);
and U13773 (N_13773,N_13168,N_13135);
nand U13774 (N_13774,N_13333,N_13272);
nand U13775 (N_13775,N_13181,N_13150);
or U13776 (N_13776,N_13308,N_13418);
nand U13777 (N_13777,N_13115,N_13190);
xor U13778 (N_13778,N_13335,N_13428);
nand U13779 (N_13779,N_13122,N_13084);
xnor U13780 (N_13780,N_13080,N_13262);
nor U13781 (N_13781,N_13248,N_13349);
or U13782 (N_13782,N_13387,N_13053);
and U13783 (N_13783,N_13353,N_13130);
xor U13784 (N_13784,N_13127,N_13440);
nand U13785 (N_13785,N_13334,N_13118);
nand U13786 (N_13786,N_13242,N_13192);
nand U13787 (N_13787,N_13370,N_13235);
nand U13788 (N_13788,N_13400,N_13210);
nand U13789 (N_13789,N_13101,N_13355);
nor U13790 (N_13790,N_13347,N_13402);
or U13791 (N_13791,N_13220,N_13325);
xor U13792 (N_13792,N_13160,N_13145);
and U13793 (N_13793,N_13493,N_13051);
xor U13794 (N_13794,N_13002,N_13131);
and U13795 (N_13795,N_13354,N_13133);
and U13796 (N_13796,N_13296,N_13179);
nand U13797 (N_13797,N_13404,N_13156);
or U13798 (N_13798,N_13078,N_13222);
or U13799 (N_13799,N_13491,N_13353);
xnor U13800 (N_13800,N_13306,N_13116);
xor U13801 (N_13801,N_13340,N_13139);
or U13802 (N_13802,N_13010,N_13211);
nor U13803 (N_13803,N_13016,N_13165);
xor U13804 (N_13804,N_13158,N_13088);
nor U13805 (N_13805,N_13337,N_13067);
nor U13806 (N_13806,N_13088,N_13115);
nor U13807 (N_13807,N_13189,N_13071);
and U13808 (N_13808,N_13449,N_13334);
nor U13809 (N_13809,N_13393,N_13147);
and U13810 (N_13810,N_13451,N_13346);
nand U13811 (N_13811,N_13209,N_13106);
and U13812 (N_13812,N_13493,N_13135);
nand U13813 (N_13813,N_13202,N_13309);
nor U13814 (N_13814,N_13221,N_13301);
xnor U13815 (N_13815,N_13153,N_13159);
xnor U13816 (N_13816,N_13252,N_13091);
nor U13817 (N_13817,N_13191,N_13324);
nor U13818 (N_13818,N_13034,N_13053);
or U13819 (N_13819,N_13022,N_13406);
nand U13820 (N_13820,N_13414,N_13310);
nor U13821 (N_13821,N_13258,N_13494);
or U13822 (N_13822,N_13373,N_13302);
nor U13823 (N_13823,N_13105,N_13429);
nor U13824 (N_13824,N_13060,N_13383);
and U13825 (N_13825,N_13203,N_13050);
nor U13826 (N_13826,N_13279,N_13250);
or U13827 (N_13827,N_13404,N_13415);
and U13828 (N_13828,N_13083,N_13069);
and U13829 (N_13829,N_13412,N_13359);
nor U13830 (N_13830,N_13388,N_13399);
nor U13831 (N_13831,N_13010,N_13386);
nand U13832 (N_13832,N_13220,N_13466);
xor U13833 (N_13833,N_13356,N_13345);
xnor U13834 (N_13834,N_13037,N_13225);
nor U13835 (N_13835,N_13206,N_13356);
nand U13836 (N_13836,N_13285,N_13484);
xnor U13837 (N_13837,N_13296,N_13113);
or U13838 (N_13838,N_13258,N_13203);
nand U13839 (N_13839,N_13449,N_13006);
xor U13840 (N_13840,N_13212,N_13146);
nor U13841 (N_13841,N_13136,N_13123);
or U13842 (N_13842,N_13127,N_13303);
or U13843 (N_13843,N_13280,N_13263);
nor U13844 (N_13844,N_13387,N_13350);
and U13845 (N_13845,N_13066,N_13459);
or U13846 (N_13846,N_13139,N_13377);
xor U13847 (N_13847,N_13298,N_13338);
xor U13848 (N_13848,N_13043,N_13313);
xnor U13849 (N_13849,N_13374,N_13044);
nand U13850 (N_13850,N_13117,N_13123);
nand U13851 (N_13851,N_13092,N_13148);
nand U13852 (N_13852,N_13008,N_13136);
or U13853 (N_13853,N_13013,N_13039);
or U13854 (N_13854,N_13243,N_13185);
nor U13855 (N_13855,N_13145,N_13370);
and U13856 (N_13856,N_13335,N_13458);
or U13857 (N_13857,N_13490,N_13416);
nand U13858 (N_13858,N_13469,N_13025);
xor U13859 (N_13859,N_13237,N_13343);
nand U13860 (N_13860,N_13239,N_13440);
or U13861 (N_13861,N_13270,N_13241);
or U13862 (N_13862,N_13269,N_13043);
xor U13863 (N_13863,N_13155,N_13066);
nor U13864 (N_13864,N_13113,N_13121);
xor U13865 (N_13865,N_13064,N_13439);
xnor U13866 (N_13866,N_13310,N_13053);
nand U13867 (N_13867,N_13004,N_13002);
and U13868 (N_13868,N_13404,N_13114);
or U13869 (N_13869,N_13084,N_13261);
or U13870 (N_13870,N_13393,N_13306);
and U13871 (N_13871,N_13100,N_13462);
nand U13872 (N_13872,N_13388,N_13319);
nor U13873 (N_13873,N_13069,N_13392);
xnor U13874 (N_13874,N_13205,N_13460);
nor U13875 (N_13875,N_13131,N_13098);
xor U13876 (N_13876,N_13290,N_13237);
and U13877 (N_13877,N_13066,N_13055);
or U13878 (N_13878,N_13415,N_13034);
nand U13879 (N_13879,N_13432,N_13063);
and U13880 (N_13880,N_13297,N_13163);
xor U13881 (N_13881,N_13422,N_13159);
or U13882 (N_13882,N_13459,N_13464);
or U13883 (N_13883,N_13304,N_13430);
nor U13884 (N_13884,N_13367,N_13148);
or U13885 (N_13885,N_13306,N_13488);
or U13886 (N_13886,N_13064,N_13225);
xnor U13887 (N_13887,N_13323,N_13350);
xnor U13888 (N_13888,N_13083,N_13336);
xor U13889 (N_13889,N_13056,N_13378);
xnor U13890 (N_13890,N_13001,N_13028);
nand U13891 (N_13891,N_13402,N_13342);
nor U13892 (N_13892,N_13171,N_13270);
or U13893 (N_13893,N_13226,N_13135);
and U13894 (N_13894,N_13381,N_13443);
xor U13895 (N_13895,N_13321,N_13065);
xor U13896 (N_13896,N_13025,N_13402);
xnor U13897 (N_13897,N_13437,N_13447);
or U13898 (N_13898,N_13007,N_13214);
and U13899 (N_13899,N_13188,N_13258);
and U13900 (N_13900,N_13262,N_13339);
xor U13901 (N_13901,N_13436,N_13043);
nor U13902 (N_13902,N_13211,N_13224);
nor U13903 (N_13903,N_13319,N_13324);
nand U13904 (N_13904,N_13030,N_13110);
or U13905 (N_13905,N_13159,N_13092);
or U13906 (N_13906,N_13290,N_13203);
nand U13907 (N_13907,N_13323,N_13081);
and U13908 (N_13908,N_13314,N_13456);
xor U13909 (N_13909,N_13212,N_13282);
or U13910 (N_13910,N_13274,N_13313);
nor U13911 (N_13911,N_13186,N_13404);
and U13912 (N_13912,N_13437,N_13182);
nand U13913 (N_13913,N_13235,N_13103);
or U13914 (N_13914,N_13302,N_13333);
nand U13915 (N_13915,N_13053,N_13457);
nand U13916 (N_13916,N_13448,N_13414);
nor U13917 (N_13917,N_13009,N_13472);
xnor U13918 (N_13918,N_13300,N_13067);
nor U13919 (N_13919,N_13369,N_13153);
nor U13920 (N_13920,N_13228,N_13453);
xnor U13921 (N_13921,N_13142,N_13472);
nor U13922 (N_13922,N_13109,N_13296);
and U13923 (N_13923,N_13319,N_13490);
nand U13924 (N_13924,N_13105,N_13236);
or U13925 (N_13925,N_13322,N_13259);
nor U13926 (N_13926,N_13283,N_13434);
nand U13927 (N_13927,N_13043,N_13213);
and U13928 (N_13928,N_13460,N_13188);
nand U13929 (N_13929,N_13222,N_13159);
nand U13930 (N_13930,N_13088,N_13036);
and U13931 (N_13931,N_13119,N_13335);
or U13932 (N_13932,N_13368,N_13080);
or U13933 (N_13933,N_13370,N_13317);
nor U13934 (N_13934,N_13464,N_13333);
and U13935 (N_13935,N_13386,N_13462);
and U13936 (N_13936,N_13240,N_13299);
nand U13937 (N_13937,N_13173,N_13063);
or U13938 (N_13938,N_13341,N_13055);
nor U13939 (N_13939,N_13170,N_13103);
nand U13940 (N_13940,N_13479,N_13065);
nor U13941 (N_13941,N_13324,N_13225);
xnor U13942 (N_13942,N_13345,N_13093);
nor U13943 (N_13943,N_13233,N_13399);
and U13944 (N_13944,N_13352,N_13193);
xnor U13945 (N_13945,N_13443,N_13071);
nand U13946 (N_13946,N_13031,N_13456);
or U13947 (N_13947,N_13436,N_13037);
xnor U13948 (N_13948,N_13087,N_13280);
nand U13949 (N_13949,N_13282,N_13178);
and U13950 (N_13950,N_13338,N_13481);
nor U13951 (N_13951,N_13022,N_13279);
nor U13952 (N_13952,N_13135,N_13148);
nand U13953 (N_13953,N_13221,N_13384);
nand U13954 (N_13954,N_13295,N_13073);
and U13955 (N_13955,N_13213,N_13020);
or U13956 (N_13956,N_13161,N_13224);
or U13957 (N_13957,N_13432,N_13195);
nand U13958 (N_13958,N_13425,N_13059);
or U13959 (N_13959,N_13147,N_13405);
nor U13960 (N_13960,N_13399,N_13479);
nor U13961 (N_13961,N_13428,N_13065);
xnor U13962 (N_13962,N_13099,N_13152);
nand U13963 (N_13963,N_13449,N_13236);
and U13964 (N_13964,N_13491,N_13216);
and U13965 (N_13965,N_13396,N_13110);
xnor U13966 (N_13966,N_13164,N_13038);
nor U13967 (N_13967,N_13073,N_13099);
and U13968 (N_13968,N_13085,N_13142);
nand U13969 (N_13969,N_13309,N_13469);
or U13970 (N_13970,N_13222,N_13029);
and U13971 (N_13971,N_13047,N_13234);
nand U13972 (N_13972,N_13219,N_13203);
xnor U13973 (N_13973,N_13419,N_13260);
and U13974 (N_13974,N_13190,N_13240);
or U13975 (N_13975,N_13181,N_13417);
nor U13976 (N_13976,N_13061,N_13351);
nor U13977 (N_13977,N_13398,N_13351);
nand U13978 (N_13978,N_13301,N_13401);
and U13979 (N_13979,N_13208,N_13128);
xnor U13980 (N_13980,N_13332,N_13449);
nand U13981 (N_13981,N_13414,N_13297);
or U13982 (N_13982,N_13041,N_13240);
and U13983 (N_13983,N_13045,N_13468);
or U13984 (N_13984,N_13096,N_13258);
nand U13985 (N_13985,N_13211,N_13330);
xnor U13986 (N_13986,N_13478,N_13122);
and U13987 (N_13987,N_13476,N_13113);
nor U13988 (N_13988,N_13408,N_13197);
xor U13989 (N_13989,N_13327,N_13279);
or U13990 (N_13990,N_13491,N_13015);
xnor U13991 (N_13991,N_13190,N_13077);
nand U13992 (N_13992,N_13135,N_13331);
nor U13993 (N_13993,N_13033,N_13142);
or U13994 (N_13994,N_13319,N_13234);
nor U13995 (N_13995,N_13290,N_13388);
and U13996 (N_13996,N_13171,N_13168);
xor U13997 (N_13997,N_13421,N_13266);
nand U13998 (N_13998,N_13319,N_13328);
nand U13999 (N_13999,N_13262,N_13186);
nor U14000 (N_14000,N_13585,N_13559);
or U14001 (N_14001,N_13506,N_13829);
xnor U14002 (N_14002,N_13670,N_13894);
xnor U14003 (N_14003,N_13715,N_13796);
nand U14004 (N_14004,N_13648,N_13930);
and U14005 (N_14005,N_13754,N_13953);
xor U14006 (N_14006,N_13693,N_13553);
xnor U14007 (N_14007,N_13826,N_13816);
or U14008 (N_14008,N_13925,N_13575);
and U14009 (N_14009,N_13966,N_13918);
nand U14010 (N_14010,N_13602,N_13781);
and U14011 (N_14011,N_13561,N_13740);
and U14012 (N_14012,N_13827,N_13954);
and U14013 (N_14013,N_13980,N_13872);
xor U14014 (N_14014,N_13916,N_13775);
or U14015 (N_14015,N_13712,N_13755);
nor U14016 (N_14016,N_13586,N_13505);
or U14017 (N_14017,N_13937,N_13919);
xnor U14018 (N_14018,N_13650,N_13717);
and U14019 (N_14019,N_13676,N_13870);
nor U14020 (N_14020,N_13901,N_13514);
nor U14021 (N_14021,N_13612,N_13519);
or U14022 (N_14022,N_13532,N_13965);
and U14023 (N_14023,N_13773,N_13944);
and U14024 (N_14024,N_13964,N_13524);
and U14025 (N_14025,N_13782,N_13959);
and U14026 (N_14026,N_13578,N_13613);
xnor U14027 (N_14027,N_13579,N_13713);
nand U14028 (N_14028,N_13837,N_13511);
xnor U14029 (N_14029,N_13991,N_13839);
nor U14030 (N_14030,N_13685,N_13683);
or U14031 (N_14031,N_13596,N_13656);
nand U14032 (N_14032,N_13800,N_13748);
xnor U14033 (N_14033,N_13645,N_13619);
nor U14034 (N_14034,N_13635,N_13507);
nor U14035 (N_14035,N_13525,N_13832);
and U14036 (N_14036,N_13622,N_13743);
or U14037 (N_14037,N_13897,N_13787);
or U14038 (N_14038,N_13828,N_13523);
and U14039 (N_14039,N_13794,N_13709);
nor U14040 (N_14040,N_13915,N_13732);
xor U14041 (N_14041,N_13746,N_13988);
nand U14042 (N_14042,N_13632,N_13616);
or U14043 (N_14043,N_13863,N_13821);
or U14044 (N_14044,N_13889,N_13730);
and U14045 (N_14045,N_13694,N_13544);
or U14046 (N_14046,N_13878,N_13929);
xor U14047 (N_14047,N_13690,N_13719);
xnor U14048 (N_14048,N_13677,N_13567);
xnor U14049 (N_14049,N_13842,N_13577);
nand U14050 (N_14050,N_13593,N_13984);
or U14051 (N_14051,N_13531,N_13974);
nand U14052 (N_14052,N_13551,N_13735);
or U14053 (N_14053,N_13806,N_13851);
nand U14054 (N_14054,N_13776,N_13741);
nor U14055 (N_14055,N_13571,N_13687);
nand U14056 (N_14056,N_13810,N_13949);
nand U14057 (N_14057,N_13757,N_13910);
and U14058 (N_14058,N_13812,N_13627);
nand U14059 (N_14059,N_13873,N_13900);
nand U14060 (N_14060,N_13550,N_13720);
and U14061 (N_14061,N_13983,N_13729);
and U14062 (N_14062,N_13856,N_13945);
xor U14063 (N_14063,N_13665,N_13847);
nor U14064 (N_14064,N_13722,N_13912);
xnor U14065 (N_14065,N_13589,N_13660);
nand U14066 (N_14066,N_13814,N_13688);
nand U14067 (N_14067,N_13633,N_13750);
nor U14068 (N_14068,N_13601,N_13646);
nand U14069 (N_14069,N_13769,N_13533);
nand U14070 (N_14070,N_13970,N_13811);
xor U14071 (N_14071,N_13540,N_13914);
nor U14072 (N_14072,N_13887,N_13555);
or U14073 (N_14073,N_13600,N_13946);
or U14074 (N_14074,N_13907,N_13809);
nor U14075 (N_14075,N_13948,N_13788);
and U14076 (N_14076,N_13819,N_13671);
xnor U14077 (N_14077,N_13536,N_13584);
nor U14078 (N_14078,N_13998,N_13591);
nor U14079 (N_14079,N_13695,N_13611);
and U14080 (N_14080,N_13513,N_13568);
nor U14081 (N_14081,N_13768,N_13880);
and U14082 (N_14082,N_13744,N_13637);
nand U14083 (N_14083,N_13888,N_13977);
nand U14084 (N_14084,N_13512,N_13858);
nand U14085 (N_14085,N_13831,N_13904);
xnor U14086 (N_14086,N_13640,N_13699);
and U14087 (N_14087,N_13967,N_13803);
nand U14088 (N_14088,N_13902,N_13700);
or U14089 (N_14089,N_13994,N_13905);
and U14090 (N_14090,N_13997,N_13569);
xor U14091 (N_14091,N_13799,N_13588);
xnor U14092 (N_14092,N_13868,N_13557);
or U14093 (N_14093,N_13751,N_13598);
nor U14094 (N_14094,N_13728,N_13978);
xor U14095 (N_14095,N_13960,N_13716);
or U14096 (N_14096,N_13864,N_13834);
and U14097 (N_14097,N_13556,N_13583);
nand U14098 (N_14098,N_13982,N_13824);
nor U14099 (N_14099,N_13893,N_13807);
and U14100 (N_14100,N_13668,N_13539);
and U14101 (N_14101,N_13552,N_13922);
or U14102 (N_14102,N_13835,N_13767);
xor U14103 (N_14103,N_13825,N_13770);
or U14104 (N_14104,N_13724,N_13943);
and U14105 (N_14105,N_13667,N_13651);
nand U14106 (N_14106,N_13517,N_13989);
and U14107 (N_14107,N_13830,N_13845);
nand U14108 (N_14108,N_13500,N_13617);
nand U14109 (N_14109,N_13502,N_13662);
and U14110 (N_14110,N_13529,N_13815);
xor U14111 (N_14111,N_13817,N_13779);
and U14112 (N_14112,N_13681,N_13697);
and U14113 (N_14113,N_13976,N_13756);
or U14114 (N_14114,N_13594,N_13638);
and U14115 (N_14115,N_13874,N_13990);
or U14116 (N_14116,N_13917,N_13896);
nand U14117 (N_14117,N_13886,N_13860);
nand U14118 (N_14118,N_13765,N_13985);
nor U14119 (N_14119,N_13762,N_13789);
xor U14120 (N_14120,N_13706,N_13672);
or U14121 (N_14121,N_13698,N_13790);
xor U14122 (N_14122,N_13726,N_13657);
or U14123 (N_14123,N_13626,N_13503);
xnor U14124 (N_14124,N_13913,N_13521);
xor U14125 (N_14125,N_13603,N_13639);
or U14126 (N_14126,N_13747,N_13924);
and U14127 (N_14127,N_13802,N_13701);
nand U14128 (N_14128,N_13636,N_13582);
and U14129 (N_14129,N_13962,N_13666);
nand U14130 (N_14130,N_13642,N_13574);
xor U14131 (N_14131,N_13752,N_13804);
nor U14132 (N_14132,N_13961,N_13703);
nand U14133 (N_14133,N_13771,N_13624);
or U14134 (N_14134,N_13778,N_13931);
nor U14135 (N_14135,N_13761,N_13623);
nand U14136 (N_14136,N_13908,N_13869);
and U14137 (N_14137,N_13801,N_13963);
nor U14138 (N_14138,N_13721,N_13675);
and U14139 (N_14139,N_13508,N_13659);
and U14140 (N_14140,N_13597,N_13655);
nand U14141 (N_14141,N_13705,N_13823);
nor U14142 (N_14142,N_13766,N_13971);
nor U14143 (N_14143,N_13879,N_13999);
nand U14144 (N_14144,N_13509,N_13899);
and U14145 (N_14145,N_13947,N_13620);
xor U14146 (N_14146,N_13956,N_13867);
nand U14147 (N_14147,N_13711,N_13714);
nor U14148 (N_14148,N_13684,N_13760);
xor U14149 (N_14149,N_13680,N_13951);
nand U14150 (N_14150,N_13798,N_13504);
nor U14151 (N_14151,N_13836,N_13822);
or U14152 (N_14152,N_13933,N_13973);
nand U14153 (N_14153,N_13840,N_13883);
nand U14154 (N_14154,N_13727,N_13805);
nand U14155 (N_14155,N_13673,N_13647);
nand U14156 (N_14156,N_13759,N_13573);
and U14157 (N_14157,N_13877,N_13926);
or U14158 (N_14158,N_13604,N_13610);
nor U14159 (N_14159,N_13534,N_13691);
xnor U14160 (N_14160,N_13526,N_13774);
or U14161 (N_14161,N_13981,N_13618);
or U14162 (N_14162,N_13696,N_13793);
or U14163 (N_14163,N_13590,N_13621);
or U14164 (N_14164,N_13848,N_13562);
nand U14165 (N_14165,N_13609,N_13891);
or U14166 (N_14166,N_13634,N_13758);
nor U14167 (N_14167,N_13707,N_13643);
or U14168 (N_14168,N_13975,N_13846);
nor U14169 (N_14169,N_13733,N_13849);
or U14170 (N_14170,N_13795,N_13565);
or U14171 (N_14171,N_13935,N_13841);
nand U14172 (N_14172,N_13663,N_13576);
nor U14173 (N_14173,N_13535,N_13784);
xor U14174 (N_14174,N_13547,N_13736);
and U14175 (N_14175,N_13686,N_13942);
nand U14176 (N_14176,N_13852,N_13838);
or U14177 (N_14177,N_13987,N_13853);
or U14178 (N_14178,N_13518,N_13969);
and U14179 (N_14179,N_13857,N_13629);
or U14180 (N_14180,N_13543,N_13996);
xor U14181 (N_14181,N_13797,N_13530);
nand U14182 (N_14182,N_13928,N_13510);
or U14183 (N_14183,N_13844,N_13850);
or U14184 (N_14184,N_13738,N_13678);
or U14185 (N_14185,N_13725,N_13866);
xnor U14186 (N_14186,N_13932,N_13772);
xnor U14187 (N_14187,N_13921,N_13558);
or U14188 (N_14188,N_13560,N_13861);
xnor U14189 (N_14189,N_13895,N_13545);
or U14190 (N_14190,N_13911,N_13516);
or U14191 (N_14191,N_13661,N_13906);
nor U14192 (N_14192,N_13763,N_13527);
and U14193 (N_14193,N_13792,N_13689);
or U14194 (N_14194,N_13674,N_13936);
and U14195 (N_14195,N_13958,N_13679);
nor U14196 (N_14196,N_13538,N_13742);
xor U14197 (N_14197,N_13731,N_13615);
and U14198 (N_14198,N_13520,N_13702);
or U14199 (N_14199,N_13764,N_13554);
nor U14200 (N_14200,N_13813,N_13876);
nand U14201 (N_14201,N_13934,N_13808);
nand U14202 (N_14202,N_13909,N_13938);
nor U14203 (N_14203,N_13952,N_13882);
nand U14204 (N_14204,N_13992,N_13979);
xor U14205 (N_14205,N_13780,N_13957);
nand U14206 (N_14206,N_13941,N_13630);
and U14207 (N_14207,N_13570,N_13708);
and U14208 (N_14208,N_13820,N_13881);
xor U14209 (N_14209,N_13972,N_13605);
xor U14210 (N_14210,N_13572,N_13739);
or U14211 (N_14211,N_13875,N_13892);
or U14212 (N_14212,N_13542,N_13898);
nor U14213 (N_14213,N_13608,N_13749);
nand U14214 (N_14214,N_13993,N_13692);
or U14215 (N_14215,N_13537,N_13777);
xor U14216 (N_14216,N_13682,N_13607);
and U14217 (N_14217,N_13791,N_13625);
or U14218 (N_14218,N_13871,N_13753);
and U14219 (N_14219,N_13885,N_13606);
xor U14220 (N_14220,N_13920,N_13541);
xnor U14221 (N_14221,N_13785,N_13854);
nand U14222 (N_14222,N_13986,N_13939);
nor U14223 (N_14223,N_13734,N_13704);
xnor U14224 (N_14224,N_13669,N_13501);
nand U14225 (N_14225,N_13890,N_13923);
nand U14226 (N_14226,N_13843,N_13718);
or U14227 (N_14227,N_13745,N_13546);
xnor U14228 (N_14228,N_13581,N_13595);
nand U14229 (N_14229,N_13940,N_13723);
nor U14230 (N_14230,N_13710,N_13903);
and U14231 (N_14231,N_13566,N_13833);
xnor U14232 (N_14232,N_13783,N_13995);
and U14233 (N_14233,N_13652,N_13950);
xor U14234 (N_14234,N_13587,N_13884);
and U14235 (N_14235,N_13644,N_13865);
nand U14236 (N_14236,N_13515,N_13522);
xnor U14237 (N_14237,N_13641,N_13592);
and U14238 (N_14238,N_13528,N_13549);
xnor U14239 (N_14239,N_13599,N_13859);
nor U14240 (N_14240,N_13580,N_13649);
and U14241 (N_14241,N_13653,N_13786);
xnor U14242 (N_14242,N_13855,N_13654);
and U14243 (N_14243,N_13631,N_13818);
xor U14244 (N_14244,N_13563,N_13862);
xnor U14245 (N_14245,N_13658,N_13955);
or U14246 (N_14246,N_13564,N_13614);
nor U14247 (N_14247,N_13548,N_13737);
and U14248 (N_14248,N_13968,N_13664);
xnor U14249 (N_14249,N_13628,N_13927);
nand U14250 (N_14250,N_13749,N_13780);
xor U14251 (N_14251,N_13502,N_13604);
or U14252 (N_14252,N_13701,N_13861);
nor U14253 (N_14253,N_13947,N_13617);
nand U14254 (N_14254,N_13983,N_13864);
xnor U14255 (N_14255,N_13740,N_13904);
and U14256 (N_14256,N_13784,N_13885);
nand U14257 (N_14257,N_13835,N_13516);
and U14258 (N_14258,N_13608,N_13787);
nand U14259 (N_14259,N_13521,N_13944);
and U14260 (N_14260,N_13890,N_13971);
nor U14261 (N_14261,N_13598,N_13582);
nor U14262 (N_14262,N_13606,N_13714);
xnor U14263 (N_14263,N_13653,N_13919);
nor U14264 (N_14264,N_13581,N_13630);
or U14265 (N_14265,N_13939,N_13883);
nand U14266 (N_14266,N_13612,N_13960);
nand U14267 (N_14267,N_13634,N_13728);
or U14268 (N_14268,N_13803,N_13684);
xor U14269 (N_14269,N_13655,N_13806);
nor U14270 (N_14270,N_13810,N_13618);
xnor U14271 (N_14271,N_13707,N_13564);
or U14272 (N_14272,N_13959,N_13891);
or U14273 (N_14273,N_13610,N_13586);
nor U14274 (N_14274,N_13511,N_13815);
nor U14275 (N_14275,N_13826,N_13790);
xor U14276 (N_14276,N_13614,N_13822);
and U14277 (N_14277,N_13815,N_13950);
nand U14278 (N_14278,N_13782,N_13775);
nand U14279 (N_14279,N_13930,N_13921);
and U14280 (N_14280,N_13796,N_13879);
nand U14281 (N_14281,N_13720,N_13892);
and U14282 (N_14282,N_13801,N_13926);
and U14283 (N_14283,N_13637,N_13918);
and U14284 (N_14284,N_13585,N_13955);
xor U14285 (N_14285,N_13732,N_13989);
and U14286 (N_14286,N_13870,N_13707);
and U14287 (N_14287,N_13890,N_13995);
or U14288 (N_14288,N_13978,N_13824);
and U14289 (N_14289,N_13621,N_13746);
or U14290 (N_14290,N_13653,N_13588);
nand U14291 (N_14291,N_13930,N_13922);
and U14292 (N_14292,N_13646,N_13589);
and U14293 (N_14293,N_13946,N_13755);
xnor U14294 (N_14294,N_13937,N_13668);
nand U14295 (N_14295,N_13515,N_13680);
and U14296 (N_14296,N_13594,N_13528);
and U14297 (N_14297,N_13953,N_13637);
nor U14298 (N_14298,N_13576,N_13504);
nor U14299 (N_14299,N_13946,N_13575);
nand U14300 (N_14300,N_13771,N_13775);
nand U14301 (N_14301,N_13877,N_13993);
or U14302 (N_14302,N_13828,N_13716);
nand U14303 (N_14303,N_13679,N_13592);
nor U14304 (N_14304,N_13862,N_13794);
and U14305 (N_14305,N_13994,N_13589);
nor U14306 (N_14306,N_13775,N_13922);
xnor U14307 (N_14307,N_13829,N_13988);
nor U14308 (N_14308,N_13550,N_13631);
xor U14309 (N_14309,N_13897,N_13700);
xnor U14310 (N_14310,N_13899,N_13936);
and U14311 (N_14311,N_13681,N_13617);
and U14312 (N_14312,N_13957,N_13619);
and U14313 (N_14313,N_13650,N_13762);
nand U14314 (N_14314,N_13584,N_13630);
nor U14315 (N_14315,N_13500,N_13683);
or U14316 (N_14316,N_13508,N_13720);
xor U14317 (N_14317,N_13517,N_13727);
nand U14318 (N_14318,N_13933,N_13603);
nand U14319 (N_14319,N_13808,N_13813);
nor U14320 (N_14320,N_13770,N_13691);
or U14321 (N_14321,N_13786,N_13754);
and U14322 (N_14322,N_13836,N_13859);
nor U14323 (N_14323,N_13993,N_13641);
xnor U14324 (N_14324,N_13852,N_13707);
xor U14325 (N_14325,N_13820,N_13733);
nor U14326 (N_14326,N_13566,N_13999);
or U14327 (N_14327,N_13548,N_13947);
nor U14328 (N_14328,N_13859,N_13621);
or U14329 (N_14329,N_13583,N_13863);
and U14330 (N_14330,N_13689,N_13731);
nand U14331 (N_14331,N_13738,N_13758);
nor U14332 (N_14332,N_13710,N_13664);
xor U14333 (N_14333,N_13707,N_13968);
nor U14334 (N_14334,N_13783,N_13676);
nor U14335 (N_14335,N_13746,N_13612);
and U14336 (N_14336,N_13519,N_13570);
xor U14337 (N_14337,N_13960,N_13802);
nand U14338 (N_14338,N_13946,N_13728);
nand U14339 (N_14339,N_13942,N_13739);
nand U14340 (N_14340,N_13530,N_13870);
nor U14341 (N_14341,N_13593,N_13711);
or U14342 (N_14342,N_13785,N_13847);
or U14343 (N_14343,N_13873,N_13696);
nor U14344 (N_14344,N_13707,N_13721);
and U14345 (N_14345,N_13504,N_13627);
xor U14346 (N_14346,N_13723,N_13897);
nand U14347 (N_14347,N_13895,N_13959);
nand U14348 (N_14348,N_13932,N_13964);
nand U14349 (N_14349,N_13825,N_13660);
xor U14350 (N_14350,N_13766,N_13826);
and U14351 (N_14351,N_13670,N_13924);
and U14352 (N_14352,N_13811,N_13539);
and U14353 (N_14353,N_13838,N_13794);
nand U14354 (N_14354,N_13758,N_13856);
xor U14355 (N_14355,N_13990,N_13713);
xor U14356 (N_14356,N_13986,N_13853);
or U14357 (N_14357,N_13564,N_13523);
xor U14358 (N_14358,N_13906,N_13880);
xnor U14359 (N_14359,N_13897,N_13859);
xor U14360 (N_14360,N_13533,N_13644);
or U14361 (N_14361,N_13539,N_13918);
xnor U14362 (N_14362,N_13573,N_13800);
nor U14363 (N_14363,N_13961,N_13707);
nor U14364 (N_14364,N_13574,N_13828);
nor U14365 (N_14365,N_13778,N_13766);
nor U14366 (N_14366,N_13979,N_13558);
xnor U14367 (N_14367,N_13999,N_13735);
nor U14368 (N_14368,N_13539,N_13680);
or U14369 (N_14369,N_13680,N_13511);
or U14370 (N_14370,N_13571,N_13718);
nand U14371 (N_14371,N_13837,N_13588);
xor U14372 (N_14372,N_13525,N_13739);
and U14373 (N_14373,N_13974,N_13726);
nor U14374 (N_14374,N_13549,N_13931);
xnor U14375 (N_14375,N_13583,N_13683);
nand U14376 (N_14376,N_13804,N_13776);
nor U14377 (N_14377,N_13896,N_13587);
nor U14378 (N_14378,N_13748,N_13752);
or U14379 (N_14379,N_13966,N_13733);
or U14380 (N_14380,N_13806,N_13774);
xnor U14381 (N_14381,N_13542,N_13643);
and U14382 (N_14382,N_13651,N_13859);
xor U14383 (N_14383,N_13843,N_13768);
xor U14384 (N_14384,N_13832,N_13961);
or U14385 (N_14385,N_13877,N_13819);
nor U14386 (N_14386,N_13516,N_13910);
and U14387 (N_14387,N_13819,N_13563);
nor U14388 (N_14388,N_13889,N_13946);
and U14389 (N_14389,N_13582,N_13859);
xnor U14390 (N_14390,N_13749,N_13997);
and U14391 (N_14391,N_13732,N_13542);
xnor U14392 (N_14392,N_13999,N_13898);
nor U14393 (N_14393,N_13756,N_13511);
nand U14394 (N_14394,N_13625,N_13631);
or U14395 (N_14395,N_13823,N_13990);
xnor U14396 (N_14396,N_13868,N_13502);
xor U14397 (N_14397,N_13673,N_13590);
or U14398 (N_14398,N_13617,N_13912);
and U14399 (N_14399,N_13944,N_13796);
nand U14400 (N_14400,N_13748,N_13910);
and U14401 (N_14401,N_13748,N_13965);
xor U14402 (N_14402,N_13512,N_13930);
xnor U14403 (N_14403,N_13636,N_13825);
xor U14404 (N_14404,N_13519,N_13902);
or U14405 (N_14405,N_13835,N_13915);
xnor U14406 (N_14406,N_13693,N_13983);
nor U14407 (N_14407,N_13808,N_13653);
xnor U14408 (N_14408,N_13868,N_13749);
and U14409 (N_14409,N_13854,N_13616);
and U14410 (N_14410,N_13976,N_13935);
xor U14411 (N_14411,N_13665,N_13650);
or U14412 (N_14412,N_13994,N_13582);
or U14413 (N_14413,N_13899,N_13561);
xor U14414 (N_14414,N_13815,N_13603);
or U14415 (N_14415,N_13916,N_13783);
and U14416 (N_14416,N_13543,N_13889);
nor U14417 (N_14417,N_13664,N_13882);
and U14418 (N_14418,N_13895,N_13734);
and U14419 (N_14419,N_13770,N_13802);
or U14420 (N_14420,N_13683,N_13863);
xnor U14421 (N_14421,N_13837,N_13845);
and U14422 (N_14422,N_13851,N_13514);
xnor U14423 (N_14423,N_13991,N_13953);
and U14424 (N_14424,N_13807,N_13633);
xnor U14425 (N_14425,N_13974,N_13898);
nor U14426 (N_14426,N_13609,N_13826);
nand U14427 (N_14427,N_13525,N_13996);
or U14428 (N_14428,N_13804,N_13501);
or U14429 (N_14429,N_13649,N_13634);
and U14430 (N_14430,N_13859,N_13816);
nand U14431 (N_14431,N_13948,N_13917);
xor U14432 (N_14432,N_13969,N_13709);
and U14433 (N_14433,N_13660,N_13645);
or U14434 (N_14434,N_13900,N_13968);
nor U14435 (N_14435,N_13630,N_13914);
and U14436 (N_14436,N_13745,N_13815);
nor U14437 (N_14437,N_13872,N_13646);
nor U14438 (N_14438,N_13742,N_13570);
xnor U14439 (N_14439,N_13999,N_13660);
and U14440 (N_14440,N_13813,N_13985);
nor U14441 (N_14441,N_13669,N_13649);
and U14442 (N_14442,N_13619,N_13840);
or U14443 (N_14443,N_13560,N_13656);
or U14444 (N_14444,N_13979,N_13539);
and U14445 (N_14445,N_13836,N_13844);
xor U14446 (N_14446,N_13762,N_13683);
or U14447 (N_14447,N_13965,N_13997);
and U14448 (N_14448,N_13878,N_13745);
nand U14449 (N_14449,N_13678,N_13560);
nor U14450 (N_14450,N_13507,N_13600);
nand U14451 (N_14451,N_13558,N_13813);
or U14452 (N_14452,N_13940,N_13730);
and U14453 (N_14453,N_13506,N_13861);
and U14454 (N_14454,N_13900,N_13532);
or U14455 (N_14455,N_13753,N_13591);
or U14456 (N_14456,N_13548,N_13593);
or U14457 (N_14457,N_13656,N_13744);
xnor U14458 (N_14458,N_13540,N_13793);
nand U14459 (N_14459,N_13816,N_13674);
or U14460 (N_14460,N_13890,N_13771);
nor U14461 (N_14461,N_13733,N_13788);
and U14462 (N_14462,N_13719,N_13834);
xnor U14463 (N_14463,N_13669,N_13633);
nor U14464 (N_14464,N_13910,N_13943);
and U14465 (N_14465,N_13727,N_13855);
nor U14466 (N_14466,N_13670,N_13881);
nand U14467 (N_14467,N_13930,N_13977);
or U14468 (N_14468,N_13684,N_13508);
or U14469 (N_14469,N_13522,N_13649);
xnor U14470 (N_14470,N_13535,N_13670);
or U14471 (N_14471,N_13641,N_13719);
xnor U14472 (N_14472,N_13725,N_13571);
nor U14473 (N_14473,N_13939,N_13902);
nor U14474 (N_14474,N_13751,N_13950);
or U14475 (N_14475,N_13797,N_13884);
or U14476 (N_14476,N_13845,N_13806);
nor U14477 (N_14477,N_13800,N_13923);
nor U14478 (N_14478,N_13792,N_13816);
and U14479 (N_14479,N_13622,N_13662);
nor U14480 (N_14480,N_13805,N_13874);
or U14481 (N_14481,N_13951,N_13843);
or U14482 (N_14482,N_13699,N_13585);
nor U14483 (N_14483,N_13801,N_13766);
xor U14484 (N_14484,N_13891,N_13661);
or U14485 (N_14485,N_13779,N_13946);
and U14486 (N_14486,N_13685,N_13562);
and U14487 (N_14487,N_13605,N_13771);
nor U14488 (N_14488,N_13555,N_13831);
xnor U14489 (N_14489,N_13912,N_13747);
xor U14490 (N_14490,N_13787,N_13794);
xnor U14491 (N_14491,N_13897,N_13777);
or U14492 (N_14492,N_13774,N_13926);
xnor U14493 (N_14493,N_13876,N_13526);
nand U14494 (N_14494,N_13538,N_13808);
nand U14495 (N_14495,N_13569,N_13846);
xor U14496 (N_14496,N_13662,N_13598);
nor U14497 (N_14497,N_13849,N_13800);
or U14498 (N_14498,N_13565,N_13597);
and U14499 (N_14499,N_13678,N_13621);
nand U14500 (N_14500,N_14210,N_14289);
and U14501 (N_14501,N_14452,N_14010);
xnor U14502 (N_14502,N_14440,N_14005);
or U14503 (N_14503,N_14132,N_14253);
xor U14504 (N_14504,N_14081,N_14110);
nand U14505 (N_14505,N_14209,N_14281);
nor U14506 (N_14506,N_14157,N_14406);
nand U14507 (N_14507,N_14314,N_14280);
or U14508 (N_14508,N_14198,N_14468);
and U14509 (N_14509,N_14290,N_14355);
or U14510 (N_14510,N_14238,N_14484);
nand U14511 (N_14511,N_14014,N_14218);
nor U14512 (N_14512,N_14271,N_14203);
and U14513 (N_14513,N_14294,N_14035);
or U14514 (N_14514,N_14177,N_14013);
and U14515 (N_14515,N_14404,N_14167);
and U14516 (N_14516,N_14023,N_14477);
or U14517 (N_14517,N_14220,N_14067);
nand U14518 (N_14518,N_14188,N_14058);
nand U14519 (N_14519,N_14375,N_14141);
nor U14520 (N_14520,N_14305,N_14117);
nand U14521 (N_14521,N_14265,N_14018);
nand U14522 (N_14522,N_14399,N_14287);
xnor U14523 (N_14523,N_14015,N_14046);
xnor U14524 (N_14524,N_14300,N_14261);
nand U14525 (N_14525,N_14017,N_14324);
xnor U14526 (N_14526,N_14411,N_14283);
nor U14527 (N_14527,N_14200,N_14487);
nor U14528 (N_14528,N_14488,N_14431);
or U14529 (N_14529,N_14070,N_14266);
or U14530 (N_14530,N_14219,N_14007);
xor U14531 (N_14531,N_14252,N_14096);
xnor U14532 (N_14532,N_14449,N_14093);
or U14533 (N_14533,N_14390,N_14293);
or U14534 (N_14534,N_14473,N_14426);
nor U14535 (N_14535,N_14403,N_14367);
xnor U14536 (N_14536,N_14376,N_14444);
nor U14537 (N_14537,N_14429,N_14085);
or U14538 (N_14538,N_14465,N_14088);
xnor U14539 (N_14539,N_14483,N_14105);
or U14540 (N_14540,N_14454,N_14469);
and U14541 (N_14541,N_14437,N_14194);
nor U14542 (N_14542,N_14301,N_14049);
nand U14543 (N_14543,N_14274,N_14201);
xor U14544 (N_14544,N_14226,N_14299);
nor U14545 (N_14545,N_14133,N_14224);
nand U14546 (N_14546,N_14215,N_14338);
or U14547 (N_14547,N_14378,N_14345);
xor U14548 (N_14548,N_14052,N_14165);
nor U14549 (N_14549,N_14244,N_14351);
nor U14550 (N_14550,N_14171,N_14024);
nand U14551 (N_14551,N_14340,N_14392);
nand U14552 (N_14552,N_14192,N_14292);
nand U14553 (N_14553,N_14172,N_14428);
nor U14554 (N_14554,N_14489,N_14108);
and U14555 (N_14555,N_14382,N_14059);
and U14556 (N_14556,N_14447,N_14222);
or U14557 (N_14557,N_14205,N_14317);
nor U14558 (N_14558,N_14051,N_14277);
nand U14559 (N_14559,N_14118,N_14459);
or U14560 (N_14560,N_14396,N_14464);
and U14561 (N_14561,N_14354,N_14229);
nor U14562 (N_14562,N_14400,N_14236);
or U14563 (N_14563,N_14125,N_14401);
xnor U14564 (N_14564,N_14490,N_14264);
xnor U14565 (N_14565,N_14311,N_14333);
nand U14566 (N_14566,N_14031,N_14098);
nor U14567 (N_14567,N_14328,N_14372);
or U14568 (N_14568,N_14159,N_14418);
nand U14569 (N_14569,N_14069,N_14421);
or U14570 (N_14570,N_14275,N_14021);
and U14571 (N_14571,N_14288,N_14457);
xor U14572 (N_14572,N_14416,N_14006);
nor U14573 (N_14573,N_14148,N_14255);
xor U14574 (N_14574,N_14258,N_14185);
nand U14575 (N_14575,N_14412,N_14267);
and U14576 (N_14576,N_14012,N_14455);
or U14577 (N_14577,N_14128,N_14458);
xnor U14578 (N_14578,N_14116,N_14291);
or U14579 (N_14579,N_14094,N_14028);
nor U14580 (N_14580,N_14388,N_14441);
xor U14581 (N_14581,N_14104,N_14425);
nand U14582 (N_14582,N_14214,N_14475);
nor U14583 (N_14583,N_14158,N_14086);
or U14584 (N_14584,N_14254,N_14410);
nand U14585 (N_14585,N_14415,N_14145);
and U14586 (N_14586,N_14498,N_14076);
xor U14587 (N_14587,N_14045,N_14217);
nor U14588 (N_14588,N_14270,N_14150);
xor U14589 (N_14589,N_14033,N_14335);
nand U14590 (N_14590,N_14466,N_14184);
nor U14591 (N_14591,N_14004,N_14161);
xor U14592 (N_14592,N_14334,N_14387);
and U14593 (N_14593,N_14307,N_14371);
and U14594 (N_14594,N_14246,N_14163);
nand U14595 (N_14595,N_14260,N_14155);
and U14596 (N_14596,N_14494,N_14446);
xnor U14597 (N_14597,N_14082,N_14089);
or U14598 (N_14598,N_14040,N_14496);
xnor U14599 (N_14599,N_14306,N_14499);
and U14600 (N_14600,N_14186,N_14336);
nand U14601 (N_14601,N_14002,N_14001);
or U14602 (N_14602,N_14420,N_14379);
and U14603 (N_14603,N_14233,N_14369);
or U14604 (N_14604,N_14039,N_14208);
or U14605 (N_14605,N_14124,N_14343);
nand U14606 (N_14606,N_14239,N_14330);
nor U14607 (N_14607,N_14251,N_14230);
nor U14608 (N_14608,N_14309,N_14385);
nand U14609 (N_14609,N_14269,N_14303);
or U14610 (N_14610,N_14072,N_14310);
nor U14611 (N_14611,N_14380,N_14140);
or U14612 (N_14612,N_14216,N_14199);
nand U14613 (N_14613,N_14029,N_14248);
and U14614 (N_14614,N_14383,N_14302);
or U14615 (N_14615,N_14176,N_14472);
and U14616 (N_14616,N_14478,N_14273);
xor U14617 (N_14617,N_14213,N_14022);
or U14618 (N_14618,N_14337,N_14249);
nor U14619 (N_14619,N_14471,N_14223);
xor U14620 (N_14620,N_14296,N_14268);
xnor U14621 (N_14621,N_14481,N_14180);
or U14622 (N_14622,N_14344,N_14057);
nand U14623 (N_14623,N_14139,N_14443);
or U14624 (N_14624,N_14111,N_14102);
xnor U14625 (N_14625,N_14331,N_14424);
nor U14626 (N_14626,N_14242,N_14342);
and U14627 (N_14627,N_14146,N_14231);
and U14628 (N_14628,N_14467,N_14099);
xor U14629 (N_14629,N_14181,N_14075);
or U14630 (N_14630,N_14065,N_14276);
or U14631 (N_14631,N_14027,N_14435);
xnor U14632 (N_14632,N_14136,N_14365);
nor U14633 (N_14633,N_14386,N_14134);
nor U14634 (N_14634,N_14092,N_14347);
and U14635 (N_14635,N_14063,N_14129);
and U14636 (N_14636,N_14361,N_14243);
xnor U14637 (N_14637,N_14329,N_14016);
xor U14638 (N_14638,N_14256,N_14346);
xor U14639 (N_14639,N_14316,N_14448);
nor U14640 (N_14640,N_14204,N_14189);
and U14641 (N_14641,N_14038,N_14056);
nand U14642 (N_14642,N_14112,N_14107);
or U14643 (N_14643,N_14060,N_14357);
nand U14644 (N_14644,N_14413,N_14087);
nand U14645 (N_14645,N_14197,N_14349);
or U14646 (N_14646,N_14362,N_14041);
or U14647 (N_14647,N_14393,N_14391);
xnor U14648 (N_14648,N_14234,N_14491);
xor U14649 (N_14649,N_14272,N_14325);
and U14650 (N_14650,N_14240,N_14263);
or U14651 (N_14651,N_14083,N_14257);
or U14652 (N_14652,N_14164,N_14373);
nor U14653 (N_14653,N_14245,N_14348);
and U14654 (N_14654,N_14127,N_14407);
xor U14655 (N_14655,N_14339,N_14154);
nor U14656 (N_14656,N_14166,N_14225);
xor U14657 (N_14657,N_14077,N_14320);
or U14658 (N_14658,N_14368,N_14438);
nand U14659 (N_14659,N_14241,N_14476);
nor U14660 (N_14660,N_14062,N_14323);
and U14661 (N_14661,N_14153,N_14008);
or U14662 (N_14662,N_14486,N_14054);
nand U14663 (N_14663,N_14235,N_14285);
nor U14664 (N_14664,N_14151,N_14169);
xor U14665 (N_14665,N_14363,N_14480);
nor U14666 (N_14666,N_14119,N_14011);
xor U14667 (N_14667,N_14482,N_14170);
or U14668 (N_14668,N_14389,N_14183);
and U14669 (N_14669,N_14460,N_14193);
nor U14670 (N_14670,N_14298,N_14034);
xnor U14671 (N_14671,N_14162,N_14114);
and U14672 (N_14672,N_14174,N_14326);
or U14673 (N_14673,N_14135,N_14071);
nor U14674 (N_14674,N_14147,N_14126);
or U14675 (N_14675,N_14073,N_14360);
or U14676 (N_14676,N_14179,N_14470);
and U14677 (N_14677,N_14453,N_14191);
nand U14678 (N_14678,N_14422,N_14282);
xnor U14679 (N_14679,N_14394,N_14398);
xnor U14680 (N_14680,N_14304,N_14123);
nor U14681 (N_14681,N_14079,N_14091);
xor U14682 (N_14682,N_14495,N_14278);
and U14683 (N_14683,N_14182,N_14374);
nand U14684 (N_14684,N_14284,N_14423);
and U14685 (N_14685,N_14211,N_14434);
xor U14686 (N_14686,N_14084,N_14436);
or U14687 (N_14687,N_14442,N_14395);
xnor U14688 (N_14688,N_14493,N_14120);
nand U14689 (N_14689,N_14417,N_14202);
xor U14690 (N_14690,N_14327,N_14318);
xnor U14691 (N_14691,N_14103,N_14456);
and U14692 (N_14692,N_14036,N_14462);
nand U14693 (N_14693,N_14350,N_14149);
and U14694 (N_14694,N_14101,N_14352);
and U14695 (N_14695,N_14143,N_14384);
and U14696 (N_14696,N_14356,N_14227);
and U14697 (N_14697,N_14364,N_14237);
nor U14698 (N_14698,N_14144,N_14190);
xnor U14699 (N_14699,N_14100,N_14195);
and U14700 (N_14700,N_14009,N_14321);
and U14701 (N_14701,N_14297,N_14232);
or U14702 (N_14702,N_14461,N_14152);
nand U14703 (N_14703,N_14131,N_14173);
and U14704 (N_14704,N_14050,N_14228);
xnor U14705 (N_14705,N_14212,N_14427);
nand U14706 (N_14706,N_14078,N_14207);
xnor U14707 (N_14707,N_14439,N_14295);
and U14708 (N_14708,N_14130,N_14402);
and U14709 (N_14709,N_14286,N_14479);
or U14710 (N_14710,N_14113,N_14221);
xnor U14711 (N_14711,N_14381,N_14095);
and U14712 (N_14712,N_14068,N_14122);
nor U14713 (N_14713,N_14097,N_14414);
nor U14714 (N_14714,N_14175,N_14168);
or U14715 (N_14715,N_14397,N_14322);
or U14716 (N_14716,N_14109,N_14451);
or U14717 (N_14717,N_14313,N_14156);
nor U14718 (N_14718,N_14474,N_14247);
and U14719 (N_14719,N_14030,N_14066);
xnor U14720 (N_14720,N_14121,N_14279);
or U14721 (N_14721,N_14259,N_14485);
xnor U14722 (N_14722,N_14138,N_14020);
nor U14723 (N_14723,N_14450,N_14206);
and U14724 (N_14724,N_14025,N_14312);
xor U14725 (N_14725,N_14003,N_14043);
nor U14726 (N_14726,N_14055,N_14000);
nand U14727 (N_14727,N_14080,N_14359);
nand U14728 (N_14728,N_14106,N_14366);
nor U14729 (N_14729,N_14178,N_14419);
or U14730 (N_14730,N_14196,N_14409);
xnor U14731 (N_14731,N_14044,N_14064);
xor U14732 (N_14732,N_14432,N_14160);
nand U14733 (N_14733,N_14463,N_14042);
or U14734 (N_14734,N_14370,N_14037);
nor U14735 (N_14735,N_14019,N_14315);
xor U14736 (N_14736,N_14137,N_14090);
xnor U14737 (N_14737,N_14492,N_14433);
nor U14738 (N_14738,N_14430,N_14262);
nand U14739 (N_14739,N_14250,N_14115);
nor U14740 (N_14740,N_14061,N_14053);
nor U14741 (N_14741,N_14074,N_14408);
or U14742 (N_14742,N_14319,N_14358);
xor U14743 (N_14743,N_14142,N_14445);
nand U14744 (N_14744,N_14341,N_14332);
xor U14745 (N_14745,N_14048,N_14026);
and U14746 (N_14746,N_14353,N_14497);
or U14747 (N_14747,N_14308,N_14377);
nand U14748 (N_14748,N_14405,N_14047);
xor U14749 (N_14749,N_14032,N_14187);
nand U14750 (N_14750,N_14000,N_14416);
nor U14751 (N_14751,N_14494,N_14334);
xor U14752 (N_14752,N_14408,N_14109);
nor U14753 (N_14753,N_14141,N_14422);
nor U14754 (N_14754,N_14234,N_14150);
xor U14755 (N_14755,N_14231,N_14458);
or U14756 (N_14756,N_14333,N_14002);
nor U14757 (N_14757,N_14253,N_14319);
nand U14758 (N_14758,N_14159,N_14161);
or U14759 (N_14759,N_14499,N_14200);
and U14760 (N_14760,N_14114,N_14171);
and U14761 (N_14761,N_14138,N_14028);
and U14762 (N_14762,N_14330,N_14085);
and U14763 (N_14763,N_14135,N_14187);
nor U14764 (N_14764,N_14257,N_14456);
and U14765 (N_14765,N_14201,N_14303);
nor U14766 (N_14766,N_14171,N_14011);
nand U14767 (N_14767,N_14348,N_14367);
nand U14768 (N_14768,N_14214,N_14194);
and U14769 (N_14769,N_14464,N_14193);
or U14770 (N_14770,N_14235,N_14237);
nor U14771 (N_14771,N_14341,N_14199);
xnor U14772 (N_14772,N_14357,N_14433);
xnor U14773 (N_14773,N_14223,N_14151);
xor U14774 (N_14774,N_14429,N_14301);
or U14775 (N_14775,N_14255,N_14469);
or U14776 (N_14776,N_14188,N_14165);
or U14777 (N_14777,N_14469,N_14133);
and U14778 (N_14778,N_14149,N_14003);
or U14779 (N_14779,N_14348,N_14338);
nand U14780 (N_14780,N_14242,N_14198);
and U14781 (N_14781,N_14352,N_14413);
nor U14782 (N_14782,N_14353,N_14286);
or U14783 (N_14783,N_14332,N_14026);
xnor U14784 (N_14784,N_14129,N_14159);
nor U14785 (N_14785,N_14452,N_14224);
or U14786 (N_14786,N_14257,N_14182);
nand U14787 (N_14787,N_14083,N_14346);
and U14788 (N_14788,N_14425,N_14292);
xnor U14789 (N_14789,N_14271,N_14342);
or U14790 (N_14790,N_14388,N_14239);
and U14791 (N_14791,N_14114,N_14128);
and U14792 (N_14792,N_14045,N_14279);
xor U14793 (N_14793,N_14056,N_14219);
and U14794 (N_14794,N_14007,N_14325);
nand U14795 (N_14795,N_14202,N_14183);
and U14796 (N_14796,N_14115,N_14305);
nand U14797 (N_14797,N_14420,N_14443);
nor U14798 (N_14798,N_14165,N_14261);
nand U14799 (N_14799,N_14237,N_14198);
nand U14800 (N_14800,N_14120,N_14354);
xor U14801 (N_14801,N_14147,N_14036);
or U14802 (N_14802,N_14396,N_14061);
and U14803 (N_14803,N_14368,N_14379);
nand U14804 (N_14804,N_14188,N_14450);
and U14805 (N_14805,N_14060,N_14276);
nor U14806 (N_14806,N_14086,N_14369);
xor U14807 (N_14807,N_14067,N_14212);
and U14808 (N_14808,N_14093,N_14152);
and U14809 (N_14809,N_14204,N_14080);
nor U14810 (N_14810,N_14234,N_14269);
or U14811 (N_14811,N_14094,N_14033);
or U14812 (N_14812,N_14164,N_14466);
and U14813 (N_14813,N_14229,N_14152);
or U14814 (N_14814,N_14130,N_14002);
and U14815 (N_14815,N_14047,N_14458);
nand U14816 (N_14816,N_14198,N_14269);
and U14817 (N_14817,N_14304,N_14248);
nand U14818 (N_14818,N_14339,N_14425);
nor U14819 (N_14819,N_14006,N_14109);
xor U14820 (N_14820,N_14300,N_14231);
nand U14821 (N_14821,N_14367,N_14227);
nor U14822 (N_14822,N_14208,N_14335);
xnor U14823 (N_14823,N_14310,N_14363);
and U14824 (N_14824,N_14496,N_14095);
xnor U14825 (N_14825,N_14223,N_14445);
and U14826 (N_14826,N_14204,N_14422);
nand U14827 (N_14827,N_14378,N_14270);
nor U14828 (N_14828,N_14281,N_14283);
or U14829 (N_14829,N_14112,N_14305);
nor U14830 (N_14830,N_14258,N_14427);
nand U14831 (N_14831,N_14104,N_14083);
and U14832 (N_14832,N_14276,N_14190);
and U14833 (N_14833,N_14209,N_14378);
or U14834 (N_14834,N_14148,N_14245);
nand U14835 (N_14835,N_14481,N_14457);
and U14836 (N_14836,N_14113,N_14238);
and U14837 (N_14837,N_14290,N_14025);
nand U14838 (N_14838,N_14023,N_14115);
or U14839 (N_14839,N_14348,N_14173);
or U14840 (N_14840,N_14142,N_14378);
nand U14841 (N_14841,N_14043,N_14079);
and U14842 (N_14842,N_14200,N_14251);
and U14843 (N_14843,N_14416,N_14011);
xor U14844 (N_14844,N_14256,N_14499);
nand U14845 (N_14845,N_14068,N_14470);
and U14846 (N_14846,N_14031,N_14004);
and U14847 (N_14847,N_14103,N_14043);
or U14848 (N_14848,N_14441,N_14121);
xnor U14849 (N_14849,N_14165,N_14437);
or U14850 (N_14850,N_14033,N_14158);
and U14851 (N_14851,N_14364,N_14478);
nand U14852 (N_14852,N_14058,N_14372);
or U14853 (N_14853,N_14338,N_14123);
and U14854 (N_14854,N_14189,N_14129);
nor U14855 (N_14855,N_14025,N_14320);
nand U14856 (N_14856,N_14363,N_14112);
xor U14857 (N_14857,N_14448,N_14089);
or U14858 (N_14858,N_14237,N_14165);
or U14859 (N_14859,N_14122,N_14367);
or U14860 (N_14860,N_14107,N_14062);
nand U14861 (N_14861,N_14265,N_14332);
xor U14862 (N_14862,N_14029,N_14469);
nor U14863 (N_14863,N_14231,N_14322);
xor U14864 (N_14864,N_14179,N_14209);
nor U14865 (N_14865,N_14205,N_14112);
or U14866 (N_14866,N_14084,N_14325);
nand U14867 (N_14867,N_14187,N_14383);
xor U14868 (N_14868,N_14141,N_14084);
or U14869 (N_14869,N_14231,N_14395);
nor U14870 (N_14870,N_14345,N_14038);
and U14871 (N_14871,N_14242,N_14284);
nor U14872 (N_14872,N_14118,N_14390);
xnor U14873 (N_14873,N_14111,N_14171);
nand U14874 (N_14874,N_14153,N_14333);
nor U14875 (N_14875,N_14434,N_14174);
xor U14876 (N_14876,N_14229,N_14250);
and U14877 (N_14877,N_14001,N_14085);
nand U14878 (N_14878,N_14097,N_14019);
nor U14879 (N_14879,N_14339,N_14443);
or U14880 (N_14880,N_14059,N_14198);
and U14881 (N_14881,N_14151,N_14247);
and U14882 (N_14882,N_14146,N_14453);
or U14883 (N_14883,N_14285,N_14447);
nand U14884 (N_14884,N_14261,N_14314);
nand U14885 (N_14885,N_14101,N_14110);
and U14886 (N_14886,N_14082,N_14123);
and U14887 (N_14887,N_14434,N_14338);
xnor U14888 (N_14888,N_14011,N_14408);
nor U14889 (N_14889,N_14436,N_14328);
and U14890 (N_14890,N_14380,N_14268);
and U14891 (N_14891,N_14488,N_14070);
nor U14892 (N_14892,N_14415,N_14200);
nor U14893 (N_14893,N_14311,N_14397);
nor U14894 (N_14894,N_14256,N_14355);
nand U14895 (N_14895,N_14002,N_14166);
nor U14896 (N_14896,N_14158,N_14325);
or U14897 (N_14897,N_14446,N_14390);
nor U14898 (N_14898,N_14264,N_14286);
nor U14899 (N_14899,N_14317,N_14401);
and U14900 (N_14900,N_14433,N_14053);
and U14901 (N_14901,N_14407,N_14028);
or U14902 (N_14902,N_14334,N_14225);
and U14903 (N_14903,N_14192,N_14373);
nor U14904 (N_14904,N_14205,N_14016);
xor U14905 (N_14905,N_14290,N_14401);
or U14906 (N_14906,N_14214,N_14156);
or U14907 (N_14907,N_14086,N_14132);
nand U14908 (N_14908,N_14288,N_14111);
and U14909 (N_14909,N_14475,N_14420);
nor U14910 (N_14910,N_14024,N_14223);
nand U14911 (N_14911,N_14360,N_14167);
and U14912 (N_14912,N_14365,N_14110);
nand U14913 (N_14913,N_14302,N_14351);
and U14914 (N_14914,N_14356,N_14364);
and U14915 (N_14915,N_14058,N_14158);
nor U14916 (N_14916,N_14365,N_14154);
and U14917 (N_14917,N_14414,N_14326);
xor U14918 (N_14918,N_14069,N_14031);
nand U14919 (N_14919,N_14168,N_14126);
nor U14920 (N_14920,N_14074,N_14238);
nand U14921 (N_14921,N_14459,N_14044);
or U14922 (N_14922,N_14054,N_14216);
nor U14923 (N_14923,N_14039,N_14426);
or U14924 (N_14924,N_14401,N_14321);
nand U14925 (N_14925,N_14480,N_14019);
and U14926 (N_14926,N_14402,N_14242);
xor U14927 (N_14927,N_14189,N_14260);
nand U14928 (N_14928,N_14042,N_14462);
and U14929 (N_14929,N_14440,N_14432);
xnor U14930 (N_14930,N_14061,N_14431);
and U14931 (N_14931,N_14061,N_14372);
and U14932 (N_14932,N_14036,N_14443);
or U14933 (N_14933,N_14353,N_14480);
or U14934 (N_14934,N_14340,N_14239);
or U14935 (N_14935,N_14002,N_14326);
nand U14936 (N_14936,N_14232,N_14105);
xnor U14937 (N_14937,N_14145,N_14242);
xor U14938 (N_14938,N_14161,N_14208);
xnor U14939 (N_14939,N_14229,N_14401);
xor U14940 (N_14940,N_14437,N_14198);
nand U14941 (N_14941,N_14399,N_14188);
and U14942 (N_14942,N_14224,N_14034);
xnor U14943 (N_14943,N_14411,N_14469);
nand U14944 (N_14944,N_14470,N_14187);
nor U14945 (N_14945,N_14343,N_14013);
or U14946 (N_14946,N_14183,N_14431);
or U14947 (N_14947,N_14340,N_14116);
or U14948 (N_14948,N_14415,N_14057);
nor U14949 (N_14949,N_14159,N_14169);
xnor U14950 (N_14950,N_14475,N_14216);
and U14951 (N_14951,N_14413,N_14025);
nor U14952 (N_14952,N_14130,N_14355);
and U14953 (N_14953,N_14303,N_14336);
and U14954 (N_14954,N_14417,N_14249);
and U14955 (N_14955,N_14249,N_14259);
nand U14956 (N_14956,N_14376,N_14075);
xnor U14957 (N_14957,N_14011,N_14041);
or U14958 (N_14958,N_14430,N_14181);
nor U14959 (N_14959,N_14216,N_14211);
xnor U14960 (N_14960,N_14489,N_14170);
nand U14961 (N_14961,N_14493,N_14362);
or U14962 (N_14962,N_14207,N_14408);
and U14963 (N_14963,N_14475,N_14295);
or U14964 (N_14964,N_14215,N_14000);
and U14965 (N_14965,N_14279,N_14391);
or U14966 (N_14966,N_14186,N_14130);
xor U14967 (N_14967,N_14124,N_14360);
nor U14968 (N_14968,N_14022,N_14100);
nor U14969 (N_14969,N_14241,N_14159);
nor U14970 (N_14970,N_14082,N_14282);
and U14971 (N_14971,N_14340,N_14359);
nand U14972 (N_14972,N_14067,N_14252);
nand U14973 (N_14973,N_14258,N_14340);
nor U14974 (N_14974,N_14295,N_14247);
or U14975 (N_14975,N_14147,N_14249);
nand U14976 (N_14976,N_14183,N_14265);
nand U14977 (N_14977,N_14177,N_14134);
nand U14978 (N_14978,N_14191,N_14427);
and U14979 (N_14979,N_14225,N_14285);
or U14980 (N_14980,N_14327,N_14044);
or U14981 (N_14981,N_14378,N_14139);
nor U14982 (N_14982,N_14459,N_14325);
nor U14983 (N_14983,N_14345,N_14287);
xnor U14984 (N_14984,N_14310,N_14286);
or U14985 (N_14985,N_14017,N_14458);
nor U14986 (N_14986,N_14447,N_14299);
nand U14987 (N_14987,N_14267,N_14031);
nor U14988 (N_14988,N_14117,N_14375);
or U14989 (N_14989,N_14378,N_14293);
nand U14990 (N_14990,N_14347,N_14014);
or U14991 (N_14991,N_14199,N_14206);
nand U14992 (N_14992,N_14437,N_14405);
nand U14993 (N_14993,N_14266,N_14316);
and U14994 (N_14994,N_14466,N_14285);
nor U14995 (N_14995,N_14272,N_14041);
xnor U14996 (N_14996,N_14397,N_14105);
xnor U14997 (N_14997,N_14463,N_14091);
nor U14998 (N_14998,N_14344,N_14067);
xor U14999 (N_14999,N_14306,N_14049);
nor U15000 (N_15000,N_14860,N_14974);
and U15001 (N_15001,N_14889,N_14983);
xor U15002 (N_15002,N_14547,N_14909);
or U15003 (N_15003,N_14811,N_14642);
nand U15004 (N_15004,N_14794,N_14644);
nand U15005 (N_15005,N_14548,N_14767);
xor U15006 (N_15006,N_14904,N_14741);
nor U15007 (N_15007,N_14653,N_14559);
xnor U15008 (N_15008,N_14978,N_14806);
or U15009 (N_15009,N_14919,N_14914);
nor U15010 (N_15010,N_14798,N_14938);
or U15011 (N_15011,N_14869,N_14501);
nand U15012 (N_15012,N_14527,N_14722);
and U15013 (N_15013,N_14640,N_14759);
xnor U15014 (N_15014,N_14577,N_14557);
and U15015 (N_15015,N_14606,N_14922);
and U15016 (N_15016,N_14701,N_14920);
nand U15017 (N_15017,N_14998,N_14778);
nor U15018 (N_15018,N_14967,N_14886);
or U15019 (N_15019,N_14768,N_14829);
nand U15020 (N_15020,N_14892,N_14815);
xnor U15021 (N_15021,N_14664,N_14776);
and U15022 (N_15022,N_14881,N_14990);
xnor U15023 (N_15023,N_14887,N_14666);
xor U15024 (N_15024,N_14962,N_14808);
or U15025 (N_15025,N_14697,N_14681);
xor U15026 (N_15026,N_14943,N_14911);
or U15027 (N_15027,N_14803,N_14634);
and U15028 (N_15028,N_14940,N_14894);
nand U15029 (N_15029,N_14582,N_14790);
and U15030 (N_15030,N_14639,N_14730);
nor U15031 (N_15031,N_14858,N_14927);
or U15032 (N_15032,N_14874,N_14515);
and U15033 (N_15033,N_14960,N_14952);
and U15034 (N_15034,N_14930,N_14752);
nor U15035 (N_15035,N_14826,N_14643);
or U15036 (N_15036,N_14864,N_14549);
xor U15037 (N_15037,N_14857,N_14706);
and U15038 (N_15038,N_14964,N_14901);
xor U15039 (N_15039,N_14529,N_14546);
or U15040 (N_15040,N_14777,N_14866);
and U15041 (N_15041,N_14812,N_14562);
nand U15042 (N_15042,N_14956,N_14840);
or U15043 (N_15043,N_14786,N_14635);
or U15044 (N_15044,N_14769,N_14797);
or U15045 (N_15045,N_14912,N_14539);
xor U15046 (N_15046,N_14800,N_14626);
and U15047 (N_15047,N_14550,N_14695);
or U15048 (N_15048,N_14804,N_14890);
nor U15049 (N_15049,N_14714,N_14718);
nand U15050 (N_15050,N_14856,N_14788);
and U15051 (N_15051,N_14760,N_14944);
and U15052 (N_15052,N_14824,N_14744);
nor U15053 (N_15053,N_14850,N_14791);
and U15054 (N_15054,N_14843,N_14727);
and U15055 (N_15055,N_14668,N_14523);
nand U15056 (N_15056,N_14963,N_14705);
or U15057 (N_15057,N_14957,N_14598);
nand U15058 (N_15058,N_14876,N_14817);
or U15059 (N_15059,N_14608,N_14721);
or U15060 (N_15060,N_14891,N_14870);
or U15061 (N_15061,N_14561,N_14970);
nor U15062 (N_15062,N_14540,N_14703);
nor U15063 (N_15063,N_14775,N_14878);
and U15064 (N_15064,N_14578,N_14558);
nor U15065 (N_15065,N_14787,N_14596);
nor U15066 (N_15066,N_14875,N_14810);
xnor U15067 (N_15067,N_14543,N_14765);
and U15068 (N_15068,N_14845,N_14923);
and U15069 (N_15069,N_14719,N_14672);
xor U15070 (N_15070,N_14616,N_14884);
nor U15071 (N_15071,N_14763,N_14696);
or U15072 (N_15072,N_14945,N_14575);
nand U15073 (N_15073,N_14942,N_14888);
and U15074 (N_15074,N_14902,N_14936);
and U15075 (N_15075,N_14819,N_14551);
nor U15076 (N_15076,N_14740,N_14896);
xor U15077 (N_15077,N_14537,N_14690);
xnor U15078 (N_15078,N_14764,N_14801);
and U15079 (N_15079,N_14620,N_14645);
nor U15080 (N_15080,N_14656,N_14841);
xnor U15081 (N_15081,N_14785,N_14906);
nand U15082 (N_15082,N_14599,N_14805);
or U15083 (N_15083,N_14822,N_14700);
xor U15084 (N_15084,N_14565,N_14855);
nor U15085 (N_15085,N_14683,N_14617);
and U15086 (N_15086,N_14795,N_14834);
and U15087 (N_15087,N_14746,N_14939);
xnor U15088 (N_15088,N_14580,N_14994);
xor U15089 (N_15089,N_14986,N_14519);
nor U15090 (N_15090,N_14848,N_14632);
and U15091 (N_15091,N_14508,N_14749);
and U15092 (N_15092,N_14615,N_14854);
and U15093 (N_15093,N_14569,N_14789);
and U15094 (N_15094,N_14979,N_14937);
and U15095 (N_15095,N_14553,N_14753);
nand U15096 (N_15096,N_14900,N_14574);
nand U15097 (N_15097,N_14882,N_14915);
and U15098 (N_15098,N_14851,N_14755);
and U15099 (N_15099,N_14799,N_14959);
nor U15100 (N_15100,N_14717,N_14732);
nand U15101 (N_15101,N_14720,N_14657);
and U15102 (N_15102,N_14835,N_14908);
or U15103 (N_15103,N_14742,N_14627);
nand U15104 (N_15104,N_14977,N_14989);
or U15105 (N_15105,N_14600,N_14509);
or U15106 (N_15106,N_14512,N_14506);
xor U15107 (N_15107,N_14623,N_14981);
and U15108 (N_15108,N_14552,N_14507);
xnor U15109 (N_15109,N_14674,N_14893);
xnor U15110 (N_15110,N_14916,N_14587);
nand U15111 (N_15111,N_14663,N_14739);
or U15112 (N_15112,N_14877,N_14976);
nor U15113 (N_15113,N_14522,N_14682);
nand U15114 (N_15114,N_14505,N_14511);
nand U15115 (N_15115,N_14712,N_14583);
nor U15116 (N_15116,N_14535,N_14796);
and U15117 (N_15117,N_14734,N_14648);
xor U15118 (N_15118,N_14932,N_14733);
nand U15119 (N_15119,N_14605,N_14542);
and U15120 (N_15120,N_14560,N_14715);
or U15121 (N_15121,N_14868,N_14729);
and U15122 (N_15122,N_14530,N_14832);
and U15123 (N_15123,N_14638,N_14883);
or U15124 (N_15124,N_14594,N_14590);
and U15125 (N_15125,N_14567,N_14670);
nand U15126 (N_15126,N_14984,N_14846);
nand U15127 (N_15127,N_14947,N_14871);
or U15128 (N_15128,N_14757,N_14807);
or U15129 (N_15129,N_14809,N_14693);
xnor U15130 (N_15130,N_14968,N_14735);
xnor U15131 (N_15131,N_14711,N_14602);
and U15132 (N_15132,N_14743,N_14774);
and U15133 (N_15133,N_14779,N_14581);
xnor U15134 (N_15134,N_14636,N_14750);
xor U15135 (N_15135,N_14773,N_14844);
nand U15136 (N_15136,N_14633,N_14934);
and U15137 (N_15137,N_14646,N_14500);
nor U15138 (N_15138,N_14710,N_14597);
and U15139 (N_15139,N_14667,N_14905);
or U15140 (N_15140,N_14589,N_14708);
and U15141 (N_15141,N_14953,N_14526);
nand U15142 (N_15142,N_14641,N_14991);
or U15143 (N_15143,N_14736,N_14903);
nor U15144 (N_15144,N_14737,N_14525);
nor U15145 (N_15145,N_14770,N_14725);
or U15146 (N_15146,N_14879,N_14745);
or U15147 (N_15147,N_14849,N_14781);
xor U15148 (N_15148,N_14772,N_14709);
and U15149 (N_15149,N_14658,N_14830);
xnor U15150 (N_15150,N_14756,N_14687);
or U15151 (N_15151,N_14685,N_14669);
nor U15152 (N_15152,N_14595,N_14880);
and U15153 (N_15153,N_14992,N_14586);
nand U15154 (N_15154,N_14630,N_14649);
and U15155 (N_15155,N_14662,N_14813);
nand U15156 (N_15156,N_14655,N_14654);
nor U15157 (N_15157,N_14973,N_14514);
nor U15158 (N_15158,N_14584,N_14573);
nand U15159 (N_15159,N_14782,N_14766);
and U15160 (N_15160,N_14895,N_14647);
or U15161 (N_15161,N_14613,N_14524);
and U15162 (N_15162,N_14593,N_14694);
or U15163 (N_15163,N_14861,N_14929);
xor U15164 (N_15164,N_14702,N_14571);
nand U15165 (N_15165,N_14771,N_14686);
or U15166 (N_15166,N_14821,N_14603);
nor U15167 (N_15167,N_14554,N_14585);
or U15168 (N_15168,N_14564,N_14521);
or U15169 (N_15169,N_14975,N_14762);
nor U15170 (N_15170,N_14680,N_14999);
nand U15171 (N_15171,N_14954,N_14637);
nor U15172 (N_15172,N_14997,N_14847);
or U15173 (N_15173,N_14955,N_14748);
xnor U15174 (N_15174,N_14754,N_14533);
and U15175 (N_15175,N_14622,N_14897);
xor U15176 (N_15176,N_14652,N_14814);
nor U15177 (N_15177,N_14541,N_14780);
and U15178 (N_15178,N_14572,N_14607);
and U15179 (N_15179,N_14563,N_14873);
and U15180 (N_15180,N_14924,N_14833);
nor U15181 (N_15181,N_14579,N_14917);
xor U15182 (N_15182,N_14863,N_14982);
nand U15183 (N_15183,N_14570,N_14661);
nor U15184 (N_15184,N_14950,N_14628);
or U15185 (N_15185,N_14842,N_14513);
or U15186 (N_15186,N_14610,N_14621);
xor U15187 (N_15187,N_14928,N_14671);
and U15188 (N_15188,N_14951,N_14996);
or U15189 (N_15189,N_14926,N_14612);
xnor U15190 (N_15190,N_14831,N_14629);
nor U15191 (N_15191,N_14918,N_14684);
and U15192 (N_15192,N_14948,N_14704);
nor U15193 (N_15193,N_14961,N_14601);
nor U15194 (N_15194,N_14836,N_14816);
xnor U15195 (N_15195,N_14837,N_14985);
and U15196 (N_15196,N_14913,N_14531);
or U15197 (N_15197,N_14673,N_14679);
and U15198 (N_15198,N_14969,N_14827);
or U15199 (N_15199,N_14698,N_14910);
nand U15200 (N_15200,N_14619,N_14716);
nor U15201 (N_15201,N_14958,N_14988);
xnor U15202 (N_15202,N_14689,N_14591);
xnor U15203 (N_15203,N_14872,N_14907);
or U15204 (N_15204,N_14568,N_14818);
xor U15205 (N_15205,N_14520,N_14823);
xor U15206 (N_15206,N_14931,N_14972);
or U15207 (N_15207,N_14536,N_14802);
nand U15208 (N_15208,N_14691,N_14899);
nor U15209 (N_15209,N_14987,N_14751);
or U15210 (N_15210,N_14933,N_14865);
xnor U15211 (N_15211,N_14838,N_14971);
nand U15212 (N_15212,N_14935,N_14604);
and U15213 (N_15213,N_14761,N_14545);
or U15214 (N_15214,N_14980,N_14576);
nand U15215 (N_15215,N_14665,N_14949);
nor U15216 (N_15216,N_14783,N_14692);
nand U15217 (N_15217,N_14517,N_14614);
or U15218 (N_15218,N_14544,N_14707);
or U15219 (N_15219,N_14713,N_14625);
or U15220 (N_15220,N_14618,N_14502);
nor U15221 (N_15221,N_14966,N_14995);
or U15222 (N_15222,N_14867,N_14588);
nand U15223 (N_15223,N_14859,N_14898);
xor U15224 (N_15224,N_14504,N_14946);
and U15225 (N_15225,N_14675,N_14747);
nor U15226 (N_15226,N_14839,N_14728);
nand U15227 (N_15227,N_14885,N_14677);
nor U15228 (N_15228,N_14828,N_14793);
and U15229 (N_15229,N_14965,N_14538);
xnor U15230 (N_15230,N_14738,N_14516);
and U15231 (N_15231,N_14820,N_14503);
and U15232 (N_15232,N_14659,N_14731);
and U15233 (N_15233,N_14678,N_14784);
and U15234 (N_15234,N_14518,N_14792);
xor U15235 (N_15235,N_14724,N_14592);
nand U15236 (N_15236,N_14853,N_14528);
or U15237 (N_15237,N_14825,N_14941);
or U15238 (N_15238,N_14852,N_14631);
nor U15239 (N_15239,N_14534,N_14566);
or U15240 (N_15240,N_14555,N_14609);
or U15241 (N_15241,N_14532,N_14650);
nor U15242 (N_15242,N_14921,N_14510);
nor U15243 (N_15243,N_14624,N_14556);
xnor U15244 (N_15244,N_14688,N_14723);
and U15245 (N_15245,N_14611,N_14925);
or U15246 (N_15246,N_14862,N_14726);
or U15247 (N_15247,N_14660,N_14651);
and U15248 (N_15248,N_14993,N_14676);
or U15249 (N_15249,N_14758,N_14699);
and U15250 (N_15250,N_14630,N_14786);
nor U15251 (N_15251,N_14924,N_14744);
nor U15252 (N_15252,N_14635,N_14732);
nand U15253 (N_15253,N_14764,N_14580);
nand U15254 (N_15254,N_14838,N_14841);
nand U15255 (N_15255,N_14698,N_14671);
and U15256 (N_15256,N_14618,N_14532);
and U15257 (N_15257,N_14601,N_14855);
and U15258 (N_15258,N_14664,N_14545);
nand U15259 (N_15259,N_14740,N_14978);
xnor U15260 (N_15260,N_14868,N_14682);
nor U15261 (N_15261,N_14510,N_14981);
nand U15262 (N_15262,N_14576,N_14841);
or U15263 (N_15263,N_14591,N_14974);
nand U15264 (N_15264,N_14846,N_14863);
nor U15265 (N_15265,N_14994,N_14583);
xor U15266 (N_15266,N_14520,N_14915);
nand U15267 (N_15267,N_14558,N_14598);
and U15268 (N_15268,N_14677,N_14990);
nand U15269 (N_15269,N_14777,N_14966);
and U15270 (N_15270,N_14595,N_14937);
and U15271 (N_15271,N_14547,N_14634);
and U15272 (N_15272,N_14516,N_14812);
nor U15273 (N_15273,N_14789,N_14570);
or U15274 (N_15274,N_14923,N_14776);
nand U15275 (N_15275,N_14669,N_14895);
or U15276 (N_15276,N_14943,N_14778);
nor U15277 (N_15277,N_14857,N_14624);
or U15278 (N_15278,N_14721,N_14874);
nor U15279 (N_15279,N_14541,N_14572);
nor U15280 (N_15280,N_14870,N_14619);
xnor U15281 (N_15281,N_14769,N_14891);
and U15282 (N_15282,N_14518,N_14858);
or U15283 (N_15283,N_14534,N_14892);
nand U15284 (N_15284,N_14588,N_14562);
nand U15285 (N_15285,N_14808,N_14951);
and U15286 (N_15286,N_14527,N_14861);
or U15287 (N_15287,N_14908,N_14684);
nor U15288 (N_15288,N_14569,N_14717);
nand U15289 (N_15289,N_14582,N_14575);
or U15290 (N_15290,N_14502,N_14530);
or U15291 (N_15291,N_14679,N_14925);
and U15292 (N_15292,N_14984,N_14541);
or U15293 (N_15293,N_14557,N_14747);
and U15294 (N_15294,N_14981,N_14908);
nor U15295 (N_15295,N_14716,N_14760);
xor U15296 (N_15296,N_14565,N_14612);
xor U15297 (N_15297,N_14691,N_14962);
or U15298 (N_15298,N_14854,N_14697);
nand U15299 (N_15299,N_14578,N_14756);
xnor U15300 (N_15300,N_14653,N_14548);
nand U15301 (N_15301,N_14601,N_14726);
nor U15302 (N_15302,N_14501,N_14529);
nand U15303 (N_15303,N_14927,N_14511);
nand U15304 (N_15304,N_14760,N_14663);
nand U15305 (N_15305,N_14824,N_14589);
nor U15306 (N_15306,N_14860,N_14901);
or U15307 (N_15307,N_14885,N_14635);
and U15308 (N_15308,N_14631,N_14587);
xnor U15309 (N_15309,N_14760,N_14778);
nor U15310 (N_15310,N_14860,N_14576);
nor U15311 (N_15311,N_14860,N_14631);
and U15312 (N_15312,N_14885,N_14889);
nand U15313 (N_15313,N_14712,N_14679);
nand U15314 (N_15314,N_14955,N_14904);
nand U15315 (N_15315,N_14719,N_14815);
or U15316 (N_15316,N_14852,N_14875);
and U15317 (N_15317,N_14717,N_14792);
nand U15318 (N_15318,N_14675,N_14887);
xnor U15319 (N_15319,N_14874,N_14989);
xnor U15320 (N_15320,N_14674,N_14774);
xnor U15321 (N_15321,N_14852,N_14508);
nand U15322 (N_15322,N_14890,N_14694);
nor U15323 (N_15323,N_14703,N_14743);
nand U15324 (N_15324,N_14770,N_14629);
xnor U15325 (N_15325,N_14811,N_14849);
xor U15326 (N_15326,N_14753,N_14649);
or U15327 (N_15327,N_14515,N_14544);
nor U15328 (N_15328,N_14782,N_14628);
xnor U15329 (N_15329,N_14527,N_14603);
nor U15330 (N_15330,N_14948,N_14879);
nor U15331 (N_15331,N_14751,N_14654);
or U15332 (N_15332,N_14980,N_14658);
nand U15333 (N_15333,N_14818,N_14968);
or U15334 (N_15334,N_14838,N_14751);
nand U15335 (N_15335,N_14862,N_14659);
or U15336 (N_15336,N_14927,N_14521);
nand U15337 (N_15337,N_14522,N_14898);
and U15338 (N_15338,N_14850,N_14534);
or U15339 (N_15339,N_14560,N_14568);
nand U15340 (N_15340,N_14717,N_14678);
and U15341 (N_15341,N_14576,N_14848);
nor U15342 (N_15342,N_14823,N_14810);
and U15343 (N_15343,N_14634,N_14990);
xor U15344 (N_15344,N_14673,N_14792);
xnor U15345 (N_15345,N_14585,N_14787);
and U15346 (N_15346,N_14984,N_14947);
and U15347 (N_15347,N_14805,N_14593);
nand U15348 (N_15348,N_14964,N_14937);
or U15349 (N_15349,N_14519,N_14958);
nand U15350 (N_15350,N_14752,N_14721);
nand U15351 (N_15351,N_14559,N_14898);
or U15352 (N_15352,N_14759,N_14502);
nand U15353 (N_15353,N_14698,N_14781);
and U15354 (N_15354,N_14873,N_14741);
and U15355 (N_15355,N_14521,N_14589);
nor U15356 (N_15356,N_14771,N_14920);
and U15357 (N_15357,N_14963,N_14946);
and U15358 (N_15358,N_14941,N_14611);
nand U15359 (N_15359,N_14504,N_14749);
xnor U15360 (N_15360,N_14614,N_14961);
or U15361 (N_15361,N_14651,N_14948);
and U15362 (N_15362,N_14859,N_14740);
nor U15363 (N_15363,N_14719,N_14874);
xor U15364 (N_15364,N_14965,N_14994);
and U15365 (N_15365,N_14502,N_14882);
nor U15366 (N_15366,N_14672,N_14999);
or U15367 (N_15367,N_14695,N_14987);
nand U15368 (N_15368,N_14956,N_14762);
and U15369 (N_15369,N_14644,N_14675);
xnor U15370 (N_15370,N_14586,N_14999);
nand U15371 (N_15371,N_14897,N_14996);
and U15372 (N_15372,N_14935,N_14671);
xor U15373 (N_15373,N_14588,N_14915);
nor U15374 (N_15374,N_14645,N_14664);
nand U15375 (N_15375,N_14675,N_14955);
and U15376 (N_15376,N_14867,N_14845);
nor U15377 (N_15377,N_14800,N_14720);
nor U15378 (N_15378,N_14797,N_14585);
xor U15379 (N_15379,N_14807,N_14591);
or U15380 (N_15380,N_14602,N_14508);
or U15381 (N_15381,N_14763,N_14511);
xor U15382 (N_15382,N_14784,N_14551);
xnor U15383 (N_15383,N_14507,N_14666);
or U15384 (N_15384,N_14987,N_14734);
and U15385 (N_15385,N_14711,N_14967);
and U15386 (N_15386,N_14929,N_14892);
or U15387 (N_15387,N_14568,N_14863);
and U15388 (N_15388,N_14621,N_14966);
or U15389 (N_15389,N_14850,N_14651);
xnor U15390 (N_15390,N_14928,N_14516);
or U15391 (N_15391,N_14608,N_14885);
or U15392 (N_15392,N_14797,N_14805);
or U15393 (N_15393,N_14730,N_14612);
nor U15394 (N_15394,N_14798,N_14652);
nand U15395 (N_15395,N_14692,N_14691);
and U15396 (N_15396,N_14689,N_14618);
xor U15397 (N_15397,N_14814,N_14970);
nor U15398 (N_15398,N_14663,N_14960);
and U15399 (N_15399,N_14972,N_14653);
or U15400 (N_15400,N_14978,N_14761);
nand U15401 (N_15401,N_14879,N_14651);
xor U15402 (N_15402,N_14996,N_14547);
xnor U15403 (N_15403,N_14809,N_14671);
xnor U15404 (N_15404,N_14583,N_14532);
xnor U15405 (N_15405,N_14671,N_14868);
nor U15406 (N_15406,N_14737,N_14780);
and U15407 (N_15407,N_14645,N_14991);
xor U15408 (N_15408,N_14781,N_14801);
nand U15409 (N_15409,N_14937,N_14532);
and U15410 (N_15410,N_14530,N_14961);
nor U15411 (N_15411,N_14926,N_14595);
and U15412 (N_15412,N_14793,N_14583);
or U15413 (N_15413,N_14521,N_14528);
and U15414 (N_15414,N_14713,N_14894);
nor U15415 (N_15415,N_14948,N_14527);
nand U15416 (N_15416,N_14539,N_14685);
nand U15417 (N_15417,N_14753,N_14578);
or U15418 (N_15418,N_14563,N_14894);
or U15419 (N_15419,N_14817,N_14681);
nand U15420 (N_15420,N_14945,N_14861);
nand U15421 (N_15421,N_14661,N_14682);
nor U15422 (N_15422,N_14501,N_14833);
xor U15423 (N_15423,N_14968,N_14984);
xnor U15424 (N_15424,N_14731,N_14808);
and U15425 (N_15425,N_14708,N_14765);
or U15426 (N_15426,N_14995,N_14877);
nand U15427 (N_15427,N_14828,N_14775);
nand U15428 (N_15428,N_14718,N_14962);
xor U15429 (N_15429,N_14683,N_14932);
or U15430 (N_15430,N_14891,N_14582);
nor U15431 (N_15431,N_14813,N_14741);
or U15432 (N_15432,N_14834,N_14759);
or U15433 (N_15433,N_14686,N_14513);
xor U15434 (N_15434,N_14528,N_14962);
and U15435 (N_15435,N_14510,N_14571);
and U15436 (N_15436,N_14701,N_14713);
nand U15437 (N_15437,N_14619,N_14671);
or U15438 (N_15438,N_14617,N_14872);
nor U15439 (N_15439,N_14569,N_14500);
nand U15440 (N_15440,N_14645,N_14955);
xnor U15441 (N_15441,N_14546,N_14822);
xor U15442 (N_15442,N_14642,N_14828);
and U15443 (N_15443,N_14737,N_14577);
or U15444 (N_15444,N_14655,N_14775);
or U15445 (N_15445,N_14645,N_14931);
nand U15446 (N_15446,N_14528,N_14737);
xnor U15447 (N_15447,N_14850,N_14961);
or U15448 (N_15448,N_14832,N_14821);
and U15449 (N_15449,N_14920,N_14636);
xor U15450 (N_15450,N_14845,N_14908);
and U15451 (N_15451,N_14946,N_14784);
xor U15452 (N_15452,N_14640,N_14794);
nand U15453 (N_15453,N_14956,N_14542);
nand U15454 (N_15454,N_14754,N_14770);
or U15455 (N_15455,N_14794,N_14953);
xor U15456 (N_15456,N_14933,N_14506);
nor U15457 (N_15457,N_14730,N_14744);
and U15458 (N_15458,N_14753,N_14907);
xnor U15459 (N_15459,N_14564,N_14523);
nand U15460 (N_15460,N_14500,N_14600);
nand U15461 (N_15461,N_14774,N_14540);
and U15462 (N_15462,N_14807,N_14577);
and U15463 (N_15463,N_14715,N_14902);
nor U15464 (N_15464,N_14507,N_14550);
nor U15465 (N_15465,N_14858,N_14923);
nor U15466 (N_15466,N_14590,N_14598);
nor U15467 (N_15467,N_14783,N_14958);
nor U15468 (N_15468,N_14636,N_14835);
nor U15469 (N_15469,N_14930,N_14632);
xnor U15470 (N_15470,N_14774,N_14798);
xor U15471 (N_15471,N_14927,N_14538);
nor U15472 (N_15472,N_14968,N_14728);
nand U15473 (N_15473,N_14776,N_14613);
or U15474 (N_15474,N_14950,N_14691);
and U15475 (N_15475,N_14528,N_14690);
and U15476 (N_15476,N_14853,N_14991);
and U15477 (N_15477,N_14517,N_14743);
or U15478 (N_15478,N_14838,N_14551);
and U15479 (N_15479,N_14757,N_14911);
and U15480 (N_15480,N_14814,N_14958);
nor U15481 (N_15481,N_14748,N_14711);
nor U15482 (N_15482,N_14847,N_14763);
xor U15483 (N_15483,N_14991,N_14771);
nand U15484 (N_15484,N_14697,N_14757);
nor U15485 (N_15485,N_14767,N_14826);
xnor U15486 (N_15486,N_14931,N_14737);
nor U15487 (N_15487,N_14540,N_14937);
nand U15488 (N_15488,N_14917,N_14594);
and U15489 (N_15489,N_14975,N_14960);
nor U15490 (N_15490,N_14574,N_14820);
nor U15491 (N_15491,N_14836,N_14734);
nor U15492 (N_15492,N_14655,N_14964);
xnor U15493 (N_15493,N_14556,N_14839);
nand U15494 (N_15494,N_14808,N_14803);
xor U15495 (N_15495,N_14510,N_14602);
nand U15496 (N_15496,N_14823,N_14995);
xor U15497 (N_15497,N_14759,N_14724);
or U15498 (N_15498,N_14856,N_14814);
or U15499 (N_15499,N_14991,N_14987);
and U15500 (N_15500,N_15440,N_15072);
and U15501 (N_15501,N_15117,N_15376);
or U15502 (N_15502,N_15348,N_15118);
nor U15503 (N_15503,N_15341,N_15446);
or U15504 (N_15504,N_15154,N_15041);
nor U15505 (N_15505,N_15488,N_15207);
xor U15506 (N_15506,N_15085,N_15024);
and U15507 (N_15507,N_15125,N_15356);
or U15508 (N_15508,N_15051,N_15453);
nor U15509 (N_15509,N_15156,N_15296);
and U15510 (N_15510,N_15078,N_15475);
xor U15511 (N_15511,N_15236,N_15160);
xnor U15512 (N_15512,N_15365,N_15015);
or U15513 (N_15513,N_15326,N_15169);
xor U15514 (N_15514,N_15403,N_15439);
nor U15515 (N_15515,N_15380,N_15077);
nor U15516 (N_15516,N_15094,N_15484);
and U15517 (N_15517,N_15229,N_15412);
nor U15518 (N_15518,N_15227,N_15260);
and U15519 (N_15519,N_15174,N_15026);
or U15520 (N_15520,N_15496,N_15471);
nand U15521 (N_15521,N_15009,N_15131);
and U15522 (N_15522,N_15478,N_15287);
nand U15523 (N_15523,N_15003,N_15122);
nor U15524 (N_15524,N_15144,N_15007);
xor U15525 (N_15525,N_15302,N_15162);
xor U15526 (N_15526,N_15237,N_15235);
nand U15527 (N_15527,N_15418,N_15383);
xnor U15528 (N_15528,N_15479,N_15048);
or U15529 (N_15529,N_15275,N_15220);
xor U15530 (N_15530,N_15022,N_15395);
xnor U15531 (N_15531,N_15212,N_15289);
and U15532 (N_15532,N_15301,N_15385);
nand U15533 (N_15533,N_15194,N_15422);
and U15534 (N_15534,N_15210,N_15185);
or U15535 (N_15535,N_15037,N_15001);
and U15536 (N_15536,N_15043,N_15280);
nor U15537 (N_15537,N_15164,N_15355);
nor U15538 (N_15538,N_15312,N_15066);
xnor U15539 (N_15539,N_15253,N_15276);
nor U15540 (N_15540,N_15406,N_15255);
nor U15541 (N_15541,N_15433,N_15423);
xnor U15542 (N_15542,N_15106,N_15054);
nor U15543 (N_15543,N_15069,N_15483);
and U15544 (N_15544,N_15163,N_15278);
nand U15545 (N_15545,N_15334,N_15092);
or U15546 (N_15546,N_15145,N_15062);
and U15547 (N_15547,N_15161,N_15130);
nor U15548 (N_15548,N_15112,N_15076);
xor U15549 (N_15549,N_15120,N_15384);
or U15550 (N_15550,N_15300,N_15434);
or U15551 (N_15551,N_15338,N_15485);
xnor U15552 (N_15552,N_15225,N_15052);
and U15553 (N_15553,N_15084,N_15230);
nand U15554 (N_15554,N_15082,N_15240);
and U15555 (N_15555,N_15400,N_15409);
nor U15556 (N_15556,N_15201,N_15399);
or U15557 (N_15557,N_15294,N_15187);
nor U15558 (N_15558,N_15397,N_15272);
or U15559 (N_15559,N_15067,N_15426);
and U15560 (N_15560,N_15215,N_15004);
nand U15561 (N_15561,N_15298,N_15257);
nand U15562 (N_15562,N_15316,N_15079);
nor U15563 (N_15563,N_15452,N_15467);
and U15564 (N_15564,N_15482,N_15317);
or U15565 (N_15565,N_15027,N_15039);
xnor U15566 (N_15566,N_15168,N_15088);
or U15567 (N_15567,N_15497,N_15038);
nand U15568 (N_15568,N_15116,N_15103);
and U15569 (N_15569,N_15345,N_15408);
and U15570 (N_15570,N_15029,N_15391);
or U15571 (N_15571,N_15310,N_15304);
xnor U15572 (N_15572,N_15273,N_15492);
xor U15573 (N_15573,N_15315,N_15241);
nor U15574 (N_15574,N_15013,N_15340);
nand U15575 (N_15575,N_15068,N_15246);
and U15576 (N_15576,N_15353,N_15364);
xor U15577 (N_15577,N_15321,N_15374);
nor U15578 (N_15578,N_15286,N_15336);
nor U15579 (N_15579,N_15019,N_15307);
nor U15580 (N_15580,N_15173,N_15424);
nor U15581 (N_15581,N_15233,N_15167);
xor U15582 (N_15582,N_15073,N_15093);
and U15583 (N_15583,N_15295,N_15098);
and U15584 (N_15584,N_15271,N_15104);
xor U15585 (N_15585,N_15010,N_15137);
or U15586 (N_15586,N_15197,N_15059);
or U15587 (N_15587,N_15363,N_15318);
or U15588 (N_15588,N_15299,N_15204);
and U15589 (N_15589,N_15107,N_15309);
or U15590 (N_15590,N_15128,N_15105);
nand U15591 (N_15591,N_15176,N_15211);
and U15592 (N_15592,N_15311,N_15214);
nor U15593 (N_15593,N_15328,N_15244);
and U15594 (N_15594,N_15420,N_15110);
nor U15595 (N_15595,N_15046,N_15159);
and U15596 (N_15596,N_15460,N_15186);
nor U15597 (N_15597,N_15429,N_15404);
nand U15598 (N_15598,N_15008,N_15249);
xnor U15599 (N_15599,N_15322,N_15323);
xnor U15600 (N_15600,N_15021,N_15189);
or U15601 (N_15601,N_15443,N_15431);
or U15602 (N_15602,N_15113,N_15126);
xor U15603 (N_15603,N_15480,N_15080);
nand U15604 (N_15604,N_15421,N_15075);
and U15605 (N_15605,N_15277,N_15147);
nor U15606 (N_15606,N_15196,N_15123);
and U15607 (N_15607,N_15011,N_15361);
nor U15608 (N_15608,N_15158,N_15442);
nor U15609 (N_15609,N_15306,N_15358);
and U15610 (N_15610,N_15266,N_15115);
and U15611 (N_15611,N_15202,N_15370);
or U15612 (N_15612,N_15382,N_15091);
nor U15613 (N_15613,N_15350,N_15329);
nand U15614 (N_15614,N_15044,N_15034);
nor U15615 (N_15615,N_15148,N_15258);
xor U15616 (N_15616,N_15047,N_15221);
nand U15617 (N_15617,N_15245,N_15477);
nor U15618 (N_15618,N_15297,N_15468);
or U15619 (N_15619,N_15136,N_15050);
nand U15620 (N_15620,N_15247,N_15184);
and U15621 (N_15621,N_15143,N_15057);
xnor U15622 (N_15622,N_15405,N_15188);
nand U15623 (N_15623,N_15209,N_15064);
nor U15624 (N_15624,N_15121,N_15149);
nor U15625 (N_15625,N_15461,N_15430);
nand U15626 (N_15626,N_15371,N_15058);
xnor U15627 (N_15627,N_15360,N_15462);
xnor U15628 (N_15628,N_15263,N_15135);
xor U15629 (N_15629,N_15081,N_15331);
nor U15630 (N_15630,N_15285,N_15179);
nor U15631 (N_15631,N_15109,N_15252);
and U15632 (N_15632,N_15262,N_15055);
and U15633 (N_15633,N_15265,N_15012);
nand U15634 (N_15634,N_15219,N_15320);
or U15635 (N_15635,N_15427,N_15466);
nor U15636 (N_15636,N_15335,N_15448);
and U15637 (N_15637,N_15213,N_15359);
xnor U15638 (N_15638,N_15469,N_15387);
or U15639 (N_15639,N_15239,N_15119);
xor U15640 (N_15640,N_15146,N_15472);
and U15641 (N_15641,N_15234,N_15206);
nor U15642 (N_15642,N_15305,N_15319);
xnor U15643 (N_15643,N_15375,N_15166);
nand U15644 (N_15644,N_15449,N_15268);
nand U15645 (N_15645,N_15362,N_15368);
nor U15646 (N_15646,N_15254,N_15099);
and U15647 (N_15647,N_15413,N_15463);
and U15648 (N_15648,N_15416,N_15170);
nor U15649 (N_15649,N_15308,N_15250);
nor U15650 (N_15650,N_15401,N_15325);
xnor U15651 (N_15651,N_15017,N_15398);
xor U15652 (N_15652,N_15490,N_15417);
nand U15653 (N_15653,N_15108,N_15005);
or U15654 (N_15654,N_15470,N_15349);
nor U15655 (N_15655,N_15279,N_15023);
nand U15656 (N_15656,N_15251,N_15366);
and U15657 (N_15657,N_15083,N_15437);
or U15658 (N_15658,N_15114,N_15373);
nand U15659 (N_15659,N_15040,N_15372);
or U15660 (N_15660,N_15491,N_15242);
and U15661 (N_15661,N_15134,N_15291);
xor U15662 (N_15662,N_15151,N_15248);
nand U15663 (N_15663,N_15025,N_15070);
xnor U15664 (N_15664,N_15428,N_15457);
nand U15665 (N_15665,N_15392,N_15016);
nor U15666 (N_15666,N_15261,N_15198);
and U15667 (N_15667,N_15381,N_15473);
xor U15668 (N_15668,N_15465,N_15282);
xor U15669 (N_15669,N_15256,N_15343);
or U15670 (N_15670,N_15445,N_15139);
nor U15671 (N_15671,N_15342,N_15053);
and U15672 (N_15672,N_15056,N_15152);
nor U15673 (N_15673,N_15191,N_15124);
nor U15674 (N_15674,N_15000,N_15216);
nor U15675 (N_15675,N_15127,N_15419);
xor U15676 (N_15676,N_15346,N_15327);
or U15677 (N_15677,N_15006,N_15288);
or U15678 (N_15678,N_15087,N_15063);
xor U15679 (N_15679,N_15486,N_15474);
nor U15680 (N_15680,N_15270,N_15100);
xor U15681 (N_15681,N_15208,N_15031);
nand U15682 (N_15682,N_15498,N_15357);
and U15683 (N_15683,N_15324,N_15458);
or U15684 (N_15684,N_15264,N_15464);
nor U15685 (N_15685,N_15410,N_15495);
nor U15686 (N_15686,N_15447,N_15223);
nand U15687 (N_15687,N_15232,N_15330);
and U15688 (N_15688,N_15142,N_15192);
nor U15689 (N_15689,N_15089,N_15178);
and U15690 (N_15690,N_15481,N_15111);
xor U15691 (N_15691,N_15436,N_15203);
nor U15692 (N_15692,N_15035,N_15333);
nand U15693 (N_15693,N_15030,N_15284);
or U15694 (N_15694,N_15378,N_15444);
xnor U15695 (N_15695,N_15224,N_15182);
xor U15696 (N_15696,N_15476,N_15243);
or U15697 (N_15697,N_15002,N_15267);
and U15698 (N_15698,N_15132,N_15493);
or U15699 (N_15699,N_15238,N_15071);
xnor U15700 (N_15700,N_15183,N_15344);
or U15701 (N_15701,N_15415,N_15150);
xor U15702 (N_15702,N_15172,N_15065);
xor U15703 (N_15703,N_15332,N_15045);
xnor U15704 (N_15704,N_15129,N_15388);
nand U15705 (N_15705,N_15205,N_15281);
xor U15706 (N_15706,N_15018,N_15097);
nand U15707 (N_15707,N_15190,N_15060);
or U15708 (N_15708,N_15394,N_15141);
nand U15709 (N_15709,N_15407,N_15379);
and U15710 (N_15710,N_15438,N_15425);
nor U15711 (N_15711,N_15102,N_15402);
xnor U15712 (N_15712,N_15432,N_15133);
and U15713 (N_15713,N_15435,N_15269);
and U15714 (N_15714,N_15351,N_15155);
nand U15715 (N_15715,N_15061,N_15157);
or U15716 (N_15716,N_15274,N_15441);
nor U15717 (N_15717,N_15290,N_15411);
xnor U15718 (N_15718,N_15228,N_15014);
and U15719 (N_15719,N_15259,N_15171);
and U15720 (N_15720,N_15028,N_15386);
or U15721 (N_15721,N_15314,N_15020);
or U15722 (N_15722,N_15292,N_15389);
xor U15723 (N_15723,N_15451,N_15218);
nand U15724 (N_15724,N_15153,N_15499);
nor U15725 (N_15725,N_15140,N_15354);
and U15726 (N_15726,N_15086,N_15042);
nand U15727 (N_15727,N_15459,N_15033);
and U15728 (N_15728,N_15293,N_15489);
or U15729 (N_15729,N_15283,N_15036);
nor U15730 (N_15730,N_15032,N_15181);
xnor U15731 (N_15731,N_15193,N_15377);
or U15732 (N_15732,N_15101,N_15096);
nand U15733 (N_15733,N_15303,N_15454);
nand U15734 (N_15734,N_15138,N_15414);
nand U15735 (N_15735,N_15177,N_15450);
or U15736 (N_15736,N_15396,N_15226);
nand U15737 (N_15737,N_15347,N_15352);
xnor U15738 (N_15738,N_15339,N_15494);
and U15739 (N_15739,N_15165,N_15199);
nand U15740 (N_15740,N_15195,N_15095);
and U15741 (N_15741,N_15180,N_15090);
and U15742 (N_15742,N_15337,N_15049);
nor U15743 (N_15743,N_15456,N_15217);
and U15744 (N_15744,N_15200,N_15369);
nand U15745 (N_15745,N_15367,N_15231);
xor U15746 (N_15746,N_15455,N_15393);
nor U15747 (N_15747,N_15390,N_15074);
nor U15748 (N_15748,N_15313,N_15487);
xnor U15749 (N_15749,N_15222,N_15175);
and U15750 (N_15750,N_15079,N_15127);
nand U15751 (N_15751,N_15319,N_15237);
or U15752 (N_15752,N_15471,N_15141);
and U15753 (N_15753,N_15280,N_15236);
xnor U15754 (N_15754,N_15397,N_15408);
or U15755 (N_15755,N_15032,N_15076);
or U15756 (N_15756,N_15426,N_15455);
xnor U15757 (N_15757,N_15312,N_15176);
and U15758 (N_15758,N_15031,N_15234);
or U15759 (N_15759,N_15157,N_15356);
or U15760 (N_15760,N_15388,N_15460);
or U15761 (N_15761,N_15382,N_15324);
xnor U15762 (N_15762,N_15375,N_15380);
or U15763 (N_15763,N_15268,N_15224);
nand U15764 (N_15764,N_15036,N_15375);
xor U15765 (N_15765,N_15482,N_15084);
xor U15766 (N_15766,N_15158,N_15499);
nand U15767 (N_15767,N_15206,N_15120);
xor U15768 (N_15768,N_15034,N_15442);
nor U15769 (N_15769,N_15402,N_15474);
xor U15770 (N_15770,N_15261,N_15212);
and U15771 (N_15771,N_15219,N_15017);
or U15772 (N_15772,N_15329,N_15083);
nor U15773 (N_15773,N_15323,N_15460);
nand U15774 (N_15774,N_15428,N_15375);
nand U15775 (N_15775,N_15039,N_15431);
or U15776 (N_15776,N_15308,N_15137);
or U15777 (N_15777,N_15268,N_15433);
or U15778 (N_15778,N_15186,N_15180);
and U15779 (N_15779,N_15106,N_15182);
nor U15780 (N_15780,N_15208,N_15137);
and U15781 (N_15781,N_15259,N_15141);
xnor U15782 (N_15782,N_15125,N_15016);
nand U15783 (N_15783,N_15249,N_15458);
or U15784 (N_15784,N_15060,N_15003);
or U15785 (N_15785,N_15476,N_15405);
xnor U15786 (N_15786,N_15149,N_15403);
nand U15787 (N_15787,N_15294,N_15353);
nand U15788 (N_15788,N_15230,N_15116);
nor U15789 (N_15789,N_15472,N_15238);
or U15790 (N_15790,N_15291,N_15156);
nand U15791 (N_15791,N_15059,N_15350);
or U15792 (N_15792,N_15271,N_15469);
xor U15793 (N_15793,N_15397,N_15409);
nand U15794 (N_15794,N_15049,N_15355);
xor U15795 (N_15795,N_15419,N_15309);
or U15796 (N_15796,N_15430,N_15093);
nand U15797 (N_15797,N_15473,N_15277);
nand U15798 (N_15798,N_15341,N_15449);
nand U15799 (N_15799,N_15012,N_15106);
nor U15800 (N_15800,N_15255,N_15385);
nor U15801 (N_15801,N_15098,N_15403);
nor U15802 (N_15802,N_15260,N_15418);
nor U15803 (N_15803,N_15208,N_15335);
xnor U15804 (N_15804,N_15026,N_15207);
xor U15805 (N_15805,N_15245,N_15127);
nor U15806 (N_15806,N_15043,N_15489);
nand U15807 (N_15807,N_15044,N_15385);
and U15808 (N_15808,N_15387,N_15467);
or U15809 (N_15809,N_15228,N_15439);
and U15810 (N_15810,N_15417,N_15385);
xnor U15811 (N_15811,N_15097,N_15440);
nand U15812 (N_15812,N_15135,N_15099);
or U15813 (N_15813,N_15173,N_15056);
and U15814 (N_15814,N_15355,N_15432);
and U15815 (N_15815,N_15185,N_15002);
xor U15816 (N_15816,N_15311,N_15410);
and U15817 (N_15817,N_15088,N_15300);
nor U15818 (N_15818,N_15382,N_15313);
nor U15819 (N_15819,N_15498,N_15135);
nor U15820 (N_15820,N_15397,N_15396);
nand U15821 (N_15821,N_15225,N_15134);
nor U15822 (N_15822,N_15272,N_15338);
xor U15823 (N_15823,N_15212,N_15404);
nand U15824 (N_15824,N_15092,N_15099);
nand U15825 (N_15825,N_15335,N_15255);
nand U15826 (N_15826,N_15446,N_15072);
nor U15827 (N_15827,N_15182,N_15344);
or U15828 (N_15828,N_15054,N_15177);
or U15829 (N_15829,N_15145,N_15305);
xor U15830 (N_15830,N_15426,N_15361);
nor U15831 (N_15831,N_15496,N_15185);
nand U15832 (N_15832,N_15227,N_15127);
nor U15833 (N_15833,N_15493,N_15270);
or U15834 (N_15834,N_15062,N_15152);
xnor U15835 (N_15835,N_15004,N_15245);
nand U15836 (N_15836,N_15451,N_15021);
xor U15837 (N_15837,N_15158,N_15413);
nand U15838 (N_15838,N_15355,N_15188);
nand U15839 (N_15839,N_15258,N_15264);
nor U15840 (N_15840,N_15212,N_15320);
xor U15841 (N_15841,N_15112,N_15440);
and U15842 (N_15842,N_15381,N_15277);
or U15843 (N_15843,N_15466,N_15161);
nor U15844 (N_15844,N_15097,N_15496);
and U15845 (N_15845,N_15390,N_15356);
nand U15846 (N_15846,N_15404,N_15413);
nand U15847 (N_15847,N_15405,N_15057);
nor U15848 (N_15848,N_15092,N_15231);
xor U15849 (N_15849,N_15398,N_15303);
or U15850 (N_15850,N_15111,N_15470);
nand U15851 (N_15851,N_15117,N_15057);
and U15852 (N_15852,N_15435,N_15482);
and U15853 (N_15853,N_15101,N_15406);
and U15854 (N_15854,N_15096,N_15059);
or U15855 (N_15855,N_15268,N_15435);
or U15856 (N_15856,N_15263,N_15209);
nand U15857 (N_15857,N_15184,N_15499);
xor U15858 (N_15858,N_15237,N_15107);
and U15859 (N_15859,N_15012,N_15082);
or U15860 (N_15860,N_15395,N_15094);
and U15861 (N_15861,N_15497,N_15199);
xnor U15862 (N_15862,N_15331,N_15204);
or U15863 (N_15863,N_15421,N_15095);
nand U15864 (N_15864,N_15258,N_15245);
or U15865 (N_15865,N_15072,N_15299);
xor U15866 (N_15866,N_15440,N_15101);
nor U15867 (N_15867,N_15108,N_15186);
nand U15868 (N_15868,N_15212,N_15005);
and U15869 (N_15869,N_15391,N_15352);
nor U15870 (N_15870,N_15433,N_15204);
or U15871 (N_15871,N_15206,N_15412);
xor U15872 (N_15872,N_15322,N_15124);
nand U15873 (N_15873,N_15393,N_15368);
and U15874 (N_15874,N_15261,N_15184);
and U15875 (N_15875,N_15191,N_15387);
nand U15876 (N_15876,N_15425,N_15003);
or U15877 (N_15877,N_15100,N_15150);
nand U15878 (N_15878,N_15269,N_15303);
nand U15879 (N_15879,N_15313,N_15064);
nor U15880 (N_15880,N_15242,N_15286);
nand U15881 (N_15881,N_15159,N_15242);
nor U15882 (N_15882,N_15145,N_15020);
nand U15883 (N_15883,N_15280,N_15122);
and U15884 (N_15884,N_15486,N_15203);
or U15885 (N_15885,N_15390,N_15472);
or U15886 (N_15886,N_15279,N_15312);
or U15887 (N_15887,N_15391,N_15082);
or U15888 (N_15888,N_15198,N_15295);
and U15889 (N_15889,N_15235,N_15492);
or U15890 (N_15890,N_15415,N_15120);
and U15891 (N_15891,N_15191,N_15395);
xor U15892 (N_15892,N_15442,N_15361);
nor U15893 (N_15893,N_15375,N_15424);
xnor U15894 (N_15894,N_15410,N_15069);
nand U15895 (N_15895,N_15113,N_15291);
nand U15896 (N_15896,N_15037,N_15410);
xor U15897 (N_15897,N_15155,N_15083);
or U15898 (N_15898,N_15461,N_15054);
and U15899 (N_15899,N_15314,N_15228);
xnor U15900 (N_15900,N_15042,N_15274);
and U15901 (N_15901,N_15108,N_15144);
xnor U15902 (N_15902,N_15455,N_15103);
nor U15903 (N_15903,N_15236,N_15400);
or U15904 (N_15904,N_15467,N_15078);
or U15905 (N_15905,N_15400,N_15383);
and U15906 (N_15906,N_15289,N_15135);
and U15907 (N_15907,N_15232,N_15299);
or U15908 (N_15908,N_15189,N_15367);
or U15909 (N_15909,N_15133,N_15090);
and U15910 (N_15910,N_15033,N_15397);
xor U15911 (N_15911,N_15189,N_15232);
or U15912 (N_15912,N_15334,N_15142);
nand U15913 (N_15913,N_15092,N_15121);
and U15914 (N_15914,N_15435,N_15490);
nor U15915 (N_15915,N_15224,N_15063);
nand U15916 (N_15916,N_15107,N_15394);
or U15917 (N_15917,N_15327,N_15168);
and U15918 (N_15918,N_15460,N_15442);
or U15919 (N_15919,N_15005,N_15262);
xnor U15920 (N_15920,N_15165,N_15262);
nor U15921 (N_15921,N_15498,N_15296);
and U15922 (N_15922,N_15486,N_15025);
nor U15923 (N_15923,N_15118,N_15291);
and U15924 (N_15924,N_15091,N_15482);
and U15925 (N_15925,N_15350,N_15020);
and U15926 (N_15926,N_15056,N_15361);
xor U15927 (N_15927,N_15129,N_15100);
and U15928 (N_15928,N_15316,N_15231);
and U15929 (N_15929,N_15417,N_15022);
xnor U15930 (N_15930,N_15171,N_15028);
xor U15931 (N_15931,N_15313,N_15267);
and U15932 (N_15932,N_15146,N_15296);
xor U15933 (N_15933,N_15020,N_15262);
or U15934 (N_15934,N_15090,N_15336);
nor U15935 (N_15935,N_15121,N_15417);
xnor U15936 (N_15936,N_15403,N_15143);
xnor U15937 (N_15937,N_15259,N_15257);
nor U15938 (N_15938,N_15106,N_15456);
nand U15939 (N_15939,N_15163,N_15323);
or U15940 (N_15940,N_15489,N_15092);
xor U15941 (N_15941,N_15140,N_15168);
or U15942 (N_15942,N_15038,N_15098);
nand U15943 (N_15943,N_15373,N_15289);
or U15944 (N_15944,N_15080,N_15465);
xnor U15945 (N_15945,N_15357,N_15096);
or U15946 (N_15946,N_15174,N_15140);
or U15947 (N_15947,N_15437,N_15499);
nand U15948 (N_15948,N_15175,N_15152);
and U15949 (N_15949,N_15353,N_15286);
or U15950 (N_15950,N_15089,N_15313);
nor U15951 (N_15951,N_15004,N_15156);
and U15952 (N_15952,N_15049,N_15250);
nand U15953 (N_15953,N_15458,N_15462);
nor U15954 (N_15954,N_15389,N_15010);
and U15955 (N_15955,N_15058,N_15204);
nand U15956 (N_15956,N_15212,N_15083);
nor U15957 (N_15957,N_15012,N_15345);
nand U15958 (N_15958,N_15413,N_15487);
xor U15959 (N_15959,N_15381,N_15221);
and U15960 (N_15960,N_15245,N_15248);
nor U15961 (N_15961,N_15022,N_15178);
or U15962 (N_15962,N_15446,N_15346);
xnor U15963 (N_15963,N_15163,N_15042);
or U15964 (N_15964,N_15059,N_15008);
xor U15965 (N_15965,N_15295,N_15233);
or U15966 (N_15966,N_15193,N_15466);
nand U15967 (N_15967,N_15167,N_15370);
or U15968 (N_15968,N_15479,N_15365);
xnor U15969 (N_15969,N_15391,N_15196);
nor U15970 (N_15970,N_15274,N_15452);
nand U15971 (N_15971,N_15135,N_15440);
xor U15972 (N_15972,N_15336,N_15381);
and U15973 (N_15973,N_15341,N_15115);
nor U15974 (N_15974,N_15121,N_15390);
and U15975 (N_15975,N_15306,N_15191);
nor U15976 (N_15976,N_15311,N_15213);
xor U15977 (N_15977,N_15432,N_15059);
or U15978 (N_15978,N_15320,N_15099);
nand U15979 (N_15979,N_15081,N_15271);
xor U15980 (N_15980,N_15149,N_15439);
or U15981 (N_15981,N_15427,N_15065);
or U15982 (N_15982,N_15386,N_15319);
nand U15983 (N_15983,N_15186,N_15010);
xor U15984 (N_15984,N_15086,N_15327);
nand U15985 (N_15985,N_15283,N_15160);
xor U15986 (N_15986,N_15444,N_15345);
or U15987 (N_15987,N_15362,N_15152);
and U15988 (N_15988,N_15011,N_15033);
nor U15989 (N_15989,N_15494,N_15087);
and U15990 (N_15990,N_15271,N_15432);
nand U15991 (N_15991,N_15352,N_15133);
or U15992 (N_15992,N_15282,N_15218);
and U15993 (N_15993,N_15354,N_15416);
or U15994 (N_15994,N_15340,N_15068);
or U15995 (N_15995,N_15369,N_15119);
and U15996 (N_15996,N_15104,N_15186);
xor U15997 (N_15997,N_15097,N_15201);
xor U15998 (N_15998,N_15022,N_15066);
nand U15999 (N_15999,N_15030,N_15407);
and U16000 (N_16000,N_15804,N_15813);
or U16001 (N_16001,N_15961,N_15985);
nor U16002 (N_16002,N_15958,N_15762);
nor U16003 (N_16003,N_15755,N_15527);
nor U16004 (N_16004,N_15725,N_15971);
xor U16005 (N_16005,N_15710,N_15796);
or U16006 (N_16006,N_15614,N_15878);
xor U16007 (N_16007,N_15953,N_15950);
nand U16008 (N_16008,N_15895,N_15835);
nand U16009 (N_16009,N_15972,N_15545);
or U16010 (N_16010,N_15609,N_15967);
nand U16011 (N_16011,N_15921,N_15868);
nor U16012 (N_16012,N_15862,N_15896);
nand U16013 (N_16013,N_15687,N_15949);
and U16014 (N_16014,N_15936,N_15881);
xor U16015 (N_16015,N_15800,N_15860);
nand U16016 (N_16016,N_15552,N_15660);
xor U16017 (N_16017,N_15995,N_15621);
nand U16018 (N_16018,N_15884,N_15988);
or U16019 (N_16019,N_15951,N_15651);
nor U16020 (N_16020,N_15797,N_15992);
nor U16021 (N_16021,N_15587,N_15541);
or U16022 (N_16022,N_15544,N_15724);
xor U16023 (N_16023,N_15897,N_15954);
nor U16024 (N_16024,N_15568,N_15761);
xor U16025 (N_16025,N_15662,N_15583);
or U16026 (N_16026,N_15556,N_15639);
or U16027 (N_16027,N_15723,N_15682);
nor U16028 (N_16028,N_15877,N_15716);
nor U16029 (N_16029,N_15848,N_15839);
xor U16030 (N_16030,N_15941,N_15880);
nand U16031 (N_16031,N_15719,N_15928);
nand U16032 (N_16032,N_15751,N_15650);
and U16033 (N_16033,N_15667,N_15994);
nor U16034 (N_16034,N_15749,N_15989);
or U16035 (N_16035,N_15592,N_15817);
xor U16036 (N_16036,N_15643,N_15826);
xnor U16037 (N_16037,N_15520,N_15542);
or U16038 (N_16038,N_15634,N_15876);
nor U16039 (N_16039,N_15979,N_15511);
xor U16040 (N_16040,N_15501,N_15683);
or U16041 (N_16041,N_15686,N_15938);
xnor U16042 (N_16042,N_15624,N_15810);
and U16043 (N_16043,N_15676,N_15512);
xnor U16044 (N_16044,N_15866,N_15604);
xnor U16045 (N_16045,N_15806,N_15616);
nand U16046 (N_16046,N_15730,N_15608);
xnor U16047 (N_16047,N_15658,N_15769);
nor U16048 (N_16048,N_15756,N_15818);
nand U16049 (N_16049,N_15704,N_15932);
or U16050 (N_16050,N_15517,N_15875);
or U16051 (N_16051,N_15709,N_15939);
and U16052 (N_16052,N_15691,N_15648);
or U16053 (N_16053,N_15955,N_15846);
and U16054 (N_16054,N_15534,N_15693);
xnor U16055 (N_16055,N_15638,N_15622);
xnor U16056 (N_16056,N_15526,N_15873);
and U16057 (N_16057,N_15681,N_15504);
or U16058 (N_16058,N_15990,N_15991);
xor U16059 (N_16059,N_15692,N_15564);
nand U16060 (N_16060,N_15523,N_15849);
nor U16061 (N_16061,N_15959,N_15633);
nand U16062 (N_16062,N_15580,N_15904);
xor U16063 (N_16063,N_15976,N_15906);
nand U16064 (N_16064,N_15503,N_15940);
nand U16065 (N_16065,N_15659,N_15822);
and U16066 (N_16066,N_15879,N_15783);
and U16067 (N_16067,N_15828,N_15737);
and U16068 (N_16068,N_15701,N_15854);
and U16069 (N_16069,N_15726,N_15948);
xor U16070 (N_16070,N_15907,N_15857);
xnor U16071 (N_16071,N_15942,N_15698);
xnor U16072 (N_16072,N_15969,N_15790);
and U16073 (N_16073,N_15700,N_15766);
or U16074 (N_16074,N_15827,N_15833);
or U16075 (N_16075,N_15689,N_15760);
nand U16076 (N_16076,N_15842,N_15588);
nand U16077 (N_16077,N_15772,N_15718);
and U16078 (N_16078,N_15536,N_15562);
and U16079 (N_16079,N_15602,N_15944);
and U16080 (N_16080,N_15533,N_15712);
nand U16081 (N_16081,N_15539,N_15661);
xnor U16082 (N_16082,N_15641,N_15620);
nor U16083 (N_16083,N_15898,N_15981);
nor U16084 (N_16084,N_15585,N_15531);
or U16085 (N_16085,N_15763,N_15966);
nand U16086 (N_16086,N_15745,N_15522);
or U16087 (N_16087,N_15919,N_15851);
nand U16088 (N_16088,N_15853,N_15535);
nand U16089 (N_16089,N_15720,N_15986);
nor U16090 (N_16090,N_15657,N_15798);
and U16091 (N_16091,N_15613,N_15632);
xnor U16092 (N_16092,N_15599,N_15572);
xor U16093 (N_16093,N_15934,N_15836);
or U16094 (N_16094,N_15812,N_15560);
xnor U16095 (N_16095,N_15708,N_15765);
nand U16096 (N_16096,N_15780,N_15824);
nor U16097 (N_16097,N_15987,N_15838);
or U16098 (N_16098,N_15914,N_15586);
xnor U16099 (N_16099,N_15680,N_15841);
nor U16100 (N_16100,N_15980,N_15722);
nand U16101 (N_16101,N_15637,N_15665);
xnor U16102 (N_16102,N_15867,N_15802);
or U16103 (N_16103,N_15732,N_15548);
nor U16104 (N_16104,N_15628,N_15711);
xnor U16105 (N_16105,N_15820,N_15815);
nand U16106 (N_16106,N_15601,N_15508);
xor U16107 (N_16107,N_15740,N_15748);
xnor U16108 (N_16108,N_15502,N_15540);
and U16109 (N_16109,N_15837,N_15823);
or U16110 (N_16110,N_15964,N_15874);
and U16111 (N_16111,N_15754,N_15774);
or U16112 (N_16112,N_15612,N_15509);
and U16113 (N_16113,N_15594,N_15695);
or U16114 (N_16114,N_15669,N_15819);
nor U16115 (N_16115,N_15629,N_15734);
xor U16116 (N_16116,N_15529,N_15753);
and U16117 (N_16117,N_15935,N_15524);
or U16118 (N_16118,N_15767,N_15702);
or U16119 (N_16119,N_15727,N_15674);
nor U16120 (N_16120,N_15558,N_15644);
xor U16121 (N_16121,N_15821,N_15902);
and U16122 (N_16122,N_15965,N_15844);
or U16123 (N_16123,N_15924,N_15909);
nand U16124 (N_16124,N_15832,N_15752);
xnor U16125 (N_16125,N_15619,N_15561);
or U16126 (N_16126,N_15591,N_15889);
xor U16127 (N_16127,N_15926,N_15997);
nor U16128 (N_16128,N_15703,N_15506);
and U16129 (N_16129,N_15892,N_15672);
nand U16130 (N_16130,N_15746,N_15597);
nand U16131 (N_16131,N_15855,N_15673);
xnor U16132 (N_16132,N_15912,N_15782);
nand U16133 (N_16133,N_15625,N_15685);
nand U16134 (N_16134,N_15890,N_15525);
or U16135 (N_16135,N_15847,N_15910);
xnor U16136 (N_16136,N_15963,N_15956);
and U16137 (N_16137,N_15915,N_15929);
nand U16138 (N_16138,N_15707,N_15553);
xor U16139 (N_16139,N_15596,N_15789);
nor U16140 (N_16140,N_15678,N_15688);
xnor U16141 (N_16141,N_15858,N_15576);
nor U16142 (N_16142,N_15668,N_15977);
nand U16143 (N_16143,N_15581,N_15792);
and U16144 (N_16144,N_15786,N_15829);
nor U16145 (N_16145,N_15869,N_15664);
and U16146 (N_16146,N_15984,N_15584);
nor U16147 (N_16147,N_15758,N_15610);
nand U16148 (N_16148,N_15776,N_15831);
xnor U16149 (N_16149,N_15735,N_15946);
and U16150 (N_16150,N_15656,N_15647);
or U16151 (N_16151,N_15917,N_15952);
nand U16152 (N_16152,N_15960,N_15805);
and U16153 (N_16153,N_15787,N_15808);
xnor U16154 (N_16154,N_15652,N_15739);
nand U16155 (N_16155,N_15903,N_15670);
nor U16156 (N_16156,N_15861,N_15883);
nand U16157 (N_16157,N_15887,N_15554);
xnor U16158 (N_16158,N_15923,N_15882);
and U16159 (N_16159,N_15742,N_15566);
and U16160 (N_16160,N_15801,N_15825);
or U16161 (N_16161,N_15916,N_15738);
or U16162 (N_16162,N_15514,N_15671);
xor U16163 (N_16163,N_15532,N_15507);
or U16164 (N_16164,N_15615,N_15705);
xor U16165 (N_16165,N_15519,N_15918);
xnor U16166 (N_16166,N_15713,N_15894);
nand U16167 (N_16167,N_15649,N_15537);
xnor U16168 (N_16168,N_15970,N_15595);
and U16169 (N_16169,N_15996,N_15764);
nor U16170 (N_16170,N_15856,N_15654);
nand U16171 (N_16171,N_15925,N_15603);
xnor U16172 (N_16172,N_15922,N_15741);
or U16173 (N_16173,N_15975,N_15973);
nand U16174 (N_16174,N_15546,N_15515);
and U16175 (N_16175,N_15559,N_15843);
or U16176 (N_16176,N_15888,N_15781);
nand U16177 (N_16177,N_15850,N_15530);
or U16178 (N_16178,N_15978,N_15598);
and U16179 (N_16179,N_15589,N_15768);
nor U16180 (N_16180,N_15690,N_15500);
nor U16181 (N_16181,N_15807,N_15635);
nor U16182 (N_16182,N_15655,N_15777);
and U16183 (N_16183,N_15794,N_15518);
xnor U16184 (N_16184,N_15911,N_15640);
xnor U16185 (N_16185,N_15575,N_15570);
and U16186 (N_16186,N_15627,N_15791);
and U16187 (N_16187,N_15770,N_15731);
nor U16188 (N_16188,N_15666,N_15646);
nand U16189 (N_16189,N_15947,N_15814);
nand U16190 (N_16190,N_15549,N_15505);
nor U16191 (N_16191,N_15573,N_15779);
nand U16192 (N_16192,N_15771,N_15998);
nand U16193 (N_16193,N_15577,N_15582);
nand U16194 (N_16194,N_15611,N_15852);
nor U16195 (N_16195,N_15927,N_15795);
nor U16196 (N_16196,N_15901,N_15793);
and U16197 (N_16197,N_15571,N_15905);
nand U16198 (N_16198,N_15893,N_15697);
xnor U16199 (N_16199,N_15679,N_15528);
and U16200 (N_16200,N_15677,N_15943);
or U16201 (N_16201,N_15663,N_15579);
or U16202 (N_16202,N_15871,N_15908);
or U16203 (N_16203,N_15930,N_15605);
xnor U16204 (N_16204,N_15645,N_15773);
or U16205 (N_16205,N_15617,N_15945);
nor U16206 (N_16206,N_15993,N_15865);
nor U16207 (N_16207,N_15626,N_15717);
xnor U16208 (N_16208,N_15606,N_15982);
or U16209 (N_16209,N_15569,N_15631);
xnor U16210 (N_16210,N_15600,N_15642);
xnor U16211 (N_16211,N_15636,N_15729);
or U16212 (N_16212,N_15593,N_15983);
xor U16213 (N_16213,N_15968,N_15872);
xnor U16214 (N_16214,N_15788,N_15785);
nor U16215 (N_16215,N_15778,N_15538);
nand U16216 (N_16216,N_15757,N_15607);
and U16217 (N_16217,N_15784,N_15590);
xnor U16218 (N_16218,N_15962,N_15937);
or U16219 (N_16219,N_15543,N_15574);
and U16220 (N_16220,N_15863,N_15900);
and U16221 (N_16221,N_15759,N_15744);
xnor U16222 (N_16222,N_15999,N_15834);
nand U16223 (N_16223,N_15721,N_15675);
and U16224 (N_16224,N_15957,N_15920);
xnor U16225 (N_16225,N_15859,N_15696);
or U16226 (N_16226,N_15885,N_15811);
or U16227 (N_16227,N_15891,N_15551);
or U16228 (N_16228,N_15931,N_15567);
xor U16229 (N_16229,N_15510,N_15513);
or U16230 (N_16230,N_15699,N_15733);
and U16231 (N_16231,N_15618,N_15684);
nand U16232 (N_16232,N_15840,N_15565);
xnor U16233 (N_16233,N_15816,N_15555);
xnor U16234 (N_16234,N_15694,N_15747);
nand U16235 (N_16235,N_15706,N_15728);
xnor U16236 (N_16236,N_15550,N_15870);
or U16237 (N_16237,N_15743,N_15803);
nand U16238 (N_16238,N_15799,N_15714);
xor U16239 (N_16239,N_15736,N_15913);
nand U16240 (N_16240,N_15557,N_15563);
and U16241 (N_16241,N_15630,N_15715);
nand U16242 (N_16242,N_15623,N_15653);
and U16243 (N_16243,N_15809,N_15886);
nand U16244 (N_16244,N_15830,N_15775);
nand U16245 (N_16245,N_15750,N_15845);
nor U16246 (N_16246,N_15864,N_15516);
and U16247 (N_16247,N_15578,N_15899);
and U16248 (N_16248,N_15521,N_15547);
nor U16249 (N_16249,N_15933,N_15974);
and U16250 (N_16250,N_15930,N_15691);
nor U16251 (N_16251,N_15891,N_15757);
nand U16252 (N_16252,N_15790,N_15745);
nor U16253 (N_16253,N_15750,N_15819);
xor U16254 (N_16254,N_15716,N_15543);
nand U16255 (N_16255,N_15640,N_15928);
or U16256 (N_16256,N_15734,N_15676);
nor U16257 (N_16257,N_15666,N_15761);
xor U16258 (N_16258,N_15725,N_15530);
nand U16259 (N_16259,N_15960,N_15938);
or U16260 (N_16260,N_15660,N_15935);
or U16261 (N_16261,N_15610,N_15845);
and U16262 (N_16262,N_15623,N_15535);
nand U16263 (N_16263,N_15852,N_15579);
nand U16264 (N_16264,N_15789,N_15995);
or U16265 (N_16265,N_15749,N_15832);
nor U16266 (N_16266,N_15755,N_15607);
xnor U16267 (N_16267,N_15708,N_15633);
nor U16268 (N_16268,N_15950,N_15931);
nor U16269 (N_16269,N_15902,N_15934);
nor U16270 (N_16270,N_15763,N_15952);
nor U16271 (N_16271,N_15935,N_15837);
xnor U16272 (N_16272,N_15907,N_15786);
or U16273 (N_16273,N_15681,N_15945);
nor U16274 (N_16274,N_15592,N_15713);
nor U16275 (N_16275,N_15864,N_15847);
and U16276 (N_16276,N_15694,N_15966);
nand U16277 (N_16277,N_15609,N_15682);
nor U16278 (N_16278,N_15670,N_15711);
or U16279 (N_16279,N_15879,N_15652);
nor U16280 (N_16280,N_15891,N_15594);
or U16281 (N_16281,N_15703,N_15842);
and U16282 (N_16282,N_15510,N_15816);
nand U16283 (N_16283,N_15923,N_15601);
and U16284 (N_16284,N_15548,N_15872);
nand U16285 (N_16285,N_15707,N_15979);
nand U16286 (N_16286,N_15642,N_15707);
nand U16287 (N_16287,N_15525,N_15965);
nand U16288 (N_16288,N_15781,N_15672);
nor U16289 (N_16289,N_15876,N_15820);
nand U16290 (N_16290,N_15747,N_15922);
nand U16291 (N_16291,N_15821,N_15929);
or U16292 (N_16292,N_15575,N_15746);
nand U16293 (N_16293,N_15788,N_15868);
nor U16294 (N_16294,N_15810,N_15546);
or U16295 (N_16295,N_15712,N_15823);
nand U16296 (N_16296,N_15657,N_15661);
or U16297 (N_16297,N_15807,N_15525);
nand U16298 (N_16298,N_15906,N_15839);
or U16299 (N_16299,N_15729,N_15638);
or U16300 (N_16300,N_15782,N_15751);
xor U16301 (N_16301,N_15720,N_15894);
and U16302 (N_16302,N_15628,N_15724);
or U16303 (N_16303,N_15825,N_15979);
xor U16304 (N_16304,N_15770,N_15805);
nand U16305 (N_16305,N_15921,N_15824);
nand U16306 (N_16306,N_15525,N_15612);
nand U16307 (N_16307,N_15893,N_15904);
or U16308 (N_16308,N_15614,N_15771);
xnor U16309 (N_16309,N_15565,N_15791);
xor U16310 (N_16310,N_15631,N_15614);
or U16311 (N_16311,N_15631,N_15573);
and U16312 (N_16312,N_15655,N_15651);
xor U16313 (N_16313,N_15859,N_15600);
xnor U16314 (N_16314,N_15823,N_15820);
nand U16315 (N_16315,N_15829,N_15750);
nand U16316 (N_16316,N_15782,N_15722);
and U16317 (N_16317,N_15678,N_15823);
xor U16318 (N_16318,N_15874,N_15888);
xor U16319 (N_16319,N_15813,N_15690);
or U16320 (N_16320,N_15777,N_15897);
and U16321 (N_16321,N_15642,N_15911);
nor U16322 (N_16322,N_15758,N_15712);
xnor U16323 (N_16323,N_15786,N_15818);
nand U16324 (N_16324,N_15715,N_15743);
and U16325 (N_16325,N_15787,N_15886);
nand U16326 (N_16326,N_15905,N_15609);
xnor U16327 (N_16327,N_15948,N_15887);
nand U16328 (N_16328,N_15769,N_15818);
or U16329 (N_16329,N_15781,N_15843);
nand U16330 (N_16330,N_15575,N_15948);
xor U16331 (N_16331,N_15723,N_15666);
xor U16332 (N_16332,N_15981,N_15765);
xnor U16333 (N_16333,N_15604,N_15560);
nand U16334 (N_16334,N_15531,N_15882);
or U16335 (N_16335,N_15692,N_15555);
and U16336 (N_16336,N_15703,N_15713);
xor U16337 (N_16337,N_15778,N_15880);
and U16338 (N_16338,N_15515,N_15796);
or U16339 (N_16339,N_15690,N_15674);
xnor U16340 (N_16340,N_15946,N_15525);
xor U16341 (N_16341,N_15595,N_15659);
nor U16342 (N_16342,N_15679,N_15964);
xor U16343 (N_16343,N_15716,N_15558);
nand U16344 (N_16344,N_15896,N_15563);
or U16345 (N_16345,N_15779,N_15569);
nor U16346 (N_16346,N_15781,N_15762);
nand U16347 (N_16347,N_15958,N_15934);
and U16348 (N_16348,N_15706,N_15972);
or U16349 (N_16349,N_15515,N_15870);
nor U16350 (N_16350,N_15677,N_15734);
nand U16351 (N_16351,N_15506,N_15508);
nor U16352 (N_16352,N_15933,N_15991);
nand U16353 (N_16353,N_15732,N_15906);
nand U16354 (N_16354,N_15628,N_15697);
nand U16355 (N_16355,N_15961,N_15799);
and U16356 (N_16356,N_15626,N_15709);
nand U16357 (N_16357,N_15575,N_15815);
xor U16358 (N_16358,N_15953,N_15879);
nand U16359 (N_16359,N_15892,N_15947);
nand U16360 (N_16360,N_15869,N_15566);
and U16361 (N_16361,N_15738,N_15615);
nand U16362 (N_16362,N_15993,N_15987);
nand U16363 (N_16363,N_15666,N_15997);
nor U16364 (N_16364,N_15722,N_15766);
and U16365 (N_16365,N_15840,N_15516);
or U16366 (N_16366,N_15988,N_15501);
or U16367 (N_16367,N_15761,N_15659);
or U16368 (N_16368,N_15650,N_15864);
nor U16369 (N_16369,N_15857,N_15776);
or U16370 (N_16370,N_15565,N_15843);
and U16371 (N_16371,N_15504,N_15755);
xor U16372 (N_16372,N_15656,N_15953);
xor U16373 (N_16373,N_15751,N_15841);
xor U16374 (N_16374,N_15682,N_15511);
or U16375 (N_16375,N_15922,N_15972);
nor U16376 (N_16376,N_15824,N_15947);
xnor U16377 (N_16377,N_15920,N_15611);
and U16378 (N_16378,N_15976,N_15740);
xor U16379 (N_16379,N_15953,N_15520);
nor U16380 (N_16380,N_15523,N_15897);
or U16381 (N_16381,N_15997,N_15593);
nor U16382 (N_16382,N_15713,N_15880);
xnor U16383 (N_16383,N_15608,N_15767);
or U16384 (N_16384,N_15625,N_15715);
nand U16385 (N_16385,N_15617,N_15507);
xnor U16386 (N_16386,N_15910,N_15647);
xor U16387 (N_16387,N_15636,N_15603);
xor U16388 (N_16388,N_15668,N_15580);
or U16389 (N_16389,N_15651,N_15607);
nor U16390 (N_16390,N_15765,N_15930);
or U16391 (N_16391,N_15784,N_15828);
xnor U16392 (N_16392,N_15674,N_15656);
nand U16393 (N_16393,N_15549,N_15646);
or U16394 (N_16394,N_15985,N_15722);
and U16395 (N_16395,N_15562,N_15509);
or U16396 (N_16396,N_15897,N_15822);
xnor U16397 (N_16397,N_15792,N_15880);
and U16398 (N_16398,N_15655,N_15682);
and U16399 (N_16399,N_15787,N_15753);
or U16400 (N_16400,N_15982,N_15742);
nor U16401 (N_16401,N_15921,N_15567);
and U16402 (N_16402,N_15666,N_15715);
or U16403 (N_16403,N_15665,N_15654);
nor U16404 (N_16404,N_15926,N_15815);
nor U16405 (N_16405,N_15922,N_15772);
nand U16406 (N_16406,N_15966,N_15698);
nand U16407 (N_16407,N_15731,N_15844);
and U16408 (N_16408,N_15717,N_15634);
and U16409 (N_16409,N_15758,N_15754);
and U16410 (N_16410,N_15520,N_15573);
nand U16411 (N_16411,N_15709,N_15677);
or U16412 (N_16412,N_15626,N_15584);
and U16413 (N_16413,N_15924,N_15511);
nand U16414 (N_16414,N_15561,N_15952);
nor U16415 (N_16415,N_15891,N_15880);
nor U16416 (N_16416,N_15680,N_15888);
or U16417 (N_16417,N_15544,N_15675);
nor U16418 (N_16418,N_15900,N_15690);
nor U16419 (N_16419,N_15994,N_15553);
nand U16420 (N_16420,N_15980,N_15671);
and U16421 (N_16421,N_15729,N_15899);
or U16422 (N_16422,N_15546,N_15746);
nor U16423 (N_16423,N_15662,N_15988);
xor U16424 (N_16424,N_15858,N_15723);
and U16425 (N_16425,N_15811,N_15924);
and U16426 (N_16426,N_15584,N_15756);
or U16427 (N_16427,N_15508,N_15615);
or U16428 (N_16428,N_15988,N_15847);
or U16429 (N_16429,N_15626,N_15528);
or U16430 (N_16430,N_15937,N_15765);
xnor U16431 (N_16431,N_15944,N_15807);
xor U16432 (N_16432,N_15938,N_15874);
xnor U16433 (N_16433,N_15917,N_15691);
nor U16434 (N_16434,N_15808,N_15985);
nor U16435 (N_16435,N_15556,N_15570);
and U16436 (N_16436,N_15582,N_15664);
and U16437 (N_16437,N_15957,N_15869);
or U16438 (N_16438,N_15512,N_15802);
and U16439 (N_16439,N_15858,N_15931);
nand U16440 (N_16440,N_15595,N_15837);
xor U16441 (N_16441,N_15606,N_15519);
and U16442 (N_16442,N_15579,N_15666);
nor U16443 (N_16443,N_15579,N_15948);
and U16444 (N_16444,N_15770,N_15906);
nand U16445 (N_16445,N_15800,N_15963);
xor U16446 (N_16446,N_15616,N_15725);
and U16447 (N_16447,N_15712,N_15971);
nand U16448 (N_16448,N_15533,N_15902);
xnor U16449 (N_16449,N_15935,N_15758);
nor U16450 (N_16450,N_15619,N_15535);
xnor U16451 (N_16451,N_15546,N_15518);
nor U16452 (N_16452,N_15726,N_15694);
nor U16453 (N_16453,N_15778,N_15810);
xnor U16454 (N_16454,N_15752,N_15978);
xor U16455 (N_16455,N_15736,N_15737);
and U16456 (N_16456,N_15805,N_15992);
xor U16457 (N_16457,N_15950,N_15515);
or U16458 (N_16458,N_15513,N_15929);
nand U16459 (N_16459,N_15612,N_15575);
or U16460 (N_16460,N_15526,N_15715);
nor U16461 (N_16461,N_15946,N_15762);
nor U16462 (N_16462,N_15623,N_15532);
or U16463 (N_16463,N_15599,N_15632);
and U16464 (N_16464,N_15911,N_15517);
or U16465 (N_16465,N_15586,N_15969);
and U16466 (N_16466,N_15563,N_15955);
nor U16467 (N_16467,N_15704,N_15761);
or U16468 (N_16468,N_15822,N_15718);
nor U16469 (N_16469,N_15631,N_15557);
nor U16470 (N_16470,N_15922,N_15994);
xnor U16471 (N_16471,N_15950,N_15639);
nor U16472 (N_16472,N_15770,N_15723);
nand U16473 (N_16473,N_15786,N_15777);
and U16474 (N_16474,N_15823,N_15657);
or U16475 (N_16475,N_15849,N_15625);
nand U16476 (N_16476,N_15562,N_15736);
and U16477 (N_16477,N_15932,N_15652);
and U16478 (N_16478,N_15634,N_15939);
nand U16479 (N_16479,N_15898,N_15712);
xnor U16480 (N_16480,N_15787,N_15696);
nand U16481 (N_16481,N_15776,N_15766);
or U16482 (N_16482,N_15688,N_15605);
nor U16483 (N_16483,N_15931,N_15619);
nand U16484 (N_16484,N_15854,N_15623);
xor U16485 (N_16485,N_15662,N_15612);
and U16486 (N_16486,N_15922,N_15528);
xor U16487 (N_16487,N_15751,N_15851);
or U16488 (N_16488,N_15502,N_15762);
nor U16489 (N_16489,N_15901,N_15584);
xnor U16490 (N_16490,N_15583,N_15585);
or U16491 (N_16491,N_15607,N_15962);
xnor U16492 (N_16492,N_15974,N_15804);
nor U16493 (N_16493,N_15794,N_15618);
and U16494 (N_16494,N_15910,N_15885);
or U16495 (N_16495,N_15610,N_15823);
or U16496 (N_16496,N_15959,N_15833);
xnor U16497 (N_16497,N_15868,N_15630);
and U16498 (N_16498,N_15746,N_15695);
xnor U16499 (N_16499,N_15757,N_15513);
and U16500 (N_16500,N_16030,N_16202);
nor U16501 (N_16501,N_16133,N_16099);
or U16502 (N_16502,N_16003,N_16112);
and U16503 (N_16503,N_16461,N_16225);
or U16504 (N_16504,N_16093,N_16022);
and U16505 (N_16505,N_16032,N_16113);
or U16506 (N_16506,N_16242,N_16345);
or U16507 (N_16507,N_16415,N_16498);
and U16508 (N_16508,N_16340,N_16495);
xnor U16509 (N_16509,N_16066,N_16426);
and U16510 (N_16510,N_16147,N_16352);
or U16511 (N_16511,N_16275,N_16063);
and U16512 (N_16512,N_16119,N_16135);
nor U16513 (N_16513,N_16049,N_16251);
nand U16514 (N_16514,N_16467,N_16444);
xor U16515 (N_16515,N_16273,N_16075);
or U16516 (N_16516,N_16156,N_16189);
or U16517 (N_16517,N_16392,N_16236);
nand U16518 (N_16518,N_16141,N_16097);
xnor U16519 (N_16519,N_16404,N_16262);
and U16520 (N_16520,N_16304,N_16215);
or U16521 (N_16521,N_16442,N_16435);
and U16522 (N_16522,N_16471,N_16419);
and U16523 (N_16523,N_16186,N_16449);
xor U16524 (N_16524,N_16343,N_16443);
nor U16525 (N_16525,N_16402,N_16493);
nor U16526 (N_16526,N_16428,N_16098);
and U16527 (N_16527,N_16420,N_16111);
nor U16528 (N_16528,N_16146,N_16137);
nor U16529 (N_16529,N_16168,N_16394);
and U16530 (N_16530,N_16438,N_16458);
or U16531 (N_16531,N_16332,N_16474);
and U16532 (N_16532,N_16244,N_16488);
or U16533 (N_16533,N_16058,N_16121);
nor U16534 (N_16534,N_16054,N_16026);
nand U16535 (N_16535,N_16334,N_16257);
or U16536 (N_16536,N_16092,N_16487);
nor U16537 (N_16537,N_16480,N_16131);
and U16538 (N_16538,N_16071,N_16292);
or U16539 (N_16539,N_16170,N_16452);
or U16540 (N_16540,N_16078,N_16395);
nand U16541 (N_16541,N_16329,N_16101);
and U16542 (N_16542,N_16199,N_16248);
xor U16543 (N_16543,N_16268,N_16254);
nor U16544 (N_16544,N_16413,N_16446);
and U16545 (N_16545,N_16211,N_16416);
xnor U16546 (N_16546,N_16074,N_16051);
nand U16547 (N_16547,N_16057,N_16210);
nand U16548 (N_16548,N_16103,N_16110);
or U16549 (N_16549,N_16319,N_16400);
or U16550 (N_16550,N_16497,N_16323);
or U16551 (N_16551,N_16441,N_16204);
nor U16552 (N_16552,N_16486,N_16020);
nor U16553 (N_16553,N_16264,N_16348);
xor U16554 (N_16554,N_16263,N_16157);
nand U16555 (N_16555,N_16360,N_16270);
xnor U16556 (N_16556,N_16277,N_16298);
nor U16557 (N_16557,N_16029,N_16371);
nor U16558 (N_16558,N_16172,N_16318);
nand U16559 (N_16559,N_16109,N_16280);
and U16560 (N_16560,N_16291,N_16485);
and U16561 (N_16561,N_16370,N_16136);
and U16562 (N_16562,N_16321,N_16408);
xor U16563 (N_16563,N_16207,N_16489);
xor U16564 (N_16564,N_16269,N_16007);
nor U16565 (N_16565,N_16324,N_16350);
xor U16566 (N_16566,N_16469,N_16399);
nor U16567 (N_16567,N_16261,N_16125);
or U16568 (N_16568,N_16123,N_16366);
xnor U16569 (N_16569,N_16358,N_16148);
nand U16570 (N_16570,N_16256,N_16312);
and U16571 (N_16571,N_16173,N_16266);
nor U16572 (N_16572,N_16140,N_16061);
xnor U16573 (N_16573,N_16044,N_16373);
xnor U16574 (N_16574,N_16245,N_16363);
or U16575 (N_16575,N_16466,N_16430);
xnor U16576 (N_16576,N_16201,N_16023);
or U16577 (N_16577,N_16187,N_16293);
or U16578 (N_16578,N_16359,N_16166);
and U16579 (N_16579,N_16265,N_16152);
nand U16580 (N_16580,N_16445,N_16299);
nand U16581 (N_16581,N_16039,N_16380);
nor U16582 (N_16582,N_16305,N_16214);
or U16583 (N_16583,N_16138,N_16302);
nand U16584 (N_16584,N_16209,N_16388);
nor U16585 (N_16585,N_16116,N_16376);
xor U16586 (N_16586,N_16234,N_16038);
nand U16587 (N_16587,N_16255,N_16353);
and U16588 (N_16588,N_16468,N_16374);
nor U16589 (N_16589,N_16190,N_16258);
nor U16590 (N_16590,N_16182,N_16027);
or U16591 (N_16591,N_16477,N_16288);
nand U16592 (N_16592,N_16117,N_16375);
or U16593 (N_16593,N_16118,N_16317);
nand U16594 (N_16594,N_16001,N_16224);
nor U16595 (N_16595,N_16046,N_16300);
and U16596 (N_16596,N_16000,N_16424);
and U16597 (N_16597,N_16231,N_16129);
xnor U16598 (N_16598,N_16412,N_16155);
nand U16599 (N_16599,N_16179,N_16378);
nand U16600 (N_16600,N_16176,N_16218);
nor U16601 (N_16601,N_16069,N_16114);
and U16602 (N_16602,N_16494,N_16278);
or U16603 (N_16603,N_16055,N_16087);
and U16604 (N_16604,N_16240,N_16169);
or U16605 (N_16605,N_16397,N_16200);
nor U16606 (N_16606,N_16437,N_16162);
xnor U16607 (N_16607,N_16223,N_16349);
and U16608 (N_16608,N_16188,N_16154);
or U16609 (N_16609,N_16130,N_16230);
nor U16610 (N_16610,N_16473,N_16427);
and U16611 (N_16611,N_16396,N_16060);
and U16612 (N_16612,N_16422,N_16167);
nor U16613 (N_16613,N_16213,N_16227);
nand U16614 (N_16614,N_16237,N_16279);
and U16615 (N_16615,N_16401,N_16433);
and U16616 (N_16616,N_16357,N_16386);
and U16617 (N_16617,N_16481,N_16295);
nand U16618 (N_16618,N_16195,N_16206);
nand U16619 (N_16619,N_16341,N_16301);
or U16620 (N_16620,N_16381,N_16454);
or U16621 (N_16621,N_16105,N_16226);
nor U16622 (N_16622,N_16409,N_16077);
or U16623 (N_16623,N_16490,N_16184);
xor U16624 (N_16624,N_16034,N_16239);
nor U16625 (N_16625,N_16017,N_16120);
nor U16626 (N_16626,N_16456,N_16059);
and U16627 (N_16627,N_16271,N_16342);
xnor U16628 (N_16628,N_16390,N_16475);
nor U16629 (N_16629,N_16483,N_16222);
or U16630 (N_16630,N_16434,N_16042);
xor U16631 (N_16631,N_16096,N_16217);
or U16632 (N_16632,N_16124,N_16286);
nand U16633 (N_16633,N_16250,N_16016);
nor U16634 (N_16634,N_16315,N_16079);
nor U16635 (N_16635,N_16457,N_16432);
or U16636 (N_16636,N_16149,N_16073);
xor U16637 (N_16637,N_16372,N_16090);
nor U16638 (N_16638,N_16327,N_16128);
xnor U16639 (N_16639,N_16142,N_16134);
xor U16640 (N_16640,N_16013,N_16339);
nor U16641 (N_16641,N_16122,N_16229);
xnor U16642 (N_16642,N_16355,N_16008);
or U16643 (N_16643,N_16153,N_16132);
and U16644 (N_16644,N_16283,N_16065);
xor U16645 (N_16645,N_16083,N_16330);
and U16646 (N_16646,N_16084,N_16068);
nand U16647 (N_16647,N_16450,N_16150);
nor U16648 (N_16648,N_16335,N_16285);
xnor U16649 (N_16649,N_16080,N_16064);
nor U16650 (N_16650,N_16043,N_16499);
or U16651 (N_16651,N_16484,N_16476);
and U16652 (N_16652,N_16470,N_16391);
nor U16653 (N_16653,N_16205,N_16050);
nor U16654 (N_16654,N_16235,N_16455);
or U16655 (N_16655,N_16451,N_16462);
nor U16656 (N_16656,N_16056,N_16383);
nor U16657 (N_16657,N_16398,N_16326);
xnor U16658 (N_16658,N_16294,N_16151);
xor U16659 (N_16659,N_16439,N_16070);
nor U16660 (N_16660,N_16431,N_16037);
nor U16661 (N_16661,N_16320,N_16067);
nor U16662 (N_16662,N_16407,N_16482);
nor U16663 (N_16663,N_16004,N_16336);
nand U16664 (N_16664,N_16178,N_16405);
xor U16665 (N_16665,N_16351,N_16423);
xnor U16666 (N_16666,N_16108,N_16448);
nand U16667 (N_16667,N_16344,N_16382);
nor U16668 (N_16668,N_16192,N_16379);
and U16669 (N_16669,N_16024,N_16102);
nor U16670 (N_16670,N_16233,N_16181);
xnor U16671 (N_16671,N_16281,N_16310);
and U16672 (N_16672,N_16272,N_16085);
nand U16673 (N_16673,N_16425,N_16472);
nor U16674 (N_16674,N_16328,N_16316);
and U16675 (N_16675,N_16246,N_16354);
xnor U16676 (N_16676,N_16249,N_16440);
nor U16677 (N_16677,N_16021,N_16377);
or U16678 (N_16678,N_16158,N_16290);
xor U16679 (N_16679,N_16282,N_16459);
nand U16680 (N_16680,N_16018,N_16238);
nor U16681 (N_16681,N_16106,N_16091);
xnor U16682 (N_16682,N_16252,N_16465);
xnor U16683 (N_16683,N_16002,N_16198);
or U16684 (N_16684,N_16010,N_16447);
and U16685 (N_16685,N_16127,N_16019);
nor U16686 (N_16686,N_16347,N_16139);
nand U16687 (N_16687,N_16062,N_16296);
nand U16688 (N_16688,N_16389,N_16314);
nor U16689 (N_16689,N_16191,N_16417);
nand U16690 (N_16690,N_16196,N_16479);
xor U16691 (N_16691,N_16175,N_16356);
xor U16692 (N_16692,N_16194,N_16009);
xor U16693 (N_16693,N_16040,N_16011);
and U16694 (N_16694,N_16276,N_16309);
nor U16695 (N_16695,N_16367,N_16185);
nand U16696 (N_16696,N_16403,N_16333);
nand U16697 (N_16697,N_16308,N_16460);
and U16698 (N_16698,N_16174,N_16267);
and U16699 (N_16699,N_16163,N_16406);
and U16700 (N_16700,N_16159,N_16035);
xor U16701 (N_16701,N_16274,N_16247);
nor U16702 (N_16702,N_16107,N_16387);
nand U16703 (N_16703,N_16165,N_16453);
nor U16704 (N_16704,N_16411,N_16052);
and U16705 (N_16705,N_16464,N_16418);
or U16706 (N_16706,N_16492,N_16033);
nand U16707 (N_16707,N_16082,N_16015);
nand U16708 (N_16708,N_16197,N_16284);
or U16709 (N_16709,N_16053,N_16145);
and U16710 (N_16710,N_16421,N_16311);
nor U16711 (N_16711,N_16414,N_16385);
and U16712 (N_16712,N_16219,N_16289);
or U16713 (N_16713,N_16143,N_16126);
or U16714 (N_16714,N_16221,N_16307);
nor U16715 (N_16715,N_16243,N_16005);
xor U16716 (N_16716,N_16095,N_16331);
nor U16717 (N_16717,N_16429,N_16478);
or U16718 (N_16718,N_16361,N_16384);
or U16719 (N_16719,N_16094,N_16088);
xor U16720 (N_16720,N_16161,N_16436);
xor U16721 (N_16721,N_16228,N_16259);
and U16722 (N_16722,N_16303,N_16260);
and U16723 (N_16723,N_16496,N_16076);
or U16724 (N_16724,N_16047,N_16086);
and U16725 (N_16725,N_16253,N_16208);
nand U16726 (N_16726,N_16183,N_16369);
or U16727 (N_16727,N_16362,N_16012);
nand U16728 (N_16728,N_16180,N_16100);
or U16729 (N_16729,N_16164,N_16014);
xor U16730 (N_16730,N_16193,N_16393);
nor U16731 (N_16731,N_16463,N_16346);
and U16732 (N_16732,N_16297,N_16081);
or U16733 (N_16733,N_16337,N_16232);
and U16734 (N_16734,N_16072,N_16364);
xnor U16735 (N_16735,N_16368,N_16338);
xor U16736 (N_16736,N_16203,N_16220);
nand U16737 (N_16737,N_16031,N_16313);
and U16738 (N_16738,N_16036,N_16410);
nand U16739 (N_16739,N_16171,N_16144);
nor U16740 (N_16740,N_16491,N_16115);
nor U16741 (N_16741,N_16089,N_16028);
xor U16742 (N_16742,N_16241,N_16006);
and U16743 (N_16743,N_16048,N_16365);
and U16744 (N_16744,N_16041,N_16045);
or U16745 (N_16745,N_16177,N_16287);
xor U16746 (N_16746,N_16025,N_16322);
nor U16747 (N_16747,N_16306,N_16325);
nor U16748 (N_16748,N_16216,N_16160);
nor U16749 (N_16749,N_16104,N_16212);
nand U16750 (N_16750,N_16343,N_16473);
nand U16751 (N_16751,N_16266,N_16195);
nand U16752 (N_16752,N_16289,N_16304);
xnor U16753 (N_16753,N_16042,N_16268);
and U16754 (N_16754,N_16068,N_16229);
nand U16755 (N_16755,N_16473,N_16117);
nor U16756 (N_16756,N_16025,N_16081);
nand U16757 (N_16757,N_16475,N_16354);
or U16758 (N_16758,N_16431,N_16343);
nor U16759 (N_16759,N_16121,N_16274);
nand U16760 (N_16760,N_16049,N_16133);
nand U16761 (N_16761,N_16365,N_16215);
nand U16762 (N_16762,N_16065,N_16317);
nand U16763 (N_16763,N_16158,N_16463);
xor U16764 (N_16764,N_16386,N_16416);
and U16765 (N_16765,N_16396,N_16415);
and U16766 (N_16766,N_16013,N_16152);
nand U16767 (N_16767,N_16352,N_16209);
nor U16768 (N_16768,N_16238,N_16231);
or U16769 (N_16769,N_16202,N_16242);
nand U16770 (N_16770,N_16398,N_16336);
or U16771 (N_16771,N_16333,N_16214);
nand U16772 (N_16772,N_16185,N_16196);
or U16773 (N_16773,N_16274,N_16186);
nor U16774 (N_16774,N_16351,N_16132);
or U16775 (N_16775,N_16398,N_16374);
nand U16776 (N_16776,N_16423,N_16275);
and U16777 (N_16777,N_16144,N_16161);
nand U16778 (N_16778,N_16074,N_16321);
xor U16779 (N_16779,N_16119,N_16260);
xnor U16780 (N_16780,N_16001,N_16331);
nor U16781 (N_16781,N_16417,N_16148);
nor U16782 (N_16782,N_16175,N_16037);
and U16783 (N_16783,N_16163,N_16491);
nor U16784 (N_16784,N_16030,N_16213);
and U16785 (N_16785,N_16239,N_16161);
nor U16786 (N_16786,N_16323,N_16496);
nor U16787 (N_16787,N_16267,N_16414);
and U16788 (N_16788,N_16489,N_16195);
nand U16789 (N_16789,N_16428,N_16039);
or U16790 (N_16790,N_16149,N_16249);
xor U16791 (N_16791,N_16062,N_16144);
xnor U16792 (N_16792,N_16315,N_16078);
and U16793 (N_16793,N_16082,N_16447);
nand U16794 (N_16794,N_16094,N_16466);
or U16795 (N_16795,N_16214,N_16497);
xor U16796 (N_16796,N_16111,N_16103);
nor U16797 (N_16797,N_16053,N_16113);
and U16798 (N_16798,N_16050,N_16495);
xor U16799 (N_16799,N_16404,N_16373);
nor U16800 (N_16800,N_16221,N_16425);
nor U16801 (N_16801,N_16103,N_16362);
or U16802 (N_16802,N_16396,N_16067);
nand U16803 (N_16803,N_16077,N_16097);
nand U16804 (N_16804,N_16170,N_16302);
nand U16805 (N_16805,N_16097,N_16197);
or U16806 (N_16806,N_16325,N_16099);
nand U16807 (N_16807,N_16238,N_16245);
and U16808 (N_16808,N_16226,N_16254);
xnor U16809 (N_16809,N_16050,N_16371);
nor U16810 (N_16810,N_16334,N_16273);
or U16811 (N_16811,N_16495,N_16481);
and U16812 (N_16812,N_16286,N_16061);
or U16813 (N_16813,N_16400,N_16264);
and U16814 (N_16814,N_16150,N_16003);
xor U16815 (N_16815,N_16393,N_16050);
nand U16816 (N_16816,N_16342,N_16057);
and U16817 (N_16817,N_16154,N_16357);
xnor U16818 (N_16818,N_16445,N_16377);
and U16819 (N_16819,N_16046,N_16114);
and U16820 (N_16820,N_16247,N_16296);
or U16821 (N_16821,N_16086,N_16053);
xnor U16822 (N_16822,N_16256,N_16475);
nand U16823 (N_16823,N_16453,N_16355);
nor U16824 (N_16824,N_16222,N_16323);
xnor U16825 (N_16825,N_16400,N_16224);
nor U16826 (N_16826,N_16408,N_16496);
or U16827 (N_16827,N_16059,N_16151);
and U16828 (N_16828,N_16383,N_16191);
nor U16829 (N_16829,N_16495,N_16447);
nor U16830 (N_16830,N_16020,N_16274);
nor U16831 (N_16831,N_16065,N_16150);
and U16832 (N_16832,N_16399,N_16039);
xnor U16833 (N_16833,N_16341,N_16179);
and U16834 (N_16834,N_16113,N_16447);
or U16835 (N_16835,N_16323,N_16298);
and U16836 (N_16836,N_16398,N_16012);
and U16837 (N_16837,N_16412,N_16355);
nor U16838 (N_16838,N_16413,N_16177);
nor U16839 (N_16839,N_16475,N_16012);
and U16840 (N_16840,N_16246,N_16466);
nor U16841 (N_16841,N_16276,N_16471);
nor U16842 (N_16842,N_16399,N_16226);
and U16843 (N_16843,N_16464,N_16397);
nor U16844 (N_16844,N_16097,N_16110);
nor U16845 (N_16845,N_16135,N_16410);
nor U16846 (N_16846,N_16084,N_16203);
xnor U16847 (N_16847,N_16051,N_16349);
nor U16848 (N_16848,N_16069,N_16334);
nand U16849 (N_16849,N_16394,N_16337);
nor U16850 (N_16850,N_16057,N_16025);
nand U16851 (N_16851,N_16139,N_16446);
xnor U16852 (N_16852,N_16407,N_16247);
or U16853 (N_16853,N_16020,N_16064);
or U16854 (N_16854,N_16337,N_16275);
and U16855 (N_16855,N_16048,N_16409);
and U16856 (N_16856,N_16190,N_16073);
xor U16857 (N_16857,N_16065,N_16437);
nor U16858 (N_16858,N_16374,N_16179);
nor U16859 (N_16859,N_16486,N_16078);
and U16860 (N_16860,N_16379,N_16168);
xor U16861 (N_16861,N_16097,N_16050);
nand U16862 (N_16862,N_16277,N_16096);
xnor U16863 (N_16863,N_16092,N_16258);
xor U16864 (N_16864,N_16325,N_16269);
xor U16865 (N_16865,N_16325,N_16158);
and U16866 (N_16866,N_16049,N_16298);
nor U16867 (N_16867,N_16382,N_16017);
nor U16868 (N_16868,N_16087,N_16371);
xor U16869 (N_16869,N_16041,N_16175);
or U16870 (N_16870,N_16317,N_16172);
or U16871 (N_16871,N_16319,N_16378);
nor U16872 (N_16872,N_16448,N_16326);
nor U16873 (N_16873,N_16307,N_16360);
xor U16874 (N_16874,N_16275,N_16244);
xnor U16875 (N_16875,N_16490,N_16480);
or U16876 (N_16876,N_16387,N_16184);
nand U16877 (N_16877,N_16172,N_16323);
nor U16878 (N_16878,N_16118,N_16357);
nor U16879 (N_16879,N_16369,N_16256);
xor U16880 (N_16880,N_16081,N_16288);
xnor U16881 (N_16881,N_16338,N_16405);
nor U16882 (N_16882,N_16123,N_16152);
nand U16883 (N_16883,N_16114,N_16291);
nor U16884 (N_16884,N_16126,N_16213);
or U16885 (N_16885,N_16221,N_16156);
xnor U16886 (N_16886,N_16043,N_16445);
or U16887 (N_16887,N_16142,N_16312);
nand U16888 (N_16888,N_16021,N_16341);
nand U16889 (N_16889,N_16492,N_16027);
and U16890 (N_16890,N_16317,N_16253);
xnor U16891 (N_16891,N_16133,N_16316);
xnor U16892 (N_16892,N_16419,N_16424);
nor U16893 (N_16893,N_16262,N_16162);
xnor U16894 (N_16894,N_16343,N_16302);
nand U16895 (N_16895,N_16361,N_16033);
nand U16896 (N_16896,N_16453,N_16231);
or U16897 (N_16897,N_16454,N_16201);
nand U16898 (N_16898,N_16487,N_16041);
xnor U16899 (N_16899,N_16499,N_16292);
nor U16900 (N_16900,N_16244,N_16031);
or U16901 (N_16901,N_16305,N_16210);
nor U16902 (N_16902,N_16219,N_16361);
nor U16903 (N_16903,N_16484,N_16344);
nor U16904 (N_16904,N_16011,N_16170);
nand U16905 (N_16905,N_16175,N_16233);
xor U16906 (N_16906,N_16384,N_16050);
nor U16907 (N_16907,N_16254,N_16107);
or U16908 (N_16908,N_16155,N_16226);
xnor U16909 (N_16909,N_16416,N_16457);
or U16910 (N_16910,N_16307,N_16342);
nor U16911 (N_16911,N_16266,N_16274);
and U16912 (N_16912,N_16089,N_16002);
xnor U16913 (N_16913,N_16325,N_16138);
nor U16914 (N_16914,N_16069,N_16058);
and U16915 (N_16915,N_16195,N_16090);
nor U16916 (N_16916,N_16475,N_16254);
and U16917 (N_16917,N_16443,N_16329);
nand U16918 (N_16918,N_16012,N_16218);
nand U16919 (N_16919,N_16274,N_16001);
xor U16920 (N_16920,N_16483,N_16323);
or U16921 (N_16921,N_16011,N_16067);
xor U16922 (N_16922,N_16211,N_16049);
and U16923 (N_16923,N_16405,N_16123);
or U16924 (N_16924,N_16389,N_16074);
xor U16925 (N_16925,N_16493,N_16118);
nand U16926 (N_16926,N_16120,N_16421);
and U16927 (N_16927,N_16058,N_16335);
and U16928 (N_16928,N_16151,N_16002);
or U16929 (N_16929,N_16123,N_16048);
xnor U16930 (N_16930,N_16030,N_16375);
nand U16931 (N_16931,N_16335,N_16304);
and U16932 (N_16932,N_16019,N_16015);
xor U16933 (N_16933,N_16428,N_16182);
or U16934 (N_16934,N_16135,N_16127);
or U16935 (N_16935,N_16339,N_16226);
nand U16936 (N_16936,N_16012,N_16084);
xnor U16937 (N_16937,N_16250,N_16117);
and U16938 (N_16938,N_16358,N_16337);
or U16939 (N_16939,N_16160,N_16081);
or U16940 (N_16940,N_16361,N_16059);
and U16941 (N_16941,N_16125,N_16012);
nand U16942 (N_16942,N_16383,N_16073);
xnor U16943 (N_16943,N_16499,N_16449);
or U16944 (N_16944,N_16391,N_16203);
and U16945 (N_16945,N_16064,N_16140);
nand U16946 (N_16946,N_16330,N_16166);
or U16947 (N_16947,N_16046,N_16493);
nand U16948 (N_16948,N_16043,N_16333);
or U16949 (N_16949,N_16232,N_16457);
or U16950 (N_16950,N_16348,N_16088);
nand U16951 (N_16951,N_16005,N_16230);
or U16952 (N_16952,N_16327,N_16124);
xor U16953 (N_16953,N_16078,N_16403);
nor U16954 (N_16954,N_16418,N_16499);
and U16955 (N_16955,N_16473,N_16120);
nor U16956 (N_16956,N_16261,N_16124);
nor U16957 (N_16957,N_16119,N_16092);
or U16958 (N_16958,N_16124,N_16282);
or U16959 (N_16959,N_16105,N_16355);
nand U16960 (N_16960,N_16347,N_16182);
and U16961 (N_16961,N_16027,N_16060);
or U16962 (N_16962,N_16027,N_16444);
nor U16963 (N_16963,N_16434,N_16157);
xor U16964 (N_16964,N_16185,N_16066);
or U16965 (N_16965,N_16057,N_16267);
xor U16966 (N_16966,N_16309,N_16107);
xor U16967 (N_16967,N_16120,N_16460);
and U16968 (N_16968,N_16468,N_16325);
xnor U16969 (N_16969,N_16311,N_16204);
nand U16970 (N_16970,N_16197,N_16460);
or U16971 (N_16971,N_16491,N_16391);
nand U16972 (N_16972,N_16029,N_16305);
xnor U16973 (N_16973,N_16378,N_16347);
and U16974 (N_16974,N_16203,N_16334);
nor U16975 (N_16975,N_16459,N_16208);
or U16976 (N_16976,N_16051,N_16287);
xnor U16977 (N_16977,N_16224,N_16012);
nor U16978 (N_16978,N_16094,N_16487);
nor U16979 (N_16979,N_16369,N_16050);
or U16980 (N_16980,N_16226,N_16241);
nand U16981 (N_16981,N_16408,N_16282);
xor U16982 (N_16982,N_16392,N_16499);
nor U16983 (N_16983,N_16007,N_16430);
nor U16984 (N_16984,N_16243,N_16175);
xnor U16985 (N_16985,N_16291,N_16011);
xor U16986 (N_16986,N_16348,N_16254);
or U16987 (N_16987,N_16167,N_16296);
or U16988 (N_16988,N_16126,N_16480);
and U16989 (N_16989,N_16251,N_16102);
or U16990 (N_16990,N_16153,N_16103);
or U16991 (N_16991,N_16332,N_16340);
xor U16992 (N_16992,N_16246,N_16162);
or U16993 (N_16993,N_16349,N_16296);
or U16994 (N_16994,N_16077,N_16225);
or U16995 (N_16995,N_16337,N_16081);
and U16996 (N_16996,N_16422,N_16220);
or U16997 (N_16997,N_16196,N_16180);
xnor U16998 (N_16998,N_16173,N_16391);
and U16999 (N_16999,N_16477,N_16364);
nand U17000 (N_17000,N_16963,N_16820);
nor U17001 (N_17001,N_16573,N_16922);
nor U17002 (N_17002,N_16890,N_16586);
nor U17003 (N_17003,N_16635,N_16813);
nor U17004 (N_17004,N_16726,N_16897);
or U17005 (N_17005,N_16787,N_16530);
and U17006 (N_17006,N_16574,N_16692);
nand U17007 (N_17007,N_16524,N_16699);
nor U17008 (N_17008,N_16650,N_16878);
nor U17009 (N_17009,N_16625,N_16522);
and U17010 (N_17010,N_16601,N_16976);
and U17011 (N_17011,N_16604,N_16858);
nand U17012 (N_17012,N_16546,N_16771);
nor U17013 (N_17013,N_16549,N_16844);
nor U17014 (N_17014,N_16930,N_16893);
and U17015 (N_17015,N_16600,N_16747);
xnor U17016 (N_17016,N_16543,N_16717);
nand U17017 (N_17017,N_16784,N_16521);
xor U17018 (N_17018,N_16518,N_16665);
or U17019 (N_17019,N_16672,N_16687);
and U17020 (N_17020,N_16989,N_16746);
nor U17021 (N_17021,N_16789,N_16790);
and U17022 (N_17022,N_16733,N_16594);
nand U17023 (N_17023,N_16811,N_16636);
nor U17024 (N_17024,N_16805,N_16690);
or U17025 (N_17025,N_16520,N_16760);
and U17026 (N_17026,N_16732,N_16857);
xnor U17027 (N_17027,N_16532,N_16703);
or U17028 (N_17028,N_16835,N_16599);
or U17029 (N_17029,N_16583,N_16705);
or U17030 (N_17030,N_16507,N_16580);
nor U17031 (N_17031,N_16772,N_16848);
nor U17032 (N_17032,N_16653,N_16924);
nand U17033 (N_17033,N_16548,N_16889);
or U17034 (N_17034,N_16998,N_16560);
and U17035 (N_17035,N_16801,N_16983);
and U17036 (N_17036,N_16707,N_16730);
or U17037 (N_17037,N_16553,N_16879);
nand U17038 (N_17038,N_16934,N_16807);
nand U17039 (N_17039,N_16777,N_16613);
nor U17040 (N_17040,N_16788,N_16815);
nor U17041 (N_17041,N_16585,N_16929);
and U17042 (N_17042,N_16993,N_16756);
and U17043 (N_17043,N_16939,N_16693);
nor U17044 (N_17044,N_16729,N_16723);
nor U17045 (N_17045,N_16995,N_16617);
or U17046 (N_17046,N_16947,N_16905);
or U17047 (N_17047,N_16849,N_16626);
or U17048 (N_17048,N_16716,N_16712);
xor U17049 (N_17049,N_16839,N_16821);
nand U17050 (N_17050,N_16845,N_16688);
nand U17051 (N_17051,N_16903,N_16972);
or U17052 (N_17052,N_16644,N_16851);
nand U17053 (N_17053,N_16720,N_16736);
nor U17054 (N_17054,N_16658,N_16834);
and U17055 (N_17055,N_16779,N_16647);
nand U17056 (N_17056,N_16673,N_16555);
nor U17057 (N_17057,N_16973,N_16966);
nor U17058 (N_17058,N_16804,N_16775);
and U17059 (N_17059,N_16540,N_16591);
xor U17060 (N_17060,N_16798,N_16877);
nor U17061 (N_17061,N_16757,N_16765);
xor U17062 (N_17062,N_16984,N_16533);
and U17063 (N_17063,N_16501,N_16944);
xor U17064 (N_17064,N_16901,N_16609);
nor U17065 (N_17065,N_16826,N_16861);
or U17066 (N_17066,N_16975,N_16842);
or U17067 (N_17067,N_16515,N_16809);
or U17068 (N_17068,N_16734,N_16743);
nand U17069 (N_17069,N_16867,N_16981);
nor U17070 (N_17070,N_16702,N_16968);
and U17071 (N_17071,N_16987,N_16920);
or U17072 (N_17072,N_16959,N_16711);
nor U17073 (N_17073,N_16564,N_16847);
nor U17074 (N_17074,N_16923,N_16953);
xor U17075 (N_17075,N_16950,N_16916);
xor U17076 (N_17076,N_16892,N_16886);
and U17077 (N_17077,N_16742,N_16952);
nor U17078 (N_17078,N_16840,N_16683);
nand U17079 (N_17079,N_16651,N_16529);
xnor U17080 (N_17080,N_16869,N_16718);
and U17081 (N_17081,N_16608,N_16750);
and U17082 (N_17082,N_16830,N_16744);
and U17083 (N_17083,N_16855,N_16865);
nor U17084 (N_17084,N_16631,N_16969);
or U17085 (N_17085,N_16517,N_16866);
or U17086 (N_17086,N_16514,N_16639);
xnor U17087 (N_17087,N_16587,N_16510);
xor U17088 (N_17088,N_16691,N_16713);
nor U17089 (N_17089,N_16628,N_16979);
and U17090 (N_17090,N_16856,N_16676);
or U17091 (N_17091,N_16695,N_16971);
nand U17092 (N_17092,N_16577,N_16803);
nand U17093 (N_17093,N_16814,N_16662);
or U17094 (N_17094,N_16942,N_16921);
or U17095 (N_17095,N_16933,N_16843);
xnor U17096 (N_17096,N_16547,N_16937);
and U17097 (N_17097,N_16770,N_16774);
xnor U17098 (N_17098,N_16967,N_16722);
nand U17099 (N_17099,N_16895,N_16649);
xnor U17100 (N_17100,N_16806,N_16951);
and U17101 (N_17101,N_16566,N_16738);
nand U17102 (N_17102,N_16615,N_16563);
nand U17103 (N_17103,N_16641,N_16838);
xor U17104 (N_17104,N_16519,N_16970);
xnor U17105 (N_17105,N_16876,N_16748);
xnor U17106 (N_17106,N_16629,N_16768);
or U17107 (N_17107,N_16926,N_16614);
or U17108 (N_17108,N_16864,N_16709);
nand U17109 (N_17109,N_16595,N_16525);
nor U17110 (N_17110,N_16887,N_16539);
or U17111 (N_17111,N_16696,N_16643);
xnor U17112 (N_17112,N_16745,N_16831);
nor U17113 (N_17113,N_16909,N_16816);
and U17114 (N_17114,N_16528,N_16759);
or U17115 (N_17115,N_16582,N_16607);
xor U17116 (N_17116,N_16885,N_16850);
xor U17117 (N_17117,N_16764,N_16940);
xnor U17118 (N_17118,N_16965,N_16818);
nor U17119 (N_17119,N_16541,N_16556);
and U17120 (N_17120,N_16990,N_16700);
or U17121 (N_17121,N_16915,N_16648);
nand U17122 (N_17122,N_16630,N_16754);
xnor U17123 (N_17123,N_16516,N_16872);
xnor U17124 (N_17124,N_16841,N_16616);
nor U17125 (N_17125,N_16502,N_16946);
nor U17126 (N_17126,N_16557,N_16881);
and U17127 (N_17127,N_16802,N_16982);
nand U17128 (N_17128,N_16682,N_16545);
xor U17129 (N_17129,N_16785,N_16656);
and U17130 (N_17130,N_16677,N_16668);
and U17131 (N_17131,N_16810,N_16646);
xnor U17132 (N_17132,N_16860,N_16581);
and U17133 (N_17133,N_16936,N_16898);
or U17134 (N_17134,N_16906,N_16919);
or U17135 (N_17135,N_16602,N_16783);
nor U17136 (N_17136,N_16761,N_16578);
nand U17137 (N_17137,N_16910,N_16731);
or U17138 (N_17138,N_16917,N_16884);
nor U17139 (N_17139,N_16911,N_16506);
nand U17140 (N_17140,N_16531,N_16657);
and U17141 (N_17141,N_16766,N_16606);
or U17142 (N_17142,N_16523,N_16735);
and U17143 (N_17143,N_16776,N_16852);
and U17144 (N_17144,N_16812,N_16535);
and U17145 (N_17145,N_16576,N_16554);
and U17146 (N_17146,N_16584,N_16786);
or U17147 (N_17147,N_16873,N_16503);
nor U17148 (N_17148,N_16710,N_16755);
and U17149 (N_17149,N_16882,N_16961);
nand U17150 (N_17150,N_16935,N_16661);
xor U17151 (N_17151,N_16931,N_16862);
nor U17152 (N_17152,N_16561,N_16592);
nor U17153 (N_17153,N_16603,N_16896);
and U17154 (N_17154,N_16589,N_16827);
nand U17155 (N_17155,N_16945,N_16902);
nand U17156 (N_17156,N_16833,N_16596);
and U17157 (N_17157,N_16575,N_16751);
nor U17158 (N_17158,N_16778,N_16551);
and U17159 (N_17159,N_16954,N_16612);
xnor U17160 (N_17160,N_16621,N_16899);
nor U17161 (N_17161,N_16670,N_16654);
nor U17162 (N_17162,N_16708,N_16704);
nor U17163 (N_17163,N_16509,N_16763);
and U17164 (N_17164,N_16664,N_16978);
nor U17165 (N_17165,N_16832,N_16634);
and U17166 (N_17166,N_16590,N_16666);
and U17167 (N_17167,N_16627,N_16997);
nand U17168 (N_17168,N_16598,N_16562);
or U17169 (N_17169,N_16991,N_16859);
nand U17170 (N_17170,N_16620,N_16558);
or U17171 (N_17171,N_16537,N_16640);
and U17172 (N_17172,N_16660,N_16846);
xnor U17173 (N_17173,N_16674,N_16829);
xnor U17174 (N_17174,N_16956,N_16671);
and U17175 (N_17175,N_16828,N_16655);
nand U17176 (N_17176,N_16526,N_16863);
and U17177 (N_17177,N_16588,N_16943);
nand U17178 (N_17178,N_16891,N_16737);
and U17179 (N_17179,N_16955,N_16837);
nand U17180 (N_17180,N_16753,N_16883);
or U17181 (N_17181,N_16611,N_16977);
or U17182 (N_17182,N_16605,N_16619);
or U17183 (N_17183,N_16793,N_16888);
and U17184 (N_17184,N_16675,N_16853);
xor U17185 (N_17185,N_16534,N_16685);
and U17186 (N_17186,N_16697,N_16918);
or U17187 (N_17187,N_16679,N_16957);
or U17188 (N_17188,N_16941,N_16767);
xor U17189 (N_17189,N_16569,N_16868);
xnor U17190 (N_17190,N_16728,N_16727);
nor U17191 (N_17191,N_16706,N_16938);
nor U17192 (N_17192,N_16715,N_16571);
and U17193 (N_17193,N_16913,N_16962);
or U17194 (N_17194,N_16817,N_16663);
or U17195 (N_17195,N_16854,N_16752);
xor U17196 (N_17196,N_16544,N_16799);
xor U17197 (N_17197,N_16513,N_16570);
and U17198 (N_17198,N_16652,N_16637);
or U17199 (N_17199,N_16508,N_16659);
nor U17200 (N_17200,N_16536,N_16928);
or U17201 (N_17201,N_16638,N_16678);
nand U17202 (N_17202,N_16684,N_16932);
xor U17203 (N_17203,N_16741,N_16996);
nor U17204 (N_17204,N_16870,N_16681);
and U17205 (N_17205,N_16622,N_16568);
or U17206 (N_17206,N_16822,N_16958);
and U17207 (N_17207,N_16904,N_16819);
and U17208 (N_17208,N_16797,N_16511);
xor U17209 (N_17209,N_16550,N_16632);
xnor U17210 (N_17210,N_16624,N_16875);
and U17211 (N_17211,N_16565,N_16642);
nand U17212 (N_17212,N_16758,N_16504);
nor U17213 (N_17213,N_16894,N_16986);
or U17214 (N_17214,N_16773,N_16999);
xor U17215 (N_17215,N_16988,N_16908);
nand U17216 (N_17216,N_16721,N_16974);
nand U17217 (N_17217,N_16597,N_16762);
nand U17218 (N_17218,N_16552,N_16694);
and U17219 (N_17219,N_16980,N_16572);
nand U17220 (N_17220,N_16714,N_16680);
xor U17221 (N_17221,N_16542,N_16964);
and U17222 (N_17222,N_16960,N_16538);
or U17223 (N_17223,N_16800,N_16836);
xnor U17224 (N_17224,N_16701,N_16782);
or U17225 (N_17225,N_16880,N_16725);
or U17226 (N_17226,N_16985,N_16739);
or U17227 (N_17227,N_16780,N_16900);
and U17228 (N_17228,N_16795,N_16825);
xnor U17229 (N_17229,N_16912,N_16992);
and U17230 (N_17230,N_16667,N_16874);
nand U17231 (N_17231,N_16505,N_16740);
and U17232 (N_17232,N_16769,N_16669);
nand U17233 (N_17233,N_16567,N_16633);
and U17234 (N_17234,N_16610,N_16618);
xnor U17235 (N_17235,N_16794,N_16623);
xnor U17236 (N_17236,N_16871,N_16593);
nor U17237 (N_17237,N_16796,N_16698);
xor U17238 (N_17238,N_16792,N_16948);
and U17239 (N_17239,N_16994,N_16914);
or U17240 (N_17240,N_16500,N_16823);
nand U17241 (N_17241,N_16824,N_16689);
and U17242 (N_17242,N_16645,N_16949);
nor U17243 (N_17243,N_16781,N_16749);
xnor U17244 (N_17244,N_16791,N_16925);
nor U17245 (N_17245,N_16579,N_16724);
nor U17246 (N_17246,N_16808,N_16927);
nor U17247 (N_17247,N_16512,N_16719);
xor U17248 (N_17248,N_16907,N_16559);
and U17249 (N_17249,N_16686,N_16527);
and U17250 (N_17250,N_16926,N_16786);
nand U17251 (N_17251,N_16949,N_16948);
xnor U17252 (N_17252,N_16654,N_16752);
or U17253 (N_17253,N_16692,N_16891);
and U17254 (N_17254,N_16983,N_16738);
xor U17255 (N_17255,N_16731,N_16696);
or U17256 (N_17256,N_16592,N_16549);
xnor U17257 (N_17257,N_16969,N_16922);
and U17258 (N_17258,N_16536,N_16921);
nor U17259 (N_17259,N_16990,N_16806);
or U17260 (N_17260,N_16784,N_16730);
nand U17261 (N_17261,N_16906,N_16822);
and U17262 (N_17262,N_16869,N_16688);
or U17263 (N_17263,N_16802,N_16746);
xor U17264 (N_17264,N_16891,N_16768);
nand U17265 (N_17265,N_16992,N_16677);
and U17266 (N_17266,N_16544,N_16926);
and U17267 (N_17267,N_16762,N_16683);
or U17268 (N_17268,N_16977,N_16789);
xor U17269 (N_17269,N_16698,N_16995);
nand U17270 (N_17270,N_16991,N_16976);
or U17271 (N_17271,N_16771,N_16665);
nor U17272 (N_17272,N_16862,N_16702);
nor U17273 (N_17273,N_16870,N_16718);
nor U17274 (N_17274,N_16942,N_16956);
and U17275 (N_17275,N_16693,N_16837);
nand U17276 (N_17276,N_16909,N_16915);
or U17277 (N_17277,N_16973,N_16778);
nor U17278 (N_17278,N_16902,N_16670);
nand U17279 (N_17279,N_16528,N_16560);
or U17280 (N_17280,N_16724,N_16752);
xor U17281 (N_17281,N_16818,N_16919);
xor U17282 (N_17282,N_16525,N_16640);
nor U17283 (N_17283,N_16723,N_16934);
and U17284 (N_17284,N_16698,N_16555);
and U17285 (N_17285,N_16870,N_16753);
or U17286 (N_17286,N_16539,N_16868);
nand U17287 (N_17287,N_16684,N_16885);
or U17288 (N_17288,N_16623,N_16950);
or U17289 (N_17289,N_16877,N_16700);
nand U17290 (N_17290,N_16601,N_16858);
or U17291 (N_17291,N_16689,N_16770);
and U17292 (N_17292,N_16858,N_16637);
xor U17293 (N_17293,N_16977,N_16912);
nor U17294 (N_17294,N_16880,N_16858);
nor U17295 (N_17295,N_16855,N_16640);
or U17296 (N_17296,N_16979,N_16608);
nor U17297 (N_17297,N_16805,N_16507);
xnor U17298 (N_17298,N_16520,N_16601);
nor U17299 (N_17299,N_16932,N_16941);
xor U17300 (N_17300,N_16939,N_16918);
nand U17301 (N_17301,N_16997,N_16932);
or U17302 (N_17302,N_16789,N_16707);
nor U17303 (N_17303,N_16857,N_16615);
and U17304 (N_17304,N_16613,N_16810);
and U17305 (N_17305,N_16939,N_16694);
and U17306 (N_17306,N_16999,N_16771);
and U17307 (N_17307,N_16929,N_16644);
or U17308 (N_17308,N_16929,N_16834);
nand U17309 (N_17309,N_16976,N_16577);
xnor U17310 (N_17310,N_16697,N_16879);
nand U17311 (N_17311,N_16739,N_16660);
nand U17312 (N_17312,N_16902,N_16887);
xnor U17313 (N_17313,N_16960,N_16657);
xnor U17314 (N_17314,N_16639,N_16947);
or U17315 (N_17315,N_16853,N_16934);
nand U17316 (N_17316,N_16915,N_16615);
nand U17317 (N_17317,N_16943,N_16793);
or U17318 (N_17318,N_16791,N_16559);
or U17319 (N_17319,N_16725,N_16836);
and U17320 (N_17320,N_16986,N_16735);
nor U17321 (N_17321,N_16642,N_16922);
nand U17322 (N_17322,N_16986,N_16965);
nor U17323 (N_17323,N_16516,N_16684);
nand U17324 (N_17324,N_16528,N_16732);
and U17325 (N_17325,N_16620,N_16697);
nand U17326 (N_17326,N_16943,N_16743);
nor U17327 (N_17327,N_16668,N_16728);
xor U17328 (N_17328,N_16615,N_16659);
and U17329 (N_17329,N_16739,N_16696);
nand U17330 (N_17330,N_16933,N_16890);
nand U17331 (N_17331,N_16969,N_16671);
or U17332 (N_17332,N_16777,N_16556);
nor U17333 (N_17333,N_16627,N_16582);
xor U17334 (N_17334,N_16969,N_16583);
nor U17335 (N_17335,N_16759,N_16548);
and U17336 (N_17336,N_16869,N_16753);
nor U17337 (N_17337,N_16812,N_16902);
xor U17338 (N_17338,N_16875,N_16882);
and U17339 (N_17339,N_16643,N_16542);
nor U17340 (N_17340,N_16849,N_16860);
or U17341 (N_17341,N_16801,N_16854);
xor U17342 (N_17342,N_16915,N_16598);
and U17343 (N_17343,N_16507,N_16965);
nand U17344 (N_17344,N_16993,N_16926);
xor U17345 (N_17345,N_16780,N_16636);
nand U17346 (N_17346,N_16956,N_16528);
and U17347 (N_17347,N_16728,N_16814);
xnor U17348 (N_17348,N_16891,N_16585);
and U17349 (N_17349,N_16613,N_16950);
xnor U17350 (N_17350,N_16917,N_16792);
or U17351 (N_17351,N_16753,N_16990);
nand U17352 (N_17352,N_16619,N_16635);
nor U17353 (N_17353,N_16509,N_16588);
or U17354 (N_17354,N_16985,N_16526);
xor U17355 (N_17355,N_16789,N_16832);
nand U17356 (N_17356,N_16589,N_16612);
or U17357 (N_17357,N_16798,N_16576);
nor U17358 (N_17358,N_16763,N_16603);
xnor U17359 (N_17359,N_16956,N_16831);
or U17360 (N_17360,N_16954,N_16966);
or U17361 (N_17361,N_16751,N_16847);
xor U17362 (N_17362,N_16954,N_16773);
nand U17363 (N_17363,N_16827,N_16814);
and U17364 (N_17364,N_16671,N_16814);
nand U17365 (N_17365,N_16856,N_16532);
nor U17366 (N_17366,N_16571,N_16786);
nor U17367 (N_17367,N_16965,N_16875);
or U17368 (N_17368,N_16693,N_16752);
nor U17369 (N_17369,N_16815,N_16680);
or U17370 (N_17370,N_16701,N_16566);
nand U17371 (N_17371,N_16623,N_16592);
and U17372 (N_17372,N_16719,N_16811);
nor U17373 (N_17373,N_16798,N_16651);
or U17374 (N_17374,N_16900,N_16655);
nor U17375 (N_17375,N_16920,N_16509);
nand U17376 (N_17376,N_16994,N_16946);
nand U17377 (N_17377,N_16645,N_16513);
nor U17378 (N_17378,N_16623,N_16649);
or U17379 (N_17379,N_16904,N_16811);
xor U17380 (N_17380,N_16908,N_16798);
and U17381 (N_17381,N_16767,N_16749);
nor U17382 (N_17382,N_16951,N_16553);
and U17383 (N_17383,N_16688,N_16886);
nand U17384 (N_17384,N_16515,N_16549);
nand U17385 (N_17385,N_16572,N_16965);
nand U17386 (N_17386,N_16653,N_16507);
nor U17387 (N_17387,N_16894,N_16832);
and U17388 (N_17388,N_16704,N_16811);
and U17389 (N_17389,N_16587,N_16650);
nand U17390 (N_17390,N_16691,N_16715);
and U17391 (N_17391,N_16779,N_16834);
nand U17392 (N_17392,N_16887,N_16780);
nor U17393 (N_17393,N_16573,N_16652);
or U17394 (N_17394,N_16657,N_16923);
or U17395 (N_17395,N_16967,N_16609);
or U17396 (N_17396,N_16748,N_16519);
nand U17397 (N_17397,N_16969,N_16837);
xnor U17398 (N_17398,N_16744,N_16716);
and U17399 (N_17399,N_16733,N_16881);
xor U17400 (N_17400,N_16726,N_16760);
or U17401 (N_17401,N_16693,N_16940);
nor U17402 (N_17402,N_16570,N_16543);
nand U17403 (N_17403,N_16503,N_16592);
nor U17404 (N_17404,N_16669,N_16815);
or U17405 (N_17405,N_16704,N_16554);
xnor U17406 (N_17406,N_16870,N_16964);
or U17407 (N_17407,N_16698,N_16966);
and U17408 (N_17408,N_16855,N_16963);
xnor U17409 (N_17409,N_16796,N_16890);
or U17410 (N_17410,N_16863,N_16994);
nor U17411 (N_17411,N_16696,N_16629);
or U17412 (N_17412,N_16600,N_16779);
nand U17413 (N_17413,N_16638,N_16586);
nand U17414 (N_17414,N_16655,N_16891);
and U17415 (N_17415,N_16693,N_16567);
xnor U17416 (N_17416,N_16789,N_16628);
xor U17417 (N_17417,N_16631,N_16799);
nand U17418 (N_17418,N_16543,N_16657);
nor U17419 (N_17419,N_16698,N_16518);
xor U17420 (N_17420,N_16855,N_16944);
nor U17421 (N_17421,N_16749,N_16680);
nor U17422 (N_17422,N_16903,N_16796);
nand U17423 (N_17423,N_16789,N_16831);
nand U17424 (N_17424,N_16841,N_16843);
nand U17425 (N_17425,N_16812,N_16619);
and U17426 (N_17426,N_16526,N_16979);
nor U17427 (N_17427,N_16518,N_16620);
nand U17428 (N_17428,N_16730,N_16768);
and U17429 (N_17429,N_16793,N_16912);
nand U17430 (N_17430,N_16792,N_16974);
xor U17431 (N_17431,N_16737,N_16823);
or U17432 (N_17432,N_16983,N_16811);
nand U17433 (N_17433,N_16810,N_16606);
xnor U17434 (N_17434,N_16919,N_16557);
and U17435 (N_17435,N_16658,N_16588);
xor U17436 (N_17436,N_16848,N_16829);
or U17437 (N_17437,N_16526,N_16660);
or U17438 (N_17438,N_16886,N_16503);
or U17439 (N_17439,N_16706,N_16649);
xor U17440 (N_17440,N_16563,N_16817);
xnor U17441 (N_17441,N_16759,N_16510);
and U17442 (N_17442,N_16986,N_16626);
xor U17443 (N_17443,N_16673,N_16620);
nor U17444 (N_17444,N_16860,N_16750);
xor U17445 (N_17445,N_16949,N_16848);
or U17446 (N_17446,N_16764,N_16679);
or U17447 (N_17447,N_16718,N_16970);
or U17448 (N_17448,N_16933,N_16619);
nand U17449 (N_17449,N_16727,N_16575);
or U17450 (N_17450,N_16591,N_16542);
xnor U17451 (N_17451,N_16862,N_16753);
and U17452 (N_17452,N_16681,N_16863);
nor U17453 (N_17453,N_16795,N_16621);
nor U17454 (N_17454,N_16987,N_16703);
or U17455 (N_17455,N_16591,N_16734);
and U17456 (N_17456,N_16694,N_16735);
nor U17457 (N_17457,N_16584,N_16962);
nor U17458 (N_17458,N_16650,N_16505);
or U17459 (N_17459,N_16924,N_16776);
and U17460 (N_17460,N_16595,N_16532);
nand U17461 (N_17461,N_16574,N_16959);
nand U17462 (N_17462,N_16636,N_16767);
xnor U17463 (N_17463,N_16873,N_16874);
or U17464 (N_17464,N_16825,N_16512);
or U17465 (N_17465,N_16972,N_16719);
or U17466 (N_17466,N_16585,N_16640);
nor U17467 (N_17467,N_16860,N_16874);
xor U17468 (N_17468,N_16738,N_16559);
nand U17469 (N_17469,N_16534,N_16773);
or U17470 (N_17470,N_16840,N_16648);
and U17471 (N_17471,N_16886,N_16980);
nor U17472 (N_17472,N_16614,N_16852);
nand U17473 (N_17473,N_16669,N_16998);
xor U17474 (N_17474,N_16722,N_16796);
and U17475 (N_17475,N_16760,N_16586);
nor U17476 (N_17476,N_16503,N_16993);
xnor U17477 (N_17477,N_16515,N_16964);
or U17478 (N_17478,N_16678,N_16820);
and U17479 (N_17479,N_16835,N_16994);
and U17480 (N_17480,N_16965,N_16950);
and U17481 (N_17481,N_16756,N_16525);
nand U17482 (N_17482,N_16755,N_16782);
nor U17483 (N_17483,N_16703,N_16742);
nand U17484 (N_17484,N_16761,N_16992);
and U17485 (N_17485,N_16847,N_16858);
nand U17486 (N_17486,N_16812,N_16610);
or U17487 (N_17487,N_16690,N_16622);
xor U17488 (N_17488,N_16723,N_16514);
or U17489 (N_17489,N_16976,N_16589);
or U17490 (N_17490,N_16610,N_16937);
nor U17491 (N_17491,N_16691,N_16932);
and U17492 (N_17492,N_16756,N_16924);
nor U17493 (N_17493,N_16955,N_16853);
xor U17494 (N_17494,N_16705,N_16617);
and U17495 (N_17495,N_16557,N_16918);
or U17496 (N_17496,N_16899,N_16871);
and U17497 (N_17497,N_16633,N_16927);
nand U17498 (N_17498,N_16637,N_16846);
or U17499 (N_17499,N_16911,N_16960);
xor U17500 (N_17500,N_17217,N_17480);
nor U17501 (N_17501,N_17485,N_17095);
nand U17502 (N_17502,N_17055,N_17072);
nand U17503 (N_17503,N_17474,N_17331);
xnor U17504 (N_17504,N_17461,N_17394);
or U17505 (N_17505,N_17092,N_17449);
nor U17506 (N_17506,N_17407,N_17154);
nand U17507 (N_17507,N_17245,N_17191);
or U17508 (N_17508,N_17110,N_17412);
or U17509 (N_17509,N_17174,N_17113);
nand U17510 (N_17510,N_17439,N_17307);
or U17511 (N_17511,N_17128,N_17020);
nor U17512 (N_17512,N_17280,N_17123);
xnor U17513 (N_17513,N_17047,N_17045);
nor U17514 (N_17514,N_17012,N_17002);
xnor U17515 (N_17515,N_17211,N_17473);
nor U17516 (N_17516,N_17108,N_17301);
and U17517 (N_17517,N_17175,N_17414);
and U17518 (N_17518,N_17443,N_17308);
or U17519 (N_17519,N_17263,N_17456);
xor U17520 (N_17520,N_17167,N_17494);
nand U17521 (N_17521,N_17492,N_17448);
or U17522 (N_17522,N_17000,N_17185);
nor U17523 (N_17523,N_17080,N_17305);
and U17524 (N_17524,N_17006,N_17145);
and U17525 (N_17525,N_17415,N_17352);
and U17526 (N_17526,N_17322,N_17106);
nor U17527 (N_17527,N_17489,N_17139);
or U17528 (N_17528,N_17481,N_17083);
nand U17529 (N_17529,N_17382,N_17342);
or U17530 (N_17530,N_17241,N_17436);
and U17531 (N_17531,N_17287,N_17255);
xor U17532 (N_17532,N_17440,N_17058);
nand U17533 (N_17533,N_17484,N_17249);
xor U17534 (N_17534,N_17432,N_17441);
nor U17535 (N_17535,N_17413,N_17476);
and U17536 (N_17536,N_17446,N_17265);
or U17537 (N_17537,N_17435,N_17300);
or U17538 (N_17538,N_17437,N_17035);
and U17539 (N_17539,N_17262,N_17355);
nor U17540 (N_17540,N_17163,N_17421);
and U17541 (N_17541,N_17470,N_17096);
xnor U17542 (N_17542,N_17099,N_17483);
or U17543 (N_17543,N_17017,N_17289);
xor U17544 (N_17544,N_17431,N_17014);
xnor U17545 (N_17545,N_17335,N_17324);
and U17546 (N_17546,N_17445,N_17268);
nand U17547 (N_17547,N_17015,N_17100);
and U17548 (N_17548,N_17345,N_17024);
xor U17549 (N_17549,N_17005,N_17029);
nor U17550 (N_17550,N_17030,N_17019);
nand U17551 (N_17551,N_17471,N_17210);
or U17552 (N_17552,N_17201,N_17087);
and U17553 (N_17553,N_17061,N_17349);
and U17554 (N_17554,N_17142,N_17409);
and U17555 (N_17555,N_17433,N_17351);
and U17556 (N_17556,N_17276,N_17309);
nor U17557 (N_17557,N_17232,N_17404);
nor U17558 (N_17558,N_17057,N_17267);
nor U17559 (N_17559,N_17453,N_17042);
xnor U17560 (N_17560,N_17283,N_17156);
or U17561 (N_17561,N_17097,N_17078);
or U17562 (N_17562,N_17273,N_17266);
nand U17563 (N_17563,N_17358,N_17297);
nand U17564 (N_17564,N_17424,N_17229);
and U17565 (N_17565,N_17274,N_17281);
or U17566 (N_17566,N_17135,N_17009);
xor U17567 (N_17567,N_17094,N_17104);
or U17568 (N_17568,N_17391,N_17194);
or U17569 (N_17569,N_17395,N_17200);
xor U17570 (N_17570,N_17004,N_17271);
or U17571 (N_17571,N_17244,N_17362);
xnor U17572 (N_17572,N_17168,N_17296);
and U17573 (N_17573,N_17402,N_17184);
nand U17574 (N_17574,N_17220,N_17215);
xor U17575 (N_17575,N_17098,N_17170);
xnor U17576 (N_17576,N_17236,N_17347);
xnor U17577 (N_17577,N_17226,N_17089);
or U17578 (N_17578,N_17277,N_17288);
nand U17579 (N_17579,N_17121,N_17203);
xnor U17580 (N_17580,N_17105,N_17270);
xnor U17581 (N_17581,N_17356,N_17199);
or U17582 (N_17582,N_17176,N_17146);
xor U17583 (N_17583,N_17008,N_17482);
nor U17584 (N_17584,N_17472,N_17173);
xnor U17585 (N_17585,N_17411,N_17326);
xnor U17586 (N_17586,N_17137,N_17093);
and U17587 (N_17587,N_17187,N_17233);
or U17588 (N_17588,N_17148,N_17216);
nand U17589 (N_17589,N_17385,N_17074);
xor U17590 (N_17590,N_17278,N_17026);
nor U17591 (N_17591,N_17181,N_17333);
or U17592 (N_17592,N_17180,N_17069);
nor U17593 (N_17593,N_17272,N_17400);
and U17594 (N_17594,N_17222,N_17038);
or U17595 (N_17595,N_17380,N_17343);
nor U17596 (N_17596,N_17334,N_17041);
nand U17597 (N_17597,N_17299,N_17493);
or U17598 (N_17598,N_17423,N_17465);
xor U17599 (N_17599,N_17158,N_17136);
or U17600 (N_17600,N_17430,N_17021);
and U17601 (N_17601,N_17022,N_17348);
and U17602 (N_17602,N_17496,N_17040);
xor U17603 (N_17603,N_17056,N_17240);
nand U17604 (N_17604,N_17116,N_17112);
and U17605 (N_17605,N_17237,N_17235);
nor U17606 (N_17606,N_17328,N_17033);
xnor U17607 (N_17607,N_17081,N_17102);
and U17608 (N_17608,N_17279,N_17111);
and U17609 (N_17609,N_17457,N_17298);
nor U17610 (N_17610,N_17238,N_17143);
or U17611 (N_17611,N_17066,N_17067);
nand U17612 (N_17612,N_17442,N_17160);
xnor U17613 (N_17613,N_17486,N_17188);
nand U17614 (N_17614,N_17007,N_17150);
or U17615 (N_17615,N_17193,N_17312);
or U17616 (N_17616,N_17386,N_17250);
nand U17617 (N_17617,N_17153,N_17344);
or U17618 (N_17618,N_17214,N_17371);
nand U17619 (N_17619,N_17314,N_17016);
nor U17620 (N_17620,N_17151,N_17044);
nor U17621 (N_17621,N_17129,N_17257);
xnor U17622 (N_17622,N_17189,N_17183);
nand U17623 (N_17623,N_17406,N_17182);
or U17624 (N_17624,N_17479,N_17118);
and U17625 (N_17625,N_17375,N_17313);
xnor U17626 (N_17626,N_17316,N_17085);
nor U17627 (N_17627,N_17082,N_17219);
nand U17628 (N_17628,N_17339,N_17256);
xor U17629 (N_17629,N_17101,N_17392);
nor U17630 (N_17630,N_17107,N_17132);
nand U17631 (N_17631,N_17490,N_17252);
nand U17632 (N_17632,N_17166,N_17357);
or U17633 (N_17633,N_17310,N_17013);
nor U17634 (N_17634,N_17049,N_17125);
nand U17635 (N_17635,N_17171,N_17077);
or U17636 (N_17636,N_17463,N_17467);
xnor U17637 (N_17637,N_17259,N_17025);
and U17638 (N_17638,N_17155,N_17192);
xnor U17639 (N_17639,N_17388,N_17353);
nor U17640 (N_17640,N_17495,N_17018);
and U17641 (N_17641,N_17346,N_17379);
and U17642 (N_17642,N_17370,N_17223);
or U17643 (N_17643,N_17064,N_17198);
xor U17644 (N_17644,N_17294,N_17491);
nor U17645 (N_17645,N_17149,N_17381);
xnor U17646 (N_17646,N_17032,N_17140);
nor U17647 (N_17647,N_17464,N_17372);
and U17648 (N_17648,N_17043,N_17246);
xnor U17649 (N_17649,N_17239,N_17037);
or U17650 (N_17650,N_17084,N_17258);
nand U17651 (N_17651,N_17365,N_17039);
nor U17652 (N_17652,N_17213,N_17396);
nor U17653 (N_17653,N_17329,N_17420);
and U17654 (N_17654,N_17230,N_17304);
or U17655 (N_17655,N_17318,N_17152);
xor U17656 (N_17656,N_17050,N_17204);
or U17657 (N_17657,N_17419,N_17377);
or U17658 (N_17658,N_17186,N_17062);
or U17659 (N_17659,N_17434,N_17458);
nor U17660 (N_17660,N_17405,N_17315);
nand U17661 (N_17661,N_17410,N_17428);
or U17662 (N_17662,N_17251,N_17399);
nor U17663 (N_17663,N_17462,N_17284);
xor U17664 (N_17664,N_17207,N_17243);
xnor U17665 (N_17665,N_17059,N_17197);
or U17666 (N_17666,N_17374,N_17282);
xor U17667 (N_17667,N_17398,N_17133);
and U17668 (N_17668,N_17079,N_17206);
xnor U17669 (N_17669,N_17438,N_17141);
nor U17670 (N_17670,N_17427,N_17231);
or U17671 (N_17671,N_17366,N_17027);
or U17672 (N_17672,N_17401,N_17468);
and U17673 (N_17673,N_17360,N_17338);
or U17674 (N_17674,N_17327,N_17090);
and U17675 (N_17675,N_17368,N_17034);
nand U17676 (N_17676,N_17364,N_17103);
nor U17677 (N_17677,N_17162,N_17051);
nor U17678 (N_17678,N_17031,N_17383);
and U17679 (N_17679,N_17429,N_17450);
xnor U17680 (N_17680,N_17317,N_17178);
or U17681 (N_17681,N_17416,N_17403);
and U17682 (N_17682,N_17075,N_17157);
nor U17683 (N_17683,N_17264,N_17052);
nor U17684 (N_17684,N_17253,N_17086);
nor U17685 (N_17685,N_17247,N_17306);
xnor U17686 (N_17686,N_17295,N_17367);
and U17687 (N_17687,N_17109,N_17393);
and U17688 (N_17688,N_17293,N_17003);
and U17689 (N_17689,N_17350,N_17261);
nand U17690 (N_17690,N_17269,N_17378);
or U17691 (N_17691,N_17124,N_17088);
nor U17692 (N_17692,N_17028,N_17455);
nor U17693 (N_17693,N_17254,N_17466);
xor U17694 (N_17694,N_17275,N_17134);
xnor U17695 (N_17695,N_17397,N_17320);
nor U17696 (N_17696,N_17418,N_17321);
nor U17697 (N_17697,N_17422,N_17114);
xor U17698 (N_17698,N_17212,N_17475);
or U17699 (N_17699,N_17228,N_17389);
or U17700 (N_17700,N_17076,N_17303);
or U17701 (N_17701,N_17001,N_17387);
xor U17702 (N_17702,N_17070,N_17195);
and U17703 (N_17703,N_17202,N_17063);
xor U17704 (N_17704,N_17127,N_17209);
or U17705 (N_17705,N_17337,N_17459);
xnor U17706 (N_17706,N_17286,N_17292);
nor U17707 (N_17707,N_17488,N_17224);
and U17708 (N_17708,N_17115,N_17311);
and U17709 (N_17709,N_17060,N_17477);
and U17710 (N_17710,N_17454,N_17363);
nor U17711 (N_17711,N_17172,N_17319);
xor U17712 (N_17712,N_17497,N_17447);
and U17713 (N_17713,N_17384,N_17147);
xor U17714 (N_17714,N_17164,N_17165);
or U17715 (N_17715,N_17323,N_17190);
or U17716 (N_17716,N_17117,N_17159);
nor U17717 (N_17717,N_17120,N_17248);
xor U17718 (N_17718,N_17126,N_17179);
or U17719 (N_17719,N_17065,N_17291);
and U17720 (N_17720,N_17048,N_17130);
and U17721 (N_17721,N_17340,N_17499);
xnor U17722 (N_17722,N_17036,N_17260);
nor U17723 (N_17723,N_17071,N_17225);
nand U17724 (N_17724,N_17361,N_17138);
nor U17725 (N_17725,N_17373,N_17444);
nand U17726 (N_17726,N_17091,N_17046);
and U17727 (N_17727,N_17073,N_17119);
xnor U17728 (N_17728,N_17290,N_17478);
or U17729 (N_17729,N_17390,N_17053);
and U17730 (N_17730,N_17376,N_17336);
nand U17731 (N_17731,N_17023,N_17417);
or U17732 (N_17732,N_17196,N_17242);
nand U17733 (N_17733,N_17068,N_17054);
nand U17734 (N_17734,N_17451,N_17408);
xnor U17735 (N_17735,N_17487,N_17234);
nor U17736 (N_17736,N_17122,N_17144);
nand U17737 (N_17737,N_17460,N_17205);
or U17738 (N_17738,N_17369,N_17498);
and U17739 (N_17739,N_17452,N_17425);
and U17740 (N_17740,N_17285,N_17169);
nor U17741 (N_17741,N_17177,N_17227);
nor U17742 (N_17742,N_17161,N_17426);
nor U17743 (N_17743,N_17341,N_17221);
nand U17744 (N_17744,N_17330,N_17469);
nor U17745 (N_17745,N_17218,N_17302);
nand U17746 (N_17746,N_17325,N_17332);
nand U17747 (N_17747,N_17131,N_17359);
xor U17748 (N_17748,N_17010,N_17354);
nand U17749 (N_17749,N_17011,N_17208);
nand U17750 (N_17750,N_17155,N_17374);
or U17751 (N_17751,N_17285,N_17243);
and U17752 (N_17752,N_17148,N_17190);
xnor U17753 (N_17753,N_17245,N_17457);
and U17754 (N_17754,N_17035,N_17369);
or U17755 (N_17755,N_17100,N_17188);
nor U17756 (N_17756,N_17272,N_17161);
xor U17757 (N_17757,N_17119,N_17288);
or U17758 (N_17758,N_17108,N_17123);
nor U17759 (N_17759,N_17464,N_17425);
or U17760 (N_17760,N_17234,N_17125);
or U17761 (N_17761,N_17109,N_17474);
xnor U17762 (N_17762,N_17137,N_17141);
and U17763 (N_17763,N_17474,N_17296);
or U17764 (N_17764,N_17077,N_17317);
nor U17765 (N_17765,N_17015,N_17400);
and U17766 (N_17766,N_17354,N_17418);
nor U17767 (N_17767,N_17059,N_17056);
xnor U17768 (N_17768,N_17204,N_17189);
nand U17769 (N_17769,N_17091,N_17387);
or U17770 (N_17770,N_17095,N_17060);
nand U17771 (N_17771,N_17457,N_17297);
or U17772 (N_17772,N_17481,N_17176);
nor U17773 (N_17773,N_17121,N_17039);
nand U17774 (N_17774,N_17179,N_17425);
nand U17775 (N_17775,N_17288,N_17279);
or U17776 (N_17776,N_17160,N_17359);
and U17777 (N_17777,N_17207,N_17388);
and U17778 (N_17778,N_17075,N_17278);
and U17779 (N_17779,N_17240,N_17205);
and U17780 (N_17780,N_17287,N_17219);
xnor U17781 (N_17781,N_17436,N_17097);
nor U17782 (N_17782,N_17322,N_17108);
and U17783 (N_17783,N_17387,N_17190);
or U17784 (N_17784,N_17113,N_17239);
nor U17785 (N_17785,N_17150,N_17076);
nor U17786 (N_17786,N_17312,N_17232);
or U17787 (N_17787,N_17171,N_17060);
or U17788 (N_17788,N_17336,N_17120);
and U17789 (N_17789,N_17301,N_17430);
and U17790 (N_17790,N_17171,N_17494);
xor U17791 (N_17791,N_17407,N_17280);
nor U17792 (N_17792,N_17012,N_17117);
and U17793 (N_17793,N_17158,N_17384);
nor U17794 (N_17794,N_17098,N_17394);
xnor U17795 (N_17795,N_17404,N_17405);
nor U17796 (N_17796,N_17364,N_17067);
nand U17797 (N_17797,N_17416,N_17344);
and U17798 (N_17798,N_17075,N_17248);
nor U17799 (N_17799,N_17003,N_17000);
nor U17800 (N_17800,N_17018,N_17324);
nand U17801 (N_17801,N_17436,N_17492);
xor U17802 (N_17802,N_17082,N_17189);
or U17803 (N_17803,N_17437,N_17141);
nor U17804 (N_17804,N_17090,N_17407);
or U17805 (N_17805,N_17247,N_17310);
nor U17806 (N_17806,N_17109,N_17230);
or U17807 (N_17807,N_17292,N_17404);
xnor U17808 (N_17808,N_17140,N_17061);
nand U17809 (N_17809,N_17411,N_17317);
and U17810 (N_17810,N_17485,N_17430);
or U17811 (N_17811,N_17312,N_17023);
xnor U17812 (N_17812,N_17168,N_17460);
nor U17813 (N_17813,N_17471,N_17259);
nand U17814 (N_17814,N_17419,N_17489);
or U17815 (N_17815,N_17075,N_17273);
nor U17816 (N_17816,N_17403,N_17060);
nand U17817 (N_17817,N_17367,N_17247);
nor U17818 (N_17818,N_17019,N_17231);
and U17819 (N_17819,N_17314,N_17264);
and U17820 (N_17820,N_17143,N_17250);
xnor U17821 (N_17821,N_17056,N_17355);
and U17822 (N_17822,N_17003,N_17431);
nor U17823 (N_17823,N_17445,N_17237);
or U17824 (N_17824,N_17239,N_17042);
nor U17825 (N_17825,N_17115,N_17331);
or U17826 (N_17826,N_17224,N_17482);
or U17827 (N_17827,N_17371,N_17000);
and U17828 (N_17828,N_17249,N_17256);
or U17829 (N_17829,N_17462,N_17482);
or U17830 (N_17830,N_17098,N_17403);
and U17831 (N_17831,N_17074,N_17162);
xor U17832 (N_17832,N_17233,N_17153);
or U17833 (N_17833,N_17398,N_17387);
or U17834 (N_17834,N_17076,N_17015);
or U17835 (N_17835,N_17454,N_17271);
and U17836 (N_17836,N_17317,N_17367);
and U17837 (N_17837,N_17353,N_17270);
and U17838 (N_17838,N_17475,N_17347);
or U17839 (N_17839,N_17288,N_17325);
xnor U17840 (N_17840,N_17295,N_17147);
xnor U17841 (N_17841,N_17232,N_17362);
nor U17842 (N_17842,N_17285,N_17469);
xnor U17843 (N_17843,N_17257,N_17258);
or U17844 (N_17844,N_17347,N_17254);
xor U17845 (N_17845,N_17087,N_17061);
nor U17846 (N_17846,N_17107,N_17306);
nor U17847 (N_17847,N_17432,N_17004);
or U17848 (N_17848,N_17133,N_17391);
xor U17849 (N_17849,N_17108,N_17197);
nor U17850 (N_17850,N_17343,N_17312);
nand U17851 (N_17851,N_17011,N_17280);
xnor U17852 (N_17852,N_17269,N_17438);
or U17853 (N_17853,N_17379,N_17319);
xor U17854 (N_17854,N_17457,N_17123);
and U17855 (N_17855,N_17380,N_17348);
or U17856 (N_17856,N_17221,N_17269);
nor U17857 (N_17857,N_17009,N_17301);
and U17858 (N_17858,N_17465,N_17480);
and U17859 (N_17859,N_17433,N_17073);
and U17860 (N_17860,N_17259,N_17289);
nand U17861 (N_17861,N_17445,N_17291);
nor U17862 (N_17862,N_17365,N_17326);
xnor U17863 (N_17863,N_17010,N_17002);
or U17864 (N_17864,N_17402,N_17117);
nand U17865 (N_17865,N_17178,N_17242);
or U17866 (N_17866,N_17308,N_17086);
nor U17867 (N_17867,N_17435,N_17384);
or U17868 (N_17868,N_17347,N_17239);
nand U17869 (N_17869,N_17068,N_17237);
or U17870 (N_17870,N_17095,N_17051);
or U17871 (N_17871,N_17086,N_17374);
and U17872 (N_17872,N_17402,N_17370);
or U17873 (N_17873,N_17307,N_17075);
nor U17874 (N_17874,N_17240,N_17176);
nor U17875 (N_17875,N_17288,N_17225);
nand U17876 (N_17876,N_17164,N_17349);
nand U17877 (N_17877,N_17292,N_17310);
xor U17878 (N_17878,N_17419,N_17037);
or U17879 (N_17879,N_17195,N_17474);
nor U17880 (N_17880,N_17421,N_17310);
xor U17881 (N_17881,N_17059,N_17209);
and U17882 (N_17882,N_17493,N_17050);
nand U17883 (N_17883,N_17083,N_17064);
nor U17884 (N_17884,N_17258,N_17372);
xnor U17885 (N_17885,N_17276,N_17148);
xnor U17886 (N_17886,N_17100,N_17294);
and U17887 (N_17887,N_17211,N_17136);
nor U17888 (N_17888,N_17370,N_17178);
or U17889 (N_17889,N_17269,N_17076);
nand U17890 (N_17890,N_17388,N_17468);
xor U17891 (N_17891,N_17195,N_17265);
or U17892 (N_17892,N_17171,N_17217);
xnor U17893 (N_17893,N_17189,N_17446);
or U17894 (N_17894,N_17149,N_17123);
xor U17895 (N_17895,N_17290,N_17264);
or U17896 (N_17896,N_17244,N_17030);
nand U17897 (N_17897,N_17169,N_17211);
and U17898 (N_17898,N_17054,N_17234);
and U17899 (N_17899,N_17029,N_17193);
and U17900 (N_17900,N_17170,N_17376);
or U17901 (N_17901,N_17155,N_17299);
nor U17902 (N_17902,N_17236,N_17391);
or U17903 (N_17903,N_17403,N_17239);
nor U17904 (N_17904,N_17104,N_17425);
or U17905 (N_17905,N_17290,N_17100);
xor U17906 (N_17906,N_17007,N_17031);
nor U17907 (N_17907,N_17069,N_17109);
nand U17908 (N_17908,N_17328,N_17087);
nand U17909 (N_17909,N_17371,N_17109);
or U17910 (N_17910,N_17236,N_17048);
nand U17911 (N_17911,N_17158,N_17014);
nor U17912 (N_17912,N_17412,N_17373);
nor U17913 (N_17913,N_17311,N_17167);
and U17914 (N_17914,N_17025,N_17146);
nand U17915 (N_17915,N_17009,N_17251);
and U17916 (N_17916,N_17308,N_17077);
xor U17917 (N_17917,N_17184,N_17102);
nand U17918 (N_17918,N_17097,N_17403);
and U17919 (N_17919,N_17351,N_17423);
nor U17920 (N_17920,N_17032,N_17317);
nor U17921 (N_17921,N_17178,N_17268);
xor U17922 (N_17922,N_17464,N_17097);
and U17923 (N_17923,N_17364,N_17037);
and U17924 (N_17924,N_17151,N_17333);
and U17925 (N_17925,N_17442,N_17143);
nor U17926 (N_17926,N_17426,N_17402);
nand U17927 (N_17927,N_17411,N_17338);
nand U17928 (N_17928,N_17258,N_17111);
or U17929 (N_17929,N_17288,N_17188);
and U17930 (N_17930,N_17132,N_17035);
and U17931 (N_17931,N_17433,N_17375);
nand U17932 (N_17932,N_17147,N_17441);
xnor U17933 (N_17933,N_17042,N_17379);
nand U17934 (N_17934,N_17303,N_17160);
nand U17935 (N_17935,N_17241,N_17120);
xnor U17936 (N_17936,N_17077,N_17141);
nand U17937 (N_17937,N_17372,N_17025);
or U17938 (N_17938,N_17300,N_17478);
nor U17939 (N_17939,N_17343,N_17168);
and U17940 (N_17940,N_17003,N_17401);
and U17941 (N_17941,N_17326,N_17247);
xnor U17942 (N_17942,N_17264,N_17468);
or U17943 (N_17943,N_17168,N_17341);
nor U17944 (N_17944,N_17116,N_17354);
nor U17945 (N_17945,N_17039,N_17186);
and U17946 (N_17946,N_17268,N_17278);
or U17947 (N_17947,N_17297,N_17480);
nor U17948 (N_17948,N_17395,N_17084);
nand U17949 (N_17949,N_17396,N_17172);
or U17950 (N_17950,N_17438,N_17337);
and U17951 (N_17951,N_17186,N_17076);
and U17952 (N_17952,N_17136,N_17032);
nand U17953 (N_17953,N_17317,N_17283);
xnor U17954 (N_17954,N_17245,N_17039);
xor U17955 (N_17955,N_17114,N_17071);
nor U17956 (N_17956,N_17190,N_17171);
xor U17957 (N_17957,N_17406,N_17437);
or U17958 (N_17958,N_17491,N_17448);
xnor U17959 (N_17959,N_17400,N_17082);
xor U17960 (N_17960,N_17229,N_17434);
nor U17961 (N_17961,N_17392,N_17313);
nand U17962 (N_17962,N_17131,N_17171);
nand U17963 (N_17963,N_17273,N_17348);
nand U17964 (N_17964,N_17026,N_17311);
or U17965 (N_17965,N_17248,N_17119);
or U17966 (N_17966,N_17348,N_17250);
or U17967 (N_17967,N_17232,N_17343);
and U17968 (N_17968,N_17453,N_17062);
or U17969 (N_17969,N_17295,N_17085);
xor U17970 (N_17970,N_17204,N_17456);
nor U17971 (N_17971,N_17071,N_17302);
and U17972 (N_17972,N_17365,N_17396);
nand U17973 (N_17973,N_17287,N_17224);
xnor U17974 (N_17974,N_17273,N_17419);
xor U17975 (N_17975,N_17226,N_17154);
nand U17976 (N_17976,N_17359,N_17050);
xor U17977 (N_17977,N_17106,N_17242);
nor U17978 (N_17978,N_17385,N_17445);
nand U17979 (N_17979,N_17316,N_17255);
nor U17980 (N_17980,N_17398,N_17353);
and U17981 (N_17981,N_17060,N_17011);
and U17982 (N_17982,N_17343,N_17154);
or U17983 (N_17983,N_17085,N_17384);
or U17984 (N_17984,N_17299,N_17157);
nor U17985 (N_17985,N_17487,N_17316);
or U17986 (N_17986,N_17288,N_17075);
and U17987 (N_17987,N_17331,N_17489);
or U17988 (N_17988,N_17351,N_17371);
nand U17989 (N_17989,N_17276,N_17395);
xnor U17990 (N_17990,N_17185,N_17007);
nand U17991 (N_17991,N_17284,N_17408);
or U17992 (N_17992,N_17067,N_17429);
xnor U17993 (N_17993,N_17245,N_17067);
and U17994 (N_17994,N_17159,N_17076);
and U17995 (N_17995,N_17064,N_17282);
xor U17996 (N_17996,N_17415,N_17083);
or U17997 (N_17997,N_17059,N_17472);
xor U17998 (N_17998,N_17220,N_17168);
xnor U17999 (N_17999,N_17444,N_17217);
xnor U18000 (N_18000,N_17692,N_17500);
xor U18001 (N_18001,N_17633,N_17975);
xor U18002 (N_18002,N_17932,N_17835);
and U18003 (N_18003,N_17760,N_17985);
or U18004 (N_18004,N_17501,N_17657);
nor U18005 (N_18005,N_17684,N_17524);
xor U18006 (N_18006,N_17590,N_17928);
nand U18007 (N_18007,N_17822,N_17648);
xor U18008 (N_18008,N_17614,N_17768);
and U18009 (N_18009,N_17634,N_17509);
nor U18010 (N_18010,N_17960,N_17737);
and U18011 (N_18011,N_17586,N_17974);
or U18012 (N_18012,N_17749,N_17560);
or U18013 (N_18013,N_17956,N_17693);
and U18014 (N_18014,N_17718,N_17802);
nand U18015 (N_18015,N_17886,N_17854);
nand U18016 (N_18016,N_17784,N_17631);
and U18017 (N_18017,N_17627,N_17608);
or U18018 (N_18018,N_17907,N_17548);
or U18019 (N_18019,N_17970,N_17998);
nand U18020 (N_18020,N_17504,N_17740);
or U18021 (N_18021,N_17581,N_17545);
xor U18022 (N_18022,N_17644,N_17685);
xnor U18023 (N_18023,N_17893,N_17966);
or U18024 (N_18024,N_17994,N_17541);
and U18025 (N_18025,N_17579,N_17773);
or U18026 (N_18026,N_17521,N_17971);
nand U18027 (N_18027,N_17831,N_17688);
and U18028 (N_18028,N_17779,N_17803);
and U18029 (N_18029,N_17572,N_17729);
nor U18030 (N_18030,N_17777,N_17515);
nor U18031 (N_18031,N_17630,N_17576);
xnor U18032 (N_18032,N_17559,N_17787);
nand U18033 (N_18033,N_17896,N_17655);
xnor U18034 (N_18034,N_17722,N_17591);
or U18035 (N_18035,N_17786,N_17708);
and U18036 (N_18036,N_17616,N_17789);
or U18037 (N_18037,N_17588,N_17759);
and U18038 (N_18038,N_17810,N_17875);
xor U18039 (N_18039,N_17554,N_17561);
xnor U18040 (N_18040,N_17715,N_17719);
xnor U18041 (N_18041,N_17671,N_17938);
nor U18042 (N_18042,N_17701,N_17919);
nand U18043 (N_18043,N_17700,N_17852);
xnor U18044 (N_18044,N_17632,N_17703);
and U18045 (N_18045,N_17678,N_17646);
xnor U18046 (N_18046,N_17776,N_17796);
xor U18047 (N_18047,N_17834,N_17964);
and U18048 (N_18048,N_17664,N_17574);
or U18049 (N_18049,N_17731,N_17566);
xnor U18050 (N_18050,N_17819,N_17676);
xnor U18051 (N_18051,N_17531,N_17903);
and U18052 (N_18052,N_17544,N_17795);
xnor U18053 (N_18053,N_17871,N_17766);
nor U18054 (N_18054,N_17750,N_17533);
xnor U18055 (N_18055,N_17889,N_17818);
nor U18056 (N_18056,N_17681,N_17954);
and U18057 (N_18057,N_17969,N_17730);
nor U18058 (N_18058,N_17667,N_17883);
or U18059 (N_18059,N_17965,N_17535);
nand U18060 (N_18060,N_17930,N_17727);
xnor U18061 (N_18061,N_17536,N_17872);
nor U18062 (N_18062,N_17649,N_17526);
and U18063 (N_18063,N_17611,N_17884);
or U18064 (N_18064,N_17902,N_17552);
nand U18065 (N_18065,N_17816,N_17546);
xnor U18066 (N_18066,N_17650,N_17885);
or U18067 (N_18067,N_17949,N_17702);
and U18068 (N_18068,N_17943,N_17656);
or U18069 (N_18069,N_17625,N_17859);
or U18070 (N_18070,N_17673,N_17542);
and U18071 (N_18071,N_17944,N_17543);
and U18072 (N_18072,N_17506,N_17597);
or U18073 (N_18073,N_17939,N_17940);
nand U18074 (N_18074,N_17799,N_17774);
nor U18075 (N_18075,N_17840,N_17647);
xnor U18076 (N_18076,N_17739,N_17563);
xnor U18077 (N_18077,N_17710,N_17629);
nand U18078 (N_18078,N_17758,N_17780);
nand U18079 (N_18079,N_17841,N_17848);
or U18080 (N_18080,N_17920,N_17751);
nand U18081 (N_18081,N_17997,N_17661);
nand U18082 (N_18082,N_17658,N_17988);
nor U18083 (N_18083,N_17717,N_17516);
or U18084 (N_18084,N_17508,N_17880);
xor U18085 (N_18085,N_17585,N_17674);
and U18086 (N_18086,N_17899,N_17596);
nor U18087 (N_18087,N_17771,N_17520);
nor U18088 (N_18088,N_17558,N_17926);
and U18089 (N_18089,N_17617,N_17892);
or U18090 (N_18090,N_17951,N_17677);
and U18091 (N_18091,N_17514,N_17555);
xnor U18092 (N_18092,N_17947,N_17817);
nand U18093 (N_18093,N_17811,N_17675);
nor U18094 (N_18094,N_17663,N_17993);
xnor U18095 (N_18095,N_17618,N_17550);
nand U18096 (N_18096,N_17679,N_17946);
nand U18097 (N_18097,N_17842,N_17711);
xnor U18098 (N_18098,N_17979,N_17936);
nor U18099 (N_18099,N_17553,N_17910);
xor U18100 (N_18100,N_17977,N_17837);
and U18101 (N_18101,N_17788,N_17670);
xnor U18102 (N_18102,N_17532,N_17522);
and U18103 (N_18103,N_17824,N_17921);
and U18104 (N_18104,N_17748,N_17991);
nor U18105 (N_18105,N_17900,N_17615);
or U18106 (N_18106,N_17623,N_17726);
and U18107 (N_18107,N_17704,N_17912);
nand U18108 (N_18108,N_17955,N_17732);
xnor U18109 (N_18109,N_17849,N_17976);
xnor U18110 (N_18110,N_17598,N_17530);
or U18111 (N_18111,N_17851,N_17838);
xnor U18112 (N_18112,N_17933,N_17924);
and U18113 (N_18113,N_17950,N_17980);
and U18114 (N_18114,N_17793,N_17782);
or U18115 (N_18115,N_17867,N_17698);
nand U18116 (N_18116,N_17745,N_17741);
nand U18117 (N_18117,N_17728,N_17682);
xnor U18118 (N_18118,N_17525,N_17645);
nand U18119 (N_18119,N_17705,N_17984);
nor U18120 (N_18120,N_17813,N_17791);
and U18121 (N_18121,N_17747,N_17589);
xor U18122 (N_18122,N_17833,N_17913);
or U18123 (N_18123,N_17669,N_17894);
nor U18124 (N_18124,N_17662,N_17820);
xor U18125 (N_18125,N_17914,N_17952);
xnor U18126 (N_18126,N_17551,N_17918);
nor U18127 (N_18127,N_17781,N_17957);
or U18128 (N_18128,N_17942,N_17503);
xor U18129 (N_18129,N_17861,N_17735);
and U18130 (N_18130,N_17996,N_17850);
or U18131 (N_18131,N_17755,N_17839);
or U18132 (N_18132,N_17635,N_17564);
nor U18133 (N_18133,N_17517,N_17593);
xor U18134 (N_18134,N_17978,N_17606);
nor U18135 (N_18135,N_17602,N_17990);
or U18136 (N_18136,N_17601,N_17734);
nor U18137 (N_18137,N_17808,N_17761);
nand U18138 (N_18138,N_17573,N_17651);
and U18139 (N_18139,N_17866,N_17832);
nor U18140 (N_18140,N_17511,N_17643);
or U18141 (N_18141,N_17959,N_17805);
and U18142 (N_18142,N_17724,N_17580);
nor U18143 (N_18143,N_17931,N_17668);
and U18144 (N_18144,N_17595,N_17605);
xor U18145 (N_18145,N_17887,N_17807);
nor U18146 (N_18146,N_17821,N_17778);
or U18147 (N_18147,N_17857,N_17765);
nor U18148 (N_18148,N_17916,N_17764);
or U18149 (N_18149,N_17540,N_17638);
and U18150 (N_18150,N_17736,N_17733);
nand U18151 (N_18151,N_17981,N_17923);
and U18152 (N_18152,N_17637,N_17763);
and U18153 (N_18153,N_17707,N_17538);
nand U18154 (N_18154,N_17876,N_17502);
and U18155 (N_18155,N_17527,N_17666);
nor U18156 (N_18156,N_17529,N_17699);
or U18157 (N_18157,N_17641,N_17587);
or U18158 (N_18158,N_17672,N_17697);
nor U18159 (N_18159,N_17706,N_17856);
or U18160 (N_18160,N_17995,N_17756);
or U18161 (N_18161,N_17583,N_17694);
nor U18162 (N_18162,N_17860,N_17642);
nor U18163 (N_18163,N_17915,N_17891);
or U18164 (N_18164,N_17754,N_17604);
nand U18165 (N_18165,N_17571,N_17743);
xnor U18166 (N_18166,N_17652,N_17770);
nand U18167 (N_18167,N_17953,N_17738);
xnor U18168 (N_18168,N_17830,N_17895);
or U18169 (N_18169,N_17603,N_17716);
xnor U18170 (N_18170,N_17610,N_17826);
or U18171 (N_18171,N_17686,N_17567);
or U18172 (N_18172,N_17855,N_17695);
xnor U18173 (N_18173,N_17654,N_17945);
nand U18174 (N_18174,N_17846,N_17626);
nor U18175 (N_18175,N_17844,N_17687);
nor U18176 (N_18176,N_17523,N_17827);
and U18177 (N_18177,N_17723,N_17815);
nor U18178 (N_18178,N_17636,N_17941);
or U18179 (N_18179,N_17639,N_17612);
nand U18180 (N_18180,N_17853,N_17792);
xnor U18181 (N_18181,N_17987,N_17691);
nand U18182 (N_18182,N_17547,N_17518);
or U18183 (N_18183,N_17801,N_17513);
nor U18184 (N_18184,N_17878,N_17609);
and U18185 (N_18185,N_17983,N_17982);
xor U18186 (N_18186,N_17881,N_17869);
and U18187 (N_18187,N_17565,N_17539);
and U18188 (N_18188,N_17569,N_17898);
nand U18189 (N_18189,N_17613,N_17690);
xnor U18190 (N_18190,N_17742,N_17962);
nor U18191 (N_18191,N_17804,N_17549);
nor U18192 (N_18192,N_17972,N_17534);
and U18193 (N_18193,N_17556,N_17659);
nor U18194 (N_18194,N_17794,N_17689);
and U18195 (N_18195,N_17825,N_17653);
xnor U18196 (N_18196,N_17911,N_17906);
xnor U18197 (N_18197,N_17709,N_17680);
nand U18198 (N_18198,N_17870,N_17973);
nor U18199 (N_18199,N_17783,N_17696);
nand U18200 (N_18200,N_17762,N_17829);
and U18201 (N_18201,N_17628,N_17927);
nor U18202 (N_18202,N_17901,N_17683);
and U18203 (N_18203,N_17963,N_17917);
or U18204 (N_18204,N_17578,N_17519);
nand U18205 (N_18205,N_17570,N_17934);
nand U18206 (N_18206,N_17619,N_17752);
and U18207 (N_18207,N_17909,N_17935);
nor U18208 (N_18208,N_17845,N_17864);
nand U18209 (N_18209,N_17961,N_17512);
nor U18210 (N_18210,N_17828,N_17660);
or U18211 (N_18211,N_17753,N_17790);
nand U18212 (N_18212,N_17713,N_17863);
or U18213 (N_18213,N_17897,N_17562);
and U18214 (N_18214,N_17868,N_17757);
or U18215 (N_18215,N_17721,N_17624);
xor U18216 (N_18216,N_17621,N_17775);
xor U18217 (N_18217,N_17537,N_17858);
xnor U18218 (N_18218,N_17592,N_17890);
xor U18219 (N_18219,N_17847,N_17725);
nor U18220 (N_18220,N_17712,N_17797);
or U18221 (N_18221,N_17785,N_17568);
and U18222 (N_18222,N_17772,N_17843);
or U18223 (N_18223,N_17986,N_17809);
and U18224 (N_18224,N_17879,N_17967);
and U18225 (N_18225,N_17607,N_17948);
nor U18226 (N_18226,N_17746,N_17575);
nand U18227 (N_18227,N_17800,N_17812);
and U18228 (N_18228,N_17992,N_17744);
xor U18229 (N_18229,N_17882,N_17577);
nand U18230 (N_18230,N_17584,N_17767);
and U18231 (N_18231,N_17622,N_17925);
and U18232 (N_18232,N_17877,N_17888);
xnor U18233 (N_18233,N_17999,N_17873);
xor U18234 (N_18234,N_17665,N_17929);
or U18235 (N_18235,N_17557,N_17798);
nand U18236 (N_18236,N_17836,N_17505);
nand U18237 (N_18237,N_17806,N_17989);
nand U18238 (N_18238,N_17908,N_17594);
or U18239 (N_18239,N_17582,N_17528);
nand U18240 (N_18240,N_17814,N_17968);
nand U18241 (N_18241,N_17720,N_17904);
nor U18242 (N_18242,N_17922,N_17640);
and U18243 (N_18243,N_17874,N_17937);
nand U18244 (N_18244,N_17958,N_17823);
or U18245 (N_18245,N_17865,N_17620);
nand U18246 (N_18246,N_17600,N_17510);
nor U18247 (N_18247,N_17862,N_17905);
and U18248 (N_18248,N_17769,N_17507);
nand U18249 (N_18249,N_17714,N_17599);
and U18250 (N_18250,N_17993,N_17872);
nor U18251 (N_18251,N_17959,N_17629);
xor U18252 (N_18252,N_17664,N_17610);
xnor U18253 (N_18253,N_17604,N_17593);
and U18254 (N_18254,N_17643,N_17622);
xor U18255 (N_18255,N_17911,N_17690);
nand U18256 (N_18256,N_17502,N_17855);
xor U18257 (N_18257,N_17652,N_17590);
xor U18258 (N_18258,N_17658,N_17946);
xor U18259 (N_18259,N_17595,N_17915);
nor U18260 (N_18260,N_17710,N_17914);
nor U18261 (N_18261,N_17988,N_17509);
and U18262 (N_18262,N_17850,N_17902);
nand U18263 (N_18263,N_17623,N_17664);
and U18264 (N_18264,N_17895,N_17778);
or U18265 (N_18265,N_17581,N_17784);
and U18266 (N_18266,N_17517,N_17860);
or U18267 (N_18267,N_17576,N_17647);
xnor U18268 (N_18268,N_17595,N_17807);
xnor U18269 (N_18269,N_17615,N_17709);
nand U18270 (N_18270,N_17949,N_17617);
and U18271 (N_18271,N_17966,N_17933);
nand U18272 (N_18272,N_17554,N_17869);
xor U18273 (N_18273,N_17677,N_17617);
xor U18274 (N_18274,N_17526,N_17921);
or U18275 (N_18275,N_17514,N_17936);
nand U18276 (N_18276,N_17891,N_17910);
nor U18277 (N_18277,N_17857,N_17752);
xnor U18278 (N_18278,N_17935,N_17824);
nand U18279 (N_18279,N_17577,N_17556);
or U18280 (N_18280,N_17680,N_17784);
nor U18281 (N_18281,N_17608,N_17798);
nor U18282 (N_18282,N_17667,N_17998);
nor U18283 (N_18283,N_17894,N_17691);
xor U18284 (N_18284,N_17968,N_17791);
nor U18285 (N_18285,N_17642,N_17826);
xor U18286 (N_18286,N_17545,N_17528);
or U18287 (N_18287,N_17984,N_17757);
nor U18288 (N_18288,N_17625,N_17708);
and U18289 (N_18289,N_17918,N_17720);
xnor U18290 (N_18290,N_17826,N_17950);
nand U18291 (N_18291,N_17672,N_17623);
or U18292 (N_18292,N_17785,N_17640);
and U18293 (N_18293,N_17952,N_17751);
nand U18294 (N_18294,N_17850,N_17539);
and U18295 (N_18295,N_17647,N_17939);
and U18296 (N_18296,N_17594,N_17802);
and U18297 (N_18297,N_17850,N_17657);
nor U18298 (N_18298,N_17942,N_17640);
or U18299 (N_18299,N_17916,N_17714);
and U18300 (N_18300,N_17830,N_17776);
nor U18301 (N_18301,N_17764,N_17729);
nand U18302 (N_18302,N_17701,N_17841);
nor U18303 (N_18303,N_17573,N_17921);
xnor U18304 (N_18304,N_17611,N_17599);
or U18305 (N_18305,N_17645,N_17963);
nor U18306 (N_18306,N_17601,N_17674);
and U18307 (N_18307,N_17912,N_17723);
xnor U18308 (N_18308,N_17710,N_17559);
nand U18309 (N_18309,N_17629,N_17936);
or U18310 (N_18310,N_17689,N_17638);
and U18311 (N_18311,N_17767,N_17646);
nor U18312 (N_18312,N_17628,N_17892);
or U18313 (N_18313,N_17856,N_17757);
nand U18314 (N_18314,N_17615,N_17986);
nor U18315 (N_18315,N_17852,N_17611);
nor U18316 (N_18316,N_17983,N_17675);
or U18317 (N_18317,N_17837,N_17538);
nor U18318 (N_18318,N_17596,N_17843);
nor U18319 (N_18319,N_17778,N_17573);
xor U18320 (N_18320,N_17829,N_17880);
and U18321 (N_18321,N_17643,N_17768);
nor U18322 (N_18322,N_17523,N_17533);
or U18323 (N_18323,N_17845,N_17801);
or U18324 (N_18324,N_17788,N_17527);
or U18325 (N_18325,N_17869,N_17991);
and U18326 (N_18326,N_17583,N_17712);
and U18327 (N_18327,N_17685,N_17512);
and U18328 (N_18328,N_17801,N_17762);
nor U18329 (N_18329,N_17690,N_17771);
and U18330 (N_18330,N_17541,N_17529);
xor U18331 (N_18331,N_17902,N_17870);
and U18332 (N_18332,N_17903,N_17644);
or U18333 (N_18333,N_17503,N_17991);
nand U18334 (N_18334,N_17973,N_17504);
nor U18335 (N_18335,N_17854,N_17902);
or U18336 (N_18336,N_17897,N_17529);
nor U18337 (N_18337,N_17974,N_17658);
nor U18338 (N_18338,N_17748,N_17971);
and U18339 (N_18339,N_17514,N_17774);
nor U18340 (N_18340,N_17678,N_17673);
and U18341 (N_18341,N_17677,N_17620);
nor U18342 (N_18342,N_17869,N_17781);
nand U18343 (N_18343,N_17748,N_17936);
nand U18344 (N_18344,N_17801,N_17593);
nand U18345 (N_18345,N_17839,N_17624);
nand U18346 (N_18346,N_17870,N_17990);
or U18347 (N_18347,N_17984,N_17889);
nor U18348 (N_18348,N_17783,N_17805);
xnor U18349 (N_18349,N_17913,N_17515);
nor U18350 (N_18350,N_17650,N_17609);
nor U18351 (N_18351,N_17654,N_17992);
and U18352 (N_18352,N_17927,N_17782);
nor U18353 (N_18353,N_17733,N_17881);
or U18354 (N_18354,N_17879,N_17728);
nand U18355 (N_18355,N_17911,N_17795);
and U18356 (N_18356,N_17577,N_17646);
or U18357 (N_18357,N_17911,N_17663);
or U18358 (N_18358,N_17573,N_17872);
xor U18359 (N_18359,N_17810,N_17659);
nor U18360 (N_18360,N_17757,N_17677);
nand U18361 (N_18361,N_17824,N_17583);
or U18362 (N_18362,N_17825,N_17665);
and U18363 (N_18363,N_17991,N_17770);
nor U18364 (N_18364,N_17747,N_17845);
and U18365 (N_18365,N_17815,N_17984);
or U18366 (N_18366,N_17809,N_17877);
nor U18367 (N_18367,N_17738,N_17992);
or U18368 (N_18368,N_17729,N_17510);
and U18369 (N_18369,N_17638,N_17952);
nor U18370 (N_18370,N_17864,N_17978);
or U18371 (N_18371,N_17981,N_17543);
and U18372 (N_18372,N_17900,N_17730);
and U18373 (N_18373,N_17713,N_17644);
or U18374 (N_18374,N_17757,N_17997);
nor U18375 (N_18375,N_17911,N_17685);
and U18376 (N_18376,N_17857,N_17736);
or U18377 (N_18377,N_17635,N_17814);
nor U18378 (N_18378,N_17829,N_17870);
and U18379 (N_18379,N_17750,N_17818);
and U18380 (N_18380,N_17877,N_17517);
xnor U18381 (N_18381,N_17922,N_17524);
and U18382 (N_18382,N_17894,N_17557);
nor U18383 (N_18383,N_17636,N_17990);
nand U18384 (N_18384,N_17541,N_17937);
and U18385 (N_18385,N_17661,N_17560);
nor U18386 (N_18386,N_17913,N_17571);
or U18387 (N_18387,N_17931,N_17633);
nand U18388 (N_18388,N_17832,N_17994);
xor U18389 (N_18389,N_17589,N_17500);
nor U18390 (N_18390,N_17569,N_17888);
and U18391 (N_18391,N_17845,N_17632);
xor U18392 (N_18392,N_17954,N_17709);
nand U18393 (N_18393,N_17865,N_17933);
nand U18394 (N_18394,N_17683,N_17594);
and U18395 (N_18395,N_17675,N_17697);
nor U18396 (N_18396,N_17508,N_17592);
and U18397 (N_18397,N_17999,N_17756);
xnor U18398 (N_18398,N_17686,N_17907);
and U18399 (N_18399,N_17951,N_17878);
xor U18400 (N_18400,N_17732,N_17547);
nand U18401 (N_18401,N_17829,N_17770);
nor U18402 (N_18402,N_17953,N_17580);
nand U18403 (N_18403,N_17643,N_17537);
and U18404 (N_18404,N_17955,N_17733);
xor U18405 (N_18405,N_17903,N_17744);
or U18406 (N_18406,N_17538,N_17527);
nor U18407 (N_18407,N_17733,N_17796);
and U18408 (N_18408,N_17588,N_17981);
xnor U18409 (N_18409,N_17539,N_17872);
or U18410 (N_18410,N_17810,N_17692);
and U18411 (N_18411,N_17843,N_17783);
xor U18412 (N_18412,N_17685,N_17923);
or U18413 (N_18413,N_17975,N_17520);
or U18414 (N_18414,N_17691,N_17709);
nor U18415 (N_18415,N_17629,N_17620);
or U18416 (N_18416,N_17961,N_17995);
nand U18417 (N_18417,N_17992,N_17529);
nor U18418 (N_18418,N_17925,N_17975);
nor U18419 (N_18419,N_17524,N_17845);
xor U18420 (N_18420,N_17790,N_17988);
nand U18421 (N_18421,N_17680,N_17662);
and U18422 (N_18422,N_17586,N_17845);
xor U18423 (N_18423,N_17963,N_17511);
and U18424 (N_18424,N_17547,N_17737);
xnor U18425 (N_18425,N_17832,N_17541);
nand U18426 (N_18426,N_17505,N_17709);
or U18427 (N_18427,N_17638,N_17561);
xor U18428 (N_18428,N_17842,N_17577);
xor U18429 (N_18429,N_17726,N_17752);
xor U18430 (N_18430,N_17857,N_17864);
xor U18431 (N_18431,N_17831,N_17651);
xor U18432 (N_18432,N_17984,N_17502);
nand U18433 (N_18433,N_17706,N_17739);
or U18434 (N_18434,N_17714,N_17612);
nand U18435 (N_18435,N_17524,N_17728);
nand U18436 (N_18436,N_17853,N_17688);
nand U18437 (N_18437,N_17732,N_17696);
nor U18438 (N_18438,N_17928,N_17723);
nor U18439 (N_18439,N_17727,N_17544);
and U18440 (N_18440,N_17506,N_17559);
nor U18441 (N_18441,N_17695,N_17721);
and U18442 (N_18442,N_17743,N_17971);
and U18443 (N_18443,N_17593,N_17759);
nand U18444 (N_18444,N_17627,N_17591);
and U18445 (N_18445,N_17724,N_17821);
or U18446 (N_18446,N_17965,N_17979);
xor U18447 (N_18447,N_17839,N_17709);
or U18448 (N_18448,N_17850,N_17707);
nor U18449 (N_18449,N_17568,N_17968);
and U18450 (N_18450,N_17627,N_17740);
or U18451 (N_18451,N_17555,N_17813);
nor U18452 (N_18452,N_17937,N_17540);
nand U18453 (N_18453,N_17619,N_17938);
nor U18454 (N_18454,N_17767,N_17805);
xor U18455 (N_18455,N_17674,N_17664);
and U18456 (N_18456,N_17879,N_17625);
nand U18457 (N_18457,N_17638,N_17852);
and U18458 (N_18458,N_17609,N_17818);
and U18459 (N_18459,N_17571,N_17935);
xnor U18460 (N_18460,N_17674,N_17955);
xnor U18461 (N_18461,N_17532,N_17842);
and U18462 (N_18462,N_17554,N_17716);
nor U18463 (N_18463,N_17638,N_17570);
and U18464 (N_18464,N_17754,N_17662);
nand U18465 (N_18465,N_17967,N_17849);
nor U18466 (N_18466,N_17857,N_17663);
and U18467 (N_18467,N_17919,N_17931);
xor U18468 (N_18468,N_17638,N_17879);
xnor U18469 (N_18469,N_17883,N_17559);
or U18470 (N_18470,N_17673,N_17593);
nand U18471 (N_18471,N_17749,N_17854);
xor U18472 (N_18472,N_17635,N_17827);
and U18473 (N_18473,N_17866,N_17789);
nor U18474 (N_18474,N_17860,N_17976);
and U18475 (N_18475,N_17601,N_17745);
nor U18476 (N_18476,N_17806,N_17860);
or U18477 (N_18477,N_17629,N_17542);
xor U18478 (N_18478,N_17911,N_17669);
and U18479 (N_18479,N_17769,N_17723);
nand U18480 (N_18480,N_17976,N_17728);
nor U18481 (N_18481,N_17972,N_17557);
or U18482 (N_18482,N_17822,N_17984);
or U18483 (N_18483,N_17978,N_17905);
and U18484 (N_18484,N_17913,N_17953);
nand U18485 (N_18485,N_17619,N_17921);
xor U18486 (N_18486,N_17716,N_17669);
nor U18487 (N_18487,N_17583,N_17632);
nand U18488 (N_18488,N_17529,N_17510);
and U18489 (N_18489,N_17690,N_17580);
and U18490 (N_18490,N_17883,N_17513);
and U18491 (N_18491,N_17752,N_17808);
and U18492 (N_18492,N_17681,N_17594);
nor U18493 (N_18493,N_17507,N_17566);
nor U18494 (N_18494,N_17952,N_17728);
nor U18495 (N_18495,N_17842,N_17913);
nor U18496 (N_18496,N_17771,N_17816);
xor U18497 (N_18497,N_17731,N_17621);
and U18498 (N_18498,N_17992,N_17705);
or U18499 (N_18499,N_17510,N_17909);
nor U18500 (N_18500,N_18078,N_18070);
or U18501 (N_18501,N_18200,N_18216);
and U18502 (N_18502,N_18479,N_18049);
nand U18503 (N_18503,N_18444,N_18489);
or U18504 (N_18504,N_18313,N_18298);
nor U18505 (N_18505,N_18483,N_18055);
or U18506 (N_18506,N_18320,N_18353);
and U18507 (N_18507,N_18182,N_18114);
xor U18508 (N_18508,N_18415,N_18021);
and U18509 (N_18509,N_18001,N_18317);
and U18510 (N_18510,N_18029,N_18421);
and U18511 (N_18511,N_18426,N_18172);
nor U18512 (N_18512,N_18458,N_18199);
nor U18513 (N_18513,N_18097,N_18263);
and U18514 (N_18514,N_18052,N_18328);
nor U18515 (N_18515,N_18314,N_18079);
and U18516 (N_18516,N_18424,N_18252);
nor U18517 (N_18517,N_18311,N_18043);
or U18518 (N_18518,N_18019,N_18150);
xnor U18519 (N_18519,N_18187,N_18084);
nor U18520 (N_18520,N_18454,N_18253);
nand U18521 (N_18521,N_18026,N_18155);
nand U18522 (N_18522,N_18148,N_18181);
nor U18523 (N_18523,N_18041,N_18406);
and U18524 (N_18524,N_18160,N_18117);
xor U18525 (N_18525,N_18345,N_18350);
and U18526 (N_18526,N_18237,N_18467);
nand U18527 (N_18527,N_18214,N_18105);
or U18528 (N_18528,N_18198,N_18032);
nor U18529 (N_18529,N_18095,N_18057);
and U18530 (N_18530,N_18101,N_18228);
and U18531 (N_18531,N_18207,N_18254);
nor U18532 (N_18532,N_18081,N_18390);
or U18533 (N_18533,N_18433,N_18071);
nor U18534 (N_18534,N_18290,N_18280);
and U18535 (N_18535,N_18235,N_18189);
and U18536 (N_18536,N_18028,N_18186);
nor U18537 (N_18537,N_18144,N_18436);
nor U18538 (N_18538,N_18146,N_18289);
xnor U18539 (N_18539,N_18062,N_18086);
or U18540 (N_18540,N_18219,N_18131);
nor U18541 (N_18541,N_18268,N_18245);
and U18542 (N_18542,N_18309,N_18145);
nor U18543 (N_18543,N_18104,N_18173);
nand U18544 (N_18544,N_18225,N_18283);
or U18545 (N_18545,N_18073,N_18069);
nor U18546 (N_18546,N_18325,N_18492);
or U18547 (N_18547,N_18474,N_18377);
xor U18548 (N_18548,N_18499,N_18323);
or U18549 (N_18549,N_18293,N_18119);
and U18550 (N_18550,N_18396,N_18184);
nor U18551 (N_18551,N_18464,N_18372);
xnor U18552 (N_18552,N_18036,N_18016);
or U18553 (N_18553,N_18209,N_18411);
xor U18554 (N_18554,N_18395,N_18151);
nor U18555 (N_18555,N_18429,N_18135);
and U18556 (N_18556,N_18238,N_18080);
or U18557 (N_18557,N_18083,N_18142);
nand U18558 (N_18558,N_18304,N_18420);
nor U18559 (N_18559,N_18352,N_18213);
and U18560 (N_18560,N_18059,N_18451);
xor U18561 (N_18561,N_18491,N_18175);
or U18562 (N_18562,N_18141,N_18301);
or U18563 (N_18563,N_18413,N_18099);
nand U18564 (N_18564,N_18264,N_18365);
or U18565 (N_18565,N_18360,N_18493);
xor U18566 (N_18566,N_18153,N_18110);
nand U18567 (N_18567,N_18262,N_18013);
xnor U18568 (N_18568,N_18340,N_18256);
nand U18569 (N_18569,N_18497,N_18361);
or U18570 (N_18570,N_18414,N_18337);
nor U18571 (N_18571,N_18241,N_18358);
or U18572 (N_18572,N_18408,N_18488);
xnor U18573 (N_18573,N_18351,N_18407);
nor U18574 (N_18574,N_18039,N_18346);
and U18575 (N_18575,N_18065,N_18296);
nor U18576 (N_18576,N_18106,N_18208);
xnor U18577 (N_18577,N_18286,N_18011);
nand U18578 (N_18578,N_18089,N_18217);
nor U18579 (N_18579,N_18326,N_18487);
nand U18580 (N_18580,N_18248,N_18077);
nor U18581 (N_18581,N_18321,N_18005);
and U18582 (N_18582,N_18432,N_18387);
xnor U18583 (N_18583,N_18018,N_18166);
xor U18584 (N_18584,N_18197,N_18473);
and U18585 (N_18585,N_18438,N_18127);
xor U18586 (N_18586,N_18193,N_18452);
nor U18587 (N_18587,N_18123,N_18076);
and U18588 (N_18588,N_18418,N_18191);
nand U18589 (N_18589,N_18221,N_18265);
nand U18590 (N_18590,N_18103,N_18220);
xor U18591 (N_18591,N_18072,N_18354);
or U18592 (N_18592,N_18470,N_18128);
and U18593 (N_18593,N_18056,N_18234);
nand U18594 (N_18594,N_18177,N_18383);
xor U18595 (N_18595,N_18068,N_18102);
nor U18596 (N_18596,N_18215,N_18136);
nand U18597 (N_18597,N_18394,N_18137);
nor U18598 (N_18598,N_18381,N_18440);
or U18599 (N_18599,N_18302,N_18004);
nand U18600 (N_18600,N_18098,N_18174);
or U18601 (N_18601,N_18210,N_18416);
nand U18602 (N_18602,N_18267,N_18138);
and U18603 (N_18603,N_18091,N_18205);
nor U18604 (N_18604,N_18211,N_18066);
nor U18605 (N_18605,N_18061,N_18038);
or U18606 (N_18606,N_18045,N_18125);
and U18607 (N_18607,N_18425,N_18255);
and U18608 (N_18608,N_18419,N_18085);
and U18609 (N_18609,N_18450,N_18259);
nand U18610 (N_18610,N_18303,N_18437);
or U18611 (N_18611,N_18342,N_18258);
nor U18612 (N_18612,N_18261,N_18275);
and U18613 (N_18613,N_18266,N_18385);
nor U18614 (N_18614,N_18475,N_18087);
or U18615 (N_18615,N_18109,N_18453);
xnor U18616 (N_18616,N_18130,N_18349);
nand U18617 (N_18617,N_18369,N_18287);
nor U18618 (N_18618,N_18042,N_18176);
nand U18619 (N_18619,N_18333,N_18201);
and U18620 (N_18620,N_18405,N_18336);
nand U18621 (N_18621,N_18339,N_18271);
xnor U18622 (N_18622,N_18270,N_18392);
nor U18623 (N_18623,N_18161,N_18058);
xnor U18624 (N_18624,N_18292,N_18455);
or U18625 (N_18625,N_18251,N_18410);
nand U18626 (N_18626,N_18388,N_18364);
nand U18627 (N_18627,N_18096,N_18107);
xor U18628 (N_18628,N_18164,N_18288);
and U18629 (N_18629,N_18122,N_18156);
xor U18630 (N_18630,N_18037,N_18315);
or U18631 (N_18631,N_18356,N_18284);
and U18632 (N_18632,N_18391,N_18115);
or U18633 (N_18633,N_18023,N_18064);
or U18634 (N_18634,N_18053,N_18082);
nor U18635 (N_18635,N_18249,N_18461);
xnor U18636 (N_18636,N_18422,N_18129);
and U18637 (N_18637,N_18375,N_18158);
or U18638 (N_18638,N_18009,N_18456);
or U18639 (N_18639,N_18463,N_18423);
nor U18640 (N_18640,N_18183,N_18498);
nand U18641 (N_18641,N_18357,N_18247);
nand U18642 (N_18642,N_18338,N_18374);
or U18643 (N_18643,N_18471,N_18134);
nor U18644 (N_18644,N_18478,N_18469);
and U18645 (N_18645,N_18273,N_18344);
and U18646 (N_18646,N_18250,N_18386);
or U18647 (N_18647,N_18482,N_18431);
xor U18648 (N_18648,N_18285,N_18294);
xnor U18649 (N_18649,N_18040,N_18243);
xor U18650 (N_18650,N_18165,N_18163);
nor U18651 (N_18651,N_18465,N_18012);
nor U18652 (N_18652,N_18030,N_18008);
nor U18653 (N_18653,N_18007,N_18476);
or U18654 (N_18654,N_18240,N_18472);
xnor U18655 (N_18655,N_18443,N_18003);
nor U18656 (N_18656,N_18132,N_18147);
nor U18657 (N_18657,N_18015,N_18341);
nor U18658 (N_18658,N_18113,N_18496);
and U18659 (N_18659,N_18307,N_18179);
or U18660 (N_18660,N_18490,N_18382);
xor U18661 (N_18661,N_18212,N_18299);
or U18662 (N_18662,N_18121,N_18196);
nor U18663 (N_18663,N_18378,N_18014);
or U18664 (N_18664,N_18457,N_18154);
and U18665 (N_18665,N_18143,N_18033);
nand U18666 (N_18666,N_18445,N_18171);
or U18667 (N_18667,N_18093,N_18466);
or U18668 (N_18668,N_18169,N_18100);
or U18669 (N_18669,N_18277,N_18276);
xor U18670 (N_18670,N_18278,N_18446);
and U18671 (N_18671,N_18495,N_18244);
or U18672 (N_18672,N_18133,N_18291);
and U18673 (N_18673,N_18047,N_18157);
xnor U18674 (N_18674,N_18046,N_18195);
nand U18675 (N_18675,N_18318,N_18020);
xor U18676 (N_18676,N_18116,N_18060);
xor U18677 (N_18677,N_18319,N_18332);
or U18678 (N_18678,N_18218,N_18035);
and U18679 (N_18679,N_18376,N_18355);
xor U18680 (N_18680,N_18439,N_18025);
nand U18681 (N_18681,N_18484,N_18260);
and U18682 (N_18682,N_18000,N_18305);
xor U18683 (N_18683,N_18233,N_18139);
nand U18684 (N_18684,N_18362,N_18379);
nand U18685 (N_18685,N_18002,N_18112);
and U18686 (N_18686,N_18159,N_18111);
or U18687 (N_18687,N_18389,N_18366);
and U18688 (N_18688,N_18222,N_18017);
nor U18689 (N_18689,N_18092,N_18359);
and U18690 (N_18690,N_18306,N_18027);
nor U18691 (N_18691,N_18409,N_18434);
or U18692 (N_18692,N_18242,N_18239);
nand U18693 (N_18693,N_18152,N_18312);
or U18694 (N_18694,N_18435,N_18236);
xnor U18695 (N_18695,N_18367,N_18272);
xor U18696 (N_18696,N_18108,N_18399);
xor U18697 (N_18697,N_18404,N_18269);
or U18698 (N_18698,N_18051,N_18063);
or U18699 (N_18699,N_18430,N_18485);
xnor U18700 (N_18700,N_18226,N_18246);
or U18701 (N_18701,N_18010,N_18428);
xor U18702 (N_18702,N_18192,N_18295);
and U18703 (N_18703,N_18370,N_18441);
or U18704 (N_18704,N_18334,N_18067);
nor U18705 (N_18705,N_18180,N_18401);
and U18706 (N_18706,N_18094,N_18462);
and U18707 (N_18707,N_18203,N_18188);
nor U18708 (N_18708,N_18257,N_18459);
nor U18709 (N_18709,N_18168,N_18329);
and U18710 (N_18710,N_18447,N_18024);
nand U18711 (N_18711,N_18316,N_18044);
nor U18712 (N_18712,N_18281,N_18442);
and U18713 (N_18713,N_18331,N_18402);
and U18714 (N_18714,N_18384,N_18477);
nand U18715 (N_18715,N_18371,N_18178);
nor U18716 (N_18716,N_18417,N_18363);
and U18717 (N_18717,N_18310,N_18048);
or U18718 (N_18718,N_18223,N_18393);
xnor U18719 (N_18719,N_18090,N_18088);
and U18720 (N_18720,N_18054,N_18224);
or U18721 (N_18721,N_18330,N_18124);
xnor U18722 (N_18722,N_18075,N_18324);
xnor U18723 (N_18723,N_18449,N_18232);
nand U18724 (N_18724,N_18322,N_18202);
and U18725 (N_18725,N_18162,N_18140);
xor U18726 (N_18726,N_18480,N_18308);
nor U18727 (N_18727,N_18494,N_18380);
xor U18728 (N_18728,N_18031,N_18204);
nand U18729 (N_18729,N_18190,N_18400);
xnor U18730 (N_18730,N_18412,N_18297);
and U18731 (N_18731,N_18120,N_18231);
or U18732 (N_18732,N_18206,N_18397);
xnor U18733 (N_18733,N_18126,N_18167);
nand U18734 (N_18734,N_18347,N_18170);
and U18735 (N_18735,N_18335,N_18230);
xnor U18736 (N_18736,N_18481,N_18194);
and U18737 (N_18737,N_18118,N_18282);
and U18738 (N_18738,N_18373,N_18398);
or U18739 (N_18739,N_18229,N_18279);
or U18740 (N_18740,N_18006,N_18050);
or U18741 (N_18741,N_18034,N_18149);
or U18742 (N_18742,N_18343,N_18074);
xor U18743 (N_18743,N_18486,N_18274);
or U18744 (N_18744,N_18403,N_18468);
nand U18745 (N_18745,N_18327,N_18448);
xnor U18746 (N_18746,N_18368,N_18427);
or U18747 (N_18747,N_18460,N_18022);
and U18748 (N_18748,N_18185,N_18227);
xor U18749 (N_18749,N_18348,N_18300);
or U18750 (N_18750,N_18121,N_18173);
nor U18751 (N_18751,N_18193,N_18219);
nor U18752 (N_18752,N_18357,N_18153);
nor U18753 (N_18753,N_18287,N_18458);
xor U18754 (N_18754,N_18144,N_18160);
nor U18755 (N_18755,N_18133,N_18245);
xor U18756 (N_18756,N_18272,N_18241);
xor U18757 (N_18757,N_18268,N_18242);
xnor U18758 (N_18758,N_18348,N_18424);
nor U18759 (N_18759,N_18289,N_18362);
xor U18760 (N_18760,N_18016,N_18094);
nand U18761 (N_18761,N_18040,N_18200);
nor U18762 (N_18762,N_18310,N_18490);
and U18763 (N_18763,N_18270,N_18183);
or U18764 (N_18764,N_18022,N_18326);
nand U18765 (N_18765,N_18050,N_18343);
and U18766 (N_18766,N_18000,N_18094);
or U18767 (N_18767,N_18076,N_18172);
or U18768 (N_18768,N_18051,N_18173);
and U18769 (N_18769,N_18433,N_18499);
or U18770 (N_18770,N_18306,N_18273);
nor U18771 (N_18771,N_18186,N_18207);
xnor U18772 (N_18772,N_18371,N_18036);
nand U18773 (N_18773,N_18260,N_18292);
nand U18774 (N_18774,N_18332,N_18048);
nand U18775 (N_18775,N_18202,N_18029);
xnor U18776 (N_18776,N_18456,N_18439);
nor U18777 (N_18777,N_18481,N_18434);
xor U18778 (N_18778,N_18242,N_18149);
nand U18779 (N_18779,N_18028,N_18285);
and U18780 (N_18780,N_18060,N_18042);
xor U18781 (N_18781,N_18483,N_18434);
nor U18782 (N_18782,N_18162,N_18315);
xnor U18783 (N_18783,N_18021,N_18254);
and U18784 (N_18784,N_18251,N_18305);
or U18785 (N_18785,N_18400,N_18322);
nor U18786 (N_18786,N_18047,N_18113);
xor U18787 (N_18787,N_18405,N_18225);
nand U18788 (N_18788,N_18033,N_18135);
or U18789 (N_18789,N_18478,N_18179);
nand U18790 (N_18790,N_18386,N_18235);
xnor U18791 (N_18791,N_18228,N_18334);
or U18792 (N_18792,N_18105,N_18147);
xor U18793 (N_18793,N_18416,N_18333);
xor U18794 (N_18794,N_18375,N_18141);
and U18795 (N_18795,N_18267,N_18089);
xnor U18796 (N_18796,N_18266,N_18142);
nor U18797 (N_18797,N_18146,N_18006);
nor U18798 (N_18798,N_18252,N_18113);
nand U18799 (N_18799,N_18263,N_18185);
nand U18800 (N_18800,N_18312,N_18432);
and U18801 (N_18801,N_18471,N_18184);
nand U18802 (N_18802,N_18480,N_18338);
nand U18803 (N_18803,N_18207,N_18118);
and U18804 (N_18804,N_18122,N_18489);
or U18805 (N_18805,N_18083,N_18066);
nor U18806 (N_18806,N_18491,N_18226);
xnor U18807 (N_18807,N_18310,N_18329);
or U18808 (N_18808,N_18359,N_18245);
nand U18809 (N_18809,N_18451,N_18301);
nand U18810 (N_18810,N_18426,N_18011);
nor U18811 (N_18811,N_18378,N_18465);
or U18812 (N_18812,N_18115,N_18062);
xnor U18813 (N_18813,N_18428,N_18432);
and U18814 (N_18814,N_18336,N_18263);
nor U18815 (N_18815,N_18294,N_18117);
and U18816 (N_18816,N_18394,N_18022);
nor U18817 (N_18817,N_18220,N_18151);
and U18818 (N_18818,N_18357,N_18318);
or U18819 (N_18819,N_18437,N_18253);
and U18820 (N_18820,N_18187,N_18240);
or U18821 (N_18821,N_18133,N_18010);
or U18822 (N_18822,N_18264,N_18212);
xor U18823 (N_18823,N_18072,N_18303);
and U18824 (N_18824,N_18379,N_18132);
nand U18825 (N_18825,N_18039,N_18001);
or U18826 (N_18826,N_18232,N_18114);
xor U18827 (N_18827,N_18032,N_18476);
nand U18828 (N_18828,N_18272,N_18461);
and U18829 (N_18829,N_18395,N_18054);
and U18830 (N_18830,N_18402,N_18159);
nor U18831 (N_18831,N_18417,N_18251);
and U18832 (N_18832,N_18182,N_18211);
and U18833 (N_18833,N_18236,N_18325);
xor U18834 (N_18834,N_18362,N_18356);
nor U18835 (N_18835,N_18495,N_18012);
and U18836 (N_18836,N_18157,N_18229);
nor U18837 (N_18837,N_18316,N_18085);
nand U18838 (N_18838,N_18130,N_18213);
or U18839 (N_18839,N_18215,N_18056);
nor U18840 (N_18840,N_18294,N_18154);
or U18841 (N_18841,N_18287,N_18246);
or U18842 (N_18842,N_18262,N_18023);
and U18843 (N_18843,N_18064,N_18455);
or U18844 (N_18844,N_18231,N_18124);
or U18845 (N_18845,N_18037,N_18246);
xor U18846 (N_18846,N_18296,N_18212);
and U18847 (N_18847,N_18483,N_18440);
xor U18848 (N_18848,N_18221,N_18145);
nor U18849 (N_18849,N_18360,N_18129);
xnor U18850 (N_18850,N_18126,N_18040);
xor U18851 (N_18851,N_18200,N_18160);
xnor U18852 (N_18852,N_18473,N_18117);
and U18853 (N_18853,N_18460,N_18395);
nor U18854 (N_18854,N_18209,N_18195);
nor U18855 (N_18855,N_18282,N_18210);
or U18856 (N_18856,N_18187,N_18017);
nor U18857 (N_18857,N_18035,N_18354);
or U18858 (N_18858,N_18384,N_18114);
and U18859 (N_18859,N_18486,N_18280);
nor U18860 (N_18860,N_18050,N_18126);
or U18861 (N_18861,N_18144,N_18441);
xnor U18862 (N_18862,N_18212,N_18290);
or U18863 (N_18863,N_18122,N_18172);
and U18864 (N_18864,N_18008,N_18443);
nand U18865 (N_18865,N_18253,N_18101);
or U18866 (N_18866,N_18169,N_18172);
nand U18867 (N_18867,N_18323,N_18009);
or U18868 (N_18868,N_18107,N_18029);
or U18869 (N_18869,N_18043,N_18224);
and U18870 (N_18870,N_18439,N_18322);
or U18871 (N_18871,N_18153,N_18162);
xnor U18872 (N_18872,N_18130,N_18119);
nor U18873 (N_18873,N_18136,N_18183);
nor U18874 (N_18874,N_18378,N_18334);
and U18875 (N_18875,N_18164,N_18078);
xnor U18876 (N_18876,N_18177,N_18308);
xnor U18877 (N_18877,N_18090,N_18408);
nor U18878 (N_18878,N_18408,N_18295);
xnor U18879 (N_18879,N_18354,N_18116);
nor U18880 (N_18880,N_18034,N_18191);
xnor U18881 (N_18881,N_18030,N_18022);
nor U18882 (N_18882,N_18171,N_18290);
nor U18883 (N_18883,N_18440,N_18252);
nor U18884 (N_18884,N_18463,N_18387);
and U18885 (N_18885,N_18264,N_18225);
xor U18886 (N_18886,N_18416,N_18435);
nor U18887 (N_18887,N_18425,N_18162);
xor U18888 (N_18888,N_18266,N_18448);
or U18889 (N_18889,N_18392,N_18251);
nor U18890 (N_18890,N_18047,N_18191);
or U18891 (N_18891,N_18024,N_18430);
nand U18892 (N_18892,N_18381,N_18186);
xnor U18893 (N_18893,N_18182,N_18219);
nor U18894 (N_18894,N_18174,N_18313);
or U18895 (N_18895,N_18323,N_18468);
nand U18896 (N_18896,N_18177,N_18297);
nand U18897 (N_18897,N_18481,N_18131);
or U18898 (N_18898,N_18016,N_18490);
nor U18899 (N_18899,N_18038,N_18126);
xor U18900 (N_18900,N_18402,N_18451);
xor U18901 (N_18901,N_18306,N_18460);
and U18902 (N_18902,N_18298,N_18300);
xor U18903 (N_18903,N_18475,N_18458);
nor U18904 (N_18904,N_18375,N_18205);
and U18905 (N_18905,N_18476,N_18059);
xnor U18906 (N_18906,N_18322,N_18099);
nor U18907 (N_18907,N_18136,N_18102);
xor U18908 (N_18908,N_18325,N_18409);
and U18909 (N_18909,N_18047,N_18494);
xor U18910 (N_18910,N_18080,N_18049);
nand U18911 (N_18911,N_18345,N_18038);
nand U18912 (N_18912,N_18105,N_18257);
nor U18913 (N_18913,N_18057,N_18357);
xor U18914 (N_18914,N_18113,N_18162);
or U18915 (N_18915,N_18488,N_18494);
nor U18916 (N_18916,N_18233,N_18260);
xnor U18917 (N_18917,N_18096,N_18234);
or U18918 (N_18918,N_18236,N_18060);
nor U18919 (N_18919,N_18369,N_18405);
nand U18920 (N_18920,N_18337,N_18464);
and U18921 (N_18921,N_18391,N_18431);
or U18922 (N_18922,N_18461,N_18170);
nand U18923 (N_18923,N_18100,N_18416);
xor U18924 (N_18924,N_18298,N_18291);
and U18925 (N_18925,N_18312,N_18135);
nand U18926 (N_18926,N_18400,N_18401);
nand U18927 (N_18927,N_18453,N_18391);
xnor U18928 (N_18928,N_18235,N_18411);
nor U18929 (N_18929,N_18222,N_18094);
xor U18930 (N_18930,N_18341,N_18250);
nand U18931 (N_18931,N_18455,N_18374);
xor U18932 (N_18932,N_18065,N_18222);
and U18933 (N_18933,N_18228,N_18110);
or U18934 (N_18934,N_18233,N_18177);
and U18935 (N_18935,N_18331,N_18434);
xor U18936 (N_18936,N_18128,N_18416);
nand U18937 (N_18937,N_18420,N_18079);
and U18938 (N_18938,N_18250,N_18434);
and U18939 (N_18939,N_18325,N_18400);
or U18940 (N_18940,N_18068,N_18111);
xnor U18941 (N_18941,N_18073,N_18245);
xnor U18942 (N_18942,N_18213,N_18459);
and U18943 (N_18943,N_18076,N_18345);
and U18944 (N_18944,N_18330,N_18290);
xor U18945 (N_18945,N_18083,N_18433);
xor U18946 (N_18946,N_18422,N_18248);
and U18947 (N_18947,N_18466,N_18162);
and U18948 (N_18948,N_18387,N_18413);
and U18949 (N_18949,N_18100,N_18466);
or U18950 (N_18950,N_18301,N_18388);
nor U18951 (N_18951,N_18450,N_18418);
xor U18952 (N_18952,N_18082,N_18209);
and U18953 (N_18953,N_18226,N_18046);
nor U18954 (N_18954,N_18125,N_18359);
and U18955 (N_18955,N_18375,N_18441);
nor U18956 (N_18956,N_18040,N_18017);
or U18957 (N_18957,N_18151,N_18327);
or U18958 (N_18958,N_18133,N_18012);
or U18959 (N_18959,N_18265,N_18048);
xnor U18960 (N_18960,N_18396,N_18062);
or U18961 (N_18961,N_18139,N_18003);
xor U18962 (N_18962,N_18493,N_18412);
nor U18963 (N_18963,N_18444,N_18071);
nand U18964 (N_18964,N_18102,N_18224);
or U18965 (N_18965,N_18024,N_18176);
nor U18966 (N_18966,N_18436,N_18019);
and U18967 (N_18967,N_18089,N_18285);
xor U18968 (N_18968,N_18304,N_18121);
nor U18969 (N_18969,N_18003,N_18234);
xnor U18970 (N_18970,N_18188,N_18285);
and U18971 (N_18971,N_18305,N_18247);
nor U18972 (N_18972,N_18351,N_18316);
or U18973 (N_18973,N_18015,N_18348);
and U18974 (N_18974,N_18279,N_18410);
and U18975 (N_18975,N_18075,N_18015);
xor U18976 (N_18976,N_18243,N_18370);
or U18977 (N_18977,N_18488,N_18289);
or U18978 (N_18978,N_18270,N_18208);
nand U18979 (N_18979,N_18097,N_18201);
and U18980 (N_18980,N_18094,N_18267);
nand U18981 (N_18981,N_18391,N_18498);
xnor U18982 (N_18982,N_18090,N_18052);
xnor U18983 (N_18983,N_18260,N_18022);
or U18984 (N_18984,N_18337,N_18098);
xor U18985 (N_18985,N_18055,N_18227);
or U18986 (N_18986,N_18082,N_18294);
nor U18987 (N_18987,N_18196,N_18212);
nand U18988 (N_18988,N_18426,N_18288);
nand U18989 (N_18989,N_18006,N_18444);
nor U18990 (N_18990,N_18497,N_18368);
nor U18991 (N_18991,N_18252,N_18262);
or U18992 (N_18992,N_18427,N_18151);
nand U18993 (N_18993,N_18174,N_18298);
or U18994 (N_18994,N_18179,N_18249);
nor U18995 (N_18995,N_18019,N_18396);
or U18996 (N_18996,N_18152,N_18375);
and U18997 (N_18997,N_18054,N_18108);
and U18998 (N_18998,N_18275,N_18417);
xor U18999 (N_18999,N_18218,N_18257);
nor U19000 (N_19000,N_18662,N_18739);
xnor U19001 (N_19001,N_18899,N_18584);
and U19002 (N_19002,N_18588,N_18842);
xnor U19003 (N_19003,N_18620,N_18952);
nand U19004 (N_19004,N_18691,N_18696);
or U19005 (N_19005,N_18617,N_18796);
nor U19006 (N_19006,N_18536,N_18520);
xor U19007 (N_19007,N_18532,N_18797);
nor U19008 (N_19008,N_18704,N_18506);
nand U19009 (N_19009,N_18823,N_18909);
nand U19010 (N_19010,N_18604,N_18992);
or U19011 (N_19011,N_18846,N_18986);
and U19012 (N_19012,N_18757,N_18682);
xnor U19013 (N_19013,N_18503,N_18512);
xor U19014 (N_19014,N_18871,N_18660);
and U19015 (N_19015,N_18609,N_18802);
nand U19016 (N_19016,N_18791,N_18607);
and U19017 (N_19017,N_18752,N_18780);
xor U19018 (N_19018,N_18618,N_18999);
or U19019 (N_19019,N_18528,N_18870);
and U19020 (N_19020,N_18906,N_18931);
xnor U19021 (N_19021,N_18991,N_18817);
nor U19022 (N_19022,N_18844,N_18728);
nand U19023 (N_19023,N_18854,N_18695);
nor U19024 (N_19024,N_18983,N_18515);
xor U19025 (N_19025,N_18897,N_18563);
xnor U19026 (N_19026,N_18890,N_18573);
nand U19027 (N_19027,N_18812,N_18546);
or U19028 (N_19028,N_18645,N_18876);
and U19029 (N_19029,N_18631,N_18715);
nand U19030 (N_19030,N_18664,N_18592);
xnor U19031 (N_19031,N_18501,N_18815);
xnor U19032 (N_19032,N_18552,N_18807);
nor U19033 (N_19033,N_18805,N_18527);
xor U19034 (N_19034,N_18721,N_18539);
xor U19035 (N_19035,N_18927,N_18700);
nor U19036 (N_19036,N_18788,N_18647);
xnor U19037 (N_19037,N_18549,N_18827);
or U19038 (N_19038,N_18679,N_18648);
nor U19039 (N_19039,N_18698,N_18525);
nor U19040 (N_19040,N_18951,N_18663);
or U19041 (N_19041,N_18633,N_18710);
nor U19042 (N_19042,N_18575,N_18530);
and U19043 (N_19043,N_18861,N_18673);
xor U19044 (N_19044,N_18705,N_18782);
nor U19045 (N_19045,N_18859,N_18767);
xor U19046 (N_19046,N_18712,N_18564);
or U19047 (N_19047,N_18824,N_18658);
nand U19048 (N_19048,N_18787,N_18774);
nand U19049 (N_19049,N_18683,N_18943);
or U19050 (N_19050,N_18822,N_18765);
and U19051 (N_19051,N_18891,N_18944);
nand U19052 (N_19052,N_18623,N_18533);
xor U19053 (N_19053,N_18930,N_18975);
nand U19054 (N_19054,N_18641,N_18997);
nand U19055 (N_19055,N_18600,N_18762);
xnor U19056 (N_19056,N_18914,N_18919);
nand U19057 (N_19057,N_18542,N_18880);
xor U19058 (N_19058,N_18723,N_18675);
nor U19059 (N_19059,N_18836,N_18887);
nor U19060 (N_19060,N_18925,N_18789);
or U19061 (N_19061,N_18534,N_18865);
or U19062 (N_19062,N_18889,N_18513);
or U19063 (N_19063,N_18637,N_18708);
and U19064 (N_19064,N_18508,N_18769);
xnor U19065 (N_19065,N_18640,N_18654);
and U19066 (N_19066,N_18760,N_18595);
or U19067 (N_19067,N_18521,N_18741);
nand U19068 (N_19068,N_18722,N_18835);
nor U19069 (N_19069,N_18763,N_18872);
or U19070 (N_19070,N_18751,N_18868);
and U19071 (N_19071,N_18828,N_18852);
or U19072 (N_19072,N_18671,N_18838);
or U19073 (N_19073,N_18699,N_18910);
and U19074 (N_19074,N_18717,N_18882);
xnor U19075 (N_19075,N_18599,N_18840);
or U19076 (N_19076,N_18616,N_18583);
nor U19077 (N_19077,N_18970,N_18858);
xnor U19078 (N_19078,N_18892,N_18638);
xor U19079 (N_19079,N_18979,N_18651);
nor U19080 (N_19080,N_18924,N_18626);
nand U19081 (N_19081,N_18684,N_18681);
and U19082 (N_19082,N_18581,N_18984);
or U19083 (N_19083,N_18948,N_18772);
nand U19084 (N_19084,N_18511,N_18524);
nand U19085 (N_19085,N_18510,N_18603);
xor U19086 (N_19086,N_18567,N_18736);
nor U19087 (N_19087,N_18937,N_18756);
xor U19088 (N_19088,N_18518,N_18965);
nand U19089 (N_19089,N_18622,N_18773);
nor U19090 (N_19090,N_18685,N_18707);
xnor U19091 (N_19091,N_18896,N_18820);
and U19092 (N_19092,N_18934,N_18571);
nor U19093 (N_19093,N_18938,N_18940);
nor U19094 (N_19094,N_18996,N_18953);
or U19095 (N_19095,N_18568,N_18956);
nor U19096 (N_19096,N_18737,N_18966);
xor U19097 (N_19097,N_18611,N_18916);
xor U19098 (N_19098,N_18615,N_18821);
nand U19099 (N_19099,N_18547,N_18507);
nor U19100 (N_19100,N_18971,N_18572);
xor U19101 (N_19101,N_18517,N_18636);
and U19102 (N_19102,N_18977,N_18540);
or U19103 (N_19103,N_18731,N_18727);
nor U19104 (N_19104,N_18693,N_18867);
or U19105 (N_19105,N_18976,N_18566);
nor U19106 (N_19106,N_18702,N_18918);
or U19107 (N_19107,N_18726,N_18612);
or U19108 (N_19108,N_18669,N_18701);
nor U19109 (N_19109,N_18509,N_18894);
or U19110 (N_19110,N_18809,N_18577);
xor U19111 (N_19111,N_18885,N_18941);
and U19112 (N_19112,N_18585,N_18869);
and U19113 (N_19113,N_18829,N_18988);
or U19114 (N_19114,N_18677,N_18987);
or U19115 (N_19115,N_18732,N_18804);
nand U19116 (N_19116,N_18900,N_18516);
nand U19117 (N_19117,N_18946,N_18863);
and U19118 (N_19118,N_18628,N_18839);
nand U19119 (N_19119,N_18860,N_18667);
or U19120 (N_19120,N_18692,N_18606);
nor U19121 (N_19121,N_18743,N_18888);
or U19122 (N_19122,N_18895,N_18740);
and U19123 (N_19123,N_18596,N_18619);
or U19124 (N_19124,N_18922,N_18911);
nand U19125 (N_19125,N_18850,N_18879);
or U19126 (N_19126,N_18605,N_18792);
and U19127 (N_19127,N_18504,N_18886);
xnor U19128 (N_19128,N_18770,N_18907);
nand U19129 (N_19129,N_18553,N_18978);
and U19130 (N_19130,N_18808,N_18947);
nand U19131 (N_19131,N_18936,N_18845);
or U19132 (N_19132,N_18557,N_18800);
or U19133 (N_19133,N_18548,N_18855);
nand U19134 (N_19134,N_18561,N_18985);
and U19135 (N_19135,N_18875,N_18634);
nor U19136 (N_19136,N_18522,N_18825);
xnor U19137 (N_19137,N_18803,N_18653);
and U19138 (N_19138,N_18874,N_18657);
nand U19139 (N_19139,N_18877,N_18519);
nor U19140 (N_19140,N_18678,N_18629);
or U19141 (N_19141,N_18958,N_18851);
nor U19142 (N_19142,N_18776,N_18543);
and U19143 (N_19143,N_18652,N_18531);
nand U19144 (N_19144,N_18714,N_18703);
nor U19145 (N_19145,N_18560,N_18690);
or U19146 (N_19146,N_18974,N_18642);
or U19147 (N_19147,N_18697,N_18841);
nand U19148 (N_19148,N_18848,N_18758);
and U19149 (N_19149,N_18749,N_18742);
nor U19150 (N_19150,N_18768,N_18748);
and U19151 (N_19151,N_18689,N_18593);
nor U19152 (N_19152,N_18643,N_18798);
nor U19153 (N_19153,N_18706,N_18720);
or U19154 (N_19154,N_18738,N_18541);
nor U19155 (N_19155,N_18917,N_18569);
xor U19156 (N_19156,N_18908,N_18687);
and U19157 (N_19157,N_18993,N_18830);
and U19158 (N_19158,N_18903,N_18810);
nand U19159 (N_19159,N_18613,N_18955);
nand U19160 (N_19160,N_18602,N_18562);
nand U19161 (N_19161,N_18949,N_18814);
nor U19162 (N_19162,N_18582,N_18793);
nor U19163 (N_19163,N_18579,N_18901);
xor U19164 (N_19164,N_18935,N_18990);
xnor U19165 (N_19165,N_18957,N_18973);
or U19166 (N_19166,N_18849,N_18995);
nand U19167 (N_19167,N_18537,N_18719);
nor U19168 (N_19168,N_18694,N_18847);
and U19169 (N_19169,N_18594,N_18811);
xor U19170 (N_19170,N_18672,N_18538);
and U19171 (N_19171,N_18725,N_18964);
nand U19172 (N_19172,N_18656,N_18790);
xor U19173 (N_19173,N_18688,N_18686);
and U19174 (N_19174,N_18665,N_18580);
nand U19175 (N_19175,N_18853,N_18754);
nand U19176 (N_19176,N_18959,N_18778);
nor U19177 (N_19177,N_18556,N_18545);
nor U19178 (N_19178,N_18905,N_18939);
nand U19179 (N_19179,N_18529,N_18576);
nand U19180 (N_19180,N_18711,N_18550);
nand U19181 (N_19181,N_18915,N_18961);
xnor U19182 (N_19182,N_18608,N_18967);
or U19183 (N_19183,N_18832,N_18866);
and U19184 (N_19184,N_18590,N_18818);
nand U19185 (N_19185,N_18801,N_18639);
nor U19186 (N_19186,N_18856,N_18873);
xor U19187 (N_19187,N_18929,N_18718);
nand U19188 (N_19188,N_18972,N_18837);
xor U19189 (N_19189,N_18932,N_18969);
nand U19190 (N_19190,N_18777,N_18551);
xor U19191 (N_19191,N_18659,N_18601);
nor U19192 (N_19192,N_18730,N_18666);
and U19193 (N_19193,N_18761,N_18942);
or U19194 (N_19194,N_18674,N_18668);
or U19195 (N_19195,N_18926,N_18650);
and U19196 (N_19196,N_18624,N_18933);
or U19197 (N_19197,N_18597,N_18826);
and U19198 (N_19198,N_18998,N_18898);
nor U19199 (N_19199,N_18555,N_18591);
xnor U19200 (N_19200,N_18745,N_18644);
nand U19201 (N_19201,N_18729,N_18716);
and U19202 (N_19202,N_18912,N_18980);
nand U19203 (N_19203,N_18733,N_18785);
or U19204 (N_19204,N_18735,N_18968);
and U19205 (N_19205,N_18746,N_18862);
nor U19206 (N_19206,N_18632,N_18630);
xnor U19207 (N_19207,N_18831,N_18535);
nand U19208 (N_19208,N_18502,N_18954);
or U19209 (N_19209,N_18813,N_18755);
or U19210 (N_19210,N_18989,N_18744);
or U19211 (N_19211,N_18794,N_18806);
and U19212 (N_19212,N_18570,N_18819);
and U19213 (N_19213,N_18923,N_18981);
and U19214 (N_19214,N_18913,N_18554);
or U19215 (N_19215,N_18565,N_18661);
nor U19216 (N_19216,N_18816,N_18621);
nand U19217 (N_19217,N_18881,N_18784);
and U19218 (N_19218,N_18878,N_18614);
xnor U19219 (N_19219,N_18625,N_18963);
nand U19220 (N_19220,N_18734,N_18982);
and U19221 (N_19221,N_18775,N_18893);
and U19222 (N_19222,N_18587,N_18500);
or U19223 (N_19223,N_18635,N_18884);
nor U19224 (N_19224,N_18526,N_18574);
and U19225 (N_19225,N_18883,N_18902);
xnor U19226 (N_19226,N_18960,N_18680);
nand U19227 (N_19227,N_18578,N_18558);
nand U19228 (N_19228,N_18786,N_18928);
or U19229 (N_19229,N_18857,N_18834);
or U19230 (N_19230,N_18781,N_18962);
nand U19231 (N_19231,N_18586,N_18589);
and U19232 (N_19232,N_18795,N_18904);
xor U19233 (N_19233,N_18724,N_18649);
xnor U19234 (N_19234,N_18994,N_18598);
nor U19235 (N_19235,N_18713,N_18523);
or U19236 (N_19236,N_18779,N_18646);
and U19237 (N_19237,N_18610,N_18753);
or U19238 (N_19238,N_18544,N_18945);
or U19239 (N_19239,N_18759,N_18833);
xnor U19240 (N_19240,N_18747,N_18514);
nand U19241 (N_19241,N_18559,N_18766);
and U19242 (N_19242,N_18799,N_18750);
or U19243 (N_19243,N_18670,N_18783);
or U19244 (N_19244,N_18655,N_18505);
nand U19245 (N_19245,N_18709,N_18920);
nand U19246 (N_19246,N_18627,N_18843);
and U19247 (N_19247,N_18764,N_18771);
and U19248 (N_19248,N_18950,N_18864);
nand U19249 (N_19249,N_18676,N_18921);
and U19250 (N_19250,N_18883,N_18517);
and U19251 (N_19251,N_18781,N_18918);
nand U19252 (N_19252,N_18739,N_18895);
and U19253 (N_19253,N_18611,N_18836);
or U19254 (N_19254,N_18944,N_18816);
nand U19255 (N_19255,N_18717,N_18720);
or U19256 (N_19256,N_18532,N_18504);
nand U19257 (N_19257,N_18769,N_18605);
xor U19258 (N_19258,N_18829,N_18951);
or U19259 (N_19259,N_18955,N_18575);
xor U19260 (N_19260,N_18782,N_18886);
or U19261 (N_19261,N_18718,N_18637);
xor U19262 (N_19262,N_18790,N_18817);
or U19263 (N_19263,N_18528,N_18773);
xnor U19264 (N_19264,N_18854,N_18732);
or U19265 (N_19265,N_18589,N_18547);
xnor U19266 (N_19266,N_18685,N_18718);
xor U19267 (N_19267,N_18999,N_18629);
nand U19268 (N_19268,N_18731,N_18997);
nor U19269 (N_19269,N_18783,N_18712);
nand U19270 (N_19270,N_18613,N_18890);
nand U19271 (N_19271,N_18981,N_18594);
nand U19272 (N_19272,N_18531,N_18809);
xor U19273 (N_19273,N_18613,N_18577);
or U19274 (N_19274,N_18827,N_18942);
and U19275 (N_19275,N_18634,N_18738);
or U19276 (N_19276,N_18872,N_18980);
and U19277 (N_19277,N_18633,N_18900);
xor U19278 (N_19278,N_18749,N_18607);
xnor U19279 (N_19279,N_18550,N_18610);
or U19280 (N_19280,N_18953,N_18697);
nor U19281 (N_19281,N_18952,N_18713);
nand U19282 (N_19282,N_18519,N_18871);
nand U19283 (N_19283,N_18511,N_18726);
or U19284 (N_19284,N_18660,N_18941);
and U19285 (N_19285,N_18844,N_18642);
or U19286 (N_19286,N_18935,N_18991);
or U19287 (N_19287,N_18541,N_18723);
nor U19288 (N_19288,N_18594,N_18921);
and U19289 (N_19289,N_18907,N_18510);
and U19290 (N_19290,N_18544,N_18777);
nand U19291 (N_19291,N_18714,N_18790);
nor U19292 (N_19292,N_18754,N_18863);
xnor U19293 (N_19293,N_18995,N_18657);
nor U19294 (N_19294,N_18932,N_18683);
nand U19295 (N_19295,N_18567,N_18530);
or U19296 (N_19296,N_18871,N_18795);
and U19297 (N_19297,N_18619,N_18577);
or U19298 (N_19298,N_18862,N_18707);
or U19299 (N_19299,N_18943,N_18661);
xnor U19300 (N_19300,N_18505,N_18802);
xnor U19301 (N_19301,N_18738,N_18548);
nor U19302 (N_19302,N_18549,N_18808);
xnor U19303 (N_19303,N_18669,N_18927);
xor U19304 (N_19304,N_18932,N_18894);
and U19305 (N_19305,N_18672,N_18512);
and U19306 (N_19306,N_18516,N_18973);
nor U19307 (N_19307,N_18822,N_18838);
nor U19308 (N_19308,N_18808,N_18803);
or U19309 (N_19309,N_18813,N_18867);
and U19310 (N_19310,N_18579,N_18898);
xor U19311 (N_19311,N_18744,N_18758);
xnor U19312 (N_19312,N_18977,N_18971);
and U19313 (N_19313,N_18501,N_18646);
xor U19314 (N_19314,N_18952,N_18533);
and U19315 (N_19315,N_18692,N_18565);
nand U19316 (N_19316,N_18931,N_18776);
and U19317 (N_19317,N_18618,N_18974);
nor U19318 (N_19318,N_18703,N_18926);
and U19319 (N_19319,N_18973,N_18576);
and U19320 (N_19320,N_18924,N_18976);
or U19321 (N_19321,N_18986,N_18634);
or U19322 (N_19322,N_18972,N_18517);
nand U19323 (N_19323,N_18952,N_18813);
or U19324 (N_19324,N_18879,N_18618);
and U19325 (N_19325,N_18984,N_18695);
xor U19326 (N_19326,N_18752,N_18728);
or U19327 (N_19327,N_18604,N_18575);
nor U19328 (N_19328,N_18633,N_18821);
xor U19329 (N_19329,N_18863,N_18675);
nand U19330 (N_19330,N_18674,N_18706);
nand U19331 (N_19331,N_18850,N_18714);
and U19332 (N_19332,N_18771,N_18712);
or U19333 (N_19333,N_18815,N_18666);
nand U19334 (N_19334,N_18629,N_18516);
or U19335 (N_19335,N_18896,N_18871);
nand U19336 (N_19336,N_18794,N_18949);
nand U19337 (N_19337,N_18770,N_18859);
nor U19338 (N_19338,N_18702,N_18876);
nand U19339 (N_19339,N_18571,N_18523);
nor U19340 (N_19340,N_18743,N_18893);
or U19341 (N_19341,N_18557,N_18743);
nand U19342 (N_19342,N_18906,N_18968);
nor U19343 (N_19343,N_18618,N_18920);
or U19344 (N_19344,N_18984,N_18762);
xnor U19345 (N_19345,N_18882,N_18532);
nand U19346 (N_19346,N_18532,N_18650);
and U19347 (N_19347,N_18752,N_18832);
xor U19348 (N_19348,N_18668,N_18926);
nand U19349 (N_19349,N_18606,N_18893);
nand U19350 (N_19350,N_18648,N_18622);
and U19351 (N_19351,N_18690,N_18781);
nand U19352 (N_19352,N_18945,N_18763);
and U19353 (N_19353,N_18570,N_18876);
and U19354 (N_19354,N_18911,N_18811);
or U19355 (N_19355,N_18530,N_18725);
nand U19356 (N_19356,N_18517,N_18709);
and U19357 (N_19357,N_18672,N_18915);
xor U19358 (N_19358,N_18685,N_18643);
nand U19359 (N_19359,N_18955,N_18974);
and U19360 (N_19360,N_18786,N_18530);
and U19361 (N_19361,N_18961,N_18802);
nor U19362 (N_19362,N_18882,N_18853);
nand U19363 (N_19363,N_18787,N_18851);
nand U19364 (N_19364,N_18950,N_18628);
nor U19365 (N_19365,N_18701,N_18607);
xnor U19366 (N_19366,N_18848,N_18529);
nor U19367 (N_19367,N_18503,N_18702);
or U19368 (N_19368,N_18990,N_18693);
or U19369 (N_19369,N_18578,N_18826);
xnor U19370 (N_19370,N_18672,N_18957);
xor U19371 (N_19371,N_18753,N_18928);
and U19372 (N_19372,N_18815,N_18598);
or U19373 (N_19373,N_18899,N_18845);
xor U19374 (N_19374,N_18961,N_18600);
xnor U19375 (N_19375,N_18803,N_18918);
or U19376 (N_19376,N_18603,N_18560);
or U19377 (N_19377,N_18984,N_18628);
nand U19378 (N_19378,N_18872,N_18770);
xor U19379 (N_19379,N_18637,N_18651);
and U19380 (N_19380,N_18566,N_18868);
and U19381 (N_19381,N_18614,N_18617);
nor U19382 (N_19382,N_18693,N_18603);
xor U19383 (N_19383,N_18881,N_18680);
nor U19384 (N_19384,N_18975,N_18915);
xor U19385 (N_19385,N_18988,N_18927);
and U19386 (N_19386,N_18546,N_18588);
nand U19387 (N_19387,N_18548,N_18917);
xor U19388 (N_19388,N_18638,N_18938);
nor U19389 (N_19389,N_18946,N_18942);
nor U19390 (N_19390,N_18788,N_18917);
or U19391 (N_19391,N_18692,N_18704);
nand U19392 (N_19392,N_18919,N_18755);
and U19393 (N_19393,N_18539,N_18602);
xnor U19394 (N_19394,N_18627,N_18743);
nand U19395 (N_19395,N_18794,N_18542);
or U19396 (N_19396,N_18713,N_18631);
nand U19397 (N_19397,N_18812,N_18750);
nand U19398 (N_19398,N_18696,N_18602);
and U19399 (N_19399,N_18608,N_18508);
xnor U19400 (N_19400,N_18770,N_18740);
and U19401 (N_19401,N_18967,N_18624);
xor U19402 (N_19402,N_18948,N_18739);
and U19403 (N_19403,N_18779,N_18631);
xor U19404 (N_19404,N_18723,N_18741);
or U19405 (N_19405,N_18583,N_18560);
xor U19406 (N_19406,N_18593,N_18592);
nand U19407 (N_19407,N_18776,N_18628);
or U19408 (N_19408,N_18817,N_18533);
nand U19409 (N_19409,N_18630,N_18987);
nor U19410 (N_19410,N_18631,N_18799);
nor U19411 (N_19411,N_18586,N_18696);
xor U19412 (N_19412,N_18584,N_18784);
xor U19413 (N_19413,N_18996,N_18959);
or U19414 (N_19414,N_18680,N_18749);
xnor U19415 (N_19415,N_18749,N_18555);
nand U19416 (N_19416,N_18512,N_18612);
xnor U19417 (N_19417,N_18924,N_18583);
xor U19418 (N_19418,N_18892,N_18748);
and U19419 (N_19419,N_18906,N_18678);
nor U19420 (N_19420,N_18632,N_18555);
or U19421 (N_19421,N_18561,N_18618);
xor U19422 (N_19422,N_18833,N_18539);
or U19423 (N_19423,N_18585,N_18704);
nor U19424 (N_19424,N_18598,N_18829);
xnor U19425 (N_19425,N_18715,N_18898);
xor U19426 (N_19426,N_18913,N_18924);
nand U19427 (N_19427,N_18827,N_18575);
nand U19428 (N_19428,N_18766,N_18556);
or U19429 (N_19429,N_18682,N_18680);
xnor U19430 (N_19430,N_18969,N_18707);
nor U19431 (N_19431,N_18922,N_18675);
or U19432 (N_19432,N_18986,N_18636);
nor U19433 (N_19433,N_18817,N_18504);
nand U19434 (N_19434,N_18812,N_18841);
nor U19435 (N_19435,N_18518,N_18682);
xnor U19436 (N_19436,N_18527,N_18638);
xor U19437 (N_19437,N_18561,N_18879);
xor U19438 (N_19438,N_18615,N_18834);
or U19439 (N_19439,N_18597,N_18544);
nor U19440 (N_19440,N_18797,N_18873);
or U19441 (N_19441,N_18654,N_18673);
nand U19442 (N_19442,N_18948,N_18634);
or U19443 (N_19443,N_18613,N_18960);
nand U19444 (N_19444,N_18613,N_18707);
and U19445 (N_19445,N_18641,N_18608);
or U19446 (N_19446,N_18692,N_18505);
or U19447 (N_19447,N_18601,N_18758);
xnor U19448 (N_19448,N_18569,N_18963);
xor U19449 (N_19449,N_18829,N_18554);
xor U19450 (N_19450,N_18980,N_18918);
nor U19451 (N_19451,N_18702,N_18964);
or U19452 (N_19452,N_18558,N_18734);
nand U19453 (N_19453,N_18798,N_18686);
xnor U19454 (N_19454,N_18831,N_18794);
or U19455 (N_19455,N_18852,N_18887);
nor U19456 (N_19456,N_18527,N_18778);
nor U19457 (N_19457,N_18761,N_18790);
nor U19458 (N_19458,N_18723,N_18603);
nand U19459 (N_19459,N_18555,N_18694);
xor U19460 (N_19460,N_18944,N_18529);
and U19461 (N_19461,N_18837,N_18815);
and U19462 (N_19462,N_18773,N_18740);
nand U19463 (N_19463,N_18581,N_18530);
xor U19464 (N_19464,N_18729,N_18551);
xnor U19465 (N_19465,N_18516,N_18778);
nand U19466 (N_19466,N_18537,N_18559);
or U19467 (N_19467,N_18522,N_18749);
nand U19468 (N_19468,N_18673,N_18794);
or U19469 (N_19469,N_18640,N_18568);
or U19470 (N_19470,N_18539,N_18752);
nand U19471 (N_19471,N_18703,N_18572);
nor U19472 (N_19472,N_18526,N_18620);
nor U19473 (N_19473,N_18923,N_18841);
or U19474 (N_19474,N_18837,N_18751);
and U19475 (N_19475,N_18551,N_18686);
nand U19476 (N_19476,N_18663,N_18841);
or U19477 (N_19477,N_18927,N_18506);
or U19478 (N_19478,N_18656,N_18769);
nand U19479 (N_19479,N_18528,N_18806);
nand U19480 (N_19480,N_18614,N_18639);
and U19481 (N_19481,N_18641,N_18850);
and U19482 (N_19482,N_18849,N_18916);
xor U19483 (N_19483,N_18787,N_18748);
and U19484 (N_19484,N_18524,N_18724);
and U19485 (N_19485,N_18828,N_18568);
and U19486 (N_19486,N_18500,N_18841);
and U19487 (N_19487,N_18503,N_18603);
and U19488 (N_19488,N_18876,N_18932);
or U19489 (N_19489,N_18603,N_18700);
or U19490 (N_19490,N_18980,N_18950);
xnor U19491 (N_19491,N_18695,N_18939);
and U19492 (N_19492,N_18943,N_18637);
xor U19493 (N_19493,N_18794,N_18644);
or U19494 (N_19494,N_18520,N_18942);
and U19495 (N_19495,N_18959,N_18618);
and U19496 (N_19496,N_18810,N_18590);
or U19497 (N_19497,N_18716,N_18601);
xnor U19498 (N_19498,N_18714,N_18764);
nor U19499 (N_19499,N_18701,N_18766);
xnor U19500 (N_19500,N_19477,N_19068);
or U19501 (N_19501,N_19087,N_19111);
xnor U19502 (N_19502,N_19061,N_19108);
and U19503 (N_19503,N_19252,N_19251);
xor U19504 (N_19504,N_19362,N_19323);
nor U19505 (N_19505,N_19003,N_19352);
and U19506 (N_19506,N_19194,N_19160);
and U19507 (N_19507,N_19063,N_19272);
nand U19508 (N_19508,N_19257,N_19421);
nand U19509 (N_19509,N_19171,N_19036);
nor U19510 (N_19510,N_19426,N_19298);
nand U19511 (N_19511,N_19007,N_19196);
nand U19512 (N_19512,N_19079,N_19182);
or U19513 (N_19513,N_19231,N_19057);
and U19514 (N_19514,N_19374,N_19330);
and U19515 (N_19515,N_19453,N_19433);
and U19516 (N_19516,N_19254,N_19150);
nor U19517 (N_19517,N_19456,N_19205);
nor U19518 (N_19518,N_19176,N_19288);
nand U19519 (N_19519,N_19100,N_19186);
xor U19520 (N_19520,N_19371,N_19417);
nor U19521 (N_19521,N_19141,N_19005);
nor U19522 (N_19522,N_19071,N_19134);
xor U19523 (N_19523,N_19304,N_19183);
nor U19524 (N_19524,N_19066,N_19219);
nand U19525 (N_19525,N_19064,N_19101);
xnor U19526 (N_19526,N_19173,N_19048);
xor U19527 (N_19527,N_19436,N_19415);
nor U19528 (N_19528,N_19490,N_19399);
nor U19529 (N_19529,N_19314,N_19143);
nand U19530 (N_19530,N_19412,N_19070);
nor U19531 (N_19531,N_19130,N_19318);
and U19532 (N_19532,N_19457,N_19467);
nor U19533 (N_19533,N_19306,N_19215);
nand U19534 (N_19534,N_19309,N_19259);
nor U19535 (N_19535,N_19075,N_19497);
and U19536 (N_19536,N_19459,N_19460);
nand U19537 (N_19537,N_19326,N_19225);
or U19538 (N_19538,N_19166,N_19344);
xnor U19539 (N_19539,N_19378,N_19324);
nor U19540 (N_19540,N_19043,N_19207);
or U19541 (N_19541,N_19125,N_19010);
and U19542 (N_19542,N_19368,N_19062);
xor U19543 (N_19543,N_19138,N_19423);
or U19544 (N_19544,N_19103,N_19494);
or U19545 (N_19545,N_19076,N_19422);
nand U19546 (N_19546,N_19105,N_19132);
nand U19547 (N_19547,N_19046,N_19136);
and U19548 (N_19548,N_19384,N_19260);
nor U19549 (N_19549,N_19340,N_19290);
nand U19550 (N_19550,N_19157,N_19337);
nor U19551 (N_19551,N_19303,N_19473);
xnor U19552 (N_19552,N_19077,N_19409);
nand U19553 (N_19553,N_19414,N_19250);
nand U19554 (N_19554,N_19404,N_19391);
nand U19555 (N_19555,N_19156,N_19109);
nand U19556 (N_19556,N_19275,N_19220);
and U19557 (N_19557,N_19223,N_19310);
nor U19558 (N_19558,N_19090,N_19361);
and U19559 (N_19559,N_19491,N_19055);
xnor U19560 (N_19560,N_19214,N_19284);
nand U19561 (N_19561,N_19047,N_19406);
xor U19562 (N_19562,N_19307,N_19359);
nand U19563 (N_19563,N_19299,N_19441);
nor U19564 (N_19564,N_19442,N_19488);
or U19565 (N_19565,N_19073,N_19475);
nor U19566 (N_19566,N_19249,N_19216);
nand U19567 (N_19567,N_19451,N_19319);
nand U19568 (N_19568,N_19386,N_19498);
and U19569 (N_19569,N_19294,N_19327);
nor U19570 (N_19570,N_19271,N_19499);
xor U19571 (N_19571,N_19121,N_19006);
and U19572 (N_19572,N_19458,N_19293);
and U19573 (N_19573,N_19235,N_19218);
or U19574 (N_19574,N_19316,N_19280);
or U19575 (N_19575,N_19297,N_19363);
nor U19576 (N_19576,N_19440,N_19204);
nor U19577 (N_19577,N_19434,N_19067);
xor U19578 (N_19578,N_19405,N_19237);
and U19579 (N_19579,N_19487,N_19408);
and U19580 (N_19580,N_19169,N_19276);
and U19581 (N_19581,N_19081,N_19206);
xnor U19582 (N_19582,N_19245,N_19479);
or U19583 (N_19583,N_19455,N_19263);
nand U19584 (N_19584,N_19325,N_19483);
xor U19585 (N_19585,N_19334,N_19202);
nand U19586 (N_19586,N_19292,N_19261);
or U19587 (N_19587,N_19464,N_19198);
xor U19588 (N_19588,N_19354,N_19140);
nand U19589 (N_19589,N_19184,N_19001);
xnor U19590 (N_19590,N_19112,N_19088);
xor U19591 (N_19591,N_19239,N_19044);
nand U19592 (N_19592,N_19230,N_19084);
nor U19593 (N_19593,N_19233,N_19489);
nor U19594 (N_19594,N_19031,N_19102);
or U19595 (N_19595,N_19347,N_19339);
xnor U19596 (N_19596,N_19411,N_19170);
nor U19597 (N_19597,N_19356,N_19152);
and U19598 (N_19598,N_19387,N_19364);
xnor U19599 (N_19599,N_19097,N_19353);
xnor U19600 (N_19600,N_19454,N_19165);
nand U19601 (N_19601,N_19243,N_19045);
xnor U19602 (N_19602,N_19246,N_19013);
and U19603 (N_19603,N_19056,N_19060);
and U19604 (N_19604,N_19129,N_19258);
nand U19605 (N_19605,N_19366,N_19492);
xnor U19606 (N_19606,N_19311,N_19039);
nand U19607 (N_19607,N_19383,N_19117);
xor U19608 (N_19608,N_19278,N_19486);
and U19609 (N_19609,N_19248,N_19450);
or U19610 (N_19610,N_19301,N_19159);
nand U19611 (N_19611,N_19098,N_19185);
nand U19612 (N_19612,N_19015,N_19443);
nand U19613 (N_19613,N_19395,N_19179);
nor U19614 (N_19614,N_19192,N_19190);
xor U19615 (N_19615,N_19026,N_19094);
nor U19616 (N_19616,N_19267,N_19470);
nor U19617 (N_19617,N_19093,N_19148);
nand U19618 (N_19618,N_19131,N_19480);
nand U19619 (N_19619,N_19322,N_19213);
nor U19620 (N_19620,N_19191,N_19282);
or U19621 (N_19621,N_19123,N_19266);
or U19622 (N_19622,N_19168,N_19200);
nand U19623 (N_19623,N_19242,N_19004);
xnor U19624 (N_19624,N_19446,N_19462);
or U19625 (N_19625,N_19028,N_19270);
or U19626 (N_19626,N_19020,N_19142);
or U19627 (N_19627,N_19493,N_19447);
and U19628 (N_19628,N_19424,N_19355);
xor U19629 (N_19629,N_19244,N_19277);
and U19630 (N_19630,N_19208,N_19124);
nand U19631 (N_19631,N_19420,N_19402);
nor U19632 (N_19632,N_19014,N_19413);
or U19633 (N_19633,N_19153,N_19040);
nor U19634 (N_19634,N_19343,N_19178);
or U19635 (N_19635,N_19471,N_19034);
nand U19636 (N_19636,N_19401,N_19195);
xor U19637 (N_19637,N_19320,N_19137);
xor U19638 (N_19638,N_19285,N_19188);
xor U19639 (N_19639,N_19133,N_19177);
or U19640 (N_19640,N_19086,N_19238);
xor U19641 (N_19641,N_19351,N_19002);
xor U19642 (N_19642,N_19114,N_19050);
and U19643 (N_19643,N_19172,N_19255);
or U19644 (N_19644,N_19315,N_19011);
nand U19645 (N_19645,N_19174,N_19302);
nor U19646 (N_19646,N_19381,N_19438);
and U19647 (N_19647,N_19146,N_19078);
and U19648 (N_19648,N_19052,N_19466);
nand U19649 (N_19649,N_19432,N_19469);
nand U19650 (N_19650,N_19478,N_19211);
nor U19651 (N_19651,N_19106,N_19122);
nand U19652 (N_19652,N_19264,N_19396);
nor U19653 (N_19653,N_19126,N_19080);
xnor U19654 (N_19654,N_19448,N_19189);
or U19655 (N_19655,N_19041,N_19092);
and U19656 (N_19656,N_19342,N_19328);
and U19657 (N_19657,N_19350,N_19127);
nand U19658 (N_19658,N_19449,N_19300);
nor U19659 (N_19659,N_19358,N_19388);
xor U19660 (N_19660,N_19229,N_19461);
and U19661 (N_19661,N_19379,N_19147);
xor U19662 (N_19662,N_19030,N_19308);
xor U19663 (N_19663,N_19390,N_19472);
and U19664 (N_19664,N_19145,N_19104);
nand U19665 (N_19665,N_19349,N_19181);
nor U19666 (N_19666,N_19279,N_19096);
nor U19667 (N_19667,N_19369,N_19370);
nand U19668 (N_19668,N_19289,N_19445);
nor U19669 (N_19669,N_19203,N_19268);
nand U19670 (N_19670,N_19247,N_19021);
or U19671 (N_19671,N_19099,N_19049);
nand U19672 (N_19672,N_19348,N_19199);
or U19673 (N_19673,N_19033,N_19212);
nor U19674 (N_19674,N_19485,N_19341);
or U19675 (N_19675,N_19017,N_19089);
nand U19676 (N_19676,N_19042,N_19222);
xnor U19677 (N_19677,N_19221,N_19385);
or U19678 (N_19678,N_19241,N_19360);
and U19679 (N_19679,N_19435,N_19180);
nor U19680 (N_19680,N_19025,N_19425);
nor U19681 (N_19681,N_19397,N_19407);
and U19682 (N_19682,N_19167,N_19365);
nor U19683 (N_19683,N_19269,N_19008);
nand U19684 (N_19684,N_19429,N_19256);
or U19685 (N_19685,N_19481,N_19154);
or U19686 (N_19686,N_19135,N_19286);
xor U19687 (N_19687,N_19474,N_19296);
nand U19688 (N_19688,N_19305,N_19037);
xor U19689 (N_19689,N_19430,N_19476);
or U19690 (N_19690,N_19382,N_19463);
nand U19691 (N_19691,N_19394,N_19163);
or U19692 (N_19692,N_19035,N_19149);
and U19693 (N_19693,N_19016,N_19465);
or U19694 (N_19694,N_19074,N_19346);
nand U19695 (N_19695,N_19444,N_19051);
xnor U19696 (N_19696,N_19228,N_19317);
or U19697 (N_19697,N_19437,N_19357);
or U19698 (N_19698,N_19119,N_19291);
and U19699 (N_19699,N_19193,N_19265);
or U19700 (N_19700,N_19377,N_19253);
xnor U19701 (N_19701,N_19018,N_19336);
or U19702 (N_19702,N_19439,N_19116);
or U19703 (N_19703,N_19333,N_19329);
and U19704 (N_19704,N_19029,N_19283);
nor U19705 (N_19705,N_19226,N_19452);
or U19706 (N_19706,N_19162,N_19115);
xor U19707 (N_19707,N_19495,N_19287);
nor U19708 (N_19708,N_19000,N_19083);
and U19709 (N_19709,N_19331,N_19120);
xnor U19710 (N_19710,N_19038,N_19091);
or U19711 (N_19711,N_19095,N_19295);
and U19712 (N_19712,N_19058,N_19022);
nand U19713 (N_19713,N_19069,N_19321);
nand U19714 (N_19714,N_19032,N_19201);
xnor U19715 (N_19715,N_19164,N_19155);
xor U19716 (N_19716,N_19151,N_19427);
nor U19717 (N_19717,N_19054,N_19376);
nor U19718 (N_19718,N_19281,N_19273);
or U19719 (N_19719,N_19367,N_19012);
nor U19720 (N_19720,N_19161,N_19335);
nor U19721 (N_19721,N_19082,N_19338);
and U19722 (N_19722,N_19113,N_19240);
nor U19723 (N_19723,N_19024,N_19065);
nor U19724 (N_19724,N_19389,N_19234);
nand U19725 (N_19725,N_19175,N_19232);
nor U19726 (N_19726,N_19009,N_19053);
and U19727 (N_19727,N_19375,N_19236);
nor U19728 (N_19728,N_19345,N_19313);
and U19729 (N_19729,N_19393,N_19428);
nor U19730 (N_19730,N_19410,N_19118);
or U19731 (N_19731,N_19400,N_19372);
nand U19732 (N_19732,N_19332,N_19380);
or U19733 (N_19733,N_19392,N_19027);
and U19734 (N_19734,N_19210,N_19059);
nor U19735 (N_19735,N_19482,N_19023);
and U19736 (N_19736,N_19416,N_19139);
xnor U19737 (N_19737,N_19262,N_19403);
nand U19738 (N_19738,N_19468,N_19110);
xor U19739 (N_19739,N_19274,N_19197);
xor U19740 (N_19740,N_19224,N_19496);
or U19741 (N_19741,N_19107,N_19227);
and U19742 (N_19742,N_19187,N_19085);
xor U19743 (N_19743,N_19217,N_19144);
or U19744 (N_19744,N_19431,N_19312);
nor U19745 (N_19745,N_19128,N_19484);
and U19746 (N_19746,N_19418,N_19158);
and U19747 (N_19747,N_19072,N_19398);
xnor U19748 (N_19748,N_19419,N_19373);
or U19749 (N_19749,N_19209,N_19019);
nand U19750 (N_19750,N_19223,N_19047);
or U19751 (N_19751,N_19145,N_19196);
nand U19752 (N_19752,N_19397,N_19320);
nor U19753 (N_19753,N_19409,N_19282);
and U19754 (N_19754,N_19260,N_19264);
xor U19755 (N_19755,N_19272,N_19089);
or U19756 (N_19756,N_19417,N_19492);
nor U19757 (N_19757,N_19010,N_19064);
and U19758 (N_19758,N_19342,N_19099);
nor U19759 (N_19759,N_19418,N_19256);
nor U19760 (N_19760,N_19326,N_19125);
or U19761 (N_19761,N_19358,N_19251);
nand U19762 (N_19762,N_19280,N_19432);
and U19763 (N_19763,N_19188,N_19235);
and U19764 (N_19764,N_19315,N_19362);
or U19765 (N_19765,N_19337,N_19391);
nor U19766 (N_19766,N_19158,N_19435);
nand U19767 (N_19767,N_19340,N_19343);
or U19768 (N_19768,N_19477,N_19226);
nand U19769 (N_19769,N_19298,N_19162);
nand U19770 (N_19770,N_19472,N_19334);
or U19771 (N_19771,N_19060,N_19221);
and U19772 (N_19772,N_19173,N_19097);
xor U19773 (N_19773,N_19072,N_19235);
or U19774 (N_19774,N_19027,N_19371);
or U19775 (N_19775,N_19493,N_19023);
and U19776 (N_19776,N_19271,N_19360);
xor U19777 (N_19777,N_19243,N_19216);
xnor U19778 (N_19778,N_19273,N_19402);
and U19779 (N_19779,N_19398,N_19052);
or U19780 (N_19780,N_19317,N_19150);
nor U19781 (N_19781,N_19179,N_19154);
xor U19782 (N_19782,N_19114,N_19362);
and U19783 (N_19783,N_19237,N_19327);
nor U19784 (N_19784,N_19409,N_19005);
or U19785 (N_19785,N_19124,N_19219);
and U19786 (N_19786,N_19283,N_19416);
or U19787 (N_19787,N_19270,N_19193);
nand U19788 (N_19788,N_19199,N_19268);
and U19789 (N_19789,N_19041,N_19487);
and U19790 (N_19790,N_19336,N_19189);
or U19791 (N_19791,N_19087,N_19003);
nand U19792 (N_19792,N_19056,N_19009);
nand U19793 (N_19793,N_19070,N_19402);
xor U19794 (N_19794,N_19459,N_19351);
nand U19795 (N_19795,N_19096,N_19034);
and U19796 (N_19796,N_19425,N_19034);
nand U19797 (N_19797,N_19227,N_19079);
xnor U19798 (N_19798,N_19163,N_19124);
nor U19799 (N_19799,N_19159,N_19470);
xnor U19800 (N_19800,N_19027,N_19425);
or U19801 (N_19801,N_19068,N_19401);
nand U19802 (N_19802,N_19330,N_19409);
nand U19803 (N_19803,N_19395,N_19459);
nor U19804 (N_19804,N_19039,N_19093);
and U19805 (N_19805,N_19350,N_19381);
xor U19806 (N_19806,N_19406,N_19213);
nand U19807 (N_19807,N_19097,N_19319);
or U19808 (N_19808,N_19435,N_19339);
xor U19809 (N_19809,N_19359,N_19015);
xor U19810 (N_19810,N_19046,N_19202);
and U19811 (N_19811,N_19257,N_19031);
or U19812 (N_19812,N_19273,N_19303);
or U19813 (N_19813,N_19104,N_19418);
nand U19814 (N_19814,N_19024,N_19263);
xnor U19815 (N_19815,N_19080,N_19045);
nand U19816 (N_19816,N_19105,N_19160);
and U19817 (N_19817,N_19006,N_19204);
nand U19818 (N_19818,N_19276,N_19170);
nand U19819 (N_19819,N_19244,N_19273);
or U19820 (N_19820,N_19443,N_19075);
nor U19821 (N_19821,N_19138,N_19222);
nand U19822 (N_19822,N_19099,N_19320);
and U19823 (N_19823,N_19340,N_19203);
xnor U19824 (N_19824,N_19197,N_19083);
xor U19825 (N_19825,N_19064,N_19082);
nand U19826 (N_19826,N_19228,N_19319);
nor U19827 (N_19827,N_19445,N_19226);
and U19828 (N_19828,N_19477,N_19070);
or U19829 (N_19829,N_19382,N_19285);
nand U19830 (N_19830,N_19327,N_19205);
and U19831 (N_19831,N_19480,N_19002);
nand U19832 (N_19832,N_19043,N_19245);
and U19833 (N_19833,N_19166,N_19219);
nor U19834 (N_19834,N_19427,N_19165);
and U19835 (N_19835,N_19463,N_19352);
nand U19836 (N_19836,N_19169,N_19199);
or U19837 (N_19837,N_19036,N_19149);
xor U19838 (N_19838,N_19424,N_19002);
nand U19839 (N_19839,N_19416,N_19441);
nand U19840 (N_19840,N_19493,N_19184);
nand U19841 (N_19841,N_19072,N_19007);
xor U19842 (N_19842,N_19470,N_19005);
xor U19843 (N_19843,N_19307,N_19018);
xor U19844 (N_19844,N_19111,N_19086);
and U19845 (N_19845,N_19404,N_19227);
nor U19846 (N_19846,N_19373,N_19473);
nand U19847 (N_19847,N_19205,N_19219);
nand U19848 (N_19848,N_19344,N_19479);
nand U19849 (N_19849,N_19394,N_19165);
nor U19850 (N_19850,N_19476,N_19436);
nand U19851 (N_19851,N_19200,N_19190);
xor U19852 (N_19852,N_19116,N_19121);
nand U19853 (N_19853,N_19045,N_19322);
nor U19854 (N_19854,N_19108,N_19039);
or U19855 (N_19855,N_19485,N_19307);
or U19856 (N_19856,N_19361,N_19460);
and U19857 (N_19857,N_19249,N_19212);
and U19858 (N_19858,N_19350,N_19035);
xnor U19859 (N_19859,N_19472,N_19252);
nand U19860 (N_19860,N_19057,N_19160);
nand U19861 (N_19861,N_19128,N_19074);
or U19862 (N_19862,N_19344,N_19084);
and U19863 (N_19863,N_19314,N_19195);
and U19864 (N_19864,N_19370,N_19015);
and U19865 (N_19865,N_19460,N_19385);
nand U19866 (N_19866,N_19310,N_19228);
nand U19867 (N_19867,N_19226,N_19361);
or U19868 (N_19868,N_19024,N_19171);
and U19869 (N_19869,N_19130,N_19166);
or U19870 (N_19870,N_19404,N_19302);
nor U19871 (N_19871,N_19254,N_19241);
and U19872 (N_19872,N_19026,N_19239);
nand U19873 (N_19873,N_19379,N_19273);
xor U19874 (N_19874,N_19308,N_19189);
and U19875 (N_19875,N_19150,N_19365);
and U19876 (N_19876,N_19306,N_19025);
or U19877 (N_19877,N_19430,N_19144);
xor U19878 (N_19878,N_19405,N_19447);
nor U19879 (N_19879,N_19389,N_19100);
nor U19880 (N_19880,N_19266,N_19401);
nand U19881 (N_19881,N_19220,N_19172);
nand U19882 (N_19882,N_19393,N_19260);
xnor U19883 (N_19883,N_19095,N_19196);
or U19884 (N_19884,N_19412,N_19461);
nor U19885 (N_19885,N_19002,N_19014);
or U19886 (N_19886,N_19497,N_19060);
nor U19887 (N_19887,N_19161,N_19251);
and U19888 (N_19888,N_19467,N_19339);
xor U19889 (N_19889,N_19026,N_19266);
nand U19890 (N_19890,N_19338,N_19351);
nor U19891 (N_19891,N_19378,N_19142);
nand U19892 (N_19892,N_19040,N_19471);
and U19893 (N_19893,N_19052,N_19397);
xor U19894 (N_19894,N_19438,N_19316);
and U19895 (N_19895,N_19204,N_19484);
and U19896 (N_19896,N_19023,N_19029);
and U19897 (N_19897,N_19126,N_19369);
nor U19898 (N_19898,N_19114,N_19333);
and U19899 (N_19899,N_19394,N_19159);
xnor U19900 (N_19900,N_19112,N_19189);
nor U19901 (N_19901,N_19369,N_19104);
nand U19902 (N_19902,N_19316,N_19379);
or U19903 (N_19903,N_19418,N_19007);
xor U19904 (N_19904,N_19217,N_19095);
xnor U19905 (N_19905,N_19036,N_19452);
nor U19906 (N_19906,N_19276,N_19188);
nor U19907 (N_19907,N_19130,N_19116);
nand U19908 (N_19908,N_19481,N_19466);
or U19909 (N_19909,N_19058,N_19367);
xnor U19910 (N_19910,N_19294,N_19367);
or U19911 (N_19911,N_19338,N_19116);
or U19912 (N_19912,N_19474,N_19235);
nor U19913 (N_19913,N_19156,N_19267);
nand U19914 (N_19914,N_19217,N_19350);
and U19915 (N_19915,N_19035,N_19398);
nor U19916 (N_19916,N_19024,N_19418);
nor U19917 (N_19917,N_19045,N_19073);
nand U19918 (N_19918,N_19068,N_19000);
nand U19919 (N_19919,N_19102,N_19411);
xnor U19920 (N_19920,N_19296,N_19054);
nor U19921 (N_19921,N_19288,N_19192);
xnor U19922 (N_19922,N_19486,N_19282);
and U19923 (N_19923,N_19399,N_19069);
or U19924 (N_19924,N_19219,N_19317);
and U19925 (N_19925,N_19184,N_19326);
or U19926 (N_19926,N_19005,N_19485);
nor U19927 (N_19927,N_19158,N_19411);
or U19928 (N_19928,N_19270,N_19345);
xor U19929 (N_19929,N_19350,N_19191);
or U19930 (N_19930,N_19416,N_19217);
xnor U19931 (N_19931,N_19125,N_19232);
and U19932 (N_19932,N_19013,N_19388);
and U19933 (N_19933,N_19137,N_19007);
xor U19934 (N_19934,N_19371,N_19232);
nand U19935 (N_19935,N_19170,N_19161);
xnor U19936 (N_19936,N_19171,N_19231);
xnor U19937 (N_19937,N_19210,N_19297);
xor U19938 (N_19938,N_19349,N_19313);
or U19939 (N_19939,N_19230,N_19093);
nand U19940 (N_19940,N_19135,N_19485);
nand U19941 (N_19941,N_19455,N_19019);
nand U19942 (N_19942,N_19487,N_19039);
xnor U19943 (N_19943,N_19300,N_19298);
nand U19944 (N_19944,N_19255,N_19106);
or U19945 (N_19945,N_19228,N_19320);
and U19946 (N_19946,N_19071,N_19347);
nor U19947 (N_19947,N_19383,N_19133);
or U19948 (N_19948,N_19450,N_19108);
or U19949 (N_19949,N_19067,N_19389);
or U19950 (N_19950,N_19486,N_19178);
xnor U19951 (N_19951,N_19180,N_19304);
nor U19952 (N_19952,N_19121,N_19144);
nand U19953 (N_19953,N_19008,N_19031);
or U19954 (N_19954,N_19389,N_19479);
or U19955 (N_19955,N_19173,N_19222);
nor U19956 (N_19956,N_19093,N_19168);
xor U19957 (N_19957,N_19294,N_19444);
nand U19958 (N_19958,N_19453,N_19490);
or U19959 (N_19959,N_19386,N_19119);
and U19960 (N_19960,N_19188,N_19198);
or U19961 (N_19961,N_19374,N_19390);
and U19962 (N_19962,N_19384,N_19236);
nor U19963 (N_19963,N_19125,N_19031);
or U19964 (N_19964,N_19282,N_19398);
or U19965 (N_19965,N_19002,N_19069);
nor U19966 (N_19966,N_19161,N_19457);
and U19967 (N_19967,N_19415,N_19240);
nand U19968 (N_19968,N_19000,N_19318);
xor U19969 (N_19969,N_19208,N_19220);
or U19970 (N_19970,N_19016,N_19024);
nor U19971 (N_19971,N_19415,N_19461);
or U19972 (N_19972,N_19309,N_19401);
nor U19973 (N_19973,N_19312,N_19145);
or U19974 (N_19974,N_19228,N_19298);
nor U19975 (N_19975,N_19351,N_19309);
xnor U19976 (N_19976,N_19000,N_19073);
nand U19977 (N_19977,N_19054,N_19460);
xnor U19978 (N_19978,N_19334,N_19243);
or U19979 (N_19979,N_19123,N_19052);
xor U19980 (N_19980,N_19487,N_19007);
xnor U19981 (N_19981,N_19406,N_19223);
nor U19982 (N_19982,N_19198,N_19325);
xor U19983 (N_19983,N_19035,N_19384);
xor U19984 (N_19984,N_19148,N_19303);
and U19985 (N_19985,N_19321,N_19013);
or U19986 (N_19986,N_19428,N_19496);
xor U19987 (N_19987,N_19281,N_19041);
or U19988 (N_19988,N_19290,N_19071);
or U19989 (N_19989,N_19133,N_19376);
nand U19990 (N_19990,N_19002,N_19339);
nor U19991 (N_19991,N_19118,N_19144);
and U19992 (N_19992,N_19080,N_19429);
and U19993 (N_19993,N_19199,N_19306);
nand U19994 (N_19994,N_19194,N_19053);
or U19995 (N_19995,N_19065,N_19364);
or U19996 (N_19996,N_19214,N_19354);
or U19997 (N_19997,N_19434,N_19017);
xor U19998 (N_19998,N_19355,N_19028);
xnor U19999 (N_19999,N_19060,N_19237);
or U20000 (N_20000,N_19661,N_19803);
xor U20001 (N_20001,N_19630,N_19825);
or U20002 (N_20002,N_19995,N_19504);
and U20003 (N_20003,N_19889,N_19758);
nor U20004 (N_20004,N_19975,N_19546);
nor U20005 (N_20005,N_19823,N_19943);
nand U20006 (N_20006,N_19531,N_19977);
xnor U20007 (N_20007,N_19936,N_19719);
and U20008 (N_20008,N_19533,N_19515);
xor U20009 (N_20009,N_19767,N_19784);
nand U20010 (N_20010,N_19513,N_19932);
nand U20011 (N_20011,N_19848,N_19904);
xor U20012 (N_20012,N_19739,N_19846);
and U20013 (N_20013,N_19884,N_19723);
nand U20014 (N_20014,N_19711,N_19587);
xnor U20015 (N_20015,N_19981,N_19813);
nor U20016 (N_20016,N_19576,N_19826);
nand U20017 (N_20017,N_19686,N_19987);
or U20018 (N_20018,N_19658,N_19636);
nand U20019 (N_20019,N_19725,N_19754);
nand U20020 (N_20020,N_19600,N_19616);
and U20021 (N_20021,N_19738,N_19762);
and U20022 (N_20022,N_19613,N_19831);
xnor U20023 (N_20023,N_19898,N_19949);
nor U20024 (N_20024,N_19908,N_19860);
nand U20025 (N_20025,N_19522,N_19935);
xnor U20026 (N_20026,N_19525,N_19700);
xor U20027 (N_20027,N_19964,N_19907);
or U20028 (N_20028,N_19714,N_19772);
xor U20029 (N_20029,N_19953,N_19957);
nand U20030 (N_20030,N_19877,N_19956);
or U20031 (N_20031,N_19548,N_19588);
or U20032 (N_20032,N_19891,N_19693);
or U20033 (N_20033,N_19972,N_19742);
and U20034 (N_20034,N_19748,N_19926);
xor U20035 (N_20035,N_19500,N_19992);
xor U20036 (N_20036,N_19710,N_19996);
or U20037 (N_20037,N_19580,N_19890);
and U20038 (N_20038,N_19555,N_19905);
or U20039 (N_20039,N_19578,N_19712);
xnor U20040 (N_20040,N_19770,N_19925);
nor U20041 (N_20041,N_19735,N_19763);
or U20042 (N_20042,N_19607,N_19844);
xor U20043 (N_20043,N_19947,N_19968);
nand U20044 (N_20044,N_19573,N_19961);
or U20045 (N_20045,N_19629,N_19717);
or U20046 (N_20046,N_19986,N_19800);
nand U20047 (N_20047,N_19539,N_19791);
nor U20048 (N_20048,N_19866,N_19785);
and U20049 (N_20049,N_19796,N_19871);
nor U20050 (N_20050,N_19601,N_19535);
or U20051 (N_20051,N_19773,N_19617);
or U20052 (N_20052,N_19612,N_19918);
xor U20053 (N_20053,N_19523,N_19635);
or U20054 (N_20054,N_19856,N_19776);
nor U20055 (N_20055,N_19683,N_19520);
nand U20056 (N_20056,N_19798,N_19913);
or U20057 (N_20057,N_19816,N_19955);
or U20058 (N_20058,N_19879,N_19868);
or U20059 (N_20059,N_19506,N_19649);
and U20060 (N_20060,N_19878,N_19537);
or U20061 (N_20061,N_19627,N_19745);
and U20062 (N_20062,N_19808,N_19632);
nand U20063 (N_20063,N_19978,N_19579);
or U20064 (N_20064,N_19792,N_19900);
nor U20065 (N_20065,N_19863,N_19609);
or U20066 (N_20066,N_19849,N_19509);
xor U20067 (N_20067,N_19681,N_19512);
nand U20068 (N_20068,N_19611,N_19851);
xnor U20069 (N_20069,N_19646,N_19881);
xnor U20070 (N_20070,N_19916,N_19757);
xor U20071 (N_20071,N_19931,N_19702);
nor U20072 (N_20072,N_19669,N_19603);
and U20073 (N_20073,N_19673,N_19641);
nor U20074 (N_20074,N_19944,N_19586);
nor U20075 (N_20075,N_19809,N_19746);
or U20076 (N_20076,N_19760,N_19692);
nand U20077 (N_20077,N_19701,N_19960);
or U20078 (N_20078,N_19511,N_19761);
and U20079 (N_20079,N_19648,N_19730);
xor U20080 (N_20080,N_19678,N_19790);
and U20081 (N_20081,N_19885,N_19778);
nand U20082 (N_20082,N_19680,N_19793);
nand U20083 (N_20083,N_19747,N_19989);
and U20084 (N_20084,N_19510,N_19843);
nor U20085 (N_20085,N_19842,N_19556);
nor U20086 (N_20086,N_19896,N_19590);
or U20087 (N_20087,N_19728,N_19558);
and U20088 (N_20088,N_19861,N_19945);
nor U20089 (N_20089,N_19715,N_19724);
xor U20090 (N_20090,N_19937,N_19731);
and U20091 (N_20091,N_19857,N_19503);
or U20092 (N_20092,N_19815,N_19619);
nand U20093 (N_20093,N_19951,N_19922);
xor U20094 (N_20094,N_19672,N_19838);
nand U20095 (N_20095,N_19777,N_19565);
nand U20096 (N_20096,N_19709,N_19832);
or U20097 (N_20097,N_19697,N_19532);
nor U20098 (N_20098,N_19568,N_19502);
or U20099 (N_20099,N_19705,N_19530);
xnor U20100 (N_20100,N_19862,N_19551);
or U20101 (N_20101,N_19850,N_19915);
nor U20102 (N_20102,N_19963,N_19560);
and U20103 (N_20103,N_19651,N_19519);
xnor U20104 (N_20104,N_19804,N_19542);
nand U20105 (N_20105,N_19897,N_19819);
or U20106 (N_20106,N_19536,N_19787);
and U20107 (N_20107,N_19950,N_19704);
or U20108 (N_20108,N_19892,N_19764);
xnor U20109 (N_20109,N_19771,N_19737);
xor U20110 (N_20110,N_19999,N_19736);
or U20111 (N_20111,N_19733,N_19883);
nand U20112 (N_20112,N_19911,N_19562);
nor U20113 (N_20113,N_19682,N_19855);
or U20114 (N_20114,N_19822,N_19633);
nor U20115 (N_20115,N_19969,N_19841);
and U20116 (N_20116,N_19817,N_19694);
nor U20117 (N_20117,N_19979,N_19874);
or U20118 (N_20118,N_19655,N_19666);
or U20119 (N_20119,N_19508,N_19782);
nand U20120 (N_20120,N_19656,N_19990);
xnor U20121 (N_20121,N_19599,N_19584);
or U20122 (N_20122,N_19959,N_19631);
nor U20123 (N_20123,N_19988,N_19594);
nand U20124 (N_20124,N_19740,N_19775);
nand U20125 (N_20125,N_19893,N_19623);
or U20126 (N_20126,N_19732,N_19596);
and U20127 (N_20127,N_19854,N_19867);
and U20128 (N_20128,N_19514,N_19769);
and U20129 (N_20129,N_19653,N_19726);
nor U20130 (N_20130,N_19563,N_19518);
xor U20131 (N_20131,N_19597,N_19722);
or U20132 (N_20132,N_19835,N_19781);
or U20133 (N_20133,N_19924,N_19820);
and U20134 (N_20134,N_19708,N_19783);
nor U20135 (N_20135,N_19983,N_19824);
and U20136 (N_20136,N_19938,N_19605);
or U20137 (N_20137,N_19637,N_19802);
xor U20138 (N_20138,N_19741,N_19582);
or U20139 (N_20139,N_19834,N_19642);
and U20140 (N_20140,N_19828,N_19997);
and U20141 (N_20141,N_19665,N_19774);
nor U20142 (N_20142,N_19865,N_19667);
or U20143 (N_20143,N_19880,N_19592);
nor U20144 (N_20144,N_19698,N_19994);
xor U20145 (N_20145,N_19887,N_19766);
nor U20146 (N_20146,N_19618,N_19652);
xnor U20147 (N_20147,N_19829,N_19827);
nor U20148 (N_20148,N_19654,N_19625);
or U20149 (N_20149,N_19688,N_19837);
xnor U20150 (N_20150,N_19575,N_19557);
nor U20151 (N_20151,N_19713,N_19647);
nor U20152 (N_20152,N_19799,N_19657);
or U20153 (N_20153,N_19901,N_19734);
nand U20154 (N_20154,N_19780,N_19952);
or U20155 (N_20155,N_19691,N_19662);
or U20156 (N_20156,N_19663,N_19721);
xnor U20157 (N_20157,N_19801,N_19752);
nand U20158 (N_20158,N_19689,N_19870);
and U20159 (N_20159,N_19830,N_19869);
and U20160 (N_20160,N_19930,N_19606);
or U20161 (N_20161,N_19521,N_19706);
xor U20162 (N_20162,N_19640,N_19695);
or U20163 (N_20163,N_19797,N_19684);
and U20164 (N_20164,N_19707,N_19679);
or U20165 (N_20165,N_19690,N_19628);
xnor U20166 (N_20166,N_19895,N_19971);
nor U20167 (N_20167,N_19967,N_19602);
nand U20168 (N_20168,N_19902,N_19676);
nand U20169 (N_20169,N_19914,N_19614);
nand U20170 (N_20170,N_19561,N_19720);
nand U20171 (N_20171,N_19577,N_19768);
nand U20172 (N_20172,N_19659,N_19644);
nand U20173 (N_20173,N_19507,N_19786);
or U20174 (N_20174,N_19677,N_19671);
xor U20175 (N_20175,N_19622,N_19564);
nor U20176 (N_20176,N_19821,N_19552);
or U20177 (N_20177,N_19872,N_19970);
nor U20178 (N_20178,N_19554,N_19593);
and U20179 (N_20179,N_19941,N_19567);
xor U20180 (N_20180,N_19976,N_19942);
and U20181 (N_20181,N_19524,N_19670);
nor U20182 (N_20182,N_19910,N_19974);
xor U20183 (N_20183,N_19727,N_19544);
or U20184 (N_20184,N_19965,N_19598);
nor U20185 (N_20185,N_19864,N_19559);
or U20186 (N_20186,N_19675,N_19984);
nor U20187 (N_20187,N_19753,N_19589);
or U20188 (N_20188,N_19553,N_19624);
nand U20189 (N_20189,N_19756,N_19985);
or U20190 (N_20190,N_19873,N_19545);
xor U20191 (N_20191,N_19566,N_19810);
nor U20192 (N_20192,N_19550,N_19859);
nand U20193 (N_20193,N_19853,N_19958);
nor U20194 (N_20194,N_19643,N_19534);
or U20195 (N_20195,N_19934,N_19993);
nor U20196 (N_20196,N_19634,N_19538);
nor U20197 (N_20197,N_19716,N_19571);
or U20198 (N_20198,N_19755,N_19699);
and U20199 (N_20199,N_19759,N_19585);
xnor U20200 (N_20200,N_19674,N_19948);
and U20201 (N_20201,N_19876,N_19807);
nor U20202 (N_20202,N_19795,N_19928);
nor U20203 (N_20203,N_19845,N_19882);
or U20204 (N_20204,N_19687,N_19650);
or U20205 (N_20205,N_19920,N_19912);
xor U20206 (N_20206,N_19909,N_19572);
or U20207 (N_20207,N_19501,N_19569);
and U20208 (N_20208,N_19696,N_19541);
nor U20209 (N_20209,N_19917,N_19921);
xor U20210 (N_20210,N_19664,N_19933);
nand U20211 (N_20211,N_19811,N_19668);
and U20212 (N_20212,N_19888,N_19903);
xnor U20213 (N_20213,N_19847,N_19973);
xor U20214 (N_20214,N_19581,N_19660);
nor U20215 (N_20215,N_19608,N_19894);
xor U20216 (N_20216,N_19789,N_19982);
xnor U20217 (N_20217,N_19615,N_19645);
and U20218 (N_20218,N_19833,N_19639);
nand U20219 (N_20219,N_19858,N_19749);
xor U20220 (N_20220,N_19543,N_19743);
nor U20221 (N_20221,N_19685,N_19840);
xor U20222 (N_20222,N_19899,N_19991);
or U20223 (N_20223,N_19547,N_19610);
and U20224 (N_20224,N_19788,N_19805);
and U20225 (N_20225,N_19744,N_19751);
and U20226 (N_20226,N_19529,N_19954);
and U20227 (N_20227,N_19980,N_19549);
nor U20228 (N_20228,N_19527,N_19583);
or U20229 (N_20229,N_19886,N_19505);
nor U20230 (N_20230,N_19703,N_19750);
nand U20231 (N_20231,N_19906,N_19998);
or U20232 (N_20232,N_19574,N_19794);
xor U20233 (N_20233,N_19814,N_19940);
nor U20234 (N_20234,N_19526,N_19962);
nand U20235 (N_20235,N_19927,N_19729);
xnor U20236 (N_20236,N_19836,N_19570);
or U20237 (N_20237,N_19839,N_19946);
and U20238 (N_20238,N_19919,N_19812);
and U20239 (N_20239,N_19765,N_19620);
and U20240 (N_20240,N_19875,N_19591);
and U20241 (N_20241,N_19818,N_19517);
xor U20242 (N_20242,N_19966,N_19626);
xnor U20243 (N_20243,N_19540,N_19528);
nor U20244 (N_20244,N_19604,N_19595);
nand U20245 (N_20245,N_19516,N_19718);
nor U20246 (N_20246,N_19939,N_19779);
xnor U20247 (N_20247,N_19638,N_19929);
nand U20248 (N_20248,N_19621,N_19852);
and U20249 (N_20249,N_19806,N_19923);
nand U20250 (N_20250,N_19523,N_19804);
and U20251 (N_20251,N_19787,N_19743);
and U20252 (N_20252,N_19516,N_19740);
nand U20253 (N_20253,N_19889,N_19990);
or U20254 (N_20254,N_19541,N_19970);
nand U20255 (N_20255,N_19596,N_19779);
nor U20256 (N_20256,N_19989,N_19888);
or U20257 (N_20257,N_19509,N_19590);
xor U20258 (N_20258,N_19807,N_19541);
nand U20259 (N_20259,N_19597,N_19979);
and U20260 (N_20260,N_19546,N_19925);
and U20261 (N_20261,N_19508,N_19753);
and U20262 (N_20262,N_19578,N_19754);
nand U20263 (N_20263,N_19923,N_19607);
xor U20264 (N_20264,N_19787,N_19840);
and U20265 (N_20265,N_19610,N_19626);
or U20266 (N_20266,N_19953,N_19918);
xnor U20267 (N_20267,N_19827,N_19653);
xnor U20268 (N_20268,N_19744,N_19645);
nand U20269 (N_20269,N_19969,N_19903);
xor U20270 (N_20270,N_19779,N_19609);
nand U20271 (N_20271,N_19834,N_19757);
xnor U20272 (N_20272,N_19738,N_19745);
or U20273 (N_20273,N_19626,N_19851);
xnor U20274 (N_20274,N_19870,N_19918);
xor U20275 (N_20275,N_19834,N_19979);
nand U20276 (N_20276,N_19508,N_19867);
xnor U20277 (N_20277,N_19500,N_19995);
nand U20278 (N_20278,N_19932,N_19824);
xnor U20279 (N_20279,N_19625,N_19827);
or U20280 (N_20280,N_19677,N_19840);
nor U20281 (N_20281,N_19995,N_19714);
or U20282 (N_20282,N_19589,N_19805);
or U20283 (N_20283,N_19701,N_19691);
nand U20284 (N_20284,N_19711,N_19892);
and U20285 (N_20285,N_19511,N_19838);
and U20286 (N_20286,N_19895,N_19540);
and U20287 (N_20287,N_19562,N_19923);
and U20288 (N_20288,N_19581,N_19841);
nand U20289 (N_20289,N_19637,N_19614);
nand U20290 (N_20290,N_19721,N_19639);
and U20291 (N_20291,N_19926,N_19614);
nor U20292 (N_20292,N_19672,N_19929);
and U20293 (N_20293,N_19936,N_19671);
and U20294 (N_20294,N_19673,N_19980);
nand U20295 (N_20295,N_19856,N_19710);
nand U20296 (N_20296,N_19916,N_19874);
nand U20297 (N_20297,N_19866,N_19601);
and U20298 (N_20298,N_19792,N_19987);
nor U20299 (N_20299,N_19829,N_19571);
or U20300 (N_20300,N_19898,N_19513);
xor U20301 (N_20301,N_19975,N_19550);
nor U20302 (N_20302,N_19775,N_19715);
nand U20303 (N_20303,N_19914,N_19768);
and U20304 (N_20304,N_19770,N_19542);
and U20305 (N_20305,N_19525,N_19592);
or U20306 (N_20306,N_19974,N_19751);
nand U20307 (N_20307,N_19947,N_19641);
nand U20308 (N_20308,N_19633,N_19785);
nor U20309 (N_20309,N_19562,N_19555);
and U20310 (N_20310,N_19553,N_19646);
nand U20311 (N_20311,N_19958,N_19605);
or U20312 (N_20312,N_19747,N_19624);
and U20313 (N_20313,N_19955,N_19636);
or U20314 (N_20314,N_19896,N_19889);
and U20315 (N_20315,N_19507,N_19813);
and U20316 (N_20316,N_19975,N_19751);
and U20317 (N_20317,N_19853,N_19911);
nor U20318 (N_20318,N_19883,N_19996);
and U20319 (N_20319,N_19679,N_19947);
and U20320 (N_20320,N_19638,N_19938);
and U20321 (N_20321,N_19817,N_19743);
or U20322 (N_20322,N_19613,N_19846);
nand U20323 (N_20323,N_19807,N_19782);
xor U20324 (N_20324,N_19551,N_19678);
nand U20325 (N_20325,N_19688,N_19906);
xor U20326 (N_20326,N_19956,N_19826);
nand U20327 (N_20327,N_19666,N_19711);
nand U20328 (N_20328,N_19822,N_19783);
xnor U20329 (N_20329,N_19798,N_19857);
nand U20330 (N_20330,N_19567,N_19789);
nand U20331 (N_20331,N_19946,N_19762);
or U20332 (N_20332,N_19882,N_19836);
xnor U20333 (N_20333,N_19545,N_19939);
and U20334 (N_20334,N_19692,N_19604);
and U20335 (N_20335,N_19527,N_19980);
nand U20336 (N_20336,N_19874,N_19744);
or U20337 (N_20337,N_19856,N_19920);
xor U20338 (N_20338,N_19707,N_19525);
nor U20339 (N_20339,N_19963,N_19993);
nand U20340 (N_20340,N_19601,N_19690);
and U20341 (N_20341,N_19684,N_19915);
nor U20342 (N_20342,N_19733,N_19594);
and U20343 (N_20343,N_19902,N_19683);
xor U20344 (N_20344,N_19661,N_19960);
or U20345 (N_20345,N_19857,N_19617);
xnor U20346 (N_20346,N_19758,N_19757);
nand U20347 (N_20347,N_19783,N_19592);
xor U20348 (N_20348,N_19567,N_19587);
nor U20349 (N_20349,N_19617,N_19804);
or U20350 (N_20350,N_19618,N_19686);
xnor U20351 (N_20351,N_19838,N_19896);
nand U20352 (N_20352,N_19957,N_19502);
nor U20353 (N_20353,N_19703,N_19682);
nor U20354 (N_20354,N_19644,N_19524);
nand U20355 (N_20355,N_19685,N_19866);
xor U20356 (N_20356,N_19730,N_19537);
nor U20357 (N_20357,N_19831,N_19837);
xnor U20358 (N_20358,N_19520,N_19958);
and U20359 (N_20359,N_19676,N_19888);
nand U20360 (N_20360,N_19597,N_19589);
and U20361 (N_20361,N_19956,N_19791);
or U20362 (N_20362,N_19823,N_19718);
or U20363 (N_20363,N_19758,N_19953);
nand U20364 (N_20364,N_19560,N_19931);
or U20365 (N_20365,N_19866,N_19748);
nand U20366 (N_20366,N_19872,N_19960);
or U20367 (N_20367,N_19858,N_19986);
nor U20368 (N_20368,N_19987,N_19638);
nor U20369 (N_20369,N_19766,N_19636);
nor U20370 (N_20370,N_19762,N_19773);
or U20371 (N_20371,N_19694,N_19811);
or U20372 (N_20372,N_19949,N_19694);
nand U20373 (N_20373,N_19683,N_19969);
nor U20374 (N_20374,N_19815,N_19534);
and U20375 (N_20375,N_19674,N_19708);
and U20376 (N_20376,N_19922,N_19582);
nand U20377 (N_20377,N_19805,N_19900);
or U20378 (N_20378,N_19769,N_19813);
nand U20379 (N_20379,N_19576,N_19986);
xnor U20380 (N_20380,N_19773,N_19643);
nor U20381 (N_20381,N_19820,N_19752);
nand U20382 (N_20382,N_19569,N_19685);
nand U20383 (N_20383,N_19805,N_19978);
xor U20384 (N_20384,N_19635,N_19922);
nor U20385 (N_20385,N_19700,N_19878);
or U20386 (N_20386,N_19731,N_19716);
nor U20387 (N_20387,N_19775,N_19765);
nor U20388 (N_20388,N_19913,N_19593);
or U20389 (N_20389,N_19671,N_19780);
nand U20390 (N_20390,N_19679,N_19977);
xnor U20391 (N_20391,N_19919,N_19567);
nor U20392 (N_20392,N_19973,N_19941);
nand U20393 (N_20393,N_19544,N_19598);
and U20394 (N_20394,N_19657,N_19572);
xor U20395 (N_20395,N_19638,N_19507);
or U20396 (N_20396,N_19511,N_19969);
xor U20397 (N_20397,N_19883,N_19919);
or U20398 (N_20398,N_19943,N_19924);
nand U20399 (N_20399,N_19781,N_19608);
xor U20400 (N_20400,N_19733,N_19937);
or U20401 (N_20401,N_19943,N_19803);
xnor U20402 (N_20402,N_19640,N_19668);
or U20403 (N_20403,N_19519,N_19565);
and U20404 (N_20404,N_19942,N_19818);
and U20405 (N_20405,N_19945,N_19868);
and U20406 (N_20406,N_19789,N_19521);
nand U20407 (N_20407,N_19944,N_19942);
and U20408 (N_20408,N_19821,N_19748);
or U20409 (N_20409,N_19821,N_19840);
nand U20410 (N_20410,N_19573,N_19933);
or U20411 (N_20411,N_19637,N_19968);
nor U20412 (N_20412,N_19680,N_19754);
and U20413 (N_20413,N_19753,N_19905);
and U20414 (N_20414,N_19775,N_19746);
and U20415 (N_20415,N_19954,N_19581);
or U20416 (N_20416,N_19919,N_19699);
nor U20417 (N_20417,N_19759,N_19634);
xor U20418 (N_20418,N_19953,N_19951);
nor U20419 (N_20419,N_19696,N_19726);
nand U20420 (N_20420,N_19849,N_19942);
nand U20421 (N_20421,N_19750,N_19999);
nor U20422 (N_20422,N_19557,N_19882);
or U20423 (N_20423,N_19840,N_19511);
nand U20424 (N_20424,N_19537,N_19865);
or U20425 (N_20425,N_19959,N_19870);
nor U20426 (N_20426,N_19672,N_19610);
or U20427 (N_20427,N_19583,N_19956);
xnor U20428 (N_20428,N_19980,N_19833);
and U20429 (N_20429,N_19716,N_19605);
xor U20430 (N_20430,N_19705,N_19670);
nor U20431 (N_20431,N_19806,N_19972);
xnor U20432 (N_20432,N_19876,N_19742);
and U20433 (N_20433,N_19609,N_19667);
and U20434 (N_20434,N_19869,N_19701);
nand U20435 (N_20435,N_19782,N_19704);
nor U20436 (N_20436,N_19960,N_19603);
nor U20437 (N_20437,N_19609,N_19807);
xor U20438 (N_20438,N_19900,N_19720);
nor U20439 (N_20439,N_19604,N_19981);
nand U20440 (N_20440,N_19593,N_19826);
and U20441 (N_20441,N_19940,N_19671);
and U20442 (N_20442,N_19777,N_19981);
and U20443 (N_20443,N_19933,N_19976);
xnor U20444 (N_20444,N_19854,N_19959);
nor U20445 (N_20445,N_19515,N_19798);
and U20446 (N_20446,N_19924,N_19743);
or U20447 (N_20447,N_19982,N_19543);
nor U20448 (N_20448,N_19908,N_19952);
nand U20449 (N_20449,N_19822,N_19839);
nand U20450 (N_20450,N_19826,N_19854);
nand U20451 (N_20451,N_19997,N_19635);
xor U20452 (N_20452,N_19908,N_19560);
and U20453 (N_20453,N_19548,N_19631);
and U20454 (N_20454,N_19728,N_19520);
nor U20455 (N_20455,N_19666,N_19733);
and U20456 (N_20456,N_19959,N_19581);
nor U20457 (N_20457,N_19963,N_19703);
nor U20458 (N_20458,N_19940,N_19685);
xnor U20459 (N_20459,N_19828,N_19804);
or U20460 (N_20460,N_19750,N_19570);
or U20461 (N_20461,N_19725,N_19897);
or U20462 (N_20462,N_19606,N_19665);
or U20463 (N_20463,N_19858,N_19569);
or U20464 (N_20464,N_19663,N_19801);
nand U20465 (N_20465,N_19768,N_19643);
and U20466 (N_20466,N_19984,N_19804);
or U20467 (N_20467,N_19919,N_19799);
nand U20468 (N_20468,N_19695,N_19869);
or U20469 (N_20469,N_19978,N_19847);
or U20470 (N_20470,N_19965,N_19751);
or U20471 (N_20471,N_19999,N_19764);
nor U20472 (N_20472,N_19802,N_19815);
nor U20473 (N_20473,N_19525,N_19554);
nand U20474 (N_20474,N_19798,N_19555);
or U20475 (N_20475,N_19514,N_19855);
nor U20476 (N_20476,N_19651,N_19663);
and U20477 (N_20477,N_19578,N_19987);
nor U20478 (N_20478,N_19696,N_19995);
nor U20479 (N_20479,N_19673,N_19923);
and U20480 (N_20480,N_19730,N_19887);
nand U20481 (N_20481,N_19612,N_19807);
nor U20482 (N_20482,N_19661,N_19507);
and U20483 (N_20483,N_19894,N_19679);
xnor U20484 (N_20484,N_19747,N_19891);
or U20485 (N_20485,N_19686,N_19865);
or U20486 (N_20486,N_19577,N_19956);
nand U20487 (N_20487,N_19994,N_19586);
or U20488 (N_20488,N_19732,N_19542);
and U20489 (N_20489,N_19512,N_19766);
xor U20490 (N_20490,N_19808,N_19807);
and U20491 (N_20491,N_19836,N_19707);
xnor U20492 (N_20492,N_19995,N_19510);
nand U20493 (N_20493,N_19899,N_19742);
xnor U20494 (N_20494,N_19590,N_19846);
nor U20495 (N_20495,N_19941,N_19625);
xnor U20496 (N_20496,N_19955,N_19676);
nor U20497 (N_20497,N_19921,N_19817);
and U20498 (N_20498,N_19596,N_19767);
or U20499 (N_20499,N_19815,N_19687);
xnor U20500 (N_20500,N_20214,N_20055);
nor U20501 (N_20501,N_20353,N_20082);
and U20502 (N_20502,N_20089,N_20039);
xor U20503 (N_20503,N_20139,N_20418);
nand U20504 (N_20504,N_20152,N_20229);
nand U20505 (N_20505,N_20157,N_20330);
xor U20506 (N_20506,N_20107,N_20026);
and U20507 (N_20507,N_20452,N_20344);
nor U20508 (N_20508,N_20073,N_20154);
or U20509 (N_20509,N_20168,N_20226);
nor U20510 (N_20510,N_20274,N_20318);
or U20511 (N_20511,N_20467,N_20027);
or U20512 (N_20512,N_20036,N_20394);
or U20513 (N_20513,N_20132,N_20174);
and U20514 (N_20514,N_20429,N_20448);
nor U20515 (N_20515,N_20205,N_20077);
xnor U20516 (N_20516,N_20068,N_20075);
and U20517 (N_20517,N_20167,N_20419);
xnor U20518 (N_20518,N_20001,N_20314);
and U20519 (N_20519,N_20123,N_20013);
nor U20520 (N_20520,N_20308,N_20494);
nand U20521 (N_20521,N_20170,N_20297);
or U20522 (N_20522,N_20112,N_20334);
xor U20523 (N_20523,N_20118,N_20322);
nor U20524 (N_20524,N_20413,N_20285);
nor U20525 (N_20525,N_20440,N_20213);
nand U20526 (N_20526,N_20007,N_20052);
or U20527 (N_20527,N_20309,N_20053);
nor U20528 (N_20528,N_20067,N_20304);
nand U20529 (N_20529,N_20141,N_20146);
nor U20530 (N_20530,N_20142,N_20444);
nand U20531 (N_20531,N_20499,N_20283);
nor U20532 (N_20532,N_20269,N_20338);
xor U20533 (N_20533,N_20371,N_20130);
and U20534 (N_20534,N_20465,N_20387);
nor U20535 (N_20535,N_20177,N_20323);
xor U20536 (N_20536,N_20015,N_20165);
xor U20537 (N_20537,N_20171,N_20201);
nor U20538 (N_20538,N_20151,N_20085);
xnor U20539 (N_20539,N_20405,N_20311);
xor U20540 (N_20540,N_20328,N_20219);
xor U20541 (N_20541,N_20277,N_20349);
nand U20542 (N_20542,N_20270,N_20094);
and U20543 (N_20543,N_20292,N_20096);
nand U20544 (N_20544,N_20182,N_20124);
and U20545 (N_20545,N_20497,N_20351);
nor U20546 (N_20546,N_20233,N_20479);
nor U20547 (N_20547,N_20066,N_20296);
nand U20548 (N_20548,N_20261,N_20163);
nand U20549 (N_20549,N_20207,N_20358);
xnor U20550 (N_20550,N_20372,N_20000);
nand U20551 (N_20551,N_20332,N_20251);
nor U20552 (N_20552,N_20042,N_20291);
xnor U20553 (N_20553,N_20469,N_20202);
or U20554 (N_20554,N_20008,N_20169);
nand U20555 (N_20555,N_20020,N_20212);
and U20556 (N_20556,N_20102,N_20050);
xor U20557 (N_20557,N_20136,N_20453);
or U20558 (N_20558,N_20069,N_20295);
nand U20559 (N_20559,N_20149,N_20159);
and U20560 (N_20560,N_20040,N_20282);
or U20561 (N_20561,N_20215,N_20091);
xor U20562 (N_20562,N_20006,N_20129);
xor U20563 (N_20563,N_20327,N_20442);
nand U20564 (N_20564,N_20478,N_20048);
xnor U20565 (N_20565,N_20148,N_20342);
xor U20566 (N_20566,N_20254,N_20051);
nand U20567 (N_20567,N_20428,N_20389);
and U20568 (N_20568,N_20003,N_20238);
nand U20569 (N_20569,N_20115,N_20074);
nand U20570 (N_20570,N_20305,N_20211);
or U20571 (N_20571,N_20087,N_20128);
and U20572 (N_20572,N_20218,N_20266);
xor U20573 (N_20573,N_20301,N_20280);
and U20574 (N_20574,N_20360,N_20045);
nand U20575 (N_20575,N_20432,N_20464);
nor U20576 (N_20576,N_20268,N_20242);
nor U20577 (N_20577,N_20273,N_20176);
or U20578 (N_20578,N_20293,N_20443);
and U20579 (N_20579,N_20310,N_20400);
xnor U20580 (N_20580,N_20247,N_20289);
or U20581 (N_20581,N_20359,N_20320);
xor U20582 (N_20582,N_20175,N_20433);
or U20583 (N_20583,N_20184,N_20290);
or U20584 (N_20584,N_20350,N_20143);
nor U20585 (N_20585,N_20046,N_20031);
nand U20586 (N_20586,N_20376,N_20030);
and U20587 (N_20587,N_20461,N_20117);
nand U20588 (N_20588,N_20252,N_20120);
xor U20589 (N_20589,N_20487,N_20185);
xnor U20590 (N_20590,N_20411,N_20361);
xor U20591 (N_20591,N_20454,N_20057);
and U20592 (N_20592,N_20475,N_20485);
and U20593 (N_20593,N_20455,N_20206);
nor U20594 (N_20594,N_20262,N_20106);
xor U20595 (N_20595,N_20179,N_20147);
nor U20596 (N_20596,N_20223,N_20125);
and U20597 (N_20597,N_20186,N_20278);
nand U20598 (N_20598,N_20072,N_20017);
nor U20599 (N_20599,N_20383,N_20284);
xor U20600 (N_20600,N_20401,N_20476);
or U20601 (N_20601,N_20249,N_20380);
and U20602 (N_20602,N_20257,N_20299);
or U20603 (N_20603,N_20386,N_20445);
nand U20604 (N_20604,N_20144,N_20495);
and U20605 (N_20605,N_20220,N_20191);
xnor U20606 (N_20606,N_20166,N_20347);
and U20607 (N_20607,N_20098,N_20435);
and U20608 (N_20608,N_20420,N_20390);
xor U20609 (N_20609,N_20246,N_20023);
nor U20610 (N_20610,N_20183,N_20321);
or U20611 (N_20611,N_20391,N_20434);
nand U20612 (N_20612,N_20195,N_20329);
and U20613 (N_20613,N_20355,N_20181);
nor U20614 (N_20614,N_20488,N_20234);
xor U20615 (N_20615,N_20034,N_20402);
nor U20616 (N_20616,N_20192,N_20150);
and U20617 (N_20617,N_20399,N_20496);
and U20618 (N_20618,N_20111,N_20172);
or U20619 (N_20619,N_20339,N_20189);
nand U20620 (N_20620,N_20037,N_20019);
nor U20621 (N_20621,N_20180,N_20025);
nand U20622 (N_20622,N_20070,N_20362);
xnor U20623 (N_20623,N_20375,N_20236);
nor U20624 (N_20624,N_20054,N_20307);
and U20625 (N_20625,N_20121,N_20244);
nor U20626 (N_20626,N_20024,N_20188);
nor U20627 (N_20627,N_20281,N_20325);
xnor U20628 (N_20628,N_20256,N_20288);
nor U20629 (N_20629,N_20286,N_20462);
nand U20630 (N_20630,N_20114,N_20460);
nand U20631 (N_20631,N_20199,N_20248);
and U20632 (N_20632,N_20490,N_20367);
nand U20633 (N_20633,N_20103,N_20187);
and U20634 (N_20634,N_20081,N_20265);
and U20635 (N_20635,N_20415,N_20374);
xor U20636 (N_20636,N_20193,N_20313);
or U20637 (N_20637,N_20416,N_20065);
xnor U20638 (N_20638,N_20457,N_20047);
nor U20639 (N_20639,N_20385,N_20439);
and U20640 (N_20640,N_20241,N_20404);
xnor U20641 (N_20641,N_20231,N_20135);
nor U20642 (N_20642,N_20459,N_20451);
xnor U20643 (N_20643,N_20090,N_20426);
or U20644 (N_20644,N_20255,N_20368);
and U20645 (N_20645,N_20410,N_20263);
or U20646 (N_20646,N_20450,N_20064);
nand U20647 (N_20647,N_20011,N_20486);
nand U20648 (N_20648,N_20110,N_20108);
or U20649 (N_20649,N_20002,N_20472);
or U20650 (N_20650,N_20210,N_20092);
nand U20651 (N_20651,N_20080,N_20382);
xor U20652 (N_20652,N_20131,N_20153);
nand U20653 (N_20653,N_20044,N_20437);
xnor U20654 (N_20654,N_20458,N_20196);
and U20655 (N_20655,N_20498,N_20204);
and U20656 (N_20656,N_20431,N_20474);
xnor U20657 (N_20657,N_20369,N_20378);
or U20658 (N_20658,N_20446,N_20018);
or U20659 (N_20659,N_20060,N_20071);
or U20660 (N_20660,N_20312,N_20161);
and U20661 (N_20661,N_20333,N_20224);
or U20662 (N_20662,N_20403,N_20119);
nor U20663 (N_20663,N_20470,N_20164);
xnor U20664 (N_20664,N_20354,N_20370);
xor U20665 (N_20665,N_20477,N_20449);
nand U20666 (N_20666,N_20331,N_20253);
xor U20667 (N_20667,N_20237,N_20221);
nor U20668 (N_20668,N_20337,N_20137);
and U20669 (N_20669,N_20414,N_20095);
xor U20670 (N_20670,N_20272,N_20029);
xor U20671 (N_20671,N_20463,N_20340);
and U20672 (N_20672,N_20438,N_20287);
nand U20673 (N_20673,N_20260,N_20471);
and U20674 (N_20674,N_20373,N_20028);
nand U20675 (N_20675,N_20088,N_20227);
nor U20676 (N_20676,N_20162,N_20468);
nor U20677 (N_20677,N_20352,N_20489);
xnor U20678 (N_20678,N_20436,N_20127);
nand U20679 (N_20679,N_20407,N_20365);
and U20680 (N_20680,N_20294,N_20232);
and U20681 (N_20681,N_20134,N_20208);
nor U20682 (N_20682,N_20319,N_20412);
and U20683 (N_20683,N_20480,N_20492);
or U20684 (N_20684,N_20259,N_20493);
nand U20685 (N_20685,N_20086,N_20379);
nor U20686 (N_20686,N_20225,N_20363);
or U20687 (N_20687,N_20104,N_20335);
or U20688 (N_20688,N_20217,N_20364);
nand U20689 (N_20689,N_20158,N_20316);
or U20690 (N_20690,N_20194,N_20447);
nand U20691 (N_20691,N_20456,N_20388);
nand U20692 (N_20692,N_20156,N_20357);
nand U20693 (N_20693,N_20406,N_20398);
nor U20694 (N_20694,N_20366,N_20076);
and U20695 (N_20695,N_20105,N_20133);
nor U20696 (N_20696,N_20491,N_20424);
xnor U20697 (N_20697,N_20009,N_20343);
xnor U20698 (N_20698,N_20303,N_20138);
nand U20699 (N_20699,N_20056,N_20063);
nor U20700 (N_20700,N_20228,N_20271);
nor U20701 (N_20701,N_20300,N_20209);
nand U20702 (N_20702,N_20356,N_20155);
and U20703 (N_20703,N_20083,N_20381);
xnor U20704 (N_20704,N_20005,N_20062);
xnor U20705 (N_20705,N_20021,N_20061);
nand U20706 (N_20706,N_20317,N_20484);
xnor U20707 (N_20707,N_20466,N_20481);
nand U20708 (N_20708,N_20482,N_20409);
nor U20709 (N_20709,N_20267,N_20396);
xnor U20710 (N_20710,N_20345,N_20324);
xnor U20711 (N_20711,N_20230,N_20016);
xnor U20712 (N_20712,N_20203,N_20239);
or U20713 (N_20713,N_20441,N_20035);
xor U20714 (N_20714,N_20377,N_20058);
xor U20715 (N_20715,N_20427,N_20041);
or U20716 (N_20716,N_20145,N_20043);
nand U20717 (N_20717,N_20395,N_20099);
xor U20718 (N_20718,N_20084,N_20264);
xor U20719 (N_20719,N_20078,N_20032);
nand U20720 (N_20720,N_20341,N_20392);
and U20721 (N_20721,N_20250,N_20302);
and U20722 (N_20722,N_20004,N_20306);
xor U20723 (N_20723,N_20116,N_20038);
and U20724 (N_20724,N_20101,N_20417);
or U20725 (N_20725,N_20198,N_20097);
nand U20726 (N_20726,N_20245,N_20276);
nor U20727 (N_20727,N_20059,N_20079);
xnor U20728 (N_20728,N_20178,N_20222);
xnor U20729 (N_20729,N_20010,N_20421);
and U20730 (N_20730,N_20190,N_20258);
xnor U20731 (N_20731,N_20012,N_20408);
xor U20732 (N_20732,N_20423,N_20326);
and U20733 (N_20733,N_20393,N_20033);
nand U20734 (N_20734,N_20275,N_20315);
nor U20735 (N_20735,N_20346,N_20298);
nand U20736 (N_20736,N_20235,N_20160);
xnor U20737 (N_20737,N_20243,N_20422);
nor U20738 (N_20738,N_20430,N_20483);
or U20739 (N_20739,N_20240,N_20022);
and U20740 (N_20740,N_20279,N_20126);
nor U20741 (N_20741,N_20100,N_20140);
nor U20742 (N_20742,N_20473,N_20093);
or U20743 (N_20743,N_20122,N_20425);
xor U20744 (N_20744,N_20049,N_20216);
nor U20745 (N_20745,N_20173,N_20197);
and U20746 (N_20746,N_20336,N_20113);
or U20747 (N_20747,N_20200,N_20384);
nand U20748 (N_20748,N_20348,N_20109);
xor U20749 (N_20749,N_20014,N_20397);
nor U20750 (N_20750,N_20479,N_20392);
xnor U20751 (N_20751,N_20231,N_20090);
nand U20752 (N_20752,N_20396,N_20000);
nor U20753 (N_20753,N_20008,N_20114);
and U20754 (N_20754,N_20376,N_20177);
nor U20755 (N_20755,N_20219,N_20435);
or U20756 (N_20756,N_20143,N_20100);
nand U20757 (N_20757,N_20460,N_20250);
and U20758 (N_20758,N_20275,N_20010);
nor U20759 (N_20759,N_20299,N_20397);
and U20760 (N_20760,N_20095,N_20083);
nor U20761 (N_20761,N_20487,N_20154);
xnor U20762 (N_20762,N_20471,N_20139);
or U20763 (N_20763,N_20179,N_20477);
nor U20764 (N_20764,N_20478,N_20357);
and U20765 (N_20765,N_20050,N_20326);
nor U20766 (N_20766,N_20170,N_20211);
nand U20767 (N_20767,N_20377,N_20341);
nand U20768 (N_20768,N_20123,N_20482);
nand U20769 (N_20769,N_20352,N_20432);
and U20770 (N_20770,N_20478,N_20209);
nand U20771 (N_20771,N_20132,N_20079);
and U20772 (N_20772,N_20189,N_20259);
xnor U20773 (N_20773,N_20174,N_20016);
or U20774 (N_20774,N_20451,N_20291);
and U20775 (N_20775,N_20076,N_20246);
xnor U20776 (N_20776,N_20136,N_20295);
and U20777 (N_20777,N_20329,N_20234);
or U20778 (N_20778,N_20345,N_20416);
and U20779 (N_20779,N_20352,N_20053);
nor U20780 (N_20780,N_20043,N_20364);
or U20781 (N_20781,N_20205,N_20357);
nand U20782 (N_20782,N_20396,N_20188);
or U20783 (N_20783,N_20133,N_20104);
and U20784 (N_20784,N_20220,N_20209);
xnor U20785 (N_20785,N_20119,N_20122);
xnor U20786 (N_20786,N_20290,N_20380);
nor U20787 (N_20787,N_20201,N_20479);
nor U20788 (N_20788,N_20360,N_20006);
and U20789 (N_20789,N_20486,N_20479);
and U20790 (N_20790,N_20116,N_20414);
or U20791 (N_20791,N_20262,N_20309);
xor U20792 (N_20792,N_20143,N_20113);
xnor U20793 (N_20793,N_20266,N_20430);
xor U20794 (N_20794,N_20368,N_20165);
nand U20795 (N_20795,N_20313,N_20221);
nor U20796 (N_20796,N_20458,N_20129);
xnor U20797 (N_20797,N_20105,N_20318);
nand U20798 (N_20798,N_20285,N_20083);
nand U20799 (N_20799,N_20202,N_20203);
or U20800 (N_20800,N_20272,N_20088);
nand U20801 (N_20801,N_20426,N_20268);
nand U20802 (N_20802,N_20181,N_20212);
nand U20803 (N_20803,N_20184,N_20468);
and U20804 (N_20804,N_20371,N_20425);
or U20805 (N_20805,N_20469,N_20413);
nand U20806 (N_20806,N_20259,N_20478);
and U20807 (N_20807,N_20251,N_20378);
nand U20808 (N_20808,N_20419,N_20123);
nand U20809 (N_20809,N_20076,N_20024);
xnor U20810 (N_20810,N_20444,N_20474);
nand U20811 (N_20811,N_20034,N_20128);
xor U20812 (N_20812,N_20466,N_20317);
and U20813 (N_20813,N_20024,N_20411);
or U20814 (N_20814,N_20112,N_20224);
or U20815 (N_20815,N_20315,N_20299);
nand U20816 (N_20816,N_20238,N_20080);
nor U20817 (N_20817,N_20401,N_20186);
nand U20818 (N_20818,N_20251,N_20142);
or U20819 (N_20819,N_20463,N_20401);
xor U20820 (N_20820,N_20420,N_20188);
xor U20821 (N_20821,N_20239,N_20050);
nor U20822 (N_20822,N_20425,N_20402);
nand U20823 (N_20823,N_20302,N_20403);
or U20824 (N_20824,N_20395,N_20420);
nand U20825 (N_20825,N_20316,N_20425);
nand U20826 (N_20826,N_20093,N_20490);
xor U20827 (N_20827,N_20103,N_20202);
and U20828 (N_20828,N_20332,N_20377);
and U20829 (N_20829,N_20358,N_20222);
and U20830 (N_20830,N_20297,N_20084);
nand U20831 (N_20831,N_20152,N_20158);
nand U20832 (N_20832,N_20350,N_20056);
nand U20833 (N_20833,N_20371,N_20307);
nor U20834 (N_20834,N_20358,N_20120);
and U20835 (N_20835,N_20402,N_20102);
or U20836 (N_20836,N_20060,N_20491);
nor U20837 (N_20837,N_20409,N_20437);
xnor U20838 (N_20838,N_20370,N_20424);
and U20839 (N_20839,N_20084,N_20415);
nand U20840 (N_20840,N_20424,N_20104);
and U20841 (N_20841,N_20423,N_20059);
and U20842 (N_20842,N_20213,N_20447);
xnor U20843 (N_20843,N_20472,N_20068);
nor U20844 (N_20844,N_20019,N_20245);
nand U20845 (N_20845,N_20260,N_20313);
or U20846 (N_20846,N_20247,N_20358);
xnor U20847 (N_20847,N_20429,N_20483);
or U20848 (N_20848,N_20216,N_20274);
or U20849 (N_20849,N_20011,N_20221);
or U20850 (N_20850,N_20016,N_20200);
and U20851 (N_20851,N_20169,N_20308);
or U20852 (N_20852,N_20349,N_20034);
nor U20853 (N_20853,N_20435,N_20097);
or U20854 (N_20854,N_20405,N_20252);
and U20855 (N_20855,N_20450,N_20239);
nand U20856 (N_20856,N_20377,N_20195);
nor U20857 (N_20857,N_20067,N_20305);
or U20858 (N_20858,N_20499,N_20088);
or U20859 (N_20859,N_20294,N_20283);
or U20860 (N_20860,N_20408,N_20441);
or U20861 (N_20861,N_20230,N_20049);
nand U20862 (N_20862,N_20075,N_20423);
nor U20863 (N_20863,N_20469,N_20393);
xnor U20864 (N_20864,N_20014,N_20069);
nor U20865 (N_20865,N_20212,N_20277);
or U20866 (N_20866,N_20166,N_20003);
and U20867 (N_20867,N_20286,N_20272);
xnor U20868 (N_20868,N_20271,N_20182);
or U20869 (N_20869,N_20087,N_20392);
nand U20870 (N_20870,N_20217,N_20473);
nor U20871 (N_20871,N_20351,N_20350);
nor U20872 (N_20872,N_20468,N_20377);
and U20873 (N_20873,N_20021,N_20250);
and U20874 (N_20874,N_20302,N_20404);
xnor U20875 (N_20875,N_20498,N_20133);
nand U20876 (N_20876,N_20422,N_20330);
xor U20877 (N_20877,N_20462,N_20095);
xor U20878 (N_20878,N_20406,N_20216);
and U20879 (N_20879,N_20035,N_20437);
or U20880 (N_20880,N_20149,N_20392);
xnor U20881 (N_20881,N_20347,N_20321);
nand U20882 (N_20882,N_20495,N_20157);
nand U20883 (N_20883,N_20307,N_20275);
xor U20884 (N_20884,N_20339,N_20292);
and U20885 (N_20885,N_20410,N_20193);
xor U20886 (N_20886,N_20480,N_20328);
nor U20887 (N_20887,N_20458,N_20011);
nand U20888 (N_20888,N_20112,N_20369);
nand U20889 (N_20889,N_20435,N_20049);
and U20890 (N_20890,N_20451,N_20362);
xnor U20891 (N_20891,N_20335,N_20122);
or U20892 (N_20892,N_20160,N_20289);
xnor U20893 (N_20893,N_20482,N_20324);
nor U20894 (N_20894,N_20449,N_20471);
or U20895 (N_20895,N_20024,N_20470);
nor U20896 (N_20896,N_20132,N_20186);
xor U20897 (N_20897,N_20010,N_20216);
nand U20898 (N_20898,N_20329,N_20452);
nand U20899 (N_20899,N_20357,N_20264);
xor U20900 (N_20900,N_20030,N_20171);
nand U20901 (N_20901,N_20097,N_20020);
or U20902 (N_20902,N_20329,N_20231);
nor U20903 (N_20903,N_20057,N_20480);
nand U20904 (N_20904,N_20397,N_20278);
nand U20905 (N_20905,N_20363,N_20181);
or U20906 (N_20906,N_20442,N_20260);
nand U20907 (N_20907,N_20240,N_20387);
or U20908 (N_20908,N_20437,N_20119);
nor U20909 (N_20909,N_20064,N_20045);
nor U20910 (N_20910,N_20055,N_20130);
or U20911 (N_20911,N_20343,N_20392);
and U20912 (N_20912,N_20495,N_20493);
xnor U20913 (N_20913,N_20176,N_20333);
xor U20914 (N_20914,N_20038,N_20487);
nor U20915 (N_20915,N_20358,N_20405);
nand U20916 (N_20916,N_20405,N_20157);
xor U20917 (N_20917,N_20240,N_20282);
xor U20918 (N_20918,N_20056,N_20001);
nor U20919 (N_20919,N_20119,N_20112);
nor U20920 (N_20920,N_20298,N_20252);
nor U20921 (N_20921,N_20269,N_20034);
xnor U20922 (N_20922,N_20086,N_20242);
or U20923 (N_20923,N_20349,N_20292);
or U20924 (N_20924,N_20369,N_20340);
and U20925 (N_20925,N_20351,N_20444);
xnor U20926 (N_20926,N_20152,N_20401);
and U20927 (N_20927,N_20204,N_20184);
and U20928 (N_20928,N_20012,N_20398);
or U20929 (N_20929,N_20497,N_20205);
nor U20930 (N_20930,N_20120,N_20442);
xor U20931 (N_20931,N_20146,N_20464);
nor U20932 (N_20932,N_20099,N_20468);
or U20933 (N_20933,N_20031,N_20371);
and U20934 (N_20934,N_20250,N_20402);
nor U20935 (N_20935,N_20185,N_20145);
or U20936 (N_20936,N_20186,N_20017);
and U20937 (N_20937,N_20176,N_20217);
or U20938 (N_20938,N_20021,N_20107);
and U20939 (N_20939,N_20095,N_20379);
and U20940 (N_20940,N_20402,N_20192);
nor U20941 (N_20941,N_20389,N_20117);
nand U20942 (N_20942,N_20212,N_20017);
xnor U20943 (N_20943,N_20114,N_20083);
or U20944 (N_20944,N_20090,N_20050);
nor U20945 (N_20945,N_20136,N_20430);
nand U20946 (N_20946,N_20483,N_20172);
and U20947 (N_20947,N_20456,N_20046);
or U20948 (N_20948,N_20423,N_20462);
or U20949 (N_20949,N_20184,N_20106);
nand U20950 (N_20950,N_20083,N_20347);
nor U20951 (N_20951,N_20218,N_20061);
or U20952 (N_20952,N_20252,N_20009);
nor U20953 (N_20953,N_20274,N_20033);
nor U20954 (N_20954,N_20441,N_20060);
nor U20955 (N_20955,N_20492,N_20001);
nor U20956 (N_20956,N_20346,N_20437);
or U20957 (N_20957,N_20015,N_20335);
or U20958 (N_20958,N_20304,N_20359);
or U20959 (N_20959,N_20342,N_20191);
and U20960 (N_20960,N_20488,N_20106);
xnor U20961 (N_20961,N_20421,N_20134);
and U20962 (N_20962,N_20092,N_20137);
and U20963 (N_20963,N_20272,N_20256);
or U20964 (N_20964,N_20213,N_20394);
xnor U20965 (N_20965,N_20259,N_20204);
and U20966 (N_20966,N_20236,N_20006);
nand U20967 (N_20967,N_20148,N_20343);
and U20968 (N_20968,N_20208,N_20423);
xnor U20969 (N_20969,N_20466,N_20161);
and U20970 (N_20970,N_20431,N_20441);
nor U20971 (N_20971,N_20446,N_20030);
and U20972 (N_20972,N_20176,N_20170);
nand U20973 (N_20973,N_20274,N_20262);
nand U20974 (N_20974,N_20357,N_20473);
nor U20975 (N_20975,N_20229,N_20082);
and U20976 (N_20976,N_20415,N_20273);
nand U20977 (N_20977,N_20057,N_20018);
nand U20978 (N_20978,N_20337,N_20028);
nand U20979 (N_20979,N_20388,N_20016);
nor U20980 (N_20980,N_20156,N_20178);
nand U20981 (N_20981,N_20262,N_20137);
and U20982 (N_20982,N_20258,N_20421);
xor U20983 (N_20983,N_20226,N_20338);
xor U20984 (N_20984,N_20415,N_20363);
and U20985 (N_20985,N_20087,N_20138);
nor U20986 (N_20986,N_20421,N_20268);
xnor U20987 (N_20987,N_20464,N_20317);
nor U20988 (N_20988,N_20194,N_20218);
nor U20989 (N_20989,N_20386,N_20376);
or U20990 (N_20990,N_20403,N_20453);
nand U20991 (N_20991,N_20297,N_20446);
and U20992 (N_20992,N_20246,N_20397);
nor U20993 (N_20993,N_20246,N_20445);
nor U20994 (N_20994,N_20065,N_20220);
nand U20995 (N_20995,N_20401,N_20096);
nor U20996 (N_20996,N_20178,N_20028);
nor U20997 (N_20997,N_20461,N_20357);
nand U20998 (N_20998,N_20200,N_20086);
or U20999 (N_20999,N_20191,N_20479);
nor U21000 (N_21000,N_20560,N_20880);
nand U21001 (N_21001,N_20850,N_20636);
xnor U21002 (N_21002,N_20816,N_20710);
xor U21003 (N_21003,N_20901,N_20932);
and U21004 (N_21004,N_20762,N_20944);
nor U21005 (N_21005,N_20564,N_20565);
nor U21006 (N_21006,N_20555,N_20703);
nand U21007 (N_21007,N_20732,N_20735);
and U21008 (N_21008,N_20609,N_20958);
nor U21009 (N_21009,N_20552,N_20993);
nor U21010 (N_21010,N_20844,N_20787);
nor U21011 (N_21011,N_20695,N_20957);
and U21012 (N_21012,N_20667,N_20856);
nand U21013 (N_21013,N_20991,N_20502);
nor U21014 (N_21014,N_20683,N_20939);
or U21015 (N_21015,N_20650,N_20888);
or U21016 (N_21016,N_20890,N_20677);
or U21017 (N_21017,N_20734,N_20883);
nand U21018 (N_21018,N_20862,N_20923);
or U21019 (N_21019,N_20898,N_20847);
nand U21020 (N_21020,N_20928,N_20934);
xnor U21021 (N_21021,N_20573,N_20871);
or U21022 (N_21022,N_20861,N_20521);
or U21023 (N_21023,N_20809,N_20680);
nand U21024 (N_21024,N_20532,N_20828);
xor U21025 (N_21025,N_20902,N_20661);
or U21026 (N_21026,N_20924,N_20571);
or U21027 (N_21027,N_20618,N_20972);
or U21028 (N_21028,N_20853,N_20772);
nand U21029 (N_21029,N_20500,N_20831);
xor U21030 (N_21030,N_20791,N_20886);
xnor U21031 (N_21031,N_20654,N_20637);
and U21032 (N_21032,N_20812,N_20725);
or U21033 (N_21033,N_20910,N_20549);
nand U21034 (N_21034,N_20887,N_20520);
and U21035 (N_21035,N_20839,N_20742);
or U21036 (N_21036,N_20501,N_20929);
or U21037 (N_21037,N_20822,N_20523);
nand U21038 (N_21038,N_20505,N_20785);
or U21039 (N_21039,N_20952,N_20859);
nand U21040 (N_21040,N_20651,N_20863);
or U21041 (N_21041,N_20876,N_20986);
and U21042 (N_21042,N_20955,N_20867);
or U21043 (N_21043,N_20835,N_20987);
nor U21044 (N_21044,N_20529,N_20534);
xor U21045 (N_21045,N_20558,N_20761);
and U21046 (N_21046,N_20796,N_20753);
and U21047 (N_21047,N_20894,N_20919);
nand U21048 (N_21048,N_20884,N_20801);
and U21049 (N_21049,N_20586,N_20595);
xor U21050 (N_21050,N_20702,N_20855);
and U21051 (N_21051,N_20617,N_20656);
nor U21052 (N_21052,N_20716,N_20748);
nor U21053 (N_21053,N_20941,N_20613);
nor U21054 (N_21054,N_20629,N_20782);
nor U21055 (N_21055,N_20525,N_20969);
nand U21056 (N_21056,N_20692,N_20547);
and U21057 (N_21057,N_20877,N_20663);
nand U21058 (N_21058,N_20569,N_20764);
nand U21059 (N_21059,N_20626,N_20604);
nor U21060 (N_21060,N_20795,N_20786);
or U21061 (N_21061,N_20630,N_20930);
and U21062 (N_21062,N_20503,N_20580);
nand U21063 (N_21063,N_20897,N_20597);
xnor U21064 (N_21064,N_20974,N_20953);
or U21065 (N_21065,N_20945,N_20647);
nor U21066 (N_21066,N_20829,N_20633);
nand U21067 (N_21067,N_20625,N_20802);
and U21068 (N_21068,N_20992,N_20908);
and U21069 (N_21069,N_20538,N_20895);
xor U21070 (N_21070,N_20550,N_20904);
or U21071 (N_21071,N_20653,N_20673);
nand U21072 (N_21072,N_20510,N_20834);
or U21073 (N_21073,N_20838,N_20504);
and U21074 (N_21074,N_20907,N_20607);
nor U21075 (N_21075,N_20589,N_20775);
or U21076 (N_21076,N_20804,N_20817);
and U21077 (N_21077,N_20705,N_20708);
xnor U21078 (N_21078,N_20837,N_20783);
nand U21079 (N_21079,N_20964,N_20836);
and U21080 (N_21080,N_20864,N_20798);
and U21081 (N_21081,N_20925,N_20612);
and U21082 (N_21082,N_20587,N_20697);
xor U21083 (N_21083,N_20514,N_20519);
or U21084 (N_21084,N_20590,N_20594);
or U21085 (N_21085,N_20541,N_20687);
xor U21086 (N_21086,N_20691,N_20781);
nor U21087 (N_21087,N_20956,N_20686);
xnor U21088 (N_21088,N_20778,N_20631);
and U21089 (N_21089,N_20739,N_20843);
nand U21090 (N_21090,N_20540,N_20535);
nand U21091 (N_21091,N_20803,N_20711);
xnor U21092 (N_21092,N_20615,N_20982);
and U21093 (N_21093,N_20996,N_20757);
or U21094 (N_21094,N_20507,N_20873);
nor U21095 (N_21095,N_20881,N_20526);
nand U21096 (N_21096,N_20750,N_20766);
xor U21097 (N_21097,N_20582,N_20852);
nor U21098 (N_21098,N_20811,N_20818);
and U21099 (N_21099,N_20726,N_20967);
nor U21100 (N_21100,N_20522,N_20690);
xor U21101 (N_21101,N_20506,N_20537);
xor U21102 (N_21102,N_20738,N_20649);
or U21103 (N_21103,N_20596,N_20730);
nand U21104 (N_21104,N_20563,N_20662);
or U21105 (N_21105,N_20693,N_20813);
xnor U21106 (N_21106,N_20997,N_20698);
and U21107 (N_21107,N_20511,N_20515);
xnor U21108 (N_21108,N_20639,N_20759);
or U21109 (N_21109,N_20842,N_20906);
nand U21110 (N_21110,N_20752,N_20810);
nor U21111 (N_21111,N_20970,N_20567);
or U21112 (N_21112,N_20696,N_20670);
and U21113 (N_21113,N_20727,N_20724);
or U21114 (N_21114,N_20624,N_20728);
nand U21115 (N_21115,N_20914,N_20528);
and U21116 (N_21116,N_20933,N_20920);
nand U21117 (N_21117,N_20833,N_20794);
nor U21118 (N_21118,N_20893,N_20721);
xor U21119 (N_21119,N_20988,N_20682);
or U21120 (N_21120,N_20998,N_20978);
xor U21121 (N_21121,N_20875,N_20891);
or U21122 (N_21122,N_20985,N_20701);
nor U21123 (N_21123,N_20882,N_20961);
nand U21124 (N_21124,N_20554,N_20575);
nor U21125 (N_21125,N_20968,N_20975);
xor U21126 (N_21126,N_20745,N_20780);
nor U21127 (N_21127,N_20593,N_20548);
or U21128 (N_21128,N_20741,N_20527);
and U21129 (N_21129,N_20840,N_20545);
nor U21130 (N_21130,N_20557,N_20591);
nor U21131 (N_21131,N_20707,N_20905);
nand U21132 (N_21132,N_20747,N_20938);
xnor U21133 (N_21133,N_20755,N_20806);
nand U21134 (N_21134,N_20603,N_20576);
and U21135 (N_21135,N_20900,N_20616);
or U21136 (N_21136,N_20733,N_20743);
and U21137 (N_21137,N_20872,N_20681);
xnor U21138 (N_21138,N_20513,N_20994);
xor U21139 (N_21139,N_20879,N_20566);
nand U21140 (N_21140,N_20942,N_20799);
nand U21141 (N_21141,N_20931,N_20823);
nor U21142 (N_21142,N_20641,N_20768);
xor U21143 (N_21143,N_20713,N_20645);
nand U21144 (N_21144,N_20832,N_20574);
nor U21145 (N_21145,N_20678,N_20827);
or U21146 (N_21146,N_20611,N_20553);
nor U21147 (N_21147,N_20679,N_20562);
and U21148 (N_21148,N_20767,N_20911);
and U21149 (N_21149,N_20760,N_20694);
and U21150 (N_21150,N_20583,N_20773);
nor U21151 (N_21151,N_20866,N_20826);
and U21152 (N_21152,N_20638,N_20717);
and U21153 (N_21153,N_20777,N_20599);
nand U21154 (N_21154,N_20524,N_20722);
xor U21155 (N_21155,N_20556,N_20784);
nand U21156 (N_21156,N_20935,N_20765);
or U21157 (N_21157,N_20614,N_20723);
xnor U21158 (N_21158,N_20605,N_20621);
nor U21159 (N_21159,N_20666,N_20643);
and U21160 (N_21160,N_20660,N_20676);
nand U21161 (N_21161,N_20963,N_20921);
nand U21162 (N_21162,N_20845,N_20789);
nand U21163 (N_21163,N_20685,N_20688);
nand U21164 (N_21164,N_20706,N_20918);
or U21165 (N_21165,N_20814,N_20937);
xor U21166 (N_21166,N_20860,N_20858);
and U21167 (N_21167,N_20909,N_20983);
or U21168 (N_21168,N_20830,N_20530);
or U21169 (N_21169,N_20628,N_20704);
nor U21170 (N_21170,N_20684,N_20776);
nand U21171 (N_21171,N_20973,N_20579);
nand U21172 (N_21172,N_20770,N_20868);
nand U21173 (N_21173,N_20592,N_20940);
nand U21174 (N_21174,N_20990,N_20546);
nor U21175 (N_21175,N_20652,N_20543);
or U21176 (N_21176,N_20674,N_20620);
and U21177 (N_21177,N_20749,N_20754);
nor U21178 (N_21178,N_20606,N_20610);
nor U21179 (N_21179,N_20714,N_20960);
or U21180 (N_21180,N_20899,N_20658);
and U21181 (N_21181,N_20965,N_20771);
or U21182 (N_21182,N_20954,N_20870);
or U21183 (N_21183,N_20917,N_20800);
xnor U21184 (N_21184,N_20962,N_20841);
xor U21185 (N_21185,N_20807,N_20646);
xor U21186 (N_21186,N_20989,N_20675);
xnor U21187 (N_21187,N_20946,N_20719);
and U21188 (N_21188,N_20869,N_20632);
and U21189 (N_21189,N_20619,N_20865);
nor U21190 (N_21190,N_20774,N_20668);
and U21191 (N_21191,N_20737,N_20769);
nor U21192 (N_21192,N_20846,N_20977);
nand U21193 (N_21193,N_20665,N_20622);
nand U21194 (N_21194,N_20634,N_20715);
xnor U21195 (N_21195,N_20508,N_20926);
or U21196 (N_21196,N_20793,N_20578);
or U21197 (N_21197,N_20949,N_20874);
xnor U21198 (N_21198,N_20878,N_20700);
or U21199 (N_21199,N_20539,N_20916);
nor U21200 (N_21200,N_20581,N_20903);
nor U21201 (N_21201,N_20976,N_20551);
nand U21202 (N_21202,N_20792,N_20825);
and U21203 (N_21203,N_20518,N_20857);
nand U21204 (N_21204,N_20815,N_20598);
nand U21205 (N_21205,N_20588,N_20999);
or U21206 (N_21206,N_20544,N_20779);
nand U21207 (N_21207,N_20533,N_20947);
xnor U21208 (N_21208,N_20570,N_20943);
and U21209 (N_21209,N_20851,N_20889);
nor U21210 (N_21210,N_20659,N_20892);
or U21211 (N_21211,N_20797,N_20689);
xor U21212 (N_21212,N_20731,N_20971);
xor U21213 (N_21213,N_20655,N_20623);
or U21214 (N_21214,N_20635,N_20984);
and U21215 (N_21215,N_20763,N_20854);
and U21216 (N_21216,N_20608,N_20517);
xnor U21217 (N_21217,N_20995,N_20981);
or U21218 (N_21218,N_20712,N_20729);
nand U21219 (N_21219,N_20927,N_20512);
nor U21220 (N_21220,N_20951,N_20820);
nor U21221 (N_21221,N_20819,N_20531);
nor U21222 (N_21222,N_20913,N_20516);
xor U21223 (N_21223,N_20585,N_20758);
or U21224 (N_21224,N_20627,N_20642);
and U21225 (N_21225,N_20718,N_20736);
nor U21226 (N_21226,N_20805,N_20720);
nand U21227 (N_21227,N_20542,N_20657);
or U21228 (N_21228,N_20896,N_20980);
xnor U21229 (N_21229,N_20959,N_20561);
and U21230 (N_21230,N_20671,N_20746);
nand U21231 (N_21231,N_20936,N_20640);
nand U21232 (N_21232,N_20948,N_20669);
nor U21233 (N_21233,N_20922,N_20644);
nand U21234 (N_21234,N_20559,N_20648);
xor U21235 (N_21235,N_20849,N_20672);
xor U21236 (N_21236,N_20509,N_20950);
or U21237 (N_21237,N_20602,N_20744);
and U21238 (N_21238,N_20824,N_20885);
nor U21239 (N_21239,N_20915,N_20664);
nand U21240 (N_21240,N_20568,N_20912);
nor U21241 (N_21241,N_20979,N_20699);
nand U21242 (N_21242,N_20756,N_20584);
nor U21243 (N_21243,N_20601,N_20848);
nor U21244 (N_21244,N_20821,N_20788);
or U21245 (N_21245,N_20790,N_20808);
nor U21246 (N_21246,N_20577,N_20572);
nor U21247 (N_21247,N_20740,N_20709);
or U21248 (N_21248,N_20536,N_20966);
or U21249 (N_21249,N_20751,N_20600);
or U21250 (N_21250,N_20686,N_20774);
or U21251 (N_21251,N_20676,N_20903);
nor U21252 (N_21252,N_20940,N_20651);
nor U21253 (N_21253,N_20510,N_20644);
and U21254 (N_21254,N_20580,N_20957);
nor U21255 (N_21255,N_20819,N_20837);
xor U21256 (N_21256,N_20895,N_20600);
nand U21257 (N_21257,N_20936,N_20595);
or U21258 (N_21258,N_20672,N_20571);
and U21259 (N_21259,N_20951,N_20684);
nor U21260 (N_21260,N_20690,N_20852);
or U21261 (N_21261,N_20620,N_20600);
nand U21262 (N_21262,N_20580,N_20782);
nand U21263 (N_21263,N_20708,N_20930);
xor U21264 (N_21264,N_20622,N_20775);
nand U21265 (N_21265,N_20778,N_20909);
nor U21266 (N_21266,N_20702,N_20695);
and U21267 (N_21267,N_20579,N_20775);
xnor U21268 (N_21268,N_20635,N_20644);
xor U21269 (N_21269,N_20813,N_20683);
and U21270 (N_21270,N_20719,N_20681);
nand U21271 (N_21271,N_20720,N_20844);
and U21272 (N_21272,N_20743,N_20728);
nand U21273 (N_21273,N_20866,N_20766);
or U21274 (N_21274,N_20875,N_20568);
nor U21275 (N_21275,N_20813,N_20548);
nor U21276 (N_21276,N_20997,N_20651);
xor U21277 (N_21277,N_20558,N_20620);
and U21278 (N_21278,N_20657,N_20905);
nand U21279 (N_21279,N_20884,N_20665);
nand U21280 (N_21280,N_20603,N_20510);
xnor U21281 (N_21281,N_20944,N_20546);
xnor U21282 (N_21282,N_20704,N_20978);
or U21283 (N_21283,N_20895,N_20722);
nand U21284 (N_21284,N_20891,N_20584);
and U21285 (N_21285,N_20608,N_20815);
nor U21286 (N_21286,N_20892,N_20867);
or U21287 (N_21287,N_20892,N_20657);
or U21288 (N_21288,N_20541,N_20981);
or U21289 (N_21289,N_20762,N_20881);
and U21290 (N_21290,N_20551,N_20536);
or U21291 (N_21291,N_20720,N_20663);
xnor U21292 (N_21292,N_20515,N_20818);
and U21293 (N_21293,N_20872,N_20576);
nand U21294 (N_21294,N_20739,N_20560);
nor U21295 (N_21295,N_20664,N_20791);
or U21296 (N_21296,N_20882,N_20866);
xor U21297 (N_21297,N_20537,N_20750);
xnor U21298 (N_21298,N_20819,N_20783);
xor U21299 (N_21299,N_20845,N_20502);
or U21300 (N_21300,N_20643,N_20910);
or U21301 (N_21301,N_20953,N_20576);
nand U21302 (N_21302,N_20578,N_20503);
xnor U21303 (N_21303,N_20972,N_20785);
and U21304 (N_21304,N_20911,N_20604);
nor U21305 (N_21305,N_20637,N_20524);
nor U21306 (N_21306,N_20681,N_20566);
or U21307 (N_21307,N_20796,N_20856);
nor U21308 (N_21308,N_20567,N_20767);
xor U21309 (N_21309,N_20626,N_20606);
or U21310 (N_21310,N_20814,N_20736);
xor U21311 (N_21311,N_20941,N_20849);
nand U21312 (N_21312,N_20968,N_20504);
nor U21313 (N_21313,N_20995,N_20809);
or U21314 (N_21314,N_20840,N_20766);
or U21315 (N_21315,N_20557,N_20749);
or U21316 (N_21316,N_20658,N_20641);
nand U21317 (N_21317,N_20652,N_20582);
nor U21318 (N_21318,N_20812,N_20876);
and U21319 (N_21319,N_20662,N_20700);
nor U21320 (N_21320,N_20832,N_20834);
nor U21321 (N_21321,N_20597,N_20950);
or U21322 (N_21322,N_20946,N_20616);
nor U21323 (N_21323,N_20533,N_20531);
nand U21324 (N_21324,N_20603,N_20643);
xnor U21325 (N_21325,N_20757,N_20728);
nand U21326 (N_21326,N_20764,N_20703);
nor U21327 (N_21327,N_20987,N_20803);
or U21328 (N_21328,N_20620,N_20753);
nor U21329 (N_21329,N_20557,N_20561);
and U21330 (N_21330,N_20585,N_20968);
and U21331 (N_21331,N_20989,N_20918);
and U21332 (N_21332,N_20666,N_20574);
and U21333 (N_21333,N_20837,N_20933);
xor U21334 (N_21334,N_20655,N_20868);
or U21335 (N_21335,N_20564,N_20833);
nor U21336 (N_21336,N_20947,N_20740);
nor U21337 (N_21337,N_20782,N_20725);
or U21338 (N_21338,N_20644,N_20684);
or U21339 (N_21339,N_20898,N_20881);
nor U21340 (N_21340,N_20911,N_20814);
and U21341 (N_21341,N_20891,N_20861);
and U21342 (N_21342,N_20599,N_20978);
or U21343 (N_21343,N_20554,N_20543);
nand U21344 (N_21344,N_20909,N_20896);
or U21345 (N_21345,N_20913,N_20613);
or U21346 (N_21346,N_20953,N_20870);
and U21347 (N_21347,N_20818,N_20572);
xor U21348 (N_21348,N_20573,N_20626);
or U21349 (N_21349,N_20661,N_20536);
nand U21350 (N_21350,N_20629,N_20675);
or U21351 (N_21351,N_20761,N_20909);
nor U21352 (N_21352,N_20593,N_20918);
or U21353 (N_21353,N_20658,N_20521);
and U21354 (N_21354,N_20519,N_20827);
nor U21355 (N_21355,N_20743,N_20647);
nor U21356 (N_21356,N_20849,N_20841);
or U21357 (N_21357,N_20828,N_20620);
nand U21358 (N_21358,N_20776,N_20913);
xor U21359 (N_21359,N_20739,N_20646);
nor U21360 (N_21360,N_20777,N_20517);
or U21361 (N_21361,N_20604,N_20602);
xnor U21362 (N_21362,N_20803,N_20939);
and U21363 (N_21363,N_20983,N_20837);
xnor U21364 (N_21364,N_20576,N_20623);
nor U21365 (N_21365,N_20505,N_20501);
xor U21366 (N_21366,N_20962,N_20747);
and U21367 (N_21367,N_20998,N_20727);
xor U21368 (N_21368,N_20854,N_20538);
xnor U21369 (N_21369,N_20716,N_20994);
nand U21370 (N_21370,N_20756,N_20571);
xnor U21371 (N_21371,N_20619,N_20912);
nand U21372 (N_21372,N_20518,N_20925);
nor U21373 (N_21373,N_20703,N_20745);
nand U21374 (N_21374,N_20683,N_20532);
and U21375 (N_21375,N_20533,N_20512);
xnor U21376 (N_21376,N_20829,N_20507);
or U21377 (N_21377,N_20998,N_20995);
and U21378 (N_21378,N_20843,N_20559);
or U21379 (N_21379,N_20518,N_20551);
xnor U21380 (N_21380,N_20817,N_20783);
xor U21381 (N_21381,N_20766,N_20519);
nor U21382 (N_21382,N_20650,N_20628);
xnor U21383 (N_21383,N_20680,N_20754);
nor U21384 (N_21384,N_20512,N_20656);
nand U21385 (N_21385,N_20953,N_20607);
or U21386 (N_21386,N_20680,N_20737);
xnor U21387 (N_21387,N_20654,N_20784);
xor U21388 (N_21388,N_20971,N_20602);
xnor U21389 (N_21389,N_20765,N_20796);
or U21390 (N_21390,N_20584,N_20946);
nor U21391 (N_21391,N_20656,N_20937);
or U21392 (N_21392,N_20552,N_20743);
nand U21393 (N_21393,N_20812,N_20552);
or U21394 (N_21394,N_20820,N_20858);
nor U21395 (N_21395,N_20710,N_20577);
or U21396 (N_21396,N_20573,N_20782);
nor U21397 (N_21397,N_20878,N_20642);
and U21398 (N_21398,N_20588,N_20662);
nand U21399 (N_21399,N_20924,N_20735);
nand U21400 (N_21400,N_20548,N_20840);
and U21401 (N_21401,N_20546,N_20579);
xnor U21402 (N_21402,N_20669,N_20887);
nand U21403 (N_21403,N_20999,N_20593);
xor U21404 (N_21404,N_20731,N_20584);
or U21405 (N_21405,N_20559,N_20674);
nor U21406 (N_21406,N_20778,N_20512);
nor U21407 (N_21407,N_20930,N_20821);
nand U21408 (N_21408,N_20577,N_20889);
nand U21409 (N_21409,N_20802,N_20565);
nand U21410 (N_21410,N_20612,N_20713);
nor U21411 (N_21411,N_20834,N_20563);
and U21412 (N_21412,N_20816,N_20579);
nand U21413 (N_21413,N_20852,N_20801);
xor U21414 (N_21414,N_20822,N_20930);
xor U21415 (N_21415,N_20728,N_20694);
and U21416 (N_21416,N_20541,N_20742);
nand U21417 (N_21417,N_20705,N_20884);
and U21418 (N_21418,N_20884,N_20847);
nand U21419 (N_21419,N_20881,N_20537);
xor U21420 (N_21420,N_20513,N_20719);
xor U21421 (N_21421,N_20996,N_20709);
nor U21422 (N_21422,N_20721,N_20852);
and U21423 (N_21423,N_20969,N_20875);
nor U21424 (N_21424,N_20979,N_20600);
xnor U21425 (N_21425,N_20566,N_20707);
or U21426 (N_21426,N_20713,N_20671);
and U21427 (N_21427,N_20780,N_20864);
nor U21428 (N_21428,N_20901,N_20805);
nor U21429 (N_21429,N_20899,N_20552);
xnor U21430 (N_21430,N_20825,N_20642);
nor U21431 (N_21431,N_20767,N_20704);
and U21432 (N_21432,N_20668,N_20509);
xnor U21433 (N_21433,N_20742,N_20862);
nand U21434 (N_21434,N_20935,N_20595);
nor U21435 (N_21435,N_20878,N_20580);
xnor U21436 (N_21436,N_20921,N_20741);
and U21437 (N_21437,N_20593,N_20888);
nand U21438 (N_21438,N_20565,N_20727);
and U21439 (N_21439,N_20691,N_20800);
or U21440 (N_21440,N_20734,N_20862);
and U21441 (N_21441,N_20813,N_20734);
and U21442 (N_21442,N_20676,N_20929);
and U21443 (N_21443,N_20944,N_20896);
or U21444 (N_21444,N_20708,N_20618);
nor U21445 (N_21445,N_20786,N_20956);
nor U21446 (N_21446,N_20576,N_20694);
or U21447 (N_21447,N_20578,N_20785);
xnor U21448 (N_21448,N_20944,N_20551);
and U21449 (N_21449,N_20862,N_20570);
nor U21450 (N_21450,N_20560,N_20539);
nand U21451 (N_21451,N_20682,N_20872);
nand U21452 (N_21452,N_20726,N_20593);
or U21453 (N_21453,N_20702,N_20585);
nand U21454 (N_21454,N_20523,N_20565);
nand U21455 (N_21455,N_20987,N_20652);
or U21456 (N_21456,N_20541,N_20856);
nor U21457 (N_21457,N_20932,N_20686);
and U21458 (N_21458,N_20824,N_20682);
or U21459 (N_21459,N_20589,N_20539);
nor U21460 (N_21460,N_20501,N_20728);
nor U21461 (N_21461,N_20589,N_20755);
nor U21462 (N_21462,N_20953,N_20691);
nor U21463 (N_21463,N_20799,N_20696);
or U21464 (N_21464,N_20552,N_20628);
nand U21465 (N_21465,N_20700,N_20680);
xnor U21466 (N_21466,N_20707,N_20683);
xnor U21467 (N_21467,N_20874,N_20927);
and U21468 (N_21468,N_20785,N_20544);
xor U21469 (N_21469,N_20550,N_20766);
xor U21470 (N_21470,N_20862,N_20811);
xor U21471 (N_21471,N_20698,N_20843);
nor U21472 (N_21472,N_20553,N_20600);
nor U21473 (N_21473,N_20729,N_20652);
or U21474 (N_21474,N_20777,N_20507);
nand U21475 (N_21475,N_20744,N_20563);
or U21476 (N_21476,N_20651,N_20720);
nor U21477 (N_21477,N_20781,N_20810);
xor U21478 (N_21478,N_20896,N_20528);
nor U21479 (N_21479,N_20833,N_20882);
and U21480 (N_21480,N_20622,N_20869);
or U21481 (N_21481,N_20628,N_20919);
nand U21482 (N_21482,N_20705,N_20535);
nand U21483 (N_21483,N_20675,N_20693);
xnor U21484 (N_21484,N_20611,N_20511);
xor U21485 (N_21485,N_20921,N_20634);
xor U21486 (N_21486,N_20587,N_20769);
nor U21487 (N_21487,N_20503,N_20954);
nor U21488 (N_21488,N_20877,N_20597);
xor U21489 (N_21489,N_20547,N_20744);
xor U21490 (N_21490,N_20947,N_20917);
xor U21491 (N_21491,N_20931,N_20517);
nor U21492 (N_21492,N_20560,N_20548);
nand U21493 (N_21493,N_20616,N_20829);
and U21494 (N_21494,N_20821,N_20968);
and U21495 (N_21495,N_20948,N_20978);
or U21496 (N_21496,N_20902,N_20538);
and U21497 (N_21497,N_20946,N_20679);
nand U21498 (N_21498,N_20606,N_20864);
nand U21499 (N_21499,N_20518,N_20944);
and U21500 (N_21500,N_21455,N_21153);
xnor U21501 (N_21501,N_21255,N_21196);
or U21502 (N_21502,N_21338,N_21052);
nor U21503 (N_21503,N_21224,N_21361);
nand U21504 (N_21504,N_21206,N_21216);
nand U21505 (N_21505,N_21372,N_21069);
xor U21506 (N_21506,N_21482,N_21440);
xor U21507 (N_21507,N_21312,N_21250);
nor U21508 (N_21508,N_21335,N_21443);
xnor U21509 (N_21509,N_21063,N_21041);
nor U21510 (N_21510,N_21367,N_21138);
nand U21511 (N_21511,N_21141,N_21350);
or U21512 (N_21512,N_21476,N_21266);
xor U21513 (N_21513,N_21466,N_21131);
xor U21514 (N_21514,N_21129,N_21448);
or U21515 (N_21515,N_21225,N_21371);
and U21516 (N_21516,N_21008,N_21322);
xor U21517 (N_21517,N_21092,N_21495);
nor U21518 (N_21518,N_21125,N_21184);
or U21519 (N_21519,N_21114,N_21182);
and U21520 (N_21520,N_21435,N_21139);
or U21521 (N_21521,N_21029,N_21379);
xor U21522 (N_21522,N_21079,N_21073);
nor U21523 (N_21523,N_21414,N_21486);
nor U21524 (N_21524,N_21144,N_21161);
nor U21525 (N_21525,N_21178,N_21355);
nand U21526 (N_21526,N_21168,N_21028);
nor U21527 (N_21527,N_21413,N_21269);
and U21528 (N_21528,N_21354,N_21062);
nand U21529 (N_21529,N_21391,N_21475);
nor U21530 (N_21530,N_21427,N_21296);
nand U21531 (N_21531,N_21356,N_21242);
nand U21532 (N_21532,N_21202,N_21173);
nand U21533 (N_21533,N_21383,N_21002);
xnor U21534 (N_21534,N_21319,N_21246);
nor U21535 (N_21535,N_21146,N_21169);
or U21536 (N_21536,N_21290,N_21087);
nor U21537 (N_21537,N_21472,N_21232);
nor U21538 (N_21538,N_21439,N_21497);
or U21539 (N_21539,N_21108,N_21357);
or U21540 (N_21540,N_21452,N_21288);
xnor U21541 (N_21541,N_21263,N_21085);
and U21542 (N_21542,N_21267,N_21336);
and U21543 (N_21543,N_21033,N_21035);
and U21544 (N_21544,N_21285,N_21140);
or U21545 (N_21545,N_21396,N_21183);
or U21546 (N_21546,N_21309,N_21281);
or U21547 (N_21547,N_21223,N_21037);
or U21548 (N_21548,N_21284,N_21231);
and U21549 (N_21549,N_21077,N_21294);
and U21550 (N_21550,N_21226,N_21038);
and U21551 (N_21551,N_21351,N_21326);
or U21552 (N_21552,N_21289,N_21292);
nand U21553 (N_21553,N_21245,N_21420);
nor U21554 (N_21554,N_21042,N_21494);
or U21555 (N_21555,N_21148,N_21253);
and U21556 (N_21556,N_21270,N_21323);
nor U21557 (N_21557,N_21282,N_21445);
nand U21558 (N_21558,N_21074,N_21358);
nand U21559 (N_21559,N_21009,N_21498);
nand U21560 (N_21560,N_21278,N_21024);
nor U21561 (N_21561,N_21080,N_21101);
xnor U21562 (N_21562,N_21421,N_21327);
nand U21563 (N_21563,N_21104,N_21329);
or U21564 (N_21564,N_21291,N_21053);
xnor U21565 (N_21565,N_21280,N_21318);
nor U21566 (N_21566,N_21341,N_21166);
xor U21567 (N_21567,N_21469,N_21483);
nor U21568 (N_21568,N_21222,N_21429);
or U21569 (N_21569,N_21147,N_21411);
nor U21570 (N_21570,N_21212,N_21170);
or U21571 (N_21571,N_21057,N_21404);
and U21572 (N_21572,N_21164,N_21082);
xnor U21573 (N_21573,N_21259,N_21369);
xor U21574 (N_21574,N_21091,N_21172);
nand U21575 (N_21575,N_21333,N_21463);
xor U21576 (N_21576,N_21058,N_21401);
nor U21577 (N_21577,N_21247,N_21377);
or U21578 (N_21578,N_21484,N_21459);
xor U21579 (N_21579,N_21218,N_21115);
and U21580 (N_21580,N_21229,N_21477);
nand U21581 (N_21581,N_21103,N_21393);
and U21582 (N_21582,N_21145,N_21277);
nor U21583 (N_21583,N_21493,N_21241);
nand U21584 (N_21584,N_21437,N_21228);
nor U21585 (N_21585,N_21339,N_21415);
or U21586 (N_21586,N_21464,N_21344);
nor U21587 (N_21587,N_21100,N_21286);
nor U21588 (N_21588,N_21478,N_21258);
or U21589 (N_21589,N_21032,N_21456);
xnor U21590 (N_21590,N_21066,N_21378);
nand U21591 (N_21591,N_21113,N_21015);
nor U21592 (N_21592,N_21382,N_21394);
nor U21593 (N_21593,N_21025,N_21340);
nor U21594 (N_21594,N_21175,N_21198);
nor U21595 (N_21595,N_21210,N_21126);
or U21596 (N_21596,N_21021,N_21449);
nor U21597 (N_21597,N_21380,N_21174);
and U21598 (N_21598,N_21201,N_21217);
nand U21599 (N_21599,N_21271,N_21432);
and U21600 (N_21600,N_21458,N_21013);
nor U21601 (N_21601,N_21177,N_21499);
and U21602 (N_21602,N_21390,N_21248);
or U21603 (N_21603,N_21107,N_21330);
nand U21604 (N_21604,N_21453,N_21023);
xnor U21605 (N_21605,N_21306,N_21213);
xor U21606 (N_21606,N_21111,N_21046);
or U21607 (N_21607,N_21214,N_21417);
xor U21608 (N_21608,N_21098,N_21007);
and U21609 (N_21609,N_21190,N_21020);
xor U21610 (N_21610,N_21334,N_21345);
nor U21611 (N_21611,N_21157,N_21311);
and U21612 (N_21612,N_21055,N_21352);
nand U21613 (N_21613,N_21343,N_21095);
nor U21614 (N_21614,N_21457,N_21049);
xor U21615 (N_21615,N_21374,N_21447);
or U21616 (N_21616,N_21363,N_21233);
and U21617 (N_21617,N_21385,N_21188);
nor U21618 (N_21618,N_21436,N_21237);
nand U21619 (N_21619,N_21451,N_21460);
xor U21620 (N_21620,N_21328,N_21018);
xor U21621 (N_21621,N_21011,N_21122);
xor U21622 (N_21622,N_21155,N_21130);
or U21623 (N_21623,N_21254,N_21102);
and U21624 (N_21624,N_21219,N_21299);
xor U21625 (N_21625,N_21488,N_21158);
or U21626 (N_21626,N_21489,N_21264);
xnor U21627 (N_21627,N_21422,N_21310);
xor U21628 (N_21628,N_21181,N_21403);
and U21629 (N_21629,N_21252,N_21321);
xor U21630 (N_21630,N_21315,N_21121);
and U21631 (N_21631,N_21471,N_21428);
xor U21632 (N_21632,N_21465,N_21287);
nor U21633 (N_21633,N_21165,N_21362);
xnor U21634 (N_21634,N_21234,N_21434);
nand U21635 (N_21635,N_21059,N_21143);
or U21636 (N_21636,N_21416,N_21016);
or U21637 (N_21637,N_21093,N_21308);
xor U21638 (N_21638,N_21039,N_21200);
or U21639 (N_21639,N_21105,N_21425);
nor U21640 (N_21640,N_21159,N_21019);
xor U21641 (N_21641,N_21342,N_21000);
and U21642 (N_21642,N_21468,N_21313);
nor U21643 (N_21643,N_21317,N_21185);
xnor U21644 (N_21644,N_21127,N_21251);
nand U21645 (N_21645,N_21387,N_21208);
and U21646 (N_21646,N_21090,N_21106);
or U21647 (N_21647,N_21441,N_21189);
and U21648 (N_21648,N_21368,N_21419);
or U21649 (N_21649,N_21300,N_21167);
nor U21650 (N_21650,N_21444,N_21081);
xor U21651 (N_21651,N_21076,N_21179);
xnor U21652 (N_21652,N_21137,N_21423);
nand U21653 (N_21653,N_21275,N_21261);
nor U21654 (N_21654,N_21132,N_21227);
or U21655 (N_21655,N_21418,N_21118);
xor U21656 (N_21656,N_21487,N_21431);
or U21657 (N_21657,N_21112,N_21134);
nand U21658 (N_21658,N_21462,N_21197);
or U21659 (N_21659,N_21154,N_21221);
or U21660 (N_21660,N_21078,N_21051);
nand U21661 (N_21661,N_21301,N_21133);
and U21662 (N_21662,N_21410,N_21470);
nand U21663 (N_21663,N_21324,N_21479);
and U21664 (N_21664,N_21316,N_21381);
nor U21665 (N_21665,N_21050,N_21065);
nor U21666 (N_21666,N_21480,N_21490);
and U21667 (N_21667,N_21260,N_21293);
nand U21668 (N_21668,N_21392,N_21454);
and U21669 (N_21669,N_21012,N_21194);
nor U21670 (N_21670,N_21359,N_21240);
nand U21671 (N_21671,N_21320,N_21060);
and U21672 (N_21672,N_21207,N_21388);
xor U21673 (N_21673,N_21407,N_21047);
xor U21674 (N_21674,N_21083,N_21048);
nor U21675 (N_21675,N_21384,N_21027);
nand U21676 (N_21676,N_21474,N_21199);
and U21677 (N_21677,N_21203,N_21176);
xnor U21678 (N_21678,N_21373,N_21068);
xnor U21679 (N_21679,N_21249,N_21473);
nand U21680 (N_21680,N_21446,N_21239);
and U21681 (N_21681,N_21283,N_21257);
or U21682 (N_21682,N_21005,N_21119);
and U21683 (N_21683,N_21337,N_21142);
and U21684 (N_21684,N_21180,N_21209);
nand U21685 (N_21685,N_21001,N_21043);
nand U21686 (N_21686,N_21215,N_21135);
xor U21687 (N_21687,N_21022,N_21353);
and U21688 (N_21688,N_21297,N_21268);
or U21689 (N_21689,N_21097,N_21128);
or U21690 (N_21690,N_21109,N_21156);
or U21691 (N_21691,N_21163,N_21072);
nor U21692 (N_21692,N_21204,N_21070);
nand U21693 (N_21693,N_21365,N_21056);
xor U21694 (N_21694,N_21405,N_21150);
or U21695 (N_21695,N_21347,N_21193);
nor U21696 (N_21696,N_21366,N_21014);
or U21697 (N_21697,N_21348,N_21044);
xor U21698 (N_21698,N_21116,N_21205);
nor U21699 (N_21699,N_21084,N_21026);
or U21700 (N_21700,N_21430,N_21243);
or U21701 (N_21701,N_21017,N_21149);
and U21702 (N_21702,N_21426,N_21433);
nand U21703 (N_21703,N_21450,N_21152);
nand U21704 (N_21704,N_21325,N_21461);
nor U21705 (N_21705,N_21364,N_21235);
nor U21706 (N_21706,N_21096,N_21398);
or U21707 (N_21707,N_21003,N_21136);
nor U21708 (N_21708,N_21467,N_21031);
xnor U21709 (N_21709,N_21370,N_21346);
and U21710 (N_21710,N_21304,N_21438);
or U21711 (N_21711,N_21064,N_21220);
xor U21712 (N_21712,N_21303,N_21279);
nor U21713 (N_21713,N_21397,N_21086);
nor U21714 (N_21714,N_21195,N_21067);
or U21715 (N_21715,N_21402,N_21412);
or U21716 (N_21716,N_21492,N_21302);
xnor U21717 (N_21717,N_21399,N_21481);
xnor U21718 (N_21718,N_21191,N_21307);
nand U21719 (N_21719,N_21262,N_21314);
xor U21720 (N_21720,N_21376,N_21117);
xor U21721 (N_21721,N_21094,N_21061);
xor U21722 (N_21722,N_21409,N_21265);
nand U21723 (N_21723,N_21036,N_21406);
xnor U21724 (N_21724,N_21295,N_21071);
nand U21725 (N_21725,N_21276,N_21120);
or U21726 (N_21726,N_21273,N_21360);
xnor U21727 (N_21727,N_21230,N_21331);
or U21728 (N_21728,N_21124,N_21045);
nand U21729 (N_21729,N_21408,N_21004);
nand U21730 (N_21730,N_21395,N_21192);
nor U21731 (N_21731,N_21375,N_21110);
nand U21732 (N_21732,N_21099,N_21030);
and U21733 (N_21733,N_21160,N_21332);
nand U21734 (N_21734,N_21491,N_21089);
nand U21735 (N_21735,N_21040,N_21123);
nor U21736 (N_21736,N_21171,N_21034);
or U21737 (N_21737,N_21424,N_21010);
nor U21738 (N_21738,N_21386,N_21442);
nand U21739 (N_21739,N_21298,N_21187);
or U21740 (N_21740,N_21006,N_21400);
nand U21741 (N_21741,N_21211,N_21162);
or U21742 (N_21742,N_21349,N_21054);
nor U21743 (N_21743,N_21186,N_21389);
or U21744 (N_21744,N_21075,N_21272);
and U21745 (N_21745,N_21151,N_21256);
or U21746 (N_21746,N_21274,N_21238);
nand U21747 (N_21747,N_21236,N_21485);
xnor U21748 (N_21748,N_21305,N_21088);
nand U21749 (N_21749,N_21244,N_21496);
nor U21750 (N_21750,N_21174,N_21128);
nand U21751 (N_21751,N_21052,N_21415);
nor U21752 (N_21752,N_21393,N_21128);
nor U21753 (N_21753,N_21166,N_21348);
and U21754 (N_21754,N_21022,N_21468);
and U21755 (N_21755,N_21189,N_21113);
nor U21756 (N_21756,N_21217,N_21338);
xnor U21757 (N_21757,N_21498,N_21315);
and U21758 (N_21758,N_21289,N_21157);
and U21759 (N_21759,N_21368,N_21135);
or U21760 (N_21760,N_21480,N_21089);
or U21761 (N_21761,N_21081,N_21276);
and U21762 (N_21762,N_21196,N_21483);
nand U21763 (N_21763,N_21082,N_21369);
xnor U21764 (N_21764,N_21387,N_21450);
and U21765 (N_21765,N_21057,N_21117);
and U21766 (N_21766,N_21179,N_21429);
nor U21767 (N_21767,N_21051,N_21248);
or U21768 (N_21768,N_21153,N_21476);
xnor U21769 (N_21769,N_21238,N_21078);
nand U21770 (N_21770,N_21185,N_21295);
nand U21771 (N_21771,N_21293,N_21323);
nand U21772 (N_21772,N_21339,N_21241);
nand U21773 (N_21773,N_21017,N_21179);
nand U21774 (N_21774,N_21215,N_21226);
xnor U21775 (N_21775,N_21138,N_21241);
and U21776 (N_21776,N_21209,N_21341);
xnor U21777 (N_21777,N_21106,N_21317);
and U21778 (N_21778,N_21129,N_21004);
nor U21779 (N_21779,N_21191,N_21337);
nand U21780 (N_21780,N_21274,N_21292);
nor U21781 (N_21781,N_21480,N_21020);
nand U21782 (N_21782,N_21389,N_21469);
nand U21783 (N_21783,N_21072,N_21068);
nor U21784 (N_21784,N_21476,N_21224);
xnor U21785 (N_21785,N_21092,N_21362);
nand U21786 (N_21786,N_21254,N_21381);
or U21787 (N_21787,N_21454,N_21098);
nor U21788 (N_21788,N_21233,N_21325);
and U21789 (N_21789,N_21019,N_21089);
nor U21790 (N_21790,N_21189,N_21446);
xnor U21791 (N_21791,N_21038,N_21193);
nor U21792 (N_21792,N_21156,N_21401);
nor U21793 (N_21793,N_21133,N_21041);
nor U21794 (N_21794,N_21270,N_21035);
or U21795 (N_21795,N_21457,N_21090);
and U21796 (N_21796,N_21205,N_21241);
nand U21797 (N_21797,N_21210,N_21157);
or U21798 (N_21798,N_21333,N_21424);
and U21799 (N_21799,N_21372,N_21138);
nor U21800 (N_21800,N_21453,N_21008);
nand U21801 (N_21801,N_21287,N_21058);
nand U21802 (N_21802,N_21401,N_21380);
nand U21803 (N_21803,N_21400,N_21357);
nor U21804 (N_21804,N_21345,N_21198);
nor U21805 (N_21805,N_21295,N_21377);
nor U21806 (N_21806,N_21416,N_21440);
nor U21807 (N_21807,N_21279,N_21102);
and U21808 (N_21808,N_21276,N_21485);
xor U21809 (N_21809,N_21397,N_21415);
nor U21810 (N_21810,N_21301,N_21008);
nand U21811 (N_21811,N_21443,N_21285);
xor U21812 (N_21812,N_21394,N_21100);
and U21813 (N_21813,N_21228,N_21043);
xnor U21814 (N_21814,N_21102,N_21272);
nor U21815 (N_21815,N_21104,N_21477);
nand U21816 (N_21816,N_21126,N_21427);
nor U21817 (N_21817,N_21097,N_21116);
xnor U21818 (N_21818,N_21154,N_21155);
and U21819 (N_21819,N_21035,N_21286);
or U21820 (N_21820,N_21318,N_21370);
nand U21821 (N_21821,N_21418,N_21406);
xnor U21822 (N_21822,N_21261,N_21288);
and U21823 (N_21823,N_21497,N_21232);
or U21824 (N_21824,N_21414,N_21068);
nor U21825 (N_21825,N_21154,N_21030);
and U21826 (N_21826,N_21039,N_21497);
xor U21827 (N_21827,N_21105,N_21493);
or U21828 (N_21828,N_21060,N_21002);
or U21829 (N_21829,N_21430,N_21272);
nor U21830 (N_21830,N_21494,N_21379);
nand U21831 (N_21831,N_21496,N_21079);
nand U21832 (N_21832,N_21043,N_21338);
xnor U21833 (N_21833,N_21473,N_21281);
and U21834 (N_21834,N_21197,N_21378);
and U21835 (N_21835,N_21357,N_21284);
xor U21836 (N_21836,N_21440,N_21368);
nor U21837 (N_21837,N_21065,N_21033);
nand U21838 (N_21838,N_21157,N_21222);
nand U21839 (N_21839,N_21247,N_21046);
and U21840 (N_21840,N_21469,N_21214);
nand U21841 (N_21841,N_21292,N_21184);
xor U21842 (N_21842,N_21479,N_21125);
and U21843 (N_21843,N_21078,N_21358);
xnor U21844 (N_21844,N_21250,N_21431);
or U21845 (N_21845,N_21121,N_21255);
xor U21846 (N_21846,N_21347,N_21020);
nor U21847 (N_21847,N_21441,N_21222);
nand U21848 (N_21848,N_21235,N_21445);
or U21849 (N_21849,N_21223,N_21338);
or U21850 (N_21850,N_21219,N_21199);
and U21851 (N_21851,N_21409,N_21364);
or U21852 (N_21852,N_21161,N_21469);
xor U21853 (N_21853,N_21437,N_21260);
nor U21854 (N_21854,N_21398,N_21347);
and U21855 (N_21855,N_21055,N_21013);
or U21856 (N_21856,N_21242,N_21179);
nand U21857 (N_21857,N_21133,N_21326);
xnor U21858 (N_21858,N_21255,N_21167);
or U21859 (N_21859,N_21348,N_21289);
and U21860 (N_21860,N_21396,N_21059);
nor U21861 (N_21861,N_21492,N_21258);
nor U21862 (N_21862,N_21107,N_21487);
or U21863 (N_21863,N_21363,N_21263);
and U21864 (N_21864,N_21313,N_21291);
nor U21865 (N_21865,N_21275,N_21051);
or U21866 (N_21866,N_21014,N_21181);
and U21867 (N_21867,N_21023,N_21128);
nor U21868 (N_21868,N_21156,N_21187);
or U21869 (N_21869,N_21111,N_21117);
nand U21870 (N_21870,N_21436,N_21148);
nor U21871 (N_21871,N_21042,N_21467);
or U21872 (N_21872,N_21040,N_21472);
or U21873 (N_21873,N_21222,N_21075);
nor U21874 (N_21874,N_21433,N_21079);
nor U21875 (N_21875,N_21156,N_21293);
nor U21876 (N_21876,N_21438,N_21272);
xnor U21877 (N_21877,N_21323,N_21220);
nand U21878 (N_21878,N_21476,N_21060);
xnor U21879 (N_21879,N_21256,N_21191);
or U21880 (N_21880,N_21006,N_21458);
or U21881 (N_21881,N_21458,N_21199);
or U21882 (N_21882,N_21474,N_21008);
and U21883 (N_21883,N_21001,N_21347);
xnor U21884 (N_21884,N_21453,N_21373);
and U21885 (N_21885,N_21236,N_21101);
and U21886 (N_21886,N_21088,N_21001);
and U21887 (N_21887,N_21205,N_21272);
or U21888 (N_21888,N_21215,N_21095);
and U21889 (N_21889,N_21370,N_21461);
nor U21890 (N_21890,N_21240,N_21081);
and U21891 (N_21891,N_21195,N_21315);
and U21892 (N_21892,N_21125,N_21062);
or U21893 (N_21893,N_21334,N_21085);
nor U21894 (N_21894,N_21213,N_21197);
or U21895 (N_21895,N_21037,N_21200);
or U21896 (N_21896,N_21357,N_21089);
or U21897 (N_21897,N_21374,N_21149);
and U21898 (N_21898,N_21488,N_21430);
nor U21899 (N_21899,N_21411,N_21403);
xnor U21900 (N_21900,N_21440,N_21210);
and U21901 (N_21901,N_21253,N_21135);
or U21902 (N_21902,N_21297,N_21181);
or U21903 (N_21903,N_21320,N_21360);
nand U21904 (N_21904,N_21082,N_21138);
xnor U21905 (N_21905,N_21374,N_21288);
and U21906 (N_21906,N_21294,N_21422);
nor U21907 (N_21907,N_21032,N_21374);
or U21908 (N_21908,N_21185,N_21269);
and U21909 (N_21909,N_21038,N_21013);
and U21910 (N_21910,N_21483,N_21038);
xnor U21911 (N_21911,N_21319,N_21067);
xnor U21912 (N_21912,N_21026,N_21205);
nor U21913 (N_21913,N_21026,N_21250);
and U21914 (N_21914,N_21328,N_21100);
nand U21915 (N_21915,N_21179,N_21240);
nand U21916 (N_21916,N_21366,N_21438);
xnor U21917 (N_21917,N_21266,N_21100);
xnor U21918 (N_21918,N_21062,N_21370);
xor U21919 (N_21919,N_21332,N_21322);
nor U21920 (N_21920,N_21113,N_21106);
and U21921 (N_21921,N_21311,N_21139);
nand U21922 (N_21922,N_21386,N_21028);
nand U21923 (N_21923,N_21108,N_21302);
nor U21924 (N_21924,N_21215,N_21230);
or U21925 (N_21925,N_21426,N_21148);
and U21926 (N_21926,N_21474,N_21164);
xor U21927 (N_21927,N_21093,N_21409);
xnor U21928 (N_21928,N_21378,N_21284);
nand U21929 (N_21929,N_21283,N_21373);
nor U21930 (N_21930,N_21378,N_21345);
or U21931 (N_21931,N_21176,N_21139);
xor U21932 (N_21932,N_21173,N_21070);
nor U21933 (N_21933,N_21129,N_21440);
xnor U21934 (N_21934,N_21298,N_21285);
and U21935 (N_21935,N_21218,N_21092);
xnor U21936 (N_21936,N_21033,N_21102);
xor U21937 (N_21937,N_21456,N_21308);
xnor U21938 (N_21938,N_21030,N_21497);
nand U21939 (N_21939,N_21135,N_21059);
and U21940 (N_21940,N_21473,N_21413);
and U21941 (N_21941,N_21012,N_21063);
nand U21942 (N_21942,N_21140,N_21064);
nand U21943 (N_21943,N_21145,N_21054);
and U21944 (N_21944,N_21361,N_21210);
nor U21945 (N_21945,N_21344,N_21198);
nand U21946 (N_21946,N_21075,N_21035);
xnor U21947 (N_21947,N_21041,N_21243);
and U21948 (N_21948,N_21463,N_21427);
or U21949 (N_21949,N_21020,N_21452);
and U21950 (N_21950,N_21271,N_21066);
or U21951 (N_21951,N_21474,N_21243);
nand U21952 (N_21952,N_21465,N_21200);
nand U21953 (N_21953,N_21070,N_21294);
and U21954 (N_21954,N_21277,N_21324);
or U21955 (N_21955,N_21158,N_21397);
nand U21956 (N_21956,N_21207,N_21296);
and U21957 (N_21957,N_21494,N_21008);
and U21958 (N_21958,N_21030,N_21038);
nand U21959 (N_21959,N_21259,N_21420);
nand U21960 (N_21960,N_21049,N_21356);
or U21961 (N_21961,N_21000,N_21304);
nor U21962 (N_21962,N_21041,N_21342);
and U21963 (N_21963,N_21055,N_21316);
nand U21964 (N_21964,N_21291,N_21471);
nand U21965 (N_21965,N_21212,N_21195);
xnor U21966 (N_21966,N_21220,N_21228);
or U21967 (N_21967,N_21290,N_21197);
nor U21968 (N_21968,N_21368,N_21340);
xnor U21969 (N_21969,N_21321,N_21258);
and U21970 (N_21970,N_21346,N_21394);
and U21971 (N_21971,N_21484,N_21201);
nand U21972 (N_21972,N_21226,N_21160);
nor U21973 (N_21973,N_21070,N_21392);
and U21974 (N_21974,N_21412,N_21400);
nand U21975 (N_21975,N_21207,N_21170);
nor U21976 (N_21976,N_21498,N_21419);
nor U21977 (N_21977,N_21210,N_21476);
or U21978 (N_21978,N_21112,N_21453);
nand U21979 (N_21979,N_21275,N_21024);
nor U21980 (N_21980,N_21145,N_21484);
nand U21981 (N_21981,N_21461,N_21298);
nand U21982 (N_21982,N_21346,N_21292);
nor U21983 (N_21983,N_21089,N_21050);
xor U21984 (N_21984,N_21448,N_21482);
or U21985 (N_21985,N_21076,N_21335);
nand U21986 (N_21986,N_21036,N_21111);
xor U21987 (N_21987,N_21064,N_21053);
xnor U21988 (N_21988,N_21401,N_21000);
or U21989 (N_21989,N_21173,N_21439);
xor U21990 (N_21990,N_21016,N_21232);
nand U21991 (N_21991,N_21380,N_21018);
xor U21992 (N_21992,N_21211,N_21169);
xnor U21993 (N_21993,N_21086,N_21490);
nand U21994 (N_21994,N_21336,N_21121);
or U21995 (N_21995,N_21336,N_21466);
and U21996 (N_21996,N_21225,N_21086);
nor U21997 (N_21997,N_21054,N_21453);
xor U21998 (N_21998,N_21017,N_21289);
nor U21999 (N_21999,N_21415,N_21211);
nand U22000 (N_22000,N_21655,N_21537);
xor U22001 (N_22001,N_21595,N_21778);
xor U22002 (N_22002,N_21749,N_21626);
nor U22003 (N_22003,N_21757,N_21692);
nand U22004 (N_22004,N_21905,N_21989);
and U22005 (N_22005,N_21566,N_21616);
nor U22006 (N_22006,N_21715,N_21853);
nor U22007 (N_22007,N_21928,N_21795);
nor U22008 (N_22008,N_21503,N_21697);
or U22009 (N_22009,N_21636,N_21965);
nor U22010 (N_22010,N_21777,N_21885);
and U22011 (N_22011,N_21984,N_21577);
nand U22012 (N_22012,N_21745,N_21890);
nand U22013 (N_22013,N_21953,N_21546);
nor U22014 (N_22014,N_21824,N_21644);
xnor U22015 (N_22015,N_21932,N_21833);
and U22016 (N_22016,N_21855,N_21772);
xor U22017 (N_22017,N_21531,N_21719);
xor U22018 (N_22018,N_21962,N_21542);
and U22019 (N_22019,N_21527,N_21549);
xor U22020 (N_22020,N_21797,N_21633);
and U22021 (N_22021,N_21974,N_21760);
and U22022 (N_22022,N_21957,N_21599);
nor U22023 (N_22023,N_21500,N_21718);
xnor U22024 (N_22024,N_21608,N_21679);
xor U22025 (N_22025,N_21628,N_21893);
nand U22026 (N_22026,N_21758,N_21627);
nor U22027 (N_22027,N_21548,N_21975);
and U22028 (N_22028,N_21638,N_21743);
or U22029 (N_22029,N_21530,N_21843);
xor U22030 (N_22030,N_21731,N_21686);
nand U22031 (N_22031,N_21898,N_21774);
nor U22032 (N_22032,N_21553,N_21990);
nand U22033 (N_22033,N_21755,N_21683);
or U22034 (N_22034,N_21939,N_21820);
xnor U22035 (N_22035,N_21654,N_21819);
xor U22036 (N_22036,N_21884,N_21763);
nand U22037 (N_22037,N_21732,N_21609);
xor U22038 (N_22038,N_21541,N_21986);
xor U22039 (N_22039,N_21594,N_21648);
or U22040 (N_22040,N_21647,N_21614);
or U22041 (N_22041,N_21729,N_21867);
nand U22042 (N_22042,N_21872,N_21857);
nor U22043 (N_22043,N_21769,N_21761);
nor U22044 (N_22044,N_21680,N_21925);
nand U22045 (N_22045,N_21949,N_21904);
nor U22046 (N_22046,N_21800,N_21584);
xnor U22047 (N_22047,N_21994,N_21750);
and U22048 (N_22048,N_21726,N_21524);
and U22049 (N_22049,N_21883,N_21722);
and U22050 (N_22050,N_21702,N_21910);
xor U22051 (N_22051,N_21861,N_21678);
nor U22052 (N_22052,N_21543,N_21799);
nand U22053 (N_22053,N_21838,N_21913);
nand U22054 (N_22054,N_21987,N_21656);
xnor U22055 (N_22055,N_21779,N_21600);
or U22056 (N_22056,N_21725,N_21922);
nand U22057 (N_22057,N_21730,N_21558);
xnor U22058 (N_22058,N_21512,N_21555);
nand U22059 (N_22059,N_21878,N_21788);
nor U22060 (N_22060,N_21746,N_21534);
nand U22061 (N_22061,N_21858,N_21579);
xnor U22062 (N_22062,N_21752,N_21552);
or U22063 (N_22063,N_21604,N_21593);
and U22064 (N_22064,N_21508,N_21864);
nand U22065 (N_22065,N_21682,N_21873);
or U22066 (N_22066,N_21773,N_21581);
nor U22067 (N_22067,N_21734,N_21635);
nor U22068 (N_22068,N_21787,N_21741);
and U22069 (N_22069,N_21879,N_21618);
and U22070 (N_22070,N_21801,N_21946);
nor U22071 (N_22071,N_21501,N_21621);
or U22072 (N_22072,N_21658,N_21909);
nand U22073 (N_22073,N_21972,N_21899);
nand U22074 (N_22074,N_21916,N_21607);
nor U22075 (N_22075,N_21963,N_21802);
and U22076 (N_22076,N_21559,N_21640);
or U22077 (N_22077,N_21659,N_21908);
and U22078 (N_22078,N_21970,N_21580);
xor U22079 (N_22079,N_21936,N_21666);
xnor U22080 (N_22080,N_21798,N_21631);
nand U22081 (N_22081,N_21918,N_21886);
xor U22082 (N_22082,N_21923,N_21516);
and U22083 (N_22083,N_21547,N_21874);
xnor U22084 (N_22084,N_21737,N_21529);
or U22085 (N_22085,N_21903,N_21863);
xor U22086 (N_22086,N_21954,N_21575);
xnor U22087 (N_22087,N_21673,N_21785);
xor U22088 (N_22088,N_21515,N_21625);
and U22089 (N_22089,N_21776,N_21652);
xnor U22090 (N_22090,N_21591,N_21597);
nor U22091 (N_22091,N_21921,N_21504);
nor U22092 (N_22092,N_21567,N_21703);
and U22093 (N_22093,N_21670,N_21997);
and U22094 (N_22094,N_21929,N_21792);
xnor U22095 (N_22095,N_21933,N_21582);
or U22096 (N_22096,N_21842,N_21624);
and U22097 (N_22097,N_21805,N_21944);
nor U22098 (N_22098,N_21556,N_21945);
xor U22099 (N_22099,N_21894,N_21937);
nand U22100 (N_22100,N_21630,N_21610);
xor U22101 (N_22101,N_21869,N_21612);
xnor U22102 (N_22102,N_21781,N_21605);
nand U22103 (N_22103,N_21533,N_21907);
xnor U22104 (N_22104,N_21808,N_21711);
and U22105 (N_22105,N_21619,N_21783);
or U22106 (N_22106,N_21796,N_21634);
nand U22107 (N_22107,N_21513,N_21868);
and U22108 (N_22108,N_21822,N_21667);
or U22109 (N_22109,N_21767,N_21789);
nor U22110 (N_22110,N_21510,N_21526);
or U22111 (N_22111,N_21598,N_21739);
or U22112 (N_22112,N_21828,N_21756);
nand U22113 (N_22113,N_21617,N_21714);
nor U22114 (N_22114,N_21506,N_21875);
and U22115 (N_22115,N_21943,N_21709);
or U22116 (N_22116,N_21791,N_21985);
and U22117 (N_22117,N_21880,N_21539);
and U22118 (N_22118,N_21601,N_21536);
xnor U22119 (N_22119,N_21852,N_21834);
nand U22120 (N_22120,N_21724,N_21952);
xor U22121 (N_22121,N_21704,N_21817);
or U22122 (N_22122,N_21771,N_21964);
nor U22123 (N_22123,N_21522,N_21941);
nor U22124 (N_22124,N_21554,N_21716);
nor U22125 (N_22125,N_21550,N_21803);
and U22126 (N_22126,N_21759,N_21979);
and U22127 (N_22127,N_21602,N_21780);
and U22128 (N_22128,N_21511,N_21764);
nand U22129 (N_22129,N_21671,N_21538);
or U22130 (N_22130,N_21813,N_21959);
or U22131 (N_22131,N_21977,N_21578);
nor U22132 (N_22132,N_21955,N_21973);
nand U22133 (N_22133,N_21717,N_21646);
nor U22134 (N_22134,N_21762,N_21999);
nor U22135 (N_22135,N_21958,N_21728);
nor U22136 (N_22136,N_21681,N_21821);
nand U22137 (N_22137,N_21850,N_21685);
nand U22138 (N_22138,N_21915,N_21695);
or U22139 (N_22139,N_21514,N_21948);
xnor U22140 (N_22140,N_21969,N_21653);
or U22141 (N_22141,N_21881,N_21562);
nand U22142 (N_22142,N_21924,N_21865);
nor U22143 (N_22143,N_21815,N_21926);
and U22144 (N_22144,N_21611,N_21691);
nor U22145 (N_22145,N_21661,N_21632);
or U22146 (N_22146,N_21665,N_21810);
and U22147 (N_22147,N_21811,N_21818);
xnor U22148 (N_22148,N_21814,N_21540);
nor U22149 (N_22149,N_21790,N_21896);
and U22150 (N_22150,N_21947,N_21657);
xnor U22151 (N_22151,N_21557,N_21535);
xnor U22152 (N_22152,N_21935,N_21521);
nand U22153 (N_22153,N_21641,N_21564);
nand U22154 (N_22154,N_21676,N_21862);
or U22155 (N_22155,N_21687,N_21831);
or U22156 (N_22156,N_21766,N_21827);
xor U22157 (N_22157,N_21991,N_21806);
nand U22158 (N_22158,N_21793,N_21940);
nor U22159 (N_22159,N_21849,N_21572);
and U22160 (N_22160,N_21809,N_21620);
nand U22161 (N_22161,N_21844,N_21545);
xnor U22162 (N_22162,N_21911,N_21897);
or U22163 (N_22163,N_21845,N_21690);
and U22164 (N_22164,N_21747,N_21934);
nor U22165 (N_22165,N_21889,N_21992);
xor U22166 (N_22166,N_21507,N_21830);
or U22167 (N_22167,N_21675,N_21829);
nor U22168 (N_22168,N_21668,N_21528);
nand U22169 (N_22169,N_21832,N_21931);
nand U22170 (N_22170,N_21505,N_21622);
nor U22171 (N_22171,N_21950,N_21727);
xnor U22172 (N_22172,N_21871,N_21971);
and U22173 (N_22173,N_21684,N_21740);
nand U22174 (N_22174,N_21669,N_21523);
and U22175 (N_22175,N_21919,N_21502);
nor U22176 (N_22176,N_21770,N_21887);
nand U22177 (N_22177,N_21738,N_21839);
and U22178 (N_22178,N_21723,N_21733);
nand U22179 (N_22179,N_21649,N_21856);
and U22180 (N_22180,N_21707,N_21900);
xnor U22181 (N_22181,N_21976,N_21980);
and U22182 (N_22182,N_21966,N_21882);
nor U22183 (N_22183,N_21860,N_21509);
xor U22184 (N_22184,N_21837,N_21643);
nand U22185 (N_22185,N_21700,N_21901);
xor U22186 (N_22186,N_21768,N_21891);
nand U22187 (N_22187,N_21596,N_21751);
and U22188 (N_22188,N_21587,N_21906);
nand U22189 (N_22189,N_21551,N_21920);
nand U22190 (N_22190,N_21721,N_21592);
xor U22191 (N_22191,N_21651,N_21981);
nand U22192 (N_22192,N_21637,N_21519);
xor U22193 (N_22193,N_21993,N_21960);
nand U22194 (N_22194,N_21672,N_21688);
xor U22195 (N_22195,N_21942,N_21642);
xnor U22196 (N_22196,N_21698,N_21561);
xor U22197 (N_22197,N_21854,N_21736);
or U22198 (N_22198,N_21895,N_21569);
or U22199 (N_22199,N_21995,N_21835);
or U22200 (N_22200,N_21847,N_21912);
nor U22201 (N_22201,N_21825,N_21576);
or U22202 (N_22202,N_21588,N_21876);
nor U22203 (N_22203,N_21560,N_21927);
and U22204 (N_22204,N_21967,N_21998);
nor U22205 (N_22205,N_21629,N_21851);
or U22206 (N_22206,N_21804,N_21713);
and U22207 (N_22207,N_21917,N_21693);
nor U22208 (N_22208,N_21720,N_21859);
xor U22209 (N_22209,N_21708,N_21816);
nand U22210 (N_22210,N_21961,N_21520);
nor U22211 (N_22211,N_21786,N_21877);
xor U22212 (N_22212,N_21586,N_21571);
nand U22213 (N_22213,N_21807,N_21623);
or U22214 (N_22214,N_21573,N_21748);
nand U22215 (N_22215,N_21585,N_21701);
or U22216 (N_22216,N_21705,N_21583);
and U22217 (N_22217,N_21812,N_21735);
xor U22218 (N_22218,N_21902,N_21603);
xor U22219 (N_22219,N_21823,N_21841);
nor U22220 (N_22220,N_21870,N_21951);
xnor U22221 (N_22221,N_21565,N_21775);
or U22222 (N_22222,N_21650,N_21662);
xor U22223 (N_22223,N_21968,N_21699);
or U22224 (N_22224,N_21753,N_21674);
nand U22225 (N_22225,N_21645,N_21988);
nor U22226 (N_22226,N_21848,N_21836);
nor U22227 (N_22227,N_21664,N_21517);
xnor U22228 (N_22228,N_21846,N_21689);
nor U22229 (N_22229,N_21710,N_21794);
and U22230 (N_22230,N_21544,N_21590);
or U22231 (N_22231,N_21694,N_21706);
nand U22232 (N_22232,N_21568,N_21606);
xor U22233 (N_22233,N_21744,N_21574);
or U22234 (N_22234,N_21696,N_21677);
and U22235 (N_22235,N_21532,N_21742);
and U22236 (N_22236,N_21826,N_21660);
nor U22237 (N_22237,N_21978,N_21888);
xor U22238 (N_22238,N_21938,N_21840);
nand U22239 (N_22239,N_21589,N_21563);
xor U22240 (N_22240,N_21982,N_21914);
xnor U22241 (N_22241,N_21782,N_21983);
and U22242 (N_22242,N_21930,N_21754);
nand U22243 (N_22243,N_21570,N_21613);
or U22244 (N_22244,N_21996,N_21525);
nor U22245 (N_22245,N_21615,N_21892);
nor U22246 (N_22246,N_21639,N_21866);
nor U22247 (N_22247,N_21784,N_21663);
xnor U22248 (N_22248,N_21518,N_21956);
or U22249 (N_22249,N_21712,N_21765);
and U22250 (N_22250,N_21789,N_21970);
nor U22251 (N_22251,N_21979,N_21726);
or U22252 (N_22252,N_21643,N_21845);
nor U22253 (N_22253,N_21911,N_21865);
xor U22254 (N_22254,N_21665,N_21823);
or U22255 (N_22255,N_21640,N_21703);
or U22256 (N_22256,N_21713,N_21505);
and U22257 (N_22257,N_21516,N_21795);
xor U22258 (N_22258,N_21627,N_21611);
and U22259 (N_22259,N_21619,N_21760);
and U22260 (N_22260,N_21631,N_21891);
nor U22261 (N_22261,N_21561,N_21515);
nand U22262 (N_22262,N_21686,N_21940);
nor U22263 (N_22263,N_21838,N_21973);
and U22264 (N_22264,N_21522,N_21600);
or U22265 (N_22265,N_21583,N_21928);
nand U22266 (N_22266,N_21915,N_21858);
or U22267 (N_22267,N_21852,N_21792);
and U22268 (N_22268,N_21617,N_21978);
or U22269 (N_22269,N_21623,N_21898);
and U22270 (N_22270,N_21743,N_21880);
and U22271 (N_22271,N_21942,N_21798);
and U22272 (N_22272,N_21965,N_21769);
and U22273 (N_22273,N_21776,N_21802);
nand U22274 (N_22274,N_21753,N_21836);
nor U22275 (N_22275,N_21696,N_21738);
and U22276 (N_22276,N_21710,N_21648);
or U22277 (N_22277,N_21533,N_21683);
nand U22278 (N_22278,N_21819,N_21689);
nand U22279 (N_22279,N_21814,N_21654);
nand U22280 (N_22280,N_21906,N_21633);
and U22281 (N_22281,N_21965,N_21598);
nand U22282 (N_22282,N_21519,N_21895);
nand U22283 (N_22283,N_21904,N_21955);
and U22284 (N_22284,N_21662,N_21689);
or U22285 (N_22285,N_21857,N_21946);
nand U22286 (N_22286,N_21517,N_21566);
and U22287 (N_22287,N_21639,N_21640);
or U22288 (N_22288,N_21911,N_21517);
and U22289 (N_22289,N_21959,N_21624);
nor U22290 (N_22290,N_21582,N_21809);
and U22291 (N_22291,N_21991,N_21846);
nor U22292 (N_22292,N_21798,N_21591);
xnor U22293 (N_22293,N_21524,N_21864);
or U22294 (N_22294,N_21554,N_21544);
nor U22295 (N_22295,N_21835,N_21578);
and U22296 (N_22296,N_21525,N_21920);
or U22297 (N_22297,N_21661,N_21801);
nor U22298 (N_22298,N_21939,N_21701);
and U22299 (N_22299,N_21813,N_21926);
xnor U22300 (N_22300,N_21661,N_21980);
or U22301 (N_22301,N_21590,N_21862);
nand U22302 (N_22302,N_21743,N_21613);
or U22303 (N_22303,N_21868,N_21574);
nand U22304 (N_22304,N_21971,N_21834);
and U22305 (N_22305,N_21774,N_21727);
nand U22306 (N_22306,N_21988,N_21598);
nand U22307 (N_22307,N_21848,N_21785);
or U22308 (N_22308,N_21629,N_21812);
and U22309 (N_22309,N_21624,N_21699);
xor U22310 (N_22310,N_21972,N_21778);
or U22311 (N_22311,N_21721,N_21666);
or U22312 (N_22312,N_21643,N_21977);
nor U22313 (N_22313,N_21754,N_21914);
xnor U22314 (N_22314,N_21572,N_21788);
and U22315 (N_22315,N_21894,N_21625);
xor U22316 (N_22316,N_21720,N_21925);
xor U22317 (N_22317,N_21994,N_21609);
and U22318 (N_22318,N_21701,N_21512);
nor U22319 (N_22319,N_21955,N_21978);
xnor U22320 (N_22320,N_21682,N_21950);
nor U22321 (N_22321,N_21931,N_21760);
and U22322 (N_22322,N_21751,N_21738);
xnor U22323 (N_22323,N_21806,N_21832);
and U22324 (N_22324,N_21817,N_21678);
and U22325 (N_22325,N_21930,N_21779);
and U22326 (N_22326,N_21676,N_21834);
and U22327 (N_22327,N_21733,N_21666);
or U22328 (N_22328,N_21739,N_21771);
nand U22329 (N_22329,N_21650,N_21747);
xnor U22330 (N_22330,N_21646,N_21980);
or U22331 (N_22331,N_21579,N_21680);
or U22332 (N_22332,N_21621,N_21715);
xor U22333 (N_22333,N_21876,N_21556);
xor U22334 (N_22334,N_21626,N_21568);
and U22335 (N_22335,N_21810,N_21514);
xnor U22336 (N_22336,N_21517,N_21615);
or U22337 (N_22337,N_21768,N_21631);
and U22338 (N_22338,N_21801,N_21554);
nor U22339 (N_22339,N_21596,N_21790);
xor U22340 (N_22340,N_21764,N_21959);
or U22341 (N_22341,N_21520,N_21869);
or U22342 (N_22342,N_21813,N_21762);
and U22343 (N_22343,N_21785,N_21786);
and U22344 (N_22344,N_21839,N_21773);
xor U22345 (N_22345,N_21570,N_21982);
nor U22346 (N_22346,N_21586,N_21605);
xor U22347 (N_22347,N_21850,N_21814);
xor U22348 (N_22348,N_21927,N_21711);
or U22349 (N_22349,N_21807,N_21570);
xnor U22350 (N_22350,N_21713,N_21802);
nand U22351 (N_22351,N_21734,N_21584);
nor U22352 (N_22352,N_21505,N_21978);
nor U22353 (N_22353,N_21583,N_21959);
or U22354 (N_22354,N_21650,N_21835);
and U22355 (N_22355,N_21651,N_21753);
or U22356 (N_22356,N_21777,N_21632);
or U22357 (N_22357,N_21637,N_21771);
xor U22358 (N_22358,N_21800,N_21590);
xor U22359 (N_22359,N_21995,N_21537);
xor U22360 (N_22360,N_21924,N_21991);
or U22361 (N_22361,N_21556,N_21824);
nand U22362 (N_22362,N_21944,N_21751);
xor U22363 (N_22363,N_21718,N_21636);
and U22364 (N_22364,N_21986,N_21915);
xor U22365 (N_22365,N_21650,N_21699);
nor U22366 (N_22366,N_21584,N_21842);
and U22367 (N_22367,N_21750,N_21902);
nor U22368 (N_22368,N_21758,N_21939);
xor U22369 (N_22369,N_21545,N_21624);
nand U22370 (N_22370,N_21692,N_21674);
or U22371 (N_22371,N_21758,N_21789);
nor U22372 (N_22372,N_21938,N_21714);
and U22373 (N_22373,N_21755,N_21504);
nor U22374 (N_22374,N_21864,N_21572);
or U22375 (N_22375,N_21730,N_21997);
xor U22376 (N_22376,N_21571,N_21684);
nor U22377 (N_22377,N_21813,N_21534);
nand U22378 (N_22378,N_21889,N_21620);
nand U22379 (N_22379,N_21813,N_21934);
xnor U22380 (N_22380,N_21735,N_21907);
or U22381 (N_22381,N_21629,N_21525);
nor U22382 (N_22382,N_21656,N_21549);
xnor U22383 (N_22383,N_21617,N_21719);
xor U22384 (N_22384,N_21921,N_21806);
nand U22385 (N_22385,N_21924,N_21814);
or U22386 (N_22386,N_21991,N_21810);
nand U22387 (N_22387,N_21683,N_21926);
and U22388 (N_22388,N_21941,N_21945);
and U22389 (N_22389,N_21869,N_21582);
nor U22390 (N_22390,N_21897,N_21600);
nand U22391 (N_22391,N_21871,N_21593);
xnor U22392 (N_22392,N_21770,N_21728);
nand U22393 (N_22393,N_21517,N_21955);
nor U22394 (N_22394,N_21840,N_21717);
xnor U22395 (N_22395,N_21511,N_21640);
xor U22396 (N_22396,N_21690,N_21895);
xnor U22397 (N_22397,N_21811,N_21676);
and U22398 (N_22398,N_21884,N_21942);
or U22399 (N_22399,N_21697,N_21639);
xnor U22400 (N_22400,N_21583,N_21906);
nor U22401 (N_22401,N_21733,N_21790);
and U22402 (N_22402,N_21617,N_21759);
nor U22403 (N_22403,N_21880,N_21611);
nand U22404 (N_22404,N_21930,N_21659);
xnor U22405 (N_22405,N_21559,N_21805);
and U22406 (N_22406,N_21920,N_21846);
xnor U22407 (N_22407,N_21589,N_21995);
nand U22408 (N_22408,N_21554,N_21515);
nor U22409 (N_22409,N_21515,N_21726);
xor U22410 (N_22410,N_21675,N_21857);
and U22411 (N_22411,N_21858,N_21614);
nand U22412 (N_22412,N_21610,N_21536);
or U22413 (N_22413,N_21694,N_21582);
or U22414 (N_22414,N_21942,N_21819);
and U22415 (N_22415,N_21889,N_21663);
nand U22416 (N_22416,N_21861,N_21774);
and U22417 (N_22417,N_21963,N_21732);
nor U22418 (N_22418,N_21535,N_21608);
nor U22419 (N_22419,N_21627,N_21911);
nand U22420 (N_22420,N_21638,N_21792);
or U22421 (N_22421,N_21621,N_21699);
xor U22422 (N_22422,N_21662,N_21989);
xnor U22423 (N_22423,N_21533,N_21666);
or U22424 (N_22424,N_21616,N_21940);
nor U22425 (N_22425,N_21619,N_21506);
nor U22426 (N_22426,N_21881,N_21974);
or U22427 (N_22427,N_21841,N_21762);
or U22428 (N_22428,N_21551,N_21942);
xor U22429 (N_22429,N_21940,N_21906);
nand U22430 (N_22430,N_21942,N_21684);
xnor U22431 (N_22431,N_21573,N_21934);
and U22432 (N_22432,N_21814,N_21527);
or U22433 (N_22433,N_21637,N_21860);
or U22434 (N_22434,N_21909,N_21778);
nor U22435 (N_22435,N_21521,N_21563);
nand U22436 (N_22436,N_21927,N_21912);
xor U22437 (N_22437,N_21626,N_21671);
or U22438 (N_22438,N_21984,N_21981);
or U22439 (N_22439,N_21953,N_21620);
xnor U22440 (N_22440,N_21836,N_21742);
nor U22441 (N_22441,N_21590,N_21553);
xnor U22442 (N_22442,N_21943,N_21693);
or U22443 (N_22443,N_21661,N_21887);
nand U22444 (N_22444,N_21771,N_21721);
and U22445 (N_22445,N_21811,N_21549);
xor U22446 (N_22446,N_21679,N_21843);
nor U22447 (N_22447,N_21803,N_21768);
xor U22448 (N_22448,N_21543,N_21937);
xor U22449 (N_22449,N_21942,N_21858);
nor U22450 (N_22450,N_21864,N_21700);
xor U22451 (N_22451,N_21902,N_21821);
nand U22452 (N_22452,N_21658,N_21712);
nor U22453 (N_22453,N_21590,N_21947);
xnor U22454 (N_22454,N_21954,N_21970);
or U22455 (N_22455,N_21789,N_21582);
and U22456 (N_22456,N_21620,N_21927);
or U22457 (N_22457,N_21868,N_21565);
nand U22458 (N_22458,N_21864,N_21547);
xnor U22459 (N_22459,N_21905,N_21584);
and U22460 (N_22460,N_21526,N_21578);
nand U22461 (N_22461,N_21806,N_21624);
nand U22462 (N_22462,N_21760,N_21633);
and U22463 (N_22463,N_21590,N_21914);
xor U22464 (N_22464,N_21982,N_21636);
xnor U22465 (N_22465,N_21647,N_21917);
or U22466 (N_22466,N_21739,N_21644);
or U22467 (N_22467,N_21905,N_21825);
nand U22468 (N_22468,N_21589,N_21706);
and U22469 (N_22469,N_21920,N_21910);
nor U22470 (N_22470,N_21911,N_21921);
xnor U22471 (N_22471,N_21688,N_21616);
nor U22472 (N_22472,N_21747,N_21704);
nor U22473 (N_22473,N_21766,N_21851);
or U22474 (N_22474,N_21682,N_21942);
and U22475 (N_22475,N_21763,N_21604);
or U22476 (N_22476,N_21834,N_21942);
nand U22477 (N_22477,N_21652,N_21708);
nand U22478 (N_22478,N_21573,N_21855);
xnor U22479 (N_22479,N_21942,N_21900);
nor U22480 (N_22480,N_21811,N_21581);
and U22481 (N_22481,N_21934,N_21703);
xor U22482 (N_22482,N_21951,N_21665);
nand U22483 (N_22483,N_21849,N_21786);
nand U22484 (N_22484,N_21688,N_21644);
or U22485 (N_22485,N_21960,N_21823);
and U22486 (N_22486,N_21583,N_21514);
nor U22487 (N_22487,N_21621,N_21645);
xnor U22488 (N_22488,N_21630,N_21745);
xor U22489 (N_22489,N_21780,N_21966);
xnor U22490 (N_22490,N_21826,N_21546);
xor U22491 (N_22491,N_21667,N_21634);
and U22492 (N_22492,N_21555,N_21755);
or U22493 (N_22493,N_21640,N_21861);
or U22494 (N_22494,N_21994,N_21990);
and U22495 (N_22495,N_21806,N_21973);
and U22496 (N_22496,N_21820,N_21932);
and U22497 (N_22497,N_21921,N_21874);
nor U22498 (N_22498,N_21756,N_21970);
or U22499 (N_22499,N_21858,N_21645);
nand U22500 (N_22500,N_22280,N_22107);
xnor U22501 (N_22501,N_22172,N_22297);
nand U22502 (N_22502,N_22205,N_22047);
xor U22503 (N_22503,N_22129,N_22215);
xnor U22504 (N_22504,N_22373,N_22268);
nand U22505 (N_22505,N_22244,N_22034);
nor U22506 (N_22506,N_22206,N_22353);
and U22507 (N_22507,N_22396,N_22236);
and U22508 (N_22508,N_22196,N_22421);
nor U22509 (N_22509,N_22256,N_22246);
xnor U22510 (N_22510,N_22477,N_22352);
nor U22511 (N_22511,N_22490,N_22162);
or U22512 (N_22512,N_22436,N_22422);
or U22513 (N_22513,N_22454,N_22405);
nand U22514 (N_22514,N_22263,N_22251);
or U22515 (N_22515,N_22186,N_22014);
and U22516 (N_22516,N_22059,N_22189);
xnor U22517 (N_22517,N_22223,N_22281);
xnor U22518 (N_22518,N_22293,N_22326);
nor U22519 (N_22519,N_22082,N_22394);
and U22520 (N_22520,N_22357,N_22228);
nor U22521 (N_22521,N_22245,N_22419);
nor U22522 (N_22522,N_22027,N_22305);
nand U22523 (N_22523,N_22482,N_22213);
and U22524 (N_22524,N_22457,N_22290);
xor U22525 (N_22525,N_22323,N_22267);
or U22526 (N_22526,N_22208,N_22310);
nand U22527 (N_22527,N_22056,N_22226);
nor U22528 (N_22528,N_22171,N_22092);
and U22529 (N_22529,N_22065,N_22271);
nor U22530 (N_22530,N_22466,N_22155);
nor U22531 (N_22531,N_22434,N_22319);
and U22532 (N_22532,N_22403,N_22349);
nand U22533 (N_22533,N_22242,N_22337);
or U22534 (N_22534,N_22187,N_22386);
and U22535 (N_22535,N_22125,N_22317);
nor U22536 (N_22536,N_22356,N_22073);
nand U22537 (N_22537,N_22083,N_22203);
or U22538 (N_22538,N_22066,N_22266);
xor U22539 (N_22539,N_22391,N_22063);
nand U22540 (N_22540,N_22057,N_22328);
nor U22541 (N_22541,N_22389,N_22276);
and U22542 (N_22542,N_22440,N_22109);
xnor U22543 (N_22543,N_22269,N_22295);
and U22544 (N_22544,N_22433,N_22111);
xnor U22545 (N_22545,N_22130,N_22494);
nand U22546 (N_22546,N_22167,N_22114);
xnor U22547 (N_22547,N_22332,N_22387);
xnor U22548 (N_22548,N_22483,N_22224);
and U22549 (N_22549,N_22374,N_22370);
and U22550 (N_22550,N_22103,N_22115);
xnor U22551 (N_22551,N_22153,N_22431);
and U22552 (N_22552,N_22447,N_22443);
xor U22553 (N_22553,N_22141,N_22442);
and U22554 (N_22554,N_22424,N_22283);
xnor U22555 (N_22555,N_22000,N_22498);
xnor U22556 (N_22556,N_22464,N_22197);
nand U22557 (N_22557,N_22050,N_22428);
nand U22558 (N_22558,N_22481,N_22361);
nor U22559 (N_22559,N_22028,N_22079);
or U22560 (N_22560,N_22099,N_22437);
and U22561 (N_22561,N_22045,N_22468);
nand U22562 (N_22562,N_22253,N_22488);
nor U22563 (N_22563,N_22329,N_22016);
xor U22564 (N_22564,N_22358,N_22462);
xor U22565 (N_22565,N_22006,N_22030);
or U22566 (N_22566,N_22146,N_22401);
nand U22567 (N_22567,N_22062,N_22429);
or U22568 (N_22568,N_22199,N_22087);
nor U22569 (N_22569,N_22288,N_22085);
nand U22570 (N_22570,N_22330,N_22138);
and U22571 (N_22571,N_22160,N_22119);
xnor U22572 (N_22572,N_22384,N_22300);
nor U22573 (N_22573,N_22142,N_22051);
nor U22574 (N_22574,N_22225,N_22315);
nor U22575 (N_22575,N_22219,N_22489);
or U22576 (N_22576,N_22425,N_22423);
xor U22577 (N_22577,N_22096,N_22347);
xnor U22578 (N_22578,N_22108,N_22390);
and U22579 (N_22579,N_22333,N_22180);
nor U22580 (N_22580,N_22380,N_22453);
and U22581 (N_22581,N_22472,N_22009);
nor U22582 (N_22582,N_22227,N_22249);
xnor U22583 (N_22583,N_22217,N_22089);
xnor U22584 (N_22584,N_22459,N_22334);
nor U22585 (N_22585,N_22412,N_22248);
xor U22586 (N_22586,N_22194,N_22005);
or U22587 (N_22587,N_22133,N_22233);
or U22588 (N_22588,N_22392,N_22220);
nor U22589 (N_22589,N_22169,N_22298);
or U22590 (N_22590,N_22214,N_22134);
xnor U22591 (N_22591,N_22452,N_22418);
nor U22592 (N_22592,N_22259,N_22366);
xnor U22593 (N_22593,N_22140,N_22346);
nand U22594 (N_22594,N_22149,N_22152);
nor U22595 (N_22595,N_22232,N_22094);
nand U22596 (N_22596,N_22025,N_22309);
nor U22597 (N_22597,N_22487,N_22148);
nor U22598 (N_22598,N_22032,N_22081);
and U22599 (N_22599,N_22299,N_22467);
nand U22600 (N_22600,N_22164,N_22112);
nor U22601 (N_22601,N_22053,N_22052);
and U22602 (N_22602,N_22035,N_22174);
nand U22603 (N_22603,N_22382,N_22465);
nand U22604 (N_22604,N_22026,N_22480);
xnor U22605 (N_22605,N_22350,N_22291);
xnor U22606 (N_22606,N_22024,N_22126);
nor U22607 (N_22607,N_22470,N_22069);
and U22608 (N_22608,N_22077,N_22496);
and U22609 (N_22609,N_22143,N_22183);
nor U22610 (N_22610,N_22284,N_22327);
nand U22611 (N_22611,N_22438,N_22408);
nand U22612 (N_22612,N_22414,N_22354);
nand U22613 (N_22613,N_22285,N_22071);
nor U22614 (N_22614,N_22445,N_22398);
xor U22615 (N_22615,N_22158,N_22411);
nand U22616 (N_22616,N_22397,N_22216);
xnor U22617 (N_22617,N_22257,N_22102);
or U22618 (N_22618,N_22039,N_22406);
xnor U22619 (N_22619,N_22145,N_22209);
or U22620 (N_22620,N_22336,N_22105);
and U22621 (N_22621,N_22198,N_22002);
xor U22622 (N_22622,N_22369,N_22313);
and U22623 (N_22623,N_22365,N_22368);
and U22624 (N_22624,N_22469,N_22170);
nor U22625 (N_22625,N_22168,N_22388);
or U22626 (N_22626,N_22478,N_22495);
xnor U22627 (N_22627,N_22076,N_22161);
and U22628 (N_22628,N_22007,N_22234);
or U22629 (N_22629,N_22262,N_22113);
or U22630 (N_22630,N_22318,N_22131);
xnor U22631 (N_22631,N_22497,N_22020);
nand U22632 (N_22632,N_22360,N_22275);
nand U22633 (N_22633,N_22463,N_22011);
nor U22634 (N_22634,N_22314,N_22378);
nor U22635 (N_22635,N_22230,N_22157);
and U22636 (N_22636,N_22118,N_22018);
and U22637 (N_22637,N_22448,N_22181);
xor U22638 (N_22638,N_22088,N_22240);
nand U22639 (N_22639,N_22279,N_22312);
xnor U22640 (N_22640,N_22250,N_22338);
or U22641 (N_22641,N_22342,N_22311);
nand U22642 (N_22642,N_22254,N_22121);
nand U22643 (N_22643,N_22235,N_22021);
xor U22644 (N_22644,N_22010,N_22258);
xnor U22645 (N_22645,N_22413,N_22446);
xnor U22646 (N_22646,N_22093,N_22286);
or U22647 (N_22647,N_22407,N_22191);
nor U22648 (N_22648,N_22450,N_22416);
nand U22649 (N_22649,N_22175,N_22362);
xor U22650 (N_22650,N_22132,N_22098);
nor U22651 (N_22651,N_22106,N_22184);
or U22652 (N_22652,N_22067,N_22041);
xor U22653 (N_22653,N_22128,N_22383);
xnor U22654 (N_22654,N_22212,N_22304);
nor U22655 (N_22655,N_22427,N_22479);
nor U22656 (N_22656,N_22135,N_22409);
xor U22657 (N_22657,N_22320,N_22202);
xnor U22658 (N_22658,N_22054,N_22072);
or U22659 (N_22659,N_22375,N_22159);
xor U22660 (N_22660,N_22377,N_22019);
xnor U22661 (N_22661,N_22151,N_22474);
and U22662 (N_22662,N_22272,N_22255);
nor U22663 (N_22663,N_22325,N_22176);
xor U22664 (N_22664,N_22110,N_22044);
and U22665 (N_22665,N_22473,N_22402);
nand U22666 (N_22666,N_22068,N_22435);
and U22667 (N_22667,N_22306,N_22100);
nor U22668 (N_22668,N_22185,N_22229);
nand U22669 (N_22669,N_22265,N_22475);
xnor U22670 (N_22670,N_22441,N_22393);
and U22671 (N_22671,N_22033,N_22493);
or U22672 (N_22672,N_22351,N_22173);
nor U22673 (N_22673,N_22136,N_22061);
xnor U22674 (N_22674,N_22117,N_22410);
and U22675 (N_22675,N_22322,N_22289);
and U22676 (N_22676,N_22339,N_22417);
nor U22677 (N_22677,N_22379,N_22355);
xor U22678 (N_22678,N_22335,N_22123);
or U22679 (N_22679,N_22070,N_22432);
nand U22680 (N_22680,N_22292,N_22080);
nor U22681 (N_22681,N_22426,N_22177);
and U22682 (N_22682,N_22367,N_22461);
and U22683 (N_22683,N_22456,N_22296);
xor U22684 (N_22684,N_22239,N_22144);
nor U22685 (N_22685,N_22097,N_22003);
xnor U22686 (N_22686,N_22178,N_22179);
or U22687 (N_22687,N_22091,N_22455);
xnor U22688 (N_22688,N_22400,N_22211);
nand U22689 (N_22689,N_22243,N_22486);
or U22690 (N_22690,N_22444,N_22252);
or U22691 (N_22691,N_22031,N_22491);
or U22692 (N_22692,N_22261,N_22122);
nor U22693 (N_22693,N_22078,N_22307);
nor U22694 (N_22694,N_22287,N_22359);
and U22695 (N_22695,N_22075,N_22451);
and U22696 (N_22696,N_22210,N_22017);
and U22697 (N_22697,N_22404,N_22192);
and U22698 (N_22698,N_22060,N_22104);
or U22699 (N_22699,N_22193,N_22348);
and U22700 (N_22700,N_22415,N_22471);
nand U22701 (N_22701,N_22013,N_22023);
xor U22702 (N_22702,N_22001,N_22036);
and U22703 (N_22703,N_22127,N_22086);
nand U22704 (N_22704,N_22420,N_22458);
and U22705 (N_22705,N_22043,N_22221);
xor U22706 (N_22706,N_22247,N_22015);
nor U22707 (N_22707,N_22237,N_22278);
and U22708 (N_22708,N_22163,N_22165);
or U22709 (N_22709,N_22218,N_22485);
xor U22710 (N_22710,N_22084,N_22090);
nand U22711 (N_22711,N_22124,N_22316);
nor U22712 (N_22712,N_22207,N_22046);
xor U22713 (N_22713,N_22166,N_22190);
or U22714 (N_22714,N_22260,N_22302);
nand U22715 (N_22715,N_22345,N_22188);
xor U22716 (N_22716,N_22344,N_22200);
nor U22717 (N_22717,N_22116,N_22154);
xor U22718 (N_22718,N_22231,N_22301);
and U22719 (N_22719,N_22004,N_22241);
or U22720 (N_22720,N_22273,N_22147);
nor U22721 (N_22721,N_22363,N_22395);
xor U22722 (N_22722,N_22238,N_22195);
xor U22723 (N_22723,N_22042,N_22282);
xor U22724 (N_22724,N_22476,N_22055);
xnor U22725 (N_22725,N_22182,N_22012);
or U22726 (N_22726,N_22294,N_22499);
or U22727 (N_22727,N_22364,N_22058);
or U22728 (N_22728,N_22049,N_22201);
or U22729 (N_22729,N_22376,N_22029);
and U22730 (N_22730,N_22460,N_22095);
or U22731 (N_22731,N_22222,N_22139);
or U22732 (N_22732,N_22399,N_22439);
or U22733 (N_22733,N_22277,N_22324);
or U22734 (N_22734,N_22372,N_22204);
xor U22735 (N_22735,N_22038,N_22074);
nor U22736 (N_22736,N_22385,N_22064);
and U22737 (N_22737,N_22101,N_22492);
or U22738 (N_22738,N_22008,N_22340);
and U22739 (N_22739,N_22156,N_22371);
or U22740 (N_22740,N_22270,N_22037);
nor U22741 (N_22741,N_22449,N_22137);
nand U22742 (N_22742,N_22303,N_22381);
nor U22743 (N_22743,N_22120,N_22484);
nand U22744 (N_22744,N_22341,N_22022);
and U22745 (N_22745,N_22343,N_22264);
nand U22746 (N_22746,N_22308,N_22040);
nand U22747 (N_22747,N_22321,N_22150);
xnor U22748 (N_22748,N_22274,N_22331);
nor U22749 (N_22749,N_22430,N_22048);
nand U22750 (N_22750,N_22248,N_22232);
nand U22751 (N_22751,N_22061,N_22303);
nor U22752 (N_22752,N_22410,N_22357);
and U22753 (N_22753,N_22488,N_22275);
xor U22754 (N_22754,N_22408,N_22334);
nor U22755 (N_22755,N_22391,N_22432);
or U22756 (N_22756,N_22116,N_22031);
nand U22757 (N_22757,N_22249,N_22297);
xor U22758 (N_22758,N_22148,N_22378);
xnor U22759 (N_22759,N_22117,N_22030);
or U22760 (N_22760,N_22049,N_22182);
nand U22761 (N_22761,N_22250,N_22397);
or U22762 (N_22762,N_22350,N_22084);
or U22763 (N_22763,N_22150,N_22456);
nand U22764 (N_22764,N_22266,N_22268);
and U22765 (N_22765,N_22230,N_22005);
nand U22766 (N_22766,N_22481,N_22067);
and U22767 (N_22767,N_22336,N_22092);
xnor U22768 (N_22768,N_22396,N_22292);
xor U22769 (N_22769,N_22244,N_22105);
nand U22770 (N_22770,N_22482,N_22030);
nor U22771 (N_22771,N_22107,N_22480);
nand U22772 (N_22772,N_22322,N_22363);
nor U22773 (N_22773,N_22394,N_22157);
nor U22774 (N_22774,N_22335,N_22085);
xnor U22775 (N_22775,N_22302,N_22178);
and U22776 (N_22776,N_22140,N_22199);
or U22777 (N_22777,N_22152,N_22053);
xnor U22778 (N_22778,N_22170,N_22316);
xnor U22779 (N_22779,N_22319,N_22108);
or U22780 (N_22780,N_22303,N_22433);
nand U22781 (N_22781,N_22106,N_22452);
xor U22782 (N_22782,N_22480,N_22163);
xor U22783 (N_22783,N_22423,N_22324);
or U22784 (N_22784,N_22398,N_22415);
and U22785 (N_22785,N_22423,N_22136);
nor U22786 (N_22786,N_22103,N_22383);
and U22787 (N_22787,N_22091,N_22488);
nand U22788 (N_22788,N_22166,N_22415);
nand U22789 (N_22789,N_22077,N_22008);
nor U22790 (N_22790,N_22494,N_22127);
or U22791 (N_22791,N_22374,N_22227);
nand U22792 (N_22792,N_22070,N_22207);
xor U22793 (N_22793,N_22393,N_22483);
xor U22794 (N_22794,N_22410,N_22348);
nand U22795 (N_22795,N_22349,N_22390);
xor U22796 (N_22796,N_22116,N_22323);
or U22797 (N_22797,N_22380,N_22196);
xnor U22798 (N_22798,N_22338,N_22240);
xor U22799 (N_22799,N_22315,N_22453);
or U22800 (N_22800,N_22162,N_22025);
xnor U22801 (N_22801,N_22372,N_22007);
and U22802 (N_22802,N_22438,N_22299);
or U22803 (N_22803,N_22268,N_22077);
nor U22804 (N_22804,N_22032,N_22419);
nor U22805 (N_22805,N_22420,N_22364);
and U22806 (N_22806,N_22174,N_22395);
xor U22807 (N_22807,N_22467,N_22483);
nor U22808 (N_22808,N_22111,N_22117);
nand U22809 (N_22809,N_22321,N_22359);
nor U22810 (N_22810,N_22241,N_22382);
nand U22811 (N_22811,N_22432,N_22169);
xnor U22812 (N_22812,N_22401,N_22134);
or U22813 (N_22813,N_22416,N_22063);
and U22814 (N_22814,N_22030,N_22264);
nor U22815 (N_22815,N_22029,N_22301);
or U22816 (N_22816,N_22229,N_22005);
nor U22817 (N_22817,N_22400,N_22140);
nor U22818 (N_22818,N_22231,N_22452);
nor U22819 (N_22819,N_22129,N_22259);
nand U22820 (N_22820,N_22336,N_22025);
nor U22821 (N_22821,N_22150,N_22381);
and U22822 (N_22822,N_22338,N_22308);
or U22823 (N_22823,N_22419,N_22192);
nand U22824 (N_22824,N_22099,N_22268);
xnor U22825 (N_22825,N_22409,N_22184);
and U22826 (N_22826,N_22000,N_22359);
xnor U22827 (N_22827,N_22157,N_22117);
nor U22828 (N_22828,N_22409,N_22165);
nand U22829 (N_22829,N_22145,N_22162);
or U22830 (N_22830,N_22321,N_22022);
nand U22831 (N_22831,N_22388,N_22461);
and U22832 (N_22832,N_22412,N_22024);
xor U22833 (N_22833,N_22073,N_22089);
nor U22834 (N_22834,N_22203,N_22201);
and U22835 (N_22835,N_22377,N_22352);
and U22836 (N_22836,N_22276,N_22430);
or U22837 (N_22837,N_22410,N_22334);
nor U22838 (N_22838,N_22443,N_22025);
nand U22839 (N_22839,N_22339,N_22311);
and U22840 (N_22840,N_22325,N_22082);
xnor U22841 (N_22841,N_22009,N_22034);
nand U22842 (N_22842,N_22072,N_22262);
nand U22843 (N_22843,N_22040,N_22489);
xnor U22844 (N_22844,N_22464,N_22165);
xor U22845 (N_22845,N_22205,N_22127);
or U22846 (N_22846,N_22052,N_22108);
and U22847 (N_22847,N_22446,N_22231);
xor U22848 (N_22848,N_22292,N_22256);
nand U22849 (N_22849,N_22236,N_22146);
xnor U22850 (N_22850,N_22283,N_22030);
and U22851 (N_22851,N_22193,N_22427);
or U22852 (N_22852,N_22295,N_22275);
xnor U22853 (N_22853,N_22003,N_22442);
nand U22854 (N_22854,N_22231,N_22349);
or U22855 (N_22855,N_22039,N_22414);
nor U22856 (N_22856,N_22433,N_22351);
nand U22857 (N_22857,N_22452,N_22174);
or U22858 (N_22858,N_22324,N_22318);
or U22859 (N_22859,N_22169,N_22311);
nand U22860 (N_22860,N_22336,N_22104);
xnor U22861 (N_22861,N_22448,N_22347);
or U22862 (N_22862,N_22361,N_22226);
nor U22863 (N_22863,N_22308,N_22249);
and U22864 (N_22864,N_22241,N_22216);
nand U22865 (N_22865,N_22139,N_22342);
nor U22866 (N_22866,N_22115,N_22194);
nand U22867 (N_22867,N_22255,N_22381);
or U22868 (N_22868,N_22009,N_22229);
and U22869 (N_22869,N_22076,N_22039);
and U22870 (N_22870,N_22141,N_22405);
xnor U22871 (N_22871,N_22341,N_22329);
nor U22872 (N_22872,N_22343,N_22398);
xnor U22873 (N_22873,N_22441,N_22135);
xor U22874 (N_22874,N_22349,N_22024);
and U22875 (N_22875,N_22091,N_22129);
nand U22876 (N_22876,N_22121,N_22437);
or U22877 (N_22877,N_22383,N_22044);
or U22878 (N_22878,N_22059,N_22342);
or U22879 (N_22879,N_22185,N_22453);
nand U22880 (N_22880,N_22004,N_22412);
xnor U22881 (N_22881,N_22078,N_22154);
or U22882 (N_22882,N_22143,N_22020);
nand U22883 (N_22883,N_22396,N_22448);
or U22884 (N_22884,N_22104,N_22455);
xnor U22885 (N_22885,N_22220,N_22067);
nor U22886 (N_22886,N_22152,N_22269);
and U22887 (N_22887,N_22148,N_22429);
or U22888 (N_22888,N_22210,N_22480);
and U22889 (N_22889,N_22053,N_22156);
and U22890 (N_22890,N_22296,N_22219);
and U22891 (N_22891,N_22472,N_22320);
nand U22892 (N_22892,N_22418,N_22041);
or U22893 (N_22893,N_22261,N_22088);
xor U22894 (N_22894,N_22022,N_22204);
xor U22895 (N_22895,N_22225,N_22231);
nor U22896 (N_22896,N_22283,N_22227);
nor U22897 (N_22897,N_22473,N_22446);
nor U22898 (N_22898,N_22261,N_22325);
and U22899 (N_22899,N_22026,N_22474);
nor U22900 (N_22900,N_22007,N_22221);
xnor U22901 (N_22901,N_22253,N_22302);
xor U22902 (N_22902,N_22283,N_22488);
nand U22903 (N_22903,N_22449,N_22126);
or U22904 (N_22904,N_22159,N_22301);
xor U22905 (N_22905,N_22384,N_22069);
and U22906 (N_22906,N_22329,N_22389);
or U22907 (N_22907,N_22360,N_22185);
nand U22908 (N_22908,N_22115,N_22383);
xor U22909 (N_22909,N_22445,N_22191);
or U22910 (N_22910,N_22478,N_22242);
xnor U22911 (N_22911,N_22355,N_22002);
and U22912 (N_22912,N_22300,N_22311);
and U22913 (N_22913,N_22121,N_22473);
xnor U22914 (N_22914,N_22486,N_22201);
xor U22915 (N_22915,N_22179,N_22164);
nand U22916 (N_22916,N_22365,N_22300);
nand U22917 (N_22917,N_22204,N_22059);
or U22918 (N_22918,N_22054,N_22291);
or U22919 (N_22919,N_22464,N_22019);
and U22920 (N_22920,N_22169,N_22363);
nor U22921 (N_22921,N_22179,N_22494);
nor U22922 (N_22922,N_22349,N_22056);
xnor U22923 (N_22923,N_22032,N_22117);
and U22924 (N_22924,N_22396,N_22002);
nor U22925 (N_22925,N_22020,N_22176);
or U22926 (N_22926,N_22494,N_22496);
or U22927 (N_22927,N_22051,N_22029);
and U22928 (N_22928,N_22047,N_22224);
nand U22929 (N_22929,N_22261,N_22470);
nand U22930 (N_22930,N_22406,N_22017);
and U22931 (N_22931,N_22224,N_22059);
or U22932 (N_22932,N_22211,N_22135);
xnor U22933 (N_22933,N_22170,N_22477);
or U22934 (N_22934,N_22274,N_22330);
or U22935 (N_22935,N_22450,N_22492);
and U22936 (N_22936,N_22455,N_22283);
or U22937 (N_22937,N_22211,N_22086);
or U22938 (N_22938,N_22435,N_22461);
nand U22939 (N_22939,N_22150,N_22347);
nor U22940 (N_22940,N_22415,N_22288);
nor U22941 (N_22941,N_22196,N_22051);
nor U22942 (N_22942,N_22386,N_22167);
nand U22943 (N_22943,N_22400,N_22052);
xnor U22944 (N_22944,N_22215,N_22474);
nor U22945 (N_22945,N_22018,N_22218);
xnor U22946 (N_22946,N_22498,N_22255);
and U22947 (N_22947,N_22414,N_22008);
nor U22948 (N_22948,N_22469,N_22189);
and U22949 (N_22949,N_22109,N_22162);
nand U22950 (N_22950,N_22434,N_22084);
nand U22951 (N_22951,N_22073,N_22411);
xor U22952 (N_22952,N_22474,N_22296);
nor U22953 (N_22953,N_22197,N_22246);
xnor U22954 (N_22954,N_22164,N_22430);
nand U22955 (N_22955,N_22242,N_22450);
and U22956 (N_22956,N_22483,N_22005);
or U22957 (N_22957,N_22068,N_22266);
nand U22958 (N_22958,N_22228,N_22074);
xnor U22959 (N_22959,N_22356,N_22022);
nand U22960 (N_22960,N_22015,N_22212);
or U22961 (N_22961,N_22165,N_22381);
and U22962 (N_22962,N_22405,N_22159);
xnor U22963 (N_22963,N_22450,N_22445);
xor U22964 (N_22964,N_22098,N_22224);
xnor U22965 (N_22965,N_22067,N_22441);
nand U22966 (N_22966,N_22361,N_22427);
or U22967 (N_22967,N_22330,N_22463);
nor U22968 (N_22968,N_22184,N_22070);
and U22969 (N_22969,N_22056,N_22399);
and U22970 (N_22970,N_22421,N_22298);
nand U22971 (N_22971,N_22022,N_22402);
nor U22972 (N_22972,N_22004,N_22490);
and U22973 (N_22973,N_22383,N_22285);
nand U22974 (N_22974,N_22482,N_22331);
nand U22975 (N_22975,N_22360,N_22146);
and U22976 (N_22976,N_22172,N_22280);
nand U22977 (N_22977,N_22181,N_22144);
nor U22978 (N_22978,N_22217,N_22374);
xor U22979 (N_22979,N_22051,N_22373);
and U22980 (N_22980,N_22267,N_22318);
or U22981 (N_22981,N_22189,N_22278);
or U22982 (N_22982,N_22172,N_22398);
or U22983 (N_22983,N_22367,N_22463);
nand U22984 (N_22984,N_22110,N_22193);
or U22985 (N_22985,N_22015,N_22384);
xor U22986 (N_22986,N_22318,N_22130);
and U22987 (N_22987,N_22082,N_22324);
or U22988 (N_22988,N_22415,N_22043);
or U22989 (N_22989,N_22242,N_22228);
nor U22990 (N_22990,N_22263,N_22100);
and U22991 (N_22991,N_22295,N_22239);
and U22992 (N_22992,N_22287,N_22390);
nand U22993 (N_22993,N_22264,N_22480);
and U22994 (N_22994,N_22022,N_22039);
xnor U22995 (N_22995,N_22073,N_22449);
nor U22996 (N_22996,N_22317,N_22354);
nand U22997 (N_22997,N_22411,N_22256);
nor U22998 (N_22998,N_22140,N_22250);
nand U22999 (N_22999,N_22092,N_22370);
or U23000 (N_23000,N_22569,N_22705);
or U23001 (N_23001,N_22619,N_22970);
or U23002 (N_23002,N_22693,N_22969);
and U23003 (N_23003,N_22546,N_22822);
nor U23004 (N_23004,N_22670,N_22857);
and U23005 (N_23005,N_22906,N_22729);
xnor U23006 (N_23006,N_22989,N_22695);
and U23007 (N_23007,N_22897,N_22583);
nor U23008 (N_23008,N_22701,N_22647);
nand U23009 (N_23009,N_22966,N_22743);
xor U23010 (N_23010,N_22870,N_22551);
or U23011 (N_23011,N_22652,N_22615);
and U23012 (N_23012,N_22507,N_22939);
nand U23013 (N_23013,N_22771,N_22642);
nor U23014 (N_23014,N_22678,N_22925);
nand U23015 (N_23015,N_22887,N_22818);
nand U23016 (N_23016,N_22959,N_22867);
or U23017 (N_23017,N_22508,N_22571);
xnor U23018 (N_23018,N_22892,N_22961);
nor U23019 (N_23019,N_22692,N_22839);
and U23020 (N_23020,N_22625,N_22732);
xnor U23021 (N_23021,N_22713,N_22760);
or U23022 (N_23022,N_22525,N_22724);
or U23023 (N_23023,N_22666,N_22778);
nand U23024 (N_23024,N_22862,N_22876);
nor U23025 (N_23025,N_22651,N_22834);
xor U23026 (N_23026,N_22755,N_22850);
nor U23027 (N_23027,N_22528,N_22894);
nor U23028 (N_23028,N_22980,N_22935);
xor U23029 (N_23029,N_22908,N_22503);
nand U23030 (N_23030,N_22677,N_22511);
nor U23031 (N_23031,N_22874,N_22796);
nand U23032 (N_23032,N_22792,N_22880);
xnor U23033 (N_23033,N_22654,N_22981);
xnor U23034 (N_23034,N_22769,N_22685);
nand U23035 (N_23035,N_22593,N_22514);
and U23036 (N_23036,N_22611,N_22888);
or U23037 (N_23037,N_22930,N_22937);
and U23038 (N_23038,N_22648,N_22519);
nor U23039 (N_23039,N_22725,N_22748);
or U23040 (N_23040,N_22534,N_22785);
and U23041 (N_23041,N_22533,N_22814);
nor U23042 (N_23042,N_22557,N_22919);
nand U23043 (N_23043,N_22806,N_22820);
nand U23044 (N_23044,N_22698,N_22837);
xnor U23045 (N_23045,N_22841,N_22764);
xnor U23046 (N_23046,N_22641,N_22548);
nand U23047 (N_23047,N_22621,N_22660);
nand U23048 (N_23048,N_22825,N_22680);
nor U23049 (N_23049,N_22501,N_22911);
and U23050 (N_23050,N_22573,N_22633);
or U23051 (N_23051,N_22632,N_22536);
nor U23052 (N_23052,N_22840,N_22637);
xor U23053 (N_23053,N_22535,N_22909);
or U23054 (N_23054,N_22576,N_22539);
nand U23055 (N_23055,N_22668,N_22815);
nand U23056 (N_23056,N_22864,N_22793);
and U23057 (N_23057,N_22689,N_22927);
nand U23058 (N_23058,N_22738,N_22772);
nand U23059 (N_23059,N_22851,N_22770);
xnor U23060 (N_23060,N_22700,N_22505);
nand U23061 (N_23061,N_22592,N_22631);
nand U23062 (N_23062,N_22962,N_22816);
and U23063 (N_23063,N_22750,N_22926);
or U23064 (N_23064,N_22614,N_22603);
nand U23065 (N_23065,N_22826,N_22996);
or U23066 (N_23066,N_22602,N_22940);
and U23067 (N_23067,N_22762,N_22972);
nor U23068 (N_23068,N_22594,N_22570);
or U23069 (N_23069,N_22575,N_22524);
xor U23070 (N_23070,N_22687,N_22828);
or U23071 (N_23071,N_22671,N_22786);
nor U23072 (N_23072,N_22513,N_22773);
nand U23073 (N_23073,N_22552,N_22601);
or U23074 (N_23074,N_22506,N_22684);
and U23075 (N_23075,N_22907,N_22912);
or U23076 (N_23076,N_22742,N_22986);
nor U23077 (N_23077,N_22577,N_22883);
nand U23078 (N_23078,N_22890,N_22636);
xor U23079 (N_23079,N_22676,N_22553);
xnor U23080 (N_23080,N_22717,N_22965);
xor U23081 (N_23081,N_22502,N_22805);
and U23082 (N_23082,N_22707,N_22955);
xor U23083 (N_23083,N_22902,N_22877);
xor U23084 (N_23084,N_22956,N_22538);
and U23085 (N_23085,N_22900,N_22640);
or U23086 (N_23086,N_22929,N_22564);
or U23087 (N_23087,N_22928,N_22835);
or U23088 (N_23088,N_22616,N_22672);
xnor U23089 (N_23089,N_22979,N_22596);
and U23090 (N_23090,N_22606,N_22620);
xor U23091 (N_23091,N_22715,N_22567);
nand U23092 (N_23092,N_22674,N_22774);
and U23093 (N_23093,N_22706,N_22711);
or U23094 (N_23094,N_22856,N_22974);
nand U23095 (N_23095,N_22659,N_22968);
xnor U23096 (N_23096,N_22994,N_22991);
or U23097 (N_23097,N_22587,N_22945);
nor U23098 (N_23098,N_22595,N_22628);
and U23099 (N_23099,N_22612,N_22765);
and U23100 (N_23100,N_22516,N_22817);
and U23101 (N_23101,N_22589,N_22556);
or U23102 (N_23102,N_22537,N_22657);
or U23103 (N_23103,N_22566,N_22635);
xnor U23104 (N_23104,N_22924,N_22947);
and U23105 (N_23105,N_22756,N_22798);
and U23106 (N_23106,N_22967,N_22971);
and U23107 (N_23107,N_22667,N_22931);
xor U23108 (N_23108,N_22920,N_22951);
xnor U23109 (N_23109,N_22675,N_22686);
nor U23110 (N_23110,N_22868,N_22938);
nand U23111 (N_23111,N_22872,N_22747);
nor U23112 (N_23112,N_22543,N_22544);
nand U23113 (N_23113,N_22944,N_22600);
xor U23114 (N_23114,N_22554,N_22699);
nand U23115 (N_23115,N_22895,N_22849);
nor U23116 (N_23116,N_22500,N_22752);
and U23117 (N_23117,N_22731,N_22861);
nand U23118 (N_23118,N_22901,N_22936);
and U23119 (N_23119,N_22598,N_22808);
or U23120 (N_23120,N_22812,N_22697);
and U23121 (N_23121,N_22823,N_22838);
nand U23122 (N_23122,N_22899,N_22599);
nor U23123 (N_23123,N_22722,N_22588);
nor U23124 (N_23124,N_22605,N_22757);
nand U23125 (N_23125,N_22896,N_22745);
nor U23126 (N_23126,N_22801,N_22555);
nor U23127 (N_23127,N_22885,N_22655);
nor U23128 (N_23128,N_22845,N_22561);
and U23129 (N_23129,N_22730,N_22664);
xor U23130 (N_23130,N_22682,N_22860);
or U23131 (N_23131,N_22736,N_22802);
xnor U23132 (N_23132,N_22704,N_22683);
or U23133 (N_23133,N_22993,N_22744);
nand U23134 (N_23134,N_22784,N_22572);
and U23135 (N_23135,N_22973,N_22910);
nor U23136 (N_23136,N_22703,N_22718);
or U23137 (N_23137,N_22696,N_22610);
nand U23138 (N_23138,N_22690,N_22954);
nor U23139 (N_23139,N_22727,N_22540);
xnor U23140 (N_23140,N_22597,N_22978);
and U23141 (N_23141,N_22942,N_22846);
and U23142 (N_23142,N_22775,N_22515);
xor U23143 (N_23143,N_22751,N_22905);
nor U23144 (N_23144,N_22783,N_22977);
or U23145 (N_23145,N_22761,N_22884);
and U23146 (N_23146,N_22526,N_22830);
and U23147 (N_23147,N_22915,N_22691);
and U23148 (N_23148,N_22759,N_22518);
or U23149 (N_23149,N_22809,N_22957);
or U23150 (N_23150,N_22788,N_22746);
xnor U23151 (N_23151,N_22665,N_22681);
nand U23152 (N_23152,N_22627,N_22811);
nor U23153 (N_23153,N_22800,N_22568);
nor U23154 (N_23154,N_22656,N_22853);
and U23155 (N_23155,N_22842,N_22529);
xor U23156 (N_23156,N_22558,N_22960);
and U23157 (N_23157,N_22988,N_22810);
xor U23158 (N_23158,N_22995,N_22630);
nand U23159 (N_23159,N_22658,N_22821);
nor U23160 (N_23160,N_22803,N_22848);
or U23161 (N_23161,N_22720,N_22590);
or U23162 (N_23162,N_22753,N_22559);
and U23163 (N_23163,N_22617,N_22585);
or U23164 (N_23164,N_22992,N_22943);
or U23165 (N_23165,N_22983,N_22565);
xor U23166 (N_23166,N_22714,N_22776);
xor U23167 (N_23167,N_22917,N_22807);
nor U23168 (N_23168,N_22542,N_22673);
or U23169 (N_23169,N_22854,N_22708);
nor U23170 (N_23170,N_22688,N_22694);
xor U23171 (N_23171,N_22591,N_22886);
xor U23172 (N_23172,N_22829,N_22767);
or U23173 (N_23173,N_22649,N_22547);
nand U23174 (N_23174,N_22958,N_22520);
nor U23175 (N_23175,N_22780,N_22634);
xnor U23176 (N_23176,N_22949,N_22844);
xor U23177 (N_23177,N_22530,N_22789);
nand U23178 (N_23178,N_22679,N_22608);
or U23179 (N_23179,N_22586,N_22999);
and U23180 (N_23180,N_22898,N_22824);
and U23181 (N_23181,N_22522,N_22662);
or U23182 (N_23182,N_22779,N_22661);
or U23183 (N_23183,N_22921,N_22990);
nand U23184 (N_23184,N_22952,N_22904);
or U23185 (N_23185,N_22646,N_22831);
xor U23186 (N_23186,N_22629,N_22618);
nor U23187 (N_23187,N_22881,N_22527);
xor U23188 (N_23188,N_22832,N_22532);
and U23189 (N_23189,N_22545,N_22733);
and U23190 (N_23190,N_22913,N_22563);
xor U23191 (N_23191,N_22782,N_22866);
nand U23192 (N_23192,N_22791,N_22787);
nor U23193 (N_23193,N_22950,N_22875);
xnor U23194 (N_23194,N_22948,N_22562);
nand U23195 (N_23195,N_22521,N_22914);
nor U23196 (N_23196,N_22976,N_22669);
xor U23197 (N_23197,N_22582,N_22581);
and U23198 (N_23198,N_22879,N_22878);
and U23199 (N_23199,N_22510,N_22523);
or U23200 (N_23200,N_22643,N_22893);
nand U23201 (N_23201,N_22889,N_22869);
and U23202 (N_23202,N_22833,N_22721);
nand U23203 (N_23203,N_22541,N_22710);
and U23204 (N_23204,N_22819,N_22797);
nor U23205 (N_23205,N_22863,N_22644);
xor U23206 (N_23206,N_22719,N_22638);
nor U23207 (N_23207,N_22578,N_22663);
nor U23208 (N_23208,N_22813,N_22728);
xnor U23209 (N_23209,N_22607,N_22903);
nand U23210 (N_23210,N_22763,N_22933);
nor U23211 (N_23211,N_22531,N_22998);
and U23212 (N_23212,N_22766,N_22941);
nor U23213 (N_23213,N_22723,N_22749);
xor U23214 (N_23214,N_22827,N_22716);
xnor U23215 (N_23215,N_22781,N_22726);
and U23216 (N_23216,N_22984,N_22639);
xnor U23217 (N_23217,N_22964,N_22799);
nand U23218 (N_23218,N_22891,N_22804);
nor U23219 (N_23219,N_22843,N_22918);
and U23220 (N_23220,N_22963,N_22836);
or U23221 (N_23221,N_22579,N_22865);
nor U23222 (N_23222,N_22946,N_22873);
nand U23223 (N_23223,N_22734,N_22580);
or U23224 (N_23224,N_22739,N_22650);
and U23225 (N_23225,N_22790,N_22623);
nor U23226 (N_23226,N_22997,N_22604);
or U23227 (N_23227,N_22922,N_22858);
nand U23228 (N_23228,N_22653,N_22754);
xnor U23229 (N_23229,N_22916,N_22847);
xor U23230 (N_23230,N_22795,N_22777);
and U23231 (N_23231,N_22855,N_22584);
or U23232 (N_23232,N_22923,N_22712);
nor U23233 (N_23233,N_22741,N_22574);
nor U23234 (N_23234,N_22709,N_22737);
xnor U23235 (N_23235,N_22509,N_22626);
xor U23236 (N_23236,N_22550,N_22975);
nand U23237 (N_23237,N_22740,N_22768);
and U23238 (N_23238,N_22613,N_22859);
nor U23239 (N_23239,N_22504,N_22987);
xor U23240 (N_23240,N_22645,N_22871);
nor U23241 (N_23241,N_22517,N_22934);
or U23242 (N_23242,N_22560,N_22622);
xnor U23243 (N_23243,N_22794,N_22882);
nor U23244 (N_23244,N_22982,N_22735);
nand U23245 (N_23245,N_22702,N_22985);
or U23246 (N_23246,N_22512,N_22953);
or U23247 (N_23247,N_22852,N_22549);
xor U23248 (N_23248,N_22758,N_22609);
and U23249 (N_23249,N_22624,N_22932);
nand U23250 (N_23250,N_22508,N_22842);
nor U23251 (N_23251,N_22779,N_22793);
and U23252 (N_23252,N_22994,N_22942);
and U23253 (N_23253,N_22788,N_22947);
xor U23254 (N_23254,N_22753,N_22645);
xor U23255 (N_23255,N_22584,N_22954);
nor U23256 (N_23256,N_22842,N_22832);
xor U23257 (N_23257,N_22916,N_22999);
nand U23258 (N_23258,N_22647,N_22829);
and U23259 (N_23259,N_22600,N_22647);
or U23260 (N_23260,N_22860,N_22681);
nor U23261 (N_23261,N_22507,N_22570);
or U23262 (N_23262,N_22716,N_22725);
and U23263 (N_23263,N_22707,N_22890);
nor U23264 (N_23264,N_22906,N_22892);
nand U23265 (N_23265,N_22612,N_22717);
xnor U23266 (N_23266,N_22850,N_22683);
xor U23267 (N_23267,N_22821,N_22766);
nand U23268 (N_23268,N_22602,N_22812);
and U23269 (N_23269,N_22791,N_22991);
nor U23270 (N_23270,N_22715,N_22699);
xnor U23271 (N_23271,N_22745,N_22709);
or U23272 (N_23272,N_22730,N_22649);
nand U23273 (N_23273,N_22765,N_22563);
nand U23274 (N_23274,N_22868,N_22535);
nor U23275 (N_23275,N_22742,N_22528);
or U23276 (N_23276,N_22540,N_22935);
xor U23277 (N_23277,N_22574,N_22935);
or U23278 (N_23278,N_22600,N_22932);
xnor U23279 (N_23279,N_22833,N_22940);
or U23280 (N_23280,N_22561,N_22638);
or U23281 (N_23281,N_22883,N_22529);
and U23282 (N_23282,N_22813,N_22756);
xnor U23283 (N_23283,N_22645,N_22849);
xor U23284 (N_23284,N_22661,N_22541);
nand U23285 (N_23285,N_22631,N_22682);
or U23286 (N_23286,N_22939,N_22759);
nor U23287 (N_23287,N_22550,N_22504);
and U23288 (N_23288,N_22821,N_22749);
nand U23289 (N_23289,N_22602,N_22902);
and U23290 (N_23290,N_22649,N_22703);
or U23291 (N_23291,N_22710,N_22772);
xnor U23292 (N_23292,N_22635,N_22616);
xor U23293 (N_23293,N_22893,N_22980);
nand U23294 (N_23294,N_22925,N_22649);
and U23295 (N_23295,N_22913,N_22981);
nand U23296 (N_23296,N_22714,N_22840);
nand U23297 (N_23297,N_22764,N_22532);
nand U23298 (N_23298,N_22880,N_22911);
and U23299 (N_23299,N_22533,N_22996);
xnor U23300 (N_23300,N_22974,N_22604);
xnor U23301 (N_23301,N_22537,N_22533);
and U23302 (N_23302,N_22809,N_22693);
xnor U23303 (N_23303,N_22970,N_22985);
nand U23304 (N_23304,N_22946,N_22823);
xor U23305 (N_23305,N_22703,N_22856);
xnor U23306 (N_23306,N_22837,N_22639);
nor U23307 (N_23307,N_22745,N_22506);
nor U23308 (N_23308,N_22825,N_22938);
or U23309 (N_23309,N_22970,N_22898);
nor U23310 (N_23310,N_22553,N_22763);
or U23311 (N_23311,N_22604,N_22947);
and U23312 (N_23312,N_22992,N_22839);
and U23313 (N_23313,N_22807,N_22677);
and U23314 (N_23314,N_22891,N_22794);
or U23315 (N_23315,N_22751,N_22862);
nand U23316 (N_23316,N_22775,N_22746);
nand U23317 (N_23317,N_22830,N_22528);
nand U23318 (N_23318,N_22558,N_22874);
xnor U23319 (N_23319,N_22775,N_22599);
nor U23320 (N_23320,N_22574,N_22846);
nor U23321 (N_23321,N_22954,N_22878);
nand U23322 (N_23322,N_22864,N_22531);
and U23323 (N_23323,N_22715,N_22538);
nor U23324 (N_23324,N_22528,N_22505);
or U23325 (N_23325,N_22829,N_22617);
or U23326 (N_23326,N_22665,N_22562);
and U23327 (N_23327,N_22544,N_22615);
and U23328 (N_23328,N_22987,N_22606);
or U23329 (N_23329,N_22677,N_22958);
nor U23330 (N_23330,N_22775,N_22633);
or U23331 (N_23331,N_22643,N_22738);
xor U23332 (N_23332,N_22841,N_22799);
nor U23333 (N_23333,N_22672,N_22759);
xnor U23334 (N_23334,N_22557,N_22822);
xor U23335 (N_23335,N_22514,N_22998);
and U23336 (N_23336,N_22753,N_22607);
and U23337 (N_23337,N_22549,N_22907);
and U23338 (N_23338,N_22653,N_22637);
or U23339 (N_23339,N_22584,N_22581);
nor U23340 (N_23340,N_22982,N_22952);
nor U23341 (N_23341,N_22687,N_22682);
nor U23342 (N_23342,N_22522,N_22527);
or U23343 (N_23343,N_22573,N_22882);
nor U23344 (N_23344,N_22843,N_22796);
and U23345 (N_23345,N_22778,N_22592);
nand U23346 (N_23346,N_22697,N_22507);
nor U23347 (N_23347,N_22541,N_22507);
nand U23348 (N_23348,N_22517,N_22947);
nor U23349 (N_23349,N_22868,N_22668);
xnor U23350 (N_23350,N_22735,N_22534);
xnor U23351 (N_23351,N_22874,N_22937);
nand U23352 (N_23352,N_22630,N_22726);
xnor U23353 (N_23353,N_22811,N_22654);
nand U23354 (N_23354,N_22865,N_22907);
and U23355 (N_23355,N_22781,N_22507);
and U23356 (N_23356,N_22837,N_22835);
nor U23357 (N_23357,N_22914,N_22768);
xor U23358 (N_23358,N_22903,N_22912);
and U23359 (N_23359,N_22934,N_22964);
nor U23360 (N_23360,N_22884,N_22860);
xor U23361 (N_23361,N_22515,N_22630);
and U23362 (N_23362,N_22644,N_22795);
nand U23363 (N_23363,N_22650,N_22838);
and U23364 (N_23364,N_22695,N_22504);
and U23365 (N_23365,N_22875,N_22621);
or U23366 (N_23366,N_22680,N_22644);
or U23367 (N_23367,N_22711,N_22502);
nor U23368 (N_23368,N_22800,N_22752);
nand U23369 (N_23369,N_22646,N_22611);
nand U23370 (N_23370,N_22525,N_22940);
xor U23371 (N_23371,N_22564,N_22578);
nor U23372 (N_23372,N_22829,N_22739);
or U23373 (N_23373,N_22946,N_22944);
or U23374 (N_23374,N_22655,N_22853);
nor U23375 (N_23375,N_22542,N_22718);
and U23376 (N_23376,N_22595,N_22670);
and U23377 (N_23377,N_22638,N_22627);
or U23378 (N_23378,N_22865,N_22531);
nand U23379 (N_23379,N_22992,N_22817);
nor U23380 (N_23380,N_22875,N_22519);
nor U23381 (N_23381,N_22680,N_22989);
nor U23382 (N_23382,N_22637,N_22506);
and U23383 (N_23383,N_22970,N_22745);
nor U23384 (N_23384,N_22822,N_22796);
nand U23385 (N_23385,N_22995,N_22594);
xor U23386 (N_23386,N_22750,N_22798);
or U23387 (N_23387,N_22667,N_22840);
xor U23388 (N_23388,N_22669,N_22981);
xor U23389 (N_23389,N_22788,N_22992);
and U23390 (N_23390,N_22819,N_22956);
nand U23391 (N_23391,N_22976,N_22787);
nand U23392 (N_23392,N_22866,N_22532);
nor U23393 (N_23393,N_22681,N_22515);
or U23394 (N_23394,N_22589,N_22705);
or U23395 (N_23395,N_22564,N_22840);
nor U23396 (N_23396,N_22535,N_22556);
nor U23397 (N_23397,N_22886,N_22645);
nand U23398 (N_23398,N_22990,N_22805);
and U23399 (N_23399,N_22643,N_22733);
and U23400 (N_23400,N_22921,N_22617);
xnor U23401 (N_23401,N_22850,N_22774);
nor U23402 (N_23402,N_22988,N_22545);
and U23403 (N_23403,N_22859,N_22807);
or U23404 (N_23404,N_22898,N_22799);
nor U23405 (N_23405,N_22593,N_22687);
or U23406 (N_23406,N_22636,N_22576);
nand U23407 (N_23407,N_22995,N_22745);
or U23408 (N_23408,N_22738,N_22656);
or U23409 (N_23409,N_22568,N_22934);
xnor U23410 (N_23410,N_22595,N_22744);
xor U23411 (N_23411,N_22652,N_22518);
or U23412 (N_23412,N_22664,N_22826);
or U23413 (N_23413,N_22541,N_22521);
nor U23414 (N_23414,N_22774,N_22769);
nand U23415 (N_23415,N_22910,N_22899);
xnor U23416 (N_23416,N_22636,N_22693);
nand U23417 (N_23417,N_22733,N_22793);
and U23418 (N_23418,N_22870,N_22587);
nand U23419 (N_23419,N_22516,N_22823);
or U23420 (N_23420,N_22593,N_22880);
nor U23421 (N_23421,N_22843,N_22888);
or U23422 (N_23422,N_22658,N_22720);
xnor U23423 (N_23423,N_22506,N_22726);
xnor U23424 (N_23424,N_22671,N_22926);
nor U23425 (N_23425,N_22610,N_22514);
and U23426 (N_23426,N_22830,N_22627);
xnor U23427 (N_23427,N_22795,N_22766);
nor U23428 (N_23428,N_22607,N_22749);
and U23429 (N_23429,N_22959,N_22903);
and U23430 (N_23430,N_22784,N_22756);
or U23431 (N_23431,N_22997,N_22758);
or U23432 (N_23432,N_22512,N_22517);
nor U23433 (N_23433,N_22980,N_22608);
and U23434 (N_23434,N_22878,N_22699);
or U23435 (N_23435,N_22931,N_22560);
or U23436 (N_23436,N_22742,N_22689);
nor U23437 (N_23437,N_22698,N_22802);
nor U23438 (N_23438,N_22886,N_22772);
and U23439 (N_23439,N_22664,N_22576);
or U23440 (N_23440,N_22854,N_22645);
and U23441 (N_23441,N_22599,N_22804);
nand U23442 (N_23442,N_22955,N_22935);
and U23443 (N_23443,N_22861,N_22612);
or U23444 (N_23444,N_22960,N_22778);
nand U23445 (N_23445,N_22558,N_22663);
or U23446 (N_23446,N_22532,N_22774);
xor U23447 (N_23447,N_22838,N_22821);
xor U23448 (N_23448,N_22828,N_22654);
or U23449 (N_23449,N_22642,N_22599);
and U23450 (N_23450,N_22994,N_22650);
xnor U23451 (N_23451,N_22772,N_22978);
or U23452 (N_23452,N_22857,N_22592);
nand U23453 (N_23453,N_22674,N_22783);
and U23454 (N_23454,N_22742,N_22666);
and U23455 (N_23455,N_22623,N_22714);
or U23456 (N_23456,N_22636,N_22981);
nand U23457 (N_23457,N_22841,N_22580);
nor U23458 (N_23458,N_22562,N_22551);
or U23459 (N_23459,N_22662,N_22750);
xnor U23460 (N_23460,N_22641,N_22663);
nand U23461 (N_23461,N_22501,N_22531);
or U23462 (N_23462,N_22956,N_22993);
xnor U23463 (N_23463,N_22671,N_22803);
xnor U23464 (N_23464,N_22670,N_22905);
or U23465 (N_23465,N_22574,N_22906);
xnor U23466 (N_23466,N_22936,N_22875);
or U23467 (N_23467,N_22759,N_22935);
nor U23468 (N_23468,N_22787,N_22576);
or U23469 (N_23469,N_22689,N_22637);
nor U23470 (N_23470,N_22806,N_22964);
xnor U23471 (N_23471,N_22553,N_22904);
and U23472 (N_23472,N_22907,N_22616);
and U23473 (N_23473,N_22881,N_22670);
nand U23474 (N_23474,N_22864,N_22956);
or U23475 (N_23475,N_22776,N_22566);
nand U23476 (N_23476,N_22506,N_22650);
nor U23477 (N_23477,N_22748,N_22828);
nor U23478 (N_23478,N_22940,N_22782);
and U23479 (N_23479,N_22706,N_22646);
or U23480 (N_23480,N_22544,N_22607);
nor U23481 (N_23481,N_22970,N_22742);
nor U23482 (N_23482,N_22937,N_22713);
nor U23483 (N_23483,N_22532,N_22743);
nand U23484 (N_23484,N_22635,N_22640);
or U23485 (N_23485,N_22588,N_22533);
and U23486 (N_23486,N_22759,N_22505);
nor U23487 (N_23487,N_22821,N_22514);
xnor U23488 (N_23488,N_22864,N_22827);
and U23489 (N_23489,N_22529,N_22766);
or U23490 (N_23490,N_22721,N_22530);
nor U23491 (N_23491,N_22827,N_22734);
xnor U23492 (N_23492,N_22637,N_22537);
or U23493 (N_23493,N_22595,N_22845);
or U23494 (N_23494,N_22563,N_22667);
nor U23495 (N_23495,N_22889,N_22531);
nor U23496 (N_23496,N_22974,N_22733);
and U23497 (N_23497,N_22862,N_22546);
xor U23498 (N_23498,N_22729,N_22683);
nand U23499 (N_23499,N_22710,N_22956);
nand U23500 (N_23500,N_23452,N_23049);
or U23501 (N_23501,N_23016,N_23065);
and U23502 (N_23502,N_23307,N_23328);
and U23503 (N_23503,N_23188,N_23163);
nor U23504 (N_23504,N_23475,N_23286);
nor U23505 (N_23505,N_23398,N_23006);
or U23506 (N_23506,N_23438,N_23312);
xor U23507 (N_23507,N_23074,N_23404);
nand U23508 (N_23508,N_23234,N_23171);
xnor U23509 (N_23509,N_23249,N_23124);
or U23510 (N_23510,N_23044,N_23193);
and U23511 (N_23511,N_23020,N_23268);
nand U23512 (N_23512,N_23185,N_23169);
xor U23513 (N_23513,N_23487,N_23258);
or U23514 (N_23514,N_23003,N_23410);
and U23515 (N_23515,N_23105,N_23356);
nand U23516 (N_23516,N_23116,N_23338);
nand U23517 (N_23517,N_23274,N_23181);
xor U23518 (N_23518,N_23494,N_23450);
nor U23519 (N_23519,N_23177,N_23341);
or U23520 (N_23520,N_23072,N_23265);
xor U23521 (N_23521,N_23127,N_23117);
nor U23522 (N_23522,N_23152,N_23413);
nor U23523 (N_23523,N_23189,N_23492);
or U23524 (N_23524,N_23148,N_23237);
and U23525 (N_23525,N_23203,N_23288);
xnor U23526 (N_23526,N_23036,N_23202);
nor U23527 (N_23527,N_23013,N_23473);
nand U23528 (N_23528,N_23362,N_23471);
nor U23529 (N_23529,N_23167,N_23285);
or U23530 (N_23530,N_23138,N_23088);
nor U23531 (N_23531,N_23057,N_23176);
and U23532 (N_23532,N_23370,N_23441);
xor U23533 (N_23533,N_23469,N_23140);
or U23534 (N_23534,N_23251,N_23290);
nand U23535 (N_23535,N_23392,N_23394);
nor U23536 (N_23536,N_23205,N_23159);
nand U23537 (N_23537,N_23108,N_23385);
nand U23538 (N_23538,N_23133,N_23296);
xor U23539 (N_23539,N_23309,N_23204);
or U23540 (N_23540,N_23486,N_23488);
or U23541 (N_23541,N_23464,N_23451);
and U23542 (N_23542,N_23200,N_23283);
nand U23543 (N_23543,N_23246,N_23001);
nor U23544 (N_23544,N_23078,N_23228);
xnor U23545 (N_23545,N_23231,N_23295);
or U23546 (N_23546,N_23449,N_23259);
and U23547 (N_23547,N_23018,N_23050);
or U23548 (N_23548,N_23344,N_23198);
nand U23549 (N_23549,N_23336,N_23238);
nor U23550 (N_23550,N_23150,N_23002);
and U23551 (N_23551,N_23028,N_23453);
and U23552 (N_23552,N_23120,N_23388);
or U23553 (N_23553,N_23374,N_23407);
xor U23554 (N_23554,N_23184,N_23484);
nor U23555 (N_23555,N_23023,N_23458);
and U23556 (N_23556,N_23099,N_23033);
or U23557 (N_23557,N_23254,N_23128);
or U23558 (N_23558,N_23168,N_23443);
xnor U23559 (N_23559,N_23287,N_23327);
xnor U23560 (N_23560,N_23009,N_23401);
xor U23561 (N_23561,N_23310,N_23419);
xor U23562 (N_23562,N_23257,N_23180);
xor U23563 (N_23563,N_23037,N_23495);
nand U23564 (N_23564,N_23276,N_23252);
nand U23565 (N_23565,N_23497,N_23080);
nor U23566 (N_23566,N_23051,N_23241);
or U23567 (N_23567,N_23250,N_23463);
or U23568 (N_23568,N_23048,N_23306);
and U23569 (N_23569,N_23101,N_23330);
nor U23570 (N_23570,N_23459,N_23104);
or U23571 (N_23571,N_23373,N_23420);
xnor U23572 (N_23572,N_23363,N_23481);
xor U23573 (N_23573,N_23038,N_23498);
nand U23574 (N_23574,N_23143,N_23224);
nand U23575 (N_23575,N_23151,N_23301);
nor U23576 (N_23576,N_23457,N_23027);
nand U23577 (N_23577,N_23197,N_23442);
nand U23578 (N_23578,N_23465,N_23432);
xnor U23579 (N_23579,N_23342,N_23405);
and U23580 (N_23580,N_23109,N_23055);
and U23581 (N_23581,N_23100,N_23434);
xnor U23582 (N_23582,N_23461,N_23244);
nor U23583 (N_23583,N_23262,N_23098);
nor U23584 (N_23584,N_23155,N_23218);
or U23585 (N_23585,N_23253,N_23381);
nand U23586 (N_23586,N_23162,N_23317);
and U23587 (N_23587,N_23289,N_23456);
nor U23588 (N_23588,N_23195,N_23358);
xnor U23589 (N_23589,N_23435,N_23447);
nand U23590 (N_23590,N_23364,N_23121);
nand U23591 (N_23591,N_23468,N_23216);
xor U23592 (N_23592,N_23350,N_23132);
xor U23593 (N_23593,N_23303,N_23066);
and U23594 (N_23594,N_23014,N_23446);
and U23595 (N_23595,N_23122,N_23482);
and U23596 (N_23596,N_23172,N_23382);
nand U23597 (N_23597,N_23149,N_23029);
xor U23598 (N_23598,N_23126,N_23349);
xnor U23599 (N_23599,N_23025,N_23085);
nand U23600 (N_23600,N_23247,N_23399);
xnor U23601 (N_23601,N_23470,N_23091);
or U23602 (N_23602,N_23112,N_23015);
and U23603 (N_23603,N_23368,N_23348);
or U23604 (N_23604,N_23073,N_23208);
or U23605 (N_23605,N_23190,N_23070);
and U23606 (N_23606,N_23275,N_23240);
nor U23607 (N_23607,N_23337,N_23480);
or U23608 (N_23608,N_23390,N_23056);
nor U23609 (N_23609,N_23455,N_23429);
nand U23610 (N_23610,N_23178,N_23115);
or U23611 (N_23611,N_23416,N_23479);
nor U23612 (N_23612,N_23311,N_23292);
nand U23613 (N_23613,N_23239,N_23436);
xor U23614 (N_23614,N_23041,N_23343);
nor U23615 (N_23615,N_23206,N_23192);
nor U23616 (N_23616,N_23280,N_23096);
nand U23617 (N_23617,N_23383,N_23084);
nor U23618 (N_23618,N_23145,N_23417);
or U23619 (N_23619,N_23272,N_23166);
xnor U23620 (N_23620,N_23040,N_23477);
or U23621 (N_23621,N_23094,N_23333);
xor U23622 (N_23622,N_23478,N_23110);
xor U23623 (N_23623,N_23142,N_23077);
and U23624 (N_23624,N_23427,N_23329);
xor U23625 (N_23625,N_23173,N_23229);
nand U23626 (N_23626,N_23406,N_23361);
or U23627 (N_23627,N_23075,N_23220);
nor U23628 (N_23628,N_23095,N_23485);
xnor U23629 (N_23629,N_23187,N_23087);
or U23630 (N_23630,N_23129,N_23000);
or U23631 (N_23631,N_23174,N_23313);
or U23632 (N_23632,N_23493,N_23157);
and U23633 (N_23633,N_23255,N_23294);
nand U23634 (N_23634,N_23182,N_23439);
nor U23635 (N_23635,N_23424,N_23213);
and U23636 (N_23636,N_23211,N_23011);
xor U23637 (N_23637,N_23396,N_23106);
nor U23638 (N_23638,N_23460,N_23352);
and U23639 (N_23639,N_23490,N_23378);
and U23640 (N_23640,N_23021,N_23302);
nor U23641 (N_23641,N_23466,N_23426);
or U23642 (N_23642,N_23332,N_23298);
nor U23643 (N_23643,N_23081,N_23359);
nor U23644 (N_23644,N_23153,N_23462);
nand U23645 (N_23645,N_23222,N_23403);
xnor U23646 (N_23646,N_23496,N_23499);
xor U23647 (N_23647,N_23232,N_23134);
nand U23648 (N_23648,N_23448,N_23165);
xor U23649 (N_23649,N_23347,N_23271);
xor U23650 (N_23650,N_23186,N_23007);
xnor U23651 (N_23651,N_23297,N_23273);
xnor U23652 (N_23652,N_23474,N_23137);
or U23653 (N_23653,N_23299,N_23183);
nor U23654 (N_23654,N_23305,N_23325);
and U23655 (N_23655,N_23346,N_23230);
or U23656 (N_23656,N_23141,N_23300);
and U23657 (N_23657,N_23428,N_23219);
nand U23658 (N_23658,N_23225,N_23114);
nor U23659 (N_23659,N_23256,N_23064);
or U23660 (N_23660,N_23017,N_23483);
nor U23661 (N_23661,N_23233,N_23422);
or U23662 (N_23662,N_23201,N_23054);
nor U23663 (N_23663,N_23035,N_23079);
nand U23664 (N_23664,N_23226,N_23371);
nor U23665 (N_23665,N_23334,N_23135);
or U23666 (N_23666,N_23393,N_23440);
nand U23667 (N_23667,N_23489,N_23323);
and U23668 (N_23668,N_23221,N_23067);
and U23669 (N_23669,N_23045,N_23111);
xnor U23670 (N_23670,N_23170,N_23062);
and U23671 (N_23671,N_23024,N_23278);
nand U23672 (N_23672,N_23082,N_23308);
nand U23673 (N_23673,N_23061,N_23414);
nand U23674 (N_23674,N_23318,N_23030);
and U23675 (N_23675,N_23154,N_23454);
nand U23676 (N_23676,N_23412,N_23365);
nand U23677 (N_23677,N_23353,N_23034);
xor U23678 (N_23678,N_23243,N_23076);
nand U23679 (N_23679,N_23217,N_23046);
and U23680 (N_23680,N_23042,N_23092);
and U23681 (N_23681,N_23068,N_23089);
xor U23682 (N_23682,N_23223,N_23476);
xor U23683 (N_23683,N_23131,N_23314);
nand U23684 (N_23684,N_23147,N_23093);
xnor U23685 (N_23685,N_23391,N_23158);
and U23686 (N_23686,N_23196,N_23322);
nor U23687 (N_23687,N_23026,N_23199);
or U23688 (N_23688,N_23380,N_23113);
nand U23689 (N_23689,N_23379,N_23209);
nor U23690 (N_23690,N_23063,N_23039);
nor U23691 (N_23691,N_23316,N_23384);
or U23692 (N_23692,N_23236,N_23433);
nand U23693 (N_23693,N_23005,N_23430);
or U23694 (N_23694,N_23279,N_23022);
nor U23695 (N_23695,N_23395,N_23086);
or U23696 (N_23696,N_23069,N_23212);
xor U23697 (N_23697,N_23103,N_23387);
or U23698 (N_23698,N_23340,N_23097);
or U23699 (N_23699,N_23156,N_23315);
nand U23700 (N_23700,N_23291,N_23210);
nand U23701 (N_23701,N_23418,N_23284);
xor U23702 (N_23702,N_23119,N_23397);
and U23703 (N_23703,N_23194,N_23047);
nand U23704 (N_23704,N_23031,N_23125);
xnor U23705 (N_23705,N_23375,N_23146);
or U23706 (N_23706,N_23179,N_23444);
nor U23707 (N_23707,N_23019,N_23402);
nor U23708 (N_23708,N_23389,N_23409);
nand U23709 (N_23709,N_23267,N_23372);
nand U23710 (N_23710,N_23425,N_23331);
and U23711 (N_23711,N_23052,N_23377);
nand U23712 (N_23712,N_23090,N_23386);
or U23713 (N_23713,N_23423,N_23264);
or U23714 (N_23714,N_23269,N_23281);
or U23715 (N_23715,N_23102,N_23248);
nor U23716 (N_23716,N_23277,N_23408);
xnor U23717 (N_23717,N_23130,N_23032);
or U23718 (N_23718,N_23139,N_23012);
nand U23719 (N_23719,N_23175,N_23261);
nor U23720 (N_23720,N_23369,N_23293);
nor U23721 (N_23721,N_23467,N_23367);
or U23722 (N_23722,N_23058,N_23335);
nor U23723 (N_23723,N_23160,N_23437);
or U23724 (N_23724,N_23431,N_23215);
and U23725 (N_23725,N_23136,N_23144);
nor U23726 (N_23726,N_23491,N_23242);
nor U23727 (N_23727,N_23366,N_23060);
nor U23728 (N_23728,N_23227,N_23360);
and U23729 (N_23729,N_23071,N_23083);
nand U23730 (N_23730,N_23059,N_23118);
and U23731 (N_23731,N_23266,N_23339);
and U23732 (N_23732,N_23004,N_23351);
nand U23733 (N_23733,N_23421,N_23107);
and U23734 (N_23734,N_23319,N_23376);
or U23735 (N_23735,N_23411,N_23355);
and U23736 (N_23736,N_23304,N_23164);
nor U23737 (N_23737,N_23010,N_23123);
or U23738 (N_23738,N_23400,N_23053);
and U23739 (N_23739,N_23214,N_23008);
nand U23740 (N_23740,N_23282,N_23321);
nor U23741 (N_23741,N_23263,N_23235);
or U23742 (N_23742,N_23320,N_23357);
or U23743 (N_23743,N_23270,N_23326);
and U23744 (N_23744,N_23161,N_23345);
xnor U23745 (N_23745,N_23260,N_23415);
and U23746 (N_23746,N_23207,N_23191);
or U23747 (N_23747,N_23445,N_23324);
nand U23748 (N_23748,N_23472,N_23245);
xor U23749 (N_23749,N_23043,N_23354);
xnor U23750 (N_23750,N_23468,N_23419);
nor U23751 (N_23751,N_23183,N_23212);
nand U23752 (N_23752,N_23423,N_23345);
nand U23753 (N_23753,N_23312,N_23222);
and U23754 (N_23754,N_23009,N_23253);
or U23755 (N_23755,N_23367,N_23164);
nor U23756 (N_23756,N_23420,N_23217);
nor U23757 (N_23757,N_23213,N_23281);
nand U23758 (N_23758,N_23010,N_23209);
nand U23759 (N_23759,N_23485,N_23278);
and U23760 (N_23760,N_23070,N_23069);
or U23761 (N_23761,N_23330,N_23437);
xor U23762 (N_23762,N_23008,N_23190);
nand U23763 (N_23763,N_23209,N_23140);
and U23764 (N_23764,N_23172,N_23252);
xnor U23765 (N_23765,N_23088,N_23238);
or U23766 (N_23766,N_23103,N_23129);
or U23767 (N_23767,N_23251,N_23127);
nand U23768 (N_23768,N_23446,N_23051);
xnor U23769 (N_23769,N_23049,N_23429);
or U23770 (N_23770,N_23428,N_23486);
nor U23771 (N_23771,N_23177,N_23036);
nand U23772 (N_23772,N_23449,N_23146);
and U23773 (N_23773,N_23229,N_23121);
or U23774 (N_23774,N_23327,N_23224);
nand U23775 (N_23775,N_23266,N_23239);
nand U23776 (N_23776,N_23363,N_23146);
nand U23777 (N_23777,N_23262,N_23254);
nand U23778 (N_23778,N_23067,N_23482);
or U23779 (N_23779,N_23246,N_23007);
or U23780 (N_23780,N_23030,N_23337);
xnor U23781 (N_23781,N_23355,N_23447);
or U23782 (N_23782,N_23306,N_23233);
or U23783 (N_23783,N_23457,N_23460);
and U23784 (N_23784,N_23430,N_23269);
nor U23785 (N_23785,N_23414,N_23261);
xor U23786 (N_23786,N_23098,N_23257);
xor U23787 (N_23787,N_23373,N_23022);
nor U23788 (N_23788,N_23070,N_23467);
nor U23789 (N_23789,N_23291,N_23049);
and U23790 (N_23790,N_23490,N_23000);
or U23791 (N_23791,N_23151,N_23194);
nand U23792 (N_23792,N_23263,N_23093);
nand U23793 (N_23793,N_23451,N_23373);
xor U23794 (N_23794,N_23064,N_23245);
nor U23795 (N_23795,N_23153,N_23468);
and U23796 (N_23796,N_23335,N_23411);
and U23797 (N_23797,N_23218,N_23357);
or U23798 (N_23798,N_23113,N_23131);
nor U23799 (N_23799,N_23035,N_23273);
or U23800 (N_23800,N_23083,N_23290);
xor U23801 (N_23801,N_23038,N_23306);
nor U23802 (N_23802,N_23065,N_23097);
xor U23803 (N_23803,N_23404,N_23331);
and U23804 (N_23804,N_23380,N_23066);
nor U23805 (N_23805,N_23069,N_23046);
and U23806 (N_23806,N_23346,N_23188);
xnor U23807 (N_23807,N_23166,N_23292);
and U23808 (N_23808,N_23320,N_23459);
and U23809 (N_23809,N_23047,N_23493);
and U23810 (N_23810,N_23362,N_23052);
and U23811 (N_23811,N_23369,N_23204);
nand U23812 (N_23812,N_23358,N_23204);
and U23813 (N_23813,N_23248,N_23405);
nand U23814 (N_23814,N_23034,N_23429);
nand U23815 (N_23815,N_23400,N_23390);
xnor U23816 (N_23816,N_23109,N_23053);
nand U23817 (N_23817,N_23347,N_23284);
or U23818 (N_23818,N_23283,N_23040);
nor U23819 (N_23819,N_23118,N_23375);
or U23820 (N_23820,N_23328,N_23277);
xnor U23821 (N_23821,N_23499,N_23010);
nor U23822 (N_23822,N_23333,N_23073);
nand U23823 (N_23823,N_23302,N_23441);
xnor U23824 (N_23824,N_23002,N_23256);
and U23825 (N_23825,N_23202,N_23006);
and U23826 (N_23826,N_23198,N_23029);
xnor U23827 (N_23827,N_23346,N_23450);
nand U23828 (N_23828,N_23279,N_23452);
nor U23829 (N_23829,N_23373,N_23342);
xnor U23830 (N_23830,N_23445,N_23286);
nand U23831 (N_23831,N_23240,N_23365);
or U23832 (N_23832,N_23245,N_23494);
nand U23833 (N_23833,N_23095,N_23362);
nand U23834 (N_23834,N_23348,N_23498);
and U23835 (N_23835,N_23392,N_23220);
xnor U23836 (N_23836,N_23261,N_23490);
nor U23837 (N_23837,N_23454,N_23110);
nor U23838 (N_23838,N_23332,N_23070);
and U23839 (N_23839,N_23264,N_23317);
nand U23840 (N_23840,N_23108,N_23133);
nand U23841 (N_23841,N_23031,N_23321);
nand U23842 (N_23842,N_23130,N_23492);
nor U23843 (N_23843,N_23082,N_23121);
nor U23844 (N_23844,N_23265,N_23195);
nand U23845 (N_23845,N_23059,N_23371);
nor U23846 (N_23846,N_23144,N_23484);
nand U23847 (N_23847,N_23124,N_23150);
nor U23848 (N_23848,N_23237,N_23046);
nand U23849 (N_23849,N_23115,N_23394);
xor U23850 (N_23850,N_23168,N_23208);
nor U23851 (N_23851,N_23131,N_23178);
nor U23852 (N_23852,N_23497,N_23294);
nor U23853 (N_23853,N_23327,N_23075);
or U23854 (N_23854,N_23081,N_23434);
or U23855 (N_23855,N_23157,N_23354);
nor U23856 (N_23856,N_23338,N_23402);
or U23857 (N_23857,N_23273,N_23106);
nand U23858 (N_23858,N_23046,N_23145);
xor U23859 (N_23859,N_23153,N_23002);
or U23860 (N_23860,N_23470,N_23311);
xor U23861 (N_23861,N_23068,N_23429);
nand U23862 (N_23862,N_23121,N_23477);
xor U23863 (N_23863,N_23227,N_23236);
nor U23864 (N_23864,N_23146,N_23031);
xnor U23865 (N_23865,N_23373,N_23066);
xnor U23866 (N_23866,N_23231,N_23205);
and U23867 (N_23867,N_23376,N_23344);
or U23868 (N_23868,N_23019,N_23213);
nand U23869 (N_23869,N_23261,N_23064);
and U23870 (N_23870,N_23091,N_23035);
nor U23871 (N_23871,N_23257,N_23115);
or U23872 (N_23872,N_23185,N_23040);
and U23873 (N_23873,N_23187,N_23339);
nand U23874 (N_23874,N_23119,N_23498);
xnor U23875 (N_23875,N_23375,N_23076);
nand U23876 (N_23876,N_23206,N_23412);
xnor U23877 (N_23877,N_23044,N_23228);
or U23878 (N_23878,N_23442,N_23396);
nor U23879 (N_23879,N_23438,N_23160);
or U23880 (N_23880,N_23307,N_23033);
nand U23881 (N_23881,N_23102,N_23134);
and U23882 (N_23882,N_23013,N_23486);
xor U23883 (N_23883,N_23235,N_23436);
and U23884 (N_23884,N_23454,N_23088);
and U23885 (N_23885,N_23053,N_23468);
xnor U23886 (N_23886,N_23272,N_23159);
or U23887 (N_23887,N_23488,N_23166);
or U23888 (N_23888,N_23452,N_23233);
and U23889 (N_23889,N_23264,N_23334);
xnor U23890 (N_23890,N_23218,N_23348);
nor U23891 (N_23891,N_23272,N_23210);
nor U23892 (N_23892,N_23220,N_23382);
nand U23893 (N_23893,N_23143,N_23155);
and U23894 (N_23894,N_23343,N_23380);
nor U23895 (N_23895,N_23155,N_23144);
xnor U23896 (N_23896,N_23474,N_23084);
or U23897 (N_23897,N_23384,N_23356);
nand U23898 (N_23898,N_23337,N_23262);
nand U23899 (N_23899,N_23462,N_23304);
and U23900 (N_23900,N_23469,N_23155);
and U23901 (N_23901,N_23224,N_23261);
nand U23902 (N_23902,N_23416,N_23124);
nand U23903 (N_23903,N_23191,N_23130);
or U23904 (N_23904,N_23276,N_23001);
nand U23905 (N_23905,N_23308,N_23479);
xor U23906 (N_23906,N_23471,N_23224);
nand U23907 (N_23907,N_23173,N_23338);
xor U23908 (N_23908,N_23493,N_23121);
xnor U23909 (N_23909,N_23264,N_23257);
xor U23910 (N_23910,N_23127,N_23133);
nor U23911 (N_23911,N_23244,N_23261);
nand U23912 (N_23912,N_23356,N_23144);
and U23913 (N_23913,N_23286,N_23245);
or U23914 (N_23914,N_23072,N_23338);
nor U23915 (N_23915,N_23360,N_23305);
nand U23916 (N_23916,N_23153,N_23114);
and U23917 (N_23917,N_23379,N_23251);
xor U23918 (N_23918,N_23366,N_23162);
nand U23919 (N_23919,N_23308,N_23102);
nand U23920 (N_23920,N_23286,N_23171);
xor U23921 (N_23921,N_23143,N_23341);
or U23922 (N_23922,N_23388,N_23178);
and U23923 (N_23923,N_23024,N_23169);
or U23924 (N_23924,N_23133,N_23124);
or U23925 (N_23925,N_23441,N_23348);
nand U23926 (N_23926,N_23012,N_23168);
and U23927 (N_23927,N_23483,N_23250);
or U23928 (N_23928,N_23448,N_23340);
xnor U23929 (N_23929,N_23479,N_23213);
nor U23930 (N_23930,N_23446,N_23483);
xnor U23931 (N_23931,N_23070,N_23090);
nand U23932 (N_23932,N_23072,N_23341);
nand U23933 (N_23933,N_23323,N_23189);
nand U23934 (N_23934,N_23457,N_23003);
nand U23935 (N_23935,N_23278,N_23384);
xor U23936 (N_23936,N_23455,N_23035);
and U23937 (N_23937,N_23447,N_23266);
nand U23938 (N_23938,N_23073,N_23316);
nand U23939 (N_23939,N_23496,N_23130);
nor U23940 (N_23940,N_23308,N_23087);
nand U23941 (N_23941,N_23168,N_23031);
xnor U23942 (N_23942,N_23189,N_23136);
xnor U23943 (N_23943,N_23096,N_23183);
and U23944 (N_23944,N_23409,N_23094);
nand U23945 (N_23945,N_23415,N_23249);
and U23946 (N_23946,N_23493,N_23411);
or U23947 (N_23947,N_23488,N_23230);
or U23948 (N_23948,N_23274,N_23273);
nand U23949 (N_23949,N_23378,N_23372);
xor U23950 (N_23950,N_23311,N_23293);
and U23951 (N_23951,N_23051,N_23400);
xnor U23952 (N_23952,N_23461,N_23115);
nor U23953 (N_23953,N_23167,N_23234);
nor U23954 (N_23954,N_23450,N_23047);
nand U23955 (N_23955,N_23224,N_23439);
and U23956 (N_23956,N_23139,N_23293);
and U23957 (N_23957,N_23485,N_23270);
xnor U23958 (N_23958,N_23261,N_23303);
nand U23959 (N_23959,N_23393,N_23465);
xor U23960 (N_23960,N_23237,N_23400);
xnor U23961 (N_23961,N_23202,N_23085);
nand U23962 (N_23962,N_23395,N_23417);
nor U23963 (N_23963,N_23185,N_23384);
and U23964 (N_23964,N_23288,N_23394);
nand U23965 (N_23965,N_23089,N_23177);
xnor U23966 (N_23966,N_23277,N_23478);
nor U23967 (N_23967,N_23205,N_23133);
or U23968 (N_23968,N_23138,N_23051);
nor U23969 (N_23969,N_23440,N_23442);
xor U23970 (N_23970,N_23382,N_23336);
nor U23971 (N_23971,N_23078,N_23245);
nor U23972 (N_23972,N_23469,N_23354);
or U23973 (N_23973,N_23413,N_23084);
nor U23974 (N_23974,N_23074,N_23267);
xnor U23975 (N_23975,N_23076,N_23227);
nor U23976 (N_23976,N_23324,N_23209);
and U23977 (N_23977,N_23426,N_23314);
xor U23978 (N_23978,N_23225,N_23049);
nor U23979 (N_23979,N_23432,N_23405);
nor U23980 (N_23980,N_23377,N_23261);
xor U23981 (N_23981,N_23445,N_23133);
and U23982 (N_23982,N_23158,N_23293);
nand U23983 (N_23983,N_23213,N_23499);
nand U23984 (N_23984,N_23363,N_23243);
xor U23985 (N_23985,N_23152,N_23170);
nand U23986 (N_23986,N_23202,N_23458);
and U23987 (N_23987,N_23180,N_23292);
xor U23988 (N_23988,N_23073,N_23464);
or U23989 (N_23989,N_23430,N_23290);
or U23990 (N_23990,N_23146,N_23252);
xor U23991 (N_23991,N_23069,N_23109);
nor U23992 (N_23992,N_23386,N_23240);
xnor U23993 (N_23993,N_23048,N_23185);
or U23994 (N_23994,N_23456,N_23422);
or U23995 (N_23995,N_23453,N_23244);
xor U23996 (N_23996,N_23139,N_23301);
xnor U23997 (N_23997,N_23304,N_23336);
xnor U23998 (N_23998,N_23338,N_23459);
xnor U23999 (N_23999,N_23447,N_23467);
nor U24000 (N_24000,N_23844,N_23511);
xor U24001 (N_24001,N_23822,N_23628);
or U24002 (N_24002,N_23620,N_23750);
nand U24003 (N_24003,N_23833,N_23643);
nand U24004 (N_24004,N_23885,N_23711);
or U24005 (N_24005,N_23622,N_23825);
nand U24006 (N_24006,N_23797,N_23631);
and U24007 (N_24007,N_23829,N_23910);
xor U24008 (N_24008,N_23670,N_23933);
nand U24009 (N_24009,N_23819,N_23773);
and U24010 (N_24010,N_23696,N_23506);
nor U24011 (N_24011,N_23577,N_23751);
xnor U24012 (N_24012,N_23816,N_23530);
and U24013 (N_24013,N_23972,N_23663);
or U24014 (N_24014,N_23541,N_23898);
nor U24015 (N_24015,N_23509,N_23518);
or U24016 (N_24016,N_23640,N_23945);
or U24017 (N_24017,N_23966,N_23921);
nand U24018 (N_24018,N_23948,N_23680);
nand U24019 (N_24019,N_23864,N_23882);
nand U24020 (N_24020,N_23874,N_23674);
nor U24021 (N_24021,N_23848,N_23734);
xnor U24022 (N_24022,N_23672,N_23560);
nor U24023 (N_24023,N_23960,N_23975);
nor U24024 (N_24024,N_23916,N_23986);
xor U24025 (N_24025,N_23889,N_23533);
or U24026 (N_24026,N_23562,N_23818);
xnor U24027 (N_24027,N_23770,N_23570);
nor U24028 (N_24028,N_23705,N_23956);
or U24029 (N_24029,N_23891,N_23869);
or U24030 (N_24030,N_23718,N_23744);
or U24031 (N_24031,N_23618,N_23721);
xnor U24032 (N_24032,N_23629,N_23988);
or U24033 (N_24033,N_23644,N_23505);
and U24034 (N_24034,N_23746,N_23926);
nor U24035 (N_24035,N_23676,N_23626);
or U24036 (N_24036,N_23740,N_23920);
and U24037 (N_24037,N_23504,N_23604);
nor U24038 (N_24038,N_23652,N_23636);
xnor U24039 (N_24039,N_23519,N_23995);
nand U24040 (N_24040,N_23714,N_23534);
and U24041 (N_24041,N_23856,N_23949);
nor U24042 (N_24042,N_23919,N_23908);
nand U24043 (N_24043,N_23915,N_23962);
xor U24044 (N_24044,N_23867,N_23946);
nor U24045 (N_24045,N_23897,N_23909);
xor U24046 (N_24046,N_23621,N_23662);
and U24047 (N_24047,N_23594,N_23990);
or U24048 (N_24048,N_23775,N_23608);
and U24049 (N_24049,N_23840,N_23573);
and U24050 (N_24050,N_23794,N_23880);
nor U24051 (N_24051,N_23658,N_23704);
nor U24052 (N_24052,N_23588,N_23901);
and U24053 (N_24053,N_23826,N_23851);
or U24054 (N_24054,N_23590,N_23974);
nand U24055 (N_24055,N_23963,N_23735);
and U24056 (N_24056,N_23563,N_23685);
nor U24057 (N_24057,N_23625,N_23692);
or U24058 (N_24058,N_23715,N_23655);
or U24059 (N_24059,N_23632,N_23795);
and U24060 (N_24060,N_23583,N_23970);
nor U24061 (N_24061,N_23996,N_23515);
or U24062 (N_24062,N_23838,N_23706);
and U24063 (N_24063,N_23890,N_23811);
or U24064 (N_24064,N_23717,N_23766);
nand U24065 (N_24065,N_23792,N_23599);
nand U24066 (N_24066,N_23539,N_23922);
nor U24067 (N_24067,N_23940,N_23809);
nor U24068 (N_24068,N_23774,N_23613);
nand U24069 (N_24069,N_23650,N_23913);
or U24070 (N_24070,N_23862,N_23866);
xnor U24071 (N_24071,N_23703,N_23906);
and U24072 (N_24072,N_23571,N_23860);
xor U24073 (N_24073,N_23859,N_23955);
or U24074 (N_24074,N_23536,N_23842);
nand U24075 (N_24075,N_23656,N_23884);
nand U24076 (N_24076,N_23796,N_23727);
or U24077 (N_24077,N_23540,N_23681);
and U24078 (N_24078,N_23665,N_23596);
xnor U24079 (N_24079,N_23895,N_23764);
xnor U24080 (N_24080,N_23875,N_23902);
or U24081 (N_24081,N_23538,N_23992);
and U24082 (N_24082,N_23589,N_23899);
or U24083 (N_24083,N_23623,N_23602);
or U24084 (N_24084,N_23684,N_23595);
and U24085 (N_24085,N_23660,N_23501);
and U24086 (N_24086,N_23572,N_23947);
and U24087 (N_24087,N_23785,N_23635);
nand U24088 (N_24088,N_23688,N_23689);
or U24089 (N_24089,N_23597,N_23691);
or U24090 (N_24090,N_23872,N_23549);
or U24091 (N_24091,N_23784,N_23732);
nor U24092 (N_24092,N_23847,N_23609);
or U24093 (N_24093,N_23939,N_23815);
or U24094 (N_24094,N_23837,N_23682);
xnor U24095 (N_24095,N_23556,N_23544);
nor U24096 (N_24096,N_23502,N_23935);
or U24097 (N_24097,N_23559,N_23664);
and U24098 (N_24098,N_23907,N_23925);
or U24099 (N_24099,N_23873,N_23606);
nand U24100 (N_24100,N_23722,N_23930);
or U24101 (N_24101,N_23981,N_23839);
nor U24102 (N_24102,N_23893,N_23759);
nand U24103 (N_24103,N_23987,N_23781);
or U24104 (N_24104,N_23500,N_23984);
nand U24105 (N_24105,N_23886,N_23546);
and U24106 (N_24106,N_23771,N_23836);
xnor U24107 (N_24107,N_23834,N_23931);
nor U24108 (N_24108,N_23817,N_23624);
or U24109 (N_24109,N_23950,N_23641);
and U24110 (N_24110,N_23508,N_23814);
or U24111 (N_24111,N_23593,N_23845);
xnor U24112 (N_24112,N_23651,N_23954);
xnor U24113 (N_24113,N_23580,N_23671);
nor U24114 (N_24114,N_23642,N_23661);
and U24115 (N_24115,N_23720,N_23699);
nor U24116 (N_24116,N_23953,N_23568);
or U24117 (N_24117,N_23853,N_23564);
xnor U24118 (N_24118,N_23576,N_23823);
or U24119 (N_24119,N_23638,N_23630);
and U24120 (N_24120,N_23603,N_23657);
or U24121 (N_24121,N_23969,N_23786);
nor U24122 (N_24122,N_23830,N_23605);
or U24123 (N_24123,N_23787,N_23979);
or U24124 (N_24124,N_23532,N_23654);
nor U24125 (N_24125,N_23782,N_23683);
xnor U24126 (N_24126,N_23645,N_23832);
xor U24127 (N_24127,N_23617,N_23522);
xor U24128 (N_24128,N_23978,N_23894);
or U24129 (N_24129,N_23754,N_23550);
nor U24130 (N_24130,N_23788,N_23510);
nor U24131 (N_24131,N_23776,N_23531);
or U24132 (N_24132,N_23600,N_23876);
nand U24133 (N_24133,N_23914,N_23964);
nand U24134 (N_24134,N_23611,N_23768);
or U24135 (N_24135,N_23799,N_23738);
nand U24136 (N_24136,N_23747,N_23687);
nor U24137 (N_24137,N_23578,N_23709);
nand U24138 (N_24138,N_23753,N_23615);
xnor U24139 (N_24139,N_23524,N_23765);
nand U24140 (N_24140,N_23521,N_23892);
nor U24141 (N_24141,N_23574,N_23918);
nand U24142 (N_24142,N_23726,N_23852);
and U24143 (N_24143,N_23999,N_23783);
nor U24144 (N_24144,N_23824,N_23957);
xnor U24145 (N_24145,N_23561,N_23827);
nand U24146 (N_24146,N_23835,N_23690);
nand U24147 (N_24147,N_23793,N_23639);
nand U24148 (N_24148,N_23828,N_23733);
nand U24149 (N_24149,N_23610,N_23810);
nand U24150 (N_24150,N_23723,N_23760);
nand U24151 (N_24151,N_23877,N_23742);
nand U24152 (N_24152,N_23888,N_23968);
xnor U24153 (N_24153,N_23967,N_23917);
nor U24154 (N_24154,N_23865,N_23971);
nand U24155 (N_24155,N_23512,N_23843);
nor U24156 (N_24156,N_23543,N_23545);
and U24157 (N_24157,N_23813,N_23535);
and U24158 (N_24158,N_23707,N_23737);
xor U24159 (N_24159,N_23646,N_23857);
nand U24160 (N_24160,N_23778,N_23555);
xor U24161 (N_24161,N_23552,N_23649);
and U24162 (N_24162,N_23973,N_23694);
or U24163 (N_24163,N_23517,N_23739);
or U24164 (N_24164,N_23584,N_23695);
or U24165 (N_24165,N_23542,N_23929);
and U24166 (N_24166,N_23748,N_23769);
xnor U24167 (N_24167,N_23700,N_23719);
nand U24168 (N_24168,N_23812,N_23537);
or U24169 (N_24169,N_23741,N_23686);
and U24170 (N_24170,N_23951,N_23944);
and U24171 (N_24171,N_23667,N_23807);
and U24172 (N_24172,N_23780,N_23598);
and U24173 (N_24173,N_23841,N_23881);
nor U24174 (N_24174,N_23725,N_23958);
or U24175 (N_24175,N_23959,N_23976);
nand U24176 (N_24176,N_23516,N_23547);
nor U24177 (N_24177,N_23557,N_23708);
and U24178 (N_24178,N_23757,N_23761);
and U24179 (N_24179,N_23904,N_23668);
nor U24180 (N_24180,N_23850,N_23805);
or U24181 (N_24181,N_23961,N_23566);
xnor U24182 (N_24182,N_23804,N_23755);
xor U24183 (N_24183,N_23763,N_23728);
xnor U24184 (N_24184,N_23777,N_23965);
or U24185 (N_24185,N_23591,N_23586);
nand U24186 (N_24186,N_23679,N_23697);
nand U24187 (N_24187,N_23879,N_23789);
xnor U24188 (N_24188,N_23565,N_23616);
or U24189 (N_24189,N_23942,N_23745);
nand U24190 (N_24190,N_23592,N_23503);
nand U24191 (N_24191,N_23941,N_23701);
nand U24192 (N_24192,N_23729,N_23983);
nand U24193 (N_24193,N_23912,N_23554);
xor U24194 (N_24194,N_23749,N_23994);
or U24195 (N_24195,N_23582,N_23802);
and U24196 (N_24196,N_23587,N_23526);
or U24197 (N_24197,N_23558,N_23911);
nor U24198 (N_24198,N_23575,N_23846);
nand U24199 (N_24199,N_23905,N_23779);
or U24200 (N_24200,N_23693,N_23993);
xnor U24201 (N_24201,N_23861,N_23936);
xnor U24202 (N_24202,N_23669,N_23863);
or U24203 (N_24203,N_23520,N_23619);
and U24204 (N_24204,N_23713,N_23937);
xnor U24205 (N_24205,N_23762,N_23712);
and U24206 (N_24206,N_23934,N_23938);
xor U24207 (N_24207,N_23896,N_23855);
xnor U24208 (N_24208,N_23868,N_23648);
nand U24209 (N_24209,N_23743,N_23581);
xor U24210 (N_24210,N_23831,N_23579);
xor U24211 (N_24211,N_23928,N_23614);
nand U24212 (N_24212,N_23952,N_23698);
or U24213 (N_24213,N_23527,N_23932);
nor U24214 (N_24214,N_23752,N_23806);
nor U24215 (N_24215,N_23637,N_23569);
or U24216 (N_24216,N_23924,N_23767);
and U24217 (N_24217,N_23900,N_23528);
xor U24218 (N_24218,N_23607,N_23525);
nor U24219 (N_24219,N_23982,N_23653);
or U24220 (N_24220,N_23870,N_23716);
nand U24221 (N_24221,N_23801,N_23927);
nor U24222 (N_24222,N_23977,N_23858);
nor U24223 (N_24223,N_23772,N_23883);
or U24224 (N_24224,N_23633,N_23985);
or U24225 (N_24225,N_23800,N_23514);
nor U24226 (N_24226,N_23998,N_23991);
xor U24227 (N_24227,N_23523,N_23820);
nand U24228 (N_24228,N_23627,N_23675);
xor U24229 (N_24229,N_23567,N_23710);
nand U24230 (N_24230,N_23903,N_23678);
nand U24231 (N_24231,N_23798,N_23702);
nor U24232 (N_24232,N_23758,N_23871);
or U24233 (N_24233,N_23731,N_23730);
or U24234 (N_24234,N_23553,N_23673);
xnor U24235 (N_24235,N_23980,N_23997);
and U24236 (N_24236,N_23601,N_23791);
nand U24237 (N_24237,N_23666,N_23551);
nor U24238 (N_24238,N_23634,N_23659);
or U24239 (N_24239,N_23756,N_23887);
nor U24240 (N_24240,N_23878,N_23989);
xor U24241 (N_24241,N_23736,N_23790);
nor U24242 (N_24242,N_23943,N_23647);
nor U24243 (N_24243,N_23808,N_23507);
nand U24244 (N_24244,N_23612,N_23821);
nor U24245 (N_24245,N_23849,N_23854);
nand U24246 (N_24246,N_23724,N_23529);
nand U24247 (N_24247,N_23803,N_23513);
or U24248 (N_24248,N_23548,N_23585);
xor U24249 (N_24249,N_23923,N_23677);
and U24250 (N_24250,N_23947,N_23511);
or U24251 (N_24251,N_23831,N_23824);
nand U24252 (N_24252,N_23767,N_23506);
xor U24253 (N_24253,N_23502,N_23872);
or U24254 (N_24254,N_23961,N_23875);
nand U24255 (N_24255,N_23513,N_23844);
xor U24256 (N_24256,N_23570,N_23982);
and U24257 (N_24257,N_23856,N_23848);
nand U24258 (N_24258,N_23725,N_23791);
xnor U24259 (N_24259,N_23721,N_23613);
and U24260 (N_24260,N_23937,N_23801);
and U24261 (N_24261,N_23810,N_23867);
or U24262 (N_24262,N_23667,N_23777);
or U24263 (N_24263,N_23622,N_23689);
or U24264 (N_24264,N_23676,N_23839);
xor U24265 (N_24265,N_23909,N_23523);
or U24266 (N_24266,N_23657,N_23984);
nand U24267 (N_24267,N_23669,N_23652);
nand U24268 (N_24268,N_23521,N_23869);
xnor U24269 (N_24269,N_23620,N_23622);
nor U24270 (N_24270,N_23845,N_23863);
or U24271 (N_24271,N_23901,N_23783);
nor U24272 (N_24272,N_23796,N_23753);
nand U24273 (N_24273,N_23598,N_23563);
and U24274 (N_24274,N_23964,N_23974);
nor U24275 (N_24275,N_23855,N_23959);
nor U24276 (N_24276,N_23690,N_23733);
and U24277 (N_24277,N_23770,N_23809);
or U24278 (N_24278,N_23600,N_23962);
nor U24279 (N_24279,N_23500,N_23989);
or U24280 (N_24280,N_23787,N_23653);
or U24281 (N_24281,N_23918,N_23604);
xnor U24282 (N_24282,N_23709,N_23871);
nand U24283 (N_24283,N_23580,N_23561);
xnor U24284 (N_24284,N_23819,N_23950);
nor U24285 (N_24285,N_23595,N_23782);
xor U24286 (N_24286,N_23916,N_23870);
and U24287 (N_24287,N_23551,N_23979);
xor U24288 (N_24288,N_23874,N_23776);
and U24289 (N_24289,N_23512,N_23784);
xor U24290 (N_24290,N_23958,N_23606);
xnor U24291 (N_24291,N_23991,N_23931);
xnor U24292 (N_24292,N_23892,N_23533);
nor U24293 (N_24293,N_23994,N_23697);
nand U24294 (N_24294,N_23960,N_23889);
xnor U24295 (N_24295,N_23982,N_23833);
or U24296 (N_24296,N_23566,N_23518);
nand U24297 (N_24297,N_23561,N_23529);
and U24298 (N_24298,N_23544,N_23586);
or U24299 (N_24299,N_23793,N_23635);
and U24300 (N_24300,N_23611,N_23810);
xor U24301 (N_24301,N_23820,N_23780);
or U24302 (N_24302,N_23559,N_23944);
or U24303 (N_24303,N_23675,N_23743);
nand U24304 (N_24304,N_23647,N_23546);
nand U24305 (N_24305,N_23521,N_23870);
and U24306 (N_24306,N_23643,N_23779);
or U24307 (N_24307,N_23996,N_23732);
nor U24308 (N_24308,N_23786,N_23747);
nor U24309 (N_24309,N_23894,N_23893);
xor U24310 (N_24310,N_23531,N_23522);
and U24311 (N_24311,N_23834,N_23958);
nand U24312 (N_24312,N_23923,N_23862);
xor U24313 (N_24313,N_23692,N_23513);
or U24314 (N_24314,N_23613,N_23667);
and U24315 (N_24315,N_23517,N_23744);
xor U24316 (N_24316,N_23603,N_23799);
xnor U24317 (N_24317,N_23537,N_23878);
xnor U24318 (N_24318,N_23522,N_23984);
nand U24319 (N_24319,N_23882,N_23672);
and U24320 (N_24320,N_23590,N_23799);
nor U24321 (N_24321,N_23967,N_23874);
xnor U24322 (N_24322,N_23914,N_23941);
nor U24323 (N_24323,N_23880,N_23939);
and U24324 (N_24324,N_23533,N_23847);
xnor U24325 (N_24325,N_23829,N_23721);
nor U24326 (N_24326,N_23675,N_23539);
nand U24327 (N_24327,N_23771,N_23934);
nor U24328 (N_24328,N_23671,N_23737);
xnor U24329 (N_24329,N_23858,N_23536);
nand U24330 (N_24330,N_23773,N_23521);
nor U24331 (N_24331,N_23560,N_23638);
or U24332 (N_24332,N_23598,N_23874);
or U24333 (N_24333,N_23522,N_23871);
and U24334 (N_24334,N_23794,N_23765);
nand U24335 (N_24335,N_23909,N_23815);
nand U24336 (N_24336,N_23977,N_23608);
xnor U24337 (N_24337,N_23880,N_23596);
and U24338 (N_24338,N_23587,N_23505);
nor U24339 (N_24339,N_23973,N_23756);
nor U24340 (N_24340,N_23949,N_23963);
xor U24341 (N_24341,N_23553,N_23905);
nor U24342 (N_24342,N_23734,N_23973);
and U24343 (N_24343,N_23588,N_23706);
nor U24344 (N_24344,N_23573,N_23728);
nor U24345 (N_24345,N_23546,N_23917);
xnor U24346 (N_24346,N_23735,N_23648);
nor U24347 (N_24347,N_23689,N_23839);
xnor U24348 (N_24348,N_23667,N_23730);
and U24349 (N_24349,N_23988,N_23574);
xnor U24350 (N_24350,N_23625,N_23884);
nand U24351 (N_24351,N_23798,N_23552);
and U24352 (N_24352,N_23674,N_23796);
xnor U24353 (N_24353,N_23584,N_23763);
and U24354 (N_24354,N_23578,N_23585);
or U24355 (N_24355,N_23684,N_23854);
xor U24356 (N_24356,N_23608,N_23622);
xnor U24357 (N_24357,N_23894,N_23699);
nand U24358 (N_24358,N_23828,N_23680);
or U24359 (N_24359,N_23953,N_23763);
nand U24360 (N_24360,N_23855,N_23837);
nand U24361 (N_24361,N_23796,N_23899);
nor U24362 (N_24362,N_23639,N_23570);
nor U24363 (N_24363,N_23615,N_23673);
xor U24364 (N_24364,N_23668,N_23623);
or U24365 (N_24365,N_23914,N_23540);
nor U24366 (N_24366,N_23782,N_23691);
or U24367 (N_24367,N_23831,N_23981);
xor U24368 (N_24368,N_23664,N_23581);
or U24369 (N_24369,N_23984,N_23653);
and U24370 (N_24370,N_23632,N_23912);
xor U24371 (N_24371,N_23570,N_23946);
and U24372 (N_24372,N_23601,N_23899);
nand U24373 (N_24373,N_23814,N_23569);
xor U24374 (N_24374,N_23662,N_23502);
nor U24375 (N_24375,N_23775,N_23721);
nor U24376 (N_24376,N_23634,N_23825);
nor U24377 (N_24377,N_23826,N_23571);
nor U24378 (N_24378,N_23984,N_23857);
or U24379 (N_24379,N_23849,N_23793);
or U24380 (N_24380,N_23596,N_23802);
and U24381 (N_24381,N_23522,N_23975);
nor U24382 (N_24382,N_23890,N_23711);
xor U24383 (N_24383,N_23665,N_23532);
and U24384 (N_24384,N_23918,N_23701);
xor U24385 (N_24385,N_23625,N_23839);
xnor U24386 (N_24386,N_23773,N_23794);
and U24387 (N_24387,N_23552,N_23642);
nor U24388 (N_24388,N_23601,N_23858);
nor U24389 (N_24389,N_23613,N_23675);
and U24390 (N_24390,N_23964,N_23862);
nor U24391 (N_24391,N_23888,N_23920);
and U24392 (N_24392,N_23586,N_23625);
nor U24393 (N_24393,N_23714,N_23708);
nor U24394 (N_24394,N_23798,N_23841);
or U24395 (N_24395,N_23800,N_23900);
or U24396 (N_24396,N_23697,N_23710);
and U24397 (N_24397,N_23593,N_23715);
nand U24398 (N_24398,N_23602,N_23857);
xor U24399 (N_24399,N_23593,N_23519);
or U24400 (N_24400,N_23669,N_23534);
nor U24401 (N_24401,N_23797,N_23648);
xor U24402 (N_24402,N_23654,N_23856);
nand U24403 (N_24403,N_23993,N_23671);
xnor U24404 (N_24404,N_23881,N_23983);
nand U24405 (N_24405,N_23680,N_23723);
or U24406 (N_24406,N_23907,N_23961);
nand U24407 (N_24407,N_23847,N_23984);
and U24408 (N_24408,N_23679,N_23837);
xor U24409 (N_24409,N_23726,N_23874);
xnor U24410 (N_24410,N_23524,N_23653);
or U24411 (N_24411,N_23609,N_23749);
nor U24412 (N_24412,N_23534,N_23615);
xnor U24413 (N_24413,N_23745,N_23954);
and U24414 (N_24414,N_23577,N_23570);
nand U24415 (N_24415,N_23527,N_23519);
nor U24416 (N_24416,N_23599,N_23793);
nand U24417 (N_24417,N_23895,N_23826);
nor U24418 (N_24418,N_23837,N_23728);
xnor U24419 (N_24419,N_23558,N_23991);
and U24420 (N_24420,N_23640,N_23755);
nor U24421 (N_24421,N_23994,N_23599);
and U24422 (N_24422,N_23514,N_23698);
nor U24423 (N_24423,N_23723,N_23977);
xor U24424 (N_24424,N_23659,N_23990);
xor U24425 (N_24425,N_23505,N_23695);
xnor U24426 (N_24426,N_23959,N_23653);
xnor U24427 (N_24427,N_23601,N_23605);
xor U24428 (N_24428,N_23834,N_23618);
and U24429 (N_24429,N_23659,N_23853);
nand U24430 (N_24430,N_23798,N_23531);
or U24431 (N_24431,N_23531,N_23851);
xor U24432 (N_24432,N_23541,N_23536);
or U24433 (N_24433,N_23748,N_23607);
or U24434 (N_24434,N_23751,N_23715);
or U24435 (N_24435,N_23850,N_23641);
xnor U24436 (N_24436,N_23557,N_23627);
or U24437 (N_24437,N_23526,N_23994);
nand U24438 (N_24438,N_23580,N_23931);
and U24439 (N_24439,N_23865,N_23599);
nor U24440 (N_24440,N_23529,N_23686);
nor U24441 (N_24441,N_23672,N_23913);
or U24442 (N_24442,N_23790,N_23596);
nor U24443 (N_24443,N_23853,N_23693);
xnor U24444 (N_24444,N_23916,N_23519);
xnor U24445 (N_24445,N_23881,N_23914);
nor U24446 (N_24446,N_23646,N_23574);
and U24447 (N_24447,N_23957,N_23908);
or U24448 (N_24448,N_23767,N_23818);
and U24449 (N_24449,N_23674,N_23857);
and U24450 (N_24450,N_23934,N_23552);
nand U24451 (N_24451,N_23528,N_23563);
xor U24452 (N_24452,N_23589,N_23708);
and U24453 (N_24453,N_23792,N_23702);
xnor U24454 (N_24454,N_23888,N_23862);
xor U24455 (N_24455,N_23739,N_23998);
and U24456 (N_24456,N_23844,N_23713);
or U24457 (N_24457,N_23558,N_23667);
and U24458 (N_24458,N_23962,N_23579);
nand U24459 (N_24459,N_23675,N_23651);
nand U24460 (N_24460,N_23942,N_23630);
nand U24461 (N_24461,N_23756,N_23656);
nand U24462 (N_24462,N_23544,N_23795);
xor U24463 (N_24463,N_23558,N_23959);
and U24464 (N_24464,N_23579,N_23725);
nor U24465 (N_24465,N_23692,N_23889);
nand U24466 (N_24466,N_23584,N_23598);
and U24467 (N_24467,N_23805,N_23877);
and U24468 (N_24468,N_23523,N_23898);
nand U24469 (N_24469,N_23727,N_23565);
nand U24470 (N_24470,N_23563,N_23866);
xor U24471 (N_24471,N_23510,N_23922);
nand U24472 (N_24472,N_23631,N_23551);
xnor U24473 (N_24473,N_23747,N_23586);
nand U24474 (N_24474,N_23518,N_23883);
and U24475 (N_24475,N_23553,N_23617);
nand U24476 (N_24476,N_23658,N_23919);
xnor U24477 (N_24477,N_23550,N_23518);
and U24478 (N_24478,N_23542,N_23889);
nor U24479 (N_24479,N_23935,N_23566);
or U24480 (N_24480,N_23885,N_23820);
and U24481 (N_24481,N_23756,N_23661);
or U24482 (N_24482,N_23557,N_23923);
and U24483 (N_24483,N_23540,N_23566);
and U24484 (N_24484,N_23635,N_23536);
or U24485 (N_24485,N_23947,N_23922);
and U24486 (N_24486,N_23966,N_23595);
or U24487 (N_24487,N_23823,N_23805);
and U24488 (N_24488,N_23598,N_23830);
and U24489 (N_24489,N_23591,N_23970);
or U24490 (N_24490,N_23975,N_23734);
xnor U24491 (N_24491,N_23785,N_23850);
nand U24492 (N_24492,N_23665,N_23662);
or U24493 (N_24493,N_23955,N_23775);
nand U24494 (N_24494,N_23648,N_23640);
nand U24495 (N_24495,N_23889,N_23955);
nor U24496 (N_24496,N_23865,N_23578);
nand U24497 (N_24497,N_23579,N_23699);
and U24498 (N_24498,N_23917,N_23598);
and U24499 (N_24499,N_23698,N_23671);
or U24500 (N_24500,N_24185,N_24480);
and U24501 (N_24501,N_24439,N_24253);
nor U24502 (N_24502,N_24161,N_24332);
xor U24503 (N_24503,N_24022,N_24145);
nor U24504 (N_24504,N_24306,N_24357);
nor U24505 (N_24505,N_24056,N_24125);
xnor U24506 (N_24506,N_24411,N_24017);
and U24507 (N_24507,N_24392,N_24244);
xnor U24508 (N_24508,N_24334,N_24173);
or U24509 (N_24509,N_24199,N_24212);
and U24510 (N_24510,N_24382,N_24008);
xor U24511 (N_24511,N_24363,N_24373);
nor U24512 (N_24512,N_24116,N_24147);
or U24513 (N_24513,N_24497,N_24104);
and U24514 (N_24514,N_24178,N_24101);
xnor U24515 (N_24515,N_24435,N_24027);
and U24516 (N_24516,N_24192,N_24490);
nand U24517 (N_24517,N_24406,N_24469);
and U24518 (N_24518,N_24206,N_24450);
or U24519 (N_24519,N_24217,N_24274);
or U24520 (N_24520,N_24191,N_24209);
and U24521 (N_24521,N_24169,N_24397);
xnor U24522 (N_24522,N_24075,N_24283);
and U24523 (N_24523,N_24277,N_24030);
xor U24524 (N_24524,N_24126,N_24196);
and U24525 (N_24525,N_24476,N_24092);
nand U24526 (N_24526,N_24325,N_24226);
nand U24527 (N_24527,N_24098,N_24471);
xor U24528 (N_24528,N_24082,N_24235);
nor U24529 (N_24529,N_24035,N_24317);
nand U24530 (N_24530,N_24163,N_24354);
and U24531 (N_24531,N_24390,N_24431);
xnor U24532 (N_24532,N_24204,N_24474);
and U24533 (N_24533,N_24138,N_24093);
nand U24534 (N_24534,N_24032,N_24285);
nor U24535 (N_24535,N_24364,N_24459);
and U24536 (N_24536,N_24000,N_24262);
nor U24537 (N_24537,N_24352,N_24097);
or U24538 (N_24538,N_24172,N_24110);
and U24539 (N_24539,N_24407,N_24318);
and U24540 (N_24540,N_24399,N_24242);
xnor U24541 (N_24541,N_24090,N_24333);
nand U24542 (N_24542,N_24440,N_24324);
nor U24543 (N_24543,N_24380,N_24207);
nand U24544 (N_24544,N_24310,N_24449);
nand U24545 (N_24545,N_24350,N_24498);
nand U24546 (N_24546,N_24282,N_24046);
or U24547 (N_24547,N_24443,N_24393);
or U24548 (N_24548,N_24360,N_24137);
or U24549 (N_24549,N_24456,N_24273);
nand U24550 (N_24550,N_24103,N_24409);
and U24551 (N_24551,N_24058,N_24180);
xor U24552 (N_24552,N_24111,N_24322);
nand U24553 (N_24553,N_24268,N_24297);
nor U24554 (N_24554,N_24213,N_24493);
nor U24555 (N_24555,N_24256,N_24228);
or U24556 (N_24556,N_24053,N_24372);
nand U24557 (N_24557,N_24057,N_24007);
or U24558 (N_24558,N_24410,N_24321);
or U24559 (N_24559,N_24043,N_24224);
and U24560 (N_24560,N_24341,N_24156);
nor U24561 (N_24561,N_24036,N_24420);
xnor U24562 (N_24562,N_24200,N_24488);
nor U24563 (N_24563,N_24470,N_24349);
xnor U24564 (N_24564,N_24462,N_24002);
xor U24565 (N_24565,N_24302,N_24254);
nand U24566 (N_24566,N_24233,N_24168);
nor U24567 (N_24567,N_24379,N_24401);
and U24568 (N_24568,N_24425,N_24246);
nand U24569 (N_24569,N_24141,N_24139);
and U24570 (N_24570,N_24073,N_24181);
nor U24571 (N_24571,N_24236,N_24303);
xnor U24572 (N_24572,N_24122,N_24417);
nor U24573 (N_24573,N_24491,N_24031);
and U24574 (N_24574,N_24299,N_24408);
xor U24575 (N_24575,N_24182,N_24049);
nand U24576 (N_24576,N_24121,N_24259);
and U24577 (N_24577,N_24154,N_24383);
or U24578 (N_24578,N_24086,N_24369);
nor U24579 (N_24579,N_24059,N_24143);
and U24580 (N_24580,N_24066,N_24494);
xnor U24581 (N_24581,N_24275,N_24144);
xnor U24582 (N_24582,N_24424,N_24377);
xor U24583 (N_24583,N_24359,N_24269);
nand U24584 (N_24584,N_24128,N_24020);
nor U24585 (N_24585,N_24396,N_24452);
and U24586 (N_24586,N_24064,N_24294);
or U24587 (N_24587,N_24499,N_24095);
or U24588 (N_24588,N_24475,N_24001);
nor U24589 (N_24589,N_24251,N_24131);
xnor U24590 (N_24590,N_24198,N_24429);
xnor U24591 (N_24591,N_24281,N_24258);
and U24592 (N_24592,N_24403,N_24158);
nor U24593 (N_24593,N_24433,N_24320);
nor U24594 (N_24594,N_24361,N_24211);
or U24595 (N_24595,N_24339,N_24448);
nand U24596 (N_24596,N_24089,N_24190);
nor U24597 (N_24597,N_24009,N_24427);
and U24598 (N_24598,N_24077,N_24220);
nor U24599 (N_24599,N_24065,N_24489);
or U24600 (N_24600,N_24405,N_24311);
xor U24601 (N_24601,N_24216,N_24289);
and U24602 (N_24602,N_24343,N_24391);
nor U24603 (N_24603,N_24315,N_24423);
nor U24604 (N_24604,N_24358,N_24323);
xnor U24605 (N_24605,N_24313,N_24487);
nor U24606 (N_24606,N_24400,N_24347);
nor U24607 (N_24607,N_24271,N_24042);
xor U24608 (N_24608,N_24286,N_24107);
xnor U24609 (N_24609,N_24366,N_24245);
nor U24610 (N_24610,N_24447,N_24214);
or U24611 (N_24611,N_24076,N_24413);
or U24612 (N_24612,N_24276,N_24062);
nand U24613 (N_24613,N_24378,N_24033);
nand U24614 (N_24614,N_24314,N_24016);
and U24615 (N_24615,N_24280,N_24109);
nor U24616 (N_24616,N_24164,N_24331);
nand U24617 (N_24617,N_24039,N_24142);
xor U24618 (N_24618,N_24422,N_24025);
xnor U24619 (N_24619,N_24133,N_24070);
and U24620 (N_24620,N_24255,N_24307);
nand U24621 (N_24621,N_24345,N_24451);
xnor U24622 (N_24622,N_24290,N_24485);
or U24623 (N_24623,N_24015,N_24445);
and U24624 (N_24624,N_24437,N_24461);
nand U24625 (N_24625,N_24149,N_24218);
and U24626 (N_24626,N_24084,N_24284);
nand U24627 (N_24627,N_24463,N_24301);
nor U24628 (N_24628,N_24127,N_24003);
nor U24629 (N_24629,N_24150,N_24112);
nand U24630 (N_24630,N_24052,N_24029);
nor U24631 (N_24631,N_24219,N_24458);
xor U24632 (N_24632,N_24428,N_24465);
xnor U24633 (N_24633,N_24241,N_24071);
and U24634 (N_24634,N_24415,N_24351);
nand U24635 (N_24635,N_24210,N_24266);
and U24636 (N_24636,N_24028,N_24329);
or U24637 (N_24637,N_24371,N_24130);
and U24638 (N_24638,N_24477,N_24048);
xor U24639 (N_24639,N_24041,N_24316);
nand U24640 (N_24640,N_24436,N_24419);
and U24641 (N_24641,N_24006,N_24205);
xnor U24642 (N_24642,N_24388,N_24367);
or U24643 (N_24643,N_24384,N_24478);
xor U24644 (N_24644,N_24272,N_24394);
nor U24645 (N_24645,N_24155,N_24455);
xnor U24646 (N_24646,N_24215,N_24426);
or U24647 (N_24647,N_24335,N_24287);
nor U24648 (N_24648,N_24087,N_24250);
nand U24649 (N_24649,N_24105,N_24327);
xnor U24650 (N_24650,N_24047,N_24004);
nand U24651 (N_24651,N_24136,N_24165);
nand U24652 (N_24652,N_24123,N_24454);
nand U24653 (N_24653,N_24229,N_24492);
and U24654 (N_24654,N_24100,N_24061);
nor U24655 (N_24655,N_24157,N_24102);
nand U24656 (N_24656,N_24416,N_24063);
xnor U24657 (N_24657,N_24441,N_24326);
xnor U24658 (N_24658,N_24069,N_24012);
and U24659 (N_24659,N_24026,N_24328);
xnor U24660 (N_24660,N_24362,N_24412);
nor U24661 (N_24661,N_24175,N_24124);
xor U24662 (N_24662,N_24078,N_24312);
and U24663 (N_24663,N_24252,N_24495);
nand U24664 (N_24664,N_24374,N_24291);
or U24665 (N_24665,N_24186,N_24208);
xnor U24666 (N_24666,N_24050,N_24395);
nor U24667 (N_24667,N_24202,N_24068);
and U24668 (N_24668,N_24091,N_24381);
nand U24669 (N_24669,N_24134,N_24247);
nand U24670 (N_24670,N_24464,N_24421);
xor U24671 (N_24671,N_24468,N_24278);
xor U24672 (N_24672,N_24221,N_24010);
and U24673 (N_24673,N_24188,N_24055);
or U24674 (N_24674,N_24201,N_24094);
nor U24675 (N_24675,N_24432,N_24365);
and U24676 (N_24676,N_24296,N_24227);
or U24677 (N_24677,N_24385,N_24106);
nand U24678 (N_24678,N_24166,N_24132);
xor U24679 (N_24679,N_24167,N_24486);
nor U24680 (N_24680,N_24153,N_24060);
and U24681 (N_24681,N_24442,N_24402);
nand U24682 (N_24682,N_24234,N_24170);
nor U24683 (N_24683,N_24389,N_24240);
nand U24684 (N_24684,N_24496,N_24338);
nand U24685 (N_24685,N_24453,N_24298);
nor U24686 (N_24686,N_24044,N_24305);
and U24687 (N_24687,N_24249,N_24484);
or U24688 (N_24688,N_24135,N_24187);
xnor U24689 (N_24689,N_24288,N_24483);
nor U24690 (N_24690,N_24232,N_24054);
nand U24691 (N_24691,N_24482,N_24114);
nand U24692 (N_24692,N_24120,N_24336);
nor U24693 (N_24693,N_24230,N_24353);
xnor U24694 (N_24694,N_24481,N_24151);
nor U24695 (N_24695,N_24261,N_24248);
or U24696 (N_24696,N_24300,N_24040);
xor U24697 (N_24697,N_24330,N_24080);
nand U24698 (N_24698,N_24176,N_24239);
nor U24699 (N_24699,N_24096,N_24264);
and U24700 (N_24700,N_24088,N_24013);
nor U24701 (N_24701,N_24340,N_24024);
nand U24702 (N_24702,N_24203,N_24021);
or U24703 (N_24703,N_24148,N_24238);
nand U24704 (N_24704,N_24083,N_24171);
nor U24705 (N_24705,N_24140,N_24193);
and U24706 (N_24706,N_24270,N_24348);
nor U24707 (N_24707,N_24446,N_24177);
or U24708 (N_24708,N_24376,N_24267);
or U24709 (N_24709,N_24319,N_24237);
nand U24710 (N_24710,N_24018,N_24386);
nand U24711 (N_24711,N_24146,N_24467);
or U24712 (N_24712,N_24479,N_24337);
and U24713 (N_24713,N_24257,N_24079);
nor U24714 (N_24714,N_24460,N_24197);
nor U24715 (N_24715,N_24067,N_24295);
and U24716 (N_24716,N_24344,N_24072);
and U24717 (N_24717,N_24430,N_24263);
and U24718 (N_24718,N_24243,N_24113);
xor U24719 (N_24719,N_24183,N_24260);
xnor U24720 (N_24720,N_24466,N_24045);
xnor U24721 (N_24721,N_24152,N_24184);
and U24722 (N_24722,N_24368,N_24174);
nor U24723 (N_24723,N_24037,N_24179);
nor U24724 (N_24724,N_24023,N_24005);
or U24725 (N_24725,N_24051,N_24129);
or U24726 (N_24726,N_24117,N_24279);
nor U24727 (N_24727,N_24194,N_24099);
and U24728 (N_24728,N_24355,N_24265);
xnor U24729 (N_24729,N_24444,N_24231);
and U24730 (N_24730,N_24309,N_24356);
nand U24731 (N_24731,N_24160,N_24162);
or U24732 (N_24732,N_24115,N_24085);
nor U24733 (N_24733,N_24342,N_24119);
xnor U24734 (N_24734,N_24019,N_24011);
xnor U24735 (N_24735,N_24081,N_24118);
xnor U24736 (N_24736,N_24346,N_24308);
or U24737 (N_24737,N_24472,N_24195);
nand U24738 (N_24738,N_24292,N_24473);
xor U24739 (N_24739,N_24375,N_24418);
nand U24740 (N_24740,N_24293,N_24159);
or U24741 (N_24741,N_24225,N_24304);
xor U24742 (N_24742,N_24074,N_24404);
nand U24743 (N_24743,N_24223,N_24414);
and U24744 (N_24744,N_24108,N_24222);
nand U24745 (N_24745,N_24457,N_24398);
nand U24746 (N_24746,N_24370,N_24434);
or U24747 (N_24747,N_24034,N_24038);
nor U24748 (N_24748,N_24014,N_24189);
and U24749 (N_24749,N_24438,N_24387);
nand U24750 (N_24750,N_24462,N_24283);
xnor U24751 (N_24751,N_24347,N_24174);
xnor U24752 (N_24752,N_24435,N_24105);
or U24753 (N_24753,N_24418,N_24364);
nand U24754 (N_24754,N_24209,N_24093);
nor U24755 (N_24755,N_24487,N_24004);
nor U24756 (N_24756,N_24106,N_24157);
nand U24757 (N_24757,N_24109,N_24379);
xor U24758 (N_24758,N_24403,N_24291);
nand U24759 (N_24759,N_24335,N_24364);
nor U24760 (N_24760,N_24140,N_24172);
nand U24761 (N_24761,N_24214,N_24361);
nand U24762 (N_24762,N_24059,N_24289);
nand U24763 (N_24763,N_24417,N_24392);
and U24764 (N_24764,N_24204,N_24438);
or U24765 (N_24765,N_24025,N_24319);
nand U24766 (N_24766,N_24382,N_24314);
and U24767 (N_24767,N_24273,N_24487);
and U24768 (N_24768,N_24270,N_24274);
or U24769 (N_24769,N_24385,N_24031);
and U24770 (N_24770,N_24463,N_24280);
nor U24771 (N_24771,N_24474,N_24391);
nand U24772 (N_24772,N_24374,N_24365);
xor U24773 (N_24773,N_24301,N_24289);
nand U24774 (N_24774,N_24456,N_24253);
nor U24775 (N_24775,N_24292,N_24495);
nand U24776 (N_24776,N_24163,N_24438);
nand U24777 (N_24777,N_24024,N_24420);
nand U24778 (N_24778,N_24225,N_24274);
or U24779 (N_24779,N_24237,N_24239);
or U24780 (N_24780,N_24262,N_24292);
and U24781 (N_24781,N_24158,N_24221);
nor U24782 (N_24782,N_24214,N_24245);
and U24783 (N_24783,N_24365,N_24018);
or U24784 (N_24784,N_24249,N_24100);
xor U24785 (N_24785,N_24186,N_24009);
and U24786 (N_24786,N_24137,N_24008);
or U24787 (N_24787,N_24115,N_24461);
and U24788 (N_24788,N_24463,N_24013);
nor U24789 (N_24789,N_24139,N_24176);
or U24790 (N_24790,N_24319,N_24478);
nor U24791 (N_24791,N_24108,N_24194);
or U24792 (N_24792,N_24077,N_24172);
xnor U24793 (N_24793,N_24421,N_24005);
xor U24794 (N_24794,N_24181,N_24479);
or U24795 (N_24795,N_24062,N_24407);
and U24796 (N_24796,N_24289,N_24120);
nor U24797 (N_24797,N_24386,N_24120);
nand U24798 (N_24798,N_24301,N_24344);
nand U24799 (N_24799,N_24011,N_24303);
nor U24800 (N_24800,N_24369,N_24071);
nor U24801 (N_24801,N_24185,N_24439);
xnor U24802 (N_24802,N_24030,N_24122);
and U24803 (N_24803,N_24000,N_24361);
nor U24804 (N_24804,N_24468,N_24445);
and U24805 (N_24805,N_24206,N_24408);
and U24806 (N_24806,N_24353,N_24102);
nand U24807 (N_24807,N_24407,N_24179);
nor U24808 (N_24808,N_24302,N_24015);
or U24809 (N_24809,N_24151,N_24015);
and U24810 (N_24810,N_24463,N_24089);
xor U24811 (N_24811,N_24464,N_24120);
or U24812 (N_24812,N_24427,N_24018);
or U24813 (N_24813,N_24344,N_24202);
and U24814 (N_24814,N_24384,N_24204);
or U24815 (N_24815,N_24040,N_24389);
nor U24816 (N_24816,N_24167,N_24387);
nand U24817 (N_24817,N_24344,N_24428);
xor U24818 (N_24818,N_24194,N_24246);
nor U24819 (N_24819,N_24411,N_24002);
and U24820 (N_24820,N_24137,N_24225);
and U24821 (N_24821,N_24456,N_24088);
or U24822 (N_24822,N_24202,N_24356);
xnor U24823 (N_24823,N_24430,N_24058);
and U24824 (N_24824,N_24019,N_24235);
and U24825 (N_24825,N_24017,N_24115);
or U24826 (N_24826,N_24295,N_24044);
xor U24827 (N_24827,N_24158,N_24494);
or U24828 (N_24828,N_24061,N_24488);
nor U24829 (N_24829,N_24343,N_24212);
nand U24830 (N_24830,N_24093,N_24265);
or U24831 (N_24831,N_24474,N_24161);
xor U24832 (N_24832,N_24144,N_24430);
and U24833 (N_24833,N_24333,N_24492);
or U24834 (N_24834,N_24292,N_24205);
xor U24835 (N_24835,N_24146,N_24124);
and U24836 (N_24836,N_24242,N_24184);
nor U24837 (N_24837,N_24181,N_24289);
or U24838 (N_24838,N_24169,N_24105);
xor U24839 (N_24839,N_24342,N_24192);
xor U24840 (N_24840,N_24143,N_24398);
or U24841 (N_24841,N_24443,N_24165);
nand U24842 (N_24842,N_24230,N_24389);
and U24843 (N_24843,N_24296,N_24211);
or U24844 (N_24844,N_24036,N_24287);
or U24845 (N_24845,N_24285,N_24328);
and U24846 (N_24846,N_24272,N_24156);
xor U24847 (N_24847,N_24320,N_24499);
nor U24848 (N_24848,N_24245,N_24422);
and U24849 (N_24849,N_24023,N_24447);
nand U24850 (N_24850,N_24355,N_24302);
nand U24851 (N_24851,N_24040,N_24497);
nor U24852 (N_24852,N_24018,N_24245);
nor U24853 (N_24853,N_24274,N_24243);
and U24854 (N_24854,N_24419,N_24076);
nor U24855 (N_24855,N_24405,N_24363);
nor U24856 (N_24856,N_24386,N_24141);
nor U24857 (N_24857,N_24137,N_24388);
or U24858 (N_24858,N_24029,N_24160);
or U24859 (N_24859,N_24077,N_24260);
xnor U24860 (N_24860,N_24361,N_24442);
nand U24861 (N_24861,N_24449,N_24472);
nand U24862 (N_24862,N_24196,N_24029);
nor U24863 (N_24863,N_24023,N_24025);
nand U24864 (N_24864,N_24487,N_24159);
xor U24865 (N_24865,N_24085,N_24260);
nand U24866 (N_24866,N_24254,N_24173);
xnor U24867 (N_24867,N_24412,N_24405);
xnor U24868 (N_24868,N_24368,N_24049);
and U24869 (N_24869,N_24428,N_24070);
and U24870 (N_24870,N_24101,N_24290);
or U24871 (N_24871,N_24164,N_24058);
or U24872 (N_24872,N_24015,N_24099);
xor U24873 (N_24873,N_24011,N_24430);
or U24874 (N_24874,N_24121,N_24207);
or U24875 (N_24875,N_24364,N_24149);
nor U24876 (N_24876,N_24315,N_24451);
nor U24877 (N_24877,N_24273,N_24283);
nor U24878 (N_24878,N_24402,N_24099);
or U24879 (N_24879,N_24307,N_24291);
or U24880 (N_24880,N_24254,N_24359);
xor U24881 (N_24881,N_24127,N_24485);
nor U24882 (N_24882,N_24280,N_24177);
nor U24883 (N_24883,N_24208,N_24282);
nor U24884 (N_24884,N_24116,N_24001);
xor U24885 (N_24885,N_24212,N_24094);
nand U24886 (N_24886,N_24472,N_24233);
xor U24887 (N_24887,N_24378,N_24111);
xnor U24888 (N_24888,N_24342,N_24489);
and U24889 (N_24889,N_24459,N_24238);
or U24890 (N_24890,N_24395,N_24169);
or U24891 (N_24891,N_24133,N_24054);
and U24892 (N_24892,N_24107,N_24089);
nand U24893 (N_24893,N_24355,N_24246);
nor U24894 (N_24894,N_24187,N_24431);
and U24895 (N_24895,N_24175,N_24352);
nand U24896 (N_24896,N_24240,N_24292);
nand U24897 (N_24897,N_24306,N_24056);
nor U24898 (N_24898,N_24141,N_24095);
and U24899 (N_24899,N_24323,N_24030);
and U24900 (N_24900,N_24444,N_24122);
and U24901 (N_24901,N_24155,N_24283);
nor U24902 (N_24902,N_24096,N_24494);
nand U24903 (N_24903,N_24016,N_24350);
or U24904 (N_24904,N_24165,N_24473);
and U24905 (N_24905,N_24279,N_24410);
and U24906 (N_24906,N_24224,N_24164);
xor U24907 (N_24907,N_24356,N_24038);
and U24908 (N_24908,N_24301,N_24240);
nand U24909 (N_24909,N_24001,N_24152);
nand U24910 (N_24910,N_24372,N_24333);
xor U24911 (N_24911,N_24294,N_24001);
nand U24912 (N_24912,N_24318,N_24471);
xor U24913 (N_24913,N_24061,N_24075);
nand U24914 (N_24914,N_24245,N_24216);
nand U24915 (N_24915,N_24211,N_24157);
xnor U24916 (N_24916,N_24148,N_24101);
nand U24917 (N_24917,N_24370,N_24357);
or U24918 (N_24918,N_24095,N_24130);
nor U24919 (N_24919,N_24340,N_24460);
xor U24920 (N_24920,N_24219,N_24377);
nor U24921 (N_24921,N_24042,N_24003);
and U24922 (N_24922,N_24003,N_24085);
and U24923 (N_24923,N_24153,N_24241);
nand U24924 (N_24924,N_24233,N_24350);
and U24925 (N_24925,N_24161,N_24431);
or U24926 (N_24926,N_24426,N_24285);
xnor U24927 (N_24927,N_24232,N_24435);
nor U24928 (N_24928,N_24370,N_24459);
xor U24929 (N_24929,N_24399,N_24313);
nand U24930 (N_24930,N_24456,N_24002);
xor U24931 (N_24931,N_24421,N_24497);
or U24932 (N_24932,N_24390,N_24159);
and U24933 (N_24933,N_24355,N_24028);
nand U24934 (N_24934,N_24337,N_24335);
and U24935 (N_24935,N_24328,N_24158);
or U24936 (N_24936,N_24343,N_24464);
nor U24937 (N_24937,N_24394,N_24326);
and U24938 (N_24938,N_24491,N_24140);
nand U24939 (N_24939,N_24028,N_24014);
xor U24940 (N_24940,N_24218,N_24403);
nor U24941 (N_24941,N_24465,N_24376);
nand U24942 (N_24942,N_24461,N_24442);
xor U24943 (N_24943,N_24270,N_24475);
xor U24944 (N_24944,N_24103,N_24470);
nor U24945 (N_24945,N_24191,N_24265);
and U24946 (N_24946,N_24383,N_24309);
or U24947 (N_24947,N_24403,N_24168);
nand U24948 (N_24948,N_24250,N_24200);
nor U24949 (N_24949,N_24461,N_24121);
nor U24950 (N_24950,N_24426,N_24216);
nor U24951 (N_24951,N_24479,N_24407);
nor U24952 (N_24952,N_24484,N_24372);
xor U24953 (N_24953,N_24225,N_24273);
and U24954 (N_24954,N_24491,N_24090);
nor U24955 (N_24955,N_24411,N_24145);
nand U24956 (N_24956,N_24445,N_24386);
and U24957 (N_24957,N_24085,N_24439);
nand U24958 (N_24958,N_24077,N_24390);
xnor U24959 (N_24959,N_24421,N_24040);
and U24960 (N_24960,N_24009,N_24287);
nor U24961 (N_24961,N_24101,N_24031);
nor U24962 (N_24962,N_24059,N_24176);
nor U24963 (N_24963,N_24350,N_24425);
xnor U24964 (N_24964,N_24147,N_24123);
xnor U24965 (N_24965,N_24364,N_24011);
or U24966 (N_24966,N_24385,N_24004);
xor U24967 (N_24967,N_24193,N_24445);
nor U24968 (N_24968,N_24377,N_24281);
nand U24969 (N_24969,N_24329,N_24347);
nor U24970 (N_24970,N_24381,N_24386);
nand U24971 (N_24971,N_24499,N_24094);
xnor U24972 (N_24972,N_24086,N_24472);
and U24973 (N_24973,N_24477,N_24045);
xnor U24974 (N_24974,N_24368,N_24208);
nand U24975 (N_24975,N_24085,N_24034);
nand U24976 (N_24976,N_24113,N_24293);
and U24977 (N_24977,N_24011,N_24122);
or U24978 (N_24978,N_24140,N_24199);
nand U24979 (N_24979,N_24043,N_24315);
nor U24980 (N_24980,N_24097,N_24116);
and U24981 (N_24981,N_24084,N_24417);
xnor U24982 (N_24982,N_24397,N_24392);
xor U24983 (N_24983,N_24229,N_24369);
nor U24984 (N_24984,N_24031,N_24237);
and U24985 (N_24985,N_24232,N_24188);
xor U24986 (N_24986,N_24326,N_24393);
nor U24987 (N_24987,N_24220,N_24049);
and U24988 (N_24988,N_24268,N_24464);
and U24989 (N_24989,N_24030,N_24358);
nor U24990 (N_24990,N_24274,N_24272);
xor U24991 (N_24991,N_24489,N_24005);
xnor U24992 (N_24992,N_24477,N_24276);
xor U24993 (N_24993,N_24319,N_24443);
nand U24994 (N_24994,N_24155,N_24221);
nand U24995 (N_24995,N_24445,N_24181);
or U24996 (N_24996,N_24434,N_24137);
nand U24997 (N_24997,N_24043,N_24275);
xnor U24998 (N_24998,N_24253,N_24432);
and U24999 (N_24999,N_24384,N_24356);
and U25000 (N_25000,N_24942,N_24936);
nor U25001 (N_25001,N_24678,N_24774);
xor U25002 (N_25002,N_24501,N_24656);
nand U25003 (N_25003,N_24930,N_24700);
and U25004 (N_25004,N_24816,N_24775);
nand U25005 (N_25005,N_24896,N_24741);
or U25006 (N_25006,N_24973,N_24957);
nor U25007 (N_25007,N_24803,N_24565);
or U25008 (N_25008,N_24600,N_24830);
nand U25009 (N_25009,N_24799,N_24869);
or U25010 (N_25010,N_24866,N_24745);
and U25011 (N_25011,N_24928,N_24572);
or U25012 (N_25012,N_24946,N_24829);
nor U25013 (N_25013,N_24996,N_24779);
nor U25014 (N_25014,N_24691,N_24509);
xnor U25015 (N_25015,N_24513,N_24833);
xnor U25016 (N_25016,N_24765,N_24670);
or U25017 (N_25017,N_24732,N_24521);
nand U25018 (N_25018,N_24808,N_24716);
and U25019 (N_25019,N_24648,N_24606);
nand U25020 (N_25020,N_24954,N_24603);
or U25021 (N_25021,N_24850,N_24629);
xor U25022 (N_25022,N_24882,N_24534);
and U25023 (N_25023,N_24988,N_24794);
nor U25024 (N_25024,N_24943,N_24529);
or U25025 (N_25025,N_24556,N_24544);
and U25026 (N_25026,N_24522,N_24505);
nand U25027 (N_25027,N_24562,N_24801);
or U25028 (N_25028,N_24619,N_24904);
xnor U25029 (N_25029,N_24987,N_24901);
nor U25030 (N_25030,N_24704,N_24965);
nor U25031 (N_25031,N_24555,N_24759);
and U25032 (N_25032,N_24539,N_24652);
nand U25033 (N_25033,N_24986,N_24875);
or U25034 (N_25034,N_24961,N_24587);
xnor U25035 (N_25035,N_24564,N_24827);
and U25036 (N_25036,N_24511,N_24638);
and U25037 (N_25037,N_24682,N_24674);
and U25038 (N_25038,N_24981,N_24714);
xnor U25039 (N_25039,N_24791,N_24650);
nor U25040 (N_25040,N_24624,N_24836);
xnor U25041 (N_25041,N_24586,N_24862);
and U25042 (N_25042,N_24881,N_24897);
nand U25043 (N_25043,N_24695,N_24898);
and U25044 (N_25044,N_24515,N_24694);
or U25045 (N_25045,N_24559,N_24546);
xnor U25046 (N_25046,N_24916,N_24596);
or U25047 (N_25047,N_24938,N_24860);
xnor U25048 (N_25048,N_24785,N_24669);
nor U25049 (N_25049,N_24710,N_24653);
or U25050 (N_25050,N_24931,N_24968);
nor U25051 (N_25051,N_24767,N_24811);
nand U25052 (N_25052,N_24845,N_24722);
xor U25053 (N_25053,N_24995,N_24769);
xor U25054 (N_25054,N_24991,N_24841);
and U25055 (N_25055,N_24789,N_24910);
or U25056 (N_25056,N_24729,N_24728);
xor U25057 (N_25057,N_24594,N_24771);
xnor U25058 (N_25058,N_24602,N_24639);
and U25059 (N_25059,N_24579,N_24720);
nor U25060 (N_25060,N_24786,N_24907);
or U25061 (N_25061,N_24703,N_24610);
xor U25062 (N_25062,N_24895,N_24818);
nor U25063 (N_25063,N_24846,N_24580);
nor U25064 (N_25064,N_24997,N_24667);
and U25065 (N_25065,N_24552,N_24542);
or U25066 (N_25066,N_24840,N_24683);
xor U25067 (N_25067,N_24848,N_24575);
and U25068 (N_25068,N_24698,N_24978);
nor U25069 (N_25069,N_24891,N_24854);
nor U25070 (N_25070,N_24908,N_24664);
xnor U25071 (N_25071,N_24514,N_24831);
nand U25072 (N_25072,N_24815,N_24658);
nand U25073 (N_25073,N_24813,N_24770);
nand U25074 (N_25074,N_24956,N_24566);
and U25075 (N_25075,N_24738,N_24660);
and U25076 (N_25076,N_24661,N_24758);
nor U25077 (N_25077,N_24681,N_24725);
nor U25078 (N_25078,N_24753,N_24616);
or U25079 (N_25079,N_24625,N_24984);
or U25080 (N_25080,N_24533,N_24666);
xor U25081 (N_25081,N_24512,N_24592);
nor U25082 (N_25082,N_24541,N_24859);
and U25083 (N_25083,N_24649,N_24709);
xor U25084 (N_25084,N_24689,N_24574);
and U25085 (N_25085,N_24526,N_24755);
xor U25086 (N_25086,N_24900,N_24595);
nor U25087 (N_25087,N_24510,N_24633);
nand U25088 (N_25088,N_24932,N_24518);
and U25089 (N_25089,N_24825,N_24976);
nand U25090 (N_25090,N_24640,N_24504);
and U25091 (N_25091,N_24750,N_24828);
or U25092 (N_25092,N_24591,N_24749);
and U25093 (N_25093,N_24576,N_24715);
nor U25094 (N_25094,N_24888,N_24886);
and U25095 (N_25095,N_24982,N_24913);
xor U25096 (N_25096,N_24843,N_24708);
and U25097 (N_25097,N_24821,N_24920);
nor U25098 (N_25098,N_24820,N_24571);
and U25099 (N_25099,N_24538,N_24730);
and U25100 (N_25100,N_24754,N_24819);
or U25101 (N_25101,N_24736,N_24917);
nor U25102 (N_25102,N_24560,N_24757);
nor U25103 (N_25103,N_24532,N_24974);
nor U25104 (N_25104,N_24673,N_24702);
and U25105 (N_25105,N_24746,N_24584);
nand U25106 (N_25106,N_24557,N_24773);
and U25107 (N_25107,N_24966,N_24508);
and U25108 (N_25108,N_24655,N_24525);
nor U25109 (N_25109,N_24858,N_24782);
or U25110 (N_25110,N_24783,N_24756);
nand U25111 (N_25111,N_24675,N_24537);
and U25112 (N_25112,N_24644,N_24998);
or U25113 (N_25113,N_24925,N_24953);
nand U25114 (N_25114,N_24739,N_24817);
nand U25115 (N_25115,N_24618,N_24622);
xnor U25116 (N_25116,N_24588,N_24990);
or U25117 (N_25117,N_24585,N_24797);
nand U25118 (N_25118,N_24949,N_24937);
nor U25119 (N_25119,N_24812,N_24832);
and U25120 (N_25120,N_24615,N_24583);
and U25121 (N_25121,N_24856,N_24519);
nand U25122 (N_25122,N_24731,N_24795);
nand U25123 (N_25123,N_24663,N_24964);
or U25124 (N_25124,N_24631,N_24554);
and U25125 (N_25125,N_24561,N_24582);
and U25126 (N_25126,N_24723,N_24752);
nand U25127 (N_25127,N_24989,N_24601);
xnor U25128 (N_25128,N_24573,N_24993);
and U25129 (N_25129,N_24543,N_24926);
and U25130 (N_25130,N_24923,N_24983);
and U25131 (N_25131,N_24684,N_24798);
and U25132 (N_25132,N_24810,N_24507);
or U25133 (N_25133,N_24780,N_24955);
or U25134 (N_25134,N_24550,N_24697);
nand U25135 (N_25135,N_24608,N_24726);
and U25136 (N_25136,N_24548,N_24788);
nor U25137 (N_25137,N_24871,N_24826);
xnor U25138 (N_25138,N_24878,N_24877);
and U25139 (N_25139,N_24915,N_24951);
or U25140 (N_25140,N_24911,N_24958);
nand U25141 (N_25141,N_24906,N_24711);
and U25142 (N_25142,N_24634,N_24994);
nor U25143 (N_25143,N_24659,N_24855);
nor U25144 (N_25144,N_24568,N_24924);
xor U25145 (N_25145,N_24593,N_24581);
or U25146 (N_25146,N_24849,N_24941);
and U25147 (N_25147,N_24558,N_24654);
or U25148 (N_25148,N_24887,N_24516);
nand U25149 (N_25149,N_24620,N_24646);
xor U25150 (N_25150,N_24947,N_24761);
xor U25151 (N_25151,N_24970,N_24837);
or U25152 (N_25152,N_24962,N_24824);
and U25153 (N_25153,N_24717,N_24867);
xnor U25154 (N_25154,N_24796,N_24657);
xnor U25155 (N_25155,N_24630,N_24766);
nand U25156 (N_25156,N_24642,N_24706);
or U25157 (N_25157,N_24969,N_24598);
xor U25158 (N_25158,N_24705,N_24743);
nor U25159 (N_25159,N_24677,N_24852);
and U25160 (N_25160,N_24524,N_24948);
nor U25161 (N_25161,N_24626,N_24802);
xnor U25162 (N_25162,N_24975,N_24506);
xor U25163 (N_25163,N_24612,N_24879);
or U25164 (N_25164,N_24933,N_24870);
or U25165 (N_25165,N_24536,N_24944);
and U25166 (N_25166,N_24718,N_24935);
xnor U25167 (N_25167,N_24641,N_24805);
xnor U25168 (N_25168,N_24617,N_24790);
nor U25169 (N_25169,N_24945,N_24967);
xnor U25170 (N_25170,N_24692,N_24977);
nor U25171 (N_25171,N_24742,N_24893);
or U25172 (N_25172,N_24549,N_24873);
or U25173 (N_25173,N_24523,N_24545);
nand U25174 (N_25174,N_24686,N_24971);
or U25175 (N_25175,N_24889,N_24884);
nor U25176 (N_25176,N_24853,N_24872);
or U25177 (N_25177,N_24980,N_24985);
nor U25178 (N_25178,N_24876,N_24637);
xor U25179 (N_25179,N_24747,N_24733);
nor U25180 (N_25180,N_24502,N_24777);
and U25181 (N_25181,N_24950,N_24680);
and U25182 (N_25182,N_24643,N_24822);
and U25183 (N_25183,N_24645,N_24835);
and U25184 (N_25184,N_24861,N_24927);
nand U25185 (N_25185,N_24762,N_24687);
and U25186 (N_25186,N_24918,N_24874);
nand U25187 (N_25187,N_24764,N_24563);
nor U25188 (N_25188,N_24597,N_24679);
nor U25189 (N_25189,N_24992,N_24793);
and U25190 (N_25190,N_24590,N_24701);
xor U25191 (N_25191,N_24599,N_24919);
nand U25192 (N_25192,N_24778,N_24614);
xnor U25193 (N_25193,N_24890,N_24894);
xnor U25194 (N_25194,N_24902,N_24734);
nor U25195 (N_25195,N_24809,N_24632);
xor U25196 (N_25196,N_24699,N_24912);
nand U25197 (N_25197,N_24503,N_24688);
or U25198 (N_25198,N_24922,N_24972);
nor U25199 (N_25199,N_24685,N_24690);
and U25200 (N_25200,N_24520,N_24892);
nor U25201 (N_25201,N_24740,N_24903);
and U25202 (N_25202,N_24693,N_24863);
nor U25203 (N_25203,N_24500,N_24885);
and U25204 (N_25204,N_24963,N_24999);
xor U25205 (N_25205,N_24865,N_24934);
and U25206 (N_25206,N_24929,N_24647);
nor U25207 (N_25207,N_24914,N_24607);
and U25208 (N_25208,N_24735,N_24721);
nor U25209 (N_25209,N_24959,N_24851);
nor U25210 (N_25210,N_24578,N_24589);
nor U25211 (N_25211,N_24844,N_24613);
or U25212 (N_25212,N_24567,N_24528);
xor U25213 (N_25213,N_24671,N_24621);
xor U25214 (N_25214,N_24806,N_24787);
nand U25215 (N_25215,N_24952,N_24712);
xor U25216 (N_25216,N_24713,N_24760);
and U25217 (N_25217,N_24517,N_24883);
and U25218 (N_25218,N_24662,N_24696);
nor U25219 (N_25219,N_24939,N_24531);
or U25220 (N_25220,N_24921,N_24635);
nand U25221 (N_25221,N_24569,N_24979);
nand U25222 (N_25222,N_24672,N_24744);
nor U25223 (N_25223,N_24605,N_24847);
nor U25224 (N_25224,N_24838,N_24547);
and U25225 (N_25225,N_24724,N_24604);
nand U25226 (N_25226,N_24807,N_24857);
nor U25227 (N_25227,N_24636,N_24781);
or U25228 (N_25228,N_24839,N_24792);
or U25229 (N_25229,N_24707,N_24530);
nor U25230 (N_25230,N_24627,N_24772);
or U25231 (N_25231,N_24628,N_24880);
and U25232 (N_25232,N_24623,N_24905);
xnor U25233 (N_25233,N_24540,N_24577);
xnor U25234 (N_25234,N_24960,N_24651);
and U25235 (N_25235,N_24553,N_24611);
nor U25236 (N_25236,N_24868,N_24842);
nor U25237 (N_25237,N_24751,N_24899);
xor U25238 (N_25238,N_24823,N_24940);
and U25239 (N_25239,N_24609,N_24776);
or U25240 (N_25240,N_24719,N_24748);
nor U25241 (N_25241,N_24784,N_24768);
or U25242 (N_25242,N_24527,N_24864);
xnor U25243 (N_25243,N_24551,N_24763);
or U25244 (N_25244,N_24570,N_24814);
nand U25245 (N_25245,N_24834,N_24909);
xor U25246 (N_25246,N_24800,N_24668);
or U25247 (N_25247,N_24804,N_24535);
nor U25248 (N_25248,N_24737,N_24665);
nand U25249 (N_25249,N_24676,N_24727);
and U25250 (N_25250,N_24806,N_24855);
or U25251 (N_25251,N_24676,N_24691);
and U25252 (N_25252,N_24832,N_24748);
nor U25253 (N_25253,N_24690,N_24747);
xor U25254 (N_25254,N_24683,N_24794);
and U25255 (N_25255,N_24711,N_24749);
xnor U25256 (N_25256,N_24627,N_24767);
nor U25257 (N_25257,N_24717,N_24805);
nand U25258 (N_25258,N_24590,N_24904);
or U25259 (N_25259,N_24625,N_24981);
and U25260 (N_25260,N_24634,N_24740);
nand U25261 (N_25261,N_24829,N_24727);
and U25262 (N_25262,N_24852,N_24721);
and U25263 (N_25263,N_24718,N_24970);
nor U25264 (N_25264,N_24706,N_24769);
nand U25265 (N_25265,N_24925,N_24558);
nand U25266 (N_25266,N_24976,N_24881);
xnor U25267 (N_25267,N_24530,N_24644);
nor U25268 (N_25268,N_24513,N_24776);
nand U25269 (N_25269,N_24788,N_24944);
xor U25270 (N_25270,N_24894,N_24942);
and U25271 (N_25271,N_24638,N_24987);
xor U25272 (N_25272,N_24941,N_24757);
xnor U25273 (N_25273,N_24883,N_24762);
xor U25274 (N_25274,N_24964,N_24896);
nor U25275 (N_25275,N_24727,N_24906);
or U25276 (N_25276,N_24959,N_24732);
nor U25277 (N_25277,N_24634,N_24852);
and U25278 (N_25278,N_24807,N_24620);
nor U25279 (N_25279,N_24665,N_24528);
xor U25280 (N_25280,N_24950,N_24785);
or U25281 (N_25281,N_24709,N_24510);
xnor U25282 (N_25282,N_24657,N_24505);
and U25283 (N_25283,N_24673,N_24781);
nand U25284 (N_25284,N_24987,N_24919);
or U25285 (N_25285,N_24875,N_24670);
nor U25286 (N_25286,N_24569,N_24631);
and U25287 (N_25287,N_24946,N_24866);
nand U25288 (N_25288,N_24932,N_24713);
or U25289 (N_25289,N_24967,N_24513);
nand U25290 (N_25290,N_24686,N_24650);
and U25291 (N_25291,N_24732,N_24957);
xor U25292 (N_25292,N_24651,N_24893);
or U25293 (N_25293,N_24802,N_24767);
nor U25294 (N_25294,N_24844,N_24955);
or U25295 (N_25295,N_24683,N_24992);
or U25296 (N_25296,N_24640,N_24867);
and U25297 (N_25297,N_24902,N_24617);
nor U25298 (N_25298,N_24653,N_24614);
and U25299 (N_25299,N_24847,N_24968);
and U25300 (N_25300,N_24904,N_24521);
nor U25301 (N_25301,N_24757,N_24974);
nor U25302 (N_25302,N_24997,N_24785);
nor U25303 (N_25303,N_24918,N_24706);
nand U25304 (N_25304,N_24987,N_24563);
or U25305 (N_25305,N_24954,N_24638);
or U25306 (N_25306,N_24950,N_24694);
nand U25307 (N_25307,N_24727,N_24995);
xor U25308 (N_25308,N_24799,N_24695);
nor U25309 (N_25309,N_24539,N_24605);
and U25310 (N_25310,N_24950,N_24554);
or U25311 (N_25311,N_24540,N_24735);
xor U25312 (N_25312,N_24500,N_24570);
nand U25313 (N_25313,N_24787,N_24924);
xnor U25314 (N_25314,N_24819,N_24632);
xor U25315 (N_25315,N_24966,N_24874);
nor U25316 (N_25316,N_24716,N_24721);
and U25317 (N_25317,N_24542,N_24794);
nand U25318 (N_25318,N_24715,N_24859);
and U25319 (N_25319,N_24636,N_24847);
xor U25320 (N_25320,N_24919,N_24895);
xor U25321 (N_25321,N_24737,N_24942);
nor U25322 (N_25322,N_24947,N_24677);
xnor U25323 (N_25323,N_24990,N_24915);
nand U25324 (N_25324,N_24791,N_24549);
nand U25325 (N_25325,N_24617,N_24917);
and U25326 (N_25326,N_24938,N_24934);
xnor U25327 (N_25327,N_24672,N_24979);
nor U25328 (N_25328,N_24917,N_24849);
nand U25329 (N_25329,N_24685,N_24945);
nor U25330 (N_25330,N_24834,N_24889);
nand U25331 (N_25331,N_24623,N_24987);
nand U25332 (N_25332,N_24502,N_24520);
nand U25333 (N_25333,N_24627,N_24619);
nand U25334 (N_25334,N_24859,N_24994);
nor U25335 (N_25335,N_24584,N_24745);
and U25336 (N_25336,N_24950,N_24543);
or U25337 (N_25337,N_24771,N_24899);
nand U25338 (N_25338,N_24659,N_24755);
nand U25339 (N_25339,N_24879,N_24581);
and U25340 (N_25340,N_24505,N_24979);
xnor U25341 (N_25341,N_24674,N_24921);
nand U25342 (N_25342,N_24926,N_24604);
nor U25343 (N_25343,N_24900,N_24600);
and U25344 (N_25344,N_24728,N_24786);
nor U25345 (N_25345,N_24962,N_24866);
nor U25346 (N_25346,N_24734,N_24823);
and U25347 (N_25347,N_24926,N_24762);
nand U25348 (N_25348,N_24563,N_24867);
nand U25349 (N_25349,N_24579,N_24661);
or U25350 (N_25350,N_24946,N_24789);
nand U25351 (N_25351,N_24740,N_24542);
and U25352 (N_25352,N_24570,N_24803);
and U25353 (N_25353,N_24718,N_24743);
xnor U25354 (N_25354,N_24514,N_24972);
nand U25355 (N_25355,N_24589,N_24531);
nand U25356 (N_25356,N_24569,N_24555);
and U25357 (N_25357,N_24761,N_24980);
xor U25358 (N_25358,N_24745,N_24570);
nor U25359 (N_25359,N_24696,N_24873);
nor U25360 (N_25360,N_24747,N_24705);
nand U25361 (N_25361,N_24591,N_24785);
nand U25362 (N_25362,N_24685,N_24939);
nor U25363 (N_25363,N_24535,N_24530);
nand U25364 (N_25364,N_24700,N_24622);
and U25365 (N_25365,N_24920,N_24828);
nor U25366 (N_25366,N_24697,N_24861);
and U25367 (N_25367,N_24949,N_24780);
nor U25368 (N_25368,N_24607,N_24912);
nand U25369 (N_25369,N_24601,N_24976);
xnor U25370 (N_25370,N_24791,N_24961);
nand U25371 (N_25371,N_24588,N_24572);
or U25372 (N_25372,N_24746,N_24619);
nand U25373 (N_25373,N_24876,N_24514);
or U25374 (N_25374,N_24910,N_24965);
xor U25375 (N_25375,N_24676,N_24577);
xnor U25376 (N_25376,N_24882,N_24613);
nor U25377 (N_25377,N_24739,N_24606);
nor U25378 (N_25378,N_24720,N_24643);
xor U25379 (N_25379,N_24657,N_24960);
nor U25380 (N_25380,N_24706,N_24514);
and U25381 (N_25381,N_24767,N_24852);
nor U25382 (N_25382,N_24781,N_24590);
nand U25383 (N_25383,N_24607,N_24984);
nand U25384 (N_25384,N_24935,N_24956);
nor U25385 (N_25385,N_24968,N_24699);
xnor U25386 (N_25386,N_24759,N_24676);
and U25387 (N_25387,N_24946,N_24797);
and U25388 (N_25388,N_24766,N_24675);
nand U25389 (N_25389,N_24611,N_24702);
xor U25390 (N_25390,N_24722,N_24589);
and U25391 (N_25391,N_24743,N_24906);
xor U25392 (N_25392,N_24709,N_24640);
nor U25393 (N_25393,N_24950,N_24559);
xnor U25394 (N_25394,N_24695,N_24835);
nand U25395 (N_25395,N_24502,N_24513);
or U25396 (N_25396,N_24990,N_24515);
nor U25397 (N_25397,N_24734,N_24969);
nor U25398 (N_25398,N_24917,N_24921);
nor U25399 (N_25399,N_24664,N_24766);
nor U25400 (N_25400,N_24687,N_24743);
and U25401 (N_25401,N_24953,N_24614);
or U25402 (N_25402,N_24746,N_24543);
and U25403 (N_25403,N_24874,N_24520);
nor U25404 (N_25404,N_24524,N_24870);
nand U25405 (N_25405,N_24971,N_24988);
nor U25406 (N_25406,N_24787,N_24900);
and U25407 (N_25407,N_24783,N_24837);
xnor U25408 (N_25408,N_24605,N_24650);
and U25409 (N_25409,N_24681,N_24951);
and U25410 (N_25410,N_24776,N_24957);
nor U25411 (N_25411,N_24975,N_24889);
nor U25412 (N_25412,N_24569,N_24873);
and U25413 (N_25413,N_24773,N_24869);
xor U25414 (N_25414,N_24630,N_24842);
nor U25415 (N_25415,N_24761,N_24584);
and U25416 (N_25416,N_24841,N_24811);
nor U25417 (N_25417,N_24761,N_24674);
nand U25418 (N_25418,N_24896,N_24919);
xnor U25419 (N_25419,N_24564,N_24577);
nor U25420 (N_25420,N_24526,N_24841);
nand U25421 (N_25421,N_24601,N_24944);
nand U25422 (N_25422,N_24663,N_24629);
nor U25423 (N_25423,N_24643,N_24982);
nor U25424 (N_25424,N_24797,N_24807);
xnor U25425 (N_25425,N_24911,N_24848);
nor U25426 (N_25426,N_24574,N_24643);
and U25427 (N_25427,N_24630,N_24566);
xnor U25428 (N_25428,N_24877,N_24602);
nand U25429 (N_25429,N_24836,N_24610);
nand U25430 (N_25430,N_24917,N_24685);
or U25431 (N_25431,N_24781,N_24552);
and U25432 (N_25432,N_24687,N_24766);
nor U25433 (N_25433,N_24900,N_24807);
xnor U25434 (N_25434,N_24551,N_24872);
and U25435 (N_25435,N_24844,N_24889);
or U25436 (N_25436,N_24998,N_24564);
xnor U25437 (N_25437,N_24978,N_24854);
nor U25438 (N_25438,N_24519,N_24887);
or U25439 (N_25439,N_24752,N_24685);
nand U25440 (N_25440,N_24738,N_24923);
xnor U25441 (N_25441,N_24897,N_24629);
xnor U25442 (N_25442,N_24685,N_24898);
and U25443 (N_25443,N_24898,N_24853);
or U25444 (N_25444,N_24714,N_24885);
nand U25445 (N_25445,N_24787,N_24705);
nor U25446 (N_25446,N_24543,N_24503);
or U25447 (N_25447,N_24655,N_24876);
or U25448 (N_25448,N_24652,N_24709);
or U25449 (N_25449,N_24534,N_24978);
nand U25450 (N_25450,N_24721,N_24674);
nand U25451 (N_25451,N_24528,N_24549);
or U25452 (N_25452,N_24700,N_24850);
nor U25453 (N_25453,N_24584,N_24901);
and U25454 (N_25454,N_24541,N_24801);
nand U25455 (N_25455,N_24795,N_24838);
nor U25456 (N_25456,N_24751,N_24605);
and U25457 (N_25457,N_24506,N_24661);
nand U25458 (N_25458,N_24809,N_24557);
or U25459 (N_25459,N_24915,N_24632);
xor U25460 (N_25460,N_24850,N_24659);
and U25461 (N_25461,N_24727,N_24795);
nor U25462 (N_25462,N_24800,N_24617);
nor U25463 (N_25463,N_24828,N_24911);
or U25464 (N_25464,N_24570,N_24738);
and U25465 (N_25465,N_24731,N_24602);
nor U25466 (N_25466,N_24537,N_24676);
nor U25467 (N_25467,N_24958,N_24569);
xor U25468 (N_25468,N_24841,N_24533);
nand U25469 (N_25469,N_24593,N_24827);
nand U25470 (N_25470,N_24636,N_24708);
nand U25471 (N_25471,N_24508,N_24978);
xor U25472 (N_25472,N_24670,N_24523);
nand U25473 (N_25473,N_24875,N_24921);
and U25474 (N_25474,N_24748,N_24747);
nor U25475 (N_25475,N_24771,N_24903);
xor U25476 (N_25476,N_24778,N_24747);
xnor U25477 (N_25477,N_24942,N_24574);
nand U25478 (N_25478,N_24742,N_24996);
nor U25479 (N_25479,N_24785,N_24793);
nor U25480 (N_25480,N_24711,N_24968);
or U25481 (N_25481,N_24983,N_24925);
nand U25482 (N_25482,N_24561,N_24904);
or U25483 (N_25483,N_24744,N_24843);
xnor U25484 (N_25484,N_24884,N_24689);
nor U25485 (N_25485,N_24999,N_24719);
and U25486 (N_25486,N_24850,N_24810);
and U25487 (N_25487,N_24646,N_24541);
or U25488 (N_25488,N_24848,N_24593);
xnor U25489 (N_25489,N_24890,N_24759);
nor U25490 (N_25490,N_24543,N_24937);
and U25491 (N_25491,N_24511,N_24875);
nor U25492 (N_25492,N_24633,N_24612);
and U25493 (N_25493,N_24573,N_24508);
nor U25494 (N_25494,N_24898,N_24766);
xnor U25495 (N_25495,N_24591,N_24520);
nor U25496 (N_25496,N_24544,N_24923);
nor U25497 (N_25497,N_24856,N_24729);
nand U25498 (N_25498,N_24905,N_24547);
nor U25499 (N_25499,N_24863,N_24853);
and U25500 (N_25500,N_25448,N_25061);
xnor U25501 (N_25501,N_25303,N_25484);
xor U25502 (N_25502,N_25251,N_25246);
and U25503 (N_25503,N_25310,N_25214);
nand U25504 (N_25504,N_25018,N_25488);
xnor U25505 (N_25505,N_25462,N_25150);
or U25506 (N_25506,N_25458,N_25117);
and U25507 (N_25507,N_25434,N_25299);
or U25508 (N_25508,N_25389,N_25247);
xnor U25509 (N_25509,N_25017,N_25363);
nor U25510 (N_25510,N_25210,N_25275);
or U25511 (N_25511,N_25089,N_25411);
and U25512 (N_25512,N_25444,N_25006);
and U25513 (N_25513,N_25332,N_25074);
xor U25514 (N_25514,N_25268,N_25080);
and U25515 (N_25515,N_25125,N_25273);
or U25516 (N_25516,N_25248,N_25428);
and U25517 (N_25517,N_25403,N_25239);
xor U25518 (N_25518,N_25130,N_25082);
xor U25519 (N_25519,N_25071,N_25477);
nor U25520 (N_25520,N_25054,N_25404);
xnor U25521 (N_25521,N_25168,N_25147);
nor U25522 (N_25522,N_25162,N_25029);
nor U25523 (N_25523,N_25254,N_25452);
xor U25524 (N_25524,N_25262,N_25414);
and U25525 (N_25525,N_25366,N_25371);
nand U25526 (N_25526,N_25126,N_25209);
or U25527 (N_25527,N_25266,N_25114);
and U25528 (N_25528,N_25208,N_25395);
xnor U25529 (N_25529,N_25339,N_25044);
xor U25530 (N_25530,N_25177,N_25342);
or U25531 (N_25531,N_25330,N_25486);
nor U25532 (N_25532,N_25170,N_25108);
nor U25533 (N_25533,N_25203,N_25379);
and U25534 (N_25534,N_25085,N_25010);
nand U25535 (N_25535,N_25056,N_25120);
xor U25536 (N_25536,N_25440,N_25314);
nand U25537 (N_25537,N_25109,N_25399);
nor U25538 (N_25538,N_25464,N_25043);
nand U25539 (N_25539,N_25463,N_25323);
or U25540 (N_25540,N_25350,N_25055);
xnor U25541 (N_25541,N_25346,N_25438);
nor U25542 (N_25542,N_25425,N_25137);
nor U25543 (N_25543,N_25265,N_25227);
nor U25544 (N_25544,N_25232,N_25042);
or U25545 (N_25545,N_25454,N_25338);
nand U25546 (N_25546,N_25327,N_25128);
or U25547 (N_25547,N_25317,N_25468);
or U25548 (N_25548,N_25374,N_25489);
nand U25549 (N_25549,N_25207,N_25073);
nand U25550 (N_25550,N_25381,N_25009);
xor U25551 (N_25551,N_25311,N_25383);
nor U25552 (N_25552,N_25372,N_25133);
xor U25553 (N_25553,N_25474,N_25138);
and U25554 (N_25554,N_25058,N_25026);
xnor U25555 (N_25555,N_25271,N_25118);
nor U25556 (N_25556,N_25027,N_25176);
nor U25557 (N_25557,N_25072,N_25129);
nand U25558 (N_25558,N_25278,N_25415);
nor U25559 (N_25559,N_25102,N_25478);
and U25560 (N_25560,N_25321,N_25420);
nand U25561 (N_25561,N_25124,N_25421);
nor U25562 (N_25562,N_25305,N_25164);
or U25563 (N_25563,N_25049,N_25357);
xnor U25564 (N_25564,N_25066,N_25306);
nand U25565 (N_25565,N_25450,N_25308);
or U25566 (N_25566,N_25131,N_25101);
nand U25567 (N_25567,N_25161,N_25252);
nand U25568 (N_25568,N_25361,N_25015);
nor U25569 (N_25569,N_25217,N_25030);
nor U25570 (N_25570,N_25094,N_25076);
nand U25571 (N_25571,N_25416,N_25493);
and U25572 (N_25572,N_25236,N_25112);
nand U25573 (N_25573,N_25469,N_25461);
nand U25574 (N_25574,N_25078,N_25096);
nand U25575 (N_25575,N_25188,N_25167);
nor U25576 (N_25576,N_25175,N_25183);
nand U25577 (N_25577,N_25364,N_25281);
nor U25578 (N_25578,N_25392,N_25107);
nor U25579 (N_25579,N_25304,N_25480);
or U25580 (N_25580,N_25471,N_25190);
nor U25581 (N_25581,N_25482,N_25057);
nand U25582 (N_25582,N_25380,N_25136);
nand U25583 (N_25583,N_25255,N_25077);
or U25584 (N_25584,N_25064,N_25004);
xor U25585 (N_25585,N_25436,N_25433);
nor U25586 (N_25586,N_25040,N_25290);
or U25587 (N_25587,N_25135,N_25022);
xnor U25588 (N_25588,N_25343,N_25143);
xnor U25589 (N_25589,N_25408,N_25487);
nand U25590 (N_25590,N_25050,N_25422);
nor U25591 (N_25591,N_25081,N_25391);
and U25592 (N_25592,N_25257,N_25097);
and U25593 (N_25593,N_25154,N_25231);
or U25594 (N_25594,N_25197,N_25204);
and U25595 (N_25595,N_25483,N_25142);
nand U25596 (N_25596,N_25155,N_25038);
nand U25597 (N_25597,N_25386,N_25123);
xor U25598 (N_25598,N_25238,N_25084);
xnor U25599 (N_25599,N_25243,N_25276);
xor U25600 (N_25600,N_25402,N_25002);
nand U25601 (N_25601,N_25407,N_25166);
nor U25602 (N_25602,N_25198,N_25370);
and U25603 (N_25603,N_25329,N_25473);
or U25604 (N_25604,N_25424,N_25041);
nor U25605 (N_25605,N_25351,N_25272);
nand U25606 (N_25606,N_25356,N_25410);
nor U25607 (N_25607,N_25344,N_25492);
nand U25608 (N_25608,N_25220,N_25439);
xor U25609 (N_25609,N_25035,N_25358);
nor U25610 (N_25610,N_25105,N_25348);
and U25611 (N_25611,N_25485,N_25007);
xor U25612 (N_25612,N_25079,N_25086);
or U25613 (N_25613,N_25098,N_25312);
nand U25614 (N_25614,N_25033,N_25083);
and U25615 (N_25615,N_25088,N_25229);
xnor U25616 (N_25616,N_25368,N_25333);
xor U25617 (N_25617,N_25460,N_25192);
nor U25618 (N_25618,N_25315,N_25233);
and U25619 (N_25619,N_25360,N_25387);
nor U25620 (N_25620,N_25242,N_25467);
or U25621 (N_25621,N_25378,N_25146);
or U25622 (N_25622,N_25497,N_25223);
or U25623 (N_25623,N_25261,N_25263);
and U25624 (N_25624,N_25345,N_25157);
and U25625 (N_25625,N_25226,N_25417);
and U25626 (N_25626,N_25385,N_25291);
nor U25627 (N_25627,N_25359,N_25053);
nor U25628 (N_25628,N_25185,N_25400);
nand U25629 (N_25629,N_25000,N_25277);
xor U25630 (N_25630,N_25465,N_25316);
xor U25631 (N_25631,N_25435,N_25213);
or U25632 (N_25632,N_25068,N_25234);
nor U25633 (N_25633,N_25432,N_25228);
or U25634 (N_25634,N_25090,N_25326);
nand U25635 (N_25635,N_25221,N_25062);
or U25636 (N_25636,N_25014,N_25091);
and U25637 (N_25637,N_25301,N_25498);
or U25638 (N_25638,N_25455,N_25075);
or U25639 (N_25639,N_25060,N_25196);
or U25640 (N_25640,N_25369,N_25413);
or U25641 (N_25641,N_25111,N_25219);
nor U25642 (N_25642,N_25016,N_25365);
or U25643 (N_25643,N_25087,N_25152);
xnor U25644 (N_25644,N_25110,N_25423);
nand U25645 (N_25645,N_25297,N_25045);
nor U25646 (N_25646,N_25211,N_25446);
or U25647 (N_25647,N_25051,N_25367);
nor U25648 (N_25648,N_25264,N_25334);
and U25649 (N_25649,N_25116,N_25394);
nand U25650 (N_25650,N_25382,N_25104);
and U25651 (N_25651,N_25279,N_25300);
or U25652 (N_25652,N_25249,N_25193);
and U25653 (N_25653,N_25396,N_25437);
or U25654 (N_25654,N_25459,N_25285);
nor U25655 (N_25655,N_25470,N_25354);
nor U25656 (N_25656,N_25453,N_25447);
and U25657 (N_25657,N_25148,N_25490);
xor U25658 (N_25658,N_25184,N_25186);
nor U25659 (N_25659,N_25494,N_25199);
and U25660 (N_25660,N_25335,N_25302);
and U25661 (N_25661,N_25200,N_25443);
xnor U25662 (N_25662,N_25289,N_25496);
nor U25663 (N_25663,N_25144,N_25047);
or U25664 (N_25664,N_25409,N_25241);
and U25665 (N_25665,N_25325,N_25331);
and U25666 (N_25666,N_25298,N_25194);
nand U25667 (N_25667,N_25445,N_25426);
or U25668 (N_25668,N_25294,N_25293);
or U25669 (N_25669,N_25224,N_25202);
or U25670 (N_25670,N_25495,N_25309);
or U25671 (N_25671,N_25151,N_25012);
and U25672 (N_25672,N_25284,N_25205);
xnor U25673 (N_25673,N_25149,N_25259);
xnor U25674 (N_25674,N_25412,N_25256);
nand U25675 (N_25675,N_25375,N_25222);
nand U25676 (N_25676,N_25352,N_25491);
xnor U25677 (N_25677,N_25419,N_25067);
and U25678 (N_25678,N_25373,N_25225);
xor U25679 (N_25679,N_25179,N_25398);
xor U25680 (N_25680,N_25245,N_25260);
nor U25681 (N_25681,N_25376,N_25013);
nor U25682 (N_25682,N_25286,N_25020);
nor U25683 (N_25683,N_25139,N_25165);
nor U25684 (N_25684,N_25337,N_25025);
xnor U25685 (N_25685,N_25180,N_25244);
nand U25686 (N_25686,N_25270,N_25048);
nor U25687 (N_25687,N_25274,N_25159);
and U25688 (N_25688,N_25173,N_25212);
or U25689 (N_25689,N_25295,N_25099);
and U25690 (N_25690,N_25028,N_25240);
nand U25691 (N_25691,N_25181,N_25036);
nor U25692 (N_25692,N_25427,N_25476);
xor U25693 (N_25693,N_25442,N_25172);
nor U25694 (N_25694,N_25158,N_25070);
nor U25695 (N_25695,N_25288,N_25336);
nand U25696 (N_25696,N_25092,N_25340);
and U25697 (N_25697,N_25362,N_25031);
nor U25698 (N_25698,N_25322,N_25052);
or U25699 (N_25699,N_25005,N_25341);
and U25700 (N_25700,N_25267,N_25182);
nor U25701 (N_25701,N_25481,N_25282);
and U25702 (N_25702,N_25353,N_25011);
nor U25703 (N_25703,N_25393,N_25187);
xnor U25704 (N_25704,N_25034,N_25100);
xnor U25705 (N_25705,N_25456,N_25003);
or U25706 (N_25706,N_25318,N_25441);
xor U25707 (N_25707,N_25115,N_25296);
xnor U25708 (N_25708,N_25280,N_25046);
nor U25709 (N_25709,N_25401,N_25103);
xor U25710 (N_25710,N_25106,N_25405);
nand U25711 (N_25711,N_25037,N_25258);
nor U25712 (N_25712,N_25169,N_25160);
or U25713 (N_25713,N_25140,N_25069);
nor U25714 (N_25714,N_25479,N_25451);
or U25715 (N_25715,N_25406,N_25475);
nor U25716 (N_25716,N_25320,N_25019);
and U25717 (N_25717,N_25024,N_25178);
or U25718 (N_25718,N_25127,N_25397);
and U25719 (N_25719,N_25429,N_25122);
xor U25720 (N_25720,N_25171,N_25216);
xnor U25721 (N_25721,N_25023,N_25250);
nor U25722 (N_25722,N_25499,N_25001);
and U25723 (N_25723,N_25287,N_25253);
nor U25724 (N_25724,N_25230,N_25113);
nor U25725 (N_25725,N_25059,N_25021);
and U25726 (N_25726,N_25206,N_25215);
and U25727 (N_25727,N_25377,N_25418);
and U25728 (N_25728,N_25384,N_25237);
nor U25729 (N_25729,N_25008,N_25132);
and U25730 (N_25730,N_25156,N_25328);
nor U25731 (N_25731,N_25141,N_25324);
nor U25732 (N_25732,N_25119,N_25039);
or U25733 (N_25733,N_25174,N_25449);
nor U25734 (N_25734,N_25134,N_25307);
nand U25735 (N_25735,N_25063,N_25065);
nor U25736 (N_25736,N_25431,N_25430);
nand U25737 (N_25737,N_25032,N_25457);
or U25738 (N_25738,N_25218,N_25390);
xnor U25739 (N_25739,N_25313,N_25093);
and U25740 (N_25740,N_25349,N_25347);
nor U25741 (N_25741,N_25235,N_25191);
and U25742 (N_25742,N_25163,N_25355);
xnor U25743 (N_25743,N_25189,N_25145);
or U25744 (N_25744,N_25095,N_25201);
nand U25745 (N_25745,N_25153,N_25269);
nor U25746 (N_25746,N_25121,N_25472);
xor U25747 (N_25747,N_25319,N_25292);
or U25748 (N_25748,N_25388,N_25195);
or U25749 (N_25749,N_25466,N_25283);
or U25750 (N_25750,N_25351,N_25394);
xor U25751 (N_25751,N_25128,N_25024);
nor U25752 (N_25752,N_25319,N_25412);
xor U25753 (N_25753,N_25356,N_25190);
nor U25754 (N_25754,N_25494,N_25313);
nand U25755 (N_25755,N_25231,N_25112);
or U25756 (N_25756,N_25439,N_25405);
nand U25757 (N_25757,N_25387,N_25051);
nand U25758 (N_25758,N_25476,N_25249);
xnor U25759 (N_25759,N_25186,N_25258);
or U25760 (N_25760,N_25475,N_25284);
nor U25761 (N_25761,N_25259,N_25261);
nand U25762 (N_25762,N_25493,N_25268);
or U25763 (N_25763,N_25332,N_25272);
and U25764 (N_25764,N_25202,N_25223);
and U25765 (N_25765,N_25454,N_25411);
nand U25766 (N_25766,N_25257,N_25153);
nand U25767 (N_25767,N_25204,N_25170);
or U25768 (N_25768,N_25178,N_25346);
nand U25769 (N_25769,N_25359,N_25243);
and U25770 (N_25770,N_25302,N_25223);
and U25771 (N_25771,N_25483,N_25280);
nand U25772 (N_25772,N_25162,N_25231);
or U25773 (N_25773,N_25466,N_25262);
nand U25774 (N_25774,N_25104,N_25205);
nand U25775 (N_25775,N_25427,N_25458);
xor U25776 (N_25776,N_25042,N_25467);
xor U25777 (N_25777,N_25129,N_25144);
xor U25778 (N_25778,N_25092,N_25041);
nor U25779 (N_25779,N_25487,N_25241);
xor U25780 (N_25780,N_25375,N_25201);
or U25781 (N_25781,N_25160,N_25040);
or U25782 (N_25782,N_25186,N_25464);
nand U25783 (N_25783,N_25095,N_25445);
and U25784 (N_25784,N_25381,N_25198);
or U25785 (N_25785,N_25288,N_25185);
xnor U25786 (N_25786,N_25487,N_25385);
nand U25787 (N_25787,N_25023,N_25138);
nand U25788 (N_25788,N_25304,N_25142);
or U25789 (N_25789,N_25363,N_25243);
xor U25790 (N_25790,N_25004,N_25044);
nand U25791 (N_25791,N_25279,N_25478);
xnor U25792 (N_25792,N_25377,N_25349);
and U25793 (N_25793,N_25281,N_25178);
nand U25794 (N_25794,N_25189,N_25462);
and U25795 (N_25795,N_25174,N_25384);
and U25796 (N_25796,N_25375,N_25172);
nand U25797 (N_25797,N_25145,N_25047);
nor U25798 (N_25798,N_25080,N_25194);
and U25799 (N_25799,N_25320,N_25059);
xnor U25800 (N_25800,N_25159,N_25343);
and U25801 (N_25801,N_25412,N_25073);
and U25802 (N_25802,N_25064,N_25365);
nor U25803 (N_25803,N_25390,N_25253);
nor U25804 (N_25804,N_25288,N_25405);
xnor U25805 (N_25805,N_25147,N_25442);
and U25806 (N_25806,N_25426,N_25176);
and U25807 (N_25807,N_25485,N_25113);
nor U25808 (N_25808,N_25106,N_25321);
nor U25809 (N_25809,N_25132,N_25070);
nor U25810 (N_25810,N_25078,N_25457);
or U25811 (N_25811,N_25163,N_25016);
and U25812 (N_25812,N_25000,N_25199);
and U25813 (N_25813,N_25265,N_25196);
xnor U25814 (N_25814,N_25365,N_25158);
and U25815 (N_25815,N_25253,N_25413);
and U25816 (N_25816,N_25129,N_25310);
xor U25817 (N_25817,N_25338,N_25047);
or U25818 (N_25818,N_25342,N_25227);
nor U25819 (N_25819,N_25085,N_25039);
xor U25820 (N_25820,N_25409,N_25406);
xnor U25821 (N_25821,N_25258,N_25187);
and U25822 (N_25822,N_25261,N_25024);
or U25823 (N_25823,N_25349,N_25241);
nand U25824 (N_25824,N_25386,N_25464);
nor U25825 (N_25825,N_25167,N_25465);
nand U25826 (N_25826,N_25474,N_25403);
xnor U25827 (N_25827,N_25435,N_25343);
nor U25828 (N_25828,N_25028,N_25153);
nor U25829 (N_25829,N_25003,N_25235);
nor U25830 (N_25830,N_25239,N_25164);
and U25831 (N_25831,N_25182,N_25265);
nand U25832 (N_25832,N_25395,N_25166);
and U25833 (N_25833,N_25224,N_25068);
or U25834 (N_25834,N_25020,N_25388);
xnor U25835 (N_25835,N_25035,N_25359);
xor U25836 (N_25836,N_25167,N_25495);
or U25837 (N_25837,N_25489,N_25081);
xor U25838 (N_25838,N_25272,N_25044);
xor U25839 (N_25839,N_25361,N_25275);
nand U25840 (N_25840,N_25315,N_25120);
or U25841 (N_25841,N_25002,N_25480);
nor U25842 (N_25842,N_25127,N_25031);
xnor U25843 (N_25843,N_25148,N_25466);
or U25844 (N_25844,N_25338,N_25251);
nor U25845 (N_25845,N_25194,N_25461);
or U25846 (N_25846,N_25155,N_25243);
nor U25847 (N_25847,N_25166,N_25250);
xor U25848 (N_25848,N_25105,N_25334);
xnor U25849 (N_25849,N_25073,N_25183);
and U25850 (N_25850,N_25297,N_25290);
nor U25851 (N_25851,N_25378,N_25003);
or U25852 (N_25852,N_25101,N_25121);
nand U25853 (N_25853,N_25219,N_25113);
nand U25854 (N_25854,N_25360,N_25081);
nor U25855 (N_25855,N_25128,N_25325);
xor U25856 (N_25856,N_25140,N_25087);
nor U25857 (N_25857,N_25186,N_25469);
and U25858 (N_25858,N_25405,N_25180);
or U25859 (N_25859,N_25138,N_25452);
nand U25860 (N_25860,N_25128,N_25383);
and U25861 (N_25861,N_25015,N_25211);
and U25862 (N_25862,N_25090,N_25332);
nand U25863 (N_25863,N_25466,N_25428);
and U25864 (N_25864,N_25105,N_25031);
nand U25865 (N_25865,N_25343,N_25123);
nand U25866 (N_25866,N_25478,N_25117);
or U25867 (N_25867,N_25297,N_25065);
nor U25868 (N_25868,N_25435,N_25312);
or U25869 (N_25869,N_25103,N_25106);
and U25870 (N_25870,N_25475,N_25061);
and U25871 (N_25871,N_25180,N_25226);
and U25872 (N_25872,N_25432,N_25482);
and U25873 (N_25873,N_25064,N_25392);
nand U25874 (N_25874,N_25315,N_25230);
nor U25875 (N_25875,N_25426,N_25379);
or U25876 (N_25876,N_25018,N_25394);
nor U25877 (N_25877,N_25039,N_25270);
and U25878 (N_25878,N_25281,N_25184);
or U25879 (N_25879,N_25017,N_25185);
or U25880 (N_25880,N_25259,N_25304);
and U25881 (N_25881,N_25349,N_25482);
or U25882 (N_25882,N_25242,N_25056);
or U25883 (N_25883,N_25376,N_25435);
nor U25884 (N_25884,N_25463,N_25347);
xnor U25885 (N_25885,N_25055,N_25215);
xnor U25886 (N_25886,N_25348,N_25146);
nor U25887 (N_25887,N_25000,N_25370);
nand U25888 (N_25888,N_25405,N_25376);
or U25889 (N_25889,N_25115,N_25341);
nand U25890 (N_25890,N_25219,N_25143);
and U25891 (N_25891,N_25493,N_25414);
nor U25892 (N_25892,N_25357,N_25173);
and U25893 (N_25893,N_25256,N_25358);
or U25894 (N_25894,N_25439,N_25164);
or U25895 (N_25895,N_25346,N_25169);
nand U25896 (N_25896,N_25403,N_25049);
and U25897 (N_25897,N_25473,N_25057);
and U25898 (N_25898,N_25439,N_25493);
nor U25899 (N_25899,N_25225,N_25353);
nor U25900 (N_25900,N_25155,N_25025);
or U25901 (N_25901,N_25053,N_25083);
nor U25902 (N_25902,N_25099,N_25093);
and U25903 (N_25903,N_25132,N_25184);
nor U25904 (N_25904,N_25273,N_25433);
xnor U25905 (N_25905,N_25145,N_25078);
nor U25906 (N_25906,N_25056,N_25129);
xor U25907 (N_25907,N_25260,N_25167);
and U25908 (N_25908,N_25274,N_25491);
or U25909 (N_25909,N_25373,N_25297);
nand U25910 (N_25910,N_25491,N_25424);
nand U25911 (N_25911,N_25230,N_25257);
nand U25912 (N_25912,N_25022,N_25275);
nor U25913 (N_25913,N_25148,N_25152);
or U25914 (N_25914,N_25350,N_25072);
nor U25915 (N_25915,N_25403,N_25428);
nor U25916 (N_25916,N_25141,N_25448);
nor U25917 (N_25917,N_25007,N_25442);
or U25918 (N_25918,N_25306,N_25159);
or U25919 (N_25919,N_25310,N_25264);
or U25920 (N_25920,N_25026,N_25387);
or U25921 (N_25921,N_25022,N_25270);
and U25922 (N_25922,N_25287,N_25093);
or U25923 (N_25923,N_25428,N_25172);
and U25924 (N_25924,N_25436,N_25310);
nor U25925 (N_25925,N_25067,N_25156);
xor U25926 (N_25926,N_25008,N_25186);
and U25927 (N_25927,N_25216,N_25065);
and U25928 (N_25928,N_25240,N_25130);
nand U25929 (N_25929,N_25461,N_25306);
xnor U25930 (N_25930,N_25149,N_25296);
nand U25931 (N_25931,N_25372,N_25465);
and U25932 (N_25932,N_25218,N_25055);
nand U25933 (N_25933,N_25489,N_25089);
nor U25934 (N_25934,N_25387,N_25024);
xor U25935 (N_25935,N_25180,N_25455);
and U25936 (N_25936,N_25055,N_25184);
and U25937 (N_25937,N_25017,N_25228);
or U25938 (N_25938,N_25397,N_25451);
and U25939 (N_25939,N_25478,N_25047);
xor U25940 (N_25940,N_25034,N_25060);
or U25941 (N_25941,N_25261,N_25268);
nand U25942 (N_25942,N_25461,N_25391);
or U25943 (N_25943,N_25314,N_25442);
nand U25944 (N_25944,N_25208,N_25261);
xnor U25945 (N_25945,N_25258,N_25252);
nand U25946 (N_25946,N_25101,N_25354);
and U25947 (N_25947,N_25342,N_25142);
nor U25948 (N_25948,N_25047,N_25310);
xor U25949 (N_25949,N_25447,N_25180);
and U25950 (N_25950,N_25438,N_25453);
xnor U25951 (N_25951,N_25086,N_25434);
nand U25952 (N_25952,N_25002,N_25038);
and U25953 (N_25953,N_25303,N_25029);
nor U25954 (N_25954,N_25487,N_25203);
and U25955 (N_25955,N_25051,N_25300);
xor U25956 (N_25956,N_25273,N_25055);
nand U25957 (N_25957,N_25423,N_25361);
nor U25958 (N_25958,N_25157,N_25302);
xnor U25959 (N_25959,N_25393,N_25250);
xor U25960 (N_25960,N_25034,N_25485);
xnor U25961 (N_25961,N_25462,N_25149);
or U25962 (N_25962,N_25213,N_25126);
nor U25963 (N_25963,N_25437,N_25025);
nand U25964 (N_25964,N_25223,N_25385);
or U25965 (N_25965,N_25138,N_25106);
and U25966 (N_25966,N_25160,N_25489);
and U25967 (N_25967,N_25066,N_25405);
xor U25968 (N_25968,N_25213,N_25425);
nand U25969 (N_25969,N_25123,N_25361);
nor U25970 (N_25970,N_25455,N_25280);
xor U25971 (N_25971,N_25418,N_25480);
or U25972 (N_25972,N_25198,N_25020);
nand U25973 (N_25973,N_25295,N_25458);
xnor U25974 (N_25974,N_25250,N_25213);
and U25975 (N_25975,N_25038,N_25385);
and U25976 (N_25976,N_25257,N_25488);
or U25977 (N_25977,N_25114,N_25323);
nor U25978 (N_25978,N_25312,N_25438);
nand U25979 (N_25979,N_25292,N_25148);
nor U25980 (N_25980,N_25203,N_25236);
or U25981 (N_25981,N_25497,N_25088);
xor U25982 (N_25982,N_25472,N_25193);
nand U25983 (N_25983,N_25326,N_25170);
nand U25984 (N_25984,N_25034,N_25468);
nor U25985 (N_25985,N_25062,N_25091);
nand U25986 (N_25986,N_25464,N_25183);
or U25987 (N_25987,N_25008,N_25253);
xnor U25988 (N_25988,N_25227,N_25217);
nor U25989 (N_25989,N_25466,N_25257);
and U25990 (N_25990,N_25062,N_25356);
nand U25991 (N_25991,N_25306,N_25012);
and U25992 (N_25992,N_25269,N_25329);
xnor U25993 (N_25993,N_25361,N_25286);
or U25994 (N_25994,N_25165,N_25070);
and U25995 (N_25995,N_25489,N_25397);
nor U25996 (N_25996,N_25040,N_25153);
and U25997 (N_25997,N_25125,N_25020);
and U25998 (N_25998,N_25138,N_25098);
or U25999 (N_25999,N_25477,N_25381);
and U26000 (N_26000,N_25810,N_25596);
or U26001 (N_26001,N_25694,N_25865);
nor U26002 (N_26002,N_25803,N_25580);
or U26003 (N_26003,N_25912,N_25748);
xor U26004 (N_26004,N_25907,N_25847);
or U26005 (N_26005,N_25636,N_25609);
and U26006 (N_26006,N_25549,N_25853);
nor U26007 (N_26007,N_25929,N_25544);
and U26008 (N_26008,N_25894,N_25872);
nor U26009 (N_26009,N_25736,N_25526);
nand U26010 (N_26010,N_25588,N_25584);
nor U26011 (N_26011,N_25813,N_25652);
or U26012 (N_26012,N_25574,N_25552);
nand U26013 (N_26013,N_25648,N_25505);
nor U26014 (N_26014,N_25858,N_25619);
or U26015 (N_26015,N_25524,N_25687);
and U26016 (N_26016,N_25901,N_25510);
xnor U26017 (N_26017,N_25969,N_25674);
or U26018 (N_26018,N_25825,N_25599);
nand U26019 (N_26019,N_25627,N_25991);
or U26020 (N_26020,N_25891,N_25795);
nand U26021 (N_26021,N_25954,N_25709);
and U26022 (N_26022,N_25774,N_25973);
nand U26023 (N_26023,N_25508,N_25855);
and U26024 (N_26024,N_25946,N_25521);
xnor U26025 (N_26025,N_25809,N_25911);
xor U26026 (N_26026,N_25504,N_25949);
nor U26027 (N_26027,N_25913,N_25697);
or U26028 (N_26028,N_25646,N_25644);
and U26029 (N_26029,N_25523,N_25534);
xor U26030 (N_26030,N_25728,N_25650);
nor U26031 (N_26031,N_25570,N_25689);
xor U26032 (N_26032,N_25794,N_25867);
xor U26033 (N_26033,N_25886,N_25895);
and U26034 (N_26034,N_25958,N_25616);
nor U26035 (N_26035,N_25666,N_25569);
and U26036 (N_26036,N_25718,N_25827);
xnor U26037 (N_26037,N_25525,N_25967);
or U26038 (N_26038,N_25922,N_25975);
or U26039 (N_26039,N_25793,N_25714);
xor U26040 (N_26040,N_25642,N_25920);
xnor U26041 (N_26041,N_25826,N_25581);
nand U26042 (N_26042,N_25963,N_25814);
nand U26043 (N_26043,N_25577,N_25861);
or U26044 (N_26044,N_25961,N_25928);
or U26045 (N_26045,N_25941,N_25741);
nor U26046 (N_26046,N_25818,N_25766);
and U26047 (N_26047,N_25993,N_25927);
nor U26048 (N_26048,N_25600,N_25799);
xnor U26049 (N_26049,N_25885,N_25686);
nand U26050 (N_26050,N_25702,N_25805);
and U26051 (N_26051,N_25645,N_25760);
or U26052 (N_26052,N_25880,N_25532);
xor U26053 (N_26053,N_25528,N_25535);
nand U26054 (N_26054,N_25683,N_25955);
nand U26055 (N_26055,N_25623,N_25639);
xnor U26056 (N_26056,N_25943,N_25960);
or U26057 (N_26057,N_25664,N_25789);
xnor U26058 (N_26058,N_25732,N_25801);
nor U26059 (N_26059,N_25933,N_25835);
nor U26060 (N_26060,N_25904,N_25785);
nand U26061 (N_26061,N_25918,N_25866);
xor U26062 (N_26062,N_25707,N_25703);
nand U26063 (N_26063,N_25680,N_25654);
or U26064 (N_26064,N_25565,N_25796);
and U26065 (N_26065,N_25653,N_25804);
xnor U26066 (N_26066,N_25840,N_25914);
nor U26067 (N_26067,N_25724,N_25873);
or U26068 (N_26068,N_25883,N_25613);
and U26069 (N_26069,N_25677,N_25790);
and U26070 (N_26070,N_25773,N_25690);
nor U26071 (N_26071,N_25828,N_25771);
xnor U26072 (N_26072,N_25806,N_25556);
xor U26073 (N_26073,N_25632,N_25625);
nor U26074 (N_26074,N_25781,N_25745);
xor U26075 (N_26075,N_25778,N_25529);
xor U26076 (N_26076,N_25947,N_25734);
and U26077 (N_26077,N_25667,N_25782);
nor U26078 (N_26078,N_25624,N_25746);
and U26079 (N_26079,N_25554,N_25601);
xnor U26080 (N_26080,N_25696,N_25906);
or U26081 (N_26081,N_25519,N_25550);
xnor U26082 (N_26082,N_25862,N_25669);
and U26083 (N_26083,N_25575,N_25698);
nor U26084 (N_26084,N_25989,N_25910);
nand U26085 (N_26085,N_25936,N_25889);
nand U26086 (N_26086,N_25935,N_25968);
or U26087 (N_26087,N_25990,N_25843);
nand U26088 (N_26088,N_25672,N_25731);
or U26089 (N_26089,N_25590,N_25541);
xnor U26090 (N_26090,N_25682,N_25940);
and U26091 (N_26091,N_25607,N_25545);
nand U26092 (N_26092,N_25708,N_25548);
xnor U26093 (N_26093,N_25939,N_25717);
nand U26094 (N_26094,N_25994,N_25953);
and U26095 (N_26095,N_25945,N_25573);
and U26096 (N_26096,N_25921,N_25699);
or U26097 (N_26097,N_25739,N_25908);
nor U26098 (N_26098,N_25846,N_25629);
and U26099 (N_26099,N_25950,N_25660);
or U26100 (N_26100,N_25919,N_25513);
nor U26101 (N_26101,N_25617,N_25924);
or U26102 (N_26102,N_25860,N_25807);
nor U26103 (N_26103,N_25753,N_25876);
nand U26104 (N_26104,N_25592,N_25621);
nor U26105 (N_26105,N_25610,N_25603);
and U26106 (N_26106,N_25633,N_25637);
nand U26107 (N_26107,N_25761,N_25604);
and U26108 (N_26108,N_25770,N_25563);
nand U26109 (N_26109,N_25558,N_25579);
nand U26110 (N_26110,N_25932,N_25605);
xor U26111 (N_26111,N_25859,N_25676);
or U26112 (N_26112,N_25530,N_25608);
xnor U26113 (N_26113,N_25780,N_25839);
xor U26114 (N_26114,N_25792,N_25874);
xnor U26115 (N_26115,N_25965,N_25980);
or U26116 (N_26116,N_25852,N_25663);
nand U26117 (N_26117,N_25537,N_25593);
and U26118 (N_26118,N_25899,N_25705);
nand U26119 (N_26119,N_25713,N_25546);
xnor U26120 (N_26120,N_25972,N_25767);
xor U26121 (N_26121,N_25568,N_25985);
nand U26122 (N_26122,N_25959,N_25501);
nand U26123 (N_26123,N_25995,N_25871);
or U26124 (N_26124,N_25597,N_25540);
nand U26125 (N_26125,N_25777,N_25884);
nor U26126 (N_26126,N_25834,N_25842);
and U26127 (N_26127,N_25618,N_25512);
or U26128 (N_26128,N_25916,N_25726);
nor U26129 (N_26129,N_25752,N_25854);
nand U26130 (N_26130,N_25543,N_25557);
nand U26131 (N_26131,N_25514,N_25576);
nor U26132 (N_26132,N_25509,N_25786);
and U26133 (N_26133,N_25555,N_25531);
nand U26134 (N_26134,N_25634,N_25812);
nand U26135 (N_26135,N_25668,N_25851);
or U26136 (N_26136,N_25938,N_25882);
xnor U26137 (N_26137,N_25800,N_25720);
xor U26138 (N_26138,N_25776,N_25900);
xnor U26139 (N_26139,N_25595,N_25863);
xor U26140 (N_26140,N_25520,N_25598);
nand U26141 (N_26141,N_25832,N_25542);
nand U26142 (N_26142,N_25533,N_25983);
xor U26143 (N_26143,N_25631,N_25643);
nand U26144 (N_26144,N_25749,N_25759);
nand U26145 (N_26145,N_25905,N_25561);
xor U26146 (N_26146,N_25536,N_25651);
nand U26147 (N_26147,N_25931,N_25744);
nor U26148 (N_26148,N_25925,N_25944);
or U26149 (N_26149,N_25638,N_25516);
nor U26150 (N_26150,N_25567,N_25869);
and U26151 (N_26151,N_25763,N_25611);
or U26152 (N_26152,N_25503,N_25849);
nand U26153 (N_26153,N_25999,N_25831);
and U26154 (N_26154,N_25656,N_25723);
nand U26155 (N_26155,N_25978,N_25671);
xor U26156 (N_26156,N_25845,N_25507);
nor U26157 (N_26157,N_25578,N_25754);
nor U26158 (N_26158,N_25964,N_25971);
nor U26159 (N_26159,N_25640,N_25979);
nand U26160 (N_26160,N_25691,N_25998);
nand U26161 (N_26161,N_25956,N_25517);
or U26162 (N_26162,N_25755,N_25515);
or U26163 (N_26163,N_25952,N_25737);
nand U26164 (N_26164,N_25547,N_25879);
nor U26165 (N_26165,N_25934,N_25620);
nor U26166 (N_26166,N_25583,N_25915);
nor U26167 (N_26167,N_25688,N_25791);
nor U26168 (N_26168,N_25996,N_25822);
nor U26169 (N_26169,N_25974,N_25841);
nor U26170 (N_26170,N_25711,N_25838);
xnor U26171 (N_26171,N_25875,N_25738);
xor U26172 (N_26172,N_25630,N_25909);
xnor U26173 (N_26173,N_25566,N_25772);
and U26174 (N_26174,N_25788,N_25562);
xnor U26175 (N_26175,N_25837,N_25783);
nor U26176 (N_26176,N_25977,N_25997);
nor U26177 (N_26177,N_25937,N_25787);
or U26178 (N_26178,N_25559,N_25665);
and U26179 (N_26179,N_25798,N_25779);
nor U26180 (N_26180,N_25982,N_25864);
xor U26181 (N_26181,N_25585,N_25743);
nand U26182 (N_26182,N_25701,N_25870);
and U26183 (N_26183,N_25888,N_25684);
nor U26184 (N_26184,N_25902,N_25970);
or U26185 (N_26185,N_25655,N_25661);
nor U26186 (N_26186,N_25551,N_25823);
xnor U26187 (N_26187,N_25716,N_25802);
nor U26188 (N_26188,N_25948,N_25820);
and U26189 (N_26189,N_25887,N_25729);
nor U26190 (N_26190,N_25984,N_25722);
nor U26191 (N_26191,N_25681,N_25502);
and U26192 (N_26192,N_25962,N_25976);
nand U26193 (N_26193,N_25930,N_25700);
or U26194 (N_26194,N_25710,N_25735);
or U26195 (N_26195,N_25647,N_25819);
nor U26196 (N_26196,N_25942,N_25742);
xnor U26197 (N_26197,N_25797,N_25923);
nor U26198 (N_26198,N_25612,N_25721);
nand U26199 (N_26199,N_25560,N_25527);
nand U26200 (N_26200,N_25649,N_25750);
or U26201 (N_26201,N_25951,N_25917);
nand U26202 (N_26202,N_25988,N_25641);
nand U26203 (N_26203,N_25893,N_25675);
nand U26204 (N_26204,N_25817,N_25615);
xnor U26205 (N_26205,N_25992,N_25815);
or U26206 (N_26206,N_25582,N_25733);
nand U26207 (N_26207,N_25898,N_25572);
nand U26208 (N_26208,N_25758,N_25811);
and U26209 (N_26209,N_25821,N_25719);
xnor U26210 (N_26210,N_25844,N_25829);
or U26211 (N_26211,N_25659,N_25878);
nand U26212 (N_26212,N_25606,N_25926);
or U26213 (N_26213,N_25725,N_25986);
nand U26214 (N_26214,N_25538,N_25764);
xor U26215 (N_26215,N_25727,N_25594);
or U26216 (N_26216,N_25553,N_25635);
nor U26217 (N_26217,N_25957,N_25704);
nand U26218 (N_26218,N_25903,N_25614);
nand U26219 (N_26219,N_25673,N_25981);
or U26220 (N_26220,N_25715,N_25836);
xor U26221 (N_26221,N_25518,N_25706);
xnor U26222 (N_26222,N_25877,N_25757);
and U26223 (N_26223,N_25626,N_25522);
or U26224 (N_26224,N_25587,N_25768);
nand U26225 (N_26225,N_25586,N_25564);
nor U26226 (N_26226,N_25685,N_25856);
and U26227 (N_26227,N_25657,N_25966);
and U26228 (N_26228,N_25622,N_25511);
nor U26229 (N_26229,N_25987,N_25602);
nand U26230 (N_26230,N_25775,N_25848);
xnor U26231 (N_26231,N_25881,N_25506);
and U26232 (N_26232,N_25712,N_25784);
and U26233 (N_26233,N_25695,N_25896);
nor U26234 (N_26234,N_25740,N_25892);
xnor U26235 (N_26235,N_25678,N_25658);
xor U26236 (N_26236,N_25693,N_25816);
xnor U26237 (N_26237,N_25571,N_25762);
nand U26238 (N_26238,N_25628,N_25662);
and U26239 (N_26239,N_25500,N_25591);
and U26240 (N_26240,N_25679,N_25692);
and U26241 (N_26241,N_25857,N_25824);
nand U26242 (N_26242,N_25539,N_25747);
nor U26243 (N_26243,N_25730,N_25756);
and U26244 (N_26244,N_25670,N_25769);
nor U26245 (N_26245,N_25830,N_25589);
and U26246 (N_26246,N_25765,N_25751);
nand U26247 (N_26247,N_25868,N_25850);
and U26248 (N_26248,N_25808,N_25833);
nor U26249 (N_26249,N_25897,N_25890);
nor U26250 (N_26250,N_25740,N_25711);
nor U26251 (N_26251,N_25627,N_25893);
and U26252 (N_26252,N_25589,N_25728);
and U26253 (N_26253,N_25609,N_25627);
nand U26254 (N_26254,N_25655,N_25985);
nor U26255 (N_26255,N_25893,N_25608);
and U26256 (N_26256,N_25843,N_25724);
nand U26257 (N_26257,N_25670,N_25971);
nand U26258 (N_26258,N_25671,N_25931);
or U26259 (N_26259,N_25503,N_25947);
nand U26260 (N_26260,N_25717,N_25913);
or U26261 (N_26261,N_25938,N_25809);
nand U26262 (N_26262,N_25663,N_25997);
or U26263 (N_26263,N_25925,N_25834);
nand U26264 (N_26264,N_25526,N_25834);
xor U26265 (N_26265,N_25849,N_25947);
nor U26266 (N_26266,N_25586,N_25691);
and U26267 (N_26267,N_25542,N_25734);
nor U26268 (N_26268,N_25599,N_25849);
xor U26269 (N_26269,N_25801,N_25964);
xnor U26270 (N_26270,N_25677,N_25631);
nand U26271 (N_26271,N_25812,N_25879);
and U26272 (N_26272,N_25924,N_25639);
and U26273 (N_26273,N_25896,N_25701);
or U26274 (N_26274,N_25713,N_25672);
nor U26275 (N_26275,N_25543,N_25843);
or U26276 (N_26276,N_25758,N_25656);
nor U26277 (N_26277,N_25957,N_25716);
and U26278 (N_26278,N_25883,N_25771);
or U26279 (N_26279,N_25742,N_25826);
xor U26280 (N_26280,N_25841,N_25790);
or U26281 (N_26281,N_25616,N_25874);
or U26282 (N_26282,N_25588,N_25962);
xnor U26283 (N_26283,N_25538,N_25766);
and U26284 (N_26284,N_25550,N_25602);
nand U26285 (N_26285,N_25828,N_25731);
nor U26286 (N_26286,N_25889,N_25557);
nor U26287 (N_26287,N_25625,N_25726);
and U26288 (N_26288,N_25999,N_25587);
xor U26289 (N_26289,N_25507,N_25885);
nor U26290 (N_26290,N_25551,N_25860);
and U26291 (N_26291,N_25977,N_25864);
nor U26292 (N_26292,N_25742,N_25930);
nor U26293 (N_26293,N_25700,N_25503);
nand U26294 (N_26294,N_25868,N_25694);
and U26295 (N_26295,N_25946,N_25568);
nor U26296 (N_26296,N_25957,N_25524);
or U26297 (N_26297,N_25963,N_25883);
and U26298 (N_26298,N_25913,N_25516);
or U26299 (N_26299,N_25884,N_25600);
or U26300 (N_26300,N_25762,N_25953);
and U26301 (N_26301,N_25705,N_25626);
and U26302 (N_26302,N_25865,N_25878);
nand U26303 (N_26303,N_25732,N_25879);
and U26304 (N_26304,N_25642,N_25782);
or U26305 (N_26305,N_25712,N_25672);
or U26306 (N_26306,N_25854,N_25888);
nor U26307 (N_26307,N_25858,N_25961);
and U26308 (N_26308,N_25804,N_25933);
or U26309 (N_26309,N_25981,N_25727);
nand U26310 (N_26310,N_25676,N_25609);
nor U26311 (N_26311,N_25745,N_25668);
nor U26312 (N_26312,N_25894,N_25563);
or U26313 (N_26313,N_25724,N_25635);
xor U26314 (N_26314,N_25544,N_25912);
nor U26315 (N_26315,N_25605,N_25871);
and U26316 (N_26316,N_25999,N_25656);
nor U26317 (N_26317,N_25500,N_25504);
nand U26318 (N_26318,N_25790,N_25880);
or U26319 (N_26319,N_25996,N_25670);
or U26320 (N_26320,N_25945,N_25992);
and U26321 (N_26321,N_25977,N_25646);
or U26322 (N_26322,N_25684,N_25928);
nand U26323 (N_26323,N_25828,N_25506);
nor U26324 (N_26324,N_25946,N_25507);
nor U26325 (N_26325,N_25500,N_25633);
xnor U26326 (N_26326,N_25965,N_25648);
nor U26327 (N_26327,N_25527,N_25705);
xnor U26328 (N_26328,N_25899,N_25679);
xor U26329 (N_26329,N_25504,N_25899);
nor U26330 (N_26330,N_25652,N_25922);
or U26331 (N_26331,N_25586,N_25955);
xor U26332 (N_26332,N_25862,N_25633);
or U26333 (N_26333,N_25792,N_25916);
xnor U26334 (N_26334,N_25521,N_25976);
and U26335 (N_26335,N_25604,N_25849);
nand U26336 (N_26336,N_25683,N_25566);
xnor U26337 (N_26337,N_25775,N_25890);
and U26338 (N_26338,N_25957,N_25546);
nand U26339 (N_26339,N_25840,N_25970);
nand U26340 (N_26340,N_25973,N_25806);
nor U26341 (N_26341,N_25996,N_25539);
xnor U26342 (N_26342,N_25657,N_25568);
xnor U26343 (N_26343,N_25673,N_25723);
or U26344 (N_26344,N_25833,N_25937);
and U26345 (N_26345,N_25699,N_25790);
nor U26346 (N_26346,N_25913,N_25712);
nand U26347 (N_26347,N_25619,N_25568);
nor U26348 (N_26348,N_25914,N_25568);
xnor U26349 (N_26349,N_25935,N_25956);
nand U26350 (N_26350,N_25504,N_25805);
and U26351 (N_26351,N_25663,N_25524);
nor U26352 (N_26352,N_25712,N_25703);
nor U26353 (N_26353,N_25948,N_25714);
nor U26354 (N_26354,N_25563,N_25517);
or U26355 (N_26355,N_25949,N_25853);
xor U26356 (N_26356,N_25779,N_25664);
or U26357 (N_26357,N_25831,N_25979);
and U26358 (N_26358,N_25739,N_25864);
nor U26359 (N_26359,N_25853,N_25803);
nor U26360 (N_26360,N_25614,N_25546);
nor U26361 (N_26361,N_25831,N_25951);
and U26362 (N_26362,N_25702,N_25733);
xor U26363 (N_26363,N_25988,N_25905);
xor U26364 (N_26364,N_25865,N_25743);
xnor U26365 (N_26365,N_25572,N_25975);
and U26366 (N_26366,N_25599,N_25703);
nor U26367 (N_26367,N_25816,N_25631);
nand U26368 (N_26368,N_25995,N_25854);
nand U26369 (N_26369,N_25964,N_25812);
nor U26370 (N_26370,N_25539,N_25597);
xor U26371 (N_26371,N_25568,N_25978);
and U26372 (N_26372,N_25613,N_25925);
nand U26373 (N_26373,N_25779,N_25616);
nand U26374 (N_26374,N_25685,N_25908);
nand U26375 (N_26375,N_25561,N_25568);
nand U26376 (N_26376,N_25796,N_25951);
and U26377 (N_26377,N_25675,N_25936);
nor U26378 (N_26378,N_25970,N_25720);
and U26379 (N_26379,N_25520,N_25825);
nor U26380 (N_26380,N_25938,N_25562);
nand U26381 (N_26381,N_25534,N_25944);
xor U26382 (N_26382,N_25788,N_25672);
or U26383 (N_26383,N_25768,N_25556);
xor U26384 (N_26384,N_25524,N_25629);
nand U26385 (N_26385,N_25916,N_25602);
nor U26386 (N_26386,N_25769,N_25795);
or U26387 (N_26387,N_25705,N_25500);
xnor U26388 (N_26388,N_25901,N_25852);
nor U26389 (N_26389,N_25972,N_25538);
or U26390 (N_26390,N_25868,N_25543);
xor U26391 (N_26391,N_25610,N_25706);
xnor U26392 (N_26392,N_25721,N_25889);
nor U26393 (N_26393,N_25629,N_25559);
xor U26394 (N_26394,N_25723,N_25684);
or U26395 (N_26395,N_25567,N_25727);
or U26396 (N_26396,N_25958,N_25949);
or U26397 (N_26397,N_25742,N_25642);
xnor U26398 (N_26398,N_25923,N_25824);
nor U26399 (N_26399,N_25897,N_25791);
nand U26400 (N_26400,N_25506,N_25620);
or U26401 (N_26401,N_25950,N_25612);
and U26402 (N_26402,N_25515,N_25511);
nand U26403 (N_26403,N_25709,N_25804);
or U26404 (N_26404,N_25517,N_25531);
nand U26405 (N_26405,N_25685,N_25837);
or U26406 (N_26406,N_25717,N_25843);
nand U26407 (N_26407,N_25811,N_25722);
and U26408 (N_26408,N_25520,N_25596);
and U26409 (N_26409,N_25952,N_25981);
xor U26410 (N_26410,N_25815,N_25929);
xor U26411 (N_26411,N_25771,N_25520);
nor U26412 (N_26412,N_25505,N_25625);
nand U26413 (N_26413,N_25765,N_25703);
and U26414 (N_26414,N_25728,N_25956);
or U26415 (N_26415,N_25850,N_25590);
and U26416 (N_26416,N_25931,N_25894);
nor U26417 (N_26417,N_25729,N_25614);
or U26418 (N_26418,N_25549,N_25798);
or U26419 (N_26419,N_25690,N_25863);
or U26420 (N_26420,N_25974,N_25689);
nor U26421 (N_26421,N_25686,N_25594);
nand U26422 (N_26422,N_25900,N_25864);
nor U26423 (N_26423,N_25621,N_25669);
xor U26424 (N_26424,N_25659,N_25689);
or U26425 (N_26425,N_25889,N_25582);
xor U26426 (N_26426,N_25914,N_25524);
or U26427 (N_26427,N_25535,N_25764);
nand U26428 (N_26428,N_25673,N_25953);
or U26429 (N_26429,N_25917,N_25701);
xnor U26430 (N_26430,N_25898,N_25989);
or U26431 (N_26431,N_25989,N_25506);
nand U26432 (N_26432,N_25868,N_25955);
nand U26433 (N_26433,N_25616,N_25676);
nand U26434 (N_26434,N_25902,N_25616);
xor U26435 (N_26435,N_25524,N_25871);
nand U26436 (N_26436,N_25706,N_25870);
xor U26437 (N_26437,N_25721,N_25782);
nand U26438 (N_26438,N_25592,N_25658);
nor U26439 (N_26439,N_25948,N_25823);
xnor U26440 (N_26440,N_25945,N_25644);
or U26441 (N_26441,N_25642,N_25627);
xor U26442 (N_26442,N_25798,N_25929);
nand U26443 (N_26443,N_25617,N_25879);
nand U26444 (N_26444,N_25759,N_25763);
xnor U26445 (N_26445,N_25864,N_25842);
nor U26446 (N_26446,N_25963,N_25615);
nor U26447 (N_26447,N_25573,N_25944);
and U26448 (N_26448,N_25978,N_25525);
nor U26449 (N_26449,N_25876,N_25744);
nor U26450 (N_26450,N_25825,N_25909);
and U26451 (N_26451,N_25611,N_25700);
xnor U26452 (N_26452,N_25907,N_25706);
xor U26453 (N_26453,N_25620,N_25553);
nand U26454 (N_26454,N_25725,N_25583);
or U26455 (N_26455,N_25971,N_25763);
xnor U26456 (N_26456,N_25609,N_25624);
xnor U26457 (N_26457,N_25604,N_25850);
or U26458 (N_26458,N_25598,N_25948);
nor U26459 (N_26459,N_25665,N_25697);
and U26460 (N_26460,N_25937,N_25706);
and U26461 (N_26461,N_25836,N_25608);
and U26462 (N_26462,N_25866,N_25574);
xnor U26463 (N_26463,N_25742,N_25773);
or U26464 (N_26464,N_25839,N_25657);
or U26465 (N_26465,N_25926,N_25700);
and U26466 (N_26466,N_25529,N_25670);
nand U26467 (N_26467,N_25901,N_25935);
xor U26468 (N_26468,N_25670,N_25554);
or U26469 (N_26469,N_25898,N_25530);
and U26470 (N_26470,N_25606,N_25934);
and U26471 (N_26471,N_25531,N_25699);
xor U26472 (N_26472,N_25829,N_25748);
and U26473 (N_26473,N_25997,N_25517);
nand U26474 (N_26474,N_25654,N_25965);
xor U26475 (N_26475,N_25846,N_25587);
nand U26476 (N_26476,N_25878,N_25722);
or U26477 (N_26477,N_25847,N_25716);
xor U26478 (N_26478,N_25823,N_25881);
and U26479 (N_26479,N_25681,N_25705);
xnor U26480 (N_26480,N_25982,N_25909);
or U26481 (N_26481,N_25822,N_25919);
xor U26482 (N_26482,N_25852,N_25585);
nor U26483 (N_26483,N_25872,N_25856);
nand U26484 (N_26484,N_25887,N_25575);
nor U26485 (N_26485,N_25542,N_25674);
and U26486 (N_26486,N_25949,N_25599);
nand U26487 (N_26487,N_25965,N_25807);
or U26488 (N_26488,N_25824,N_25730);
nand U26489 (N_26489,N_25691,N_25901);
and U26490 (N_26490,N_25642,N_25769);
xnor U26491 (N_26491,N_25875,N_25718);
xnor U26492 (N_26492,N_25979,N_25550);
or U26493 (N_26493,N_25530,N_25534);
or U26494 (N_26494,N_25917,N_25928);
or U26495 (N_26495,N_25552,N_25576);
and U26496 (N_26496,N_25917,N_25576);
xnor U26497 (N_26497,N_25674,N_25622);
or U26498 (N_26498,N_25795,N_25931);
nand U26499 (N_26499,N_25536,N_25574);
and U26500 (N_26500,N_26216,N_26439);
nor U26501 (N_26501,N_26332,N_26090);
nand U26502 (N_26502,N_26402,N_26247);
nor U26503 (N_26503,N_26182,N_26058);
xor U26504 (N_26504,N_26165,N_26436);
and U26505 (N_26505,N_26495,N_26110);
xor U26506 (N_26506,N_26279,N_26043);
nor U26507 (N_26507,N_26105,N_26489);
and U26508 (N_26508,N_26333,N_26361);
or U26509 (N_26509,N_26312,N_26075);
xor U26510 (N_26510,N_26128,N_26218);
nor U26511 (N_26511,N_26240,N_26106);
nor U26512 (N_26512,N_26358,N_26210);
nand U26513 (N_26513,N_26336,N_26377);
or U26514 (N_26514,N_26421,N_26063);
and U26515 (N_26515,N_26397,N_26494);
nand U26516 (N_26516,N_26153,N_26025);
or U26517 (N_26517,N_26124,N_26190);
nor U26518 (N_26518,N_26045,N_26146);
nor U26519 (N_26519,N_26398,N_26406);
and U26520 (N_26520,N_26388,N_26185);
and U26521 (N_26521,N_26301,N_26337);
nand U26522 (N_26522,N_26033,N_26446);
or U26523 (N_26523,N_26457,N_26288);
xor U26524 (N_26524,N_26444,N_26047);
nand U26525 (N_26525,N_26453,N_26331);
nand U26526 (N_26526,N_26098,N_26313);
nand U26527 (N_26527,N_26425,N_26060);
or U26528 (N_26528,N_26262,N_26347);
nor U26529 (N_26529,N_26365,N_26395);
and U26530 (N_26530,N_26121,N_26263);
nand U26531 (N_26531,N_26472,N_26345);
nand U26532 (N_26532,N_26438,N_26178);
and U26533 (N_26533,N_26448,N_26135);
or U26534 (N_26534,N_26102,N_26000);
nor U26535 (N_26535,N_26306,N_26392);
nor U26536 (N_26536,N_26481,N_26271);
or U26537 (N_26537,N_26316,N_26255);
nor U26538 (N_26538,N_26343,N_26074);
nand U26539 (N_26539,N_26173,N_26391);
nand U26540 (N_26540,N_26264,N_26295);
or U26541 (N_26541,N_26242,N_26148);
or U26542 (N_26542,N_26099,N_26249);
and U26543 (N_26543,N_26183,N_26082);
nand U26544 (N_26544,N_26052,N_26428);
nand U26545 (N_26545,N_26408,N_26385);
nand U26546 (N_26546,N_26257,N_26290);
or U26547 (N_26547,N_26204,N_26451);
nor U26548 (N_26548,N_26344,N_26096);
nand U26549 (N_26549,N_26223,N_26077);
or U26550 (N_26550,N_26215,N_26177);
nand U26551 (N_26551,N_26415,N_26433);
or U26552 (N_26552,N_26196,N_26208);
nor U26553 (N_26553,N_26467,N_26318);
nand U26554 (N_26554,N_26474,N_26141);
and U26555 (N_26555,N_26079,N_26284);
nand U26556 (N_26556,N_26325,N_26108);
or U26557 (N_26557,N_26293,N_26246);
and U26558 (N_26558,N_26368,N_26422);
nor U26559 (N_26559,N_26236,N_26285);
xor U26560 (N_26560,N_26364,N_26418);
nand U26561 (N_26561,N_26038,N_26237);
nand U26562 (N_26562,N_26034,N_26107);
and U26563 (N_26563,N_26286,N_26231);
xnor U26564 (N_26564,N_26320,N_26078);
nand U26565 (N_26565,N_26274,N_26125);
nor U26566 (N_26566,N_26412,N_26349);
and U26567 (N_26567,N_26088,N_26036);
or U26568 (N_26568,N_26468,N_26229);
nor U26569 (N_26569,N_26005,N_26241);
nor U26570 (N_26570,N_26384,N_26287);
nand U26571 (N_26571,N_26195,N_26490);
nor U26572 (N_26572,N_26441,N_26219);
or U26573 (N_26573,N_26399,N_26203);
or U26574 (N_26574,N_26035,N_26002);
nor U26575 (N_26575,N_26460,N_26405);
and U26576 (N_26576,N_26319,N_26248);
and U26577 (N_26577,N_26091,N_26134);
nor U26578 (N_26578,N_26062,N_26224);
and U26579 (N_26579,N_26465,N_26167);
or U26580 (N_26580,N_26217,N_26245);
nor U26581 (N_26581,N_26256,N_26056);
nand U26582 (N_26582,N_26054,N_26352);
xor U26583 (N_26583,N_26400,N_26488);
xor U26584 (N_26584,N_26142,N_26123);
nor U26585 (N_26585,N_26206,N_26170);
xor U26586 (N_26586,N_26181,N_26454);
and U26587 (N_26587,N_26278,N_26189);
and U26588 (N_26588,N_26169,N_26371);
xnor U26589 (N_26589,N_26046,N_26150);
or U26590 (N_26590,N_26140,N_26394);
nand U26591 (N_26591,N_26059,N_26073);
xnor U26592 (N_26592,N_26297,N_26423);
xor U26593 (N_26593,N_26314,N_26374);
nor U26594 (N_26594,N_26469,N_26303);
xnor U26595 (N_26595,N_26144,N_26087);
nand U26596 (N_26596,N_26230,N_26066);
nand U26597 (N_26597,N_26067,N_26006);
xor U26598 (N_26598,N_26341,N_26324);
xnor U26599 (N_26599,N_26276,N_26413);
and U26600 (N_26600,N_26235,N_26122);
or U26601 (N_26601,N_26298,N_26281);
and U26602 (N_26602,N_26040,N_26176);
nand U26603 (N_26603,N_26445,N_26008);
xnor U26604 (N_26604,N_26437,N_26267);
xnor U26605 (N_26605,N_26083,N_26338);
and U26606 (N_26606,N_26086,N_26273);
and U26607 (N_26607,N_26458,N_26030);
and U26608 (N_26608,N_26225,N_26021);
nor U26609 (N_26609,N_26419,N_26199);
nor U26610 (N_26610,N_26039,N_26172);
nor U26611 (N_26611,N_26012,N_26139);
nand U26612 (N_26612,N_26243,N_26113);
or U26613 (N_26613,N_26409,N_26100);
nor U26614 (N_26614,N_26156,N_26111);
nand U26615 (N_26615,N_26061,N_26227);
or U26616 (N_26616,N_26147,N_26166);
or U26617 (N_26617,N_26299,N_26456);
or U26618 (N_26618,N_26411,N_26386);
and U26619 (N_26619,N_26292,N_26342);
and U26620 (N_26620,N_26434,N_26270);
and U26621 (N_26621,N_26307,N_26372);
nor U26622 (N_26622,N_26154,N_26003);
nor U26623 (N_26623,N_26202,N_26028);
nand U26624 (N_26624,N_26259,N_26001);
nand U26625 (N_26625,N_26220,N_26127);
nor U26626 (N_26626,N_26426,N_26334);
and U26627 (N_26627,N_26093,N_26376);
nand U26628 (N_26628,N_26404,N_26053);
nand U26629 (N_26629,N_26348,N_26327);
xnor U26630 (N_26630,N_26131,N_26396);
or U26631 (N_26631,N_26390,N_26152);
xnor U26632 (N_26632,N_26353,N_26308);
or U26633 (N_26633,N_26435,N_26209);
or U26634 (N_26634,N_26076,N_26369);
nor U26635 (N_26635,N_26375,N_26023);
nand U26636 (N_26636,N_26484,N_26104);
nor U26637 (N_26637,N_26057,N_26151);
xnor U26638 (N_26638,N_26464,N_26485);
nand U26639 (N_26639,N_26432,N_26186);
or U26640 (N_26640,N_26018,N_26459);
or U26641 (N_26641,N_26269,N_26296);
and U26642 (N_26642,N_26359,N_26115);
xnor U26643 (N_26643,N_26022,N_26470);
or U26644 (N_26644,N_26380,N_26461);
nor U26645 (N_26645,N_26254,N_26410);
and U26646 (N_26646,N_26019,N_26029);
nor U26647 (N_26647,N_26119,N_26252);
nand U26648 (N_26648,N_26085,N_26471);
nand U26649 (N_26649,N_26159,N_26234);
or U26650 (N_26650,N_26447,N_26089);
nand U26651 (N_26651,N_26311,N_26389);
nand U26652 (N_26652,N_26198,N_26265);
and U26653 (N_26653,N_26321,N_26138);
xor U26654 (N_26654,N_26221,N_26226);
nand U26655 (N_26655,N_26149,N_26294);
and U26656 (N_26656,N_26232,N_26009);
nor U26657 (N_26657,N_26260,N_26476);
xnor U26658 (N_26658,N_26462,N_26212);
xnor U26659 (N_26659,N_26103,N_26109);
xor U26660 (N_26660,N_26157,N_26282);
xnor U26661 (N_26661,N_26048,N_26363);
nand U26662 (N_26662,N_26013,N_26163);
and U26663 (N_26663,N_26132,N_26027);
nor U26664 (N_26664,N_26068,N_26133);
or U26665 (N_26665,N_26031,N_26350);
nor U26666 (N_26666,N_26244,N_26486);
and U26667 (N_26667,N_26239,N_26201);
xor U26668 (N_26668,N_26137,N_26492);
or U26669 (N_26669,N_26211,N_26145);
xnor U26670 (N_26670,N_26430,N_26370);
nand U26671 (N_26671,N_26443,N_26401);
and U26672 (N_26672,N_26480,N_26381);
nand U26673 (N_26673,N_26479,N_26112);
and U26674 (N_26674,N_26431,N_26116);
and U26675 (N_26675,N_26072,N_26339);
nand U26676 (N_26676,N_26498,N_26010);
nor U26677 (N_26677,N_26016,N_26097);
or U26678 (N_26678,N_26487,N_26367);
xor U26679 (N_26679,N_26449,N_26323);
xor U26680 (N_26680,N_26362,N_26360);
and U26681 (N_26681,N_26155,N_26200);
xor U26682 (N_26682,N_26192,N_26305);
or U26683 (N_26683,N_26272,N_26483);
nor U26684 (N_26684,N_26383,N_26427);
nand U26685 (N_26685,N_26084,N_26207);
nand U26686 (N_26686,N_26024,N_26357);
nand U26687 (N_26687,N_26101,N_26064);
nor U26688 (N_26688,N_26194,N_26161);
xor U26689 (N_26689,N_26171,N_26118);
or U26690 (N_26690,N_26222,N_26499);
or U26691 (N_26691,N_26205,N_26354);
nand U26692 (N_26692,N_26014,N_26055);
and U26693 (N_26693,N_26042,N_26393);
xnor U26694 (N_26694,N_26158,N_26289);
and U26695 (N_26695,N_26180,N_26266);
or U26696 (N_26696,N_26070,N_26017);
xnor U26697 (N_26697,N_26300,N_26322);
and U26698 (N_26698,N_26482,N_26164);
or U26699 (N_26699,N_26117,N_26317);
or U26700 (N_26700,N_26065,N_26455);
nor U26701 (N_26701,N_26330,N_26114);
or U26702 (N_26702,N_26214,N_26473);
and U26703 (N_26703,N_26268,N_26387);
nand U26704 (N_26704,N_26417,N_26291);
or U26705 (N_26705,N_26261,N_26007);
and U26706 (N_26706,N_26497,N_26315);
and U26707 (N_26707,N_26496,N_26213);
and U26708 (N_26708,N_26191,N_26095);
nor U26709 (N_26709,N_26251,N_26351);
and U26710 (N_26710,N_26081,N_26335);
and U26711 (N_26711,N_26197,N_26037);
nand U26712 (N_26712,N_26463,N_26069);
xnor U26713 (N_26713,N_26094,N_26424);
nand U26714 (N_26714,N_26310,N_26407);
and U26715 (N_26715,N_26250,N_26346);
and U26716 (N_26716,N_26309,N_26340);
nor U26717 (N_26717,N_26032,N_26187);
or U26718 (N_26718,N_26302,N_26477);
and U26719 (N_26719,N_26379,N_26382);
nand U26720 (N_26720,N_26378,N_26277);
and U26721 (N_26721,N_26328,N_26071);
or U26722 (N_26722,N_26493,N_26478);
or U26723 (N_26723,N_26356,N_26026);
nor U26724 (N_26724,N_26452,N_26275);
nor U26725 (N_26725,N_26253,N_26129);
nand U26726 (N_26726,N_26442,N_26160);
or U26727 (N_26727,N_26004,N_26475);
nand U26728 (N_26728,N_26373,N_26304);
xnor U26729 (N_26729,N_26233,N_26168);
nand U26730 (N_26730,N_26403,N_26130);
nand U26731 (N_26731,N_26174,N_26228);
nand U26732 (N_26732,N_26414,N_26329);
nor U26733 (N_26733,N_26136,N_26092);
and U26734 (N_26734,N_26049,N_26193);
xor U26735 (N_26735,N_26051,N_26080);
xor U26736 (N_26736,N_26440,N_26015);
or U26737 (N_26737,N_26355,N_26466);
and U26738 (N_26738,N_26011,N_26416);
xor U26739 (N_26739,N_26280,N_26184);
and U26740 (N_26740,N_26175,N_26050);
nand U26741 (N_26741,N_26450,N_26143);
nor U26742 (N_26742,N_26366,N_26258);
nand U26743 (N_26743,N_26120,N_26126);
nand U26744 (N_26744,N_26044,N_26420);
nor U26745 (N_26745,N_26429,N_26491);
and U26746 (N_26746,N_26188,N_26283);
xnor U26747 (N_26747,N_26238,N_26179);
xor U26748 (N_26748,N_26162,N_26041);
or U26749 (N_26749,N_26020,N_26326);
nand U26750 (N_26750,N_26210,N_26309);
nor U26751 (N_26751,N_26368,N_26440);
nor U26752 (N_26752,N_26152,N_26347);
xor U26753 (N_26753,N_26371,N_26266);
xnor U26754 (N_26754,N_26469,N_26290);
and U26755 (N_26755,N_26367,N_26114);
or U26756 (N_26756,N_26149,N_26280);
nor U26757 (N_26757,N_26389,N_26449);
nand U26758 (N_26758,N_26318,N_26210);
xor U26759 (N_26759,N_26327,N_26286);
nand U26760 (N_26760,N_26363,N_26066);
xnor U26761 (N_26761,N_26013,N_26470);
nand U26762 (N_26762,N_26380,N_26238);
and U26763 (N_26763,N_26139,N_26113);
and U26764 (N_26764,N_26292,N_26472);
or U26765 (N_26765,N_26059,N_26109);
nand U26766 (N_26766,N_26253,N_26347);
nand U26767 (N_26767,N_26130,N_26171);
xnor U26768 (N_26768,N_26414,N_26092);
or U26769 (N_26769,N_26215,N_26378);
xor U26770 (N_26770,N_26257,N_26102);
xnor U26771 (N_26771,N_26109,N_26025);
nor U26772 (N_26772,N_26399,N_26330);
xnor U26773 (N_26773,N_26332,N_26129);
and U26774 (N_26774,N_26380,N_26151);
nand U26775 (N_26775,N_26468,N_26028);
nor U26776 (N_26776,N_26112,N_26331);
nand U26777 (N_26777,N_26391,N_26252);
xnor U26778 (N_26778,N_26150,N_26223);
xor U26779 (N_26779,N_26474,N_26102);
xor U26780 (N_26780,N_26086,N_26419);
and U26781 (N_26781,N_26374,N_26486);
and U26782 (N_26782,N_26334,N_26183);
xor U26783 (N_26783,N_26221,N_26394);
or U26784 (N_26784,N_26060,N_26446);
nor U26785 (N_26785,N_26368,N_26071);
nor U26786 (N_26786,N_26300,N_26067);
nand U26787 (N_26787,N_26468,N_26100);
xnor U26788 (N_26788,N_26330,N_26142);
nand U26789 (N_26789,N_26129,N_26437);
and U26790 (N_26790,N_26424,N_26180);
or U26791 (N_26791,N_26078,N_26354);
xnor U26792 (N_26792,N_26135,N_26266);
xor U26793 (N_26793,N_26219,N_26065);
xor U26794 (N_26794,N_26201,N_26164);
nand U26795 (N_26795,N_26020,N_26053);
nor U26796 (N_26796,N_26375,N_26201);
nor U26797 (N_26797,N_26451,N_26149);
nand U26798 (N_26798,N_26417,N_26352);
nand U26799 (N_26799,N_26350,N_26405);
and U26800 (N_26800,N_26462,N_26341);
xnor U26801 (N_26801,N_26354,N_26364);
nand U26802 (N_26802,N_26317,N_26052);
nor U26803 (N_26803,N_26169,N_26348);
nor U26804 (N_26804,N_26334,N_26425);
xnor U26805 (N_26805,N_26266,N_26198);
nor U26806 (N_26806,N_26394,N_26048);
nor U26807 (N_26807,N_26298,N_26442);
nand U26808 (N_26808,N_26435,N_26130);
and U26809 (N_26809,N_26269,N_26270);
nand U26810 (N_26810,N_26420,N_26356);
or U26811 (N_26811,N_26141,N_26484);
or U26812 (N_26812,N_26436,N_26005);
xor U26813 (N_26813,N_26204,N_26491);
nand U26814 (N_26814,N_26431,N_26385);
nand U26815 (N_26815,N_26257,N_26366);
xor U26816 (N_26816,N_26431,N_26241);
nor U26817 (N_26817,N_26305,N_26189);
nand U26818 (N_26818,N_26005,N_26496);
and U26819 (N_26819,N_26393,N_26022);
xnor U26820 (N_26820,N_26344,N_26120);
and U26821 (N_26821,N_26493,N_26081);
or U26822 (N_26822,N_26186,N_26226);
and U26823 (N_26823,N_26382,N_26130);
nand U26824 (N_26824,N_26188,N_26039);
and U26825 (N_26825,N_26213,N_26314);
xor U26826 (N_26826,N_26257,N_26445);
or U26827 (N_26827,N_26241,N_26415);
and U26828 (N_26828,N_26366,N_26347);
and U26829 (N_26829,N_26049,N_26489);
nor U26830 (N_26830,N_26088,N_26477);
nand U26831 (N_26831,N_26207,N_26267);
or U26832 (N_26832,N_26010,N_26263);
nand U26833 (N_26833,N_26483,N_26499);
nor U26834 (N_26834,N_26416,N_26160);
nand U26835 (N_26835,N_26410,N_26251);
or U26836 (N_26836,N_26084,N_26325);
and U26837 (N_26837,N_26138,N_26370);
and U26838 (N_26838,N_26124,N_26173);
nand U26839 (N_26839,N_26246,N_26191);
nand U26840 (N_26840,N_26129,N_26221);
or U26841 (N_26841,N_26446,N_26431);
nand U26842 (N_26842,N_26341,N_26314);
nor U26843 (N_26843,N_26464,N_26126);
nand U26844 (N_26844,N_26357,N_26420);
xor U26845 (N_26845,N_26405,N_26256);
and U26846 (N_26846,N_26356,N_26315);
and U26847 (N_26847,N_26105,N_26169);
or U26848 (N_26848,N_26288,N_26315);
or U26849 (N_26849,N_26044,N_26055);
nand U26850 (N_26850,N_26440,N_26496);
xnor U26851 (N_26851,N_26373,N_26092);
and U26852 (N_26852,N_26490,N_26291);
and U26853 (N_26853,N_26233,N_26325);
nand U26854 (N_26854,N_26237,N_26077);
or U26855 (N_26855,N_26093,N_26173);
or U26856 (N_26856,N_26179,N_26292);
nand U26857 (N_26857,N_26223,N_26060);
and U26858 (N_26858,N_26231,N_26375);
nor U26859 (N_26859,N_26338,N_26043);
xnor U26860 (N_26860,N_26359,N_26205);
nor U26861 (N_26861,N_26319,N_26405);
nand U26862 (N_26862,N_26295,N_26364);
or U26863 (N_26863,N_26310,N_26154);
xor U26864 (N_26864,N_26153,N_26088);
nor U26865 (N_26865,N_26485,N_26417);
xnor U26866 (N_26866,N_26305,N_26203);
and U26867 (N_26867,N_26353,N_26099);
nand U26868 (N_26868,N_26257,N_26295);
nor U26869 (N_26869,N_26465,N_26170);
xnor U26870 (N_26870,N_26435,N_26062);
or U26871 (N_26871,N_26314,N_26237);
nor U26872 (N_26872,N_26427,N_26238);
and U26873 (N_26873,N_26341,N_26161);
xnor U26874 (N_26874,N_26387,N_26342);
xor U26875 (N_26875,N_26190,N_26079);
nand U26876 (N_26876,N_26173,N_26435);
and U26877 (N_26877,N_26010,N_26446);
nor U26878 (N_26878,N_26412,N_26151);
nor U26879 (N_26879,N_26125,N_26091);
xnor U26880 (N_26880,N_26093,N_26265);
nor U26881 (N_26881,N_26315,N_26321);
nand U26882 (N_26882,N_26370,N_26461);
and U26883 (N_26883,N_26113,N_26479);
nand U26884 (N_26884,N_26412,N_26188);
or U26885 (N_26885,N_26265,N_26008);
or U26886 (N_26886,N_26284,N_26215);
or U26887 (N_26887,N_26312,N_26417);
nand U26888 (N_26888,N_26234,N_26035);
nand U26889 (N_26889,N_26497,N_26305);
xor U26890 (N_26890,N_26282,N_26208);
nor U26891 (N_26891,N_26070,N_26025);
nor U26892 (N_26892,N_26300,N_26039);
or U26893 (N_26893,N_26378,N_26465);
nor U26894 (N_26894,N_26057,N_26220);
nor U26895 (N_26895,N_26285,N_26408);
or U26896 (N_26896,N_26446,N_26356);
nand U26897 (N_26897,N_26272,N_26396);
nor U26898 (N_26898,N_26176,N_26295);
xor U26899 (N_26899,N_26130,N_26020);
or U26900 (N_26900,N_26149,N_26001);
nand U26901 (N_26901,N_26073,N_26383);
nor U26902 (N_26902,N_26108,N_26229);
and U26903 (N_26903,N_26076,N_26023);
and U26904 (N_26904,N_26284,N_26211);
or U26905 (N_26905,N_26212,N_26363);
or U26906 (N_26906,N_26077,N_26258);
xnor U26907 (N_26907,N_26313,N_26021);
nor U26908 (N_26908,N_26310,N_26101);
xor U26909 (N_26909,N_26176,N_26310);
nand U26910 (N_26910,N_26380,N_26318);
xor U26911 (N_26911,N_26265,N_26498);
or U26912 (N_26912,N_26152,N_26353);
or U26913 (N_26913,N_26297,N_26034);
xor U26914 (N_26914,N_26098,N_26428);
or U26915 (N_26915,N_26295,N_26307);
nor U26916 (N_26916,N_26407,N_26386);
and U26917 (N_26917,N_26109,N_26378);
nand U26918 (N_26918,N_26149,N_26299);
nor U26919 (N_26919,N_26093,N_26363);
and U26920 (N_26920,N_26245,N_26311);
nand U26921 (N_26921,N_26255,N_26020);
xor U26922 (N_26922,N_26400,N_26103);
nor U26923 (N_26923,N_26443,N_26284);
nand U26924 (N_26924,N_26105,N_26396);
nand U26925 (N_26925,N_26065,N_26348);
nand U26926 (N_26926,N_26124,N_26471);
nand U26927 (N_26927,N_26217,N_26147);
nor U26928 (N_26928,N_26367,N_26239);
and U26929 (N_26929,N_26385,N_26003);
and U26930 (N_26930,N_26253,N_26216);
nor U26931 (N_26931,N_26139,N_26401);
and U26932 (N_26932,N_26043,N_26316);
or U26933 (N_26933,N_26069,N_26318);
xnor U26934 (N_26934,N_26222,N_26064);
and U26935 (N_26935,N_26146,N_26102);
and U26936 (N_26936,N_26154,N_26467);
or U26937 (N_26937,N_26301,N_26365);
xor U26938 (N_26938,N_26366,N_26016);
xnor U26939 (N_26939,N_26161,N_26254);
nand U26940 (N_26940,N_26442,N_26495);
xor U26941 (N_26941,N_26199,N_26076);
nand U26942 (N_26942,N_26351,N_26113);
xnor U26943 (N_26943,N_26011,N_26142);
nand U26944 (N_26944,N_26415,N_26228);
or U26945 (N_26945,N_26050,N_26056);
nor U26946 (N_26946,N_26078,N_26170);
or U26947 (N_26947,N_26379,N_26361);
xor U26948 (N_26948,N_26144,N_26059);
xnor U26949 (N_26949,N_26000,N_26236);
xnor U26950 (N_26950,N_26398,N_26428);
nand U26951 (N_26951,N_26163,N_26387);
nor U26952 (N_26952,N_26358,N_26304);
or U26953 (N_26953,N_26497,N_26034);
or U26954 (N_26954,N_26438,N_26333);
and U26955 (N_26955,N_26206,N_26221);
and U26956 (N_26956,N_26467,N_26339);
nand U26957 (N_26957,N_26307,N_26347);
and U26958 (N_26958,N_26205,N_26209);
and U26959 (N_26959,N_26137,N_26220);
xor U26960 (N_26960,N_26332,N_26360);
nor U26961 (N_26961,N_26044,N_26415);
and U26962 (N_26962,N_26355,N_26459);
or U26963 (N_26963,N_26295,N_26254);
or U26964 (N_26964,N_26235,N_26211);
nor U26965 (N_26965,N_26094,N_26210);
xor U26966 (N_26966,N_26285,N_26384);
xnor U26967 (N_26967,N_26152,N_26418);
and U26968 (N_26968,N_26115,N_26113);
nor U26969 (N_26969,N_26484,N_26333);
nand U26970 (N_26970,N_26058,N_26003);
or U26971 (N_26971,N_26354,N_26118);
nor U26972 (N_26972,N_26256,N_26052);
and U26973 (N_26973,N_26325,N_26451);
nor U26974 (N_26974,N_26317,N_26478);
and U26975 (N_26975,N_26129,N_26291);
and U26976 (N_26976,N_26468,N_26417);
nor U26977 (N_26977,N_26308,N_26361);
or U26978 (N_26978,N_26437,N_26443);
nand U26979 (N_26979,N_26375,N_26075);
and U26980 (N_26980,N_26354,N_26088);
or U26981 (N_26981,N_26124,N_26118);
and U26982 (N_26982,N_26494,N_26273);
and U26983 (N_26983,N_26326,N_26319);
nand U26984 (N_26984,N_26275,N_26279);
xor U26985 (N_26985,N_26317,N_26432);
xor U26986 (N_26986,N_26297,N_26091);
or U26987 (N_26987,N_26065,N_26385);
nand U26988 (N_26988,N_26302,N_26186);
xor U26989 (N_26989,N_26261,N_26054);
xnor U26990 (N_26990,N_26304,N_26414);
and U26991 (N_26991,N_26142,N_26313);
xor U26992 (N_26992,N_26049,N_26097);
nor U26993 (N_26993,N_26360,N_26480);
nor U26994 (N_26994,N_26058,N_26091);
or U26995 (N_26995,N_26266,N_26391);
nand U26996 (N_26996,N_26452,N_26071);
nand U26997 (N_26997,N_26445,N_26277);
nand U26998 (N_26998,N_26074,N_26300);
and U26999 (N_26999,N_26003,N_26325);
or U27000 (N_27000,N_26917,N_26846);
nor U27001 (N_27001,N_26632,N_26804);
nand U27002 (N_27002,N_26955,N_26687);
nand U27003 (N_27003,N_26834,N_26784);
xnor U27004 (N_27004,N_26583,N_26680);
xor U27005 (N_27005,N_26947,N_26787);
xnor U27006 (N_27006,N_26880,N_26878);
or U27007 (N_27007,N_26888,N_26507);
nand U27008 (N_27008,N_26832,N_26890);
nand U27009 (N_27009,N_26624,N_26509);
xor U27010 (N_27010,N_26988,N_26653);
or U27011 (N_27011,N_26677,N_26548);
nor U27012 (N_27012,N_26761,N_26622);
nand U27013 (N_27013,N_26968,N_26926);
nor U27014 (N_27014,N_26969,N_26716);
nand U27015 (N_27015,N_26844,N_26875);
and U27016 (N_27016,N_26663,N_26522);
or U27017 (N_27017,N_26534,N_26764);
nand U27018 (N_27018,N_26995,N_26599);
xnor U27019 (N_27019,N_26619,N_26807);
nor U27020 (N_27020,N_26780,N_26750);
nand U27021 (N_27021,N_26506,N_26701);
nor U27022 (N_27022,N_26838,N_26965);
and U27023 (N_27023,N_26946,N_26667);
xnor U27024 (N_27024,N_26772,N_26665);
xnor U27025 (N_27025,N_26713,N_26837);
nor U27026 (N_27026,N_26670,N_26578);
or U27027 (N_27027,N_26868,N_26738);
and U27028 (N_27028,N_26524,N_26511);
xor U27029 (N_27029,N_26852,N_26860);
nor U27030 (N_27030,N_26876,N_26948);
or U27031 (N_27031,N_26513,N_26829);
nor U27032 (N_27032,N_26885,N_26603);
or U27033 (N_27033,N_26849,N_26676);
xor U27034 (N_27034,N_26997,N_26944);
nand U27035 (N_27035,N_26671,N_26637);
nor U27036 (N_27036,N_26959,N_26538);
nor U27037 (N_27037,N_26625,N_26694);
nor U27038 (N_27038,N_26999,N_26605);
nand U27039 (N_27039,N_26554,N_26618);
xor U27040 (N_27040,N_26977,N_26674);
or U27041 (N_27041,N_26759,N_26553);
nand U27042 (N_27042,N_26539,N_26596);
or U27043 (N_27043,N_26567,N_26669);
or U27044 (N_27044,N_26725,N_26769);
nor U27045 (N_27045,N_26881,N_26898);
nand U27046 (N_27046,N_26573,N_26691);
and U27047 (N_27047,N_26664,N_26980);
xnor U27048 (N_27048,N_26529,N_26666);
and U27049 (N_27049,N_26523,N_26963);
or U27050 (N_27050,N_26610,N_26773);
or U27051 (N_27051,N_26961,N_26717);
nand U27052 (N_27052,N_26648,N_26517);
or U27053 (N_27053,N_26574,N_26763);
xnor U27054 (N_27054,N_26699,N_26851);
and U27055 (N_27055,N_26649,N_26512);
and U27056 (N_27056,N_26783,N_26540);
xnor U27057 (N_27057,N_26941,N_26715);
nand U27058 (N_27058,N_26850,N_26927);
xnor U27059 (N_27059,N_26558,N_26874);
xor U27060 (N_27060,N_26733,N_26601);
or U27061 (N_27061,N_26910,N_26801);
nor U27062 (N_27062,N_26695,N_26752);
nor U27063 (N_27063,N_26613,N_26532);
nor U27064 (N_27064,N_26939,N_26704);
and U27065 (N_27065,N_26647,N_26744);
nor U27066 (N_27066,N_26604,N_26545);
nor U27067 (N_27067,N_26854,N_26818);
and U27068 (N_27068,N_26938,N_26710);
nor U27069 (N_27069,N_26933,N_26847);
nand U27070 (N_27070,N_26551,N_26835);
xnor U27071 (N_27071,N_26857,N_26819);
nor U27072 (N_27072,N_26561,N_26889);
nand U27073 (N_27073,N_26935,N_26983);
nor U27074 (N_27074,N_26905,N_26828);
and U27075 (N_27075,N_26655,N_26643);
xor U27076 (N_27076,N_26810,N_26564);
nor U27077 (N_27077,N_26753,N_26645);
and U27078 (N_27078,N_26748,N_26651);
xor U27079 (N_27079,N_26608,N_26500);
nand U27080 (N_27080,N_26901,N_26537);
xor U27081 (N_27081,N_26893,N_26747);
xnor U27082 (N_27082,N_26799,N_26689);
and U27083 (N_27083,N_26631,N_26639);
xnor U27084 (N_27084,N_26952,N_26930);
xnor U27085 (N_27085,N_26644,N_26634);
and U27086 (N_27086,N_26510,N_26755);
or U27087 (N_27087,N_26683,N_26919);
or U27088 (N_27088,N_26629,N_26731);
and U27089 (N_27089,N_26745,N_26505);
xnor U27090 (N_27090,N_26813,N_26668);
nand U27091 (N_27091,N_26929,N_26895);
nor U27092 (N_27092,N_26957,N_26730);
nand U27093 (N_27093,N_26897,N_26812);
nor U27094 (N_27094,N_26887,N_26547);
nand U27095 (N_27095,N_26729,N_26953);
and U27096 (N_27096,N_26584,N_26791);
xor U27097 (N_27097,N_26535,N_26697);
or U27098 (N_27098,N_26816,N_26956);
and U27099 (N_27099,N_26964,N_26842);
or U27100 (N_27100,N_26682,N_26552);
nor U27101 (N_27101,N_26581,N_26519);
xnor U27102 (N_27102,N_26742,N_26657);
xor U27103 (N_27103,N_26760,N_26521);
and U27104 (N_27104,N_26877,N_26626);
nor U27105 (N_27105,N_26661,N_26912);
nor U27106 (N_27106,N_26830,N_26652);
or U27107 (N_27107,N_26972,N_26673);
nand U27108 (N_27108,N_26616,N_26913);
and U27109 (N_27109,N_26908,N_26514);
or U27110 (N_27110,N_26734,N_26709);
nand U27111 (N_27111,N_26768,N_26594);
nor U27112 (N_27112,N_26916,N_26520);
nor U27113 (N_27113,N_26530,N_26967);
nor U27114 (N_27114,N_26706,N_26976);
xnor U27115 (N_27115,N_26981,N_26803);
nand U27116 (N_27116,N_26627,N_26598);
and U27117 (N_27117,N_26911,N_26903);
xnor U27118 (N_27118,N_26580,N_26686);
nor U27119 (N_27119,N_26526,N_26990);
xnor U27120 (N_27120,N_26942,N_26970);
and U27121 (N_27121,N_26568,N_26525);
nor U27122 (N_27122,N_26951,N_26588);
nor U27123 (N_27123,N_26931,N_26754);
or U27124 (N_27124,N_26718,N_26623);
and U27125 (N_27125,N_26815,N_26638);
or U27126 (N_27126,N_26576,N_26600);
xnor U27127 (N_27127,N_26612,N_26794);
nand U27128 (N_27128,N_26650,N_26918);
nand U27129 (N_27129,N_26743,N_26735);
xnor U27130 (N_27130,N_26550,N_26575);
xnor U27131 (N_27131,N_26693,N_26985);
nor U27132 (N_27132,N_26593,N_26757);
nand U27133 (N_27133,N_26630,N_26590);
nand U27134 (N_27134,N_26636,N_26698);
nand U27135 (N_27135,N_26726,N_26820);
and U27136 (N_27136,N_26770,N_26891);
nand U27137 (N_27137,N_26937,N_26789);
or U27138 (N_27138,N_26560,N_26659);
xor U27139 (N_27139,N_26595,N_26678);
nor U27140 (N_27140,N_26936,N_26658);
xnor U27141 (N_27141,N_26831,N_26504);
nor U27142 (N_27142,N_26607,N_26719);
nor U27143 (N_27143,N_26765,N_26790);
xnor U27144 (N_27144,N_26703,N_26615);
and U27145 (N_27145,N_26776,N_26902);
nand U27146 (N_27146,N_26805,N_26728);
or U27147 (N_27147,N_26797,N_26681);
or U27148 (N_27148,N_26899,N_26871);
xnor U27149 (N_27149,N_26886,N_26592);
nand U27150 (N_27150,N_26853,N_26924);
nand U27151 (N_27151,N_26823,N_26502);
or U27152 (N_27152,N_26579,N_26563);
xor U27153 (N_27153,N_26907,N_26503);
nand U27154 (N_27154,N_26587,N_26758);
nand U27155 (N_27155,N_26727,N_26786);
nand U27156 (N_27156,N_26869,N_26991);
or U27157 (N_27157,N_26708,N_26646);
or U27158 (N_27158,N_26922,N_26771);
nand U27159 (N_27159,N_26700,N_26998);
or U27160 (N_27160,N_26751,N_26739);
xnor U27161 (N_27161,N_26696,N_26900);
nor U27162 (N_27162,N_26611,N_26873);
nand U27163 (N_27163,N_26746,N_26516);
xnor U27164 (N_27164,N_26614,N_26940);
nand U27165 (N_27165,N_26542,N_26923);
and U27166 (N_27166,N_26654,N_26884);
or U27167 (N_27167,N_26802,N_26814);
or U27168 (N_27168,N_26641,N_26577);
and U27169 (N_27169,N_26870,N_26855);
nand U27170 (N_27170,N_26762,N_26732);
nand U27171 (N_27171,N_26609,N_26992);
and U27172 (N_27172,N_26856,N_26766);
nand U27173 (N_27173,N_26925,N_26958);
or U27174 (N_27174,N_26996,N_26945);
or U27175 (N_27175,N_26793,N_26571);
or U27176 (N_27176,N_26914,N_26872);
nand U27177 (N_27177,N_26882,N_26781);
xor U27178 (N_27178,N_26839,N_26987);
nor U27179 (N_27179,N_26672,N_26824);
or U27180 (N_27180,N_26896,N_26777);
nor U27181 (N_27181,N_26966,N_26556);
or U27182 (N_27182,N_26909,N_26740);
nor U27183 (N_27183,N_26642,N_26620);
xor U27184 (N_27184,N_26861,N_26690);
and U27185 (N_27185,N_26827,N_26817);
or U27186 (N_27186,N_26741,N_26994);
and U27187 (N_27187,N_26749,N_26943);
or U27188 (N_27188,N_26640,N_26660);
nor U27189 (N_27189,N_26633,N_26591);
nand U27190 (N_27190,N_26932,N_26723);
and U27191 (N_27191,N_26707,N_26606);
xnor U27192 (N_27192,N_26821,N_26788);
nor U27193 (N_27193,N_26974,N_26779);
or U27194 (N_27194,N_26962,N_26825);
xnor U27195 (N_27195,N_26792,N_26688);
and U27196 (N_27196,N_26836,N_26978);
or U27197 (N_27197,N_26971,N_26892);
or U27198 (N_27198,N_26702,N_26859);
xor U27199 (N_27199,N_26508,N_26714);
and U27200 (N_27200,N_26841,N_26555);
or U27201 (N_27201,N_26774,N_26546);
or U27202 (N_27202,N_26883,N_26848);
nand U27203 (N_27203,N_26954,N_26617);
or U27204 (N_27204,N_26767,N_26920);
or U27205 (N_27205,N_26712,N_26662);
xnor U27206 (N_27206,N_26982,N_26565);
and U27207 (N_27207,N_26656,N_26721);
or U27208 (N_27208,N_26737,N_26635);
and U27209 (N_27209,N_26973,N_26566);
nand U27210 (N_27210,N_26559,N_26543);
xor U27211 (N_27211,N_26879,N_26934);
nor U27212 (N_27212,N_26904,N_26549);
xor U27213 (N_27213,N_26527,N_26711);
nor U27214 (N_27214,N_26845,N_26684);
or U27215 (N_27215,N_26736,N_26775);
xnor U27216 (N_27216,N_26984,N_26628);
xnor U27217 (N_27217,N_26515,N_26858);
xnor U27218 (N_27218,N_26685,N_26867);
nand U27219 (N_27219,N_26811,N_26724);
nand U27220 (N_27220,N_26795,N_26975);
and U27221 (N_27221,N_26586,N_26570);
and U27222 (N_27222,N_26585,N_26501);
xnor U27223 (N_27223,N_26602,N_26778);
nand U27224 (N_27224,N_26921,N_26562);
and U27225 (N_27225,N_26979,N_26785);
or U27226 (N_27226,N_26798,N_26536);
nor U27227 (N_27227,N_26533,N_26986);
and U27228 (N_27228,N_26906,N_26569);
nand U27229 (N_27229,N_26756,N_26949);
or U27230 (N_27230,N_26528,N_26621);
or U27231 (N_27231,N_26993,N_26822);
and U27232 (N_27232,N_26862,N_26809);
nand U27233 (N_27233,N_26541,N_26894);
xor U27234 (N_27234,N_26531,N_26866);
xor U27235 (N_27235,N_26865,N_26826);
nor U27236 (N_27236,N_26597,N_26915);
or U27237 (N_27237,N_26782,N_26960);
nand U27238 (N_27238,N_26557,N_26806);
or U27239 (N_27239,N_26928,N_26840);
xor U27240 (N_27240,N_26833,N_26863);
and U27241 (N_27241,N_26796,N_26864);
nor U27242 (N_27242,N_26989,N_26582);
or U27243 (N_27243,N_26572,N_26705);
nand U27244 (N_27244,N_26675,N_26950);
or U27245 (N_27245,N_26720,N_26679);
nor U27246 (N_27246,N_26843,N_26544);
nand U27247 (N_27247,N_26722,N_26800);
nand U27248 (N_27248,N_26692,N_26808);
and U27249 (N_27249,N_26518,N_26589);
nand U27250 (N_27250,N_26616,N_26523);
xnor U27251 (N_27251,N_26688,N_26796);
or U27252 (N_27252,N_26586,N_26514);
xnor U27253 (N_27253,N_26712,N_26575);
xor U27254 (N_27254,N_26924,N_26506);
or U27255 (N_27255,N_26687,N_26690);
or U27256 (N_27256,N_26947,N_26503);
nor U27257 (N_27257,N_26537,N_26610);
xnor U27258 (N_27258,N_26633,N_26637);
nor U27259 (N_27259,N_26868,N_26991);
or U27260 (N_27260,N_26577,N_26562);
or U27261 (N_27261,N_26767,N_26898);
or U27262 (N_27262,N_26523,N_26993);
or U27263 (N_27263,N_26578,N_26979);
xnor U27264 (N_27264,N_26878,N_26709);
or U27265 (N_27265,N_26714,N_26581);
and U27266 (N_27266,N_26674,N_26777);
and U27267 (N_27267,N_26980,N_26880);
or U27268 (N_27268,N_26805,N_26770);
nand U27269 (N_27269,N_26950,N_26705);
xor U27270 (N_27270,N_26944,N_26677);
nand U27271 (N_27271,N_26652,N_26912);
and U27272 (N_27272,N_26856,N_26677);
xnor U27273 (N_27273,N_26639,N_26509);
nor U27274 (N_27274,N_26990,N_26780);
xnor U27275 (N_27275,N_26535,N_26827);
or U27276 (N_27276,N_26915,N_26689);
or U27277 (N_27277,N_26994,N_26926);
xor U27278 (N_27278,N_26684,N_26686);
nand U27279 (N_27279,N_26964,N_26657);
nand U27280 (N_27280,N_26514,N_26779);
or U27281 (N_27281,N_26875,N_26578);
or U27282 (N_27282,N_26670,N_26524);
and U27283 (N_27283,N_26707,N_26888);
xor U27284 (N_27284,N_26644,N_26622);
nor U27285 (N_27285,N_26953,N_26835);
xnor U27286 (N_27286,N_26902,N_26966);
nor U27287 (N_27287,N_26658,N_26924);
nor U27288 (N_27288,N_26642,N_26638);
or U27289 (N_27289,N_26792,N_26933);
xor U27290 (N_27290,N_26773,N_26961);
xnor U27291 (N_27291,N_26645,N_26902);
and U27292 (N_27292,N_26506,N_26903);
xnor U27293 (N_27293,N_26691,N_26603);
and U27294 (N_27294,N_26557,N_26911);
or U27295 (N_27295,N_26708,N_26559);
or U27296 (N_27296,N_26520,N_26899);
or U27297 (N_27297,N_26808,N_26560);
nor U27298 (N_27298,N_26791,N_26868);
or U27299 (N_27299,N_26641,N_26875);
and U27300 (N_27300,N_26569,N_26929);
or U27301 (N_27301,N_26536,N_26772);
xor U27302 (N_27302,N_26551,N_26887);
or U27303 (N_27303,N_26997,N_26524);
and U27304 (N_27304,N_26650,N_26723);
or U27305 (N_27305,N_26648,N_26980);
nor U27306 (N_27306,N_26549,N_26915);
or U27307 (N_27307,N_26883,N_26755);
nand U27308 (N_27308,N_26907,N_26855);
nor U27309 (N_27309,N_26752,N_26589);
or U27310 (N_27310,N_26551,N_26742);
and U27311 (N_27311,N_26871,N_26692);
nor U27312 (N_27312,N_26785,N_26719);
xor U27313 (N_27313,N_26955,N_26514);
and U27314 (N_27314,N_26797,N_26996);
or U27315 (N_27315,N_26742,N_26542);
or U27316 (N_27316,N_26975,N_26923);
and U27317 (N_27317,N_26714,N_26778);
nor U27318 (N_27318,N_26895,N_26874);
or U27319 (N_27319,N_26890,N_26792);
xor U27320 (N_27320,N_26749,N_26616);
xor U27321 (N_27321,N_26662,N_26938);
nor U27322 (N_27322,N_26657,N_26641);
or U27323 (N_27323,N_26777,N_26890);
and U27324 (N_27324,N_26563,N_26532);
nand U27325 (N_27325,N_26573,N_26527);
or U27326 (N_27326,N_26873,N_26565);
and U27327 (N_27327,N_26579,N_26735);
and U27328 (N_27328,N_26695,N_26943);
and U27329 (N_27329,N_26695,N_26817);
and U27330 (N_27330,N_26847,N_26820);
nand U27331 (N_27331,N_26660,N_26561);
or U27332 (N_27332,N_26632,N_26723);
nand U27333 (N_27333,N_26615,N_26972);
xnor U27334 (N_27334,N_26574,N_26871);
xor U27335 (N_27335,N_26911,N_26829);
xnor U27336 (N_27336,N_26558,N_26827);
or U27337 (N_27337,N_26802,N_26933);
nand U27338 (N_27338,N_26900,N_26753);
xor U27339 (N_27339,N_26808,N_26704);
xnor U27340 (N_27340,N_26656,N_26901);
nand U27341 (N_27341,N_26777,N_26863);
nand U27342 (N_27342,N_26574,N_26696);
nor U27343 (N_27343,N_26953,N_26736);
xor U27344 (N_27344,N_26955,N_26861);
nand U27345 (N_27345,N_26803,N_26520);
xor U27346 (N_27346,N_26714,N_26889);
or U27347 (N_27347,N_26765,N_26953);
and U27348 (N_27348,N_26902,N_26561);
and U27349 (N_27349,N_26598,N_26876);
xnor U27350 (N_27350,N_26730,N_26937);
nand U27351 (N_27351,N_26900,N_26657);
xnor U27352 (N_27352,N_26740,N_26823);
nand U27353 (N_27353,N_26948,N_26960);
nand U27354 (N_27354,N_26743,N_26894);
and U27355 (N_27355,N_26679,N_26848);
and U27356 (N_27356,N_26769,N_26514);
or U27357 (N_27357,N_26636,N_26943);
xor U27358 (N_27358,N_26597,N_26993);
nand U27359 (N_27359,N_26507,N_26790);
nor U27360 (N_27360,N_26779,N_26722);
xnor U27361 (N_27361,N_26560,N_26817);
xor U27362 (N_27362,N_26559,N_26972);
xnor U27363 (N_27363,N_26931,N_26651);
or U27364 (N_27364,N_26887,N_26778);
nor U27365 (N_27365,N_26771,N_26505);
or U27366 (N_27366,N_26576,N_26964);
nor U27367 (N_27367,N_26660,N_26874);
xnor U27368 (N_27368,N_26721,N_26650);
or U27369 (N_27369,N_26588,N_26675);
nand U27370 (N_27370,N_26854,N_26911);
or U27371 (N_27371,N_26833,N_26763);
xor U27372 (N_27372,N_26798,N_26838);
xor U27373 (N_27373,N_26746,N_26540);
and U27374 (N_27374,N_26638,N_26996);
xnor U27375 (N_27375,N_26922,N_26574);
xnor U27376 (N_27376,N_26631,N_26546);
or U27377 (N_27377,N_26690,N_26998);
or U27378 (N_27378,N_26516,N_26602);
nor U27379 (N_27379,N_26959,N_26996);
nand U27380 (N_27380,N_26572,N_26802);
or U27381 (N_27381,N_26983,N_26908);
nor U27382 (N_27382,N_26552,N_26764);
xnor U27383 (N_27383,N_26551,N_26899);
and U27384 (N_27384,N_26907,N_26857);
xor U27385 (N_27385,N_26799,N_26777);
or U27386 (N_27386,N_26936,N_26696);
nand U27387 (N_27387,N_26918,N_26670);
nor U27388 (N_27388,N_26638,N_26511);
nand U27389 (N_27389,N_26912,N_26529);
nand U27390 (N_27390,N_26662,N_26647);
nor U27391 (N_27391,N_26749,N_26735);
xor U27392 (N_27392,N_26688,N_26929);
xor U27393 (N_27393,N_26865,N_26994);
nand U27394 (N_27394,N_26673,N_26551);
nand U27395 (N_27395,N_26958,N_26960);
and U27396 (N_27396,N_26945,N_26894);
nand U27397 (N_27397,N_26748,N_26861);
and U27398 (N_27398,N_26607,N_26653);
xor U27399 (N_27399,N_26726,N_26502);
nor U27400 (N_27400,N_26789,N_26979);
or U27401 (N_27401,N_26985,N_26794);
or U27402 (N_27402,N_26629,N_26515);
xnor U27403 (N_27403,N_26950,N_26930);
or U27404 (N_27404,N_26832,N_26502);
nor U27405 (N_27405,N_26749,N_26561);
or U27406 (N_27406,N_26517,N_26961);
or U27407 (N_27407,N_26886,N_26507);
and U27408 (N_27408,N_26946,N_26595);
xnor U27409 (N_27409,N_26955,N_26822);
xnor U27410 (N_27410,N_26770,N_26762);
nand U27411 (N_27411,N_26868,N_26528);
and U27412 (N_27412,N_26773,N_26607);
nor U27413 (N_27413,N_26822,N_26626);
nor U27414 (N_27414,N_26992,N_26513);
or U27415 (N_27415,N_26685,N_26625);
nor U27416 (N_27416,N_26914,N_26689);
nor U27417 (N_27417,N_26654,N_26863);
and U27418 (N_27418,N_26840,N_26843);
or U27419 (N_27419,N_26943,N_26628);
and U27420 (N_27420,N_26895,N_26736);
and U27421 (N_27421,N_26803,N_26894);
xor U27422 (N_27422,N_26797,N_26641);
xor U27423 (N_27423,N_26942,N_26781);
or U27424 (N_27424,N_26763,N_26979);
and U27425 (N_27425,N_26703,N_26900);
nand U27426 (N_27426,N_26609,N_26698);
xnor U27427 (N_27427,N_26596,N_26777);
nand U27428 (N_27428,N_26887,N_26671);
and U27429 (N_27429,N_26746,N_26869);
nor U27430 (N_27430,N_26811,N_26550);
nor U27431 (N_27431,N_26728,N_26615);
xor U27432 (N_27432,N_26668,N_26539);
nand U27433 (N_27433,N_26643,N_26853);
nand U27434 (N_27434,N_26607,N_26547);
nand U27435 (N_27435,N_26821,N_26503);
or U27436 (N_27436,N_26876,N_26968);
and U27437 (N_27437,N_26738,N_26762);
or U27438 (N_27438,N_26707,N_26848);
xnor U27439 (N_27439,N_26896,N_26722);
xnor U27440 (N_27440,N_26964,N_26751);
xnor U27441 (N_27441,N_26671,N_26749);
or U27442 (N_27442,N_26746,N_26742);
or U27443 (N_27443,N_26848,N_26666);
nor U27444 (N_27444,N_26602,N_26768);
nor U27445 (N_27445,N_26507,N_26725);
xnor U27446 (N_27446,N_26828,N_26582);
and U27447 (N_27447,N_26521,N_26517);
xnor U27448 (N_27448,N_26558,N_26941);
xor U27449 (N_27449,N_26780,N_26733);
nor U27450 (N_27450,N_26652,N_26948);
nor U27451 (N_27451,N_26711,N_26912);
nor U27452 (N_27452,N_26672,N_26543);
and U27453 (N_27453,N_26700,N_26663);
and U27454 (N_27454,N_26981,N_26919);
xor U27455 (N_27455,N_26757,N_26564);
xor U27456 (N_27456,N_26813,N_26568);
or U27457 (N_27457,N_26800,N_26785);
and U27458 (N_27458,N_26748,N_26868);
nor U27459 (N_27459,N_26842,N_26617);
xnor U27460 (N_27460,N_26807,N_26723);
or U27461 (N_27461,N_26999,N_26642);
xnor U27462 (N_27462,N_26559,N_26941);
and U27463 (N_27463,N_26547,N_26671);
nand U27464 (N_27464,N_26767,N_26607);
nor U27465 (N_27465,N_26961,N_26932);
nand U27466 (N_27466,N_26968,N_26639);
nand U27467 (N_27467,N_26857,N_26995);
nor U27468 (N_27468,N_26883,N_26567);
xnor U27469 (N_27469,N_26921,N_26593);
nand U27470 (N_27470,N_26753,N_26608);
or U27471 (N_27471,N_26508,N_26733);
and U27472 (N_27472,N_26943,N_26955);
nand U27473 (N_27473,N_26576,N_26865);
nor U27474 (N_27474,N_26727,N_26993);
xnor U27475 (N_27475,N_26810,N_26848);
nand U27476 (N_27476,N_26857,N_26713);
or U27477 (N_27477,N_26873,N_26880);
nor U27478 (N_27478,N_26960,N_26649);
nor U27479 (N_27479,N_26718,N_26540);
nand U27480 (N_27480,N_26911,N_26614);
xor U27481 (N_27481,N_26764,N_26775);
and U27482 (N_27482,N_26901,N_26932);
nor U27483 (N_27483,N_26648,N_26646);
and U27484 (N_27484,N_26570,N_26807);
nor U27485 (N_27485,N_26637,N_26623);
nor U27486 (N_27486,N_26876,N_26702);
xnor U27487 (N_27487,N_26593,N_26554);
xnor U27488 (N_27488,N_26657,N_26834);
and U27489 (N_27489,N_26977,N_26806);
nand U27490 (N_27490,N_26564,N_26997);
xnor U27491 (N_27491,N_26858,N_26855);
nor U27492 (N_27492,N_26725,N_26621);
nor U27493 (N_27493,N_26839,N_26572);
nor U27494 (N_27494,N_26832,N_26948);
xor U27495 (N_27495,N_26695,N_26709);
and U27496 (N_27496,N_26897,N_26932);
nand U27497 (N_27497,N_26554,N_26749);
or U27498 (N_27498,N_26982,N_26509);
nand U27499 (N_27499,N_26912,N_26640);
xnor U27500 (N_27500,N_27084,N_27444);
nand U27501 (N_27501,N_27223,N_27023);
xnor U27502 (N_27502,N_27251,N_27157);
and U27503 (N_27503,N_27463,N_27384);
and U27504 (N_27504,N_27191,N_27380);
and U27505 (N_27505,N_27300,N_27335);
nor U27506 (N_27506,N_27214,N_27271);
nor U27507 (N_27507,N_27320,N_27123);
xor U27508 (N_27508,N_27201,N_27165);
nor U27509 (N_27509,N_27051,N_27158);
xnor U27510 (N_27510,N_27287,N_27153);
nor U27511 (N_27511,N_27053,N_27456);
nor U27512 (N_27512,N_27237,N_27050);
and U27513 (N_27513,N_27003,N_27283);
and U27514 (N_27514,N_27495,N_27074);
or U27515 (N_27515,N_27253,N_27422);
nor U27516 (N_27516,N_27092,N_27397);
and U27517 (N_27517,N_27485,N_27008);
nor U27518 (N_27518,N_27361,N_27220);
nand U27519 (N_27519,N_27405,N_27021);
nor U27520 (N_27520,N_27216,N_27160);
or U27521 (N_27521,N_27224,N_27094);
and U27522 (N_27522,N_27186,N_27403);
nor U27523 (N_27523,N_27130,N_27069);
and U27524 (N_27524,N_27337,N_27033);
and U27525 (N_27525,N_27349,N_27414);
or U27526 (N_27526,N_27228,N_27198);
or U27527 (N_27527,N_27119,N_27254);
xnor U27528 (N_27528,N_27188,N_27034);
and U27529 (N_27529,N_27281,N_27098);
nand U27530 (N_27530,N_27371,N_27260);
xnor U27531 (N_27531,N_27404,N_27221);
nor U27532 (N_27532,N_27163,N_27316);
xor U27533 (N_27533,N_27341,N_27313);
xor U27534 (N_27534,N_27409,N_27238);
xnor U27535 (N_27535,N_27464,N_27484);
or U27536 (N_27536,N_27174,N_27440);
nand U27537 (N_27537,N_27326,N_27429);
xnor U27538 (N_27538,N_27467,N_27132);
and U27539 (N_27539,N_27309,N_27466);
nand U27540 (N_27540,N_27280,N_27151);
nor U27541 (N_27541,N_27450,N_27204);
and U27542 (N_27542,N_27202,N_27244);
or U27543 (N_27543,N_27210,N_27138);
nand U27544 (N_27544,N_27412,N_27282);
and U27545 (N_27545,N_27424,N_27056);
or U27546 (N_27546,N_27116,N_27275);
nor U27547 (N_27547,N_27012,N_27332);
nor U27548 (N_27548,N_27024,N_27054);
nor U27549 (N_27549,N_27036,N_27219);
nand U27550 (N_27550,N_27112,N_27308);
xnor U27551 (N_27551,N_27070,N_27458);
and U27552 (N_27552,N_27019,N_27108);
nand U27553 (N_27553,N_27342,N_27179);
or U27554 (N_27554,N_27298,N_27078);
xor U27555 (N_27555,N_27048,N_27047);
and U27556 (N_27556,N_27460,N_27277);
nand U27557 (N_27557,N_27149,N_27076);
nand U27558 (N_27558,N_27322,N_27031);
nor U27559 (N_27559,N_27290,N_27192);
nand U27560 (N_27560,N_27242,N_27391);
nand U27561 (N_27561,N_27431,N_27468);
nand U27562 (N_27562,N_27473,N_27383);
or U27563 (N_27563,N_27410,N_27453);
or U27564 (N_27564,N_27226,N_27386);
or U27565 (N_27565,N_27490,N_27339);
nor U27566 (N_27566,N_27315,N_27285);
nor U27567 (N_27567,N_27373,N_27388);
nor U27568 (N_27568,N_27434,N_27292);
nand U27569 (N_27569,N_27338,N_27103);
and U27570 (N_27570,N_27025,N_27016);
xor U27571 (N_27571,N_27068,N_27161);
nor U27572 (N_27572,N_27369,N_27117);
or U27573 (N_27573,N_27213,N_27312);
xnor U27574 (N_27574,N_27058,N_27252);
nand U27575 (N_27575,N_27156,N_27235);
nand U27576 (N_27576,N_27042,N_27476);
nand U27577 (N_27577,N_27284,N_27364);
nor U27578 (N_27578,N_27278,N_27107);
or U27579 (N_27579,N_27407,N_27289);
nand U27580 (N_27580,N_27459,N_27328);
xor U27581 (N_27581,N_27043,N_27073);
or U27582 (N_27582,N_27137,N_27408);
nand U27583 (N_27583,N_27478,N_27131);
nor U27584 (N_27584,N_27110,N_27480);
xnor U27585 (N_27585,N_27488,N_27441);
nand U27586 (N_27586,N_27091,N_27493);
and U27587 (N_27587,N_27304,N_27154);
or U27588 (N_27588,N_27199,N_27010);
and U27589 (N_27589,N_27415,N_27295);
or U27590 (N_27590,N_27211,N_27365);
and U27591 (N_27591,N_27439,N_27225);
and U27592 (N_27592,N_27115,N_27075);
and U27593 (N_27593,N_27269,N_27207);
nor U27594 (N_27594,N_27302,N_27279);
or U27595 (N_27595,N_27370,N_27085);
and U27596 (N_27596,N_27089,N_27120);
or U27597 (N_27597,N_27258,N_27381);
xor U27598 (N_27598,N_27374,N_27134);
or U27599 (N_27599,N_27100,N_27001);
xor U27600 (N_27600,N_27105,N_27129);
nand U27601 (N_27601,N_27396,N_27368);
or U27602 (N_27602,N_27472,N_27474);
xnor U27603 (N_27603,N_27022,N_27497);
or U27604 (N_27604,N_27417,N_27243);
xor U27605 (N_27605,N_27353,N_27145);
and U27606 (N_27606,N_27081,N_27272);
nand U27607 (N_27607,N_27425,N_27419);
and U27608 (N_27608,N_27239,N_27035);
nand U27609 (N_27609,N_27475,N_27299);
nor U27610 (N_27610,N_27358,N_27379);
nand U27611 (N_27611,N_27447,N_27345);
nand U27612 (N_27612,N_27392,N_27166);
xor U27613 (N_27613,N_27127,N_27294);
nor U27614 (N_27614,N_27395,N_27125);
and U27615 (N_27615,N_27433,N_27026);
or U27616 (N_27616,N_27133,N_27323);
nor U27617 (N_27617,N_27028,N_27066);
xor U27618 (N_27618,N_27234,N_27347);
or U27619 (N_27619,N_27448,N_27005);
or U27620 (N_27620,N_27064,N_27082);
and U27621 (N_27621,N_27274,N_27147);
xnor U27622 (N_27622,N_27461,N_27393);
nor U27623 (N_27623,N_27420,N_27185);
or U27624 (N_27624,N_27443,N_27124);
nor U27625 (N_27625,N_27139,N_27004);
or U27626 (N_27626,N_27099,N_27162);
xnor U27627 (N_27627,N_27465,N_27378);
nand U27628 (N_27628,N_27215,N_27088);
or U27629 (N_27629,N_27079,N_27189);
nand U27630 (N_27630,N_27321,N_27255);
nand U27631 (N_27631,N_27457,N_27233);
nand U27632 (N_27632,N_27319,N_27265);
nor U27633 (N_27633,N_27462,N_27155);
nand U27634 (N_27634,N_27491,N_27387);
and U27635 (N_27635,N_27249,N_27122);
nand U27636 (N_27636,N_27095,N_27101);
nor U27637 (N_27637,N_27267,N_27193);
nand U27638 (N_27638,N_27044,N_27167);
nand U27639 (N_27639,N_27077,N_27090);
and U27640 (N_27640,N_27146,N_27398);
nor U27641 (N_27641,N_27229,N_27263);
or U27642 (N_27642,N_27266,N_27080);
nor U27643 (N_27643,N_27150,N_27449);
nand U27644 (N_27644,N_27032,N_27059);
and U27645 (N_27645,N_27143,N_27259);
xnor U27646 (N_27646,N_27212,N_27057);
and U27647 (N_27647,N_27187,N_27487);
xnor U27648 (N_27648,N_27218,N_27006);
nand U27649 (N_27649,N_27394,N_27482);
nand U27650 (N_27650,N_27256,N_27421);
or U27651 (N_27651,N_27486,N_27401);
xnor U27652 (N_27652,N_27045,N_27102);
xnor U27653 (N_27653,N_27144,N_27257);
nor U27654 (N_27654,N_27046,N_27331);
or U27655 (N_27655,N_27236,N_27250);
nand U27656 (N_27656,N_27027,N_27344);
xor U27657 (N_27657,N_27445,N_27087);
xnor U27658 (N_27658,N_27176,N_27061);
and U27659 (N_27659,N_27314,N_27402);
nor U27660 (N_27660,N_27411,N_27007);
nor U27661 (N_27661,N_27416,N_27303);
nor U27662 (N_27662,N_27017,N_27037);
and U27663 (N_27663,N_27232,N_27067);
or U27664 (N_27664,N_27469,N_27390);
nand U27665 (N_27665,N_27217,N_27184);
nor U27666 (N_27666,N_27360,N_27038);
xor U27667 (N_27667,N_27230,N_27307);
xnor U27668 (N_27668,N_27159,N_27114);
and U27669 (N_27669,N_27483,N_27248);
and U27670 (N_27670,N_27297,N_27432);
nand U27671 (N_27671,N_27009,N_27428);
and U27672 (N_27672,N_27039,N_27400);
nor U27673 (N_27673,N_27494,N_27301);
and U27674 (N_27674,N_27148,N_27262);
xnor U27675 (N_27675,N_27195,N_27499);
and U27676 (N_27676,N_27126,N_27013);
nand U27677 (N_27677,N_27288,N_27136);
or U27678 (N_27678,N_27000,N_27093);
and U27679 (N_27679,N_27113,N_27261);
nand U27680 (N_27680,N_27170,N_27086);
nand U27681 (N_27681,N_27455,N_27427);
nand U27682 (N_27682,N_27351,N_27111);
and U27683 (N_27683,N_27177,N_27270);
nand U27684 (N_27684,N_27072,N_27363);
and U27685 (N_27685,N_27011,N_27169);
xor U27686 (N_27686,N_27014,N_27382);
or U27687 (N_27687,N_27181,N_27172);
and U27688 (N_27688,N_27470,N_27182);
or U27689 (N_27689,N_27030,N_27438);
nor U27690 (N_27690,N_27240,N_27227);
nand U27691 (N_27691,N_27489,N_27336);
and U27692 (N_27692,N_27002,N_27442);
nor U27693 (N_27693,N_27330,N_27197);
xor U27694 (N_27694,N_27286,N_27040);
nor U27695 (N_27695,N_27273,N_27306);
nor U27696 (N_27696,N_27121,N_27247);
nand U27697 (N_27697,N_27142,N_27446);
or U27698 (N_27698,N_27208,N_27327);
nor U27699 (N_27699,N_27109,N_27346);
and U27700 (N_27700,N_27097,N_27055);
nand U27701 (N_27701,N_27362,N_27357);
nor U27702 (N_27702,N_27366,N_27071);
or U27703 (N_27703,N_27264,N_27389);
or U27704 (N_27704,N_27052,N_27479);
nor U27705 (N_27705,N_27310,N_27496);
xor U27706 (N_27706,N_27190,N_27352);
or U27707 (N_27707,N_27372,N_27311);
or U27708 (N_27708,N_27305,N_27436);
xnor U27709 (N_27709,N_27245,N_27063);
nand U27710 (N_27710,N_27276,N_27200);
or U27711 (N_27711,N_27318,N_27171);
and U27712 (N_27712,N_27222,N_27317);
nor U27713 (N_27713,N_27140,N_27477);
xnor U27714 (N_27714,N_27029,N_27206);
and U27715 (N_27715,N_27041,N_27375);
and U27716 (N_27716,N_27355,N_27385);
xnor U27717 (N_27717,N_27194,N_27152);
xnor U27718 (N_27718,N_27135,N_27451);
xnor U27719 (N_27719,N_27065,N_27128);
nor U27720 (N_27720,N_27376,N_27325);
xnor U27721 (N_27721,N_27498,N_27180);
nand U27722 (N_27722,N_27020,N_27334);
nor U27723 (N_27723,N_27062,N_27049);
nand U27724 (N_27724,N_27096,N_27104);
nor U27725 (N_27725,N_27430,N_27175);
nor U27726 (N_27726,N_27173,N_27178);
nor U27727 (N_27727,N_27015,N_27343);
and U27728 (N_27728,N_27333,N_27399);
or U27729 (N_27729,N_27492,N_27454);
nor U27730 (N_27730,N_27435,N_27437);
and U27731 (N_27731,N_27083,N_27168);
xor U27732 (N_27732,N_27329,N_27106);
or U27733 (N_27733,N_27377,N_27481);
nor U27734 (N_27734,N_27268,N_27324);
xnor U27735 (N_27735,N_27183,N_27359);
nor U27736 (N_27736,N_27426,N_27196);
or U27737 (N_27737,N_27367,N_27413);
or U27738 (N_27738,N_27291,N_27350);
nor U27739 (N_27739,N_27340,N_27471);
nor U27740 (N_27740,N_27203,N_27118);
nor U27741 (N_27741,N_27423,N_27209);
and U27742 (N_27742,N_27231,N_27348);
and U27743 (N_27743,N_27418,N_27452);
xor U27744 (N_27744,N_27406,N_27246);
and U27745 (N_27745,N_27060,N_27164);
or U27746 (N_27746,N_27296,N_27356);
nand U27747 (N_27747,N_27141,N_27205);
nand U27748 (N_27748,N_27293,N_27241);
nor U27749 (N_27749,N_27354,N_27018);
and U27750 (N_27750,N_27025,N_27033);
nor U27751 (N_27751,N_27479,N_27361);
nor U27752 (N_27752,N_27434,N_27162);
xnor U27753 (N_27753,N_27414,N_27382);
nand U27754 (N_27754,N_27053,N_27162);
nor U27755 (N_27755,N_27393,N_27094);
and U27756 (N_27756,N_27246,N_27009);
or U27757 (N_27757,N_27131,N_27181);
nand U27758 (N_27758,N_27234,N_27285);
and U27759 (N_27759,N_27284,N_27036);
nand U27760 (N_27760,N_27049,N_27124);
and U27761 (N_27761,N_27044,N_27490);
nand U27762 (N_27762,N_27143,N_27022);
nor U27763 (N_27763,N_27135,N_27437);
nor U27764 (N_27764,N_27130,N_27173);
and U27765 (N_27765,N_27234,N_27280);
nand U27766 (N_27766,N_27117,N_27399);
nor U27767 (N_27767,N_27057,N_27370);
and U27768 (N_27768,N_27071,N_27491);
nor U27769 (N_27769,N_27283,N_27050);
and U27770 (N_27770,N_27413,N_27120);
nand U27771 (N_27771,N_27183,N_27089);
nor U27772 (N_27772,N_27404,N_27235);
nand U27773 (N_27773,N_27112,N_27275);
or U27774 (N_27774,N_27172,N_27088);
xnor U27775 (N_27775,N_27255,N_27187);
or U27776 (N_27776,N_27137,N_27308);
nand U27777 (N_27777,N_27365,N_27412);
and U27778 (N_27778,N_27125,N_27256);
xnor U27779 (N_27779,N_27283,N_27186);
nor U27780 (N_27780,N_27017,N_27155);
and U27781 (N_27781,N_27272,N_27357);
and U27782 (N_27782,N_27224,N_27126);
and U27783 (N_27783,N_27375,N_27453);
nor U27784 (N_27784,N_27467,N_27050);
nand U27785 (N_27785,N_27285,N_27373);
and U27786 (N_27786,N_27050,N_27188);
xor U27787 (N_27787,N_27258,N_27284);
and U27788 (N_27788,N_27010,N_27047);
or U27789 (N_27789,N_27055,N_27347);
or U27790 (N_27790,N_27374,N_27137);
or U27791 (N_27791,N_27467,N_27472);
or U27792 (N_27792,N_27289,N_27002);
nor U27793 (N_27793,N_27322,N_27086);
nand U27794 (N_27794,N_27165,N_27054);
or U27795 (N_27795,N_27444,N_27217);
nor U27796 (N_27796,N_27122,N_27151);
nand U27797 (N_27797,N_27180,N_27255);
nand U27798 (N_27798,N_27208,N_27288);
and U27799 (N_27799,N_27302,N_27357);
nand U27800 (N_27800,N_27448,N_27445);
or U27801 (N_27801,N_27403,N_27417);
xnor U27802 (N_27802,N_27116,N_27487);
and U27803 (N_27803,N_27293,N_27493);
or U27804 (N_27804,N_27175,N_27481);
or U27805 (N_27805,N_27414,N_27194);
nor U27806 (N_27806,N_27352,N_27444);
or U27807 (N_27807,N_27442,N_27302);
nor U27808 (N_27808,N_27238,N_27282);
nand U27809 (N_27809,N_27194,N_27088);
xnor U27810 (N_27810,N_27051,N_27255);
xor U27811 (N_27811,N_27342,N_27311);
xnor U27812 (N_27812,N_27416,N_27313);
and U27813 (N_27813,N_27341,N_27254);
nand U27814 (N_27814,N_27228,N_27244);
xnor U27815 (N_27815,N_27344,N_27010);
xnor U27816 (N_27816,N_27076,N_27223);
and U27817 (N_27817,N_27101,N_27006);
or U27818 (N_27818,N_27148,N_27246);
xnor U27819 (N_27819,N_27139,N_27002);
xor U27820 (N_27820,N_27372,N_27338);
nor U27821 (N_27821,N_27315,N_27081);
or U27822 (N_27822,N_27326,N_27003);
or U27823 (N_27823,N_27172,N_27091);
nand U27824 (N_27824,N_27258,N_27218);
nand U27825 (N_27825,N_27173,N_27166);
xor U27826 (N_27826,N_27010,N_27369);
or U27827 (N_27827,N_27179,N_27336);
xor U27828 (N_27828,N_27028,N_27234);
nor U27829 (N_27829,N_27408,N_27397);
and U27830 (N_27830,N_27288,N_27194);
nand U27831 (N_27831,N_27417,N_27322);
and U27832 (N_27832,N_27340,N_27382);
xnor U27833 (N_27833,N_27311,N_27482);
nand U27834 (N_27834,N_27248,N_27455);
or U27835 (N_27835,N_27095,N_27447);
or U27836 (N_27836,N_27252,N_27428);
xor U27837 (N_27837,N_27197,N_27358);
or U27838 (N_27838,N_27261,N_27403);
nor U27839 (N_27839,N_27169,N_27004);
and U27840 (N_27840,N_27043,N_27113);
or U27841 (N_27841,N_27402,N_27254);
and U27842 (N_27842,N_27116,N_27491);
nor U27843 (N_27843,N_27404,N_27368);
and U27844 (N_27844,N_27265,N_27212);
or U27845 (N_27845,N_27280,N_27067);
nand U27846 (N_27846,N_27384,N_27363);
or U27847 (N_27847,N_27275,N_27058);
nand U27848 (N_27848,N_27369,N_27494);
and U27849 (N_27849,N_27228,N_27422);
xor U27850 (N_27850,N_27491,N_27464);
or U27851 (N_27851,N_27417,N_27429);
and U27852 (N_27852,N_27282,N_27216);
nor U27853 (N_27853,N_27444,N_27392);
nand U27854 (N_27854,N_27138,N_27276);
nor U27855 (N_27855,N_27166,N_27458);
nor U27856 (N_27856,N_27347,N_27017);
or U27857 (N_27857,N_27396,N_27036);
nor U27858 (N_27858,N_27421,N_27330);
and U27859 (N_27859,N_27350,N_27276);
xnor U27860 (N_27860,N_27352,N_27160);
xor U27861 (N_27861,N_27309,N_27495);
or U27862 (N_27862,N_27362,N_27205);
and U27863 (N_27863,N_27237,N_27007);
xnor U27864 (N_27864,N_27391,N_27160);
xor U27865 (N_27865,N_27283,N_27288);
xor U27866 (N_27866,N_27138,N_27350);
nor U27867 (N_27867,N_27357,N_27497);
xnor U27868 (N_27868,N_27352,N_27167);
and U27869 (N_27869,N_27152,N_27330);
or U27870 (N_27870,N_27096,N_27424);
or U27871 (N_27871,N_27055,N_27234);
xor U27872 (N_27872,N_27308,N_27477);
nand U27873 (N_27873,N_27497,N_27036);
and U27874 (N_27874,N_27283,N_27099);
nand U27875 (N_27875,N_27256,N_27388);
or U27876 (N_27876,N_27228,N_27433);
and U27877 (N_27877,N_27262,N_27074);
or U27878 (N_27878,N_27296,N_27318);
and U27879 (N_27879,N_27258,N_27461);
nand U27880 (N_27880,N_27459,N_27125);
or U27881 (N_27881,N_27235,N_27267);
xor U27882 (N_27882,N_27172,N_27308);
nor U27883 (N_27883,N_27415,N_27380);
or U27884 (N_27884,N_27383,N_27304);
nor U27885 (N_27885,N_27493,N_27366);
nor U27886 (N_27886,N_27040,N_27006);
or U27887 (N_27887,N_27424,N_27260);
or U27888 (N_27888,N_27108,N_27306);
and U27889 (N_27889,N_27340,N_27257);
nand U27890 (N_27890,N_27099,N_27288);
xor U27891 (N_27891,N_27022,N_27150);
and U27892 (N_27892,N_27499,N_27343);
nor U27893 (N_27893,N_27053,N_27399);
xor U27894 (N_27894,N_27011,N_27000);
or U27895 (N_27895,N_27161,N_27181);
xnor U27896 (N_27896,N_27480,N_27062);
xnor U27897 (N_27897,N_27459,N_27187);
and U27898 (N_27898,N_27099,N_27102);
nand U27899 (N_27899,N_27083,N_27470);
xor U27900 (N_27900,N_27270,N_27262);
and U27901 (N_27901,N_27390,N_27340);
or U27902 (N_27902,N_27454,N_27014);
and U27903 (N_27903,N_27438,N_27414);
xnor U27904 (N_27904,N_27476,N_27104);
or U27905 (N_27905,N_27175,N_27006);
or U27906 (N_27906,N_27323,N_27162);
or U27907 (N_27907,N_27442,N_27460);
or U27908 (N_27908,N_27015,N_27397);
or U27909 (N_27909,N_27090,N_27418);
nor U27910 (N_27910,N_27093,N_27493);
nor U27911 (N_27911,N_27407,N_27228);
nor U27912 (N_27912,N_27255,N_27220);
or U27913 (N_27913,N_27001,N_27009);
or U27914 (N_27914,N_27264,N_27139);
and U27915 (N_27915,N_27055,N_27015);
nand U27916 (N_27916,N_27347,N_27441);
nor U27917 (N_27917,N_27173,N_27407);
nand U27918 (N_27918,N_27135,N_27394);
nand U27919 (N_27919,N_27430,N_27074);
and U27920 (N_27920,N_27188,N_27067);
xnor U27921 (N_27921,N_27471,N_27118);
or U27922 (N_27922,N_27271,N_27109);
xor U27923 (N_27923,N_27308,N_27321);
or U27924 (N_27924,N_27297,N_27483);
or U27925 (N_27925,N_27095,N_27316);
nand U27926 (N_27926,N_27224,N_27175);
xor U27927 (N_27927,N_27066,N_27256);
and U27928 (N_27928,N_27447,N_27006);
or U27929 (N_27929,N_27186,N_27006);
nor U27930 (N_27930,N_27078,N_27042);
xor U27931 (N_27931,N_27070,N_27148);
or U27932 (N_27932,N_27226,N_27011);
nor U27933 (N_27933,N_27014,N_27095);
nor U27934 (N_27934,N_27416,N_27352);
and U27935 (N_27935,N_27263,N_27267);
or U27936 (N_27936,N_27390,N_27367);
nand U27937 (N_27937,N_27335,N_27240);
nand U27938 (N_27938,N_27256,N_27469);
nor U27939 (N_27939,N_27376,N_27232);
or U27940 (N_27940,N_27460,N_27453);
xor U27941 (N_27941,N_27257,N_27002);
xor U27942 (N_27942,N_27308,N_27184);
xor U27943 (N_27943,N_27302,N_27106);
nor U27944 (N_27944,N_27125,N_27243);
nand U27945 (N_27945,N_27312,N_27303);
or U27946 (N_27946,N_27167,N_27152);
and U27947 (N_27947,N_27094,N_27211);
nor U27948 (N_27948,N_27020,N_27406);
nor U27949 (N_27949,N_27325,N_27153);
or U27950 (N_27950,N_27258,N_27423);
xor U27951 (N_27951,N_27176,N_27170);
xor U27952 (N_27952,N_27480,N_27353);
or U27953 (N_27953,N_27257,N_27174);
nor U27954 (N_27954,N_27087,N_27118);
xnor U27955 (N_27955,N_27423,N_27415);
nor U27956 (N_27956,N_27098,N_27067);
nor U27957 (N_27957,N_27380,N_27175);
or U27958 (N_27958,N_27227,N_27483);
nor U27959 (N_27959,N_27013,N_27368);
xnor U27960 (N_27960,N_27042,N_27446);
nor U27961 (N_27961,N_27017,N_27117);
xor U27962 (N_27962,N_27005,N_27258);
and U27963 (N_27963,N_27435,N_27400);
or U27964 (N_27964,N_27353,N_27018);
nand U27965 (N_27965,N_27099,N_27094);
nand U27966 (N_27966,N_27473,N_27048);
nand U27967 (N_27967,N_27315,N_27316);
nand U27968 (N_27968,N_27372,N_27096);
nor U27969 (N_27969,N_27443,N_27089);
or U27970 (N_27970,N_27461,N_27159);
xor U27971 (N_27971,N_27289,N_27161);
nor U27972 (N_27972,N_27091,N_27090);
nor U27973 (N_27973,N_27054,N_27076);
nor U27974 (N_27974,N_27430,N_27028);
and U27975 (N_27975,N_27008,N_27444);
xor U27976 (N_27976,N_27369,N_27018);
or U27977 (N_27977,N_27429,N_27323);
nor U27978 (N_27978,N_27457,N_27199);
nor U27979 (N_27979,N_27360,N_27467);
nand U27980 (N_27980,N_27490,N_27165);
nor U27981 (N_27981,N_27359,N_27431);
xnor U27982 (N_27982,N_27313,N_27055);
nor U27983 (N_27983,N_27433,N_27359);
or U27984 (N_27984,N_27130,N_27190);
and U27985 (N_27985,N_27041,N_27301);
nor U27986 (N_27986,N_27297,N_27477);
nand U27987 (N_27987,N_27231,N_27490);
xor U27988 (N_27988,N_27202,N_27360);
and U27989 (N_27989,N_27494,N_27272);
or U27990 (N_27990,N_27131,N_27301);
nor U27991 (N_27991,N_27287,N_27157);
or U27992 (N_27992,N_27476,N_27436);
nand U27993 (N_27993,N_27368,N_27111);
and U27994 (N_27994,N_27298,N_27415);
and U27995 (N_27995,N_27096,N_27436);
and U27996 (N_27996,N_27426,N_27065);
xnor U27997 (N_27997,N_27018,N_27180);
or U27998 (N_27998,N_27149,N_27267);
or U27999 (N_27999,N_27455,N_27473);
nand U28000 (N_28000,N_27883,N_27932);
and U28001 (N_28001,N_27948,N_27995);
nand U28002 (N_28002,N_27787,N_27881);
nor U28003 (N_28003,N_27855,N_27928);
nand U28004 (N_28004,N_27771,N_27743);
and U28005 (N_28005,N_27974,N_27624);
xor U28006 (N_28006,N_27584,N_27651);
nor U28007 (N_28007,N_27941,N_27655);
or U28008 (N_28008,N_27814,N_27888);
nor U28009 (N_28009,N_27508,N_27964);
and U28010 (N_28010,N_27605,N_27644);
nor U28011 (N_28011,N_27671,N_27969);
or U28012 (N_28012,N_27954,N_27816);
nor U28013 (N_28013,N_27763,N_27933);
nand U28014 (N_28014,N_27632,N_27838);
and U28015 (N_28015,N_27819,N_27746);
or U28016 (N_28016,N_27502,N_27802);
nor U28017 (N_28017,N_27976,N_27693);
and U28018 (N_28018,N_27989,N_27872);
and U28019 (N_28019,N_27526,N_27772);
nand U28020 (N_28020,N_27952,N_27507);
and U28021 (N_28021,N_27768,N_27839);
xnor U28022 (N_28022,N_27524,N_27650);
or U28023 (N_28023,N_27505,N_27805);
or U28024 (N_28024,N_27596,N_27555);
xor U28025 (N_28025,N_27694,N_27984);
xor U28026 (N_28026,N_27585,N_27737);
nand U28027 (N_28027,N_27884,N_27797);
xor U28028 (N_28028,N_27527,N_27504);
nand U28029 (N_28029,N_27779,N_27593);
or U28030 (N_28030,N_27675,N_27597);
nand U28031 (N_28031,N_27638,N_27545);
or U28032 (N_28032,N_27923,N_27701);
nor U28033 (N_28033,N_27576,N_27601);
xnor U28034 (N_28034,N_27525,N_27652);
nor U28035 (N_28035,N_27854,N_27582);
nor U28036 (N_28036,N_27621,N_27868);
nor U28037 (N_28037,N_27692,N_27600);
nor U28038 (N_28038,N_27796,N_27960);
xor U28039 (N_28039,N_27702,N_27587);
or U28040 (N_28040,N_27800,N_27707);
or U28041 (N_28041,N_27871,N_27950);
xnor U28042 (N_28042,N_27677,N_27935);
and U28043 (N_28043,N_27536,N_27939);
xnor U28044 (N_28044,N_27734,N_27660);
or U28045 (N_28045,N_27942,N_27885);
xor U28046 (N_28046,N_27685,N_27682);
nor U28047 (N_28047,N_27759,N_27560);
nand U28048 (N_28048,N_27554,N_27653);
or U28049 (N_28049,N_27611,N_27519);
nor U28050 (N_28050,N_27945,N_27717);
nand U28051 (N_28051,N_27997,N_27756);
xor U28052 (N_28052,N_27637,N_27999);
nand U28053 (N_28053,N_27711,N_27781);
and U28054 (N_28054,N_27616,N_27532);
and U28055 (N_28055,N_27573,N_27609);
xor U28056 (N_28056,N_27983,N_27518);
xnor U28057 (N_28057,N_27861,N_27667);
nor U28058 (N_28058,N_27506,N_27801);
nor U28059 (N_28059,N_27808,N_27748);
nand U28060 (N_28060,N_27914,N_27846);
xor U28061 (N_28061,N_27674,N_27543);
nor U28062 (N_28062,N_27911,N_27656);
or U28063 (N_28063,N_27956,N_27835);
and U28064 (N_28064,N_27842,N_27889);
xnor U28065 (N_28065,N_27698,N_27988);
or U28066 (N_28066,N_27908,N_27934);
nor U28067 (N_28067,N_27912,N_27552);
or U28068 (N_28068,N_27864,N_27625);
and U28069 (N_28069,N_27684,N_27687);
or U28070 (N_28070,N_27982,N_27794);
and U28071 (N_28071,N_27567,N_27892);
xor U28072 (N_28072,N_27869,N_27586);
nor U28073 (N_28073,N_27641,N_27940);
nor U28074 (N_28074,N_27957,N_27930);
nor U28075 (N_28075,N_27968,N_27673);
nand U28076 (N_28076,N_27817,N_27509);
xor U28077 (N_28077,N_27810,N_27635);
and U28078 (N_28078,N_27785,N_27961);
or U28079 (N_28079,N_27870,N_27538);
xor U28080 (N_28080,N_27858,N_27548);
xor U28081 (N_28081,N_27840,N_27773);
nand U28082 (N_28082,N_27517,N_27774);
nand U28083 (N_28083,N_27708,N_27766);
and U28084 (N_28084,N_27725,N_27919);
nor U28085 (N_28085,N_27829,N_27970);
and U28086 (N_28086,N_27991,N_27521);
nor U28087 (N_28087,N_27823,N_27513);
xor U28088 (N_28088,N_27965,N_27613);
nor U28089 (N_28089,N_27683,N_27972);
and U28090 (N_28090,N_27886,N_27668);
and U28091 (N_28091,N_27583,N_27899);
xor U28092 (N_28092,N_27998,N_27818);
nand U28093 (N_28093,N_27726,N_27857);
xor U28094 (N_28094,N_27903,N_27561);
nor U28095 (N_28095,N_27845,N_27657);
and U28096 (N_28096,N_27691,N_27792);
nor U28097 (N_28097,N_27994,N_27849);
and U28098 (N_28098,N_27764,N_27672);
nor U28099 (N_28099,N_27670,N_27703);
and U28100 (N_28100,N_27880,N_27736);
or U28101 (N_28101,N_27893,N_27580);
nor U28102 (N_28102,N_27769,N_27742);
or U28103 (N_28103,N_27733,N_27966);
nor U28104 (N_28104,N_27887,N_27907);
nand U28105 (N_28105,N_27809,N_27744);
xor U28106 (N_28106,N_27806,N_27782);
nand U28107 (N_28107,N_27522,N_27891);
or U28108 (N_28108,N_27757,N_27709);
nand U28109 (N_28109,N_27859,N_27619);
or U28110 (N_28110,N_27588,N_27570);
and U28111 (N_28111,N_27865,N_27546);
xor U28112 (N_28112,N_27544,N_27550);
nand U28113 (N_28113,N_27662,N_27730);
nor U28114 (N_28114,N_27936,N_27658);
nor U28115 (N_28115,N_27535,N_27705);
nand U28116 (N_28116,N_27811,N_27804);
and U28117 (N_28117,N_27501,N_27634);
or U28118 (N_28118,N_27738,N_27761);
or U28119 (N_28119,N_27990,N_27595);
xnor U28120 (N_28120,N_27719,N_27831);
xnor U28121 (N_28121,N_27747,N_27788);
nand U28122 (N_28122,N_27847,N_27754);
nor U28123 (N_28123,N_27514,N_27944);
xnor U28124 (N_28124,N_27723,N_27803);
and U28125 (N_28125,N_27895,N_27851);
or U28126 (N_28126,N_27649,N_27610);
nand U28127 (N_28127,N_27775,N_27973);
and U28128 (N_28128,N_27876,N_27834);
or U28129 (N_28129,N_27791,N_27510);
and U28130 (N_28130,N_27700,N_27760);
xnor U28131 (N_28131,N_27607,N_27904);
or U28132 (N_28132,N_27712,N_27572);
nand U28133 (N_28133,N_27617,N_27777);
or U28134 (N_28134,N_27598,N_27790);
nor U28135 (N_28135,N_27987,N_27820);
nand U28136 (N_28136,N_27951,N_27843);
and U28137 (N_28137,N_27853,N_27530);
and U28138 (N_28138,N_27755,N_27828);
nand U28139 (N_28139,N_27537,N_27762);
and U28140 (N_28140,N_27967,N_27827);
or U28141 (N_28141,N_27955,N_27867);
and U28142 (N_28142,N_27556,N_27750);
or U28143 (N_28143,N_27993,N_27629);
nor U28144 (N_28144,N_27962,N_27647);
and U28145 (N_28145,N_27825,N_27978);
nor U28146 (N_28146,N_27837,N_27648);
xnor U28147 (N_28147,N_27699,N_27710);
nor U28148 (N_28148,N_27640,N_27614);
nor U28149 (N_28149,N_27589,N_27669);
xor U28150 (N_28150,N_27929,N_27676);
and U28151 (N_28151,N_27793,N_27542);
and U28152 (N_28152,N_27549,N_27848);
xnor U28153 (N_28153,N_27592,N_27992);
or U28154 (N_28154,N_27830,N_27778);
or U28155 (N_28155,N_27953,N_27665);
or U28156 (N_28156,N_27776,N_27630);
or U28157 (N_28157,N_27696,N_27946);
nand U28158 (N_28158,N_27566,N_27515);
nor U28159 (N_28159,N_27979,N_27666);
nand U28160 (N_28160,N_27689,N_27679);
or U28161 (N_28161,N_27645,N_27852);
or U28162 (N_28162,N_27821,N_27765);
xnor U28163 (N_28163,N_27822,N_27639);
and U28164 (N_28164,N_27716,N_27620);
xor U28165 (N_28165,N_27558,N_27623);
nand U28166 (N_28166,N_27841,N_27905);
nand U28167 (N_28167,N_27959,N_27654);
nand U28168 (N_28168,N_27815,N_27863);
nor U28169 (N_28169,N_27920,N_27915);
and U28170 (N_28170,N_27751,N_27579);
xnor U28171 (N_28171,N_27996,N_27882);
or U28172 (N_28172,N_27523,N_27900);
and U28173 (N_28173,N_27569,N_27547);
and U28174 (N_28174,N_27926,N_27896);
nor U28175 (N_28175,N_27500,N_27780);
and U28176 (N_28176,N_27874,N_27531);
nor U28177 (N_28177,N_27784,N_27836);
or U28178 (N_28178,N_27799,N_27602);
nor U28179 (N_28179,N_27807,N_27752);
xor U28180 (N_28180,N_27599,N_27947);
and U28181 (N_28181,N_27688,N_27866);
xor U28182 (N_28182,N_27590,N_27913);
or U28183 (N_28183,N_27713,N_27562);
and U28184 (N_28184,N_27875,N_27520);
xor U28185 (N_28185,N_27910,N_27690);
nor U28186 (N_28186,N_27975,N_27578);
xnor U28187 (N_28187,N_27844,N_27557);
xor U28188 (N_28188,N_27745,N_27902);
or U28189 (N_28189,N_27714,N_27606);
and U28190 (N_28190,N_27512,N_27618);
nor U28191 (N_28191,N_27581,N_27732);
nor U28192 (N_28192,N_27901,N_27938);
xnor U28193 (N_28193,N_27539,N_27873);
and U28194 (N_28194,N_27722,N_27971);
xnor U28195 (N_28195,N_27541,N_27678);
and U28196 (N_28196,N_27894,N_27642);
nand U28197 (N_28197,N_27724,N_27878);
nand U28198 (N_28198,N_27663,N_27511);
nand U28199 (N_28199,N_27856,N_27626);
or U28200 (N_28200,N_27917,N_27937);
nor U28201 (N_28201,N_27704,N_27516);
xor U28202 (N_28202,N_27718,N_27664);
xnor U28203 (N_28203,N_27628,N_27575);
nor U28204 (N_28204,N_27559,N_27798);
and U28205 (N_28205,N_27706,N_27897);
nand U28206 (N_28206,N_27720,N_27826);
nor U28207 (N_28207,N_27604,N_27949);
and U28208 (N_28208,N_27577,N_27918);
xnor U28209 (N_28209,N_27770,N_27812);
and U28210 (N_28210,N_27727,N_27922);
or U28211 (N_28211,N_27615,N_27728);
xnor U28212 (N_28212,N_27980,N_27659);
and U28213 (N_28213,N_27608,N_27563);
nor U28214 (N_28214,N_27553,N_27731);
nor U28215 (N_28215,N_27646,N_27565);
xnor U28216 (N_28216,N_27643,N_27877);
nor U28217 (N_28217,N_27833,N_27528);
xor U28218 (N_28218,N_27695,N_27977);
or U28219 (N_28219,N_27879,N_27574);
and U28220 (N_28220,N_27925,N_27749);
and U28221 (N_28221,N_27927,N_27681);
xnor U28222 (N_28222,N_27729,N_27622);
nand U28223 (N_28223,N_27850,N_27783);
xor U28224 (N_28224,N_27594,N_27862);
nand U28225 (N_28225,N_27931,N_27890);
xnor U28226 (N_28226,N_27916,N_27758);
nor U28227 (N_28227,N_27571,N_27568);
nand U28228 (N_28228,N_27981,N_27612);
or U28229 (N_28229,N_27789,N_27697);
nand U28230 (N_28230,N_27921,N_27898);
xor U28231 (N_28231,N_27603,N_27963);
xnor U28232 (N_28232,N_27721,N_27813);
or U28233 (N_28233,N_27551,N_27906);
xor U28234 (N_28234,N_27740,N_27753);
nand U28235 (N_28235,N_27786,N_27503);
and U28236 (N_28236,N_27680,N_27686);
xnor U28237 (N_28237,N_27533,N_27739);
xor U28238 (N_28238,N_27985,N_27735);
xor U28239 (N_28239,N_27924,N_27943);
xnor U28240 (N_28240,N_27529,N_27636);
or U28241 (N_28241,N_27909,N_27860);
and U28242 (N_28242,N_27795,N_27958);
or U28243 (N_28243,N_27534,N_27767);
and U28244 (N_28244,N_27564,N_27986);
nand U28245 (N_28245,N_27540,N_27591);
and U28246 (N_28246,N_27824,N_27633);
nand U28247 (N_28247,N_27741,N_27631);
and U28248 (N_28248,N_27715,N_27832);
xnor U28249 (N_28249,N_27627,N_27661);
and U28250 (N_28250,N_27781,N_27844);
and U28251 (N_28251,N_27702,N_27870);
and U28252 (N_28252,N_27902,N_27934);
nor U28253 (N_28253,N_27729,N_27735);
nor U28254 (N_28254,N_27909,N_27550);
nor U28255 (N_28255,N_27687,N_27987);
or U28256 (N_28256,N_27880,N_27826);
nand U28257 (N_28257,N_27764,N_27747);
and U28258 (N_28258,N_27598,N_27943);
nor U28259 (N_28259,N_27542,N_27676);
and U28260 (N_28260,N_27885,N_27886);
or U28261 (N_28261,N_27570,N_27799);
xor U28262 (N_28262,N_27945,N_27547);
xor U28263 (N_28263,N_27939,N_27898);
and U28264 (N_28264,N_27661,N_27519);
xor U28265 (N_28265,N_27589,N_27926);
or U28266 (N_28266,N_27573,N_27819);
and U28267 (N_28267,N_27816,N_27647);
xor U28268 (N_28268,N_27796,N_27862);
nor U28269 (N_28269,N_27760,N_27548);
nor U28270 (N_28270,N_27616,N_27650);
nor U28271 (N_28271,N_27858,N_27640);
nor U28272 (N_28272,N_27840,N_27833);
and U28273 (N_28273,N_27945,N_27736);
xnor U28274 (N_28274,N_27998,N_27844);
or U28275 (N_28275,N_27527,N_27893);
and U28276 (N_28276,N_27565,N_27622);
nor U28277 (N_28277,N_27916,N_27713);
or U28278 (N_28278,N_27551,N_27953);
and U28279 (N_28279,N_27600,N_27552);
nor U28280 (N_28280,N_27685,N_27963);
and U28281 (N_28281,N_27667,N_27733);
or U28282 (N_28282,N_27595,N_27965);
or U28283 (N_28283,N_27565,N_27634);
nor U28284 (N_28284,N_27806,N_27597);
or U28285 (N_28285,N_27536,N_27650);
xnor U28286 (N_28286,N_27574,N_27750);
and U28287 (N_28287,N_27699,N_27719);
and U28288 (N_28288,N_27692,N_27988);
or U28289 (N_28289,N_27900,N_27914);
or U28290 (N_28290,N_27925,N_27772);
nand U28291 (N_28291,N_27712,N_27705);
xor U28292 (N_28292,N_27508,N_27806);
or U28293 (N_28293,N_27748,N_27662);
or U28294 (N_28294,N_27506,N_27896);
nand U28295 (N_28295,N_27979,N_27920);
nor U28296 (N_28296,N_27736,N_27886);
or U28297 (N_28297,N_27583,N_27986);
nand U28298 (N_28298,N_27669,N_27536);
and U28299 (N_28299,N_27703,N_27511);
and U28300 (N_28300,N_27614,N_27603);
nand U28301 (N_28301,N_27868,N_27748);
xor U28302 (N_28302,N_27771,N_27585);
nand U28303 (N_28303,N_27873,N_27833);
nor U28304 (N_28304,N_27918,N_27673);
nand U28305 (N_28305,N_27658,N_27901);
or U28306 (N_28306,N_27853,N_27906);
xor U28307 (N_28307,N_27840,N_27981);
or U28308 (N_28308,N_27788,N_27783);
nand U28309 (N_28309,N_27663,N_27974);
nand U28310 (N_28310,N_27757,N_27524);
and U28311 (N_28311,N_27822,N_27504);
nand U28312 (N_28312,N_27587,N_27903);
or U28313 (N_28313,N_27656,N_27801);
nor U28314 (N_28314,N_27728,N_27962);
xnor U28315 (N_28315,N_27832,N_27525);
nor U28316 (N_28316,N_27763,N_27559);
nor U28317 (N_28317,N_27543,N_27782);
nand U28318 (N_28318,N_27689,N_27694);
and U28319 (N_28319,N_27786,N_27816);
xnor U28320 (N_28320,N_27732,N_27653);
or U28321 (N_28321,N_27852,N_27614);
nand U28322 (N_28322,N_27972,N_27529);
nand U28323 (N_28323,N_27664,N_27587);
nor U28324 (N_28324,N_27746,N_27600);
xnor U28325 (N_28325,N_27859,N_27712);
nor U28326 (N_28326,N_27690,N_27662);
nand U28327 (N_28327,N_27864,N_27651);
nand U28328 (N_28328,N_27770,N_27959);
nor U28329 (N_28329,N_27855,N_27601);
xnor U28330 (N_28330,N_27505,N_27655);
or U28331 (N_28331,N_27843,N_27887);
and U28332 (N_28332,N_27558,N_27642);
nand U28333 (N_28333,N_27720,N_27939);
xor U28334 (N_28334,N_27752,N_27798);
or U28335 (N_28335,N_27915,N_27570);
and U28336 (N_28336,N_27833,N_27737);
xor U28337 (N_28337,N_27503,N_27562);
nor U28338 (N_28338,N_27605,N_27604);
xor U28339 (N_28339,N_27562,N_27875);
or U28340 (N_28340,N_27817,N_27815);
and U28341 (N_28341,N_27604,N_27911);
or U28342 (N_28342,N_27649,N_27693);
nand U28343 (N_28343,N_27703,N_27547);
nand U28344 (N_28344,N_27696,N_27560);
nand U28345 (N_28345,N_27505,N_27929);
nand U28346 (N_28346,N_27871,N_27503);
and U28347 (N_28347,N_27818,N_27964);
nor U28348 (N_28348,N_27891,N_27948);
xor U28349 (N_28349,N_27573,N_27864);
nor U28350 (N_28350,N_27612,N_27676);
xnor U28351 (N_28351,N_27719,N_27743);
and U28352 (N_28352,N_27932,N_27800);
xnor U28353 (N_28353,N_27587,N_27721);
xor U28354 (N_28354,N_27662,N_27708);
nor U28355 (N_28355,N_27614,N_27707);
nor U28356 (N_28356,N_27649,N_27838);
and U28357 (N_28357,N_27803,N_27892);
nor U28358 (N_28358,N_27992,N_27512);
xnor U28359 (N_28359,N_27641,N_27502);
nor U28360 (N_28360,N_27821,N_27675);
or U28361 (N_28361,N_27819,N_27877);
xnor U28362 (N_28362,N_27551,N_27501);
xnor U28363 (N_28363,N_27634,N_27541);
nand U28364 (N_28364,N_27898,N_27645);
nand U28365 (N_28365,N_27724,N_27701);
nand U28366 (N_28366,N_27677,N_27748);
xor U28367 (N_28367,N_27858,N_27623);
nor U28368 (N_28368,N_27789,N_27953);
xnor U28369 (N_28369,N_27850,N_27965);
nor U28370 (N_28370,N_27689,N_27644);
nand U28371 (N_28371,N_27512,N_27561);
and U28372 (N_28372,N_27815,N_27514);
xnor U28373 (N_28373,N_27702,N_27796);
xor U28374 (N_28374,N_27999,N_27760);
and U28375 (N_28375,N_27999,N_27792);
and U28376 (N_28376,N_27771,N_27819);
and U28377 (N_28377,N_27734,N_27569);
and U28378 (N_28378,N_27990,N_27848);
nand U28379 (N_28379,N_27915,N_27643);
xnor U28380 (N_28380,N_27754,N_27846);
xor U28381 (N_28381,N_27644,N_27961);
or U28382 (N_28382,N_27534,N_27969);
nor U28383 (N_28383,N_27680,N_27581);
and U28384 (N_28384,N_27727,N_27724);
nor U28385 (N_28385,N_27849,N_27667);
nand U28386 (N_28386,N_27884,N_27616);
xor U28387 (N_28387,N_27983,N_27782);
nor U28388 (N_28388,N_27805,N_27543);
xor U28389 (N_28389,N_27574,N_27577);
and U28390 (N_28390,N_27666,N_27694);
xor U28391 (N_28391,N_27703,N_27658);
or U28392 (N_28392,N_27655,N_27631);
or U28393 (N_28393,N_27772,N_27765);
xor U28394 (N_28394,N_27542,N_27651);
or U28395 (N_28395,N_27882,N_27625);
and U28396 (N_28396,N_27644,N_27966);
or U28397 (N_28397,N_27985,N_27856);
and U28398 (N_28398,N_27572,N_27577);
xor U28399 (N_28399,N_27714,N_27987);
and U28400 (N_28400,N_27520,N_27967);
or U28401 (N_28401,N_27816,N_27743);
nand U28402 (N_28402,N_27768,N_27725);
and U28403 (N_28403,N_27514,N_27629);
or U28404 (N_28404,N_27672,N_27550);
nand U28405 (N_28405,N_27902,N_27658);
and U28406 (N_28406,N_27790,N_27945);
or U28407 (N_28407,N_27572,N_27872);
nand U28408 (N_28408,N_27653,N_27961);
and U28409 (N_28409,N_27959,N_27677);
nor U28410 (N_28410,N_27730,N_27904);
nor U28411 (N_28411,N_27720,N_27611);
nor U28412 (N_28412,N_27739,N_27577);
and U28413 (N_28413,N_27665,N_27669);
nor U28414 (N_28414,N_27996,N_27824);
nand U28415 (N_28415,N_27826,N_27730);
nor U28416 (N_28416,N_27813,N_27959);
xor U28417 (N_28417,N_27882,N_27997);
nand U28418 (N_28418,N_27928,N_27787);
xor U28419 (N_28419,N_27890,N_27703);
nand U28420 (N_28420,N_27969,N_27928);
and U28421 (N_28421,N_27507,N_27830);
and U28422 (N_28422,N_27817,N_27571);
nor U28423 (N_28423,N_27955,N_27544);
or U28424 (N_28424,N_27727,N_27735);
nand U28425 (N_28425,N_27602,N_27840);
or U28426 (N_28426,N_27698,N_27821);
nor U28427 (N_28427,N_27741,N_27889);
nand U28428 (N_28428,N_27664,N_27683);
and U28429 (N_28429,N_27710,N_27906);
and U28430 (N_28430,N_27635,N_27930);
nor U28431 (N_28431,N_27994,N_27519);
nor U28432 (N_28432,N_27549,N_27877);
nor U28433 (N_28433,N_27940,N_27535);
nor U28434 (N_28434,N_27979,N_27747);
and U28435 (N_28435,N_27891,N_27840);
and U28436 (N_28436,N_27971,N_27653);
xnor U28437 (N_28437,N_27897,N_27722);
xor U28438 (N_28438,N_27940,N_27570);
nor U28439 (N_28439,N_27811,N_27825);
and U28440 (N_28440,N_27955,N_27684);
and U28441 (N_28441,N_27731,N_27701);
nor U28442 (N_28442,N_27711,N_27681);
xnor U28443 (N_28443,N_27549,N_27759);
xor U28444 (N_28444,N_27664,N_27887);
nand U28445 (N_28445,N_27874,N_27969);
nor U28446 (N_28446,N_27932,N_27794);
xor U28447 (N_28447,N_27536,N_27503);
xnor U28448 (N_28448,N_27851,N_27592);
xnor U28449 (N_28449,N_27670,N_27734);
nand U28450 (N_28450,N_27719,N_27712);
and U28451 (N_28451,N_27736,N_27745);
nand U28452 (N_28452,N_27955,N_27548);
xor U28453 (N_28453,N_27533,N_27994);
or U28454 (N_28454,N_27722,N_27609);
or U28455 (N_28455,N_27818,N_27772);
or U28456 (N_28456,N_27852,N_27773);
nand U28457 (N_28457,N_27695,N_27664);
nand U28458 (N_28458,N_27976,N_27503);
or U28459 (N_28459,N_27603,N_27621);
xnor U28460 (N_28460,N_27603,N_27630);
nor U28461 (N_28461,N_27592,N_27612);
nand U28462 (N_28462,N_27599,N_27848);
xor U28463 (N_28463,N_27579,N_27639);
or U28464 (N_28464,N_27873,N_27642);
nand U28465 (N_28465,N_27888,N_27947);
xnor U28466 (N_28466,N_27878,N_27969);
xor U28467 (N_28467,N_27927,N_27627);
nand U28468 (N_28468,N_27997,N_27698);
nor U28469 (N_28469,N_27894,N_27870);
xnor U28470 (N_28470,N_27639,N_27502);
or U28471 (N_28471,N_27979,N_27594);
xnor U28472 (N_28472,N_27623,N_27927);
nand U28473 (N_28473,N_27555,N_27976);
xnor U28474 (N_28474,N_27620,N_27980);
and U28475 (N_28475,N_27572,N_27969);
xnor U28476 (N_28476,N_27748,N_27964);
nor U28477 (N_28477,N_27513,N_27759);
nor U28478 (N_28478,N_27505,N_27658);
xnor U28479 (N_28479,N_27595,N_27668);
nand U28480 (N_28480,N_27531,N_27815);
nand U28481 (N_28481,N_27555,N_27680);
nor U28482 (N_28482,N_27531,N_27837);
nand U28483 (N_28483,N_27841,N_27519);
or U28484 (N_28484,N_27578,N_27704);
nand U28485 (N_28485,N_27760,N_27905);
xnor U28486 (N_28486,N_27703,N_27600);
xnor U28487 (N_28487,N_27517,N_27763);
and U28488 (N_28488,N_27928,N_27846);
xnor U28489 (N_28489,N_27719,N_27794);
nand U28490 (N_28490,N_27746,N_27757);
or U28491 (N_28491,N_27686,N_27742);
and U28492 (N_28492,N_27642,N_27776);
nand U28493 (N_28493,N_27840,N_27620);
xnor U28494 (N_28494,N_27883,N_27831);
nor U28495 (N_28495,N_27938,N_27867);
or U28496 (N_28496,N_27996,N_27697);
and U28497 (N_28497,N_27680,N_27601);
xnor U28498 (N_28498,N_27946,N_27501);
nor U28499 (N_28499,N_27782,N_27545);
xnor U28500 (N_28500,N_28400,N_28456);
xor U28501 (N_28501,N_28247,N_28401);
nand U28502 (N_28502,N_28343,N_28430);
or U28503 (N_28503,N_28313,N_28054);
nor U28504 (N_28504,N_28361,N_28358);
or U28505 (N_28505,N_28292,N_28443);
nand U28506 (N_28506,N_28364,N_28248);
or U28507 (N_28507,N_28479,N_28195);
or U28508 (N_28508,N_28201,N_28229);
or U28509 (N_28509,N_28096,N_28330);
or U28510 (N_28510,N_28373,N_28387);
xnor U28511 (N_28511,N_28133,N_28246);
nor U28512 (N_28512,N_28331,N_28017);
or U28513 (N_28513,N_28356,N_28039);
xor U28514 (N_28514,N_28363,N_28434);
nor U28515 (N_28515,N_28104,N_28348);
or U28516 (N_28516,N_28350,N_28076);
or U28517 (N_28517,N_28252,N_28211);
or U28518 (N_28518,N_28110,N_28448);
nor U28519 (N_28519,N_28389,N_28203);
nor U28520 (N_28520,N_28319,N_28063);
nand U28521 (N_28521,N_28447,N_28134);
nand U28522 (N_28522,N_28200,N_28457);
xor U28523 (N_28523,N_28328,N_28438);
xnor U28524 (N_28524,N_28173,N_28181);
nor U28525 (N_28525,N_28102,N_28496);
and U28526 (N_28526,N_28029,N_28473);
nor U28527 (N_28527,N_28212,N_28235);
xor U28528 (N_28528,N_28048,N_28162);
or U28529 (N_28529,N_28130,N_28255);
xnor U28530 (N_28530,N_28368,N_28204);
xor U28531 (N_28531,N_28440,N_28494);
and U28532 (N_28532,N_28307,N_28390);
nand U28533 (N_28533,N_28106,N_28189);
nor U28534 (N_28534,N_28305,N_28274);
nor U28535 (N_28535,N_28145,N_28069);
or U28536 (N_28536,N_28199,N_28150);
and U28537 (N_28537,N_28367,N_28483);
nor U28538 (N_28538,N_28018,N_28198);
nor U28539 (N_28539,N_28414,N_28061);
nand U28540 (N_28540,N_28013,N_28462);
and U28541 (N_28541,N_28070,N_28445);
nor U28542 (N_28542,N_28410,N_28141);
or U28543 (N_28543,N_28129,N_28239);
or U28544 (N_28544,N_28399,N_28004);
and U28545 (N_28545,N_28275,N_28049);
and U28546 (N_28546,N_28327,N_28345);
or U28547 (N_28547,N_28403,N_28393);
or U28548 (N_28548,N_28135,N_28192);
and U28549 (N_28549,N_28144,N_28472);
nor U28550 (N_28550,N_28059,N_28493);
nand U28551 (N_28551,N_28458,N_28481);
xnor U28552 (N_28552,N_28253,N_28213);
xnor U28553 (N_28553,N_28273,N_28337);
xnor U28554 (N_28554,N_28044,N_28116);
or U28555 (N_28555,N_28001,N_28412);
nor U28556 (N_28556,N_28466,N_28170);
and U28557 (N_28557,N_28261,N_28371);
nand U28558 (N_28558,N_28244,N_28046);
or U28559 (N_28559,N_28446,N_28180);
xnor U28560 (N_28560,N_28107,N_28409);
xor U28561 (N_28561,N_28209,N_28224);
or U28562 (N_28562,N_28487,N_28038);
or U28563 (N_28563,N_28424,N_28171);
and U28564 (N_28564,N_28072,N_28272);
or U28565 (N_28565,N_28202,N_28220);
xnor U28566 (N_28566,N_28080,N_28178);
nand U28567 (N_28567,N_28223,N_28190);
xor U28568 (N_28568,N_28137,N_28056);
xnor U28569 (N_28569,N_28161,N_28113);
and U28570 (N_28570,N_28315,N_28222);
or U28571 (N_28571,N_28094,N_28498);
nor U28572 (N_28572,N_28378,N_28089);
xor U28573 (N_28573,N_28164,N_28084);
and U28574 (N_28574,N_28413,N_28431);
nand U28575 (N_28575,N_28152,N_28132);
nor U28576 (N_28576,N_28158,N_28475);
nand U28577 (N_28577,N_28486,N_28208);
nor U28578 (N_28578,N_28233,N_28395);
nor U28579 (N_28579,N_28035,N_28194);
nor U28580 (N_28580,N_28011,N_28021);
xor U28581 (N_28581,N_28023,N_28022);
or U28582 (N_28582,N_28338,N_28444);
or U28583 (N_28583,N_28168,N_28471);
or U28584 (N_28584,N_28346,N_28262);
and U28585 (N_28585,N_28311,N_28271);
nor U28586 (N_28586,N_28300,N_28303);
and U28587 (N_28587,N_28492,N_28482);
nand U28588 (N_28588,N_28034,N_28065);
and U28589 (N_28589,N_28126,N_28007);
xor U28590 (N_28590,N_28236,N_28344);
or U28591 (N_28591,N_28043,N_28312);
nand U28592 (N_28592,N_28058,N_28416);
xor U28593 (N_28593,N_28016,N_28377);
or U28594 (N_28594,N_28249,N_28294);
and U28595 (N_28595,N_28077,N_28382);
or U28596 (N_28596,N_28278,N_28442);
or U28597 (N_28597,N_28119,N_28226);
nor U28598 (N_28598,N_28341,N_28480);
xnor U28599 (N_28599,N_28075,N_28468);
xor U28600 (N_28600,N_28392,N_28185);
xnor U28601 (N_28601,N_28415,N_28187);
xnor U28602 (N_28602,N_28463,N_28012);
or U28603 (N_28603,N_28231,N_28225);
or U28604 (N_28604,N_28484,N_28398);
nor U28605 (N_28605,N_28435,N_28461);
xnor U28606 (N_28606,N_28386,N_28365);
nor U28607 (N_28607,N_28467,N_28335);
or U28608 (N_28608,N_28040,N_28092);
or U28609 (N_28609,N_28285,N_28301);
or U28610 (N_28610,N_28042,N_28083);
nor U28611 (N_28611,N_28250,N_28028);
xor U28612 (N_28612,N_28115,N_28297);
nand U28613 (N_28613,N_28318,N_28287);
or U28614 (N_28614,N_28347,N_28064);
nor U28615 (N_28615,N_28120,N_28339);
and U28616 (N_28616,N_28153,N_28243);
nand U28617 (N_28617,N_28136,N_28264);
or U28618 (N_28618,N_28032,N_28357);
nor U28619 (N_28619,N_28349,N_28041);
or U28620 (N_28620,N_28423,N_28497);
xor U28621 (N_28621,N_28078,N_28384);
or U28622 (N_28622,N_28045,N_28408);
nor U28623 (N_28623,N_28031,N_28406);
nor U28624 (N_28624,N_28227,N_28138);
nand U28625 (N_28625,N_28323,N_28298);
xor U28626 (N_28626,N_28026,N_28156);
and U28627 (N_28627,N_28407,N_28374);
or U28628 (N_28628,N_28429,N_28140);
nor U28629 (N_28629,N_28436,N_28266);
and U28630 (N_28630,N_28268,N_28205);
or U28631 (N_28631,N_28452,N_28030);
and U28632 (N_28632,N_28432,N_28352);
nand U28633 (N_28633,N_28093,N_28172);
and U28634 (N_28634,N_28295,N_28353);
and U28635 (N_28635,N_28299,N_28010);
and U28636 (N_28636,N_28283,N_28036);
and U28637 (N_28637,N_28169,N_28490);
and U28638 (N_28638,N_28006,N_28216);
nor U28639 (N_28639,N_28385,N_28469);
and U28640 (N_28640,N_28105,N_28183);
and U28641 (N_28641,N_28421,N_28491);
and U28642 (N_28642,N_28288,N_28428);
nand U28643 (N_28643,N_28316,N_28306);
xor U28644 (N_28644,N_28086,N_28476);
nand U28645 (N_28645,N_28304,N_28455);
xnor U28646 (N_28646,N_28279,N_28418);
nor U28647 (N_28647,N_28215,N_28351);
and U28648 (N_28648,N_28121,N_28478);
xor U28649 (N_28649,N_28114,N_28376);
xor U28650 (N_28650,N_28188,N_28117);
or U28651 (N_28651,N_28329,N_28242);
nand U28652 (N_28652,N_28334,N_28217);
nand U28653 (N_28653,N_28112,N_28474);
and U28654 (N_28654,N_28073,N_28097);
xnor U28655 (N_28655,N_28193,N_28196);
nand U28656 (N_28656,N_28459,N_28175);
xor U28657 (N_28657,N_28441,N_28057);
and U28658 (N_28658,N_28055,N_28176);
and U28659 (N_28659,N_28108,N_28100);
and U28660 (N_28660,N_28281,N_28146);
and U28661 (N_28661,N_28383,N_28047);
xor U28662 (N_28662,N_28489,N_28079);
or U28663 (N_28663,N_28182,N_28125);
nor U28664 (N_28664,N_28053,N_28427);
nor U28665 (N_28665,N_28111,N_28081);
nand U28666 (N_28666,N_28355,N_28372);
nor U28667 (N_28667,N_28286,N_28003);
nand U28668 (N_28668,N_28020,N_28166);
or U28669 (N_28669,N_28369,N_28360);
and U28670 (N_28670,N_28333,N_28437);
or U28671 (N_28671,N_28320,N_28159);
and U28672 (N_28672,N_28062,N_28477);
and U28673 (N_28673,N_28082,N_28068);
xor U28674 (N_28674,N_28426,N_28391);
or U28675 (N_28675,N_28085,N_28336);
nand U28676 (N_28676,N_28177,N_28362);
nand U28677 (N_28677,N_28232,N_28422);
and U28678 (N_28678,N_28254,N_28310);
nor U28679 (N_28679,N_28014,N_28005);
nand U28680 (N_28680,N_28263,N_28167);
and U28681 (N_28681,N_28179,N_28277);
xor U28682 (N_28682,N_28396,N_28090);
or U28683 (N_28683,N_28326,N_28375);
nand U28684 (N_28684,N_28219,N_28197);
nor U28685 (N_28685,N_28417,N_28207);
xor U28686 (N_28686,N_28131,N_28454);
or U28687 (N_28687,N_28230,N_28148);
or U28688 (N_28688,N_28381,N_28109);
or U28689 (N_28689,N_28160,N_28221);
nor U28690 (N_28690,N_28228,N_28317);
xnor U28691 (N_28691,N_28139,N_28332);
xnor U28692 (N_28692,N_28433,N_28098);
xnor U28693 (N_28693,N_28280,N_28088);
xnor U28694 (N_28694,N_28025,N_28214);
nand U28695 (N_28695,N_28124,N_28191);
xnor U28696 (N_28696,N_28397,N_28037);
and U28697 (N_28697,N_28128,N_28015);
and U28698 (N_28698,N_28050,N_28302);
nor U28699 (N_28699,N_28149,N_28122);
nor U28700 (N_28700,N_28425,N_28314);
and U28701 (N_28701,N_28103,N_28245);
or U28702 (N_28702,N_28142,N_28269);
nand U28703 (N_28703,N_28052,N_28282);
nand U28704 (N_28704,N_28309,N_28260);
xor U28705 (N_28705,N_28379,N_28450);
and U28706 (N_28706,N_28174,N_28291);
and U28707 (N_28707,N_28206,N_28118);
or U28708 (N_28708,N_28293,N_28470);
or U28709 (N_28709,N_28404,N_28165);
and U28710 (N_28710,N_28258,N_28411);
xor U28711 (N_28711,N_28289,N_28051);
xor U28712 (N_28712,N_28060,N_28002);
nand U28713 (N_28713,N_28308,N_28123);
or U28714 (N_28714,N_28066,N_28276);
xnor U28715 (N_28715,N_28256,N_28019);
or U28716 (N_28716,N_28420,N_28354);
and U28717 (N_28717,N_28067,N_28184);
nand U28718 (N_28718,N_28027,N_28465);
nand U28719 (N_28719,N_28210,N_28143);
or U28720 (N_28720,N_28074,N_28322);
or U28721 (N_28721,N_28449,N_28240);
nor U28722 (N_28722,N_28451,N_28488);
nand U28723 (N_28723,N_28151,N_28495);
nand U28724 (N_28724,N_28157,N_28237);
xnor U28725 (N_28725,N_28101,N_28325);
or U28726 (N_28726,N_28241,N_28155);
xor U28727 (N_28727,N_28405,N_28460);
and U28728 (N_28728,N_28499,N_28270);
and U28729 (N_28729,N_28259,N_28380);
nand U28730 (N_28730,N_28402,N_28284);
xor U28731 (N_28731,N_28464,N_28186);
xnor U28732 (N_28732,N_28127,N_28033);
and U28733 (N_28733,N_28267,N_28095);
or U28734 (N_28734,N_28000,N_28008);
and U28735 (N_28735,N_28394,N_28163);
and U28736 (N_28736,N_28366,N_28290);
xnor U28737 (N_28737,N_28234,N_28024);
xor U28738 (N_28738,N_28439,N_28257);
nor U28739 (N_28739,N_28218,N_28087);
nand U28740 (N_28740,N_28321,N_28419);
xnor U28741 (N_28741,N_28485,N_28359);
nor U28742 (N_28742,N_28453,N_28370);
nor U28743 (N_28743,N_28099,N_28009);
nand U28744 (N_28744,N_28324,N_28154);
or U28745 (N_28745,N_28265,N_28388);
nor U28746 (N_28746,N_28147,N_28340);
nand U28747 (N_28747,N_28071,N_28296);
nand U28748 (N_28748,N_28342,N_28238);
or U28749 (N_28749,N_28091,N_28251);
nor U28750 (N_28750,N_28031,N_28349);
and U28751 (N_28751,N_28329,N_28427);
nand U28752 (N_28752,N_28412,N_28350);
xor U28753 (N_28753,N_28280,N_28492);
xnor U28754 (N_28754,N_28299,N_28107);
nor U28755 (N_28755,N_28016,N_28199);
nand U28756 (N_28756,N_28242,N_28133);
nor U28757 (N_28757,N_28409,N_28442);
xnor U28758 (N_28758,N_28279,N_28426);
nor U28759 (N_28759,N_28009,N_28039);
and U28760 (N_28760,N_28428,N_28123);
and U28761 (N_28761,N_28194,N_28054);
or U28762 (N_28762,N_28481,N_28252);
xnor U28763 (N_28763,N_28069,N_28363);
and U28764 (N_28764,N_28244,N_28416);
xor U28765 (N_28765,N_28259,N_28451);
nor U28766 (N_28766,N_28168,N_28421);
nand U28767 (N_28767,N_28232,N_28322);
nor U28768 (N_28768,N_28261,N_28383);
nand U28769 (N_28769,N_28117,N_28031);
nor U28770 (N_28770,N_28125,N_28476);
nor U28771 (N_28771,N_28359,N_28058);
nand U28772 (N_28772,N_28341,N_28323);
and U28773 (N_28773,N_28357,N_28260);
xor U28774 (N_28774,N_28271,N_28170);
nor U28775 (N_28775,N_28181,N_28223);
and U28776 (N_28776,N_28464,N_28395);
xnor U28777 (N_28777,N_28300,N_28100);
or U28778 (N_28778,N_28009,N_28278);
xnor U28779 (N_28779,N_28112,N_28452);
nand U28780 (N_28780,N_28111,N_28171);
or U28781 (N_28781,N_28116,N_28020);
or U28782 (N_28782,N_28490,N_28143);
nor U28783 (N_28783,N_28351,N_28036);
nand U28784 (N_28784,N_28195,N_28269);
or U28785 (N_28785,N_28280,N_28276);
nand U28786 (N_28786,N_28188,N_28040);
xnor U28787 (N_28787,N_28150,N_28428);
nand U28788 (N_28788,N_28311,N_28487);
and U28789 (N_28789,N_28467,N_28149);
nor U28790 (N_28790,N_28430,N_28190);
xnor U28791 (N_28791,N_28051,N_28387);
nand U28792 (N_28792,N_28003,N_28460);
nand U28793 (N_28793,N_28061,N_28241);
xor U28794 (N_28794,N_28443,N_28410);
and U28795 (N_28795,N_28369,N_28418);
nand U28796 (N_28796,N_28449,N_28014);
or U28797 (N_28797,N_28314,N_28233);
nand U28798 (N_28798,N_28006,N_28370);
nor U28799 (N_28799,N_28201,N_28490);
or U28800 (N_28800,N_28210,N_28398);
or U28801 (N_28801,N_28222,N_28104);
xnor U28802 (N_28802,N_28107,N_28389);
or U28803 (N_28803,N_28221,N_28278);
or U28804 (N_28804,N_28328,N_28334);
nand U28805 (N_28805,N_28316,N_28495);
nor U28806 (N_28806,N_28286,N_28369);
nand U28807 (N_28807,N_28451,N_28477);
or U28808 (N_28808,N_28082,N_28483);
xnor U28809 (N_28809,N_28277,N_28249);
or U28810 (N_28810,N_28045,N_28164);
or U28811 (N_28811,N_28486,N_28222);
or U28812 (N_28812,N_28424,N_28333);
nor U28813 (N_28813,N_28139,N_28228);
or U28814 (N_28814,N_28348,N_28474);
or U28815 (N_28815,N_28467,N_28469);
nand U28816 (N_28816,N_28207,N_28014);
xnor U28817 (N_28817,N_28388,N_28293);
nor U28818 (N_28818,N_28343,N_28146);
xnor U28819 (N_28819,N_28037,N_28044);
nor U28820 (N_28820,N_28411,N_28137);
nor U28821 (N_28821,N_28269,N_28276);
or U28822 (N_28822,N_28263,N_28285);
or U28823 (N_28823,N_28215,N_28405);
and U28824 (N_28824,N_28203,N_28250);
xnor U28825 (N_28825,N_28115,N_28412);
xnor U28826 (N_28826,N_28095,N_28447);
and U28827 (N_28827,N_28141,N_28348);
nand U28828 (N_28828,N_28350,N_28131);
xor U28829 (N_28829,N_28409,N_28180);
nand U28830 (N_28830,N_28195,N_28142);
and U28831 (N_28831,N_28492,N_28323);
xor U28832 (N_28832,N_28239,N_28253);
nand U28833 (N_28833,N_28063,N_28099);
or U28834 (N_28834,N_28280,N_28113);
nand U28835 (N_28835,N_28460,N_28167);
and U28836 (N_28836,N_28243,N_28376);
or U28837 (N_28837,N_28276,N_28327);
xor U28838 (N_28838,N_28279,N_28106);
xnor U28839 (N_28839,N_28488,N_28122);
and U28840 (N_28840,N_28110,N_28128);
and U28841 (N_28841,N_28297,N_28383);
xor U28842 (N_28842,N_28091,N_28140);
and U28843 (N_28843,N_28421,N_28063);
or U28844 (N_28844,N_28227,N_28340);
xnor U28845 (N_28845,N_28221,N_28431);
nor U28846 (N_28846,N_28337,N_28496);
or U28847 (N_28847,N_28410,N_28176);
or U28848 (N_28848,N_28204,N_28374);
nor U28849 (N_28849,N_28164,N_28328);
or U28850 (N_28850,N_28308,N_28280);
nor U28851 (N_28851,N_28309,N_28330);
nor U28852 (N_28852,N_28272,N_28377);
or U28853 (N_28853,N_28231,N_28302);
or U28854 (N_28854,N_28408,N_28382);
nand U28855 (N_28855,N_28100,N_28061);
or U28856 (N_28856,N_28381,N_28188);
nor U28857 (N_28857,N_28271,N_28046);
xnor U28858 (N_28858,N_28348,N_28030);
nand U28859 (N_28859,N_28244,N_28427);
nor U28860 (N_28860,N_28156,N_28384);
xnor U28861 (N_28861,N_28292,N_28238);
nand U28862 (N_28862,N_28466,N_28378);
and U28863 (N_28863,N_28170,N_28411);
and U28864 (N_28864,N_28447,N_28365);
and U28865 (N_28865,N_28452,N_28379);
and U28866 (N_28866,N_28242,N_28468);
xor U28867 (N_28867,N_28245,N_28209);
or U28868 (N_28868,N_28263,N_28066);
xor U28869 (N_28869,N_28186,N_28487);
xnor U28870 (N_28870,N_28126,N_28176);
nand U28871 (N_28871,N_28184,N_28412);
or U28872 (N_28872,N_28327,N_28423);
or U28873 (N_28873,N_28084,N_28390);
or U28874 (N_28874,N_28072,N_28331);
xnor U28875 (N_28875,N_28069,N_28025);
nand U28876 (N_28876,N_28056,N_28001);
xor U28877 (N_28877,N_28376,N_28052);
nand U28878 (N_28878,N_28400,N_28388);
nor U28879 (N_28879,N_28235,N_28259);
nand U28880 (N_28880,N_28058,N_28009);
xnor U28881 (N_28881,N_28247,N_28207);
nor U28882 (N_28882,N_28493,N_28381);
xor U28883 (N_28883,N_28447,N_28295);
and U28884 (N_28884,N_28410,N_28211);
xor U28885 (N_28885,N_28042,N_28129);
or U28886 (N_28886,N_28416,N_28065);
nand U28887 (N_28887,N_28193,N_28416);
xnor U28888 (N_28888,N_28414,N_28297);
nand U28889 (N_28889,N_28311,N_28452);
nand U28890 (N_28890,N_28074,N_28351);
and U28891 (N_28891,N_28047,N_28338);
and U28892 (N_28892,N_28437,N_28484);
and U28893 (N_28893,N_28082,N_28366);
or U28894 (N_28894,N_28302,N_28245);
or U28895 (N_28895,N_28406,N_28332);
nand U28896 (N_28896,N_28269,N_28098);
or U28897 (N_28897,N_28285,N_28238);
or U28898 (N_28898,N_28001,N_28422);
or U28899 (N_28899,N_28157,N_28285);
nand U28900 (N_28900,N_28024,N_28238);
nor U28901 (N_28901,N_28103,N_28344);
xor U28902 (N_28902,N_28007,N_28431);
nor U28903 (N_28903,N_28420,N_28132);
or U28904 (N_28904,N_28247,N_28045);
nand U28905 (N_28905,N_28380,N_28404);
xor U28906 (N_28906,N_28016,N_28263);
nand U28907 (N_28907,N_28056,N_28299);
or U28908 (N_28908,N_28182,N_28193);
and U28909 (N_28909,N_28068,N_28190);
nand U28910 (N_28910,N_28117,N_28340);
and U28911 (N_28911,N_28189,N_28099);
nor U28912 (N_28912,N_28273,N_28394);
nor U28913 (N_28913,N_28436,N_28094);
xor U28914 (N_28914,N_28443,N_28260);
xor U28915 (N_28915,N_28479,N_28030);
nand U28916 (N_28916,N_28331,N_28226);
and U28917 (N_28917,N_28070,N_28107);
xor U28918 (N_28918,N_28273,N_28382);
or U28919 (N_28919,N_28360,N_28259);
nand U28920 (N_28920,N_28173,N_28033);
xor U28921 (N_28921,N_28395,N_28497);
nand U28922 (N_28922,N_28485,N_28401);
nand U28923 (N_28923,N_28487,N_28447);
xor U28924 (N_28924,N_28255,N_28415);
nand U28925 (N_28925,N_28153,N_28226);
and U28926 (N_28926,N_28366,N_28214);
xnor U28927 (N_28927,N_28362,N_28316);
xnor U28928 (N_28928,N_28046,N_28154);
nand U28929 (N_28929,N_28008,N_28082);
and U28930 (N_28930,N_28443,N_28143);
xor U28931 (N_28931,N_28447,N_28379);
or U28932 (N_28932,N_28210,N_28014);
nand U28933 (N_28933,N_28122,N_28212);
nor U28934 (N_28934,N_28039,N_28260);
or U28935 (N_28935,N_28386,N_28443);
nor U28936 (N_28936,N_28373,N_28153);
nand U28937 (N_28937,N_28031,N_28385);
nor U28938 (N_28938,N_28312,N_28045);
xnor U28939 (N_28939,N_28130,N_28277);
xor U28940 (N_28940,N_28156,N_28141);
xor U28941 (N_28941,N_28370,N_28223);
xor U28942 (N_28942,N_28220,N_28056);
and U28943 (N_28943,N_28302,N_28455);
xor U28944 (N_28944,N_28137,N_28232);
nand U28945 (N_28945,N_28061,N_28122);
and U28946 (N_28946,N_28436,N_28225);
nor U28947 (N_28947,N_28032,N_28111);
or U28948 (N_28948,N_28175,N_28202);
and U28949 (N_28949,N_28191,N_28018);
nand U28950 (N_28950,N_28288,N_28469);
and U28951 (N_28951,N_28347,N_28496);
or U28952 (N_28952,N_28075,N_28310);
nand U28953 (N_28953,N_28276,N_28421);
and U28954 (N_28954,N_28014,N_28138);
xnor U28955 (N_28955,N_28190,N_28488);
xnor U28956 (N_28956,N_28446,N_28121);
nand U28957 (N_28957,N_28246,N_28001);
or U28958 (N_28958,N_28411,N_28226);
and U28959 (N_28959,N_28194,N_28246);
xnor U28960 (N_28960,N_28383,N_28439);
nor U28961 (N_28961,N_28359,N_28110);
or U28962 (N_28962,N_28356,N_28145);
nand U28963 (N_28963,N_28476,N_28131);
nor U28964 (N_28964,N_28446,N_28295);
nand U28965 (N_28965,N_28051,N_28116);
nand U28966 (N_28966,N_28301,N_28218);
and U28967 (N_28967,N_28447,N_28039);
and U28968 (N_28968,N_28291,N_28242);
nand U28969 (N_28969,N_28461,N_28110);
nor U28970 (N_28970,N_28372,N_28393);
nor U28971 (N_28971,N_28393,N_28180);
nor U28972 (N_28972,N_28110,N_28346);
nand U28973 (N_28973,N_28217,N_28001);
nand U28974 (N_28974,N_28454,N_28486);
nand U28975 (N_28975,N_28055,N_28376);
or U28976 (N_28976,N_28489,N_28055);
xnor U28977 (N_28977,N_28066,N_28028);
or U28978 (N_28978,N_28357,N_28348);
nand U28979 (N_28979,N_28446,N_28265);
xnor U28980 (N_28980,N_28357,N_28408);
nor U28981 (N_28981,N_28084,N_28378);
xor U28982 (N_28982,N_28090,N_28216);
and U28983 (N_28983,N_28409,N_28013);
and U28984 (N_28984,N_28140,N_28215);
nor U28985 (N_28985,N_28370,N_28228);
nand U28986 (N_28986,N_28420,N_28049);
nor U28987 (N_28987,N_28013,N_28188);
nand U28988 (N_28988,N_28322,N_28392);
nand U28989 (N_28989,N_28364,N_28087);
nand U28990 (N_28990,N_28408,N_28107);
and U28991 (N_28991,N_28035,N_28083);
and U28992 (N_28992,N_28308,N_28216);
and U28993 (N_28993,N_28491,N_28193);
and U28994 (N_28994,N_28263,N_28441);
nor U28995 (N_28995,N_28081,N_28087);
nor U28996 (N_28996,N_28127,N_28331);
nand U28997 (N_28997,N_28234,N_28494);
nor U28998 (N_28998,N_28312,N_28002);
xor U28999 (N_28999,N_28422,N_28216);
and U29000 (N_29000,N_28917,N_28674);
and U29001 (N_29001,N_28647,N_28548);
xor U29002 (N_29002,N_28751,N_28598);
or U29003 (N_29003,N_28616,N_28824);
xnor U29004 (N_29004,N_28955,N_28989);
xor U29005 (N_29005,N_28565,N_28878);
nand U29006 (N_29006,N_28743,N_28981);
nand U29007 (N_29007,N_28819,N_28766);
nor U29008 (N_29008,N_28804,N_28756);
or U29009 (N_29009,N_28833,N_28968);
and U29010 (N_29010,N_28737,N_28563);
nor U29011 (N_29011,N_28533,N_28755);
nand U29012 (N_29012,N_28783,N_28534);
nor U29013 (N_29013,N_28599,N_28511);
or U29014 (N_29014,N_28868,N_28893);
nor U29015 (N_29015,N_28520,N_28714);
nor U29016 (N_29016,N_28600,N_28660);
or U29017 (N_29017,N_28710,N_28942);
and U29018 (N_29018,N_28627,N_28589);
nand U29019 (N_29019,N_28650,N_28770);
xnor U29020 (N_29020,N_28894,N_28898);
xnor U29021 (N_29021,N_28946,N_28601);
xnor U29022 (N_29022,N_28906,N_28842);
and U29023 (N_29023,N_28848,N_28811);
and U29024 (N_29024,N_28573,N_28654);
or U29025 (N_29025,N_28966,N_28857);
xnor U29026 (N_29026,N_28618,N_28877);
and U29027 (N_29027,N_28830,N_28813);
nand U29028 (N_29028,N_28584,N_28794);
or U29029 (N_29029,N_28869,N_28965);
xor U29030 (N_29030,N_28789,N_28772);
nor U29031 (N_29031,N_28580,N_28529);
xnor U29032 (N_29032,N_28642,N_28776);
and U29033 (N_29033,N_28542,N_28812);
and U29034 (N_29034,N_28644,N_28960);
nand U29035 (N_29035,N_28708,N_28632);
nand U29036 (N_29036,N_28577,N_28523);
xnor U29037 (N_29037,N_28684,N_28829);
or U29038 (N_29038,N_28891,N_28860);
or U29039 (N_29039,N_28676,N_28905);
and U29040 (N_29040,N_28591,N_28975);
nand U29041 (N_29041,N_28653,N_28866);
nand U29042 (N_29042,N_28793,N_28760);
xor U29043 (N_29043,N_28696,N_28913);
nand U29044 (N_29044,N_28698,N_28639);
and U29045 (N_29045,N_28953,N_28727);
xnor U29046 (N_29046,N_28980,N_28762);
and U29047 (N_29047,N_28934,N_28694);
nand U29048 (N_29048,N_28587,N_28532);
nor U29049 (N_29049,N_28515,N_28550);
and U29050 (N_29050,N_28500,N_28661);
or U29051 (N_29051,N_28881,N_28731);
and U29052 (N_29052,N_28503,N_28918);
xnor U29053 (N_29053,N_28570,N_28861);
or U29054 (N_29054,N_28741,N_28682);
nor U29055 (N_29055,N_28637,N_28739);
nor U29056 (N_29056,N_28909,N_28876);
and U29057 (N_29057,N_28991,N_28502);
and U29058 (N_29058,N_28930,N_28691);
and U29059 (N_29059,N_28662,N_28996);
nand U29060 (N_29060,N_28706,N_28705);
xnor U29061 (N_29061,N_28972,N_28843);
nand U29062 (N_29062,N_28590,N_28790);
or U29063 (N_29063,N_28971,N_28610);
or U29064 (N_29064,N_28865,N_28800);
nor U29065 (N_29065,N_28724,N_28611);
nor U29066 (N_29066,N_28801,N_28621);
nand U29067 (N_29067,N_28973,N_28779);
or U29068 (N_29068,N_28536,N_28717);
nor U29069 (N_29069,N_28720,N_28853);
or U29070 (N_29070,N_28608,N_28513);
or U29071 (N_29071,N_28579,N_28807);
nand U29072 (N_29072,N_28749,N_28753);
xnor U29073 (N_29073,N_28998,N_28867);
or U29074 (N_29074,N_28562,N_28875);
nor U29075 (N_29075,N_28940,N_28526);
or U29076 (N_29076,N_28847,N_28597);
nor U29077 (N_29077,N_28995,N_28754);
xnor U29078 (N_29078,N_28631,N_28612);
xor U29079 (N_29079,N_28667,N_28689);
nand U29080 (N_29080,N_28850,N_28954);
and U29081 (N_29081,N_28634,N_28636);
nand U29082 (N_29082,N_28773,N_28758);
or U29083 (N_29083,N_28509,N_28849);
and U29084 (N_29084,N_28796,N_28912);
nand U29085 (N_29085,N_28537,N_28982);
and U29086 (N_29086,N_28566,N_28752);
nor U29087 (N_29087,N_28962,N_28620);
nor U29088 (N_29088,N_28744,N_28643);
xnor U29089 (N_29089,N_28686,N_28927);
nor U29090 (N_29090,N_28757,N_28967);
xor U29091 (N_29091,N_28508,N_28677);
and U29092 (N_29092,N_28786,N_28568);
and U29093 (N_29093,N_28892,N_28987);
and U29094 (N_29094,N_28540,N_28816);
xor U29095 (N_29095,N_28609,N_28555);
nand U29096 (N_29096,N_28688,N_28748);
nand U29097 (N_29097,N_28514,N_28715);
nand U29098 (N_29098,N_28665,N_28655);
nor U29099 (N_29099,N_28716,N_28528);
nor U29100 (N_29100,N_28903,N_28519);
xor U29101 (N_29101,N_28675,N_28915);
nand U29102 (N_29102,N_28961,N_28896);
xor U29103 (N_29103,N_28806,N_28723);
and U29104 (N_29104,N_28922,N_28659);
xor U29105 (N_29105,N_28571,N_28984);
nand U29106 (N_29106,N_28859,N_28963);
xnor U29107 (N_29107,N_28880,N_28888);
or U29108 (N_29108,N_28864,N_28950);
or U29109 (N_29109,N_28952,N_28777);
xor U29110 (N_29110,N_28846,N_28837);
nor U29111 (N_29111,N_28552,N_28958);
nor U29112 (N_29112,N_28742,N_28551);
xnor U29113 (N_29113,N_28924,N_28910);
or U29114 (N_29114,N_28974,N_28645);
nand U29115 (N_29115,N_28932,N_28992);
and U29116 (N_29116,N_28569,N_28747);
and U29117 (N_29117,N_28535,N_28510);
nand U29118 (N_29118,N_28541,N_28628);
and U29119 (N_29119,N_28761,N_28870);
nor U29120 (N_29120,N_28718,N_28803);
and U29121 (N_29121,N_28858,N_28841);
xor U29122 (N_29122,N_28592,N_28657);
nand U29123 (N_29123,N_28840,N_28889);
nor U29124 (N_29124,N_28985,N_28944);
nand U29125 (N_29125,N_28964,N_28885);
nand U29126 (N_29126,N_28633,N_28671);
and U29127 (N_29127,N_28640,N_28656);
nand U29128 (N_29128,N_28890,N_28651);
nand U29129 (N_29129,N_28736,N_28559);
nor U29130 (N_29130,N_28933,N_28664);
and U29131 (N_29131,N_28818,N_28993);
nor U29132 (N_29132,N_28852,N_28594);
nand U29133 (N_29133,N_28873,N_28778);
and U29134 (N_29134,N_28831,N_28673);
xnor U29135 (N_29135,N_28606,N_28506);
and U29136 (N_29136,N_28521,N_28512);
and U29137 (N_29137,N_28576,N_28745);
xnor U29138 (N_29138,N_28799,N_28516);
and U29139 (N_29139,N_28856,N_28561);
nand U29140 (N_29140,N_28630,N_28554);
xnor U29141 (N_29141,N_28707,N_28558);
xor U29142 (N_29142,N_28539,N_28947);
or U29143 (N_29143,N_28504,N_28795);
nand U29144 (N_29144,N_28926,N_28615);
xnor U29145 (N_29145,N_28557,N_28525);
or U29146 (N_29146,N_28604,N_28740);
or U29147 (N_29147,N_28709,N_28701);
or U29148 (N_29148,N_28638,N_28827);
xor U29149 (N_29149,N_28788,N_28832);
nand U29150 (N_29150,N_28895,N_28919);
nor U29151 (N_29151,N_28828,N_28928);
nand U29152 (N_29152,N_28988,N_28825);
nor U29153 (N_29153,N_28994,N_28680);
or U29154 (N_29154,N_28907,N_28668);
nand U29155 (N_29155,N_28648,N_28863);
and U29156 (N_29156,N_28911,N_28595);
nor U29157 (N_29157,N_28999,N_28874);
xor U29158 (N_29158,N_28970,N_28544);
xnor U29159 (N_29159,N_28791,N_28635);
nor U29160 (N_29160,N_28871,N_28734);
nand U29161 (N_29161,N_28814,N_28602);
nor U29162 (N_29162,N_28951,N_28854);
xnor U29163 (N_29163,N_28619,N_28501);
xnor U29164 (N_29164,N_28768,N_28729);
nor U29165 (N_29165,N_28728,N_28692);
xnor U29166 (N_29166,N_28699,N_28941);
or U29167 (N_29167,N_28901,N_28518);
and U29168 (N_29168,N_28914,N_28957);
nand U29169 (N_29169,N_28738,N_28887);
or U29170 (N_29170,N_28929,N_28605);
nor U29171 (N_29171,N_28583,N_28652);
xnor U29172 (N_29172,N_28641,N_28899);
xor U29173 (N_29173,N_28969,N_28629);
nand U29174 (N_29174,N_28983,N_28826);
or U29175 (N_29175,N_28931,N_28897);
xor U29176 (N_29176,N_28785,N_28775);
nor U29177 (N_29177,N_28774,N_28693);
nand U29178 (N_29178,N_28797,N_28622);
nand U29179 (N_29179,N_28767,N_28663);
nand U29180 (N_29180,N_28530,N_28697);
xnor U29181 (N_29181,N_28531,N_28603);
nor U29182 (N_29182,N_28670,N_28979);
xnor U29183 (N_29183,N_28678,N_28549);
and U29184 (N_29184,N_28704,N_28721);
nand U29185 (N_29185,N_28959,N_28925);
nor U29186 (N_29186,N_28607,N_28582);
nor U29187 (N_29187,N_28817,N_28976);
or U29188 (N_29188,N_28585,N_28556);
nand U29189 (N_29189,N_28681,N_28862);
nor U29190 (N_29190,N_28546,N_28787);
xor U29191 (N_29191,N_28839,N_28908);
nor U29192 (N_29192,N_28527,N_28623);
or U29193 (N_29193,N_28792,N_28939);
or U29194 (N_29194,N_28725,N_28596);
and U29195 (N_29195,N_28505,N_28759);
and U29196 (N_29196,N_28997,N_28543);
xor U29197 (N_29197,N_28733,N_28886);
nor U29198 (N_29198,N_28713,N_28614);
xor U29199 (N_29199,N_28567,N_28879);
and U29200 (N_29200,N_28672,N_28695);
or U29201 (N_29201,N_28937,N_28553);
and U29202 (N_29202,N_28945,N_28820);
nor U29203 (N_29203,N_28517,N_28700);
and U29204 (N_29204,N_28711,N_28703);
nor U29205 (N_29205,N_28732,N_28798);
or U29206 (N_29206,N_28575,N_28624);
nand U29207 (N_29207,N_28572,N_28943);
nand U29208 (N_29208,N_28805,N_28902);
nand U29209 (N_29209,N_28581,N_28883);
nor U29210 (N_29210,N_28683,N_28935);
or U29211 (N_29211,N_28547,N_28834);
nor U29212 (N_29212,N_28522,N_28948);
nor U29213 (N_29213,N_28746,N_28574);
xor U29214 (N_29214,N_28763,N_28685);
or U29215 (N_29215,N_28949,N_28838);
nand U29216 (N_29216,N_28936,N_28538);
or U29217 (N_29217,N_28916,N_28586);
or U29218 (N_29218,N_28564,N_28649);
nand U29219 (N_29219,N_28956,N_28845);
xor U29220 (N_29220,N_28900,N_28750);
nand U29221 (N_29221,N_28810,N_28545);
xnor U29222 (N_29222,N_28617,N_28815);
xor U29223 (N_29223,N_28872,N_28882);
or U29224 (N_29224,N_28802,N_28990);
nand U29225 (N_29225,N_28782,N_28730);
and U29226 (N_29226,N_28822,N_28669);
or U29227 (N_29227,N_28809,N_28507);
nor U29228 (N_29228,N_28986,N_28712);
xor U29229 (N_29229,N_28844,N_28771);
nand U29230 (N_29230,N_28904,N_28524);
nand U29231 (N_29231,N_28613,N_28765);
xor U29232 (N_29232,N_28722,N_28836);
and U29233 (N_29233,N_28978,N_28808);
nor U29234 (N_29234,N_28851,N_28679);
nand U29235 (N_29235,N_28781,N_28719);
or U29236 (N_29236,N_28855,N_28764);
nor U29237 (N_29237,N_28726,N_28920);
and U29238 (N_29238,N_28658,N_28769);
xor U29239 (N_29239,N_28784,N_28593);
or U29240 (N_29240,N_28588,N_28666);
nor U29241 (N_29241,N_28835,N_28884);
nor U29242 (N_29242,N_28823,N_28938);
and U29243 (N_29243,N_28687,N_28923);
xor U29244 (N_29244,N_28578,N_28735);
and U29245 (N_29245,N_28921,N_28560);
nor U29246 (N_29246,N_28821,N_28977);
nor U29247 (N_29247,N_28690,N_28646);
or U29248 (N_29248,N_28626,N_28625);
and U29249 (N_29249,N_28780,N_28702);
nor U29250 (N_29250,N_28649,N_28863);
xnor U29251 (N_29251,N_28550,N_28903);
nor U29252 (N_29252,N_28636,N_28558);
xnor U29253 (N_29253,N_28590,N_28652);
nor U29254 (N_29254,N_28826,N_28603);
nor U29255 (N_29255,N_28980,N_28983);
and U29256 (N_29256,N_28749,N_28742);
or U29257 (N_29257,N_28940,N_28672);
or U29258 (N_29258,N_28988,N_28776);
xor U29259 (N_29259,N_28697,N_28607);
xor U29260 (N_29260,N_28516,N_28842);
nand U29261 (N_29261,N_28702,N_28594);
xnor U29262 (N_29262,N_28506,N_28754);
nand U29263 (N_29263,N_28950,N_28816);
and U29264 (N_29264,N_28534,N_28946);
xor U29265 (N_29265,N_28587,N_28849);
xor U29266 (N_29266,N_28526,N_28989);
and U29267 (N_29267,N_28667,N_28929);
or U29268 (N_29268,N_28563,N_28658);
nor U29269 (N_29269,N_28729,N_28520);
or U29270 (N_29270,N_28987,N_28743);
nand U29271 (N_29271,N_28895,N_28724);
or U29272 (N_29272,N_28892,N_28748);
nand U29273 (N_29273,N_28816,N_28897);
and U29274 (N_29274,N_28779,N_28825);
nor U29275 (N_29275,N_28509,N_28516);
or U29276 (N_29276,N_28983,N_28908);
nand U29277 (N_29277,N_28500,N_28789);
and U29278 (N_29278,N_28606,N_28579);
nor U29279 (N_29279,N_28522,N_28738);
and U29280 (N_29280,N_28506,N_28691);
nor U29281 (N_29281,N_28740,N_28522);
nor U29282 (N_29282,N_28669,N_28930);
xor U29283 (N_29283,N_28680,N_28597);
xor U29284 (N_29284,N_28974,N_28768);
and U29285 (N_29285,N_28798,N_28648);
and U29286 (N_29286,N_28527,N_28689);
and U29287 (N_29287,N_28892,N_28762);
or U29288 (N_29288,N_28621,N_28540);
and U29289 (N_29289,N_28724,N_28966);
xor U29290 (N_29290,N_28976,N_28924);
and U29291 (N_29291,N_28905,N_28826);
xnor U29292 (N_29292,N_28611,N_28741);
and U29293 (N_29293,N_28633,N_28940);
xor U29294 (N_29294,N_28852,N_28795);
nand U29295 (N_29295,N_28547,N_28971);
nor U29296 (N_29296,N_28705,N_28690);
nor U29297 (N_29297,N_28953,N_28935);
and U29298 (N_29298,N_28706,N_28642);
nor U29299 (N_29299,N_28811,N_28879);
or U29300 (N_29300,N_28601,N_28941);
or U29301 (N_29301,N_28910,N_28888);
nor U29302 (N_29302,N_28800,N_28729);
xor U29303 (N_29303,N_28777,N_28652);
and U29304 (N_29304,N_28721,N_28591);
nor U29305 (N_29305,N_28686,N_28719);
or U29306 (N_29306,N_28912,N_28777);
nor U29307 (N_29307,N_28684,N_28720);
or U29308 (N_29308,N_28941,N_28995);
or U29309 (N_29309,N_28694,N_28747);
nand U29310 (N_29310,N_28972,N_28986);
xor U29311 (N_29311,N_28955,N_28829);
xnor U29312 (N_29312,N_28825,N_28898);
nor U29313 (N_29313,N_28896,N_28516);
nand U29314 (N_29314,N_28906,N_28563);
or U29315 (N_29315,N_28877,N_28886);
nor U29316 (N_29316,N_28653,N_28989);
or U29317 (N_29317,N_28621,N_28855);
xnor U29318 (N_29318,N_28831,N_28534);
nand U29319 (N_29319,N_28987,N_28949);
xnor U29320 (N_29320,N_28513,N_28684);
xnor U29321 (N_29321,N_28802,N_28819);
or U29322 (N_29322,N_28671,N_28854);
xor U29323 (N_29323,N_28887,N_28676);
nand U29324 (N_29324,N_28613,N_28514);
xnor U29325 (N_29325,N_28832,N_28859);
and U29326 (N_29326,N_28693,N_28717);
nand U29327 (N_29327,N_28853,N_28873);
or U29328 (N_29328,N_28793,N_28637);
and U29329 (N_29329,N_28524,N_28537);
nor U29330 (N_29330,N_28685,N_28863);
xnor U29331 (N_29331,N_28624,N_28868);
nand U29332 (N_29332,N_28629,N_28931);
xnor U29333 (N_29333,N_28846,N_28649);
xnor U29334 (N_29334,N_28713,N_28949);
xor U29335 (N_29335,N_28609,N_28929);
or U29336 (N_29336,N_28728,N_28716);
xor U29337 (N_29337,N_28711,N_28743);
xor U29338 (N_29338,N_28718,N_28773);
or U29339 (N_29339,N_28811,N_28582);
nand U29340 (N_29340,N_28701,N_28954);
nor U29341 (N_29341,N_28873,N_28848);
xor U29342 (N_29342,N_28977,N_28617);
nor U29343 (N_29343,N_28599,N_28989);
or U29344 (N_29344,N_28567,N_28948);
and U29345 (N_29345,N_28598,N_28969);
nand U29346 (N_29346,N_28828,N_28968);
nand U29347 (N_29347,N_28682,N_28961);
nand U29348 (N_29348,N_28829,N_28745);
nand U29349 (N_29349,N_28770,N_28920);
nor U29350 (N_29350,N_28937,N_28708);
and U29351 (N_29351,N_28666,N_28824);
and U29352 (N_29352,N_28793,N_28942);
nor U29353 (N_29353,N_28711,N_28559);
or U29354 (N_29354,N_28875,N_28668);
and U29355 (N_29355,N_28994,N_28896);
nor U29356 (N_29356,N_28508,N_28517);
or U29357 (N_29357,N_28960,N_28802);
xor U29358 (N_29358,N_28740,N_28520);
and U29359 (N_29359,N_28821,N_28579);
nor U29360 (N_29360,N_28586,N_28998);
nor U29361 (N_29361,N_28517,N_28795);
xnor U29362 (N_29362,N_28765,N_28918);
xnor U29363 (N_29363,N_28937,N_28722);
xnor U29364 (N_29364,N_28783,N_28784);
xnor U29365 (N_29365,N_28738,N_28631);
nor U29366 (N_29366,N_28720,N_28819);
or U29367 (N_29367,N_28938,N_28999);
and U29368 (N_29368,N_28892,N_28607);
or U29369 (N_29369,N_28536,N_28638);
nor U29370 (N_29370,N_28728,N_28697);
xor U29371 (N_29371,N_28759,N_28739);
and U29372 (N_29372,N_28942,N_28825);
or U29373 (N_29373,N_28889,N_28631);
nor U29374 (N_29374,N_28949,N_28626);
nor U29375 (N_29375,N_28918,N_28673);
nand U29376 (N_29376,N_28555,N_28658);
or U29377 (N_29377,N_28567,N_28714);
nor U29378 (N_29378,N_28990,N_28624);
or U29379 (N_29379,N_28718,N_28688);
nor U29380 (N_29380,N_28695,N_28709);
xnor U29381 (N_29381,N_28546,N_28552);
and U29382 (N_29382,N_28806,N_28882);
nand U29383 (N_29383,N_28802,N_28623);
xnor U29384 (N_29384,N_28815,N_28754);
nor U29385 (N_29385,N_28600,N_28615);
nand U29386 (N_29386,N_28648,N_28935);
or U29387 (N_29387,N_28864,N_28757);
xor U29388 (N_29388,N_28527,N_28564);
nand U29389 (N_29389,N_28596,N_28801);
nand U29390 (N_29390,N_28653,N_28842);
nand U29391 (N_29391,N_28931,N_28602);
nor U29392 (N_29392,N_28722,N_28884);
and U29393 (N_29393,N_28983,N_28558);
or U29394 (N_29394,N_28783,N_28519);
and U29395 (N_29395,N_28802,N_28763);
and U29396 (N_29396,N_28929,N_28658);
nand U29397 (N_29397,N_28540,N_28631);
and U29398 (N_29398,N_28882,N_28767);
xor U29399 (N_29399,N_28649,N_28763);
and U29400 (N_29400,N_28801,N_28951);
or U29401 (N_29401,N_28890,N_28758);
nand U29402 (N_29402,N_28863,N_28710);
or U29403 (N_29403,N_28899,N_28850);
xor U29404 (N_29404,N_28507,N_28591);
nand U29405 (N_29405,N_28862,N_28738);
or U29406 (N_29406,N_28920,N_28826);
and U29407 (N_29407,N_28744,N_28751);
nor U29408 (N_29408,N_28757,N_28665);
nor U29409 (N_29409,N_28695,N_28732);
or U29410 (N_29410,N_28843,N_28689);
nand U29411 (N_29411,N_28990,N_28884);
nand U29412 (N_29412,N_28603,N_28915);
nor U29413 (N_29413,N_28742,N_28926);
and U29414 (N_29414,N_28683,N_28620);
or U29415 (N_29415,N_28614,N_28917);
or U29416 (N_29416,N_28607,N_28834);
or U29417 (N_29417,N_28883,N_28732);
nor U29418 (N_29418,N_28774,N_28741);
xor U29419 (N_29419,N_28846,N_28648);
nand U29420 (N_29420,N_28629,N_28887);
and U29421 (N_29421,N_28509,N_28505);
xor U29422 (N_29422,N_28765,N_28806);
nand U29423 (N_29423,N_28756,N_28908);
xnor U29424 (N_29424,N_28739,N_28716);
xor U29425 (N_29425,N_28728,N_28803);
and U29426 (N_29426,N_28504,N_28602);
xor U29427 (N_29427,N_28560,N_28509);
and U29428 (N_29428,N_28997,N_28939);
nand U29429 (N_29429,N_28557,N_28583);
and U29430 (N_29430,N_28875,N_28691);
and U29431 (N_29431,N_28686,N_28842);
nor U29432 (N_29432,N_28503,N_28514);
xnor U29433 (N_29433,N_28516,N_28859);
and U29434 (N_29434,N_28548,N_28683);
xor U29435 (N_29435,N_28935,N_28527);
xor U29436 (N_29436,N_28891,N_28620);
or U29437 (N_29437,N_28925,N_28612);
and U29438 (N_29438,N_28538,N_28897);
nor U29439 (N_29439,N_28587,N_28919);
or U29440 (N_29440,N_28931,N_28763);
and U29441 (N_29441,N_28770,N_28777);
nor U29442 (N_29442,N_28692,N_28786);
nand U29443 (N_29443,N_28838,N_28784);
nand U29444 (N_29444,N_28791,N_28583);
nor U29445 (N_29445,N_28554,N_28885);
xor U29446 (N_29446,N_28906,N_28869);
or U29447 (N_29447,N_28629,N_28723);
nand U29448 (N_29448,N_28767,N_28547);
nand U29449 (N_29449,N_28693,N_28753);
nor U29450 (N_29450,N_28836,N_28874);
and U29451 (N_29451,N_28519,N_28735);
nand U29452 (N_29452,N_28568,N_28815);
nand U29453 (N_29453,N_28881,N_28886);
xor U29454 (N_29454,N_28780,N_28612);
xor U29455 (N_29455,N_28872,N_28720);
or U29456 (N_29456,N_28647,N_28721);
and U29457 (N_29457,N_28759,N_28711);
or U29458 (N_29458,N_28807,N_28701);
or U29459 (N_29459,N_28752,N_28818);
nand U29460 (N_29460,N_28716,N_28614);
or U29461 (N_29461,N_28817,N_28812);
xor U29462 (N_29462,N_28943,N_28708);
nor U29463 (N_29463,N_28922,N_28526);
nand U29464 (N_29464,N_28631,N_28689);
nor U29465 (N_29465,N_28878,N_28981);
nand U29466 (N_29466,N_28652,N_28807);
xor U29467 (N_29467,N_28825,N_28841);
and U29468 (N_29468,N_28515,N_28508);
nor U29469 (N_29469,N_28964,N_28502);
nand U29470 (N_29470,N_28959,N_28665);
nor U29471 (N_29471,N_28580,N_28695);
nor U29472 (N_29472,N_28943,N_28606);
nor U29473 (N_29473,N_28848,N_28933);
and U29474 (N_29474,N_28963,N_28723);
and U29475 (N_29475,N_28852,N_28500);
and U29476 (N_29476,N_28581,N_28620);
and U29477 (N_29477,N_28740,N_28670);
or U29478 (N_29478,N_28893,N_28518);
xnor U29479 (N_29479,N_28544,N_28975);
and U29480 (N_29480,N_28692,N_28759);
or U29481 (N_29481,N_28627,N_28641);
nor U29482 (N_29482,N_28807,N_28725);
and U29483 (N_29483,N_28793,N_28775);
xnor U29484 (N_29484,N_28678,N_28751);
and U29485 (N_29485,N_28958,N_28918);
nand U29486 (N_29486,N_28715,N_28837);
xor U29487 (N_29487,N_28531,N_28557);
and U29488 (N_29488,N_28970,N_28901);
and U29489 (N_29489,N_28746,N_28675);
nor U29490 (N_29490,N_28820,N_28892);
nand U29491 (N_29491,N_28907,N_28821);
nor U29492 (N_29492,N_28641,N_28680);
xnor U29493 (N_29493,N_28877,N_28962);
xnor U29494 (N_29494,N_28760,N_28979);
or U29495 (N_29495,N_28656,N_28601);
or U29496 (N_29496,N_28698,N_28788);
nand U29497 (N_29497,N_28933,N_28949);
or U29498 (N_29498,N_28774,N_28586);
nor U29499 (N_29499,N_28816,N_28995);
nand U29500 (N_29500,N_29032,N_29487);
nor U29501 (N_29501,N_29377,N_29117);
xnor U29502 (N_29502,N_29303,N_29478);
nand U29503 (N_29503,N_29454,N_29451);
nor U29504 (N_29504,N_29205,N_29070);
and U29505 (N_29505,N_29009,N_29271);
nand U29506 (N_29506,N_29179,N_29202);
and U29507 (N_29507,N_29233,N_29291);
nor U29508 (N_29508,N_29068,N_29113);
nand U29509 (N_29509,N_29428,N_29010);
and U29510 (N_29510,N_29211,N_29056);
nand U29511 (N_29511,N_29494,N_29420);
and U29512 (N_29512,N_29363,N_29036);
and U29513 (N_29513,N_29173,N_29258);
nor U29514 (N_29514,N_29488,N_29135);
nor U29515 (N_29515,N_29256,N_29189);
and U29516 (N_29516,N_29027,N_29421);
nor U29517 (N_29517,N_29362,N_29081);
nand U29518 (N_29518,N_29355,N_29482);
nand U29519 (N_29519,N_29318,N_29358);
and U29520 (N_29520,N_29314,N_29402);
xnor U29521 (N_29521,N_29281,N_29394);
and U29522 (N_29522,N_29112,N_29090);
and U29523 (N_29523,N_29151,N_29086);
xor U29524 (N_29524,N_29197,N_29289);
xor U29525 (N_29525,N_29438,N_29134);
xor U29526 (N_29526,N_29450,N_29275);
nand U29527 (N_29527,N_29191,N_29203);
and U29528 (N_29528,N_29263,N_29097);
and U29529 (N_29529,N_29435,N_29120);
xor U29530 (N_29530,N_29472,N_29294);
and U29531 (N_29531,N_29163,N_29194);
or U29532 (N_29532,N_29092,N_29348);
nor U29533 (N_29533,N_29225,N_29388);
nor U29534 (N_29534,N_29221,N_29138);
nand U29535 (N_29535,N_29082,N_29423);
or U29536 (N_29536,N_29442,N_29433);
nand U29537 (N_29537,N_29483,N_29060);
and U29538 (N_29538,N_29003,N_29392);
and U29539 (N_29539,N_29072,N_29401);
nand U29540 (N_29540,N_29033,N_29326);
or U29541 (N_29541,N_29464,N_29150);
xor U29542 (N_29542,N_29108,N_29463);
and U29543 (N_29543,N_29440,N_29029);
xor U29544 (N_29544,N_29195,N_29201);
xnor U29545 (N_29545,N_29279,N_29424);
nand U29546 (N_29546,N_29298,N_29485);
nand U29547 (N_29547,N_29088,N_29245);
nand U29548 (N_29548,N_29218,N_29430);
xnor U29549 (N_29549,N_29213,N_29490);
nand U29550 (N_29550,N_29019,N_29302);
nor U29551 (N_29551,N_29356,N_29414);
xnor U29552 (N_29552,N_29287,N_29210);
or U29553 (N_29553,N_29322,N_29044);
xnor U29554 (N_29554,N_29146,N_29368);
xor U29555 (N_29555,N_29344,N_29354);
xor U29556 (N_29556,N_29389,N_29030);
or U29557 (N_29557,N_29058,N_29071);
xnor U29558 (N_29558,N_29077,N_29057);
xnor U29559 (N_29559,N_29069,N_29028);
xor U29560 (N_29560,N_29396,N_29319);
and U29561 (N_29561,N_29075,N_29481);
xor U29562 (N_29562,N_29361,N_29188);
or U29563 (N_29563,N_29162,N_29214);
nor U29564 (N_29564,N_29448,N_29152);
nand U29565 (N_29565,N_29331,N_29467);
or U29566 (N_29566,N_29419,N_29444);
nand U29567 (N_29567,N_29457,N_29227);
nand U29568 (N_29568,N_29296,N_29373);
or U29569 (N_29569,N_29399,N_29268);
nand U29570 (N_29570,N_29141,N_29224);
and U29571 (N_29571,N_29397,N_29270);
or U29572 (N_29572,N_29063,N_29439);
xnor U29573 (N_29573,N_29094,N_29219);
nand U29574 (N_29574,N_29237,N_29380);
xor U29575 (N_29575,N_29192,N_29048);
xnor U29576 (N_29576,N_29267,N_29431);
and U29577 (N_29577,N_29374,N_29222);
and U29578 (N_29578,N_29025,N_29290);
nor U29579 (N_29579,N_29250,N_29436);
xor U29580 (N_29580,N_29230,N_29198);
or U29581 (N_29581,N_29231,N_29144);
and U29582 (N_29582,N_29473,N_29101);
nand U29583 (N_29583,N_29052,N_29142);
or U29584 (N_29584,N_29080,N_29446);
xor U29585 (N_29585,N_29367,N_29340);
and U29586 (N_29586,N_29262,N_29441);
and U29587 (N_29587,N_29477,N_29334);
nor U29588 (N_29588,N_29257,N_29017);
nor U29589 (N_29589,N_29096,N_29172);
and U29590 (N_29590,N_29165,N_29067);
nand U29591 (N_29591,N_29333,N_29183);
and U29592 (N_29592,N_29105,N_29474);
or U29593 (N_29593,N_29199,N_29342);
nand U29594 (N_29594,N_29427,N_29486);
nand U29595 (N_29595,N_29054,N_29208);
or U29596 (N_29596,N_29286,N_29232);
nor U29597 (N_29597,N_29000,N_29182);
nand U29598 (N_29598,N_29278,N_29372);
and U29599 (N_29599,N_29297,N_29353);
or U29600 (N_29600,N_29498,N_29247);
or U29601 (N_29601,N_29200,N_29371);
or U29602 (N_29602,N_29379,N_29171);
and U29603 (N_29603,N_29242,N_29259);
nand U29604 (N_29604,N_29386,N_29416);
or U29605 (N_29605,N_29137,N_29119);
xnor U29606 (N_29606,N_29404,N_29015);
or U29607 (N_29607,N_29324,N_29468);
xnor U29608 (N_29608,N_29308,N_29492);
and U29609 (N_29609,N_29229,N_29031);
xor U29610 (N_29610,N_29418,N_29083);
xor U29611 (N_29611,N_29124,N_29223);
nand U29612 (N_29612,N_29107,N_29012);
xor U29613 (N_29613,N_29307,N_29384);
or U29614 (N_29614,N_29405,N_29313);
and U29615 (N_29615,N_29338,N_29369);
nor U29616 (N_29616,N_29042,N_29156);
and U29617 (N_29617,N_29304,N_29026);
xor U29618 (N_29618,N_29065,N_29234);
nor U29619 (N_29619,N_29282,N_29274);
or U29620 (N_29620,N_29168,N_29484);
nor U29621 (N_29621,N_29360,N_29095);
nor U29622 (N_29622,N_29206,N_29403);
and U29623 (N_29623,N_29207,N_29215);
xor U29624 (N_29624,N_29132,N_29078);
nand U29625 (N_29625,N_29260,N_29153);
or U29626 (N_29626,N_29018,N_29445);
nor U29627 (N_29627,N_29238,N_29385);
or U29628 (N_29628,N_29140,N_29046);
xnor U29629 (N_29629,N_29181,N_29240);
xnor U29630 (N_29630,N_29160,N_29317);
nor U29631 (N_29631,N_29024,N_29336);
nor U29632 (N_29632,N_29400,N_29352);
nand U29633 (N_29633,N_29013,N_29131);
nand U29634 (N_29634,N_29346,N_29395);
nor U29635 (N_29635,N_29139,N_29159);
nand U29636 (N_29636,N_29040,N_29434);
and U29637 (N_29637,N_29236,N_29111);
nand U29638 (N_29638,N_29345,N_29106);
nand U29639 (N_29639,N_29415,N_29417);
or U29640 (N_29640,N_29053,N_29043);
xor U29641 (N_29641,N_29469,N_29493);
nand U29642 (N_29642,N_29461,N_29114);
or U29643 (N_29643,N_29453,N_29320);
nor U29644 (N_29644,N_29285,N_29011);
xor U29645 (N_29645,N_29148,N_29093);
and U29646 (N_29646,N_29147,N_29128);
or U29647 (N_29647,N_29127,N_29020);
xor U29648 (N_29648,N_29016,N_29382);
nor U29649 (N_29649,N_29123,N_29253);
and U29650 (N_29650,N_29196,N_29125);
or U29651 (N_29651,N_29329,N_29426);
and U29652 (N_29652,N_29432,N_29276);
nand U29653 (N_29653,N_29204,N_29209);
and U29654 (N_29654,N_29251,N_29325);
nor U29655 (N_29655,N_29064,N_29398);
nor U29656 (N_29656,N_29180,N_29375);
and U29657 (N_29657,N_29265,N_29305);
nor U29658 (N_29658,N_29335,N_29005);
and U29659 (N_29659,N_29248,N_29295);
nor U29660 (N_29660,N_29422,N_29243);
nand U29661 (N_29661,N_29174,N_29158);
nand U29662 (N_29662,N_29050,N_29157);
and U29663 (N_29663,N_29034,N_29312);
or U29664 (N_29664,N_29491,N_29366);
or U29665 (N_29665,N_29100,N_29130);
nand U29666 (N_29666,N_29252,N_29387);
nand U29667 (N_29667,N_29184,N_29273);
xor U29668 (N_29668,N_29104,N_29412);
xor U29669 (N_29669,N_29059,N_29301);
nor U29670 (N_29670,N_29091,N_29465);
xnor U29671 (N_29671,N_29425,N_29299);
xor U29672 (N_29672,N_29118,N_29116);
and U29673 (N_29673,N_29452,N_29288);
nand U29674 (N_29674,N_29001,N_29462);
nand U29675 (N_29675,N_29178,N_29143);
or U29676 (N_29676,N_29186,N_29155);
nor U29677 (N_29677,N_29216,N_29079);
and U29678 (N_29678,N_29176,N_29272);
nand U29679 (N_29679,N_29133,N_29035);
or U29680 (N_29680,N_29084,N_29073);
nand U29681 (N_29681,N_29383,N_29039);
and U29682 (N_29682,N_29292,N_29458);
nor U29683 (N_29683,N_29087,N_29350);
or U29684 (N_29684,N_29264,N_29115);
nand U29685 (N_29685,N_29235,N_29283);
or U29686 (N_29686,N_29239,N_29332);
and U29687 (N_29687,N_29149,N_29129);
xor U29688 (N_29688,N_29376,N_29051);
nor U29689 (N_29689,N_29391,N_29408);
and U29690 (N_29690,N_29074,N_29045);
nor U29691 (N_29691,N_29055,N_29321);
nand U29692 (N_29692,N_29364,N_29455);
nor U29693 (N_29693,N_29496,N_29102);
xnor U29694 (N_29694,N_29315,N_29089);
or U29695 (N_29695,N_29351,N_29429);
xnor U29696 (N_29696,N_29246,N_29284);
and U29697 (N_29697,N_29341,N_29460);
nand U29698 (N_29698,N_29062,N_29212);
nand U29699 (N_29699,N_29443,N_29413);
xnor U29700 (N_29700,N_29047,N_29006);
xnor U29701 (N_29701,N_29456,N_29255);
and U29702 (N_29702,N_29407,N_29339);
nand U29703 (N_29703,N_29004,N_29459);
nor U29704 (N_29704,N_29476,N_29471);
nor U29705 (N_29705,N_29261,N_29122);
nor U29706 (N_29706,N_29022,N_29449);
nand U29707 (N_29707,N_29169,N_29249);
and U29708 (N_29708,N_29411,N_29293);
and U29709 (N_29709,N_29349,N_29410);
xnor U29710 (N_29710,N_29145,N_29447);
or U29711 (N_29711,N_29164,N_29126);
and U29712 (N_29712,N_29217,N_29167);
xor U29713 (N_29713,N_29337,N_29365);
nor U29714 (N_29714,N_29220,N_29110);
and U29715 (N_29715,N_29103,N_29076);
nor U29716 (N_29716,N_29038,N_29166);
nand U29717 (N_29717,N_29269,N_29499);
nand U29718 (N_29718,N_29154,N_29437);
nor U29719 (N_29719,N_29495,N_29343);
and U29720 (N_29720,N_29187,N_29466);
nor U29721 (N_29721,N_29008,N_29021);
nand U29722 (N_29722,N_29393,N_29098);
and U29723 (N_29723,N_29226,N_29161);
and U29724 (N_29724,N_29406,N_29185);
and U29725 (N_29725,N_29136,N_29280);
or U29726 (N_29726,N_29041,N_29311);
xor U29727 (N_29727,N_29470,N_29190);
nand U29728 (N_29728,N_29497,N_29378);
xnor U29729 (N_29729,N_29049,N_29266);
and U29730 (N_29730,N_29175,N_29330);
and U29731 (N_29731,N_29007,N_29357);
nand U29732 (N_29732,N_29328,N_29390);
nor U29733 (N_29733,N_29085,N_29381);
nor U29734 (N_29734,N_29170,N_29066);
or U29735 (N_29735,N_29099,N_29228);
and U29736 (N_29736,N_29300,N_29316);
nor U29737 (N_29737,N_29309,N_29480);
nor U29738 (N_29738,N_29014,N_29359);
and U29739 (N_29739,N_29327,N_29409);
xor U29740 (N_29740,N_29489,N_29037);
xnor U29741 (N_29741,N_29023,N_29306);
or U29742 (N_29742,N_29479,N_29347);
nand U29743 (N_29743,N_29177,N_29323);
or U29744 (N_29744,N_29244,N_29061);
and U29745 (N_29745,N_29277,N_29241);
nor U29746 (N_29746,N_29109,N_29475);
or U29747 (N_29747,N_29254,N_29002);
xor U29748 (N_29748,N_29370,N_29121);
nor U29749 (N_29749,N_29310,N_29193);
or U29750 (N_29750,N_29069,N_29234);
and U29751 (N_29751,N_29330,N_29098);
or U29752 (N_29752,N_29027,N_29079);
and U29753 (N_29753,N_29416,N_29465);
nand U29754 (N_29754,N_29326,N_29105);
and U29755 (N_29755,N_29000,N_29372);
or U29756 (N_29756,N_29465,N_29003);
xnor U29757 (N_29757,N_29456,N_29153);
nor U29758 (N_29758,N_29282,N_29256);
nor U29759 (N_29759,N_29312,N_29276);
and U29760 (N_29760,N_29112,N_29062);
and U29761 (N_29761,N_29207,N_29030);
or U29762 (N_29762,N_29169,N_29143);
and U29763 (N_29763,N_29391,N_29476);
nand U29764 (N_29764,N_29149,N_29305);
and U29765 (N_29765,N_29125,N_29440);
nand U29766 (N_29766,N_29214,N_29221);
and U29767 (N_29767,N_29097,N_29450);
xor U29768 (N_29768,N_29125,N_29174);
xnor U29769 (N_29769,N_29329,N_29448);
xnor U29770 (N_29770,N_29427,N_29434);
or U29771 (N_29771,N_29012,N_29150);
nand U29772 (N_29772,N_29168,N_29489);
and U29773 (N_29773,N_29364,N_29203);
xnor U29774 (N_29774,N_29252,N_29204);
and U29775 (N_29775,N_29296,N_29481);
xor U29776 (N_29776,N_29320,N_29485);
or U29777 (N_29777,N_29468,N_29227);
or U29778 (N_29778,N_29420,N_29456);
or U29779 (N_29779,N_29013,N_29122);
and U29780 (N_29780,N_29429,N_29334);
nand U29781 (N_29781,N_29424,N_29003);
xnor U29782 (N_29782,N_29087,N_29262);
nor U29783 (N_29783,N_29363,N_29399);
and U29784 (N_29784,N_29187,N_29291);
nor U29785 (N_29785,N_29367,N_29320);
and U29786 (N_29786,N_29361,N_29376);
xor U29787 (N_29787,N_29320,N_29355);
and U29788 (N_29788,N_29362,N_29353);
nor U29789 (N_29789,N_29304,N_29204);
nand U29790 (N_29790,N_29085,N_29090);
nand U29791 (N_29791,N_29178,N_29261);
and U29792 (N_29792,N_29003,N_29353);
xnor U29793 (N_29793,N_29232,N_29333);
nor U29794 (N_29794,N_29437,N_29398);
nor U29795 (N_29795,N_29095,N_29228);
or U29796 (N_29796,N_29330,N_29256);
nor U29797 (N_29797,N_29453,N_29156);
or U29798 (N_29798,N_29371,N_29341);
nand U29799 (N_29799,N_29087,N_29146);
xnor U29800 (N_29800,N_29448,N_29304);
xnor U29801 (N_29801,N_29331,N_29325);
nand U29802 (N_29802,N_29045,N_29387);
and U29803 (N_29803,N_29245,N_29059);
xor U29804 (N_29804,N_29463,N_29263);
nor U29805 (N_29805,N_29061,N_29265);
xor U29806 (N_29806,N_29153,N_29078);
or U29807 (N_29807,N_29330,N_29250);
nor U29808 (N_29808,N_29295,N_29286);
and U29809 (N_29809,N_29493,N_29497);
nand U29810 (N_29810,N_29228,N_29385);
nand U29811 (N_29811,N_29092,N_29064);
and U29812 (N_29812,N_29186,N_29138);
nor U29813 (N_29813,N_29036,N_29371);
and U29814 (N_29814,N_29328,N_29036);
nand U29815 (N_29815,N_29078,N_29089);
xnor U29816 (N_29816,N_29390,N_29273);
and U29817 (N_29817,N_29258,N_29434);
and U29818 (N_29818,N_29486,N_29328);
nand U29819 (N_29819,N_29315,N_29008);
and U29820 (N_29820,N_29053,N_29070);
and U29821 (N_29821,N_29335,N_29180);
xnor U29822 (N_29822,N_29454,N_29295);
or U29823 (N_29823,N_29403,N_29400);
or U29824 (N_29824,N_29394,N_29252);
and U29825 (N_29825,N_29427,N_29460);
nor U29826 (N_29826,N_29001,N_29097);
or U29827 (N_29827,N_29266,N_29412);
nand U29828 (N_29828,N_29358,N_29488);
and U29829 (N_29829,N_29041,N_29117);
and U29830 (N_29830,N_29231,N_29477);
nand U29831 (N_29831,N_29194,N_29219);
xnor U29832 (N_29832,N_29304,N_29253);
or U29833 (N_29833,N_29020,N_29154);
nand U29834 (N_29834,N_29195,N_29451);
nand U29835 (N_29835,N_29439,N_29083);
nand U29836 (N_29836,N_29349,N_29054);
or U29837 (N_29837,N_29242,N_29373);
nand U29838 (N_29838,N_29333,N_29331);
nor U29839 (N_29839,N_29115,N_29364);
or U29840 (N_29840,N_29287,N_29220);
xor U29841 (N_29841,N_29124,N_29180);
nor U29842 (N_29842,N_29369,N_29300);
nand U29843 (N_29843,N_29049,N_29237);
or U29844 (N_29844,N_29121,N_29391);
nor U29845 (N_29845,N_29116,N_29306);
or U29846 (N_29846,N_29068,N_29393);
or U29847 (N_29847,N_29469,N_29417);
nor U29848 (N_29848,N_29325,N_29459);
xor U29849 (N_29849,N_29178,N_29277);
nand U29850 (N_29850,N_29435,N_29457);
xor U29851 (N_29851,N_29004,N_29032);
nor U29852 (N_29852,N_29253,N_29217);
and U29853 (N_29853,N_29308,N_29331);
and U29854 (N_29854,N_29250,N_29276);
nor U29855 (N_29855,N_29391,N_29154);
xor U29856 (N_29856,N_29091,N_29437);
or U29857 (N_29857,N_29412,N_29398);
and U29858 (N_29858,N_29394,N_29174);
or U29859 (N_29859,N_29267,N_29404);
nand U29860 (N_29860,N_29242,N_29177);
or U29861 (N_29861,N_29137,N_29049);
nor U29862 (N_29862,N_29161,N_29304);
xor U29863 (N_29863,N_29460,N_29432);
and U29864 (N_29864,N_29434,N_29055);
xor U29865 (N_29865,N_29221,N_29343);
and U29866 (N_29866,N_29196,N_29129);
or U29867 (N_29867,N_29039,N_29331);
nor U29868 (N_29868,N_29110,N_29319);
and U29869 (N_29869,N_29101,N_29041);
or U29870 (N_29870,N_29231,N_29315);
and U29871 (N_29871,N_29212,N_29288);
nor U29872 (N_29872,N_29408,N_29319);
and U29873 (N_29873,N_29315,N_29103);
or U29874 (N_29874,N_29249,N_29333);
nor U29875 (N_29875,N_29110,N_29312);
xnor U29876 (N_29876,N_29404,N_29036);
xnor U29877 (N_29877,N_29377,N_29191);
or U29878 (N_29878,N_29429,N_29388);
or U29879 (N_29879,N_29344,N_29348);
nand U29880 (N_29880,N_29218,N_29193);
and U29881 (N_29881,N_29164,N_29137);
and U29882 (N_29882,N_29159,N_29164);
and U29883 (N_29883,N_29441,N_29409);
and U29884 (N_29884,N_29047,N_29255);
or U29885 (N_29885,N_29435,N_29028);
xor U29886 (N_29886,N_29456,N_29046);
nand U29887 (N_29887,N_29318,N_29335);
xnor U29888 (N_29888,N_29415,N_29308);
or U29889 (N_29889,N_29034,N_29041);
nand U29890 (N_29890,N_29456,N_29468);
nor U29891 (N_29891,N_29206,N_29335);
xor U29892 (N_29892,N_29190,N_29053);
nor U29893 (N_29893,N_29186,N_29432);
and U29894 (N_29894,N_29321,N_29265);
or U29895 (N_29895,N_29066,N_29487);
and U29896 (N_29896,N_29396,N_29144);
or U29897 (N_29897,N_29121,N_29337);
nor U29898 (N_29898,N_29303,N_29079);
and U29899 (N_29899,N_29269,N_29039);
xor U29900 (N_29900,N_29094,N_29288);
and U29901 (N_29901,N_29457,N_29247);
and U29902 (N_29902,N_29309,N_29151);
nand U29903 (N_29903,N_29116,N_29176);
and U29904 (N_29904,N_29273,N_29444);
nand U29905 (N_29905,N_29181,N_29182);
nor U29906 (N_29906,N_29232,N_29325);
nand U29907 (N_29907,N_29435,N_29254);
nor U29908 (N_29908,N_29112,N_29168);
and U29909 (N_29909,N_29280,N_29062);
and U29910 (N_29910,N_29286,N_29404);
or U29911 (N_29911,N_29124,N_29494);
nor U29912 (N_29912,N_29254,N_29222);
xnor U29913 (N_29913,N_29242,N_29107);
and U29914 (N_29914,N_29377,N_29448);
or U29915 (N_29915,N_29101,N_29392);
or U29916 (N_29916,N_29265,N_29239);
nand U29917 (N_29917,N_29394,N_29090);
or U29918 (N_29918,N_29138,N_29233);
nand U29919 (N_29919,N_29221,N_29059);
or U29920 (N_29920,N_29226,N_29315);
or U29921 (N_29921,N_29129,N_29246);
nand U29922 (N_29922,N_29309,N_29376);
nand U29923 (N_29923,N_29282,N_29111);
and U29924 (N_29924,N_29479,N_29116);
nand U29925 (N_29925,N_29067,N_29189);
nor U29926 (N_29926,N_29164,N_29011);
nor U29927 (N_29927,N_29134,N_29492);
nand U29928 (N_29928,N_29191,N_29455);
xnor U29929 (N_29929,N_29031,N_29471);
nor U29930 (N_29930,N_29212,N_29161);
xor U29931 (N_29931,N_29481,N_29108);
nand U29932 (N_29932,N_29072,N_29463);
and U29933 (N_29933,N_29090,N_29355);
nand U29934 (N_29934,N_29287,N_29462);
and U29935 (N_29935,N_29279,N_29317);
or U29936 (N_29936,N_29373,N_29202);
nor U29937 (N_29937,N_29310,N_29000);
or U29938 (N_29938,N_29419,N_29166);
and U29939 (N_29939,N_29054,N_29105);
xnor U29940 (N_29940,N_29281,N_29454);
xor U29941 (N_29941,N_29085,N_29418);
and U29942 (N_29942,N_29310,N_29041);
xnor U29943 (N_29943,N_29148,N_29197);
xor U29944 (N_29944,N_29122,N_29491);
nor U29945 (N_29945,N_29220,N_29362);
nand U29946 (N_29946,N_29160,N_29307);
and U29947 (N_29947,N_29036,N_29475);
nor U29948 (N_29948,N_29084,N_29145);
nand U29949 (N_29949,N_29289,N_29006);
and U29950 (N_29950,N_29303,N_29379);
or U29951 (N_29951,N_29109,N_29342);
nand U29952 (N_29952,N_29034,N_29264);
or U29953 (N_29953,N_29389,N_29233);
nand U29954 (N_29954,N_29283,N_29329);
or U29955 (N_29955,N_29415,N_29149);
nor U29956 (N_29956,N_29389,N_29432);
nand U29957 (N_29957,N_29288,N_29254);
nor U29958 (N_29958,N_29169,N_29429);
nand U29959 (N_29959,N_29134,N_29451);
nor U29960 (N_29960,N_29164,N_29278);
nand U29961 (N_29961,N_29021,N_29172);
nor U29962 (N_29962,N_29370,N_29468);
nor U29963 (N_29963,N_29166,N_29345);
nand U29964 (N_29964,N_29430,N_29069);
nand U29965 (N_29965,N_29391,N_29245);
and U29966 (N_29966,N_29349,N_29172);
nand U29967 (N_29967,N_29486,N_29370);
xor U29968 (N_29968,N_29281,N_29351);
nor U29969 (N_29969,N_29161,N_29224);
and U29970 (N_29970,N_29273,N_29309);
or U29971 (N_29971,N_29246,N_29132);
and U29972 (N_29972,N_29065,N_29222);
nand U29973 (N_29973,N_29214,N_29158);
nor U29974 (N_29974,N_29260,N_29005);
or U29975 (N_29975,N_29106,N_29242);
nand U29976 (N_29976,N_29439,N_29400);
nand U29977 (N_29977,N_29275,N_29182);
nand U29978 (N_29978,N_29164,N_29160);
nand U29979 (N_29979,N_29347,N_29460);
and U29980 (N_29980,N_29351,N_29448);
nand U29981 (N_29981,N_29086,N_29199);
xor U29982 (N_29982,N_29470,N_29142);
nand U29983 (N_29983,N_29279,N_29267);
and U29984 (N_29984,N_29079,N_29129);
and U29985 (N_29985,N_29024,N_29184);
nand U29986 (N_29986,N_29164,N_29452);
and U29987 (N_29987,N_29276,N_29090);
or U29988 (N_29988,N_29319,N_29145);
nand U29989 (N_29989,N_29111,N_29160);
nor U29990 (N_29990,N_29204,N_29031);
xnor U29991 (N_29991,N_29090,N_29140);
or U29992 (N_29992,N_29118,N_29483);
xnor U29993 (N_29993,N_29029,N_29127);
xnor U29994 (N_29994,N_29376,N_29294);
and U29995 (N_29995,N_29040,N_29356);
and U29996 (N_29996,N_29340,N_29006);
xor U29997 (N_29997,N_29034,N_29230);
nor U29998 (N_29998,N_29019,N_29157);
xnor U29999 (N_29999,N_29306,N_29225);
xnor UO_0 (O_0,N_29932,N_29705);
nor UO_1 (O_1,N_29970,N_29506);
nor UO_2 (O_2,N_29575,N_29867);
nor UO_3 (O_3,N_29863,N_29826);
nand UO_4 (O_4,N_29942,N_29812);
nor UO_5 (O_5,N_29721,N_29740);
and UO_6 (O_6,N_29821,N_29846);
nand UO_7 (O_7,N_29832,N_29901);
nand UO_8 (O_8,N_29574,N_29703);
and UO_9 (O_9,N_29912,N_29982);
nand UO_10 (O_10,N_29845,N_29893);
nor UO_11 (O_11,N_29690,N_29682);
or UO_12 (O_12,N_29570,N_29508);
nand UO_13 (O_13,N_29672,N_29510);
and UO_14 (O_14,N_29803,N_29828);
and UO_15 (O_15,N_29852,N_29977);
or UO_16 (O_16,N_29971,N_29567);
and UO_17 (O_17,N_29525,N_29786);
and UO_18 (O_18,N_29702,N_29571);
or UO_19 (O_19,N_29637,N_29896);
and UO_20 (O_20,N_29814,N_29646);
nor UO_21 (O_21,N_29903,N_29511);
nand UO_22 (O_22,N_29605,N_29669);
nor UO_23 (O_23,N_29757,N_29984);
nor UO_24 (O_24,N_29923,N_29878);
nor UO_25 (O_25,N_29630,N_29884);
nor UO_26 (O_26,N_29798,N_29710);
nor UO_27 (O_27,N_29563,N_29865);
nor UO_28 (O_28,N_29524,N_29914);
nand UO_29 (O_29,N_29502,N_29781);
and UO_30 (O_30,N_29770,N_29976);
or UO_31 (O_31,N_29911,N_29775);
and UO_32 (O_32,N_29674,N_29691);
or UO_33 (O_33,N_29737,N_29905);
nand UO_34 (O_34,N_29625,N_29517);
xnor UO_35 (O_35,N_29644,N_29577);
xnor UO_36 (O_36,N_29875,N_29583);
nor UO_37 (O_37,N_29729,N_29862);
nor UO_38 (O_38,N_29604,N_29993);
xor UO_39 (O_39,N_29808,N_29592);
or UO_40 (O_40,N_29753,N_29928);
or UO_41 (O_41,N_29504,N_29505);
nor UO_42 (O_42,N_29613,N_29732);
nor UO_43 (O_43,N_29658,N_29758);
nand UO_44 (O_44,N_29934,N_29909);
or UO_45 (O_45,N_29980,N_29784);
xnor UO_46 (O_46,N_29938,N_29586);
nand UO_47 (O_47,N_29981,N_29759);
or UO_48 (O_48,N_29544,N_29565);
nand UO_49 (O_49,N_29589,N_29667);
xor UO_50 (O_50,N_29720,N_29995);
or UO_51 (O_51,N_29949,N_29871);
xor UO_52 (O_52,N_29787,N_29869);
xnor UO_53 (O_53,N_29628,N_29924);
and UO_54 (O_54,N_29783,N_29640);
nand UO_55 (O_55,N_29701,N_29853);
nor UO_56 (O_56,N_29666,N_29848);
or UO_57 (O_57,N_29904,N_29989);
or UO_58 (O_58,N_29700,N_29620);
xor UO_59 (O_59,N_29925,N_29802);
and UO_60 (O_60,N_29888,N_29872);
nand UO_61 (O_61,N_29807,N_29632);
xnor UO_62 (O_62,N_29673,N_29996);
and UO_63 (O_63,N_29838,N_29785);
xor UO_64 (O_64,N_29773,N_29696);
xor UO_65 (O_65,N_29503,N_29941);
xnor UO_66 (O_66,N_29687,N_29739);
nand UO_67 (O_67,N_29889,N_29816);
nand UO_68 (O_68,N_29727,N_29873);
xnor UO_69 (O_69,N_29734,N_29522);
xor UO_70 (O_70,N_29974,N_29627);
nand UO_71 (O_71,N_29708,N_29817);
xor UO_72 (O_72,N_29518,N_29582);
nor UO_73 (O_73,N_29623,N_29764);
nand UO_74 (O_74,N_29736,N_29801);
nor UO_75 (O_75,N_29972,N_29684);
or UO_76 (O_76,N_29731,N_29986);
nand UO_77 (O_77,N_29779,N_29656);
and UO_78 (O_78,N_29899,N_29835);
xor UO_79 (O_79,N_29957,N_29561);
or UO_80 (O_80,N_29868,N_29842);
xnor UO_81 (O_81,N_29854,N_29813);
xor UO_82 (O_82,N_29594,N_29839);
nor UO_83 (O_83,N_29650,N_29664);
or UO_84 (O_84,N_29545,N_29891);
or UO_85 (O_85,N_29857,N_29782);
xnor UO_86 (O_86,N_29730,N_29678);
and UO_87 (O_87,N_29654,N_29626);
nand UO_88 (O_88,N_29738,N_29573);
xnor UO_89 (O_89,N_29704,N_29535);
and UO_90 (O_90,N_29966,N_29537);
or UO_91 (O_91,N_29799,N_29973);
or UO_92 (O_92,N_29892,N_29841);
nor UO_93 (O_93,N_29723,N_29692);
or UO_94 (O_94,N_29983,N_29937);
or UO_95 (O_95,N_29992,N_29500);
nand UO_96 (O_96,N_29509,N_29595);
or UO_97 (O_97,N_29921,N_29564);
or UO_98 (O_98,N_29890,N_29861);
xor UO_99 (O_99,N_29608,N_29772);
or UO_100 (O_100,N_29760,N_29615);
nor UO_101 (O_101,N_29952,N_29856);
nor UO_102 (O_102,N_29755,N_29585);
xnor UO_103 (O_103,N_29748,N_29943);
xnor UO_104 (O_104,N_29831,N_29750);
nand UO_105 (O_105,N_29709,N_29979);
or UO_106 (O_106,N_29836,N_29512);
nand UO_107 (O_107,N_29515,N_29693);
nand UO_108 (O_108,N_29685,N_29935);
and UO_109 (O_109,N_29645,N_29761);
nor UO_110 (O_110,N_29947,N_29699);
or UO_111 (O_111,N_29745,N_29636);
xnor UO_112 (O_112,N_29552,N_29797);
nand UO_113 (O_113,N_29837,N_29774);
and UO_114 (O_114,N_29559,N_29806);
and UO_115 (O_115,N_29689,N_29603);
nand UO_116 (O_116,N_29825,N_29767);
nand UO_117 (O_117,N_29649,N_29560);
nand UO_118 (O_118,N_29777,N_29514);
or UO_119 (O_119,N_29572,N_29765);
nor UO_120 (O_120,N_29647,N_29600);
nor UO_121 (O_121,N_29717,N_29885);
xor UO_122 (O_122,N_29752,N_29675);
nor UO_123 (O_123,N_29791,N_29963);
or UO_124 (O_124,N_29551,N_29910);
xor UO_125 (O_125,N_29619,N_29988);
xnor UO_126 (O_126,N_29516,N_29990);
or UO_127 (O_127,N_29541,N_29881);
or UO_128 (O_128,N_29733,N_29612);
or UO_129 (O_129,N_29805,N_29631);
xor UO_130 (O_130,N_29746,N_29556);
and UO_131 (O_131,N_29766,N_29829);
nor UO_132 (O_132,N_29707,N_29991);
nor UO_133 (O_133,N_29558,N_29665);
nand UO_134 (O_134,N_29531,N_29719);
or UO_135 (O_135,N_29610,N_29822);
nor UO_136 (O_136,N_29827,N_29617);
xnor UO_137 (O_137,N_29538,N_29576);
nand UO_138 (O_138,N_29894,N_29820);
nor UO_139 (O_139,N_29819,N_29680);
xor UO_140 (O_140,N_29792,N_29520);
or UO_141 (O_141,N_29599,N_29960);
nor UO_142 (O_142,N_29578,N_29621);
and UO_143 (O_143,N_29780,N_29507);
nor UO_144 (O_144,N_29931,N_29953);
xnor UO_145 (O_145,N_29994,N_29542);
nand UO_146 (O_146,N_29554,N_29501);
or UO_147 (O_147,N_29533,N_29796);
or UO_148 (O_148,N_29718,N_29858);
and UO_149 (O_149,N_29969,N_29744);
nor UO_150 (O_150,N_29956,N_29587);
and UO_151 (O_151,N_29895,N_29849);
xnor UO_152 (O_152,N_29724,N_29553);
nor UO_153 (O_153,N_29855,N_29639);
xnor UO_154 (O_154,N_29769,N_29951);
or UO_155 (O_155,N_29959,N_29548);
xnor UO_156 (O_156,N_29523,N_29534);
xnor UO_157 (O_157,N_29530,N_29778);
nand UO_158 (O_158,N_29810,N_29987);
nor UO_159 (O_159,N_29555,N_29795);
xor UO_160 (O_160,N_29940,N_29920);
xor UO_161 (O_161,N_29898,N_29527);
or UO_162 (O_162,N_29859,N_29683);
or UO_163 (O_163,N_29638,N_29844);
or UO_164 (O_164,N_29681,N_29958);
and UO_165 (O_165,N_29790,N_29866);
nor UO_166 (O_166,N_29579,N_29876);
nor UO_167 (O_167,N_29539,N_29540);
nand UO_168 (O_168,N_29962,N_29741);
nor UO_169 (O_169,N_29686,N_29804);
or UO_170 (O_170,N_29754,N_29728);
xnor UO_171 (O_171,N_29602,N_29726);
xnor UO_172 (O_172,N_29800,N_29624);
nand UO_173 (O_173,N_29950,N_29616);
or UO_174 (O_174,N_29908,N_29823);
nor UO_175 (O_175,N_29663,N_29715);
nand UO_176 (O_176,N_29590,N_29771);
xor UO_177 (O_177,N_29526,N_29581);
nand UO_178 (O_178,N_29874,N_29546);
xnor UO_179 (O_179,N_29776,N_29999);
xnor UO_180 (O_180,N_29913,N_29713);
and UO_181 (O_181,N_29641,N_29864);
and UO_182 (O_182,N_29840,N_29834);
nor UO_183 (O_183,N_29851,N_29955);
or UO_184 (O_184,N_29648,N_29521);
or UO_185 (O_185,N_29618,N_29860);
xor UO_186 (O_186,N_29850,N_29998);
and UO_187 (O_187,N_29601,N_29706);
xnor UO_188 (O_188,N_29788,N_29697);
nand UO_189 (O_189,N_29670,N_29643);
or UO_190 (O_190,N_29830,N_29939);
xnor UO_191 (O_191,N_29883,N_29562);
nor UO_192 (O_192,N_29879,N_29622);
nand UO_193 (O_193,N_29967,N_29927);
nand UO_194 (O_194,N_29597,N_29662);
nor UO_195 (O_195,N_29659,N_29596);
xor UO_196 (O_196,N_29917,N_29657);
or UO_197 (O_197,N_29532,N_29762);
nor UO_198 (O_198,N_29711,N_29965);
xnor UO_199 (O_199,N_29824,N_29930);
xnor UO_200 (O_200,N_29847,N_29529);
nand UO_201 (O_201,N_29743,N_29653);
and UO_202 (O_202,N_29818,N_29886);
nand UO_203 (O_203,N_29789,N_29676);
xor UO_204 (O_204,N_29968,N_29900);
xnor UO_205 (O_205,N_29714,N_29929);
and UO_206 (O_206,N_29936,N_29964);
or UO_207 (O_207,N_29588,N_29611);
or UO_208 (O_208,N_29528,N_29997);
nor UO_209 (O_209,N_29661,N_29742);
or UO_210 (O_210,N_29749,N_29882);
nand UO_211 (O_211,N_29961,N_29897);
nor UO_212 (O_212,N_29815,N_29671);
and UO_213 (O_213,N_29668,N_29652);
nor UO_214 (O_214,N_29591,N_29747);
nor UO_215 (O_215,N_29688,N_29598);
nor UO_216 (O_216,N_29580,N_29975);
xnor UO_217 (O_217,N_29954,N_29919);
nor UO_218 (O_218,N_29593,N_29695);
and UO_219 (O_219,N_29584,N_29763);
xor UO_220 (O_220,N_29651,N_29906);
and UO_221 (O_221,N_29547,N_29922);
or UO_222 (O_222,N_29811,N_29569);
nand UO_223 (O_223,N_29557,N_29660);
xnor UO_224 (O_224,N_29698,N_29519);
nand UO_225 (O_225,N_29809,N_29606);
nand UO_226 (O_226,N_29933,N_29833);
nor UO_227 (O_227,N_29550,N_29751);
or UO_228 (O_228,N_29712,N_29566);
nand UO_229 (O_229,N_29543,N_29642);
and UO_230 (O_230,N_29679,N_29725);
or UO_231 (O_231,N_29677,N_29549);
nand UO_232 (O_232,N_29629,N_29536);
and UO_233 (O_233,N_29945,N_29694);
nand UO_234 (O_234,N_29633,N_29607);
nand UO_235 (O_235,N_29634,N_29985);
xor UO_236 (O_236,N_29944,N_29614);
or UO_237 (O_237,N_29880,N_29568);
or UO_238 (O_238,N_29843,N_29609);
nand UO_239 (O_239,N_29735,N_29635);
nand UO_240 (O_240,N_29916,N_29948);
and UO_241 (O_241,N_29946,N_29978);
nand UO_242 (O_242,N_29902,N_29918);
nand UO_243 (O_243,N_29907,N_29513);
and UO_244 (O_244,N_29716,N_29877);
and UO_245 (O_245,N_29768,N_29655);
or UO_246 (O_246,N_29870,N_29915);
nand UO_247 (O_247,N_29722,N_29926);
or UO_248 (O_248,N_29756,N_29793);
nand UO_249 (O_249,N_29887,N_29794);
nor UO_250 (O_250,N_29851,N_29515);
and UO_251 (O_251,N_29884,N_29964);
xnor UO_252 (O_252,N_29689,N_29841);
xnor UO_253 (O_253,N_29600,N_29814);
nand UO_254 (O_254,N_29676,N_29924);
and UO_255 (O_255,N_29647,N_29636);
or UO_256 (O_256,N_29756,N_29700);
xnor UO_257 (O_257,N_29752,N_29798);
or UO_258 (O_258,N_29501,N_29675);
or UO_259 (O_259,N_29787,N_29638);
xnor UO_260 (O_260,N_29785,N_29766);
or UO_261 (O_261,N_29975,N_29705);
and UO_262 (O_262,N_29761,N_29850);
nor UO_263 (O_263,N_29968,N_29508);
and UO_264 (O_264,N_29854,N_29857);
xnor UO_265 (O_265,N_29898,N_29946);
xnor UO_266 (O_266,N_29619,N_29821);
or UO_267 (O_267,N_29711,N_29875);
and UO_268 (O_268,N_29520,N_29645);
nor UO_269 (O_269,N_29776,N_29612);
nand UO_270 (O_270,N_29928,N_29522);
and UO_271 (O_271,N_29683,N_29622);
nand UO_272 (O_272,N_29714,N_29501);
nand UO_273 (O_273,N_29969,N_29663);
nand UO_274 (O_274,N_29610,N_29750);
xnor UO_275 (O_275,N_29586,N_29983);
or UO_276 (O_276,N_29595,N_29825);
xor UO_277 (O_277,N_29550,N_29988);
xor UO_278 (O_278,N_29526,N_29557);
xnor UO_279 (O_279,N_29532,N_29998);
nor UO_280 (O_280,N_29950,N_29844);
xnor UO_281 (O_281,N_29944,N_29900);
and UO_282 (O_282,N_29595,N_29672);
or UO_283 (O_283,N_29925,N_29866);
and UO_284 (O_284,N_29924,N_29795);
xnor UO_285 (O_285,N_29758,N_29849);
nand UO_286 (O_286,N_29850,N_29557);
and UO_287 (O_287,N_29845,N_29613);
or UO_288 (O_288,N_29794,N_29771);
or UO_289 (O_289,N_29730,N_29875);
nand UO_290 (O_290,N_29636,N_29583);
and UO_291 (O_291,N_29919,N_29753);
xor UO_292 (O_292,N_29668,N_29835);
nand UO_293 (O_293,N_29548,N_29843);
nand UO_294 (O_294,N_29843,N_29641);
and UO_295 (O_295,N_29988,N_29561);
and UO_296 (O_296,N_29951,N_29587);
nor UO_297 (O_297,N_29853,N_29650);
nand UO_298 (O_298,N_29768,N_29963);
or UO_299 (O_299,N_29746,N_29840);
nand UO_300 (O_300,N_29658,N_29862);
nor UO_301 (O_301,N_29513,N_29567);
nand UO_302 (O_302,N_29783,N_29539);
nand UO_303 (O_303,N_29819,N_29755);
xor UO_304 (O_304,N_29678,N_29945);
and UO_305 (O_305,N_29916,N_29821);
and UO_306 (O_306,N_29722,N_29699);
nor UO_307 (O_307,N_29762,N_29810);
nand UO_308 (O_308,N_29922,N_29500);
nand UO_309 (O_309,N_29902,N_29670);
or UO_310 (O_310,N_29811,N_29544);
xor UO_311 (O_311,N_29562,N_29856);
or UO_312 (O_312,N_29713,N_29653);
or UO_313 (O_313,N_29889,N_29619);
xor UO_314 (O_314,N_29528,N_29794);
and UO_315 (O_315,N_29811,N_29918);
and UO_316 (O_316,N_29991,N_29592);
xnor UO_317 (O_317,N_29522,N_29636);
nor UO_318 (O_318,N_29821,N_29987);
nand UO_319 (O_319,N_29584,N_29772);
xnor UO_320 (O_320,N_29627,N_29717);
nand UO_321 (O_321,N_29769,N_29581);
xor UO_322 (O_322,N_29768,N_29714);
nor UO_323 (O_323,N_29683,N_29774);
or UO_324 (O_324,N_29983,N_29603);
or UO_325 (O_325,N_29551,N_29862);
nor UO_326 (O_326,N_29562,N_29626);
and UO_327 (O_327,N_29875,N_29772);
xor UO_328 (O_328,N_29696,N_29863);
nor UO_329 (O_329,N_29729,N_29993);
or UO_330 (O_330,N_29529,N_29536);
and UO_331 (O_331,N_29841,N_29823);
nand UO_332 (O_332,N_29782,N_29607);
nor UO_333 (O_333,N_29769,N_29630);
nor UO_334 (O_334,N_29932,N_29546);
xor UO_335 (O_335,N_29820,N_29991);
and UO_336 (O_336,N_29572,N_29630);
nand UO_337 (O_337,N_29623,N_29663);
or UO_338 (O_338,N_29729,N_29713);
or UO_339 (O_339,N_29952,N_29683);
nor UO_340 (O_340,N_29950,N_29955);
nor UO_341 (O_341,N_29695,N_29969);
xor UO_342 (O_342,N_29783,N_29895);
nor UO_343 (O_343,N_29684,N_29903);
or UO_344 (O_344,N_29638,N_29654);
nand UO_345 (O_345,N_29711,N_29557);
xnor UO_346 (O_346,N_29606,N_29897);
or UO_347 (O_347,N_29883,N_29501);
nand UO_348 (O_348,N_29656,N_29746);
xor UO_349 (O_349,N_29608,N_29834);
nor UO_350 (O_350,N_29855,N_29746);
xor UO_351 (O_351,N_29509,N_29961);
or UO_352 (O_352,N_29730,N_29889);
xnor UO_353 (O_353,N_29940,N_29915);
xnor UO_354 (O_354,N_29886,N_29637);
xnor UO_355 (O_355,N_29954,N_29692);
nor UO_356 (O_356,N_29937,N_29697);
or UO_357 (O_357,N_29798,N_29864);
or UO_358 (O_358,N_29861,N_29745);
nand UO_359 (O_359,N_29831,N_29505);
nor UO_360 (O_360,N_29533,N_29737);
nor UO_361 (O_361,N_29632,N_29846);
xnor UO_362 (O_362,N_29974,N_29948);
xor UO_363 (O_363,N_29912,N_29796);
xor UO_364 (O_364,N_29780,N_29557);
xnor UO_365 (O_365,N_29985,N_29940);
or UO_366 (O_366,N_29902,N_29925);
or UO_367 (O_367,N_29857,N_29547);
nand UO_368 (O_368,N_29989,N_29578);
xor UO_369 (O_369,N_29914,N_29994);
or UO_370 (O_370,N_29724,N_29969);
nand UO_371 (O_371,N_29849,N_29930);
nor UO_372 (O_372,N_29841,N_29995);
or UO_373 (O_373,N_29677,N_29868);
nand UO_374 (O_374,N_29867,N_29921);
nor UO_375 (O_375,N_29813,N_29865);
xor UO_376 (O_376,N_29691,N_29745);
and UO_377 (O_377,N_29722,N_29965);
xor UO_378 (O_378,N_29673,N_29777);
xor UO_379 (O_379,N_29509,N_29747);
and UO_380 (O_380,N_29509,N_29536);
nor UO_381 (O_381,N_29541,N_29675);
xor UO_382 (O_382,N_29790,N_29676);
or UO_383 (O_383,N_29635,N_29731);
xnor UO_384 (O_384,N_29854,N_29960);
nor UO_385 (O_385,N_29716,N_29802);
nor UO_386 (O_386,N_29658,N_29937);
and UO_387 (O_387,N_29738,N_29591);
nand UO_388 (O_388,N_29954,N_29991);
xor UO_389 (O_389,N_29604,N_29508);
nand UO_390 (O_390,N_29616,N_29970);
or UO_391 (O_391,N_29541,N_29606);
or UO_392 (O_392,N_29543,N_29564);
nand UO_393 (O_393,N_29779,N_29616);
and UO_394 (O_394,N_29924,N_29578);
nor UO_395 (O_395,N_29898,N_29883);
or UO_396 (O_396,N_29510,N_29902);
nand UO_397 (O_397,N_29611,N_29632);
nor UO_398 (O_398,N_29699,N_29771);
nor UO_399 (O_399,N_29626,N_29805);
xnor UO_400 (O_400,N_29707,N_29592);
nor UO_401 (O_401,N_29976,N_29767);
nand UO_402 (O_402,N_29934,N_29891);
and UO_403 (O_403,N_29641,N_29946);
and UO_404 (O_404,N_29895,N_29997);
xnor UO_405 (O_405,N_29749,N_29843);
nor UO_406 (O_406,N_29533,N_29620);
or UO_407 (O_407,N_29551,N_29613);
nand UO_408 (O_408,N_29585,N_29633);
xnor UO_409 (O_409,N_29639,N_29665);
xnor UO_410 (O_410,N_29861,N_29958);
or UO_411 (O_411,N_29691,N_29751);
xnor UO_412 (O_412,N_29966,N_29690);
xor UO_413 (O_413,N_29580,N_29794);
xnor UO_414 (O_414,N_29867,N_29591);
or UO_415 (O_415,N_29738,N_29843);
and UO_416 (O_416,N_29825,N_29964);
xor UO_417 (O_417,N_29736,N_29733);
nand UO_418 (O_418,N_29788,N_29877);
nand UO_419 (O_419,N_29952,N_29741);
and UO_420 (O_420,N_29877,N_29685);
xor UO_421 (O_421,N_29688,N_29654);
nor UO_422 (O_422,N_29809,N_29575);
or UO_423 (O_423,N_29943,N_29843);
nand UO_424 (O_424,N_29841,N_29777);
nand UO_425 (O_425,N_29753,N_29892);
nor UO_426 (O_426,N_29977,N_29733);
and UO_427 (O_427,N_29605,N_29563);
or UO_428 (O_428,N_29878,N_29987);
nor UO_429 (O_429,N_29819,N_29603);
nor UO_430 (O_430,N_29997,N_29530);
nor UO_431 (O_431,N_29606,N_29969);
and UO_432 (O_432,N_29600,N_29861);
nand UO_433 (O_433,N_29632,N_29564);
nor UO_434 (O_434,N_29894,N_29582);
xor UO_435 (O_435,N_29500,N_29561);
and UO_436 (O_436,N_29709,N_29667);
nor UO_437 (O_437,N_29760,N_29713);
nand UO_438 (O_438,N_29612,N_29754);
nor UO_439 (O_439,N_29601,N_29625);
xor UO_440 (O_440,N_29870,N_29863);
and UO_441 (O_441,N_29725,N_29604);
or UO_442 (O_442,N_29533,N_29703);
and UO_443 (O_443,N_29569,N_29788);
or UO_444 (O_444,N_29696,N_29654);
or UO_445 (O_445,N_29597,N_29637);
xnor UO_446 (O_446,N_29817,N_29733);
nand UO_447 (O_447,N_29767,N_29736);
and UO_448 (O_448,N_29556,N_29588);
nor UO_449 (O_449,N_29761,N_29606);
nor UO_450 (O_450,N_29987,N_29658);
or UO_451 (O_451,N_29818,N_29797);
and UO_452 (O_452,N_29823,N_29583);
nand UO_453 (O_453,N_29702,N_29749);
and UO_454 (O_454,N_29879,N_29991);
nand UO_455 (O_455,N_29552,N_29913);
nand UO_456 (O_456,N_29683,N_29577);
and UO_457 (O_457,N_29859,N_29879);
nor UO_458 (O_458,N_29913,N_29607);
nand UO_459 (O_459,N_29966,N_29923);
nor UO_460 (O_460,N_29595,N_29706);
and UO_461 (O_461,N_29504,N_29542);
or UO_462 (O_462,N_29623,N_29862);
xnor UO_463 (O_463,N_29971,N_29961);
and UO_464 (O_464,N_29844,N_29900);
nor UO_465 (O_465,N_29953,N_29528);
nand UO_466 (O_466,N_29794,N_29520);
and UO_467 (O_467,N_29601,N_29700);
nand UO_468 (O_468,N_29559,N_29708);
nor UO_469 (O_469,N_29890,N_29707);
nor UO_470 (O_470,N_29796,N_29749);
and UO_471 (O_471,N_29989,N_29897);
xnor UO_472 (O_472,N_29827,N_29978);
or UO_473 (O_473,N_29632,N_29691);
nor UO_474 (O_474,N_29649,N_29662);
xnor UO_475 (O_475,N_29804,N_29634);
xor UO_476 (O_476,N_29645,N_29654);
and UO_477 (O_477,N_29650,N_29788);
nand UO_478 (O_478,N_29576,N_29755);
xnor UO_479 (O_479,N_29953,N_29752);
xnor UO_480 (O_480,N_29813,N_29664);
or UO_481 (O_481,N_29867,N_29530);
and UO_482 (O_482,N_29637,N_29861);
xor UO_483 (O_483,N_29720,N_29526);
nor UO_484 (O_484,N_29793,N_29620);
xnor UO_485 (O_485,N_29816,N_29844);
xnor UO_486 (O_486,N_29522,N_29555);
and UO_487 (O_487,N_29531,N_29561);
or UO_488 (O_488,N_29990,N_29757);
or UO_489 (O_489,N_29895,N_29787);
nor UO_490 (O_490,N_29933,N_29969);
xnor UO_491 (O_491,N_29880,N_29657);
and UO_492 (O_492,N_29681,N_29873);
xor UO_493 (O_493,N_29882,N_29993);
and UO_494 (O_494,N_29600,N_29984);
or UO_495 (O_495,N_29864,N_29718);
nand UO_496 (O_496,N_29856,N_29510);
nor UO_497 (O_497,N_29940,N_29583);
nor UO_498 (O_498,N_29723,N_29613);
and UO_499 (O_499,N_29631,N_29796);
or UO_500 (O_500,N_29681,N_29684);
nand UO_501 (O_501,N_29913,N_29722);
nor UO_502 (O_502,N_29700,N_29893);
xnor UO_503 (O_503,N_29843,N_29933);
and UO_504 (O_504,N_29663,N_29762);
or UO_505 (O_505,N_29705,N_29605);
or UO_506 (O_506,N_29849,N_29966);
and UO_507 (O_507,N_29524,N_29829);
and UO_508 (O_508,N_29737,N_29853);
and UO_509 (O_509,N_29598,N_29996);
nor UO_510 (O_510,N_29618,N_29956);
nor UO_511 (O_511,N_29607,N_29808);
or UO_512 (O_512,N_29715,N_29538);
xor UO_513 (O_513,N_29705,N_29730);
or UO_514 (O_514,N_29714,N_29736);
or UO_515 (O_515,N_29780,N_29632);
or UO_516 (O_516,N_29850,N_29665);
or UO_517 (O_517,N_29738,N_29678);
nand UO_518 (O_518,N_29518,N_29941);
and UO_519 (O_519,N_29747,N_29681);
or UO_520 (O_520,N_29640,N_29651);
or UO_521 (O_521,N_29770,N_29650);
nand UO_522 (O_522,N_29640,N_29535);
xor UO_523 (O_523,N_29765,N_29864);
and UO_524 (O_524,N_29769,N_29867);
nand UO_525 (O_525,N_29933,N_29759);
nand UO_526 (O_526,N_29702,N_29532);
or UO_527 (O_527,N_29827,N_29865);
nor UO_528 (O_528,N_29992,N_29625);
nor UO_529 (O_529,N_29552,N_29825);
and UO_530 (O_530,N_29636,N_29557);
or UO_531 (O_531,N_29956,N_29722);
nor UO_532 (O_532,N_29693,N_29573);
xor UO_533 (O_533,N_29799,N_29501);
or UO_534 (O_534,N_29555,N_29671);
or UO_535 (O_535,N_29777,N_29657);
or UO_536 (O_536,N_29967,N_29891);
xor UO_537 (O_537,N_29630,N_29703);
or UO_538 (O_538,N_29939,N_29606);
nand UO_539 (O_539,N_29869,N_29537);
and UO_540 (O_540,N_29774,N_29806);
and UO_541 (O_541,N_29799,N_29676);
nand UO_542 (O_542,N_29876,N_29885);
and UO_543 (O_543,N_29617,N_29971);
nor UO_544 (O_544,N_29797,N_29596);
xnor UO_545 (O_545,N_29609,N_29672);
or UO_546 (O_546,N_29679,N_29517);
or UO_547 (O_547,N_29523,N_29839);
and UO_548 (O_548,N_29631,N_29896);
or UO_549 (O_549,N_29780,N_29906);
or UO_550 (O_550,N_29583,N_29677);
or UO_551 (O_551,N_29949,N_29629);
or UO_552 (O_552,N_29717,N_29518);
xnor UO_553 (O_553,N_29764,N_29636);
xor UO_554 (O_554,N_29933,N_29886);
or UO_555 (O_555,N_29513,N_29730);
xnor UO_556 (O_556,N_29638,N_29588);
xor UO_557 (O_557,N_29741,N_29644);
nor UO_558 (O_558,N_29504,N_29868);
xor UO_559 (O_559,N_29913,N_29702);
nor UO_560 (O_560,N_29781,N_29930);
nand UO_561 (O_561,N_29504,N_29593);
or UO_562 (O_562,N_29792,N_29761);
nor UO_563 (O_563,N_29924,N_29871);
nor UO_564 (O_564,N_29677,N_29822);
xor UO_565 (O_565,N_29530,N_29503);
nor UO_566 (O_566,N_29812,N_29901);
xor UO_567 (O_567,N_29884,N_29500);
or UO_568 (O_568,N_29820,N_29739);
nand UO_569 (O_569,N_29774,N_29860);
nand UO_570 (O_570,N_29611,N_29663);
and UO_571 (O_571,N_29666,N_29811);
and UO_572 (O_572,N_29796,N_29614);
or UO_573 (O_573,N_29702,N_29706);
xor UO_574 (O_574,N_29728,N_29996);
and UO_575 (O_575,N_29504,N_29855);
and UO_576 (O_576,N_29923,N_29700);
xnor UO_577 (O_577,N_29794,N_29541);
nor UO_578 (O_578,N_29596,N_29556);
nor UO_579 (O_579,N_29798,N_29569);
or UO_580 (O_580,N_29590,N_29550);
xnor UO_581 (O_581,N_29818,N_29555);
or UO_582 (O_582,N_29951,N_29998);
xnor UO_583 (O_583,N_29773,N_29695);
nor UO_584 (O_584,N_29570,N_29579);
nand UO_585 (O_585,N_29824,N_29725);
and UO_586 (O_586,N_29533,N_29779);
xnor UO_587 (O_587,N_29662,N_29797);
xor UO_588 (O_588,N_29598,N_29505);
nand UO_589 (O_589,N_29791,N_29896);
and UO_590 (O_590,N_29632,N_29511);
nor UO_591 (O_591,N_29811,N_29770);
or UO_592 (O_592,N_29806,N_29540);
nand UO_593 (O_593,N_29559,N_29957);
or UO_594 (O_594,N_29595,N_29807);
and UO_595 (O_595,N_29800,N_29572);
and UO_596 (O_596,N_29958,N_29840);
or UO_597 (O_597,N_29534,N_29658);
nor UO_598 (O_598,N_29586,N_29554);
nand UO_599 (O_599,N_29822,N_29557);
or UO_600 (O_600,N_29712,N_29620);
nand UO_601 (O_601,N_29936,N_29621);
or UO_602 (O_602,N_29839,N_29807);
nand UO_603 (O_603,N_29891,N_29594);
nor UO_604 (O_604,N_29949,N_29966);
or UO_605 (O_605,N_29670,N_29755);
nand UO_606 (O_606,N_29814,N_29722);
and UO_607 (O_607,N_29650,N_29841);
nor UO_608 (O_608,N_29579,N_29948);
and UO_609 (O_609,N_29780,N_29813);
nor UO_610 (O_610,N_29895,N_29847);
nand UO_611 (O_611,N_29708,N_29584);
and UO_612 (O_612,N_29658,N_29860);
nor UO_613 (O_613,N_29852,N_29569);
or UO_614 (O_614,N_29836,N_29755);
nor UO_615 (O_615,N_29574,N_29613);
nand UO_616 (O_616,N_29678,N_29826);
or UO_617 (O_617,N_29613,N_29736);
nand UO_618 (O_618,N_29724,N_29676);
xnor UO_619 (O_619,N_29829,N_29595);
nand UO_620 (O_620,N_29641,N_29801);
or UO_621 (O_621,N_29777,N_29548);
and UO_622 (O_622,N_29770,N_29637);
nor UO_623 (O_623,N_29760,N_29793);
and UO_624 (O_624,N_29508,N_29865);
and UO_625 (O_625,N_29926,N_29584);
or UO_626 (O_626,N_29994,N_29507);
xnor UO_627 (O_627,N_29562,N_29833);
and UO_628 (O_628,N_29649,N_29882);
xnor UO_629 (O_629,N_29827,N_29818);
nand UO_630 (O_630,N_29642,N_29725);
or UO_631 (O_631,N_29648,N_29912);
and UO_632 (O_632,N_29787,N_29761);
nand UO_633 (O_633,N_29962,N_29676);
or UO_634 (O_634,N_29658,N_29749);
xor UO_635 (O_635,N_29776,N_29710);
and UO_636 (O_636,N_29723,N_29649);
nand UO_637 (O_637,N_29509,N_29766);
and UO_638 (O_638,N_29824,N_29786);
nand UO_639 (O_639,N_29922,N_29944);
nor UO_640 (O_640,N_29995,N_29711);
xor UO_641 (O_641,N_29592,N_29915);
nor UO_642 (O_642,N_29709,N_29553);
and UO_643 (O_643,N_29851,N_29601);
nor UO_644 (O_644,N_29700,N_29664);
nor UO_645 (O_645,N_29974,N_29872);
xor UO_646 (O_646,N_29584,N_29563);
and UO_647 (O_647,N_29828,N_29991);
nand UO_648 (O_648,N_29732,N_29654);
nor UO_649 (O_649,N_29776,N_29602);
nand UO_650 (O_650,N_29941,N_29556);
nand UO_651 (O_651,N_29600,N_29821);
xnor UO_652 (O_652,N_29817,N_29956);
nand UO_653 (O_653,N_29926,N_29677);
nand UO_654 (O_654,N_29648,N_29757);
and UO_655 (O_655,N_29934,N_29555);
xor UO_656 (O_656,N_29609,N_29719);
and UO_657 (O_657,N_29882,N_29699);
nand UO_658 (O_658,N_29804,N_29761);
xnor UO_659 (O_659,N_29682,N_29514);
and UO_660 (O_660,N_29894,N_29934);
nand UO_661 (O_661,N_29691,N_29547);
nand UO_662 (O_662,N_29934,N_29775);
xnor UO_663 (O_663,N_29649,N_29605);
nor UO_664 (O_664,N_29969,N_29554);
and UO_665 (O_665,N_29794,N_29602);
nand UO_666 (O_666,N_29567,N_29875);
xor UO_667 (O_667,N_29798,N_29652);
and UO_668 (O_668,N_29552,N_29724);
nor UO_669 (O_669,N_29789,N_29823);
or UO_670 (O_670,N_29717,N_29512);
nor UO_671 (O_671,N_29527,N_29859);
xnor UO_672 (O_672,N_29963,N_29891);
nor UO_673 (O_673,N_29560,N_29902);
nand UO_674 (O_674,N_29846,N_29925);
and UO_675 (O_675,N_29527,N_29931);
nor UO_676 (O_676,N_29781,N_29842);
or UO_677 (O_677,N_29702,N_29625);
and UO_678 (O_678,N_29873,N_29755);
or UO_679 (O_679,N_29714,N_29943);
nor UO_680 (O_680,N_29700,N_29881);
nor UO_681 (O_681,N_29973,N_29758);
or UO_682 (O_682,N_29772,N_29640);
nor UO_683 (O_683,N_29711,N_29595);
or UO_684 (O_684,N_29949,N_29722);
nor UO_685 (O_685,N_29546,N_29862);
or UO_686 (O_686,N_29918,N_29947);
xnor UO_687 (O_687,N_29519,N_29694);
nor UO_688 (O_688,N_29859,N_29684);
xnor UO_689 (O_689,N_29733,N_29667);
nand UO_690 (O_690,N_29899,N_29813);
and UO_691 (O_691,N_29940,N_29696);
or UO_692 (O_692,N_29703,N_29539);
or UO_693 (O_693,N_29607,N_29672);
or UO_694 (O_694,N_29648,N_29544);
xnor UO_695 (O_695,N_29990,N_29833);
nand UO_696 (O_696,N_29726,N_29648);
nand UO_697 (O_697,N_29720,N_29896);
nor UO_698 (O_698,N_29622,N_29931);
nand UO_699 (O_699,N_29632,N_29639);
nor UO_700 (O_700,N_29715,N_29898);
nand UO_701 (O_701,N_29921,N_29776);
and UO_702 (O_702,N_29816,N_29934);
xor UO_703 (O_703,N_29904,N_29851);
nand UO_704 (O_704,N_29620,N_29885);
or UO_705 (O_705,N_29948,N_29631);
nor UO_706 (O_706,N_29928,N_29965);
xor UO_707 (O_707,N_29919,N_29561);
and UO_708 (O_708,N_29510,N_29617);
and UO_709 (O_709,N_29673,N_29975);
nor UO_710 (O_710,N_29746,N_29771);
xnor UO_711 (O_711,N_29786,N_29501);
and UO_712 (O_712,N_29668,N_29627);
or UO_713 (O_713,N_29822,N_29618);
nor UO_714 (O_714,N_29994,N_29714);
nand UO_715 (O_715,N_29614,N_29740);
xor UO_716 (O_716,N_29767,N_29658);
xor UO_717 (O_717,N_29951,N_29881);
or UO_718 (O_718,N_29602,N_29814);
xnor UO_719 (O_719,N_29688,N_29962);
and UO_720 (O_720,N_29501,N_29906);
and UO_721 (O_721,N_29783,N_29501);
nand UO_722 (O_722,N_29866,N_29947);
nand UO_723 (O_723,N_29692,N_29732);
nand UO_724 (O_724,N_29570,N_29902);
xor UO_725 (O_725,N_29660,N_29864);
xnor UO_726 (O_726,N_29896,N_29794);
xnor UO_727 (O_727,N_29988,N_29834);
nor UO_728 (O_728,N_29781,N_29779);
or UO_729 (O_729,N_29875,N_29817);
nor UO_730 (O_730,N_29885,N_29968);
nor UO_731 (O_731,N_29976,N_29523);
and UO_732 (O_732,N_29838,N_29607);
or UO_733 (O_733,N_29736,N_29730);
and UO_734 (O_734,N_29513,N_29590);
nor UO_735 (O_735,N_29567,N_29821);
and UO_736 (O_736,N_29753,N_29817);
nand UO_737 (O_737,N_29897,N_29693);
nor UO_738 (O_738,N_29582,N_29770);
or UO_739 (O_739,N_29758,N_29643);
nand UO_740 (O_740,N_29883,N_29721);
nand UO_741 (O_741,N_29951,N_29916);
and UO_742 (O_742,N_29613,N_29905);
xor UO_743 (O_743,N_29532,N_29937);
nor UO_744 (O_744,N_29922,N_29948);
nand UO_745 (O_745,N_29739,N_29807);
or UO_746 (O_746,N_29763,N_29955);
xor UO_747 (O_747,N_29911,N_29622);
or UO_748 (O_748,N_29625,N_29736);
nor UO_749 (O_749,N_29744,N_29524);
and UO_750 (O_750,N_29897,N_29552);
xor UO_751 (O_751,N_29954,N_29850);
or UO_752 (O_752,N_29746,N_29530);
xnor UO_753 (O_753,N_29833,N_29724);
and UO_754 (O_754,N_29750,N_29729);
or UO_755 (O_755,N_29508,N_29846);
nor UO_756 (O_756,N_29750,N_29637);
nor UO_757 (O_757,N_29914,N_29553);
nor UO_758 (O_758,N_29708,N_29859);
xor UO_759 (O_759,N_29528,N_29523);
and UO_760 (O_760,N_29803,N_29664);
nor UO_761 (O_761,N_29932,N_29626);
and UO_762 (O_762,N_29928,N_29583);
nor UO_763 (O_763,N_29943,N_29619);
or UO_764 (O_764,N_29777,N_29551);
and UO_765 (O_765,N_29832,N_29891);
and UO_766 (O_766,N_29628,N_29584);
and UO_767 (O_767,N_29816,N_29590);
nor UO_768 (O_768,N_29559,N_29995);
nor UO_769 (O_769,N_29666,N_29614);
nand UO_770 (O_770,N_29848,N_29647);
nor UO_771 (O_771,N_29937,N_29757);
xor UO_772 (O_772,N_29627,N_29942);
and UO_773 (O_773,N_29525,N_29999);
nor UO_774 (O_774,N_29506,N_29961);
or UO_775 (O_775,N_29582,N_29973);
or UO_776 (O_776,N_29847,N_29860);
xnor UO_777 (O_777,N_29887,N_29762);
nand UO_778 (O_778,N_29959,N_29524);
and UO_779 (O_779,N_29708,N_29712);
and UO_780 (O_780,N_29527,N_29541);
nor UO_781 (O_781,N_29968,N_29659);
and UO_782 (O_782,N_29807,N_29940);
nand UO_783 (O_783,N_29610,N_29915);
or UO_784 (O_784,N_29649,N_29957);
nor UO_785 (O_785,N_29606,N_29951);
nand UO_786 (O_786,N_29574,N_29542);
nand UO_787 (O_787,N_29969,N_29975);
xnor UO_788 (O_788,N_29898,N_29508);
nor UO_789 (O_789,N_29536,N_29711);
nor UO_790 (O_790,N_29883,N_29609);
and UO_791 (O_791,N_29532,N_29693);
nor UO_792 (O_792,N_29915,N_29778);
nand UO_793 (O_793,N_29520,N_29899);
nor UO_794 (O_794,N_29727,N_29721);
and UO_795 (O_795,N_29928,N_29717);
nand UO_796 (O_796,N_29633,N_29587);
nor UO_797 (O_797,N_29601,N_29738);
or UO_798 (O_798,N_29718,N_29985);
or UO_799 (O_799,N_29962,N_29863);
or UO_800 (O_800,N_29811,N_29758);
nor UO_801 (O_801,N_29912,N_29664);
and UO_802 (O_802,N_29636,N_29575);
nand UO_803 (O_803,N_29961,N_29795);
and UO_804 (O_804,N_29823,N_29884);
or UO_805 (O_805,N_29960,N_29608);
xnor UO_806 (O_806,N_29650,N_29641);
or UO_807 (O_807,N_29550,N_29601);
and UO_808 (O_808,N_29538,N_29644);
nor UO_809 (O_809,N_29687,N_29571);
nor UO_810 (O_810,N_29679,N_29522);
or UO_811 (O_811,N_29715,N_29570);
nor UO_812 (O_812,N_29752,N_29983);
or UO_813 (O_813,N_29889,N_29650);
nor UO_814 (O_814,N_29859,N_29935);
xor UO_815 (O_815,N_29919,N_29928);
or UO_816 (O_816,N_29810,N_29516);
or UO_817 (O_817,N_29641,N_29510);
nor UO_818 (O_818,N_29778,N_29507);
or UO_819 (O_819,N_29696,N_29517);
and UO_820 (O_820,N_29969,N_29559);
xor UO_821 (O_821,N_29952,N_29796);
xor UO_822 (O_822,N_29750,N_29928);
nor UO_823 (O_823,N_29610,N_29964);
nand UO_824 (O_824,N_29505,N_29602);
xnor UO_825 (O_825,N_29582,N_29855);
xor UO_826 (O_826,N_29929,N_29903);
and UO_827 (O_827,N_29526,N_29667);
nor UO_828 (O_828,N_29943,N_29693);
and UO_829 (O_829,N_29869,N_29657);
or UO_830 (O_830,N_29894,N_29811);
xnor UO_831 (O_831,N_29508,N_29755);
nand UO_832 (O_832,N_29804,N_29682);
or UO_833 (O_833,N_29799,N_29597);
nand UO_834 (O_834,N_29691,N_29560);
and UO_835 (O_835,N_29557,N_29534);
nand UO_836 (O_836,N_29517,N_29971);
nor UO_837 (O_837,N_29757,N_29796);
nand UO_838 (O_838,N_29654,N_29618);
or UO_839 (O_839,N_29647,N_29728);
xor UO_840 (O_840,N_29656,N_29922);
nand UO_841 (O_841,N_29715,N_29810);
or UO_842 (O_842,N_29958,N_29993);
nor UO_843 (O_843,N_29769,N_29793);
nor UO_844 (O_844,N_29746,N_29707);
nor UO_845 (O_845,N_29627,N_29549);
or UO_846 (O_846,N_29782,N_29995);
xor UO_847 (O_847,N_29597,N_29764);
xnor UO_848 (O_848,N_29633,N_29805);
nor UO_849 (O_849,N_29816,N_29530);
xnor UO_850 (O_850,N_29856,N_29854);
and UO_851 (O_851,N_29672,N_29959);
nand UO_852 (O_852,N_29947,N_29713);
xnor UO_853 (O_853,N_29777,N_29659);
nor UO_854 (O_854,N_29522,N_29843);
xnor UO_855 (O_855,N_29754,N_29927);
and UO_856 (O_856,N_29815,N_29626);
nor UO_857 (O_857,N_29717,N_29742);
and UO_858 (O_858,N_29585,N_29649);
nand UO_859 (O_859,N_29945,N_29511);
xor UO_860 (O_860,N_29685,N_29648);
or UO_861 (O_861,N_29917,N_29737);
nor UO_862 (O_862,N_29970,N_29733);
nor UO_863 (O_863,N_29994,N_29884);
xor UO_864 (O_864,N_29880,N_29869);
xnor UO_865 (O_865,N_29544,N_29605);
xor UO_866 (O_866,N_29639,N_29692);
nor UO_867 (O_867,N_29942,N_29989);
xnor UO_868 (O_868,N_29706,N_29705);
or UO_869 (O_869,N_29790,N_29709);
nand UO_870 (O_870,N_29965,N_29945);
nor UO_871 (O_871,N_29992,N_29513);
xor UO_872 (O_872,N_29952,N_29779);
nor UO_873 (O_873,N_29648,N_29642);
or UO_874 (O_874,N_29906,N_29666);
and UO_875 (O_875,N_29719,N_29541);
or UO_876 (O_876,N_29662,N_29616);
nand UO_877 (O_877,N_29787,N_29554);
nor UO_878 (O_878,N_29792,N_29776);
or UO_879 (O_879,N_29798,N_29739);
nor UO_880 (O_880,N_29798,N_29603);
and UO_881 (O_881,N_29948,N_29791);
or UO_882 (O_882,N_29886,N_29666);
and UO_883 (O_883,N_29992,N_29915);
or UO_884 (O_884,N_29870,N_29837);
nor UO_885 (O_885,N_29876,N_29926);
xnor UO_886 (O_886,N_29728,N_29904);
or UO_887 (O_887,N_29889,N_29665);
nor UO_888 (O_888,N_29879,N_29609);
nor UO_889 (O_889,N_29776,N_29969);
nor UO_890 (O_890,N_29927,N_29882);
nor UO_891 (O_891,N_29526,N_29921);
nand UO_892 (O_892,N_29773,N_29584);
and UO_893 (O_893,N_29919,N_29977);
nor UO_894 (O_894,N_29692,N_29684);
nor UO_895 (O_895,N_29988,N_29535);
nand UO_896 (O_896,N_29982,N_29863);
nor UO_897 (O_897,N_29765,N_29604);
nand UO_898 (O_898,N_29575,N_29661);
and UO_899 (O_899,N_29751,N_29985);
nor UO_900 (O_900,N_29879,N_29830);
xnor UO_901 (O_901,N_29691,N_29738);
nand UO_902 (O_902,N_29524,N_29557);
or UO_903 (O_903,N_29684,N_29939);
xor UO_904 (O_904,N_29791,N_29518);
nor UO_905 (O_905,N_29506,N_29500);
or UO_906 (O_906,N_29581,N_29929);
or UO_907 (O_907,N_29540,N_29781);
nand UO_908 (O_908,N_29906,N_29722);
or UO_909 (O_909,N_29904,N_29829);
nand UO_910 (O_910,N_29779,N_29941);
nand UO_911 (O_911,N_29595,N_29623);
nand UO_912 (O_912,N_29779,N_29755);
xnor UO_913 (O_913,N_29972,N_29986);
or UO_914 (O_914,N_29519,N_29942);
and UO_915 (O_915,N_29766,N_29608);
nor UO_916 (O_916,N_29607,N_29815);
or UO_917 (O_917,N_29903,N_29832);
nor UO_918 (O_918,N_29611,N_29501);
nor UO_919 (O_919,N_29602,N_29703);
and UO_920 (O_920,N_29862,N_29757);
nand UO_921 (O_921,N_29628,N_29933);
xor UO_922 (O_922,N_29844,N_29686);
nor UO_923 (O_923,N_29728,N_29655);
and UO_924 (O_924,N_29642,N_29545);
and UO_925 (O_925,N_29593,N_29834);
and UO_926 (O_926,N_29548,N_29682);
nand UO_927 (O_927,N_29987,N_29608);
nand UO_928 (O_928,N_29985,N_29612);
xnor UO_929 (O_929,N_29725,N_29503);
and UO_930 (O_930,N_29847,N_29853);
or UO_931 (O_931,N_29634,N_29854);
nand UO_932 (O_932,N_29843,N_29704);
nor UO_933 (O_933,N_29717,N_29508);
xnor UO_934 (O_934,N_29946,N_29979);
nor UO_935 (O_935,N_29925,N_29677);
or UO_936 (O_936,N_29741,N_29520);
nor UO_937 (O_937,N_29967,N_29788);
and UO_938 (O_938,N_29743,N_29845);
nor UO_939 (O_939,N_29755,N_29652);
xnor UO_940 (O_940,N_29976,N_29791);
nand UO_941 (O_941,N_29967,N_29962);
nand UO_942 (O_942,N_29588,N_29910);
or UO_943 (O_943,N_29661,N_29921);
or UO_944 (O_944,N_29986,N_29871);
and UO_945 (O_945,N_29641,N_29576);
nand UO_946 (O_946,N_29847,N_29946);
and UO_947 (O_947,N_29806,N_29502);
nor UO_948 (O_948,N_29928,N_29849);
and UO_949 (O_949,N_29835,N_29981);
or UO_950 (O_950,N_29544,N_29589);
xnor UO_951 (O_951,N_29720,N_29678);
nand UO_952 (O_952,N_29543,N_29757);
and UO_953 (O_953,N_29860,N_29601);
xnor UO_954 (O_954,N_29695,N_29548);
or UO_955 (O_955,N_29584,N_29572);
xnor UO_956 (O_956,N_29636,N_29552);
xnor UO_957 (O_957,N_29657,N_29737);
and UO_958 (O_958,N_29998,N_29826);
nand UO_959 (O_959,N_29588,N_29980);
xnor UO_960 (O_960,N_29768,N_29609);
and UO_961 (O_961,N_29776,N_29867);
or UO_962 (O_962,N_29869,N_29902);
nor UO_963 (O_963,N_29758,N_29782);
and UO_964 (O_964,N_29982,N_29854);
nand UO_965 (O_965,N_29522,N_29846);
nor UO_966 (O_966,N_29894,N_29659);
xor UO_967 (O_967,N_29920,N_29990);
xnor UO_968 (O_968,N_29586,N_29874);
xor UO_969 (O_969,N_29520,N_29844);
or UO_970 (O_970,N_29679,N_29965);
nand UO_971 (O_971,N_29884,N_29929);
and UO_972 (O_972,N_29768,N_29803);
and UO_973 (O_973,N_29883,N_29704);
xor UO_974 (O_974,N_29756,N_29670);
and UO_975 (O_975,N_29836,N_29765);
nand UO_976 (O_976,N_29902,N_29834);
nand UO_977 (O_977,N_29963,N_29747);
xnor UO_978 (O_978,N_29748,N_29954);
nand UO_979 (O_979,N_29672,N_29616);
nand UO_980 (O_980,N_29961,N_29584);
and UO_981 (O_981,N_29708,N_29601);
nand UO_982 (O_982,N_29800,N_29758);
nor UO_983 (O_983,N_29794,N_29855);
nor UO_984 (O_984,N_29602,N_29738);
and UO_985 (O_985,N_29873,N_29820);
nor UO_986 (O_986,N_29541,N_29738);
nand UO_987 (O_987,N_29563,N_29780);
nor UO_988 (O_988,N_29921,N_29821);
xnor UO_989 (O_989,N_29598,N_29600);
or UO_990 (O_990,N_29893,N_29709);
nand UO_991 (O_991,N_29946,N_29546);
or UO_992 (O_992,N_29585,N_29609);
nor UO_993 (O_993,N_29821,N_29684);
nor UO_994 (O_994,N_29657,N_29565);
nor UO_995 (O_995,N_29758,N_29578);
nand UO_996 (O_996,N_29911,N_29769);
nand UO_997 (O_997,N_29875,N_29757);
and UO_998 (O_998,N_29658,N_29874);
nor UO_999 (O_999,N_29779,N_29991);
xor UO_1000 (O_1000,N_29868,N_29922);
nor UO_1001 (O_1001,N_29545,N_29962);
nor UO_1002 (O_1002,N_29847,N_29834);
nand UO_1003 (O_1003,N_29777,N_29862);
nor UO_1004 (O_1004,N_29739,N_29941);
nor UO_1005 (O_1005,N_29977,N_29749);
nand UO_1006 (O_1006,N_29547,N_29613);
and UO_1007 (O_1007,N_29969,N_29931);
nand UO_1008 (O_1008,N_29817,N_29928);
xor UO_1009 (O_1009,N_29966,N_29789);
and UO_1010 (O_1010,N_29727,N_29739);
and UO_1011 (O_1011,N_29515,N_29664);
or UO_1012 (O_1012,N_29746,N_29958);
nand UO_1013 (O_1013,N_29872,N_29508);
nor UO_1014 (O_1014,N_29861,N_29621);
nand UO_1015 (O_1015,N_29676,N_29798);
and UO_1016 (O_1016,N_29901,N_29796);
or UO_1017 (O_1017,N_29530,N_29653);
nand UO_1018 (O_1018,N_29884,N_29904);
nor UO_1019 (O_1019,N_29567,N_29743);
and UO_1020 (O_1020,N_29550,N_29843);
nor UO_1021 (O_1021,N_29839,N_29953);
nand UO_1022 (O_1022,N_29553,N_29981);
nor UO_1023 (O_1023,N_29604,N_29892);
and UO_1024 (O_1024,N_29723,N_29898);
nand UO_1025 (O_1025,N_29954,N_29719);
and UO_1026 (O_1026,N_29566,N_29811);
xor UO_1027 (O_1027,N_29692,N_29641);
and UO_1028 (O_1028,N_29803,N_29603);
and UO_1029 (O_1029,N_29964,N_29967);
nand UO_1030 (O_1030,N_29584,N_29726);
and UO_1031 (O_1031,N_29596,N_29937);
nor UO_1032 (O_1032,N_29565,N_29634);
nor UO_1033 (O_1033,N_29643,N_29704);
and UO_1034 (O_1034,N_29888,N_29680);
and UO_1035 (O_1035,N_29995,N_29548);
nor UO_1036 (O_1036,N_29894,N_29839);
nor UO_1037 (O_1037,N_29880,N_29733);
xor UO_1038 (O_1038,N_29861,N_29670);
xnor UO_1039 (O_1039,N_29987,N_29741);
xnor UO_1040 (O_1040,N_29928,N_29609);
nand UO_1041 (O_1041,N_29601,N_29743);
nand UO_1042 (O_1042,N_29956,N_29518);
nor UO_1043 (O_1043,N_29885,N_29595);
xor UO_1044 (O_1044,N_29978,N_29906);
and UO_1045 (O_1045,N_29701,N_29984);
or UO_1046 (O_1046,N_29691,N_29914);
xor UO_1047 (O_1047,N_29762,N_29962);
and UO_1048 (O_1048,N_29744,N_29925);
nand UO_1049 (O_1049,N_29705,N_29784);
nand UO_1050 (O_1050,N_29653,N_29577);
nor UO_1051 (O_1051,N_29696,N_29726);
or UO_1052 (O_1052,N_29995,N_29545);
nor UO_1053 (O_1053,N_29910,N_29533);
or UO_1054 (O_1054,N_29523,N_29948);
and UO_1055 (O_1055,N_29533,N_29683);
xnor UO_1056 (O_1056,N_29894,N_29704);
nand UO_1057 (O_1057,N_29815,N_29836);
nand UO_1058 (O_1058,N_29666,N_29629);
or UO_1059 (O_1059,N_29871,N_29626);
xor UO_1060 (O_1060,N_29731,N_29864);
nand UO_1061 (O_1061,N_29653,N_29648);
xnor UO_1062 (O_1062,N_29551,N_29660);
or UO_1063 (O_1063,N_29882,N_29871);
xnor UO_1064 (O_1064,N_29731,N_29610);
nand UO_1065 (O_1065,N_29574,N_29985);
xnor UO_1066 (O_1066,N_29978,N_29872);
and UO_1067 (O_1067,N_29962,N_29662);
and UO_1068 (O_1068,N_29874,N_29954);
nor UO_1069 (O_1069,N_29793,N_29827);
nand UO_1070 (O_1070,N_29776,N_29645);
nor UO_1071 (O_1071,N_29613,N_29649);
nand UO_1072 (O_1072,N_29623,N_29581);
and UO_1073 (O_1073,N_29789,N_29546);
nand UO_1074 (O_1074,N_29798,N_29998);
xor UO_1075 (O_1075,N_29719,N_29627);
xnor UO_1076 (O_1076,N_29749,N_29921);
nor UO_1077 (O_1077,N_29720,N_29602);
nand UO_1078 (O_1078,N_29885,N_29879);
or UO_1079 (O_1079,N_29598,N_29579);
nor UO_1080 (O_1080,N_29870,N_29691);
and UO_1081 (O_1081,N_29595,N_29695);
xnor UO_1082 (O_1082,N_29967,N_29886);
and UO_1083 (O_1083,N_29952,N_29582);
and UO_1084 (O_1084,N_29986,N_29933);
nor UO_1085 (O_1085,N_29992,N_29999);
nor UO_1086 (O_1086,N_29899,N_29967);
and UO_1087 (O_1087,N_29593,N_29651);
or UO_1088 (O_1088,N_29698,N_29761);
nand UO_1089 (O_1089,N_29955,N_29719);
xor UO_1090 (O_1090,N_29826,N_29653);
and UO_1091 (O_1091,N_29739,N_29862);
xnor UO_1092 (O_1092,N_29989,N_29793);
or UO_1093 (O_1093,N_29720,N_29759);
xor UO_1094 (O_1094,N_29678,N_29676);
and UO_1095 (O_1095,N_29727,N_29611);
nor UO_1096 (O_1096,N_29842,N_29791);
xnor UO_1097 (O_1097,N_29678,N_29786);
or UO_1098 (O_1098,N_29964,N_29961);
nand UO_1099 (O_1099,N_29616,N_29904);
nand UO_1100 (O_1100,N_29629,N_29834);
nor UO_1101 (O_1101,N_29540,N_29522);
and UO_1102 (O_1102,N_29915,N_29539);
nand UO_1103 (O_1103,N_29799,N_29648);
or UO_1104 (O_1104,N_29791,N_29987);
xnor UO_1105 (O_1105,N_29632,N_29801);
and UO_1106 (O_1106,N_29944,N_29807);
nor UO_1107 (O_1107,N_29821,N_29629);
xnor UO_1108 (O_1108,N_29750,N_29896);
or UO_1109 (O_1109,N_29918,N_29785);
nor UO_1110 (O_1110,N_29982,N_29629);
nor UO_1111 (O_1111,N_29941,N_29504);
and UO_1112 (O_1112,N_29666,N_29867);
and UO_1113 (O_1113,N_29645,N_29755);
and UO_1114 (O_1114,N_29545,N_29898);
or UO_1115 (O_1115,N_29570,N_29829);
xor UO_1116 (O_1116,N_29806,N_29506);
xnor UO_1117 (O_1117,N_29663,N_29532);
or UO_1118 (O_1118,N_29983,N_29632);
nor UO_1119 (O_1119,N_29608,N_29768);
nor UO_1120 (O_1120,N_29973,N_29703);
or UO_1121 (O_1121,N_29671,N_29955);
xnor UO_1122 (O_1122,N_29873,N_29603);
and UO_1123 (O_1123,N_29877,N_29871);
and UO_1124 (O_1124,N_29636,N_29540);
nand UO_1125 (O_1125,N_29635,N_29761);
nand UO_1126 (O_1126,N_29696,N_29821);
xor UO_1127 (O_1127,N_29562,N_29764);
and UO_1128 (O_1128,N_29708,N_29605);
nor UO_1129 (O_1129,N_29687,N_29514);
or UO_1130 (O_1130,N_29735,N_29817);
and UO_1131 (O_1131,N_29883,N_29569);
and UO_1132 (O_1132,N_29670,N_29808);
and UO_1133 (O_1133,N_29812,N_29626);
nand UO_1134 (O_1134,N_29524,N_29795);
or UO_1135 (O_1135,N_29864,N_29929);
and UO_1136 (O_1136,N_29512,N_29979);
or UO_1137 (O_1137,N_29637,N_29941);
and UO_1138 (O_1138,N_29725,N_29955);
or UO_1139 (O_1139,N_29616,N_29981);
or UO_1140 (O_1140,N_29857,N_29574);
and UO_1141 (O_1141,N_29894,N_29628);
nor UO_1142 (O_1142,N_29774,N_29842);
nand UO_1143 (O_1143,N_29941,N_29717);
nor UO_1144 (O_1144,N_29722,N_29980);
or UO_1145 (O_1145,N_29981,N_29855);
or UO_1146 (O_1146,N_29712,N_29600);
nand UO_1147 (O_1147,N_29611,N_29502);
nand UO_1148 (O_1148,N_29658,N_29724);
or UO_1149 (O_1149,N_29748,N_29522);
nand UO_1150 (O_1150,N_29691,N_29612);
or UO_1151 (O_1151,N_29754,N_29987);
or UO_1152 (O_1152,N_29963,N_29588);
nor UO_1153 (O_1153,N_29942,N_29710);
and UO_1154 (O_1154,N_29987,N_29746);
or UO_1155 (O_1155,N_29826,N_29560);
and UO_1156 (O_1156,N_29541,N_29862);
nor UO_1157 (O_1157,N_29503,N_29505);
xor UO_1158 (O_1158,N_29802,N_29789);
nand UO_1159 (O_1159,N_29684,N_29576);
xnor UO_1160 (O_1160,N_29908,N_29611);
xor UO_1161 (O_1161,N_29616,N_29611);
and UO_1162 (O_1162,N_29807,N_29933);
xor UO_1163 (O_1163,N_29869,N_29691);
xnor UO_1164 (O_1164,N_29826,N_29952);
or UO_1165 (O_1165,N_29888,N_29594);
nor UO_1166 (O_1166,N_29602,N_29918);
nand UO_1167 (O_1167,N_29817,N_29811);
or UO_1168 (O_1168,N_29801,N_29858);
or UO_1169 (O_1169,N_29609,N_29623);
nor UO_1170 (O_1170,N_29853,N_29969);
nor UO_1171 (O_1171,N_29797,N_29540);
or UO_1172 (O_1172,N_29737,N_29563);
and UO_1173 (O_1173,N_29897,N_29674);
nor UO_1174 (O_1174,N_29573,N_29641);
xor UO_1175 (O_1175,N_29819,N_29899);
nor UO_1176 (O_1176,N_29694,N_29697);
xnor UO_1177 (O_1177,N_29753,N_29509);
nor UO_1178 (O_1178,N_29923,N_29983);
nand UO_1179 (O_1179,N_29553,N_29631);
or UO_1180 (O_1180,N_29733,N_29748);
nand UO_1181 (O_1181,N_29779,N_29548);
and UO_1182 (O_1182,N_29987,N_29916);
xnor UO_1183 (O_1183,N_29625,N_29649);
xnor UO_1184 (O_1184,N_29616,N_29708);
nor UO_1185 (O_1185,N_29568,N_29887);
nand UO_1186 (O_1186,N_29734,N_29622);
or UO_1187 (O_1187,N_29920,N_29736);
nor UO_1188 (O_1188,N_29730,N_29573);
nor UO_1189 (O_1189,N_29575,N_29715);
or UO_1190 (O_1190,N_29927,N_29988);
and UO_1191 (O_1191,N_29697,N_29656);
nor UO_1192 (O_1192,N_29971,N_29788);
nand UO_1193 (O_1193,N_29873,N_29771);
xnor UO_1194 (O_1194,N_29846,N_29723);
and UO_1195 (O_1195,N_29746,N_29600);
and UO_1196 (O_1196,N_29705,N_29979);
or UO_1197 (O_1197,N_29584,N_29974);
or UO_1198 (O_1198,N_29928,N_29905);
and UO_1199 (O_1199,N_29759,N_29551);
xor UO_1200 (O_1200,N_29983,N_29979);
nor UO_1201 (O_1201,N_29680,N_29879);
and UO_1202 (O_1202,N_29838,N_29833);
nand UO_1203 (O_1203,N_29535,N_29816);
nor UO_1204 (O_1204,N_29941,N_29850);
and UO_1205 (O_1205,N_29691,N_29780);
and UO_1206 (O_1206,N_29579,N_29721);
nand UO_1207 (O_1207,N_29893,N_29748);
and UO_1208 (O_1208,N_29551,N_29734);
nor UO_1209 (O_1209,N_29549,N_29824);
nand UO_1210 (O_1210,N_29706,N_29972);
xnor UO_1211 (O_1211,N_29857,N_29769);
nand UO_1212 (O_1212,N_29826,N_29862);
or UO_1213 (O_1213,N_29895,N_29705);
nand UO_1214 (O_1214,N_29606,N_29967);
or UO_1215 (O_1215,N_29664,N_29808);
or UO_1216 (O_1216,N_29705,N_29662);
and UO_1217 (O_1217,N_29957,N_29627);
nand UO_1218 (O_1218,N_29981,N_29815);
nand UO_1219 (O_1219,N_29780,N_29618);
nand UO_1220 (O_1220,N_29685,N_29703);
and UO_1221 (O_1221,N_29647,N_29956);
nor UO_1222 (O_1222,N_29766,N_29609);
and UO_1223 (O_1223,N_29977,N_29708);
xor UO_1224 (O_1224,N_29706,N_29578);
nor UO_1225 (O_1225,N_29682,N_29956);
or UO_1226 (O_1226,N_29758,N_29746);
nor UO_1227 (O_1227,N_29791,N_29971);
nor UO_1228 (O_1228,N_29681,N_29737);
nand UO_1229 (O_1229,N_29659,N_29501);
xnor UO_1230 (O_1230,N_29687,N_29880);
nor UO_1231 (O_1231,N_29537,N_29943);
and UO_1232 (O_1232,N_29653,N_29636);
nand UO_1233 (O_1233,N_29898,N_29600);
nand UO_1234 (O_1234,N_29599,N_29876);
nand UO_1235 (O_1235,N_29882,N_29831);
or UO_1236 (O_1236,N_29998,N_29690);
and UO_1237 (O_1237,N_29534,N_29997);
or UO_1238 (O_1238,N_29760,N_29771);
nand UO_1239 (O_1239,N_29637,N_29675);
and UO_1240 (O_1240,N_29666,N_29762);
xor UO_1241 (O_1241,N_29567,N_29950);
nand UO_1242 (O_1242,N_29925,N_29932);
nor UO_1243 (O_1243,N_29520,N_29711);
xor UO_1244 (O_1244,N_29676,N_29963);
nand UO_1245 (O_1245,N_29872,N_29750);
and UO_1246 (O_1246,N_29956,N_29670);
nand UO_1247 (O_1247,N_29567,N_29699);
and UO_1248 (O_1248,N_29691,N_29708);
nand UO_1249 (O_1249,N_29993,N_29695);
or UO_1250 (O_1250,N_29887,N_29551);
and UO_1251 (O_1251,N_29630,N_29880);
nor UO_1252 (O_1252,N_29517,N_29963);
and UO_1253 (O_1253,N_29575,N_29691);
nor UO_1254 (O_1254,N_29806,N_29650);
xnor UO_1255 (O_1255,N_29802,N_29621);
or UO_1256 (O_1256,N_29566,N_29544);
nor UO_1257 (O_1257,N_29842,N_29944);
xnor UO_1258 (O_1258,N_29635,N_29730);
and UO_1259 (O_1259,N_29977,N_29956);
and UO_1260 (O_1260,N_29689,N_29930);
or UO_1261 (O_1261,N_29868,N_29517);
nor UO_1262 (O_1262,N_29905,N_29944);
nor UO_1263 (O_1263,N_29838,N_29687);
nand UO_1264 (O_1264,N_29562,N_29553);
and UO_1265 (O_1265,N_29567,N_29787);
xor UO_1266 (O_1266,N_29598,N_29689);
nand UO_1267 (O_1267,N_29691,N_29818);
xnor UO_1268 (O_1268,N_29639,N_29613);
nand UO_1269 (O_1269,N_29757,N_29790);
nor UO_1270 (O_1270,N_29800,N_29927);
nor UO_1271 (O_1271,N_29509,N_29813);
or UO_1272 (O_1272,N_29942,N_29806);
and UO_1273 (O_1273,N_29610,N_29623);
xor UO_1274 (O_1274,N_29936,N_29558);
and UO_1275 (O_1275,N_29931,N_29608);
xor UO_1276 (O_1276,N_29660,N_29512);
xnor UO_1277 (O_1277,N_29657,N_29814);
xnor UO_1278 (O_1278,N_29918,N_29965);
xor UO_1279 (O_1279,N_29577,N_29773);
nand UO_1280 (O_1280,N_29853,N_29880);
nor UO_1281 (O_1281,N_29841,N_29552);
nand UO_1282 (O_1282,N_29991,N_29726);
or UO_1283 (O_1283,N_29983,N_29548);
xor UO_1284 (O_1284,N_29570,N_29679);
and UO_1285 (O_1285,N_29925,N_29740);
or UO_1286 (O_1286,N_29919,N_29821);
and UO_1287 (O_1287,N_29738,N_29699);
nand UO_1288 (O_1288,N_29858,N_29874);
xnor UO_1289 (O_1289,N_29993,N_29973);
xnor UO_1290 (O_1290,N_29959,N_29815);
nand UO_1291 (O_1291,N_29821,N_29588);
or UO_1292 (O_1292,N_29633,N_29870);
and UO_1293 (O_1293,N_29819,N_29782);
or UO_1294 (O_1294,N_29793,N_29997);
nand UO_1295 (O_1295,N_29554,N_29540);
xor UO_1296 (O_1296,N_29985,N_29937);
or UO_1297 (O_1297,N_29741,N_29511);
xnor UO_1298 (O_1298,N_29843,N_29817);
and UO_1299 (O_1299,N_29971,N_29859);
nor UO_1300 (O_1300,N_29596,N_29952);
nor UO_1301 (O_1301,N_29835,N_29692);
or UO_1302 (O_1302,N_29610,N_29543);
xnor UO_1303 (O_1303,N_29859,N_29773);
nand UO_1304 (O_1304,N_29843,N_29834);
xnor UO_1305 (O_1305,N_29751,N_29731);
nand UO_1306 (O_1306,N_29544,N_29549);
nand UO_1307 (O_1307,N_29947,N_29666);
xor UO_1308 (O_1308,N_29624,N_29596);
or UO_1309 (O_1309,N_29521,N_29506);
or UO_1310 (O_1310,N_29571,N_29804);
and UO_1311 (O_1311,N_29524,N_29683);
nand UO_1312 (O_1312,N_29539,N_29733);
nor UO_1313 (O_1313,N_29908,N_29909);
and UO_1314 (O_1314,N_29747,N_29993);
nand UO_1315 (O_1315,N_29976,N_29981);
xor UO_1316 (O_1316,N_29621,N_29865);
nand UO_1317 (O_1317,N_29681,N_29839);
or UO_1318 (O_1318,N_29518,N_29810);
nand UO_1319 (O_1319,N_29788,N_29637);
or UO_1320 (O_1320,N_29588,N_29820);
nor UO_1321 (O_1321,N_29672,N_29653);
and UO_1322 (O_1322,N_29994,N_29716);
or UO_1323 (O_1323,N_29891,N_29581);
xnor UO_1324 (O_1324,N_29828,N_29831);
nor UO_1325 (O_1325,N_29867,N_29541);
nor UO_1326 (O_1326,N_29867,N_29570);
nor UO_1327 (O_1327,N_29628,N_29721);
xnor UO_1328 (O_1328,N_29638,N_29793);
nand UO_1329 (O_1329,N_29716,N_29938);
xor UO_1330 (O_1330,N_29872,N_29694);
xor UO_1331 (O_1331,N_29893,N_29777);
or UO_1332 (O_1332,N_29662,N_29761);
or UO_1333 (O_1333,N_29513,N_29971);
nand UO_1334 (O_1334,N_29692,N_29579);
nor UO_1335 (O_1335,N_29713,N_29656);
and UO_1336 (O_1336,N_29782,N_29795);
or UO_1337 (O_1337,N_29555,N_29584);
and UO_1338 (O_1338,N_29894,N_29769);
nor UO_1339 (O_1339,N_29961,N_29859);
and UO_1340 (O_1340,N_29635,N_29557);
nor UO_1341 (O_1341,N_29542,N_29962);
and UO_1342 (O_1342,N_29792,N_29932);
or UO_1343 (O_1343,N_29950,N_29620);
nand UO_1344 (O_1344,N_29870,N_29879);
nand UO_1345 (O_1345,N_29618,N_29561);
xor UO_1346 (O_1346,N_29960,N_29843);
or UO_1347 (O_1347,N_29972,N_29893);
xnor UO_1348 (O_1348,N_29977,N_29582);
nand UO_1349 (O_1349,N_29767,N_29722);
xnor UO_1350 (O_1350,N_29722,N_29545);
xnor UO_1351 (O_1351,N_29507,N_29951);
and UO_1352 (O_1352,N_29520,N_29868);
or UO_1353 (O_1353,N_29958,N_29759);
or UO_1354 (O_1354,N_29708,N_29681);
nor UO_1355 (O_1355,N_29734,N_29953);
and UO_1356 (O_1356,N_29809,N_29541);
and UO_1357 (O_1357,N_29755,N_29691);
nor UO_1358 (O_1358,N_29886,N_29855);
nor UO_1359 (O_1359,N_29881,N_29517);
nand UO_1360 (O_1360,N_29733,N_29634);
or UO_1361 (O_1361,N_29788,N_29867);
nor UO_1362 (O_1362,N_29699,N_29763);
xnor UO_1363 (O_1363,N_29674,N_29704);
and UO_1364 (O_1364,N_29701,N_29966);
or UO_1365 (O_1365,N_29986,N_29527);
or UO_1366 (O_1366,N_29912,N_29993);
or UO_1367 (O_1367,N_29509,N_29994);
or UO_1368 (O_1368,N_29511,N_29831);
nor UO_1369 (O_1369,N_29604,N_29622);
and UO_1370 (O_1370,N_29898,N_29795);
and UO_1371 (O_1371,N_29955,N_29805);
nor UO_1372 (O_1372,N_29731,N_29573);
or UO_1373 (O_1373,N_29673,N_29766);
nor UO_1374 (O_1374,N_29686,N_29741);
and UO_1375 (O_1375,N_29650,N_29816);
or UO_1376 (O_1376,N_29745,N_29613);
nand UO_1377 (O_1377,N_29534,N_29852);
or UO_1378 (O_1378,N_29696,N_29923);
nand UO_1379 (O_1379,N_29843,N_29830);
and UO_1380 (O_1380,N_29505,N_29964);
and UO_1381 (O_1381,N_29564,N_29583);
or UO_1382 (O_1382,N_29953,N_29714);
or UO_1383 (O_1383,N_29784,N_29656);
and UO_1384 (O_1384,N_29980,N_29637);
nand UO_1385 (O_1385,N_29848,N_29721);
or UO_1386 (O_1386,N_29864,N_29915);
xnor UO_1387 (O_1387,N_29893,N_29586);
xnor UO_1388 (O_1388,N_29740,N_29644);
xor UO_1389 (O_1389,N_29798,N_29656);
and UO_1390 (O_1390,N_29793,N_29713);
xnor UO_1391 (O_1391,N_29611,N_29797);
and UO_1392 (O_1392,N_29500,N_29655);
and UO_1393 (O_1393,N_29886,N_29576);
and UO_1394 (O_1394,N_29874,N_29653);
or UO_1395 (O_1395,N_29536,N_29738);
or UO_1396 (O_1396,N_29630,N_29731);
or UO_1397 (O_1397,N_29673,N_29704);
nor UO_1398 (O_1398,N_29506,N_29811);
xor UO_1399 (O_1399,N_29817,N_29592);
xor UO_1400 (O_1400,N_29587,N_29799);
nand UO_1401 (O_1401,N_29831,N_29540);
nand UO_1402 (O_1402,N_29655,N_29510);
nor UO_1403 (O_1403,N_29722,N_29753);
nor UO_1404 (O_1404,N_29864,N_29542);
or UO_1405 (O_1405,N_29920,N_29800);
nor UO_1406 (O_1406,N_29937,N_29991);
nor UO_1407 (O_1407,N_29901,N_29973);
xor UO_1408 (O_1408,N_29994,N_29791);
nor UO_1409 (O_1409,N_29667,N_29679);
xor UO_1410 (O_1410,N_29903,N_29529);
xor UO_1411 (O_1411,N_29949,N_29521);
nor UO_1412 (O_1412,N_29754,N_29680);
or UO_1413 (O_1413,N_29553,N_29921);
nand UO_1414 (O_1414,N_29660,N_29582);
and UO_1415 (O_1415,N_29609,N_29690);
nor UO_1416 (O_1416,N_29935,N_29586);
nor UO_1417 (O_1417,N_29988,N_29533);
nor UO_1418 (O_1418,N_29696,N_29752);
and UO_1419 (O_1419,N_29616,N_29794);
nand UO_1420 (O_1420,N_29868,N_29857);
xor UO_1421 (O_1421,N_29853,N_29761);
and UO_1422 (O_1422,N_29803,N_29926);
xnor UO_1423 (O_1423,N_29745,N_29919);
or UO_1424 (O_1424,N_29824,N_29773);
xnor UO_1425 (O_1425,N_29529,N_29825);
nor UO_1426 (O_1426,N_29777,N_29510);
xnor UO_1427 (O_1427,N_29740,N_29685);
nor UO_1428 (O_1428,N_29602,N_29501);
and UO_1429 (O_1429,N_29581,N_29938);
or UO_1430 (O_1430,N_29573,N_29930);
nor UO_1431 (O_1431,N_29768,N_29887);
or UO_1432 (O_1432,N_29755,N_29785);
nor UO_1433 (O_1433,N_29590,N_29645);
and UO_1434 (O_1434,N_29569,N_29960);
or UO_1435 (O_1435,N_29503,N_29791);
or UO_1436 (O_1436,N_29615,N_29547);
xor UO_1437 (O_1437,N_29990,N_29718);
nor UO_1438 (O_1438,N_29571,N_29947);
or UO_1439 (O_1439,N_29880,N_29502);
or UO_1440 (O_1440,N_29963,N_29568);
and UO_1441 (O_1441,N_29588,N_29511);
and UO_1442 (O_1442,N_29618,N_29838);
nand UO_1443 (O_1443,N_29985,N_29580);
and UO_1444 (O_1444,N_29929,N_29790);
nand UO_1445 (O_1445,N_29834,N_29857);
and UO_1446 (O_1446,N_29711,N_29501);
nor UO_1447 (O_1447,N_29611,N_29525);
or UO_1448 (O_1448,N_29713,N_29999);
or UO_1449 (O_1449,N_29876,N_29700);
xnor UO_1450 (O_1450,N_29556,N_29956);
nor UO_1451 (O_1451,N_29801,N_29883);
or UO_1452 (O_1452,N_29955,N_29557);
nand UO_1453 (O_1453,N_29893,N_29970);
or UO_1454 (O_1454,N_29976,N_29992);
and UO_1455 (O_1455,N_29840,N_29653);
nor UO_1456 (O_1456,N_29718,N_29795);
nor UO_1457 (O_1457,N_29538,N_29836);
xnor UO_1458 (O_1458,N_29540,N_29962);
nand UO_1459 (O_1459,N_29749,N_29770);
xor UO_1460 (O_1460,N_29780,N_29775);
nand UO_1461 (O_1461,N_29577,N_29533);
nand UO_1462 (O_1462,N_29534,N_29824);
xnor UO_1463 (O_1463,N_29699,N_29568);
xor UO_1464 (O_1464,N_29551,N_29841);
xor UO_1465 (O_1465,N_29791,N_29866);
and UO_1466 (O_1466,N_29958,N_29687);
and UO_1467 (O_1467,N_29773,N_29616);
nand UO_1468 (O_1468,N_29643,N_29572);
nor UO_1469 (O_1469,N_29977,N_29529);
and UO_1470 (O_1470,N_29641,N_29870);
xnor UO_1471 (O_1471,N_29590,N_29622);
and UO_1472 (O_1472,N_29663,N_29767);
nand UO_1473 (O_1473,N_29900,N_29613);
or UO_1474 (O_1474,N_29677,N_29521);
nand UO_1475 (O_1475,N_29515,N_29509);
or UO_1476 (O_1476,N_29760,N_29628);
nand UO_1477 (O_1477,N_29521,N_29707);
xnor UO_1478 (O_1478,N_29610,N_29849);
or UO_1479 (O_1479,N_29950,N_29575);
nor UO_1480 (O_1480,N_29900,N_29766);
and UO_1481 (O_1481,N_29873,N_29908);
or UO_1482 (O_1482,N_29548,N_29872);
xnor UO_1483 (O_1483,N_29816,N_29717);
nor UO_1484 (O_1484,N_29951,N_29641);
or UO_1485 (O_1485,N_29759,N_29942);
or UO_1486 (O_1486,N_29646,N_29901);
xnor UO_1487 (O_1487,N_29694,N_29910);
xor UO_1488 (O_1488,N_29684,N_29674);
or UO_1489 (O_1489,N_29530,N_29948);
and UO_1490 (O_1490,N_29871,N_29609);
nor UO_1491 (O_1491,N_29804,N_29797);
xnor UO_1492 (O_1492,N_29975,N_29685);
and UO_1493 (O_1493,N_29953,N_29843);
and UO_1494 (O_1494,N_29884,N_29701);
or UO_1495 (O_1495,N_29940,N_29672);
xnor UO_1496 (O_1496,N_29831,N_29902);
nand UO_1497 (O_1497,N_29717,N_29750);
and UO_1498 (O_1498,N_29983,N_29716);
or UO_1499 (O_1499,N_29721,N_29666);
nand UO_1500 (O_1500,N_29754,N_29548);
or UO_1501 (O_1501,N_29763,N_29638);
and UO_1502 (O_1502,N_29903,N_29789);
nor UO_1503 (O_1503,N_29688,N_29553);
or UO_1504 (O_1504,N_29636,N_29666);
nor UO_1505 (O_1505,N_29945,N_29849);
or UO_1506 (O_1506,N_29849,N_29979);
xor UO_1507 (O_1507,N_29855,N_29559);
and UO_1508 (O_1508,N_29509,N_29504);
or UO_1509 (O_1509,N_29992,N_29545);
or UO_1510 (O_1510,N_29669,N_29776);
xnor UO_1511 (O_1511,N_29673,N_29835);
nor UO_1512 (O_1512,N_29870,N_29969);
nand UO_1513 (O_1513,N_29658,N_29670);
or UO_1514 (O_1514,N_29882,N_29690);
xor UO_1515 (O_1515,N_29885,N_29823);
xnor UO_1516 (O_1516,N_29935,N_29961);
nand UO_1517 (O_1517,N_29764,N_29873);
nand UO_1518 (O_1518,N_29876,N_29955);
and UO_1519 (O_1519,N_29661,N_29585);
xnor UO_1520 (O_1520,N_29526,N_29915);
and UO_1521 (O_1521,N_29551,N_29501);
nor UO_1522 (O_1522,N_29968,N_29757);
nand UO_1523 (O_1523,N_29939,N_29677);
or UO_1524 (O_1524,N_29860,N_29642);
nor UO_1525 (O_1525,N_29721,N_29594);
nand UO_1526 (O_1526,N_29871,N_29673);
nor UO_1527 (O_1527,N_29643,N_29909);
and UO_1528 (O_1528,N_29802,N_29634);
nor UO_1529 (O_1529,N_29619,N_29780);
or UO_1530 (O_1530,N_29855,N_29937);
nand UO_1531 (O_1531,N_29861,N_29964);
nand UO_1532 (O_1532,N_29792,N_29690);
xnor UO_1533 (O_1533,N_29687,N_29780);
or UO_1534 (O_1534,N_29903,N_29605);
nor UO_1535 (O_1535,N_29590,N_29585);
or UO_1536 (O_1536,N_29916,N_29720);
nor UO_1537 (O_1537,N_29846,N_29651);
or UO_1538 (O_1538,N_29841,N_29682);
nor UO_1539 (O_1539,N_29689,N_29691);
xor UO_1540 (O_1540,N_29754,N_29847);
or UO_1541 (O_1541,N_29802,N_29962);
nand UO_1542 (O_1542,N_29794,N_29734);
xor UO_1543 (O_1543,N_29545,N_29928);
nand UO_1544 (O_1544,N_29761,N_29987);
and UO_1545 (O_1545,N_29983,N_29970);
nor UO_1546 (O_1546,N_29749,N_29744);
or UO_1547 (O_1547,N_29632,N_29989);
and UO_1548 (O_1548,N_29885,N_29604);
nor UO_1549 (O_1549,N_29609,N_29740);
xnor UO_1550 (O_1550,N_29615,N_29794);
nor UO_1551 (O_1551,N_29884,N_29536);
xnor UO_1552 (O_1552,N_29942,N_29722);
or UO_1553 (O_1553,N_29831,N_29778);
nand UO_1554 (O_1554,N_29540,N_29905);
or UO_1555 (O_1555,N_29730,N_29657);
nor UO_1556 (O_1556,N_29803,N_29584);
and UO_1557 (O_1557,N_29895,N_29839);
xor UO_1558 (O_1558,N_29924,N_29866);
and UO_1559 (O_1559,N_29802,N_29806);
nand UO_1560 (O_1560,N_29666,N_29884);
and UO_1561 (O_1561,N_29596,N_29528);
or UO_1562 (O_1562,N_29571,N_29841);
or UO_1563 (O_1563,N_29715,N_29654);
xnor UO_1564 (O_1564,N_29845,N_29501);
nor UO_1565 (O_1565,N_29601,N_29698);
and UO_1566 (O_1566,N_29909,N_29963);
or UO_1567 (O_1567,N_29530,N_29533);
nor UO_1568 (O_1568,N_29570,N_29566);
or UO_1569 (O_1569,N_29809,N_29859);
or UO_1570 (O_1570,N_29588,N_29710);
nor UO_1571 (O_1571,N_29742,N_29564);
nor UO_1572 (O_1572,N_29857,N_29794);
or UO_1573 (O_1573,N_29782,N_29725);
and UO_1574 (O_1574,N_29581,N_29710);
or UO_1575 (O_1575,N_29797,N_29607);
nand UO_1576 (O_1576,N_29717,N_29649);
and UO_1577 (O_1577,N_29551,N_29981);
nand UO_1578 (O_1578,N_29749,N_29613);
nand UO_1579 (O_1579,N_29523,N_29624);
or UO_1580 (O_1580,N_29575,N_29512);
nand UO_1581 (O_1581,N_29839,N_29960);
and UO_1582 (O_1582,N_29549,N_29536);
nor UO_1583 (O_1583,N_29582,N_29745);
nand UO_1584 (O_1584,N_29963,N_29846);
or UO_1585 (O_1585,N_29539,N_29679);
and UO_1586 (O_1586,N_29617,N_29503);
xnor UO_1587 (O_1587,N_29749,N_29865);
nor UO_1588 (O_1588,N_29744,N_29891);
nor UO_1589 (O_1589,N_29704,N_29918);
xnor UO_1590 (O_1590,N_29787,N_29923);
xor UO_1591 (O_1591,N_29938,N_29868);
nand UO_1592 (O_1592,N_29651,N_29859);
nand UO_1593 (O_1593,N_29779,N_29551);
nor UO_1594 (O_1594,N_29627,N_29702);
and UO_1595 (O_1595,N_29691,N_29736);
nor UO_1596 (O_1596,N_29857,N_29987);
and UO_1597 (O_1597,N_29589,N_29637);
and UO_1598 (O_1598,N_29895,N_29802);
nand UO_1599 (O_1599,N_29849,N_29674);
nand UO_1600 (O_1600,N_29634,N_29717);
nor UO_1601 (O_1601,N_29858,N_29739);
and UO_1602 (O_1602,N_29901,N_29639);
xor UO_1603 (O_1603,N_29567,N_29874);
and UO_1604 (O_1604,N_29535,N_29511);
and UO_1605 (O_1605,N_29631,N_29974);
nand UO_1606 (O_1606,N_29590,N_29995);
and UO_1607 (O_1607,N_29799,N_29630);
nor UO_1608 (O_1608,N_29530,N_29565);
xnor UO_1609 (O_1609,N_29559,N_29537);
nand UO_1610 (O_1610,N_29817,N_29586);
nand UO_1611 (O_1611,N_29609,N_29844);
and UO_1612 (O_1612,N_29569,N_29978);
and UO_1613 (O_1613,N_29556,N_29960);
nand UO_1614 (O_1614,N_29583,N_29996);
nor UO_1615 (O_1615,N_29719,N_29684);
nand UO_1616 (O_1616,N_29737,N_29613);
and UO_1617 (O_1617,N_29794,N_29575);
and UO_1618 (O_1618,N_29947,N_29700);
xor UO_1619 (O_1619,N_29530,N_29690);
and UO_1620 (O_1620,N_29766,N_29890);
and UO_1621 (O_1621,N_29835,N_29999);
xor UO_1622 (O_1622,N_29664,N_29999);
and UO_1623 (O_1623,N_29902,N_29572);
xnor UO_1624 (O_1624,N_29883,N_29984);
nand UO_1625 (O_1625,N_29699,N_29791);
and UO_1626 (O_1626,N_29777,N_29653);
or UO_1627 (O_1627,N_29989,N_29934);
nand UO_1628 (O_1628,N_29873,N_29532);
or UO_1629 (O_1629,N_29977,N_29858);
nand UO_1630 (O_1630,N_29831,N_29723);
and UO_1631 (O_1631,N_29907,N_29642);
or UO_1632 (O_1632,N_29507,N_29844);
or UO_1633 (O_1633,N_29640,N_29779);
xor UO_1634 (O_1634,N_29528,N_29601);
nand UO_1635 (O_1635,N_29959,N_29892);
and UO_1636 (O_1636,N_29870,N_29709);
nand UO_1637 (O_1637,N_29779,N_29661);
xor UO_1638 (O_1638,N_29689,N_29511);
xor UO_1639 (O_1639,N_29588,N_29544);
nand UO_1640 (O_1640,N_29554,N_29515);
or UO_1641 (O_1641,N_29527,N_29902);
xor UO_1642 (O_1642,N_29876,N_29977);
nand UO_1643 (O_1643,N_29643,N_29517);
nor UO_1644 (O_1644,N_29827,N_29977);
or UO_1645 (O_1645,N_29599,N_29603);
nor UO_1646 (O_1646,N_29847,N_29964);
nor UO_1647 (O_1647,N_29587,N_29644);
or UO_1648 (O_1648,N_29597,N_29514);
nor UO_1649 (O_1649,N_29750,N_29706);
xor UO_1650 (O_1650,N_29524,N_29534);
nor UO_1651 (O_1651,N_29552,N_29559);
xnor UO_1652 (O_1652,N_29680,N_29951);
nand UO_1653 (O_1653,N_29834,N_29501);
xnor UO_1654 (O_1654,N_29964,N_29583);
nor UO_1655 (O_1655,N_29629,N_29841);
and UO_1656 (O_1656,N_29661,N_29936);
or UO_1657 (O_1657,N_29591,N_29650);
xnor UO_1658 (O_1658,N_29802,N_29515);
nor UO_1659 (O_1659,N_29560,N_29976);
nand UO_1660 (O_1660,N_29729,N_29664);
or UO_1661 (O_1661,N_29930,N_29503);
nand UO_1662 (O_1662,N_29806,N_29552);
and UO_1663 (O_1663,N_29960,N_29932);
nand UO_1664 (O_1664,N_29913,N_29858);
xor UO_1665 (O_1665,N_29971,N_29532);
or UO_1666 (O_1666,N_29879,N_29708);
xor UO_1667 (O_1667,N_29933,N_29869);
nand UO_1668 (O_1668,N_29749,N_29616);
nand UO_1669 (O_1669,N_29862,N_29995);
nand UO_1670 (O_1670,N_29652,N_29819);
nor UO_1671 (O_1671,N_29649,N_29987);
and UO_1672 (O_1672,N_29972,N_29720);
nor UO_1673 (O_1673,N_29892,N_29717);
xor UO_1674 (O_1674,N_29817,N_29582);
or UO_1675 (O_1675,N_29690,N_29618);
nand UO_1676 (O_1676,N_29781,N_29519);
xor UO_1677 (O_1677,N_29805,N_29569);
or UO_1678 (O_1678,N_29971,N_29641);
nor UO_1679 (O_1679,N_29638,N_29932);
nor UO_1680 (O_1680,N_29602,N_29521);
or UO_1681 (O_1681,N_29959,N_29764);
nand UO_1682 (O_1682,N_29772,N_29698);
nor UO_1683 (O_1683,N_29823,N_29722);
or UO_1684 (O_1684,N_29672,N_29868);
xnor UO_1685 (O_1685,N_29733,N_29963);
or UO_1686 (O_1686,N_29990,N_29933);
xnor UO_1687 (O_1687,N_29950,N_29762);
and UO_1688 (O_1688,N_29862,N_29919);
or UO_1689 (O_1689,N_29591,N_29850);
and UO_1690 (O_1690,N_29743,N_29838);
nand UO_1691 (O_1691,N_29759,N_29532);
and UO_1692 (O_1692,N_29836,N_29740);
and UO_1693 (O_1693,N_29737,N_29829);
and UO_1694 (O_1694,N_29686,N_29781);
xor UO_1695 (O_1695,N_29672,N_29605);
xnor UO_1696 (O_1696,N_29838,N_29772);
nor UO_1697 (O_1697,N_29813,N_29954);
xor UO_1698 (O_1698,N_29744,N_29568);
nor UO_1699 (O_1699,N_29928,N_29884);
or UO_1700 (O_1700,N_29795,N_29560);
nor UO_1701 (O_1701,N_29620,N_29986);
and UO_1702 (O_1702,N_29690,N_29834);
and UO_1703 (O_1703,N_29898,N_29807);
or UO_1704 (O_1704,N_29534,N_29895);
nor UO_1705 (O_1705,N_29967,N_29516);
or UO_1706 (O_1706,N_29758,N_29881);
and UO_1707 (O_1707,N_29869,N_29642);
or UO_1708 (O_1708,N_29656,N_29729);
or UO_1709 (O_1709,N_29767,N_29939);
or UO_1710 (O_1710,N_29631,N_29855);
and UO_1711 (O_1711,N_29697,N_29711);
xnor UO_1712 (O_1712,N_29748,N_29567);
nor UO_1713 (O_1713,N_29994,N_29779);
or UO_1714 (O_1714,N_29556,N_29574);
nor UO_1715 (O_1715,N_29927,N_29772);
xor UO_1716 (O_1716,N_29708,N_29643);
or UO_1717 (O_1717,N_29862,N_29528);
nand UO_1718 (O_1718,N_29527,N_29749);
xnor UO_1719 (O_1719,N_29949,N_29926);
nor UO_1720 (O_1720,N_29774,N_29559);
and UO_1721 (O_1721,N_29969,N_29708);
xnor UO_1722 (O_1722,N_29637,N_29960);
nand UO_1723 (O_1723,N_29710,N_29553);
nand UO_1724 (O_1724,N_29856,N_29692);
nand UO_1725 (O_1725,N_29992,N_29604);
or UO_1726 (O_1726,N_29835,N_29698);
and UO_1727 (O_1727,N_29765,N_29884);
or UO_1728 (O_1728,N_29981,N_29921);
nand UO_1729 (O_1729,N_29558,N_29877);
xnor UO_1730 (O_1730,N_29507,N_29921);
or UO_1731 (O_1731,N_29521,N_29548);
nand UO_1732 (O_1732,N_29919,N_29631);
or UO_1733 (O_1733,N_29601,N_29927);
nor UO_1734 (O_1734,N_29824,N_29820);
xor UO_1735 (O_1735,N_29938,N_29588);
nand UO_1736 (O_1736,N_29638,N_29567);
or UO_1737 (O_1737,N_29961,N_29533);
xor UO_1738 (O_1738,N_29747,N_29694);
xor UO_1739 (O_1739,N_29516,N_29686);
nor UO_1740 (O_1740,N_29545,N_29593);
nand UO_1741 (O_1741,N_29585,N_29743);
or UO_1742 (O_1742,N_29628,N_29701);
or UO_1743 (O_1743,N_29929,N_29901);
xor UO_1744 (O_1744,N_29817,N_29520);
and UO_1745 (O_1745,N_29860,N_29647);
nand UO_1746 (O_1746,N_29902,N_29866);
xnor UO_1747 (O_1747,N_29928,N_29678);
or UO_1748 (O_1748,N_29588,N_29837);
and UO_1749 (O_1749,N_29744,N_29966);
nand UO_1750 (O_1750,N_29891,N_29878);
or UO_1751 (O_1751,N_29649,N_29968);
nand UO_1752 (O_1752,N_29685,N_29946);
and UO_1753 (O_1753,N_29624,N_29851);
or UO_1754 (O_1754,N_29760,N_29885);
nor UO_1755 (O_1755,N_29758,N_29651);
or UO_1756 (O_1756,N_29740,N_29645);
nor UO_1757 (O_1757,N_29513,N_29880);
nand UO_1758 (O_1758,N_29523,N_29774);
and UO_1759 (O_1759,N_29554,N_29524);
and UO_1760 (O_1760,N_29860,N_29894);
or UO_1761 (O_1761,N_29776,N_29595);
and UO_1762 (O_1762,N_29982,N_29984);
nor UO_1763 (O_1763,N_29921,N_29625);
and UO_1764 (O_1764,N_29920,N_29903);
or UO_1765 (O_1765,N_29937,N_29642);
nand UO_1766 (O_1766,N_29553,N_29664);
xnor UO_1767 (O_1767,N_29997,N_29972);
or UO_1768 (O_1768,N_29830,N_29919);
and UO_1769 (O_1769,N_29578,N_29590);
or UO_1770 (O_1770,N_29666,N_29500);
or UO_1771 (O_1771,N_29598,N_29671);
nand UO_1772 (O_1772,N_29584,N_29719);
xnor UO_1773 (O_1773,N_29845,N_29899);
xor UO_1774 (O_1774,N_29619,N_29612);
or UO_1775 (O_1775,N_29571,N_29682);
or UO_1776 (O_1776,N_29967,N_29826);
or UO_1777 (O_1777,N_29894,N_29706);
nand UO_1778 (O_1778,N_29660,N_29734);
nand UO_1779 (O_1779,N_29792,N_29961);
or UO_1780 (O_1780,N_29934,N_29945);
and UO_1781 (O_1781,N_29533,N_29949);
xor UO_1782 (O_1782,N_29810,N_29921);
and UO_1783 (O_1783,N_29565,N_29619);
and UO_1784 (O_1784,N_29932,N_29935);
and UO_1785 (O_1785,N_29941,N_29898);
nor UO_1786 (O_1786,N_29955,N_29985);
and UO_1787 (O_1787,N_29675,N_29718);
or UO_1788 (O_1788,N_29752,N_29543);
or UO_1789 (O_1789,N_29805,N_29942);
or UO_1790 (O_1790,N_29501,N_29755);
nor UO_1791 (O_1791,N_29746,N_29936);
or UO_1792 (O_1792,N_29521,N_29735);
and UO_1793 (O_1793,N_29618,N_29837);
and UO_1794 (O_1794,N_29951,N_29990);
xor UO_1795 (O_1795,N_29916,N_29894);
nand UO_1796 (O_1796,N_29780,N_29604);
xnor UO_1797 (O_1797,N_29744,N_29702);
nand UO_1798 (O_1798,N_29529,N_29890);
nand UO_1799 (O_1799,N_29752,N_29931);
xnor UO_1800 (O_1800,N_29526,N_29719);
nor UO_1801 (O_1801,N_29715,N_29834);
xor UO_1802 (O_1802,N_29921,N_29558);
nor UO_1803 (O_1803,N_29643,N_29855);
nand UO_1804 (O_1804,N_29593,N_29527);
or UO_1805 (O_1805,N_29543,N_29753);
xor UO_1806 (O_1806,N_29550,N_29892);
nor UO_1807 (O_1807,N_29684,N_29820);
nand UO_1808 (O_1808,N_29647,N_29782);
nand UO_1809 (O_1809,N_29728,N_29649);
and UO_1810 (O_1810,N_29967,N_29622);
nor UO_1811 (O_1811,N_29570,N_29565);
and UO_1812 (O_1812,N_29767,N_29585);
or UO_1813 (O_1813,N_29866,N_29535);
or UO_1814 (O_1814,N_29735,N_29725);
nand UO_1815 (O_1815,N_29997,N_29610);
xor UO_1816 (O_1816,N_29732,N_29547);
xnor UO_1817 (O_1817,N_29751,N_29594);
xnor UO_1818 (O_1818,N_29529,N_29935);
nor UO_1819 (O_1819,N_29874,N_29996);
and UO_1820 (O_1820,N_29614,N_29694);
or UO_1821 (O_1821,N_29920,N_29936);
or UO_1822 (O_1822,N_29580,N_29638);
nor UO_1823 (O_1823,N_29763,N_29512);
nand UO_1824 (O_1824,N_29884,N_29816);
or UO_1825 (O_1825,N_29919,N_29765);
and UO_1826 (O_1826,N_29814,N_29681);
nor UO_1827 (O_1827,N_29740,N_29576);
nor UO_1828 (O_1828,N_29789,N_29893);
and UO_1829 (O_1829,N_29513,N_29932);
nor UO_1830 (O_1830,N_29545,N_29792);
nor UO_1831 (O_1831,N_29728,N_29959);
or UO_1832 (O_1832,N_29877,N_29697);
or UO_1833 (O_1833,N_29817,N_29564);
nor UO_1834 (O_1834,N_29721,N_29838);
nor UO_1835 (O_1835,N_29528,N_29520);
or UO_1836 (O_1836,N_29891,N_29587);
or UO_1837 (O_1837,N_29848,N_29883);
xnor UO_1838 (O_1838,N_29827,N_29910);
and UO_1839 (O_1839,N_29659,N_29514);
xnor UO_1840 (O_1840,N_29849,N_29755);
and UO_1841 (O_1841,N_29768,N_29966);
xnor UO_1842 (O_1842,N_29848,N_29612);
xor UO_1843 (O_1843,N_29758,N_29719);
nand UO_1844 (O_1844,N_29925,N_29941);
and UO_1845 (O_1845,N_29647,N_29824);
and UO_1846 (O_1846,N_29929,N_29507);
and UO_1847 (O_1847,N_29687,N_29898);
nor UO_1848 (O_1848,N_29872,N_29936);
nor UO_1849 (O_1849,N_29547,N_29925);
nand UO_1850 (O_1850,N_29892,N_29805);
nand UO_1851 (O_1851,N_29658,N_29888);
nand UO_1852 (O_1852,N_29558,N_29816);
or UO_1853 (O_1853,N_29862,N_29608);
xnor UO_1854 (O_1854,N_29780,N_29763);
or UO_1855 (O_1855,N_29647,N_29735);
or UO_1856 (O_1856,N_29938,N_29695);
xnor UO_1857 (O_1857,N_29726,N_29836);
nand UO_1858 (O_1858,N_29629,N_29816);
or UO_1859 (O_1859,N_29573,N_29502);
nor UO_1860 (O_1860,N_29689,N_29904);
or UO_1861 (O_1861,N_29592,N_29746);
nand UO_1862 (O_1862,N_29932,N_29677);
nor UO_1863 (O_1863,N_29567,N_29806);
xnor UO_1864 (O_1864,N_29560,N_29541);
nand UO_1865 (O_1865,N_29696,N_29723);
nor UO_1866 (O_1866,N_29754,N_29770);
and UO_1867 (O_1867,N_29839,N_29835);
or UO_1868 (O_1868,N_29716,N_29569);
xor UO_1869 (O_1869,N_29698,N_29589);
nor UO_1870 (O_1870,N_29599,N_29806);
xnor UO_1871 (O_1871,N_29638,N_29834);
nand UO_1872 (O_1872,N_29992,N_29990);
nand UO_1873 (O_1873,N_29967,N_29825);
or UO_1874 (O_1874,N_29820,N_29812);
and UO_1875 (O_1875,N_29689,N_29673);
and UO_1876 (O_1876,N_29839,N_29860);
xor UO_1877 (O_1877,N_29719,N_29909);
nand UO_1878 (O_1878,N_29882,N_29811);
nor UO_1879 (O_1879,N_29727,N_29658);
or UO_1880 (O_1880,N_29829,N_29656);
or UO_1881 (O_1881,N_29791,N_29649);
nor UO_1882 (O_1882,N_29555,N_29504);
xor UO_1883 (O_1883,N_29872,N_29854);
nand UO_1884 (O_1884,N_29723,N_29655);
or UO_1885 (O_1885,N_29753,N_29505);
nor UO_1886 (O_1886,N_29562,N_29677);
nor UO_1887 (O_1887,N_29506,N_29929);
and UO_1888 (O_1888,N_29787,N_29519);
nor UO_1889 (O_1889,N_29744,N_29643);
nor UO_1890 (O_1890,N_29970,N_29581);
nand UO_1891 (O_1891,N_29539,N_29694);
xor UO_1892 (O_1892,N_29853,N_29558);
and UO_1893 (O_1893,N_29799,N_29740);
xor UO_1894 (O_1894,N_29649,N_29534);
xnor UO_1895 (O_1895,N_29655,N_29712);
nor UO_1896 (O_1896,N_29984,N_29620);
xnor UO_1897 (O_1897,N_29626,N_29670);
nor UO_1898 (O_1898,N_29549,N_29833);
xor UO_1899 (O_1899,N_29858,N_29722);
nand UO_1900 (O_1900,N_29818,N_29848);
and UO_1901 (O_1901,N_29942,N_29643);
nor UO_1902 (O_1902,N_29984,N_29724);
nor UO_1903 (O_1903,N_29848,N_29905);
and UO_1904 (O_1904,N_29897,N_29834);
nand UO_1905 (O_1905,N_29667,N_29651);
nor UO_1906 (O_1906,N_29796,N_29683);
and UO_1907 (O_1907,N_29968,N_29950);
or UO_1908 (O_1908,N_29727,N_29659);
and UO_1909 (O_1909,N_29849,N_29585);
and UO_1910 (O_1910,N_29613,N_29839);
and UO_1911 (O_1911,N_29802,N_29636);
or UO_1912 (O_1912,N_29644,N_29758);
xor UO_1913 (O_1913,N_29770,N_29888);
xor UO_1914 (O_1914,N_29626,N_29683);
or UO_1915 (O_1915,N_29555,N_29629);
or UO_1916 (O_1916,N_29953,N_29640);
or UO_1917 (O_1917,N_29747,N_29567);
nor UO_1918 (O_1918,N_29684,N_29993);
nand UO_1919 (O_1919,N_29648,N_29539);
nor UO_1920 (O_1920,N_29745,N_29859);
nor UO_1921 (O_1921,N_29817,N_29621);
and UO_1922 (O_1922,N_29720,N_29968);
and UO_1923 (O_1923,N_29869,N_29695);
nand UO_1924 (O_1924,N_29775,N_29757);
nand UO_1925 (O_1925,N_29913,N_29911);
nand UO_1926 (O_1926,N_29984,N_29679);
xnor UO_1927 (O_1927,N_29883,N_29748);
nand UO_1928 (O_1928,N_29834,N_29925);
or UO_1929 (O_1929,N_29999,N_29832);
nor UO_1930 (O_1930,N_29784,N_29527);
xor UO_1931 (O_1931,N_29564,N_29862);
nand UO_1932 (O_1932,N_29914,N_29883);
and UO_1933 (O_1933,N_29619,N_29747);
and UO_1934 (O_1934,N_29862,N_29755);
or UO_1935 (O_1935,N_29581,N_29575);
nand UO_1936 (O_1936,N_29561,N_29576);
and UO_1937 (O_1937,N_29606,N_29653);
xnor UO_1938 (O_1938,N_29968,N_29802);
nand UO_1939 (O_1939,N_29729,N_29508);
or UO_1940 (O_1940,N_29812,N_29744);
nor UO_1941 (O_1941,N_29733,N_29585);
and UO_1942 (O_1942,N_29910,N_29721);
or UO_1943 (O_1943,N_29737,N_29520);
or UO_1944 (O_1944,N_29917,N_29925);
nor UO_1945 (O_1945,N_29786,N_29701);
nand UO_1946 (O_1946,N_29626,N_29649);
nand UO_1947 (O_1947,N_29572,N_29749);
nand UO_1948 (O_1948,N_29655,N_29996);
and UO_1949 (O_1949,N_29666,N_29850);
nor UO_1950 (O_1950,N_29750,N_29970);
and UO_1951 (O_1951,N_29869,N_29840);
xor UO_1952 (O_1952,N_29901,N_29808);
nand UO_1953 (O_1953,N_29692,N_29669);
nor UO_1954 (O_1954,N_29999,N_29794);
and UO_1955 (O_1955,N_29808,N_29926);
or UO_1956 (O_1956,N_29652,N_29839);
and UO_1957 (O_1957,N_29708,N_29669);
xnor UO_1958 (O_1958,N_29730,N_29612);
nand UO_1959 (O_1959,N_29670,N_29937);
nand UO_1960 (O_1960,N_29573,N_29596);
xor UO_1961 (O_1961,N_29835,N_29674);
nor UO_1962 (O_1962,N_29884,N_29875);
nand UO_1963 (O_1963,N_29706,N_29830);
and UO_1964 (O_1964,N_29965,N_29988);
nand UO_1965 (O_1965,N_29671,N_29697);
nor UO_1966 (O_1966,N_29598,N_29991);
nand UO_1967 (O_1967,N_29807,N_29654);
or UO_1968 (O_1968,N_29563,N_29873);
nor UO_1969 (O_1969,N_29894,N_29674);
xor UO_1970 (O_1970,N_29675,N_29507);
or UO_1971 (O_1971,N_29754,N_29800);
xor UO_1972 (O_1972,N_29751,N_29605);
or UO_1973 (O_1973,N_29840,N_29619);
and UO_1974 (O_1974,N_29976,N_29860);
and UO_1975 (O_1975,N_29870,N_29542);
or UO_1976 (O_1976,N_29807,N_29788);
or UO_1977 (O_1977,N_29941,N_29908);
or UO_1978 (O_1978,N_29900,N_29655);
and UO_1979 (O_1979,N_29859,N_29800);
nand UO_1980 (O_1980,N_29976,N_29891);
nand UO_1981 (O_1981,N_29538,N_29595);
and UO_1982 (O_1982,N_29713,N_29572);
nand UO_1983 (O_1983,N_29829,N_29989);
and UO_1984 (O_1984,N_29847,N_29988);
nand UO_1985 (O_1985,N_29579,N_29500);
and UO_1986 (O_1986,N_29534,N_29758);
nor UO_1987 (O_1987,N_29618,N_29680);
xor UO_1988 (O_1988,N_29819,N_29934);
and UO_1989 (O_1989,N_29613,N_29644);
or UO_1990 (O_1990,N_29935,N_29659);
nor UO_1991 (O_1991,N_29981,N_29649);
xnor UO_1992 (O_1992,N_29861,N_29541);
and UO_1993 (O_1993,N_29528,N_29929);
nand UO_1994 (O_1994,N_29945,N_29988);
nand UO_1995 (O_1995,N_29658,N_29620);
nor UO_1996 (O_1996,N_29606,N_29690);
or UO_1997 (O_1997,N_29588,N_29873);
and UO_1998 (O_1998,N_29708,N_29737);
nand UO_1999 (O_1999,N_29571,N_29839);
or UO_2000 (O_2000,N_29758,N_29901);
nand UO_2001 (O_2001,N_29650,N_29646);
or UO_2002 (O_2002,N_29634,N_29875);
nand UO_2003 (O_2003,N_29557,N_29933);
or UO_2004 (O_2004,N_29802,N_29765);
and UO_2005 (O_2005,N_29954,N_29596);
nor UO_2006 (O_2006,N_29722,N_29919);
or UO_2007 (O_2007,N_29687,N_29889);
or UO_2008 (O_2008,N_29916,N_29594);
and UO_2009 (O_2009,N_29542,N_29637);
nand UO_2010 (O_2010,N_29662,N_29811);
xnor UO_2011 (O_2011,N_29994,N_29675);
nor UO_2012 (O_2012,N_29857,N_29700);
and UO_2013 (O_2013,N_29999,N_29922);
xnor UO_2014 (O_2014,N_29922,N_29994);
and UO_2015 (O_2015,N_29718,N_29961);
or UO_2016 (O_2016,N_29553,N_29973);
nor UO_2017 (O_2017,N_29661,N_29866);
xor UO_2018 (O_2018,N_29762,N_29884);
or UO_2019 (O_2019,N_29649,N_29874);
xor UO_2020 (O_2020,N_29531,N_29765);
nor UO_2021 (O_2021,N_29980,N_29892);
nand UO_2022 (O_2022,N_29754,N_29818);
xor UO_2023 (O_2023,N_29911,N_29890);
nor UO_2024 (O_2024,N_29963,N_29913);
or UO_2025 (O_2025,N_29729,N_29600);
and UO_2026 (O_2026,N_29680,N_29947);
and UO_2027 (O_2027,N_29645,N_29550);
nand UO_2028 (O_2028,N_29699,N_29943);
or UO_2029 (O_2029,N_29648,N_29980);
xor UO_2030 (O_2030,N_29680,N_29758);
and UO_2031 (O_2031,N_29706,N_29575);
and UO_2032 (O_2032,N_29882,N_29505);
or UO_2033 (O_2033,N_29746,N_29821);
and UO_2034 (O_2034,N_29986,N_29996);
nor UO_2035 (O_2035,N_29667,N_29680);
nand UO_2036 (O_2036,N_29625,N_29873);
or UO_2037 (O_2037,N_29637,N_29880);
or UO_2038 (O_2038,N_29673,N_29544);
nor UO_2039 (O_2039,N_29533,N_29837);
and UO_2040 (O_2040,N_29519,N_29610);
xnor UO_2041 (O_2041,N_29726,N_29635);
nand UO_2042 (O_2042,N_29847,N_29804);
or UO_2043 (O_2043,N_29978,N_29810);
xor UO_2044 (O_2044,N_29844,N_29971);
and UO_2045 (O_2045,N_29717,N_29741);
nor UO_2046 (O_2046,N_29543,N_29776);
and UO_2047 (O_2047,N_29869,N_29770);
xor UO_2048 (O_2048,N_29671,N_29605);
nor UO_2049 (O_2049,N_29602,N_29833);
and UO_2050 (O_2050,N_29902,N_29646);
xor UO_2051 (O_2051,N_29994,N_29838);
xor UO_2052 (O_2052,N_29899,N_29659);
or UO_2053 (O_2053,N_29543,N_29555);
and UO_2054 (O_2054,N_29507,N_29761);
xnor UO_2055 (O_2055,N_29830,N_29918);
and UO_2056 (O_2056,N_29556,N_29836);
or UO_2057 (O_2057,N_29727,N_29505);
and UO_2058 (O_2058,N_29788,N_29972);
and UO_2059 (O_2059,N_29616,N_29675);
nor UO_2060 (O_2060,N_29969,N_29649);
nand UO_2061 (O_2061,N_29694,N_29758);
nor UO_2062 (O_2062,N_29534,N_29708);
and UO_2063 (O_2063,N_29771,N_29837);
xnor UO_2064 (O_2064,N_29773,N_29688);
nand UO_2065 (O_2065,N_29576,N_29759);
or UO_2066 (O_2066,N_29823,N_29725);
nor UO_2067 (O_2067,N_29646,N_29921);
and UO_2068 (O_2068,N_29776,N_29832);
or UO_2069 (O_2069,N_29727,N_29750);
nor UO_2070 (O_2070,N_29912,N_29757);
and UO_2071 (O_2071,N_29514,N_29761);
nor UO_2072 (O_2072,N_29907,N_29727);
and UO_2073 (O_2073,N_29621,N_29763);
nand UO_2074 (O_2074,N_29583,N_29598);
xor UO_2075 (O_2075,N_29996,N_29876);
nand UO_2076 (O_2076,N_29816,N_29913);
and UO_2077 (O_2077,N_29763,N_29702);
nor UO_2078 (O_2078,N_29560,N_29589);
nand UO_2079 (O_2079,N_29635,N_29757);
nand UO_2080 (O_2080,N_29631,N_29989);
xnor UO_2081 (O_2081,N_29706,N_29975);
and UO_2082 (O_2082,N_29589,N_29714);
nor UO_2083 (O_2083,N_29806,N_29550);
and UO_2084 (O_2084,N_29709,N_29658);
or UO_2085 (O_2085,N_29546,N_29841);
nand UO_2086 (O_2086,N_29633,N_29590);
nor UO_2087 (O_2087,N_29835,N_29885);
nand UO_2088 (O_2088,N_29976,N_29660);
nand UO_2089 (O_2089,N_29660,N_29910);
or UO_2090 (O_2090,N_29530,N_29612);
nor UO_2091 (O_2091,N_29672,N_29659);
xnor UO_2092 (O_2092,N_29567,N_29870);
or UO_2093 (O_2093,N_29719,N_29827);
nor UO_2094 (O_2094,N_29637,N_29704);
xnor UO_2095 (O_2095,N_29879,N_29932);
or UO_2096 (O_2096,N_29530,N_29749);
and UO_2097 (O_2097,N_29986,N_29987);
nor UO_2098 (O_2098,N_29801,N_29834);
or UO_2099 (O_2099,N_29796,N_29648);
or UO_2100 (O_2100,N_29725,N_29609);
nand UO_2101 (O_2101,N_29664,N_29505);
xor UO_2102 (O_2102,N_29733,N_29531);
or UO_2103 (O_2103,N_29928,N_29600);
and UO_2104 (O_2104,N_29991,N_29885);
nand UO_2105 (O_2105,N_29573,N_29944);
nor UO_2106 (O_2106,N_29913,N_29720);
nor UO_2107 (O_2107,N_29580,N_29509);
nand UO_2108 (O_2108,N_29613,N_29941);
nand UO_2109 (O_2109,N_29644,N_29847);
and UO_2110 (O_2110,N_29748,N_29818);
nand UO_2111 (O_2111,N_29698,N_29859);
nor UO_2112 (O_2112,N_29742,N_29781);
xor UO_2113 (O_2113,N_29741,N_29581);
nand UO_2114 (O_2114,N_29849,N_29509);
and UO_2115 (O_2115,N_29722,N_29501);
or UO_2116 (O_2116,N_29763,N_29559);
nand UO_2117 (O_2117,N_29803,N_29788);
or UO_2118 (O_2118,N_29685,N_29517);
or UO_2119 (O_2119,N_29689,N_29785);
nor UO_2120 (O_2120,N_29592,N_29587);
nand UO_2121 (O_2121,N_29866,N_29983);
or UO_2122 (O_2122,N_29833,N_29544);
nor UO_2123 (O_2123,N_29546,N_29726);
xnor UO_2124 (O_2124,N_29928,N_29693);
nand UO_2125 (O_2125,N_29664,N_29972);
and UO_2126 (O_2126,N_29829,N_29551);
and UO_2127 (O_2127,N_29552,N_29729);
nor UO_2128 (O_2128,N_29821,N_29799);
nor UO_2129 (O_2129,N_29864,N_29693);
or UO_2130 (O_2130,N_29870,N_29817);
nand UO_2131 (O_2131,N_29888,N_29790);
or UO_2132 (O_2132,N_29887,N_29552);
or UO_2133 (O_2133,N_29735,N_29698);
or UO_2134 (O_2134,N_29706,N_29909);
xor UO_2135 (O_2135,N_29553,N_29590);
xnor UO_2136 (O_2136,N_29927,N_29506);
or UO_2137 (O_2137,N_29570,N_29552);
and UO_2138 (O_2138,N_29656,N_29862);
xor UO_2139 (O_2139,N_29734,N_29737);
nor UO_2140 (O_2140,N_29882,N_29540);
nand UO_2141 (O_2141,N_29627,N_29767);
or UO_2142 (O_2142,N_29821,N_29918);
or UO_2143 (O_2143,N_29808,N_29795);
and UO_2144 (O_2144,N_29932,N_29647);
or UO_2145 (O_2145,N_29671,N_29729);
nand UO_2146 (O_2146,N_29804,N_29720);
nor UO_2147 (O_2147,N_29992,N_29613);
and UO_2148 (O_2148,N_29823,N_29818);
or UO_2149 (O_2149,N_29533,N_29978);
and UO_2150 (O_2150,N_29911,N_29633);
and UO_2151 (O_2151,N_29841,N_29849);
nand UO_2152 (O_2152,N_29792,N_29679);
nand UO_2153 (O_2153,N_29894,N_29915);
nor UO_2154 (O_2154,N_29678,N_29830);
or UO_2155 (O_2155,N_29760,N_29548);
or UO_2156 (O_2156,N_29821,N_29690);
xor UO_2157 (O_2157,N_29875,N_29564);
or UO_2158 (O_2158,N_29811,N_29762);
xor UO_2159 (O_2159,N_29961,N_29632);
nor UO_2160 (O_2160,N_29503,N_29746);
and UO_2161 (O_2161,N_29650,N_29942);
and UO_2162 (O_2162,N_29894,N_29621);
nor UO_2163 (O_2163,N_29581,N_29871);
or UO_2164 (O_2164,N_29923,N_29640);
and UO_2165 (O_2165,N_29811,N_29742);
xor UO_2166 (O_2166,N_29808,N_29861);
xor UO_2167 (O_2167,N_29728,N_29502);
xor UO_2168 (O_2168,N_29768,N_29515);
nand UO_2169 (O_2169,N_29747,N_29740);
nand UO_2170 (O_2170,N_29617,N_29562);
and UO_2171 (O_2171,N_29631,N_29934);
nand UO_2172 (O_2172,N_29851,N_29616);
and UO_2173 (O_2173,N_29856,N_29672);
nand UO_2174 (O_2174,N_29523,N_29600);
nand UO_2175 (O_2175,N_29871,N_29718);
and UO_2176 (O_2176,N_29525,N_29632);
xor UO_2177 (O_2177,N_29658,N_29549);
and UO_2178 (O_2178,N_29785,N_29609);
or UO_2179 (O_2179,N_29782,N_29853);
nor UO_2180 (O_2180,N_29670,N_29962);
and UO_2181 (O_2181,N_29763,N_29927);
or UO_2182 (O_2182,N_29599,N_29852);
and UO_2183 (O_2183,N_29589,N_29699);
and UO_2184 (O_2184,N_29913,N_29508);
xnor UO_2185 (O_2185,N_29957,N_29542);
xnor UO_2186 (O_2186,N_29859,N_29820);
nor UO_2187 (O_2187,N_29635,N_29689);
nand UO_2188 (O_2188,N_29974,N_29816);
nand UO_2189 (O_2189,N_29620,N_29827);
nor UO_2190 (O_2190,N_29588,N_29911);
and UO_2191 (O_2191,N_29724,N_29983);
nand UO_2192 (O_2192,N_29740,N_29528);
nor UO_2193 (O_2193,N_29567,N_29575);
or UO_2194 (O_2194,N_29507,N_29821);
nand UO_2195 (O_2195,N_29799,N_29716);
xnor UO_2196 (O_2196,N_29523,N_29939);
xnor UO_2197 (O_2197,N_29761,N_29909);
and UO_2198 (O_2198,N_29856,N_29779);
and UO_2199 (O_2199,N_29947,N_29585);
or UO_2200 (O_2200,N_29585,N_29978);
xor UO_2201 (O_2201,N_29515,N_29506);
nor UO_2202 (O_2202,N_29663,N_29953);
or UO_2203 (O_2203,N_29811,N_29773);
xor UO_2204 (O_2204,N_29721,N_29598);
xnor UO_2205 (O_2205,N_29679,N_29999);
nor UO_2206 (O_2206,N_29856,N_29686);
xor UO_2207 (O_2207,N_29978,N_29725);
or UO_2208 (O_2208,N_29850,N_29674);
and UO_2209 (O_2209,N_29959,N_29946);
nor UO_2210 (O_2210,N_29712,N_29874);
or UO_2211 (O_2211,N_29500,N_29817);
xnor UO_2212 (O_2212,N_29831,N_29855);
nand UO_2213 (O_2213,N_29905,N_29666);
or UO_2214 (O_2214,N_29919,N_29859);
xor UO_2215 (O_2215,N_29640,N_29977);
nor UO_2216 (O_2216,N_29952,N_29699);
or UO_2217 (O_2217,N_29863,N_29568);
xnor UO_2218 (O_2218,N_29830,N_29846);
or UO_2219 (O_2219,N_29787,N_29539);
and UO_2220 (O_2220,N_29934,N_29619);
nand UO_2221 (O_2221,N_29602,N_29783);
or UO_2222 (O_2222,N_29937,N_29720);
nand UO_2223 (O_2223,N_29509,N_29746);
nor UO_2224 (O_2224,N_29898,N_29657);
and UO_2225 (O_2225,N_29863,N_29671);
nor UO_2226 (O_2226,N_29734,N_29511);
nor UO_2227 (O_2227,N_29927,N_29778);
xor UO_2228 (O_2228,N_29548,N_29936);
xnor UO_2229 (O_2229,N_29547,N_29954);
nor UO_2230 (O_2230,N_29823,N_29997);
and UO_2231 (O_2231,N_29886,N_29805);
nor UO_2232 (O_2232,N_29591,N_29879);
xor UO_2233 (O_2233,N_29523,N_29875);
and UO_2234 (O_2234,N_29826,N_29595);
nor UO_2235 (O_2235,N_29715,N_29811);
and UO_2236 (O_2236,N_29927,N_29767);
nor UO_2237 (O_2237,N_29858,N_29681);
and UO_2238 (O_2238,N_29582,N_29829);
nor UO_2239 (O_2239,N_29527,N_29979);
xor UO_2240 (O_2240,N_29917,N_29829);
xnor UO_2241 (O_2241,N_29713,N_29521);
nand UO_2242 (O_2242,N_29565,N_29569);
nor UO_2243 (O_2243,N_29755,N_29616);
xnor UO_2244 (O_2244,N_29707,N_29517);
and UO_2245 (O_2245,N_29725,N_29624);
nor UO_2246 (O_2246,N_29843,N_29589);
or UO_2247 (O_2247,N_29617,N_29877);
xor UO_2248 (O_2248,N_29571,N_29881);
nand UO_2249 (O_2249,N_29650,N_29672);
xnor UO_2250 (O_2250,N_29688,N_29746);
nor UO_2251 (O_2251,N_29621,N_29945);
or UO_2252 (O_2252,N_29716,N_29746);
nor UO_2253 (O_2253,N_29713,N_29633);
and UO_2254 (O_2254,N_29564,N_29840);
or UO_2255 (O_2255,N_29985,N_29863);
and UO_2256 (O_2256,N_29529,N_29940);
or UO_2257 (O_2257,N_29813,N_29675);
nand UO_2258 (O_2258,N_29761,N_29813);
nand UO_2259 (O_2259,N_29801,N_29910);
nand UO_2260 (O_2260,N_29587,N_29768);
and UO_2261 (O_2261,N_29971,N_29612);
or UO_2262 (O_2262,N_29553,N_29855);
or UO_2263 (O_2263,N_29974,N_29517);
nand UO_2264 (O_2264,N_29749,N_29533);
xor UO_2265 (O_2265,N_29661,N_29897);
nand UO_2266 (O_2266,N_29824,N_29571);
and UO_2267 (O_2267,N_29553,N_29635);
or UO_2268 (O_2268,N_29714,N_29603);
xor UO_2269 (O_2269,N_29708,N_29801);
and UO_2270 (O_2270,N_29673,N_29894);
nand UO_2271 (O_2271,N_29732,N_29915);
or UO_2272 (O_2272,N_29550,N_29543);
or UO_2273 (O_2273,N_29527,N_29626);
nand UO_2274 (O_2274,N_29643,N_29521);
xor UO_2275 (O_2275,N_29950,N_29613);
nand UO_2276 (O_2276,N_29910,N_29896);
nand UO_2277 (O_2277,N_29985,N_29680);
or UO_2278 (O_2278,N_29920,N_29884);
nor UO_2279 (O_2279,N_29531,N_29646);
nand UO_2280 (O_2280,N_29809,N_29523);
or UO_2281 (O_2281,N_29949,N_29954);
and UO_2282 (O_2282,N_29792,N_29716);
xnor UO_2283 (O_2283,N_29827,N_29559);
xor UO_2284 (O_2284,N_29834,N_29900);
xor UO_2285 (O_2285,N_29593,N_29673);
xnor UO_2286 (O_2286,N_29732,N_29534);
xor UO_2287 (O_2287,N_29961,N_29769);
nor UO_2288 (O_2288,N_29828,N_29640);
or UO_2289 (O_2289,N_29512,N_29744);
nor UO_2290 (O_2290,N_29820,N_29923);
xnor UO_2291 (O_2291,N_29712,N_29766);
and UO_2292 (O_2292,N_29729,N_29740);
nor UO_2293 (O_2293,N_29682,N_29689);
xor UO_2294 (O_2294,N_29649,N_29524);
xnor UO_2295 (O_2295,N_29600,N_29973);
and UO_2296 (O_2296,N_29767,N_29837);
or UO_2297 (O_2297,N_29616,N_29994);
or UO_2298 (O_2298,N_29781,N_29684);
and UO_2299 (O_2299,N_29948,N_29739);
or UO_2300 (O_2300,N_29728,N_29635);
xor UO_2301 (O_2301,N_29597,N_29755);
xnor UO_2302 (O_2302,N_29738,N_29824);
nor UO_2303 (O_2303,N_29655,N_29914);
nand UO_2304 (O_2304,N_29753,N_29791);
or UO_2305 (O_2305,N_29966,N_29945);
xnor UO_2306 (O_2306,N_29800,N_29807);
and UO_2307 (O_2307,N_29572,N_29537);
or UO_2308 (O_2308,N_29853,N_29794);
and UO_2309 (O_2309,N_29600,N_29550);
nor UO_2310 (O_2310,N_29768,N_29566);
nor UO_2311 (O_2311,N_29872,N_29821);
nand UO_2312 (O_2312,N_29614,N_29615);
or UO_2313 (O_2313,N_29915,N_29998);
nand UO_2314 (O_2314,N_29873,N_29918);
or UO_2315 (O_2315,N_29685,N_29992);
nor UO_2316 (O_2316,N_29604,N_29918);
and UO_2317 (O_2317,N_29503,N_29901);
and UO_2318 (O_2318,N_29559,N_29728);
or UO_2319 (O_2319,N_29684,N_29875);
nor UO_2320 (O_2320,N_29583,N_29828);
nor UO_2321 (O_2321,N_29893,N_29724);
nand UO_2322 (O_2322,N_29974,N_29514);
nor UO_2323 (O_2323,N_29501,N_29903);
nand UO_2324 (O_2324,N_29731,N_29534);
xnor UO_2325 (O_2325,N_29586,N_29877);
nand UO_2326 (O_2326,N_29706,N_29517);
or UO_2327 (O_2327,N_29823,N_29708);
xnor UO_2328 (O_2328,N_29801,N_29709);
and UO_2329 (O_2329,N_29993,N_29934);
xor UO_2330 (O_2330,N_29520,N_29957);
nor UO_2331 (O_2331,N_29810,N_29544);
nand UO_2332 (O_2332,N_29955,N_29935);
xnor UO_2333 (O_2333,N_29530,N_29894);
nand UO_2334 (O_2334,N_29500,N_29509);
nor UO_2335 (O_2335,N_29588,N_29535);
xnor UO_2336 (O_2336,N_29832,N_29727);
nand UO_2337 (O_2337,N_29541,N_29846);
nor UO_2338 (O_2338,N_29635,N_29664);
or UO_2339 (O_2339,N_29570,N_29544);
or UO_2340 (O_2340,N_29591,N_29614);
nand UO_2341 (O_2341,N_29817,N_29848);
nor UO_2342 (O_2342,N_29674,N_29959);
and UO_2343 (O_2343,N_29959,N_29853);
xor UO_2344 (O_2344,N_29648,N_29869);
nand UO_2345 (O_2345,N_29755,N_29921);
or UO_2346 (O_2346,N_29572,N_29739);
nand UO_2347 (O_2347,N_29662,N_29569);
nand UO_2348 (O_2348,N_29934,N_29826);
nor UO_2349 (O_2349,N_29625,N_29934);
xor UO_2350 (O_2350,N_29568,N_29870);
or UO_2351 (O_2351,N_29983,N_29640);
and UO_2352 (O_2352,N_29524,N_29519);
xor UO_2353 (O_2353,N_29867,N_29606);
and UO_2354 (O_2354,N_29800,N_29840);
nand UO_2355 (O_2355,N_29598,N_29924);
xnor UO_2356 (O_2356,N_29956,N_29793);
xor UO_2357 (O_2357,N_29666,N_29627);
or UO_2358 (O_2358,N_29755,N_29689);
and UO_2359 (O_2359,N_29680,N_29656);
nor UO_2360 (O_2360,N_29942,N_29639);
and UO_2361 (O_2361,N_29939,N_29978);
nand UO_2362 (O_2362,N_29765,N_29876);
nor UO_2363 (O_2363,N_29502,N_29669);
nand UO_2364 (O_2364,N_29671,N_29655);
and UO_2365 (O_2365,N_29855,N_29719);
or UO_2366 (O_2366,N_29871,N_29539);
and UO_2367 (O_2367,N_29977,N_29891);
or UO_2368 (O_2368,N_29696,N_29822);
xor UO_2369 (O_2369,N_29633,N_29533);
or UO_2370 (O_2370,N_29902,N_29674);
xnor UO_2371 (O_2371,N_29715,N_29779);
nand UO_2372 (O_2372,N_29863,N_29707);
and UO_2373 (O_2373,N_29574,N_29545);
or UO_2374 (O_2374,N_29730,N_29507);
xor UO_2375 (O_2375,N_29649,N_29590);
or UO_2376 (O_2376,N_29940,N_29770);
nand UO_2377 (O_2377,N_29671,N_29905);
or UO_2378 (O_2378,N_29548,N_29747);
nor UO_2379 (O_2379,N_29804,N_29973);
nor UO_2380 (O_2380,N_29722,N_29721);
xnor UO_2381 (O_2381,N_29873,N_29583);
or UO_2382 (O_2382,N_29790,N_29839);
xor UO_2383 (O_2383,N_29745,N_29833);
and UO_2384 (O_2384,N_29537,N_29980);
xnor UO_2385 (O_2385,N_29687,N_29949);
nand UO_2386 (O_2386,N_29662,N_29555);
nor UO_2387 (O_2387,N_29849,N_29975);
and UO_2388 (O_2388,N_29998,N_29696);
nand UO_2389 (O_2389,N_29505,N_29555);
and UO_2390 (O_2390,N_29967,N_29520);
and UO_2391 (O_2391,N_29544,N_29766);
and UO_2392 (O_2392,N_29936,N_29768);
or UO_2393 (O_2393,N_29935,N_29964);
and UO_2394 (O_2394,N_29702,N_29889);
nor UO_2395 (O_2395,N_29730,N_29948);
nand UO_2396 (O_2396,N_29989,N_29993);
xor UO_2397 (O_2397,N_29826,N_29738);
xnor UO_2398 (O_2398,N_29538,N_29654);
xnor UO_2399 (O_2399,N_29825,N_29760);
nor UO_2400 (O_2400,N_29584,N_29522);
and UO_2401 (O_2401,N_29640,N_29773);
and UO_2402 (O_2402,N_29761,N_29674);
and UO_2403 (O_2403,N_29820,N_29532);
nand UO_2404 (O_2404,N_29557,N_29728);
xor UO_2405 (O_2405,N_29802,N_29668);
or UO_2406 (O_2406,N_29782,N_29699);
nor UO_2407 (O_2407,N_29961,N_29651);
xnor UO_2408 (O_2408,N_29649,N_29757);
nand UO_2409 (O_2409,N_29655,N_29843);
or UO_2410 (O_2410,N_29550,N_29609);
nand UO_2411 (O_2411,N_29911,N_29800);
or UO_2412 (O_2412,N_29518,N_29580);
and UO_2413 (O_2413,N_29765,N_29882);
nor UO_2414 (O_2414,N_29919,N_29950);
and UO_2415 (O_2415,N_29928,N_29984);
nand UO_2416 (O_2416,N_29607,N_29935);
xor UO_2417 (O_2417,N_29584,N_29552);
xnor UO_2418 (O_2418,N_29996,N_29871);
nand UO_2419 (O_2419,N_29525,N_29802);
or UO_2420 (O_2420,N_29864,N_29927);
xor UO_2421 (O_2421,N_29996,N_29559);
nand UO_2422 (O_2422,N_29723,N_29990);
or UO_2423 (O_2423,N_29614,N_29999);
nor UO_2424 (O_2424,N_29928,N_29792);
xor UO_2425 (O_2425,N_29974,N_29607);
nand UO_2426 (O_2426,N_29665,N_29934);
nand UO_2427 (O_2427,N_29955,N_29790);
nor UO_2428 (O_2428,N_29666,N_29963);
and UO_2429 (O_2429,N_29774,N_29717);
nor UO_2430 (O_2430,N_29562,N_29825);
xnor UO_2431 (O_2431,N_29577,N_29643);
xnor UO_2432 (O_2432,N_29812,N_29698);
nand UO_2433 (O_2433,N_29836,N_29594);
xnor UO_2434 (O_2434,N_29704,N_29915);
nand UO_2435 (O_2435,N_29671,N_29831);
xnor UO_2436 (O_2436,N_29673,N_29700);
and UO_2437 (O_2437,N_29568,N_29506);
nand UO_2438 (O_2438,N_29922,N_29679);
nor UO_2439 (O_2439,N_29581,N_29894);
and UO_2440 (O_2440,N_29559,N_29895);
xnor UO_2441 (O_2441,N_29508,N_29665);
xor UO_2442 (O_2442,N_29936,N_29626);
nand UO_2443 (O_2443,N_29671,N_29725);
nor UO_2444 (O_2444,N_29870,N_29995);
and UO_2445 (O_2445,N_29787,N_29910);
and UO_2446 (O_2446,N_29681,N_29780);
nor UO_2447 (O_2447,N_29885,N_29855);
or UO_2448 (O_2448,N_29811,N_29698);
nand UO_2449 (O_2449,N_29633,N_29711);
xor UO_2450 (O_2450,N_29506,N_29917);
xnor UO_2451 (O_2451,N_29519,N_29982);
nand UO_2452 (O_2452,N_29651,N_29747);
nand UO_2453 (O_2453,N_29957,N_29608);
or UO_2454 (O_2454,N_29696,N_29849);
nor UO_2455 (O_2455,N_29553,N_29946);
or UO_2456 (O_2456,N_29814,N_29887);
nand UO_2457 (O_2457,N_29668,N_29987);
or UO_2458 (O_2458,N_29558,N_29758);
and UO_2459 (O_2459,N_29707,N_29939);
or UO_2460 (O_2460,N_29813,N_29731);
xnor UO_2461 (O_2461,N_29988,N_29575);
xor UO_2462 (O_2462,N_29546,N_29502);
nor UO_2463 (O_2463,N_29869,N_29685);
xor UO_2464 (O_2464,N_29943,N_29781);
and UO_2465 (O_2465,N_29665,N_29510);
and UO_2466 (O_2466,N_29697,N_29553);
nor UO_2467 (O_2467,N_29833,N_29865);
or UO_2468 (O_2468,N_29985,N_29625);
xor UO_2469 (O_2469,N_29824,N_29945);
nor UO_2470 (O_2470,N_29951,N_29579);
xnor UO_2471 (O_2471,N_29926,N_29566);
nor UO_2472 (O_2472,N_29642,N_29804);
nor UO_2473 (O_2473,N_29837,N_29987);
and UO_2474 (O_2474,N_29506,N_29797);
xnor UO_2475 (O_2475,N_29588,N_29819);
nand UO_2476 (O_2476,N_29741,N_29564);
nand UO_2477 (O_2477,N_29752,N_29609);
and UO_2478 (O_2478,N_29748,N_29507);
nand UO_2479 (O_2479,N_29957,N_29991);
nand UO_2480 (O_2480,N_29530,N_29982);
or UO_2481 (O_2481,N_29759,N_29689);
nand UO_2482 (O_2482,N_29927,N_29641);
nor UO_2483 (O_2483,N_29533,N_29852);
nor UO_2484 (O_2484,N_29750,N_29692);
xor UO_2485 (O_2485,N_29776,N_29996);
nor UO_2486 (O_2486,N_29759,N_29555);
or UO_2487 (O_2487,N_29922,N_29781);
or UO_2488 (O_2488,N_29650,N_29637);
xor UO_2489 (O_2489,N_29896,N_29523);
xnor UO_2490 (O_2490,N_29758,N_29743);
and UO_2491 (O_2491,N_29654,N_29810);
nor UO_2492 (O_2492,N_29874,N_29989);
nand UO_2493 (O_2493,N_29701,N_29667);
or UO_2494 (O_2494,N_29754,N_29955);
nor UO_2495 (O_2495,N_29817,N_29923);
xnor UO_2496 (O_2496,N_29932,N_29672);
nor UO_2497 (O_2497,N_29895,N_29911);
nand UO_2498 (O_2498,N_29925,N_29555);
or UO_2499 (O_2499,N_29999,N_29809);
and UO_2500 (O_2500,N_29572,N_29850);
and UO_2501 (O_2501,N_29918,N_29592);
nand UO_2502 (O_2502,N_29606,N_29973);
or UO_2503 (O_2503,N_29596,N_29551);
nor UO_2504 (O_2504,N_29971,N_29837);
xor UO_2505 (O_2505,N_29523,N_29573);
and UO_2506 (O_2506,N_29679,N_29935);
xnor UO_2507 (O_2507,N_29807,N_29870);
nand UO_2508 (O_2508,N_29603,N_29728);
nand UO_2509 (O_2509,N_29783,N_29514);
and UO_2510 (O_2510,N_29668,N_29568);
nor UO_2511 (O_2511,N_29697,N_29740);
nand UO_2512 (O_2512,N_29678,N_29635);
or UO_2513 (O_2513,N_29670,N_29963);
or UO_2514 (O_2514,N_29711,N_29831);
nand UO_2515 (O_2515,N_29797,N_29587);
xor UO_2516 (O_2516,N_29807,N_29574);
xor UO_2517 (O_2517,N_29751,N_29945);
or UO_2518 (O_2518,N_29568,N_29797);
nand UO_2519 (O_2519,N_29841,N_29836);
nor UO_2520 (O_2520,N_29611,N_29959);
nand UO_2521 (O_2521,N_29760,N_29614);
nor UO_2522 (O_2522,N_29945,N_29505);
nand UO_2523 (O_2523,N_29936,N_29584);
nor UO_2524 (O_2524,N_29911,N_29834);
and UO_2525 (O_2525,N_29736,N_29980);
nor UO_2526 (O_2526,N_29684,N_29595);
or UO_2527 (O_2527,N_29702,N_29965);
xor UO_2528 (O_2528,N_29617,N_29506);
nor UO_2529 (O_2529,N_29548,N_29851);
and UO_2530 (O_2530,N_29801,N_29505);
or UO_2531 (O_2531,N_29881,N_29560);
nand UO_2532 (O_2532,N_29943,N_29780);
xnor UO_2533 (O_2533,N_29528,N_29776);
and UO_2534 (O_2534,N_29779,N_29623);
or UO_2535 (O_2535,N_29821,N_29687);
nor UO_2536 (O_2536,N_29947,N_29944);
or UO_2537 (O_2537,N_29979,N_29552);
xor UO_2538 (O_2538,N_29660,N_29669);
or UO_2539 (O_2539,N_29968,N_29628);
and UO_2540 (O_2540,N_29522,N_29731);
xor UO_2541 (O_2541,N_29962,N_29752);
or UO_2542 (O_2542,N_29665,N_29927);
xor UO_2543 (O_2543,N_29549,N_29590);
nand UO_2544 (O_2544,N_29639,N_29796);
nor UO_2545 (O_2545,N_29699,N_29945);
xor UO_2546 (O_2546,N_29543,N_29788);
nor UO_2547 (O_2547,N_29532,N_29712);
nand UO_2548 (O_2548,N_29821,N_29893);
or UO_2549 (O_2549,N_29500,N_29588);
nor UO_2550 (O_2550,N_29724,N_29843);
and UO_2551 (O_2551,N_29847,N_29810);
nand UO_2552 (O_2552,N_29730,N_29932);
and UO_2553 (O_2553,N_29569,N_29505);
nand UO_2554 (O_2554,N_29659,N_29639);
xor UO_2555 (O_2555,N_29752,N_29762);
nand UO_2556 (O_2556,N_29711,N_29757);
xnor UO_2557 (O_2557,N_29843,N_29688);
nand UO_2558 (O_2558,N_29735,N_29957);
or UO_2559 (O_2559,N_29544,N_29610);
nand UO_2560 (O_2560,N_29548,N_29734);
or UO_2561 (O_2561,N_29786,N_29508);
nand UO_2562 (O_2562,N_29541,N_29936);
or UO_2563 (O_2563,N_29755,N_29761);
nand UO_2564 (O_2564,N_29558,N_29645);
or UO_2565 (O_2565,N_29679,N_29598);
and UO_2566 (O_2566,N_29661,N_29964);
xnor UO_2567 (O_2567,N_29876,N_29900);
nand UO_2568 (O_2568,N_29958,N_29941);
and UO_2569 (O_2569,N_29605,N_29766);
xnor UO_2570 (O_2570,N_29527,N_29511);
or UO_2571 (O_2571,N_29748,N_29919);
or UO_2572 (O_2572,N_29568,N_29762);
nor UO_2573 (O_2573,N_29853,N_29789);
xor UO_2574 (O_2574,N_29948,N_29630);
or UO_2575 (O_2575,N_29610,N_29831);
nor UO_2576 (O_2576,N_29526,N_29630);
nor UO_2577 (O_2577,N_29859,N_29778);
xor UO_2578 (O_2578,N_29845,N_29561);
nor UO_2579 (O_2579,N_29918,N_29694);
nand UO_2580 (O_2580,N_29752,N_29527);
nor UO_2581 (O_2581,N_29539,N_29782);
nor UO_2582 (O_2582,N_29880,N_29759);
nand UO_2583 (O_2583,N_29957,N_29533);
nand UO_2584 (O_2584,N_29987,N_29640);
nor UO_2585 (O_2585,N_29924,N_29983);
nand UO_2586 (O_2586,N_29546,N_29957);
xor UO_2587 (O_2587,N_29850,N_29632);
nand UO_2588 (O_2588,N_29732,N_29876);
and UO_2589 (O_2589,N_29725,N_29660);
nand UO_2590 (O_2590,N_29943,N_29763);
or UO_2591 (O_2591,N_29652,N_29820);
nand UO_2592 (O_2592,N_29893,N_29986);
and UO_2593 (O_2593,N_29838,N_29761);
xor UO_2594 (O_2594,N_29760,N_29725);
and UO_2595 (O_2595,N_29516,N_29672);
nand UO_2596 (O_2596,N_29541,N_29941);
nor UO_2597 (O_2597,N_29775,N_29870);
and UO_2598 (O_2598,N_29716,N_29522);
xor UO_2599 (O_2599,N_29925,N_29645);
nand UO_2600 (O_2600,N_29978,N_29715);
xnor UO_2601 (O_2601,N_29893,N_29590);
nand UO_2602 (O_2602,N_29854,N_29564);
xnor UO_2603 (O_2603,N_29978,N_29658);
xor UO_2604 (O_2604,N_29870,N_29825);
or UO_2605 (O_2605,N_29891,N_29557);
xnor UO_2606 (O_2606,N_29669,N_29702);
or UO_2607 (O_2607,N_29637,N_29944);
or UO_2608 (O_2608,N_29830,N_29946);
xor UO_2609 (O_2609,N_29870,N_29684);
nand UO_2610 (O_2610,N_29859,N_29829);
nor UO_2611 (O_2611,N_29645,N_29509);
nor UO_2612 (O_2612,N_29748,N_29524);
nor UO_2613 (O_2613,N_29844,N_29830);
nand UO_2614 (O_2614,N_29584,N_29998);
nand UO_2615 (O_2615,N_29801,N_29972);
or UO_2616 (O_2616,N_29528,N_29801);
xnor UO_2617 (O_2617,N_29871,N_29832);
nand UO_2618 (O_2618,N_29731,N_29516);
nor UO_2619 (O_2619,N_29643,N_29967);
nand UO_2620 (O_2620,N_29992,N_29945);
and UO_2621 (O_2621,N_29874,N_29565);
or UO_2622 (O_2622,N_29935,N_29999);
and UO_2623 (O_2623,N_29515,N_29942);
or UO_2624 (O_2624,N_29941,N_29584);
and UO_2625 (O_2625,N_29711,N_29576);
nor UO_2626 (O_2626,N_29921,N_29797);
or UO_2627 (O_2627,N_29793,N_29540);
and UO_2628 (O_2628,N_29929,N_29736);
nor UO_2629 (O_2629,N_29928,N_29507);
and UO_2630 (O_2630,N_29899,N_29590);
xnor UO_2631 (O_2631,N_29622,N_29653);
and UO_2632 (O_2632,N_29659,N_29521);
or UO_2633 (O_2633,N_29767,N_29851);
and UO_2634 (O_2634,N_29830,N_29788);
and UO_2635 (O_2635,N_29592,N_29699);
and UO_2636 (O_2636,N_29746,N_29725);
and UO_2637 (O_2637,N_29743,N_29769);
xnor UO_2638 (O_2638,N_29569,N_29679);
nand UO_2639 (O_2639,N_29643,N_29811);
xnor UO_2640 (O_2640,N_29973,N_29612);
or UO_2641 (O_2641,N_29931,N_29841);
and UO_2642 (O_2642,N_29819,N_29799);
nand UO_2643 (O_2643,N_29875,N_29585);
nor UO_2644 (O_2644,N_29556,N_29798);
or UO_2645 (O_2645,N_29836,N_29980);
nand UO_2646 (O_2646,N_29906,N_29871);
nand UO_2647 (O_2647,N_29849,N_29630);
or UO_2648 (O_2648,N_29926,N_29775);
xor UO_2649 (O_2649,N_29771,N_29653);
xor UO_2650 (O_2650,N_29983,N_29560);
nor UO_2651 (O_2651,N_29910,N_29527);
xor UO_2652 (O_2652,N_29752,N_29781);
nand UO_2653 (O_2653,N_29952,N_29781);
and UO_2654 (O_2654,N_29575,N_29542);
or UO_2655 (O_2655,N_29878,N_29585);
nand UO_2656 (O_2656,N_29579,N_29938);
or UO_2657 (O_2657,N_29869,N_29773);
nor UO_2658 (O_2658,N_29556,N_29628);
xnor UO_2659 (O_2659,N_29706,N_29927);
nand UO_2660 (O_2660,N_29525,N_29931);
nand UO_2661 (O_2661,N_29673,N_29665);
xnor UO_2662 (O_2662,N_29952,N_29558);
and UO_2663 (O_2663,N_29803,N_29758);
and UO_2664 (O_2664,N_29899,N_29789);
nand UO_2665 (O_2665,N_29619,N_29843);
and UO_2666 (O_2666,N_29834,N_29757);
nand UO_2667 (O_2667,N_29776,N_29510);
and UO_2668 (O_2668,N_29799,N_29724);
nor UO_2669 (O_2669,N_29952,N_29715);
or UO_2670 (O_2670,N_29886,N_29934);
xnor UO_2671 (O_2671,N_29666,N_29667);
nor UO_2672 (O_2672,N_29607,N_29611);
and UO_2673 (O_2673,N_29859,N_29547);
xor UO_2674 (O_2674,N_29711,N_29984);
or UO_2675 (O_2675,N_29794,N_29682);
nor UO_2676 (O_2676,N_29904,N_29544);
or UO_2677 (O_2677,N_29544,N_29870);
and UO_2678 (O_2678,N_29662,N_29830);
or UO_2679 (O_2679,N_29864,N_29571);
nor UO_2680 (O_2680,N_29842,N_29921);
xnor UO_2681 (O_2681,N_29853,N_29885);
nor UO_2682 (O_2682,N_29769,N_29604);
xor UO_2683 (O_2683,N_29914,N_29657);
xnor UO_2684 (O_2684,N_29779,N_29951);
and UO_2685 (O_2685,N_29856,N_29756);
or UO_2686 (O_2686,N_29715,N_29594);
xor UO_2687 (O_2687,N_29561,N_29668);
nor UO_2688 (O_2688,N_29643,N_29805);
nor UO_2689 (O_2689,N_29987,N_29548);
or UO_2690 (O_2690,N_29506,N_29601);
and UO_2691 (O_2691,N_29719,N_29729);
and UO_2692 (O_2692,N_29704,N_29913);
or UO_2693 (O_2693,N_29579,N_29545);
nor UO_2694 (O_2694,N_29758,N_29988);
nor UO_2695 (O_2695,N_29838,N_29803);
nand UO_2696 (O_2696,N_29898,N_29604);
xor UO_2697 (O_2697,N_29560,N_29642);
xor UO_2698 (O_2698,N_29760,N_29649);
and UO_2699 (O_2699,N_29611,N_29992);
or UO_2700 (O_2700,N_29543,N_29975);
nor UO_2701 (O_2701,N_29986,N_29641);
nand UO_2702 (O_2702,N_29500,N_29845);
or UO_2703 (O_2703,N_29698,N_29762);
and UO_2704 (O_2704,N_29969,N_29970);
or UO_2705 (O_2705,N_29891,N_29648);
or UO_2706 (O_2706,N_29620,N_29674);
xor UO_2707 (O_2707,N_29959,N_29941);
nor UO_2708 (O_2708,N_29533,N_29736);
and UO_2709 (O_2709,N_29873,N_29914);
nand UO_2710 (O_2710,N_29516,N_29604);
nand UO_2711 (O_2711,N_29682,N_29792);
or UO_2712 (O_2712,N_29841,N_29704);
nand UO_2713 (O_2713,N_29580,N_29639);
nor UO_2714 (O_2714,N_29896,N_29632);
nor UO_2715 (O_2715,N_29582,N_29554);
or UO_2716 (O_2716,N_29760,N_29846);
and UO_2717 (O_2717,N_29970,N_29946);
and UO_2718 (O_2718,N_29772,N_29507);
or UO_2719 (O_2719,N_29681,N_29973);
nand UO_2720 (O_2720,N_29828,N_29798);
or UO_2721 (O_2721,N_29638,N_29974);
and UO_2722 (O_2722,N_29936,N_29520);
nor UO_2723 (O_2723,N_29882,N_29571);
xnor UO_2724 (O_2724,N_29980,N_29851);
xor UO_2725 (O_2725,N_29668,N_29548);
xnor UO_2726 (O_2726,N_29967,N_29955);
nand UO_2727 (O_2727,N_29798,N_29991);
nor UO_2728 (O_2728,N_29518,N_29586);
or UO_2729 (O_2729,N_29515,N_29599);
or UO_2730 (O_2730,N_29625,N_29672);
nand UO_2731 (O_2731,N_29989,N_29848);
nor UO_2732 (O_2732,N_29668,N_29962);
or UO_2733 (O_2733,N_29946,N_29632);
xnor UO_2734 (O_2734,N_29984,N_29733);
or UO_2735 (O_2735,N_29980,N_29812);
and UO_2736 (O_2736,N_29504,N_29598);
xor UO_2737 (O_2737,N_29901,N_29858);
or UO_2738 (O_2738,N_29702,N_29886);
and UO_2739 (O_2739,N_29873,N_29630);
xnor UO_2740 (O_2740,N_29592,N_29678);
or UO_2741 (O_2741,N_29997,N_29695);
or UO_2742 (O_2742,N_29872,N_29904);
or UO_2743 (O_2743,N_29971,N_29661);
nand UO_2744 (O_2744,N_29892,N_29629);
nand UO_2745 (O_2745,N_29705,N_29870);
or UO_2746 (O_2746,N_29678,N_29881);
or UO_2747 (O_2747,N_29889,N_29655);
nand UO_2748 (O_2748,N_29723,N_29657);
and UO_2749 (O_2749,N_29883,N_29940);
nand UO_2750 (O_2750,N_29952,N_29945);
and UO_2751 (O_2751,N_29810,N_29962);
nor UO_2752 (O_2752,N_29533,N_29820);
nor UO_2753 (O_2753,N_29700,N_29941);
nand UO_2754 (O_2754,N_29910,N_29665);
nand UO_2755 (O_2755,N_29563,N_29535);
nand UO_2756 (O_2756,N_29852,N_29949);
or UO_2757 (O_2757,N_29950,N_29953);
and UO_2758 (O_2758,N_29684,N_29554);
or UO_2759 (O_2759,N_29632,N_29887);
nor UO_2760 (O_2760,N_29907,N_29963);
or UO_2761 (O_2761,N_29674,N_29646);
nand UO_2762 (O_2762,N_29593,N_29526);
nand UO_2763 (O_2763,N_29869,N_29721);
and UO_2764 (O_2764,N_29540,N_29531);
and UO_2765 (O_2765,N_29841,N_29734);
nand UO_2766 (O_2766,N_29994,N_29530);
xor UO_2767 (O_2767,N_29706,N_29732);
nand UO_2768 (O_2768,N_29881,N_29514);
nor UO_2769 (O_2769,N_29599,N_29623);
nor UO_2770 (O_2770,N_29997,N_29794);
nand UO_2771 (O_2771,N_29950,N_29604);
or UO_2772 (O_2772,N_29760,N_29983);
or UO_2773 (O_2773,N_29739,N_29805);
nand UO_2774 (O_2774,N_29508,N_29939);
and UO_2775 (O_2775,N_29667,N_29902);
and UO_2776 (O_2776,N_29775,N_29792);
or UO_2777 (O_2777,N_29588,N_29704);
nor UO_2778 (O_2778,N_29610,N_29958);
nand UO_2779 (O_2779,N_29905,N_29984);
nor UO_2780 (O_2780,N_29860,N_29557);
and UO_2781 (O_2781,N_29785,N_29576);
or UO_2782 (O_2782,N_29897,N_29656);
nand UO_2783 (O_2783,N_29946,N_29797);
xor UO_2784 (O_2784,N_29985,N_29565);
or UO_2785 (O_2785,N_29903,N_29593);
and UO_2786 (O_2786,N_29805,N_29771);
or UO_2787 (O_2787,N_29832,N_29655);
nand UO_2788 (O_2788,N_29742,N_29646);
or UO_2789 (O_2789,N_29680,N_29921);
and UO_2790 (O_2790,N_29501,N_29835);
and UO_2791 (O_2791,N_29622,N_29889);
xor UO_2792 (O_2792,N_29780,N_29978);
nand UO_2793 (O_2793,N_29714,N_29613);
xor UO_2794 (O_2794,N_29756,N_29693);
nor UO_2795 (O_2795,N_29691,N_29902);
or UO_2796 (O_2796,N_29556,N_29717);
nor UO_2797 (O_2797,N_29935,N_29774);
and UO_2798 (O_2798,N_29986,N_29793);
or UO_2799 (O_2799,N_29772,N_29731);
xor UO_2800 (O_2800,N_29711,N_29988);
xor UO_2801 (O_2801,N_29624,N_29916);
xor UO_2802 (O_2802,N_29629,N_29643);
or UO_2803 (O_2803,N_29958,N_29961);
nor UO_2804 (O_2804,N_29671,N_29965);
nor UO_2805 (O_2805,N_29733,N_29591);
nand UO_2806 (O_2806,N_29958,N_29561);
nor UO_2807 (O_2807,N_29686,N_29771);
nand UO_2808 (O_2808,N_29738,N_29762);
or UO_2809 (O_2809,N_29662,N_29536);
or UO_2810 (O_2810,N_29629,N_29935);
and UO_2811 (O_2811,N_29936,N_29592);
or UO_2812 (O_2812,N_29695,N_29651);
xnor UO_2813 (O_2813,N_29923,N_29719);
or UO_2814 (O_2814,N_29837,N_29922);
and UO_2815 (O_2815,N_29585,N_29746);
nand UO_2816 (O_2816,N_29941,N_29609);
nor UO_2817 (O_2817,N_29505,N_29566);
or UO_2818 (O_2818,N_29585,N_29943);
or UO_2819 (O_2819,N_29976,N_29669);
and UO_2820 (O_2820,N_29755,N_29939);
or UO_2821 (O_2821,N_29914,N_29529);
xor UO_2822 (O_2822,N_29532,N_29939);
xor UO_2823 (O_2823,N_29590,N_29564);
or UO_2824 (O_2824,N_29828,N_29522);
xor UO_2825 (O_2825,N_29895,N_29520);
xnor UO_2826 (O_2826,N_29905,N_29539);
xor UO_2827 (O_2827,N_29591,N_29510);
or UO_2828 (O_2828,N_29883,N_29686);
and UO_2829 (O_2829,N_29710,N_29715);
and UO_2830 (O_2830,N_29682,N_29795);
xnor UO_2831 (O_2831,N_29607,N_29871);
nor UO_2832 (O_2832,N_29816,N_29631);
or UO_2833 (O_2833,N_29753,N_29500);
and UO_2834 (O_2834,N_29645,N_29976);
and UO_2835 (O_2835,N_29672,N_29762);
and UO_2836 (O_2836,N_29581,N_29967);
or UO_2837 (O_2837,N_29825,N_29579);
nand UO_2838 (O_2838,N_29595,N_29802);
nand UO_2839 (O_2839,N_29578,N_29885);
nand UO_2840 (O_2840,N_29873,N_29529);
nand UO_2841 (O_2841,N_29681,N_29643);
nor UO_2842 (O_2842,N_29871,N_29738);
and UO_2843 (O_2843,N_29861,N_29701);
nand UO_2844 (O_2844,N_29745,N_29889);
and UO_2845 (O_2845,N_29635,N_29684);
xor UO_2846 (O_2846,N_29951,N_29554);
and UO_2847 (O_2847,N_29681,N_29617);
nand UO_2848 (O_2848,N_29926,N_29646);
nand UO_2849 (O_2849,N_29690,N_29699);
nand UO_2850 (O_2850,N_29769,N_29631);
nand UO_2851 (O_2851,N_29556,N_29958);
nor UO_2852 (O_2852,N_29867,N_29870);
or UO_2853 (O_2853,N_29817,N_29927);
or UO_2854 (O_2854,N_29632,N_29620);
nor UO_2855 (O_2855,N_29603,N_29813);
and UO_2856 (O_2856,N_29920,N_29764);
nor UO_2857 (O_2857,N_29593,N_29745);
xor UO_2858 (O_2858,N_29976,N_29840);
or UO_2859 (O_2859,N_29887,N_29948);
and UO_2860 (O_2860,N_29612,N_29800);
and UO_2861 (O_2861,N_29569,N_29604);
xor UO_2862 (O_2862,N_29826,N_29993);
nand UO_2863 (O_2863,N_29715,N_29510);
or UO_2864 (O_2864,N_29783,N_29759);
or UO_2865 (O_2865,N_29982,N_29748);
nand UO_2866 (O_2866,N_29561,N_29579);
or UO_2867 (O_2867,N_29511,N_29813);
and UO_2868 (O_2868,N_29540,N_29772);
xor UO_2869 (O_2869,N_29556,N_29639);
nor UO_2870 (O_2870,N_29684,N_29961);
xnor UO_2871 (O_2871,N_29698,N_29962);
xor UO_2872 (O_2872,N_29528,N_29982);
xor UO_2873 (O_2873,N_29641,N_29584);
or UO_2874 (O_2874,N_29620,N_29541);
xor UO_2875 (O_2875,N_29990,N_29945);
nor UO_2876 (O_2876,N_29504,N_29568);
or UO_2877 (O_2877,N_29853,N_29861);
nor UO_2878 (O_2878,N_29733,N_29795);
and UO_2879 (O_2879,N_29673,N_29649);
xor UO_2880 (O_2880,N_29826,N_29642);
or UO_2881 (O_2881,N_29816,N_29944);
and UO_2882 (O_2882,N_29769,N_29751);
nor UO_2883 (O_2883,N_29631,N_29668);
nand UO_2884 (O_2884,N_29550,N_29974);
and UO_2885 (O_2885,N_29830,N_29688);
xor UO_2886 (O_2886,N_29580,N_29560);
nand UO_2887 (O_2887,N_29650,N_29516);
nand UO_2888 (O_2888,N_29684,N_29758);
and UO_2889 (O_2889,N_29710,N_29916);
or UO_2890 (O_2890,N_29964,N_29635);
nand UO_2891 (O_2891,N_29928,N_29563);
nor UO_2892 (O_2892,N_29536,N_29732);
xor UO_2893 (O_2893,N_29623,N_29659);
xnor UO_2894 (O_2894,N_29543,N_29773);
nor UO_2895 (O_2895,N_29660,N_29892);
and UO_2896 (O_2896,N_29517,N_29680);
or UO_2897 (O_2897,N_29616,N_29513);
nor UO_2898 (O_2898,N_29984,N_29554);
xnor UO_2899 (O_2899,N_29658,N_29790);
and UO_2900 (O_2900,N_29699,N_29707);
and UO_2901 (O_2901,N_29961,N_29713);
nand UO_2902 (O_2902,N_29776,N_29609);
and UO_2903 (O_2903,N_29549,N_29738);
and UO_2904 (O_2904,N_29830,N_29772);
nand UO_2905 (O_2905,N_29954,N_29997);
and UO_2906 (O_2906,N_29915,N_29873);
nand UO_2907 (O_2907,N_29787,N_29741);
and UO_2908 (O_2908,N_29611,N_29518);
nor UO_2909 (O_2909,N_29889,N_29554);
and UO_2910 (O_2910,N_29717,N_29694);
xnor UO_2911 (O_2911,N_29708,N_29900);
and UO_2912 (O_2912,N_29851,N_29544);
nand UO_2913 (O_2913,N_29697,N_29723);
nand UO_2914 (O_2914,N_29943,N_29912);
nor UO_2915 (O_2915,N_29754,N_29956);
or UO_2916 (O_2916,N_29554,N_29773);
xor UO_2917 (O_2917,N_29833,N_29795);
nor UO_2918 (O_2918,N_29576,N_29933);
or UO_2919 (O_2919,N_29522,N_29971);
or UO_2920 (O_2920,N_29579,N_29502);
xnor UO_2921 (O_2921,N_29680,N_29784);
and UO_2922 (O_2922,N_29921,N_29668);
nand UO_2923 (O_2923,N_29966,N_29699);
nand UO_2924 (O_2924,N_29771,N_29718);
or UO_2925 (O_2925,N_29690,N_29681);
and UO_2926 (O_2926,N_29873,N_29884);
or UO_2927 (O_2927,N_29845,N_29765);
nor UO_2928 (O_2928,N_29802,N_29690);
or UO_2929 (O_2929,N_29750,N_29628);
nand UO_2930 (O_2930,N_29647,N_29875);
xor UO_2931 (O_2931,N_29942,N_29590);
nor UO_2932 (O_2932,N_29852,N_29978);
xor UO_2933 (O_2933,N_29907,N_29939);
and UO_2934 (O_2934,N_29597,N_29749);
or UO_2935 (O_2935,N_29855,N_29977);
nand UO_2936 (O_2936,N_29946,N_29773);
or UO_2937 (O_2937,N_29595,N_29735);
nand UO_2938 (O_2938,N_29754,N_29560);
or UO_2939 (O_2939,N_29590,N_29957);
nor UO_2940 (O_2940,N_29984,N_29657);
nor UO_2941 (O_2941,N_29879,N_29589);
or UO_2942 (O_2942,N_29615,N_29922);
xor UO_2943 (O_2943,N_29948,N_29560);
and UO_2944 (O_2944,N_29943,N_29842);
and UO_2945 (O_2945,N_29965,N_29781);
nor UO_2946 (O_2946,N_29771,N_29536);
or UO_2947 (O_2947,N_29677,N_29963);
and UO_2948 (O_2948,N_29757,N_29939);
nand UO_2949 (O_2949,N_29878,N_29618);
and UO_2950 (O_2950,N_29551,N_29837);
xnor UO_2951 (O_2951,N_29661,N_29840);
and UO_2952 (O_2952,N_29808,N_29513);
nand UO_2953 (O_2953,N_29873,N_29843);
and UO_2954 (O_2954,N_29733,N_29738);
or UO_2955 (O_2955,N_29913,N_29510);
or UO_2956 (O_2956,N_29636,N_29892);
xor UO_2957 (O_2957,N_29592,N_29531);
and UO_2958 (O_2958,N_29647,N_29729);
xnor UO_2959 (O_2959,N_29985,N_29764);
nor UO_2960 (O_2960,N_29667,N_29512);
or UO_2961 (O_2961,N_29950,N_29794);
xnor UO_2962 (O_2962,N_29885,N_29969);
or UO_2963 (O_2963,N_29956,N_29865);
nand UO_2964 (O_2964,N_29766,N_29535);
nor UO_2965 (O_2965,N_29959,N_29956);
nor UO_2966 (O_2966,N_29726,N_29843);
and UO_2967 (O_2967,N_29966,N_29852);
or UO_2968 (O_2968,N_29742,N_29783);
nor UO_2969 (O_2969,N_29942,N_29513);
xor UO_2970 (O_2970,N_29816,N_29528);
and UO_2971 (O_2971,N_29543,N_29760);
and UO_2972 (O_2972,N_29727,N_29923);
xnor UO_2973 (O_2973,N_29873,N_29680);
nor UO_2974 (O_2974,N_29544,N_29862);
or UO_2975 (O_2975,N_29948,N_29618);
nor UO_2976 (O_2976,N_29809,N_29894);
and UO_2977 (O_2977,N_29732,N_29624);
nor UO_2978 (O_2978,N_29931,N_29895);
xnor UO_2979 (O_2979,N_29598,N_29626);
or UO_2980 (O_2980,N_29565,N_29537);
or UO_2981 (O_2981,N_29785,N_29841);
or UO_2982 (O_2982,N_29779,N_29961);
or UO_2983 (O_2983,N_29846,N_29756);
nand UO_2984 (O_2984,N_29807,N_29886);
and UO_2985 (O_2985,N_29996,N_29638);
xnor UO_2986 (O_2986,N_29897,N_29530);
or UO_2987 (O_2987,N_29555,N_29762);
and UO_2988 (O_2988,N_29973,N_29692);
or UO_2989 (O_2989,N_29713,N_29855);
or UO_2990 (O_2990,N_29758,N_29666);
nand UO_2991 (O_2991,N_29900,N_29571);
or UO_2992 (O_2992,N_29828,N_29690);
xor UO_2993 (O_2993,N_29967,N_29883);
or UO_2994 (O_2994,N_29642,N_29709);
nand UO_2995 (O_2995,N_29714,N_29571);
xnor UO_2996 (O_2996,N_29916,N_29878);
xnor UO_2997 (O_2997,N_29978,N_29968);
or UO_2998 (O_2998,N_29710,N_29816);
nand UO_2999 (O_2999,N_29608,N_29819);
nor UO_3000 (O_3000,N_29891,N_29547);
and UO_3001 (O_3001,N_29800,N_29638);
nand UO_3002 (O_3002,N_29940,N_29611);
xor UO_3003 (O_3003,N_29656,N_29578);
or UO_3004 (O_3004,N_29886,N_29516);
nor UO_3005 (O_3005,N_29608,N_29927);
nor UO_3006 (O_3006,N_29663,N_29686);
and UO_3007 (O_3007,N_29961,N_29606);
or UO_3008 (O_3008,N_29903,N_29583);
or UO_3009 (O_3009,N_29889,N_29749);
nor UO_3010 (O_3010,N_29836,N_29670);
nor UO_3011 (O_3011,N_29590,N_29779);
nor UO_3012 (O_3012,N_29847,N_29572);
or UO_3013 (O_3013,N_29564,N_29596);
nor UO_3014 (O_3014,N_29850,N_29977);
xor UO_3015 (O_3015,N_29507,N_29991);
nor UO_3016 (O_3016,N_29995,N_29652);
and UO_3017 (O_3017,N_29979,N_29619);
or UO_3018 (O_3018,N_29772,N_29832);
or UO_3019 (O_3019,N_29582,N_29589);
or UO_3020 (O_3020,N_29616,N_29951);
nand UO_3021 (O_3021,N_29581,N_29830);
xor UO_3022 (O_3022,N_29798,N_29520);
xnor UO_3023 (O_3023,N_29772,N_29943);
nor UO_3024 (O_3024,N_29670,N_29995);
nor UO_3025 (O_3025,N_29768,N_29734);
nor UO_3026 (O_3026,N_29800,N_29834);
xnor UO_3027 (O_3027,N_29556,N_29739);
xnor UO_3028 (O_3028,N_29534,N_29587);
nand UO_3029 (O_3029,N_29892,N_29914);
nor UO_3030 (O_3030,N_29808,N_29798);
xnor UO_3031 (O_3031,N_29659,N_29605);
nand UO_3032 (O_3032,N_29525,N_29708);
nor UO_3033 (O_3033,N_29913,N_29669);
xor UO_3034 (O_3034,N_29706,N_29994);
and UO_3035 (O_3035,N_29980,N_29660);
nor UO_3036 (O_3036,N_29642,N_29521);
nand UO_3037 (O_3037,N_29867,N_29500);
and UO_3038 (O_3038,N_29678,N_29655);
nand UO_3039 (O_3039,N_29975,N_29542);
nor UO_3040 (O_3040,N_29600,N_29751);
xor UO_3041 (O_3041,N_29502,N_29574);
nor UO_3042 (O_3042,N_29806,N_29776);
xor UO_3043 (O_3043,N_29720,N_29500);
nand UO_3044 (O_3044,N_29866,N_29616);
xor UO_3045 (O_3045,N_29665,N_29817);
xnor UO_3046 (O_3046,N_29712,N_29829);
nor UO_3047 (O_3047,N_29923,N_29970);
or UO_3048 (O_3048,N_29995,N_29717);
and UO_3049 (O_3049,N_29800,N_29775);
nor UO_3050 (O_3050,N_29508,N_29683);
or UO_3051 (O_3051,N_29982,N_29694);
nor UO_3052 (O_3052,N_29721,N_29813);
nor UO_3053 (O_3053,N_29619,N_29693);
xor UO_3054 (O_3054,N_29554,N_29731);
and UO_3055 (O_3055,N_29649,N_29592);
or UO_3056 (O_3056,N_29774,N_29670);
nor UO_3057 (O_3057,N_29690,N_29776);
and UO_3058 (O_3058,N_29578,N_29696);
and UO_3059 (O_3059,N_29855,N_29961);
nor UO_3060 (O_3060,N_29829,N_29774);
and UO_3061 (O_3061,N_29721,N_29575);
nor UO_3062 (O_3062,N_29660,N_29601);
xor UO_3063 (O_3063,N_29511,N_29703);
and UO_3064 (O_3064,N_29984,N_29791);
or UO_3065 (O_3065,N_29755,N_29972);
nand UO_3066 (O_3066,N_29546,N_29620);
nor UO_3067 (O_3067,N_29783,N_29952);
xor UO_3068 (O_3068,N_29866,N_29636);
xnor UO_3069 (O_3069,N_29684,N_29609);
nand UO_3070 (O_3070,N_29520,N_29884);
nand UO_3071 (O_3071,N_29605,N_29552);
nand UO_3072 (O_3072,N_29925,N_29518);
or UO_3073 (O_3073,N_29877,N_29982);
nand UO_3074 (O_3074,N_29994,N_29749);
nor UO_3075 (O_3075,N_29617,N_29677);
and UO_3076 (O_3076,N_29946,N_29540);
nand UO_3077 (O_3077,N_29657,N_29976);
or UO_3078 (O_3078,N_29511,N_29895);
or UO_3079 (O_3079,N_29935,N_29972);
or UO_3080 (O_3080,N_29547,N_29870);
nand UO_3081 (O_3081,N_29545,N_29680);
nor UO_3082 (O_3082,N_29556,N_29924);
nor UO_3083 (O_3083,N_29846,N_29765);
and UO_3084 (O_3084,N_29983,N_29522);
nand UO_3085 (O_3085,N_29927,N_29503);
nor UO_3086 (O_3086,N_29824,N_29912);
or UO_3087 (O_3087,N_29943,N_29617);
and UO_3088 (O_3088,N_29936,N_29598);
nor UO_3089 (O_3089,N_29702,N_29501);
nor UO_3090 (O_3090,N_29823,N_29836);
nand UO_3091 (O_3091,N_29730,N_29523);
nand UO_3092 (O_3092,N_29887,N_29905);
nand UO_3093 (O_3093,N_29716,N_29633);
nand UO_3094 (O_3094,N_29723,N_29934);
nor UO_3095 (O_3095,N_29626,N_29909);
xor UO_3096 (O_3096,N_29631,N_29807);
or UO_3097 (O_3097,N_29933,N_29698);
and UO_3098 (O_3098,N_29757,N_29707);
nor UO_3099 (O_3099,N_29546,N_29989);
and UO_3100 (O_3100,N_29874,N_29698);
and UO_3101 (O_3101,N_29809,N_29931);
nand UO_3102 (O_3102,N_29506,N_29981);
nand UO_3103 (O_3103,N_29953,N_29651);
xnor UO_3104 (O_3104,N_29599,N_29975);
xnor UO_3105 (O_3105,N_29509,N_29760);
xor UO_3106 (O_3106,N_29817,N_29684);
or UO_3107 (O_3107,N_29785,N_29645);
and UO_3108 (O_3108,N_29871,N_29720);
xnor UO_3109 (O_3109,N_29585,N_29803);
and UO_3110 (O_3110,N_29949,N_29522);
xor UO_3111 (O_3111,N_29523,N_29622);
nand UO_3112 (O_3112,N_29895,N_29701);
or UO_3113 (O_3113,N_29637,N_29582);
nor UO_3114 (O_3114,N_29677,N_29716);
nor UO_3115 (O_3115,N_29936,N_29763);
nand UO_3116 (O_3116,N_29634,N_29938);
nand UO_3117 (O_3117,N_29701,N_29557);
nor UO_3118 (O_3118,N_29671,N_29732);
nor UO_3119 (O_3119,N_29784,N_29949);
nand UO_3120 (O_3120,N_29684,N_29904);
nand UO_3121 (O_3121,N_29637,N_29610);
nand UO_3122 (O_3122,N_29995,N_29710);
nor UO_3123 (O_3123,N_29608,N_29527);
nor UO_3124 (O_3124,N_29995,N_29979);
and UO_3125 (O_3125,N_29909,N_29791);
or UO_3126 (O_3126,N_29596,N_29722);
and UO_3127 (O_3127,N_29707,N_29602);
xor UO_3128 (O_3128,N_29978,N_29506);
and UO_3129 (O_3129,N_29984,N_29639);
and UO_3130 (O_3130,N_29544,N_29654);
xor UO_3131 (O_3131,N_29918,N_29545);
nand UO_3132 (O_3132,N_29718,N_29885);
nor UO_3133 (O_3133,N_29538,N_29977);
nor UO_3134 (O_3134,N_29656,N_29519);
xnor UO_3135 (O_3135,N_29952,N_29777);
and UO_3136 (O_3136,N_29504,N_29512);
nor UO_3137 (O_3137,N_29552,N_29939);
or UO_3138 (O_3138,N_29902,N_29627);
or UO_3139 (O_3139,N_29539,N_29650);
nor UO_3140 (O_3140,N_29954,N_29717);
or UO_3141 (O_3141,N_29863,N_29799);
nor UO_3142 (O_3142,N_29677,N_29862);
or UO_3143 (O_3143,N_29568,N_29901);
and UO_3144 (O_3144,N_29865,N_29575);
xnor UO_3145 (O_3145,N_29819,N_29542);
and UO_3146 (O_3146,N_29804,N_29999);
xor UO_3147 (O_3147,N_29870,N_29666);
and UO_3148 (O_3148,N_29657,N_29739);
or UO_3149 (O_3149,N_29505,N_29850);
nand UO_3150 (O_3150,N_29885,N_29828);
nor UO_3151 (O_3151,N_29589,N_29841);
or UO_3152 (O_3152,N_29859,N_29769);
or UO_3153 (O_3153,N_29818,N_29817);
nor UO_3154 (O_3154,N_29935,N_29921);
xnor UO_3155 (O_3155,N_29510,N_29698);
or UO_3156 (O_3156,N_29522,N_29655);
and UO_3157 (O_3157,N_29823,N_29640);
nor UO_3158 (O_3158,N_29838,N_29853);
nand UO_3159 (O_3159,N_29873,N_29541);
or UO_3160 (O_3160,N_29872,N_29644);
nand UO_3161 (O_3161,N_29827,N_29813);
nor UO_3162 (O_3162,N_29835,N_29837);
xor UO_3163 (O_3163,N_29504,N_29632);
and UO_3164 (O_3164,N_29979,N_29548);
and UO_3165 (O_3165,N_29747,N_29748);
nand UO_3166 (O_3166,N_29529,N_29801);
nor UO_3167 (O_3167,N_29614,N_29767);
and UO_3168 (O_3168,N_29611,N_29579);
nand UO_3169 (O_3169,N_29827,N_29924);
or UO_3170 (O_3170,N_29927,N_29858);
xnor UO_3171 (O_3171,N_29650,N_29631);
nor UO_3172 (O_3172,N_29795,N_29501);
or UO_3173 (O_3173,N_29895,N_29677);
and UO_3174 (O_3174,N_29660,N_29702);
nor UO_3175 (O_3175,N_29920,N_29889);
nand UO_3176 (O_3176,N_29914,N_29579);
xnor UO_3177 (O_3177,N_29872,N_29760);
or UO_3178 (O_3178,N_29900,N_29500);
and UO_3179 (O_3179,N_29795,N_29515);
nand UO_3180 (O_3180,N_29665,N_29504);
and UO_3181 (O_3181,N_29587,N_29648);
xnor UO_3182 (O_3182,N_29795,N_29536);
and UO_3183 (O_3183,N_29927,N_29803);
and UO_3184 (O_3184,N_29612,N_29910);
nor UO_3185 (O_3185,N_29567,N_29753);
nand UO_3186 (O_3186,N_29650,N_29555);
and UO_3187 (O_3187,N_29579,N_29538);
nor UO_3188 (O_3188,N_29983,N_29892);
or UO_3189 (O_3189,N_29583,N_29832);
or UO_3190 (O_3190,N_29673,N_29834);
nand UO_3191 (O_3191,N_29610,N_29869);
xnor UO_3192 (O_3192,N_29994,N_29948);
or UO_3193 (O_3193,N_29692,N_29971);
and UO_3194 (O_3194,N_29713,N_29836);
and UO_3195 (O_3195,N_29565,N_29594);
xor UO_3196 (O_3196,N_29509,N_29817);
nand UO_3197 (O_3197,N_29834,N_29934);
and UO_3198 (O_3198,N_29716,N_29993);
nor UO_3199 (O_3199,N_29642,N_29537);
and UO_3200 (O_3200,N_29787,N_29568);
nand UO_3201 (O_3201,N_29893,N_29982);
nand UO_3202 (O_3202,N_29660,N_29691);
xnor UO_3203 (O_3203,N_29903,N_29840);
xor UO_3204 (O_3204,N_29627,N_29785);
xnor UO_3205 (O_3205,N_29986,N_29666);
or UO_3206 (O_3206,N_29959,N_29752);
xnor UO_3207 (O_3207,N_29907,N_29897);
or UO_3208 (O_3208,N_29779,N_29529);
xor UO_3209 (O_3209,N_29570,N_29660);
xnor UO_3210 (O_3210,N_29547,N_29982);
and UO_3211 (O_3211,N_29609,N_29822);
nand UO_3212 (O_3212,N_29888,N_29971);
xor UO_3213 (O_3213,N_29617,N_29914);
or UO_3214 (O_3214,N_29950,N_29570);
xor UO_3215 (O_3215,N_29504,N_29897);
nor UO_3216 (O_3216,N_29707,N_29884);
and UO_3217 (O_3217,N_29685,N_29714);
or UO_3218 (O_3218,N_29765,N_29592);
and UO_3219 (O_3219,N_29866,N_29943);
xnor UO_3220 (O_3220,N_29598,N_29888);
and UO_3221 (O_3221,N_29834,N_29927);
nand UO_3222 (O_3222,N_29666,N_29719);
or UO_3223 (O_3223,N_29853,N_29546);
nor UO_3224 (O_3224,N_29814,N_29553);
nor UO_3225 (O_3225,N_29509,N_29545);
or UO_3226 (O_3226,N_29515,N_29567);
nor UO_3227 (O_3227,N_29752,N_29681);
and UO_3228 (O_3228,N_29901,N_29864);
nand UO_3229 (O_3229,N_29819,N_29947);
and UO_3230 (O_3230,N_29804,N_29843);
and UO_3231 (O_3231,N_29866,N_29863);
xnor UO_3232 (O_3232,N_29519,N_29859);
nand UO_3233 (O_3233,N_29690,N_29901);
nor UO_3234 (O_3234,N_29757,N_29911);
nand UO_3235 (O_3235,N_29526,N_29993);
or UO_3236 (O_3236,N_29504,N_29526);
nand UO_3237 (O_3237,N_29793,N_29733);
xor UO_3238 (O_3238,N_29982,N_29811);
or UO_3239 (O_3239,N_29710,N_29833);
or UO_3240 (O_3240,N_29912,N_29842);
xnor UO_3241 (O_3241,N_29683,N_29659);
xor UO_3242 (O_3242,N_29557,N_29982);
nor UO_3243 (O_3243,N_29888,N_29784);
nor UO_3244 (O_3244,N_29773,N_29757);
xnor UO_3245 (O_3245,N_29525,N_29675);
xor UO_3246 (O_3246,N_29631,N_29975);
or UO_3247 (O_3247,N_29580,N_29916);
xnor UO_3248 (O_3248,N_29964,N_29845);
nand UO_3249 (O_3249,N_29941,N_29754);
and UO_3250 (O_3250,N_29931,N_29848);
xor UO_3251 (O_3251,N_29862,N_29830);
and UO_3252 (O_3252,N_29583,N_29871);
and UO_3253 (O_3253,N_29518,N_29608);
and UO_3254 (O_3254,N_29898,N_29598);
or UO_3255 (O_3255,N_29910,N_29890);
nor UO_3256 (O_3256,N_29985,N_29674);
nand UO_3257 (O_3257,N_29691,N_29610);
nand UO_3258 (O_3258,N_29650,N_29592);
nor UO_3259 (O_3259,N_29594,N_29787);
or UO_3260 (O_3260,N_29855,N_29508);
nand UO_3261 (O_3261,N_29991,N_29784);
nor UO_3262 (O_3262,N_29918,N_29927);
and UO_3263 (O_3263,N_29631,N_29995);
or UO_3264 (O_3264,N_29876,N_29994);
nor UO_3265 (O_3265,N_29671,N_29506);
nand UO_3266 (O_3266,N_29818,N_29674);
and UO_3267 (O_3267,N_29871,N_29585);
xnor UO_3268 (O_3268,N_29905,N_29882);
xnor UO_3269 (O_3269,N_29893,N_29630);
or UO_3270 (O_3270,N_29683,N_29953);
xor UO_3271 (O_3271,N_29656,N_29725);
xor UO_3272 (O_3272,N_29745,N_29952);
xnor UO_3273 (O_3273,N_29753,N_29889);
xor UO_3274 (O_3274,N_29684,N_29986);
or UO_3275 (O_3275,N_29842,N_29644);
and UO_3276 (O_3276,N_29568,N_29842);
xnor UO_3277 (O_3277,N_29660,N_29917);
and UO_3278 (O_3278,N_29900,N_29618);
xnor UO_3279 (O_3279,N_29934,N_29649);
and UO_3280 (O_3280,N_29685,N_29924);
xor UO_3281 (O_3281,N_29997,N_29785);
and UO_3282 (O_3282,N_29876,N_29997);
xnor UO_3283 (O_3283,N_29617,N_29994);
nor UO_3284 (O_3284,N_29604,N_29973);
and UO_3285 (O_3285,N_29872,N_29868);
xor UO_3286 (O_3286,N_29503,N_29918);
xnor UO_3287 (O_3287,N_29805,N_29850);
and UO_3288 (O_3288,N_29713,N_29703);
or UO_3289 (O_3289,N_29680,N_29536);
or UO_3290 (O_3290,N_29796,N_29787);
and UO_3291 (O_3291,N_29859,N_29901);
xor UO_3292 (O_3292,N_29754,N_29710);
nor UO_3293 (O_3293,N_29642,N_29527);
or UO_3294 (O_3294,N_29910,N_29556);
and UO_3295 (O_3295,N_29676,N_29941);
or UO_3296 (O_3296,N_29946,N_29629);
xor UO_3297 (O_3297,N_29938,N_29507);
nand UO_3298 (O_3298,N_29880,N_29670);
xnor UO_3299 (O_3299,N_29619,N_29594);
nand UO_3300 (O_3300,N_29699,N_29533);
or UO_3301 (O_3301,N_29657,N_29606);
xnor UO_3302 (O_3302,N_29994,N_29624);
xnor UO_3303 (O_3303,N_29996,N_29724);
and UO_3304 (O_3304,N_29849,N_29620);
xnor UO_3305 (O_3305,N_29872,N_29735);
nor UO_3306 (O_3306,N_29821,N_29999);
xnor UO_3307 (O_3307,N_29519,N_29999);
or UO_3308 (O_3308,N_29924,N_29551);
or UO_3309 (O_3309,N_29749,N_29993);
nor UO_3310 (O_3310,N_29756,N_29678);
or UO_3311 (O_3311,N_29789,N_29612);
or UO_3312 (O_3312,N_29507,N_29545);
nor UO_3313 (O_3313,N_29918,N_29999);
nand UO_3314 (O_3314,N_29668,N_29837);
nand UO_3315 (O_3315,N_29811,N_29684);
xnor UO_3316 (O_3316,N_29550,N_29824);
xnor UO_3317 (O_3317,N_29645,N_29949);
nand UO_3318 (O_3318,N_29870,N_29928);
xnor UO_3319 (O_3319,N_29969,N_29746);
and UO_3320 (O_3320,N_29852,N_29592);
or UO_3321 (O_3321,N_29585,N_29865);
nor UO_3322 (O_3322,N_29755,N_29639);
and UO_3323 (O_3323,N_29768,N_29651);
and UO_3324 (O_3324,N_29784,N_29939);
xnor UO_3325 (O_3325,N_29908,N_29518);
and UO_3326 (O_3326,N_29841,N_29579);
nand UO_3327 (O_3327,N_29792,N_29923);
nand UO_3328 (O_3328,N_29592,N_29509);
or UO_3329 (O_3329,N_29589,N_29701);
and UO_3330 (O_3330,N_29867,N_29542);
nand UO_3331 (O_3331,N_29725,N_29732);
nor UO_3332 (O_3332,N_29776,N_29630);
nand UO_3333 (O_3333,N_29512,N_29809);
xnor UO_3334 (O_3334,N_29857,N_29516);
nor UO_3335 (O_3335,N_29684,N_29725);
and UO_3336 (O_3336,N_29650,N_29939);
xnor UO_3337 (O_3337,N_29925,N_29987);
or UO_3338 (O_3338,N_29513,N_29943);
and UO_3339 (O_3339,N_29623,N_29631);
xor UO_3340 (O_3340,N_29799,N_29598);
nor UO_3341 (O_3341,N_29969,N_29731);
and UO_3342 (O_3342,N_29962,N_29827);
or UO_3343 (O_3343,N_29927,N_29871);
or UO_3344 (O_3344,N_29878,N_29601);
and UO_3345 (O_3345,N_29623,N_29593);
xnor UO_3346 (O_3346,N_29617,N_29900);
xnor UO_3347 (O_3347,N_29545,N_29552);
and UO_3348 (O_3348,N_29782,N_29531);
and UO_3349 (O_3349,N_29505,N_29637);
nand UO_3350 (O_3350,N_29924,N_29844);
xor UO_3351 (O_3351,N_29838,N_29750);
xor UO_3352 (O_3352,N_29882,N_29709);
nor UO_3353 (O_3353,N_29762,N_29880);
nor UO_3354 (O_3354,N_29881,N_29801);
xor UO_3355 (O_3355,N_29979,N_29641);
nor UO_3356 (O_3356,N_29685,N_29929);
nor UO_3357 (O_3357,N_29742,N_29740);
nor UO_3358 (O_3358,N_29656,N_29724);
xor UO_3359 (O_3359,N_29746,N_29787);
or UO_3360 (O_3360,N_29985,N_29696);
nand UO_3361 (O_3361,N_29685,N_29980);
or UO_3362 (O_3362,N_29796,N_29630);
nand UO_3363 (O_3363,N_29908,N_29707);
xor UO_3364 (O_3364,N_29841,N_29703);
nor UO_3365 (O_3365,N_29667,N_29819);
or UO_3366 (O_3366,N_29671,N_29647);
nor UO_3367 (O_3367,N_29718,N_29968);
or UO_3368 (O_3368,N_29559,N_29858);
or UO_3369 (O_3369,N_29640,N_29549);
and UO_3370 (O_3370,N_29917,N_29624);
and UO_3371 (O_3371,N_29584,N_29748);
and UO_3372 (O_3372,N_29928,N_29719);
or UO_3373 (O_3373,N_29624,N_29609);
or UO_3374 (O_3374,N_29613,N_29648);
nor UO_3375 (O_3375,N_29932,N_29528);
nand UO_3376 (O_3376,N_29604,N_29625);
nor UO_3377 (O_3377,N_29866,N_29836);
xor UO_3378 (O_3378,N_29948,N_29701);
nand UO_3379 (O_3379,N_29675,N_29732);
nand UO_3380 (O_3380,N_29721,N_29786);
nor UO_3381 (O_3381,N_29918,N_29863);
nand UO_3382 (O_3382,N_29725,N_29825);
nand UO_3383 (O_3383,N_29896,N_29505);
and UO_3384 (O_3384,N_29866,N_29887);
xor UO_3385 (O_3385,N_29955,N_29752);
xnor UO_3386 (O_3386,N_29832,N_29760);
xnor UO_3387 (O_3387,N_29535,N_29648);
and UO_3388 (O_3388,N_29647,N_29718);
or UO_3389 (O_3389,N_29726,N_29890);
xnor UO_3390 (O_3390,N_29575,N_29555);
xor UO_3391 (O_3391,N_29694,N_29912);
xor UO_3392 (O_3392,N_29898,N_29746);
or UO_3393 (O_3393,N_29513,N_29552);
or UO_3394 (O_3394,N_29846,N_29592);
xor UO_3395 (O_3395,N_29997,N_29825);
nand UO_3396 (O_3396,N_29784,N_29556);
nor UO_3397 (O_3397,N_29619,N_29584);
xor UO_3398 (O_3398,N_29758,N_29544);
nand UO_3399 (O_3399,N_29667,N_29507);
and UO_3400 (O_3400,N_29967,N_29749);
xor UO_3401 (O_3401,N_29930,N_29861);
or UO_3402 (O_3402,N_29997,N_29641);
or UO_3403 (O_3403,N_29939,N_29985);
nor UO_3404 (O_3404,N_29625,N_29929);
xnor UO_3405 (O_3405,N_29612,N_29719);
or UO_3406 (O_3406,N_29753,N_29537);
xnor UO_3407 (O_3407,N_29585,N_29986);
or UO_3408 (O_3408,N_29693,N_29834);
or UO_3409 (O_3409,N_29542,N_29640);
or UO_3410 (O_3410,N_29523,N_29677);
nand UO_3411 (O_3411,N_29681,N_29518);
or UO_3412 (O_3412,N_29917,N_29769);
xor UO_3413 (O_3413,N_29780,N_29998);
nor UO_3414 (O_3414,N_29663,N_29853);
or UO_3415 (O_3415,N_29697,N_29731);
nand UO_3416 (O_3416,N_29832,N_29990);
nand UO_3417 (O_3417,N_29901,N_29795);
nor UO_3418 (O_3418,N_29865,N_29636);
nand UO_3419 (O_3419,N_29871,N_29977);
nor UO_3420 (O_3420,N_29762,N_29818);
and UO_3421 (O_3421,N_29819,N_29887);
nand UO_3422 (O_3422,N_29563,N_29632);
and UO_3423 (O_3423,N_29990,N_29708);
nand UO_3424 (O_3424,N_29797,N_29754);
or UO_3425 (O_3425,N_29524,N_29715);
xnor UO_3426 (O_3426,N_29873,N_29635);
or UO_3427 (O_3427,N_29933,N_29795);
xor UO_3428 (O_3428,N_29812,N_29665);
and UO_3429 (O_3429,N_29784,N_29876);
nor UO_3430 (O_3430,N_29776,N_29658);
or UO_3431 (O_3431,N_29561,N_29986);
nor UO_3432 (O_3432,N_29959,N_29685);
and UO_3433 (O_3433,N_29707,N_29864);
and UO_3434 (O_3434,N_29723,N_29694);
or UO_3435 (O_3435,N_29841,N_29634);
nor UO_3436 (O_3436,N_29743,N_29610);
xnor UO_3437 (O_3437,N_29691,N_29838);
or UO_3438 (O_3438,N_29821,N_29902);
xnor UO_3439 (O_3439,N_29622,N_29972);
nand UO_3440 (O_3440,N_29705,N_29554);
or UO_3441 (O_3441,N_29670,N_29740);
or UO_3442 (O_3442,N_29991,N_29623);
and UO_3443 (O_3443,N_29729,N_29777);
or UO_3444 (O_3444,N_29600,N_29667);
and UO_3445 (O_3445,N_29998,N_29763);
xnor UO_3446 (O_3446,N_29973,N_29912);
nor UO_3447 (O_3447,N_29555,N_29674);
or UO_3448 (O_3448,N_29881,N_29637);
nand UO_3449 (O_3449,N_29758,N_29863);
and UO_3450 (O_3450,N_29766,N_29980);
xnor UO_3451 (O_3451,N_29652,N_29883);
or UO_3452 (O_3452,N_29785,N_29906);
and UO_3453 (O_3453,N_29838,N_29621);
or UO_3454 (O_3454,N_29776,N_29745);
nor UO_3455 (O_3455,N_29917,N_29721);
nor UO_3456 (O_3456,N_29568,N_29734);
xor UO_3457 (O_3457,N_29858,N_29588);
or UO_3458 (O_3458,N_29751,N_29785);
nor UO_3459 (O_3459,N_29559,N_29667);
nor UO_3460 (O_3460,N_29782,N_29601);
or UO_3461 (O_3461,N_29728,N_29822);
and UO_3462 (O_3462,N_29986,N_29780);
and UO_3463 (O_3463,N_29540,N_29888);
and UO_3464 (O_3464,N_29873,N_29787);
xnor UO_3465 (O_3465,N_29699,N_29815);
or UO_3466 (O_3466,N_29626,N_29718);
nand UO_3467 (O_3467,N_29701,N_29585);
nand UO_3468 (O_3468,N_29627,N_29900);
nand UO_3469 (O_3469,N_29941,N_29565);
and UO_3470 (O_3470,N_29987,N_29793);
and UO_3471 (O_3471,N_29747,N_29833);
xnor UO_3472 (O_3472,N_29915,N_29868);
or UO_3473 (O_3473,N_29605,N_29919);
nor UO_3474 (O_3474,N_29930,N_29872);
and UO_3475 (O_3475,N_29650,N_29611);
or UO_3476 (O_3476,N_29977,N_29615);
xnor UO_3477 (O_3477,N_29970,N_29558);
xor UO_3478 (O_3478,N_29992,N_29664);
or UO_3479 (O_3479,N_29932,N_29897);
nand UO_3480 (O_3480,N_29726,N_29650);
and UO_3481 (O_3481,N_29955,N_29515);
nor UO_3482 (O_3482,N_29790,N_29774);
nand UO_3483 (O_3483,N_29593,N_29947);
nand UO_3484 (O_3484,N_29529,N_29638);
nand UO_3485 (O_3485,N_29609,N_29993);
xor UO_3486 (O_3486,N_29700,N_29579);
and UO_3487 (O_3487,N_29518,N_29858);
nand UO_3488 (O_3488,N_29960,N_29821);
or UO_3489 (O_3489,N_29929,N_29852);
and UO_3490 (O_3490,N_29725,N_29701);
nand UO_3491 (O_3491,N_29893,N_29857);
xnor UO_3492 (O_3492,N_29595,N_29771);
nand UO_3493 (O_3493,N_29838,N_29815);
nand UO_3494 (O_3494,N_29825,N_29985);
xnor UO_3495 (O_3495,N_29577,N_29512);
xor UO_3496 (O_3496,N_29522,N_29651);
xor UO_3497 (O_3497,N_29671,N_29790);
or UO_3498 (O_3498,N_29732,N_29639);
nor UO_3499 (O_3499,N_29780,N_29873);
endmodule