module basic_1000_10000_1500_100_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_322,In_586);
nor U1 (N_1,In_506,In_926);
nor U2 (N_2,In_587,In_570);
and U3 (N_3,In_44,In_574);
or U4 (N_4,In_326,In_170);
nand U5 (N_5,In_997,In_627);
nor U6 (N_6,In_771,In_411);
and U7 (N_7,In_466,In_48);
nand U8 (N_8,In_999,In_38);
or U9 (N_9,In_367,In_550);
nand U10 (N_10,In_385,In_85);
nand U11 (N_11,In_37,In_73);
and U12 (N_12,In_118,In_484);
or U13 (N_13,In_14,In_715);
nor U14 (N_14,In_952,In_507);
or U15 (N_15,In_60,In_329);
and U16 (N_16,In_207,In_799);
nor U17 (N_17,In_689,In_16);
or U18 (N_18,In_529,In_876);
nor U19 (N_19,In_553,In_872);
or U20 (N_20,In_439,In_103);
or U21 (N_21,In_323,In_959);
nand U22 (N_22,In_998,In_815);
nor U23 (N_23,In_943,In_105);
nor U24 (N_24,In_432,In_179);
xnor U25 (N_25,In_348,In_899);
xor U26 (N_26,In_729,In_620);
nand U27 (N_27,In_679,In_781);
nand U28 (N_28,In_410,In_857);
and U29 (N_29,In_615,In_919);
and U30 (N_30,In_523,In_483);
nor U31 (N_31,In_871,In_164);
or U32 (N_32,In_23,In_752);
nor U33 (N_33,In_652,In_158);
or U34 (N_34,In_783,In_306);
nand U35 (N_35,In_903,In_624);
nor U36 (N_36,In_218,In_901);
and U37 (N_37,In_127,In_236);
and U38 (N_38,In_528,In_989);
nand U39 (N_39,In_223,In_535);
nand U40 (N_40,In_626,In_101);
nor U41 (N_41,In_55,In_547);
and U42 (N_42,In_971,In_471);
nor U43 (N_43,In_81,In_667);
and U44 (N_44,In_635,In_569);
nand U45 (N_45,In_212,In_182);
nor U46 (N_46,In_677,In_774);
xor U47 (N_47,In_548,In_109);
or U48 (N_48,In_923,In_59);
xnor U49 (N_49,In_345,In_437);
and U50 (N_50,In_246,In_925);
nor U51 (N_51,In_724,In_993);
nand U52 (N_52,In_660,In_392);
and U53 (N_53,In_585,In_363);
nand U54 (N_54,In_864,In_769);
or U55 (N_55,In_169,In_650);
nand U56 (N_56,In_451,In_247);
nor U57 (N_57,In_756,In_958);
and U58 (N_58,In_669,In_57);
nor U59 (N_59,In_922,In_195);
or U60 (N_60,In_708,In_163);
and U61 (N_61,In_690,In_65);
and U62 (N_62,In_955,In_350);
nor U63 (N_63,In_893,In_803);
and U64 (N_64,In_421,In_792);
or U65 (N_65,In_382,In_371);
and U66 (N_66,In_753,In_777);
nor U67 (N_67,In_859,In_688);
nand U68 (N_68,In_510,In_237);
nand U69 (N_69,In_716,In_456);
nor U70 (N_70,In_389,In_545);
nand U71 (N_71,In_744,In_134);
and U72 (N_72,In_53,In_987);
nand U73 (N_73,In_417,In_111);
nor U74 (N_74,In_379,In_654);
or U75 (N_75,In_469,In_914);
nor U76 (N_76,In_668,In_400);
nand U77 (N_77,In_339,In_992);
and U78 (N_78,In_3,In_242);
nor U79 (N_79,In_848,In_968);
nand U80 (N_80,In_648,In_333);
nand U81 (N_81,In_147,In_427);
or U82 (N_82,In_796,In_892);
nand U83 (N_83,In_356,In_274);
and U84 (N_84,In_67,In_413);
nor U85 (N_85,In_470,In_945);
or U86 (N_86,In_50,In_646);
nand U87 (N_87,In_167,In_593);
or U88 (N_88,In_25,In_687);
or U89 (N_89,In_36,In_184);
nand U90 (N_90,In_407,In_79);
nor U91 (N_91,In_293,In_592);
or U92 (N_92,In_283,In_558);
or U93 (N_93,In_565,In_349);
nand U94 (N_94,In_359,In_328);
nor U95 (N_95,In_622,In_80);
nor U96 (N_96,In_509,In_397);
or U97 (N_97,In_493,In_768);
nand U98 (N_98,In_970,In_860);
nor U99 (N_99,In_233,In_152);
and U100 (N_100,In_964,In_836);
xor U101 (N_101,In_807,N_96);
and U102 (N_102,In_730,In_215);
nand U103 (N_103,In_946,In_176);
nor U104 (N_104,In_633,In_994);
nand U105 (N_105,In_288,In_938);
or U106 (N_106,In_291,In_825);
or U107 (N_107,In_866,In_555);
or U108 (N_108,In_281,In_540);
nand U109 (N_109,In_880,In_542);
and U110 (N_110,In_702,In_721);
or U111 (N_111,In_598,In_108);
or U112 (N_112,In_601,In_603);
xor U113 (N_113,In_608,In_775);
or U114 (N_114,In_967,In_537);
or U115 (N_115,In_351,In_129);
and U116 (N_116,In_696,N_64);
xnor U117 (N_117,In_831,In_891);
nor U118 (N_118,In_556,In_699);
nor U119 (N_119,In_638,In_915);
and U120 (N_120,In_568,In_415);
or U121 (N_121,In_953,In_186);
and U122 (N_122,In_606,In_793);
and U123 (N_123,In_849,In_671);
nor U124 (N_124,In_957,In_941);
nor U125 (N_125,N_39,In_745);
nand U126 (N_126,In_91,In_512);
or U127 (N_127,In_643,In_858);
nand U128 (N_128,In_34,In_995);
nor U129 (N_129,In_374,In_496);
and U130 (N_130,N_28,In_227);
nand U131 (N_131,In_468,In_855);
and U132 (N_132,In_980,In_942);
nor U133 (N_133,N_9,N_59);
or U134 (N_134,In_861,In_817);
nand U135 (N_135,In_181,In_243);
nor U136 (N_136,In_431,In_444);
nor U137 (N_137,In_875,In_112);
or U138 (N_138,In_827,In_700);
or U139 (N_139,In_611,In_578);
and U140 (N_140,In_674,In_882);
or U141 (N_141,In_106,In_384);
and U142 (N_142,In_984,In_634);
and U143 (N_143,In_494,In_972);
or U144 (N_144,N_51,In_452);
nor U145 (N_145,N_43,In_114);
or U146 (N_146,In_779,N_37);
or U147 (N_147,In_697,In_965);
nand U148 (N_148,In_380,In_948);
or U149 (N_149,In_758,In_352);
nor U150 (N_150,N_94,In_904);
or U151 (N_151,In_29,In_813);
and U152 (N_152,In_762,In_124);
or U153 (N_153,In_589,In_704);
nor U154 (N_154,N_0,In_560);
and U155 (N_155,In_805,In_185);
or U156 (N_156,In_200,In_388);
nor U157 (N_157,N_46,In_364);
and U158 (N_158,In_479,In_932);
nor U159 (N_159,In_303,In_641);
and U160 (N_160,In_913,In_617);
nor U161 (N_161,N_24,In_368);
and U162 (N_162,In_950,In_712);
or U163 (N_163,In_406,In_686);
or U164 (N_164,In_433,In_773);
nand U165 (N_165,In_463,In_354);
or U166 (N_166,In_12,In_714);
nand U167 (N_167,In_8,In_40);
nor U168 (N_168,In_282,In_315);
xnor U169 (N_169,In_436,In_629);
or U170 (N_170,In_360,N_4);
nor U171 (N_171,In_180,In_647);
or U172 (N_172,N_86,In_670);
and U173 (N_173,In_318,In_273);
nand U174 (N_174,In_330,N_22);
and U175 (N_175,In_100,In_319);
nand U176 (N_176,In_564,In_69);
nor U177 (N_177,In_41,In_331);
nor U178 (N_178,In_940,In_21);
nor U179 (N_179,In_325,N_26);
or U180 (N_180,In_149,In_151);
and U181 (N_181,In_597,In_202);
nand U182 (N_182,N_89,In_344);
nand U183 (N_183,In_455,In_961);
or U184 (N_184,In_132,In_720);
xor U185 (N_185,In_187,In_511);
or U186 (N_186,In_912,In_666);
and U187 (N_187,In_599,In_743);
nor U188 (N_188,In_175,In_673);
and U189 (N_189,In_314,N_97);
or U190 (N_190,In_250,In_265);
or U191 (N_191,N_84,In_226);
xor U192 (N_192,In_458,In_517);
and U193 (N_193,N_11,In_10);
nand U194 (N_194,In_403,In_270);
nor U195 (N_195,N_13,In_557);
nor U196 (N_196,In_935,N_36);
or U197 (N_197,N_98,N_87);
nand U198 (N_198,In_962,In_676);
and U199 (N_199,In_18,In_373);
or U200 (N_200,In_188,In_695);
nand U201 (N_201,N_82,In_486);
xor U202 (N_202,N_106,N_115);
and U203 (N_203,In_56,In_54);
or U204 (N_204,In_271,N_185);
nor U205 (N_205,N_188,In_429);
nor U206 (N_206,In_430,In_409);
or U207 (N_207,N_129,In_161);
nor U208 (N_208,In_931,In_275);
nor U209 (N_209,In_257,N_147);
nor U210 (N_210,In_990,In_541);
and U211 (N_211,In_764,N_47);
and U212 (N_212,In_838,In_530);
nand U213 (N_213,In_358,N_179);
or U214 (N_214,In_304,In_513);
or U215 (N_215,In_137,In_934);
and U216 (N_216,In_881,In_613);
nand U217 (N_217,N_79,In_311);
xnor U218 (N_218,In_802,In_278);
and U219 (N_219,N_139,In_818);
nor U220 (N_220,N_85,In_165);
and U221 (N_221,In_631,In_736);
nand U222 (N_222,In_832,In_798);
or U223 (N_223,In_898,N_182);
nand U224 (N_224,In_947,In_778);
nand U225 (N_225,In_614,N_121);
nor U226 (N_226,In_27,In_300);
nor U227 (N_227,In_518,N_180);
nand U228 (N_228,In_71,N_165);
nand U229 (N_229,N_23,In_317);
or U230 (N_230,In_131,In_682);
or U231 (N_231,In_390,In_154);
or U232 (N_232,In_581,In_464);
or U233 (N_233,In_604,In_297);
nand U234 (N_234,In_795,In_692);
and U235 (N_235,In_896,In_683);
nor U236 (N_236,In_797,In_133);
nor U237 (N_237,In_765,In_809);
nor U238 (N_238,N_48,In_991);
and U239 (N_239,In_199,In_307);
and U240 (N_240,N_170,In_9);
nor U241 (N_241,In_562,In_974);
and U242 (N_242,In_378,In_96);
nand U243 (N_243,In_508,In_782);
nand U244 (N_244,In_874,N_41);
nor U245 (N_245,In_357,In_424);
and U246 (N_246,In_75,In_684);
nand U247 (N_247,In_787,N_25);
or U248 (N_248,N_159,In_301);
or U249 (N_249,In_289,In_299);
or U250 (N_250,In_693,In_873);
and U251 (N_251,In_976,In_637);
or U252 (N_252,N_137,In_728);
and U253 (N_253,N_80,In_747);
or U254 (N_254,In_482,N_162);
nand U255 (N_255,In_391,N_8);
nor U256 (N_256,In_543,In_885);
nor U257 (N_257,In_240,In_123);
and U258 (N_258,In_918,In_110);
or U259 (N_259,N_101,In_956);
nand U260 (N_260,N_160,In_70);
nand U261 (N_261,In_6,In_655);
and U262 (N_262,In_751,In_732);
or U263 (N_263,N_44,N_138);
or U264 (N_264,In_830,In_639);
xor U265 (N_265,In_534,In_750);
or U266 (N_266,N_184,N_126);
and U267 (N_267,In_495,In_895);
and U268 (N_268,N_181,In_996);
nand U269 (N_269,In_746,N_81);
or U270 (N_270,In_571,In_924);
or U271 (N_271,In_723,In_538);
nand U272 (N_272,In_183,N_93);
and U273 (N_273,N_154,In_524);
nand U274 (N_274,N_142,N_100);
or U275 (N_275,In_74,N_175);
and U276 (N_276,In_766,In_786);
nand U277 (N_277,In_381,In_710);
nor U278 (N_278,In_285,In_969);
nand U279 (N_279,In_2,In_393);
nor U280 (N_280,In_986,In_135);
or U281 (N_281,In_717,In_814);
or U282 (N_282,In_930,In_203);
nor U283 (N_283,In_840,In_31);
and U284 (N_284,N_141,In_890);
or U285 (N_285,In_536,N_54);
nor U286 (N_286,In_951,In_155);
or U287 (N_287,In_13,N_34);
nor U288 (N_288,N_15,In_168);
nor U289 (N_289,In_204,In_761);
and U290 (N_290,N_73,In_804);
nand U291 (N_291,In_425,In_93);
nor U292 (N_292,In_49,In_475);
or U293 (N_293,In_362,In_192);
or U294 (N_294,In_228,In_42);
nor U295 (N_295,N_134,In_981);
and U296 (N_296,N_19,N_151);
or U297 (N_297,N_144,In_272);
or U298 (N_298,In_691,In_78);
nor U299 (N_299,In_474,In_121);
nand U300 (N_300,In_573,In_28);
nand U301 (N_301,N_261,In_988);
or U302 (N_302,N_291,N_239);
nand U303 (N_303,In_707,In_706);
nor U304 (N_304,In_651,N_274);
and U305 (N_305,In_178,In_440);
nor U306 (N_306,N_225,N_190);
nand U307 (N_307,N_266,In_166);
nor U308 (N_308,N_247,In_286);
nor U309 (N_309,In_850,In_102);
and U310 (N_310,In_209,In_190);
and U311 (N_311,In_780,N_227);
nand U312 (N_312,N_206,In_869);
nor U313 (N_313,In_72,In_902);
or U314 (N_314,In_159,In_812);
and U315 (N_315,In_316,In_84);
and U316 (N_316,In_929,In_465);
or U317 (N_317,In_77,N_199);
or U318 (N_318,In_162,In_544);
and U319 (N_319,In_198,N_150);
or U320 (N_320,In_757,In_519);
and U321 (N_321,N_284,In_739);
or U322 (N_322,N_187,In_577);
and U323 (N_323,In_148,In_255);
nand U324 (N_324,In_321,In_395);
or U325 (N_325,In_741,N_245);
or U326 (N_326,In_143,In_98);
or U327 (N_327,In_434,In_423);
nor U328 (N_328,N_169,In_399);
and U329 (N_329,In_24,In_174);
nand U330 (N_330,In_579,In_20);
or U331 (N_331,N_168,N_265);
nand U332 (N_332,In_632,In_298);
or U333 (N_333,N_166,In_467);
nand U334 (N_334,In_933,In_454);
nor U335 (N_335,In_709,In_561);
or U336 (N_336,N_208,In_879);
and U337 (N_337,In_917,In_828);
nor U338 (N_338,In_920,In_841);
or U339 (N_339,In_435,In_334);
and U340 (N_340,In_826,In_210);
nand U341 (N_341,In_906,In_711);
or U342 (N_342,N_297,N_217);
nand U343 (N_343,In_623,In_92);
nor U344 (N_344,In_488,N_125);
nor U345 (N_345,In_816,In_894);
nand U346 (N_346,In_449,N_289);
and U347 (N_347,In_835,N_242);
nor U348 (N_348,In_794,In_126);
or U349 (N_349,In_269,In_759);
and U350 (N_350,In_921,N_83);
nor U351 (N_351,In_239,N_211);
and U352 (N_352,N_109,N_95);
and U353 (N_353,N_71,In_944);
nor U354 (N_354,In_414,In_115);
or U355 (N_355,N_228,N_62);
and U356 (N_356,In_591,N_244);
nand U357 (N_357,In_86,In_822);
and U358 (N_358,In_267,In_33);
or U359 (N_359,N_108,In_173);
and U360 (N_360,In_7,N_102);
nor U361 (N_361,In_656,In_909);
nand U362 (N_362,In_575,In_268);
nand U363 (N_363,In_563,In_229);
or U364 (N_364,In_477,In_490);
and U365 (N_365,N_7,In_338);
nor U366 (N_366,N_75,N_191);
and U367 (N_367,In_370,N_233);
and U368 (N_368,In_99,In_128);
nor U369 (N_369,In_602,In_837);
and U370 (N_370,N_249,N_212);
nand U371 (N_371,N_173,N_88);
and U372 (N_372,N_223,N_197);
and U373 (N_373,In_884,In_936);
nor U374 (N_374,In_854,N_260);
and U375 (N_375,In_749,In_680);
xor U376 (N_376,In_487,In_422);
nand U377 (N_377,In_43,In_305);
nand U378 (N_378,In_95,In_453);
nand U379 (N_379,N_280,In_788);
nand U380 (N_380,N_248,N_196);
nand U381 (N_381,In_960,In_438);
or U382 (N_382,N_153,N_61);
or U383 (N_383,In_618,N_273);
and U384 (N_384,N_278,N_72);
or U385 (N_385,In_658,In_985);
and U386 (N_386,In_302,In_90);
or U387 (N_387,In_621,N_282);
and U388 (N_388,In_785,N_292);
or U389 (N_389,In_249,In_515);
nor U390 (N_390,In_460,N_234);
nand U391 (N_391,N_112,In_46);
nand U392 (N_392,N_268,In_734);
or U393 (N_393,In_489,N_238);
nand U394 (N_394,N_178,In_402);
or U395 (N_395,N_183,In_327);
or U396 (N_396,In_824,In_979);
nand U397 (N_397,N_250,In_26);
nor U398 (N_398,In_863,N_91);
or U399 (N_399,In_220,In_258);
nor U400 (N_400,N_113,In_366);
nand U401 (N_401,In_642,In_52);
nor U402 (N_402,In_398,N_92);
and U403 (N_403,In_516,In_446);
nor U404 (N_404,In_141,N_322);
nor U405 (N_405,In_221,N_52);
nand U406 (N_406,N_343,N_210);
nor U407 (N_407,N_381,In_726);
nor U408 (N_408,In_549,N_99);
and U409 (N_409,N_65,N_334);
nand U410 (N_410,In_284,N_321);
nor U411 (N_411,In_476,In_653);
or U412 (N_412,N_345,In_313);
and U413 (N_413,In_588,N_16);
nor U414 (N_414,N_77,N_171);
or U415 (N_415,In_412,In_851);
nor U416 (N_416,In_76,N_114);
nor U417 (N_417,In_663,In_448);
xor U418 (N_418,N_246,In_865);
nand U419 (N_419,N_376,N_104);
nand U420 (N_420,In_264,N_389);
nor U421 (N_421,N_146,N_222);
nor U422 (N_422,In_526,N_257);
nand U423 (N_423,In_843,In_58);
or U424 (N_424,N_5,N_386);
nor U425 (N_425,N_226,N_241);
and U426 (N_426,N_17,N_313);
or U427 (N_427,In_485,N_374);
and U428 (N_428,In_619,In_808);
and U429 (N_429,N_269,N_213);
nor U430 (N_430,N_304,N_35);
nand U431 (N_431,N_362,In_566);
and U432 (N_432,In_262,In_790);
nor U433 (N_433,N_58,In_125);
or U434 (N_434,In_292,In_87);
nand U435 (N_435,N_21,N_349);
nand U436 (N_436,N_375,In_733);
and U437 (N_437,In_583,N_136);
nand U438 (N_438,In_441,In_612);
and U439 (N_439,In_117,N_209);
nor U440 (N_440,In_554,In_88);
nand U441 (N_441,In_616,In_294);
or U442 (N_442,In_296,In_206);
nand U443 (N_443,In_905,In_61);
nand U444 (N_444,N_368,N_359);
nand U445 (N_445,N_255,N_148);
nor U446 (N_446,In_954,In_823);
and U447 (N_447,N_366,In_145);
nor U448 (N_448,In_156,In_396);
nand U449 (N_449,In_442,N_279);
or U450 (N_450,In_657,In_644);
and U451 (N_451,N_352,N_111);
and U452 (N_452,N_336,In_630);
nor U453 (N_453,In_335,N_164);
and U454 (N_454,In_640,In_539);
nor U455 (N_455,In_63,In_461);
nand U456 (N_456,N_330,N_90);
and U457 (N_457,In_120,In_844);
nor U458 (N_458,N_306,In_32);
or U459 (N_459,In_675,In_900);
or U460 (N_460,N_218,N_326);
and U461 (N_461,In_908,In_767);
or U462 (N_462,N_276,In_551);
nand U463 (N_463,In_820,In_500);
or U464 (N_464,In_982,N_42);
and U465 (N_465,In_62,In_232);
or U466 (N_466,N_78,N_207);
or U467 (N_467,In_681,In_341);
nand U468 (N_468,N_315,In_763);
nand U469 (N_469,In_870,In_64);
or U470 (N_470,N_329,In_138);
nand U471 (N_471,N_384,In_244);
or U472 (N_472,N_385,In_191);
or U473 (N_473,In_251,In_625);
or U474 (N_474,In_238,N_117);
nor U475 (N_475,In_846,In_355);
nand U476 (N_476,In_116,In_277);
nor U477 (N_477,In_705,N_288);
nand U478 (N_478,In_83,In_829);
nor U479 (N_479,In_1,In_525);
and U480 (N_480,In_290,In_340);
nor U481 (N_481,In_552,N_320);
and U482 (N_482,N_286,In_531);
nand U483 (N_483,In_222,N_123);
nor U484 (N_484,N_29,N_333);
or U485 (N_485,N_49,In_214);
or U486 (N_486,In_737,In_386);
nor U487 (N_487,In_559,In_256);
and U488 (N_488,N_202,In_770);
nand U489 (N_489,In_201,In_231);
or U490 (N_490,N_296,In_834);
nor U491 (N_491,N_363,N_360);
nor U492 (N_492,In_791,In_372);
or U493 (N_493,N_231,In_343);
and U494 (N_494,N_355,In_819);
nor U495 (N_495,In_665,N_299);
nand U496 (N_496,In_731,N_172);
nand U497 (N_497,In_320,In_261);
nand U498 (N_498,N_232,In_722);
nand U499 (N_499,In_276,In_862);
or U500 (N_500,N_411,In_19);
and U501 (N_501,In_607,N_237);
or U502 (N_502,N_294,N_356);
or U503 (N_503,N_124,N_14);
and U504 (N_504,N_397,N_174);
or U505 (N_505,In_113,N_335);
or U506 (N_506,N_358,N_192);
or U507 (N_507,In_983,N_451);
and U508 (N_508,In_718,In_949);
nor U509 (N_509,N_462,In_939);
and U510 (N_510,In_47,In_755);
and U511 (N_511,In_784,In_480);
and U512 (N_512,N_373,N_383);
and U513 (N_513,N_413,N_69);
and U514 (N_514,N_295,In_889);
and U515 (N_515,N_470,In_89);
and U516 (N_516,N_391,N_454);
or U517 (N_517,In_975,N_444);
and U518 (N_518,In_252,In_408);
and U519 (N_519,In_609,In_977);
or U520 (N_520,N_388,In_473);
or U521 (N_521,In_595,In_230);
nor U522 (N_522,In_800,In_678);
or U523 (N_523,N_132,N_449);
and U524 (N_524,N_177,In_22);
nor U525 (N_525,N_33,N_230);
or U526 (N_526,N_493,In_418);
nand U527 (N_527,N_434,N_476);
and U528 (N_528,N_221,N_394);
nand U529 (N_529,In_194,N_40);
nor U530 (N_530,In_505,N_145);
and U531 (N_531,In_172,N_382);
nor U532 (N_532,N_157,In_39);
nor U533 (N_533,In_157,In_886);
nand U534 (N_534,N_473,N_435);
and U535 (N_535,In_789,N_203);
nor U536 (N_536,In_478,N_195);
and U537 (N_537,In_104,N_68);
or U538 (N_538,In_916,N_216);
nor U539 (N_539,In_17,N_425);
nand U540 (N_540,N_156,N_310);
and U541 (N_541,In_727,N_272);
nand U542 (N_542,In_82,N_448);
or U543 (N_543,N_364,In_346);
nand U544 (N_544,N_457,N_204);
and U545 (N_545,N_402,N_472);
or U546 (N_546,In_140,In_754);
nor U547 (N_547,N_18,N_403);
nand U548 (N_548,In_502,In_907);
and U549 (N_549,N_458,N_478);
or U550 (N_550,N_133,N_460);
nor U551 (N_551,N_423,N_452);
or U552 (N_552,N_419,In_853);
and U553 (N_553,In_821,N_420);
nand U554 (N_554,N_12,N_463);
or U555 (N_555,In_738,N_259);
and U556 (N_556,N_285,In_937);
nor U557 (N_557,N_263,In_594);
or U558 (N_558,N_465,N_371);
nand U559 (N_559,In_719,In_801);
and U560 (N_560,In_887,N_428);
and U561 (N_561,N_324,In_845);
and U562 (N_562,N_401,N_135);
nand U563 (N_563,N_287,N_131);
and U564 (N_564,In_522,In_521);
nor U565 (N_565,N_152,In_694);
nand U566 (N_566,In_309,In_501);
nand U567 (N_567,In_68,In_94);
nand U568 (N_568,In_582,In_377);
and U569 (N_569,N_293,In_426);
or U570 (N_570,N_367,In_142);
nand U571 (N_571,In_806,N_308);
nand U572 (N_572,N_283,In_600);
and U573 (N_573,N_488,In_193);
or U574 (N_574,N_392,N_468);
and U575 (N_575,In_353,N_387);
nand U576 (N_576,In_0,In_978);
nand U577 (N_577,In_878,In_649);
nor U578 (N_578,In_645,In_234);
nor U579 (N_579,N_447,In_740);
or U580 (N_580,N_490,In_742);
or U581 (N_581,N_446,N_429);
or U582 (N_582,N_353,In_927);
or U583 (N_583,N_219,In_144);
and U584 (N_584,In_661,N_317);
nor U585 (N_585,N_57,In_462);
nor U586 (N_586,In_150,N_455);
and U587 (N_587,N_267,In_225);
nor U588 (N_588,N_432,N_118);
nand U589 (N_589,N_167,In_533);
or U590 (N_590,N_10,In_546);
or U591 (N_591,N_215,N_410);
and U592 (N_592,N_379,In_295);
nor U593 (N_593,N_496,In_605);
or U594 (N_594,In_662,In_491);
and U595 (N_595,N_149,N_486);
and U596 (N_596,N_339,N_497);
nand U597 (N_597,N_254,N_412);
nor U598 (N_598,N_140,N_105);
nor U599 (N_599,In_213,N_395);
and U600 (N_600,N_243,N_404);
nand U601 (N_601,N_122,In_248);
and U602 (N_602,N_553,N_344);
xnor U603 (N_603,N_189,N_564);
xnor U604 (N_604,N_535,In_472);
nor U605 (N_605,N_487,In_208);
nor U606 (N_606,In_139,In_928);
and U607 (N_607,In_833,N_264);
and U608 (N_608,N_55,In_856);
nor U609 (N_609,In_520,N_158);
and U610 (N_610,N_258,N_281);
or U611 (N_611,N_499,N_523);
nor U612 (N_612,N_316,N_433);
and U613 (N_613,N_450,N_549);
nor U614 (N_614,N_348,N_431);
or U615 (N_615,N_60,N_396);
and U616 (N_616,N_307,In_910);
or U617 (N_617,N_116,In_443);
and U618 (N_618,In_504,N_576);
nor U619 (N_619,N_414,N_563);
and U620 (N_620,In_287,N_370);
nor U621 (N_621,In_51,N_3);
nor U622 (N_622,In_254,In_868);
or U623 (N_623,In_867,N_500);
and U624 (N_624,In_572,N_256);
nor U625 (N_625,N_533,N_398);
nand U626 (N_626,N_570,N_445);
nand U627 (N_627,N_474,In_279);
and U628 (N_628,In_659,N_438);
and U629 (N_629,N_505,In_450);
nand U630 (N_630,In_394,In_11);
xnor U631 (N_631,N_441,N_482);
nand U632 (N_632,N_597,N_45);
or U633 (N_633,N_235,N_585);
or U634 (N_634,N_526,N_541);
nor U635 (N_635,N_236,In_383);
nand U636 (N_636,In_205,In_35);
and U637 (N_637,In_725,N_558);
nor U638 (N_638,In_5,In_847);
nand U639 (N_639,N_331,N_305);
nand U640 (N_640,N_53,N_107);
nand U641 (N_641,N_592,N_544);
nand U642 (N_642,N_581,N_504);
nor U643 (N_643,N_580,N_517);
nor U644 (N_644,N_1,N_511);
nand U645 (N_645,N_38,N_303);
nor U646 (N_646,N_214,In_122);
nand U647 (N_647,N_554,N_557);
or U648 (N_648,N_354,In_963);
nand U649 (N_649,N_593,N_566);
and U650 (N_650,N_76,N_312);
nor U651 (N_651,N_2,N_378);
and U652 (N_652,In_216,N_494);
and U653 (N_653,In_211,N_338);
nand U654 (N_654,N_548,N_524);
and U655 (N_655,In_312,In_259);
nor U656 (N_656,In_877,In_160);
or U657 (N_657,In_171,N_270);
nor U658 (N_658,In_576,N_453);
nor U659 (N_659,N_155,In_457);
and U660 (N_660,N_351,N_416);
and U661 (N_661,N_596,In_196);
nand U662 (N_662,N_31,In_153);
nand U663 (N_663,N_514,N_437);
nand U664 (N_664,N_503,In_897);
or U665 (N_665,N_480,N_415);
nand U666 (N_666,In_698,N_584);
nand U667 (N_667,N_572,N_589);
and U668 (N_668,In_701,N_461);
nand U669 (N_669,N_586,N_200);
nor U670 (N_670,N_527,N_464);
nor U671 (N_671,In_107,N_63);
or U672 (N_672,In_636,N_442);
nand U673 (N_673,N_340,N_426);
and U674 (N_674,In_15,N_417);
nor U675 (N_675,N_439,In_361);
or U676 (N_676,N_128,N_271);
or U677 (N_677,In_811,In_241);
nor U678 (N_678,N_498,In_527);
and U679 (N_679,N_555,In_703);
or U680 (N_680,In_369,N_519);
and U681 (N_681,N_440,In_308);
nand U682 (N_682,N_319,N_551);
nor U683 (N_683,N_467,N_30);
nor U684 (N_684,N_127,N_194);
nand U685 (N_685,N_534,N_27);
nor U686 (N_686,N_569,In_310);
and U687 (N_687,N_300,N_357);
nand U688 (N_688,N_537,N_408);
or U689 (N_689,In_197,In_532);
and U690 (N_690,N_422,N_251);
nand U691 (N_691,In_332,In_416);
and U692 (N_692,In_342,N_332);
nand U693 (N_693,In_590,N_475);
or U694 (N_694,In_217,In_177);
nand U695 (N_695,N_318,In_428);
or U696 (N_696,N_484,N_579);
and U697 (N_697,N_545,N_599);
and U698 (N_698,N_516,N_471);
nand U699 (N_699,N_567,In_596);
nand U700 (N_700,N_634,N_528);
or U701 (N_701,N_616,N_590);
nand U702 (N_702,N_510,N_609);
nand U703 (N_703,N_314,In_146);
or U704 (N_704,N_618,N_477);
or U705 (N_705,N_481,N_67);
nor U706 (N_706,N_556,N_622);
nor U707 (N_707,N_103,N_224);
nor U708 (N_708,N_559,N_608);
and U709 (N_709,N_641,N_575);
nand U710 (N_710,N_538,In_672);
and U711 (N_711,In_584,In_280);
and U712 (N_712,N_642,N_636);
nand U713 (N_713,N_669,In_404);
nand U714 (N_714,N_466,N_603);
nand U715 (N_715,N_688,N_540);
and U716 (N_716,N_601,N_492);
or U717 (N_717,N_201,N_650);
or U718 (N_718,N_591,N_687);
nand U719 (N_719,N_604,N_529);
and U720 (N_720,In_337,In_685);
nand U721 (N_721,N_56,N_624);
and U722 (N_722,N_605,In_387);
and U723 (N_723,N_176,N_588);
nand U724 (N_724,N_681,N_518);
nand U725 (N_725,N_653,N_698);
nand U726 (N_726,N_119,N_479);
or U727 (N_727,N_6,N_509);
and U728 (N_728,In_253,N_699);
nor U729 (N_729,N_365,N_436);
or U730 (N_730,N_130,In_189);
nor U731 (N_731,N_623,N_539);
nor U732 (N_732,N_561,N_643);
and U733 (N_733,N_613,N_670);
and U734 (N_734,In_266,In_713);
nand U735 (N_735,N_512,In_136);
and U736 (N_736,N_619,N_507);
or U737 (N_737,N_672,N_685);
and U738 (N_738,In_842,N_400);
nor U739 (N_739,N_328,N_542);
and U740 (N_740,N_418,N_506);
or U741 (N_741,N_627,N_683);
nand U742 (N_742,N_369,N_347);
nand U743 (N_743,N_552,N_501);
nand U744 (N_744,N_565,In_97);
and U745 (N_745,N_667,In_405);
nor U746 (N_746,N_696,N_689);
xor U747 (N_747,N_205,N_649);
nor U748 (N_748,N_405,N_612);
nand U749 (N_749,In_459,N_677);
or U750 (N_750,N_489,N_647);
nor U751 (N_751,In_503,N_652);
nand U752 (N_752,N_676,N_302);
and U753 (N_753,N_372,In_966);
nor U754 (N_754,N_424,N_587);
nand U755 (N_755,N_32,N_323);
or U756 (N_756,N_606,N_607);
or U757 (N_757,N_409,N_684);
or U758 (N_758,In_420,N_240);
nor U759 (N_759,N_655,In_419);
nand U760 (N_760,In_883,N_495);
nor U761 (N_761,N_74,N_421);
and U762 (N_762,N_483,N_393);
nor U763 (N_763,N_678,N_50);
or U764 (N_764,N_668,N_638);
and U765 (N_765,In_445,In_119);
and U766 (N_766,N_143,N_674);
nor U767 (N_767,N_325,N_675);
nand U768 (N_768,In_567,In_888);
nand U769 (N_769,N_691,In_30);
or U770 (N_770,N_262,In_481);
or U771 (N_771,N_546,N_508);
nor U772 (N_772,In_735,N_594);
nor U773 (N_773,N_110,N_502);
nor U774 (N_774,N_380,In_224);
and U775 (N_775,N_620,N_629);
or U776 (N_776,N_161,N_543);
and U777 (N_777,N_631,N_346);
or U778 (N_778,N_513,N_562);
nor U779 (N_779,N_341,N_659);
nor U780 (N_780,N_626,N_578);
or U781 (N_781,N_645,In_497);
nand U782 (N_782,N_377,N_697);
nor U783 (N_783,N_630,N_693);
nor U784 (N_784,N_459,N_309);
and U785 (N_785,N_252,N_686);
nor U786 (N_786,N_491,N_342);
nand U787 (N_787,In_664,In_492);
or U788 (N_788,N_628,N_692);
and U789 (N_789,N_610,N_625);
or U790 (N_790,N_407,In_324);
nand U791 (N_791,N_573,In_628);
or U792 (N_792,N_680,N_666);
nor U793 (N_793,N_399,N_600);
and U794 (N_794,N_644,N_661);
and U795 (N_795,N_637,N_602);
nor U796 (N_796,N_583,N_662);
and U797 (N_797,N_66,N_651);
nor U798 (N_798,In_376,N_337);
or U799 (N_799,In_4,N_547);
nand U800 (N_800,N_361,N_621);
nor U801 (N_801,N_744,N_737);
nand U802 (N_802,N_708,N_763);
or U803 (N_803,N_791,N_783);
or U804 (N_804,N_728,N_747);
nor U805 (N_805,N_735,N_639);
nand U806 (N_806,N_633,N_784);
nand U807 (N_807,N_778,N_712);
nand U808 (N_808,N_720,In_336);
or U809 (N_809,N_617,In_610);
nand U810 (N_810,N_753,N_750);
nand U811 (N_811,In_498,N_530);
nand U812 (N_812,N_719,N_186);
or U813 (N_813,N_787,N_635);
and U814 (N_814,N_198,N_350);
nor U815 (N_815,N_704,N_574);
or U816 (N_816,N_595,N_648);
and U817 (N_817,N_700,N_710);
nand U818 (N_818,N_654,N_739);
nor U819 (N_819,N_390,N_531);
nand U820 (N_820,N_406,N_730);
nand U821 (N_821,In_760,N_752);
nor U822 (N_822,N_755,N_70);
nor U823 (N_823,In_130,N_782);
nand U824 (N_824,N_711,N_718);
nand U825 (N_825,N_797,In_852);
nand U826 (N_826,N_742,N_758);
nor U827 (N_827,N_780,N_777);
nand U828 (N_828,N_770,N_582);
nor U829 (N_829,In_401,In_365);
nand U830 (N_830,N_515,N_275);
or U831 (N_831,N_301,N_290);
or U832 (N_832,In_776,N_764);
xor U833 (N_833,N_795,N_796);
and U834 (N_834,N_701,N_456);
nor U835 (N_835,N_762,N_721);
or U836 (N_836,N_760,N_749);
nor U837 (N_837,In_514,N_658);
or U838 (N_838,N_774,In_911);
and U839 (N_839,N_20,In_839);
nand U840 (N_840,N_705,N_521);
and U841 (N_841,N_786,N_615);
xnor U842 (N_842,N_713,In_748);
nor U843 (N_843,N_731,N_729);
or U844 (N_844,N_727,N_703);
nand U845 (N_845,In_260,In_219);
nor U846 (N_846,In_973,N_550);
or U847 (N_847,In_772,N_776);
nor U848 (N_848,N_788,N_522);
and U849 (N_849,In_375,N_614);
nor U850 (N_850,N_746,N_427);
nand U851 (N_851,N_756,N_779);
nor U852 (N_852,N_430,N_785);
and U853 (N_853,N_793,In_810);
or U854 (N_854,N_560,N_679);
or U855 (N_855,N_706,In_499);
nor U856 (N_856,N_798,N_725);
nor U857 (N_857,In_235,N_657);
nor U858 (N_858,N_520,N_485);
xnor U859 (N_859,N_761,N_714);
nand U860 (N_860,In_347,N_327);
and U861 (N_861,N_740,N_664);
nor U862 (N_862,N_738,N_220);
nor U863 (N_863,N_525,N_702);
or U864 (N_864,N_671,N_775);
and U865 (N_865,N_120,N_748);
xnor U866 (N_866,In_263,N_690);
and U867 (N_867,N_768,N_726);
nor U868 (N_868,N_682,In_45);
nor U869 (N_869,N_646,N_298);
nor U870 (N_870,N_469,N_733);
nand U871 (N_871,N_741,N_722);
nor U872 (N_872,N_759,N_229);
nand U873 (N_873,In_447,N_443);
nand U874 (N_874,N_577,N_598);
and U875 (N_875,N_754,N_571);
nor U876 (N_876,N_789,N_767);
xnor U877 (N_877,N_736,N_766);
or U878 (N_878,N_568,In_580);
nand U879 (N_879,N_794,N_773);
nand U880 (N_880,N_772,N_694);
or U881 (N_881,N_757,N_536);
and U882 (N_882,N_163,In_66);
nor U883 (N_883,N_717,N_673);
xor U884 (N_884,N_724,N_765);
and U885 (N_885,N_665,N_663);
or U886 (N_886,N_695,N_311);
and U887 (N_887,N_771,N_781);
and U888 (N_888,N_769,N_745);
nand U889 (N_889,N_611,N_751);
nor U890 (N_890,N_640,N_660);
nand U891 (N_891,N_790,N_532);
nor U892 (N_892,N_799,N_716);
nor U893 (N_893,N_253,N_715);
nor U894 (N_894,In_245,N_743);
or U895 (N_895,N_193,N_277);
or U896 (N_896,N_734,N_792);
or U897 (N_897,N_707,N_709);
nand U898 (N_898,N_656,N_732);
nand U899 (N_899,N_723,N_632);
nand U900 (N_900,N_880,N_808);
nand U901 (N_901,N_865,N_806);
or U902 (N_902,N_888,N_857);
xor U903 (N_903,N_820,N_801);
or U904 (N_904,N_866,N_870);
or U905 (N_905,N_832,N_815);
or U906 (N_906,N_859,N_856);
nand U907 (N_907,N_894,N_829);
and U908 (N_908,N_884,N_879);
or U909 (N_909,N_862,N_825);
nor U910 (N_910,N_883,N_892);
or U911 (N_911,N_833,N_882);
nor U912 (N_912,N_842,N_896);
nand U913 (N_913,N_837,N_886);
or U914 (N_914,N_813,N_812);
or U915 (N_915,N_868,N_850);
or U916 (N_916,N_867,N_852);
nor U917 (N_917,N_858,N_836);
nor U918 (N_918,N_800,N_840);
nand U919 (N_919,N_847,N_811);
nand U920 (N_920,N_814,N_863);
nand U921 (N_921,N_853,N_843);
and U922 (N_922,N_838,N_891);
nor U923 (N_923,N_875,N_860);
nand U924 (N_924,N_889,N_871);
nand U925 (N_925,N_855,N_826);
and U926 (N_926,N_804,N_873);
or U927 (N_927,N_818,N_869);
nand U928 (N_928,N_827,N_823);
nand U929 (N_929,N_848,N_830);
and U930 (N_930,N_890,N_831);
and U931 (N_931,N_807,N_893);
and U932 (N_932,N_851,N_877);
nor U933 (N_933,N_803,N_817);
and U934 (N_934,N_895,N_874);
nor U935 (N_935,N_898,N_841);
nor U936 (N_936,N_897,N_899);
or U937 (N_937,N_846,N_864);
nand U938 (N_938,N_805,N_810);
or U939 (N_939,N_854,N_849);
nor U940 (N_940,N_839,N_881);
and U941 (N_941,N_824,N_861);
or U942 (N_942,N_821,N_845);
nand U943 (N_943,N_819,N_816);
nand U944 (N_944,N_887,N_802);
nor U945 (N_945,N_822,N_872);
xnor U946 (N_946,N_844,N_835);
nor U947 (N_947,N_834,N_876);
nand U948 (N_948,N_828,N_885);
xor U949 (N_949,N_878,N_809);
nand U950 (N_950,N_878,N_896);
and U951 (N_951,N_886,N_880);
nor U952 (N_952,N_896,N_894);
nand U953 (N_953,N_814,N_875);
and U954 (N_954,N_894,N_841);
nor U955 (N_955,N_822,N_847);
and U956 (N_956,N_830,N_803);
nand U957 (N_957,N_822,N_829);
and U958 (N_958,N_833,N_886);
nand U959 (N_959,N_864,N_835);
nor U960 (N_960,N_836,N_866);
or U961 (N_961,N_869,N_800);
and U962 (N_962,N_857,N_865);
nor U963 (N_963,N_875,N_802);
and U964 (N_964,N_806,N_874);
nand U965 (N_965,N_878,N_850);
nor U966 (N_966,N_890,N_851);
nor U967 (N_967,N_893,N_887);
nor U968 (N_968,N_804,N_869);
nor U969 (N_969,N_859,N_813);
and U970 (N_970,N_875,N_857);
nand U971 (N_971,N_832,N_860);
nor U972 (N_972,N_877,N_854);
or U973 (N_973,N_867,N_832);
nor U974 (N_974,N_833,N_814);
nand U975 (N_975,N_844,N_846);
nand U976 (N_976,N_879,N_802);
nor U977 (N_977,N_867,N_810);
and U978 (N_978,N_874,N_860);
nand U979 (N_979,N_834,N_848);
and U980 (N_980,N_842,N_833);
or U981 (N_981,N_838,N_883);
nand U982 (N_982,N_897,N_881);
nor U983 (N_983,N_806,N_867);
nor U984 (N_984,N_835,N_812);
nor U985 (N_985,N_885,N_847);
nand U986 (N_986,N_849,N_833);
or U987 (N_987,N_835,N_863);
and U988 (N_988,N_828,N_809);
nand U989 (N_989,N_820,N_851);
or U990 (N_990,N_876,N_845);
nand U991 (N_991,N_816,N_851);
and U992 (N_992,N_838,N_802);
nor U993 (N_993,N_881,N_858);
or U994 (N_994,N_878,N_827);
nor U995 (N_995,N_801,N_854);
or U996 (N_996,N_836,N_814);
nand U997 (N_997,N_850,N_894);
or U998 (N_998,N_815,N_800);
xnor U999 (N_999,N_881,N_899);
and U1000 (N_1000,N_980,N_990);
nor U1001 (N_1001,N_991,N_947);
nand U1002 (N_1002,N_920,N_975);
nand U1003 (N_1003,N_905,N_973);
nand U1004 (N_1004,N_908,N_928);
nand U1005 (N_1005,N_996,N_909);
or U1006 (N_1006,N_917,N_986);
and U1007 (N_1007,N_903,N_995);
and U1008 (N_1008,N_981,N_931);
nand U1009 (N_1009,N_988,N_900);
and U1010 (N_1010,N_959,N_925);
nor U1011 (N_1011,N_974,N_957);
nor U1012 (N_1012,N_923,N_932);
and U1013 (N_1013,N_967,N_960);
and U1014 (N_1014,N_944,N_936);
and U1015 (N_1015,N_982,N_979);
or U1016 (N_1016,N_910,N_939);
nand U1017 (N_1017,N_906,N_916);
or U1018 (N_1018,N_966,N_977);
and U1019 (N_1019,N_952,N_914);
nand U1020 (N_1020,N_935,N_956);
and U1021 (N_1021,N_946,N_924);
and U1022 (N_1022,N_976,N_965);
nand U1023 (N_1023,N_915,N_983);
or U1024 (N_1024,N_949,N_941);
nor U1025 (N_1025,N_942,N_971);
or U1026 (N_1026,N_969,N_902);
and U1027 (N_1027,N_921,N_972);
xnor U1028 (N_1028,N_929,N_913);
or U1029 (N_1029,N_955,N_918);
or U1030 (N_1030,N_958,N_911);
or U1031 (N_1031,N_940,N_963);
and U1032 (N_1032,N_951,N_950);
and U1033 (N_1033,N_919,N_953);
and U1034 (N_1034,N_912,N_984);
nand U1035 (N_1035,N_927,N_985);
nor U1036 (N_1036,N_943,N_998);
nor U1037 (N_1037,N_934,N_993);
or U1038 (N_1038,N_954,N_948);
nand U1039 (N_1039,N_968,N_994);
and U1040 (N_1040,N_997,N_901);
nor U1041 (N_1041,N_930,N_961);
or U1042 (N_1042,N_964,N_999);
and U1043 (N_1043,N_962,N_992);
or U1044 (N_1044,N_937,N_926);
nand U1045 (N_1045,N_987,N_945);
and U1046 (N_1046,N_922,N_907);
nand U1047 (N_1047,N_938,N_970);
and U1048 (N_1048,N_933,N_989);
or U1049 (N_1049,N_904,N_978);
nand U1050 (N_1050,N_997,N_923);
nor U1051 (N_1051,N_986,N_914);
and U1052 (N_1052,N_930,N_941);
xnor U1053 (N_1053,N_901,N_923);
or U1054 (N_1054,N_919,N_940);
nor U1055 (N_1055,N_977,N_984);
and U1056 (N_1056,N_938,N_906);
nor U1057 (N_1057,N_915,N_924);
and U1058 (N_1058,N_962,N_959);
and U1059 (N_1059,N_965,N_945);
nand U1060 (N_1060,N_918,N_927);
nor U1061 (N_1061,N_933,N_991);
nor U1062 (N_1062,N_910,N_918);
xnor U1063 (N_1063,N_954,N_943);
or U1064 (N_1064,N_974,N_927);
nand U1065 (N_1065,N_990,N_902);
nor U1066 (N_1066,N_959,N_939);
nor U1067 (N_1067,N_913,N_903);
nand U1068 (N_1068,N_997,N_942);
and U1069 (N_1069,N_999,N_977);
or U1070 (N_1070,N_932,N_935);
nand U1071 (N_1071,N_942,N_969);
or U1072 (N_1072,N_993,N_910);
and U1073 (N_1073,N_959,N_937);
and U1074 (N_1074,N_981,N_954);
nor U1075 (N_1075,N_970,N_963);
nor U1076 (N_1076,N_939,N_940);
xor U1077 (N_1077,N_968,N_955);
nand U1078 (N_1078,N_984,N_963);
or U1079 (N_1079,N_950,N_920);
nor U1080 (N_1080,N_994,N_908);
and U1081 (N_1081,N_957,N_985);
and U1082 (N_1082,N_993,N_909);
nor U1083 (N_1083,N_977,N_944);
or U1084 (N_1084,N_952,N_912);
and U1085 (N_1085,N_988,N_929);
nand U1086 (N_1086,N_960,N_983);
nor U1087 (N_1087,N_994,N_972);
nand U1088 (N_1088,N_909,N_976);
nand U1089 (N_1089,N_986,N_966);
nor U1090 (N_1090,N_933,N_915);
or U1091 (N_1091,N_906,N_994);
xnor U1092 (N_1092,N_992,N_918);
and U1093 (N_1093,N_938,N_951);
or U1094 (N_1094,N_934,N_900);
and U1095 (N_1095,N_967,N_926);
nand U1096 (N_1096,N_915,N_979);
or U1097 (N_1097,N_974,N_918);
nand U1098 (N_1098,N_904,N_966);
or U1099 (N_1099,N_946,N_991);
nor U1100 (N_1100,N_1096,N_1088);
or U1101 (N_1101,N_1087,N_1095);
or U1102 (N_1102,N_1094,N_1069);
nor U1103 (N_1103,N_1015,N_1062);
or U1104 (N_1104,N_1049,N_1039);
and U1105 (N_1105,N_1055,N_1030);
and U1106 (N_1106,N_1053,N_1078);
nand U1107 (N_1107,N_1044,N_1046);
and U1108 (N_1108,N_1074,N_1048);
nand U1109 (N_1109,N_1091,N_1014);
nand U1110 (N_1110,N_1098,N_1029);
nor U1111 (N_1111,N_1083,N_1047);
nor U1112 (N_1112,N_1082,N_1032);
and U1113 (N_1113,N_1072,N_1019);
and U1114 (N_1114,N_1061,N_1017);
xnor U1115 (N_1115,N_1067,N_1013);
nand U1116 (N_1116,N_1097,N_1085);
nand U1117 (N_1117,N_1064,N_1004);
nor U1118 (N_1118,N_1011,N_1057);
and U1119 (N_1119,N_1066,N_1002);
nor U1120 (N_1120,N_1089,N_1045);
nor U1121 (N_1121,N_1076,N_1022);
or U1122 (N_1122,N_1059,N_1028);
nand U1123 (N_1123,N_1040,N_1042);
and U1124 (N_1124,N_1036,N_1050);
and U1125 (N_1125,N_1084,N_1001);
and U1126 (N_1126,N_1023,N_1035);
or U1127 (N_1127,N_1008,N_1092);
nor U1128 (N_1128,N_1081,N_1070);
or U1129 (N_1129,N_1054,N_1007);
nor U1130 (N_1130,N_1021,N_1026);
and U1131 (N_1131,N_1003,N_1012);
and U1132 (N_1132,N_1024,N_1060);
or U1133 (N_1133,N_1058,N_1051);
and U1134 (N_1134,N_1068,N_1065);
nand U1135 (N_1135,N_1080,N_1075);
nand U1136 (N_1136,N_1031,N_1016);
xor U1137 (N_1137,N_1010,N_1000);
nor U1138 (N_1138,N_1020,N_1090);
nand U1139 (N_1139,N_1079,N_1071);
or U1140 (N_1140,N_1025,N_1038);
nor U1141 (N_1141,N_1034,N_1027);
nor U1142 (N_1142,N_1093,N_1033);
nand U1143 (N_1143,N_1037,N_1052);
nor U1144 (N_1144,N_1005,N_1086);
and U1145 (N_1145,N_1018,N_1099);
nor U1146 (N_1146,N_1077,N_1009);
and U1147 (N_1147,N_1043,N_1041);
nand U1148 (N_1148,N_1056,N_1073);
or U1149 (N_1149,N_1006,N_1063);
or U1150 (N_1150,N_1058,N_1024);
or U1151 (N_1151,N_1092,N_1061);
nor U1152 (N_1152,N_1029,N_1077);
or U1153 (N_1153,N_1072,N_1018);
nand U1154 (N_1154,N_1008,N_1030);
nand U1155 (N_1155,N_1061,N_1005);
nor U1156 (N_1156,N_1091,N_1089);
or U1157 (N_1157,N_1030,N_1044);
nand U1158 (N_1158,N_1044,N_1076);
or U1159 (N_1159,N_1008,N_1009);
nor U1160 (N_1160,N_1077,N_1038);
or U1161 (N_1161,N_1079,N_1064);
and U1162 (N_1162,N_1006,N_1002);
nor U1163 (N_1163,N_1011,N_1068);
and U1164 (N_1164,N_1034,N_1020);
or U1165 (N_1165,N_1087,N_1085);
or U1166 (N_1166,N_1006,N_1011);
or U1167 (N_1167,N_1058,N_1064);
and U1168 (N_1168,N_1042,N_1054);
and U1169 (N_1169,N_1026,N_1028);
or U1170 (N_1170,N_1001,N_1077);
nor U1171 (N_1171,N_1049,N_1014);
or U1172 (N_1172,N_1006,N_1069);
nor U1173 (N_1173,N_1029,N_1059);
or U1174 (N_1174,N_1013,N_1099);
nor U1175 (N_1175,N_1008,N_1058);
and U1176 (N_1176,N_1047,N_1072);
nand U1177 (N_1177,N_1083,N_1098);
or U1178 (N_1178,N_1054,N_1058);
or U1179 (N_1179,N_1019,N_1080);
nor U1180 (N_1180,N_1039,N_1074);
or U1181 (N_1181,N_1093,N_1066);
nand U1182 (N_1182,N_1041,N_1080);
or U1183 (N_1183,N_1096,N_1037);
and U1184 (N_1184,N_1047,N_1011);
or U1185 (N_1185,N_1068,N_1009);
nand U1186 (N_1186,N_1030,N_1099);
and U1187 (N_1187,N_1017,N_1082);
or U1188 (N_1188,N_1042,N_1022);
or U1189 (N_1189,N_1042,N_1071);
nand U1190 (N_1190,N_1065,N_1056);
or U1191 (N_1191,N_1033,N_1047);
or U1192 (N_1192,N_1095,N_1082);
and U1193 (N_1193,N_1030,N_1019);
nand U1194 (N_1194,N_1065,N_1091);
nor U1195 (N_1195,N_1031,N_1064);
nor U1196 (N_1196,N_1004,N_1017);
and U1197 (N_1197,N_1017,N_1024);
nor U1198 (N_1198,N_1070,N_1041);
or U1199 (N_1199,N_1028,N_1074);
nand U1200 (N_1200,N_1183,N_1129);
nor U1201 (N_1201,N_1135,N_1118);
nor U1202 (N_1202,N_1112,N_1159);
nand U1203 (N_1203,N_1138,N_1179);
and U1204 (N_1204,N_1160,N_1102);
or U1205 (N_1205,N_1143,N_1104);
and U1206 (N_1206,N_1165,N_1117);
nand U1207 (N_1207,N_1174,N_1126);
nor U1208 (N_1208,N_1109,N_1154);
and U1209 (N_1209,N_1161,N_1125);
xor U1210 (N_1210,N_1172,N_1144);
or U1211 (N_1211,N_1173,N_1195);
and U1212 (N_1212,N_1140,N_1127);
nor U1213 (N_1213,N_1170,N_1193);
xnor U1214 (N_1214,N_1142,N_1101);
and U1215 (N_1215,N_1194,N_1151);
and U1216 (N_1216,N_1164,N_1198);
or U1217 (N_1217,N_1175,N_1185);
or U1218 (N_1218,N_1106,N_1168);
nor U1219 (N_1219,N_1110,N_1178);
and U1220 (N_1220,N_1149,N_1136);
or U1221 (N_1221,N_1191,N_1124);
nor U1222 (N_1222,N_1116,N_1184);
or U1223 (N_1223,N_1114,N_1197);
nor U1224 (N_1224,N_1176,N_1148);
and U1225 (N_1225,N_1181,N_1177);
or U1226 (N_1226,N_1163,N_1186);
and U1227 (N_1227,N_1133,N_1108);
or U1228 (N_1228,N_1146,N_1166);
nand U1229 (N_1229,N_1100,N_1119);
nand U1230 (N_1230,N_1131,N_1162);
and U1231 (N_1231,N_1105,N_1171);
and U1232 (N_1232,N_1167,N_1115);
nand U1233 (N_1233,N_1187,N_1134);
nor U1234 (N_1234,N_1123,N_1113);
nand U1235 (N_1235,N_1111,N_1190);
nand U1236 (N_1236,N_1132,N_1130);
or U1237 (N_1237,N_1182,N_1121);
nand U1238 (N_1238,N_1152,N_1158);
or U1239 (N_1239,N_1147,N_1188);
or U1240 (N_1240,N_1155,N_1199);
and U1241 (N_1241,N_1150,N_1196);
nor U1242 (N_1242,N_1128,N_1122);
and U1243 (N_1243,N_1169,N_1157);
or U1244 (N_1244,N_1139,N_1189);
nand U1245 (N_1245,N_1145,N_1141);
nand U1246 (N_1246,N_1107,N_1137);
and U1247 (N_1247,N_1192,N_1153);
or U1248 (N_1248,N_1180,N_1120);
nand U1249 (N_1249,N_1103,N_1156);
and U1250 (N_1250,N_1165,N_1172);
xnor U1251 (N_1251,N_1173,N_1188);
nand U1252 (N_1252,N_1196,N_1119);
or U1253 (N_1253,N_1148,N_1199);
nand U1254 (N_1254,N_1126,N_1120);
or U1255 (N_1255,N_1117,N_1121);
or U1256 (N_1256,N_1158,N_1121);
or U1257 (N_1257,N_1185,N_1195);
nand U1258 (N_1258,N_1115,N_1168);
nand U1259 (N_1259,N_1145,N_1153);
and U1260 (N_1260,N_1185,N_1163);
nor U1261 (N_1261,N_1138,N_1145);
nor U1262 (N_1262,N_1189,N_1113);
nor U1263 (N_1263,N_1189,N_1178);
or U1264 (N_1264,N_1166,N_1138);
nor U1265 (N_1265,N_1106,N_1167);
nand U1266 (N_1266,N_1135,N_1191);
and U1267 (N_1267,N_1156,N_1154);
nor U1268 (N_1268,N_1191,N_1173);
and U1269 (N_1269,N_1173,N_1194);
and U1270 (N_1270,N_1101,N_1195);
and U1271 (N_1271,N_1113,N_1198);
nand U1272 (N_1272,N_1126,N_1140);
xor U1273 (N_1273,N_1118,N_1193);
xnor U1274 (N_1274,N_1139,N_1190);
nand U1275 (N_1275,N_1105,N_1186);
or U1276 (N_1276,N_1147,N_1110);
xnor U1277 (N_1277,N_1119,N_1122);
and U1278 (N_1278,N_1136,N_1193);
or U1279 (N_1279,N_1168,N_1188);
nand U1280 (N_1280,N_1166,N_1185);
nor U1281 (N_1281,N_1123,N_1127);
or U1282 (N_1282,N_1123,N_1164);
nand U1283 (N_1283,N_1137,N_1198);
and U1284 (N_1284,N_1121,N_1161);
nand U1285 (N_1285,N_1150,N_1142);
nor U1286 (N_1286,N_1150,N_1165);
nand U1287 (N_1287,N_1157,N_1193);
nand U1288 (N_1288,N_1198,N_1121);
or U1289 (N_1289,N_1176,N_1193);
or U1290 (N_1290,N_1106,N_1169);
and U1291 (N_1291,N_1113,N_1126);
nor U1292 (N_1292,N_1102,N_1161);
and U1293 (N_1293,N_1162,N_1158);
and U1294 (N_1294,N_1128,N_1142);
or U1295 (N_1295,N_1121,N_1116);
nand U1296 (N_1296,N_1104,N_1144);
nor U1297 (N_1297,N_1184,N_1113);
nand U1298 (N_1298,N_1193,N_1148);
and U1299 (N_1299,N_1164,N_1148);
or U1300 (N_1300,N_1239,N_1218);
or U1301 (N_1301,N_1261,N_1237);
nand U1302 (N_1302,N_1251,N_1270);
or U1303 (N_1303,N_1200,N_1243);
nand U1304 (N_1304,N_1230,N_1227);
nor U1305 (N_1305,N_1296,N_1273);
and U1306 (N_1306,N_1269,N_1244);
or U1307 (N_1307,N_1286,N_1284);
nand U1308 (N_1308,N_1206,N_1264);
and U1309 (N_1309,N_1258,N_1257);
nor U1310 (N_1310,N_1263,N_1246);
and U1311 (N_1311,N_1277,N_1207);
nand U1312 (N_1312,N_1201,N_1281);
nor U1313 (N_1313,N_1279,N_1225);
or U1314 (N_1314,N_1291,N_1271);
and U1315 (N_1315,N_1210,N_1240);
nor U1316 (N_1316,N_1262,N_1250);
nor U1317 (N_1317,N_1292,N_1212);
or U1318 (N_1318,N_1272,N_1252);
and U1319 (N_1319,N_1255,N_1253);
or U1320 (N_1320,N_1260,N_1290);
or U1321 (N_1321,N_1228,N_1222);
nor U1322 (N_1322,N_1268,N_1288);
nand U1323 (N_1323,N_1226,N_1229);
or U1324 (N_1324,N_1276,N_1242);
and U1325 (N_1325,N_1235,N_1204);
nor U1326 (N_1326,N_1256,N_1282);
or U1327 (N_1327,N_1298,N_1274);
and U1328 (N_1328,N_1245,N_1297);
and U1329 (N_1329,N_1259,N_1275);
or U1330 (N_1330,N_1205,N_1249);
and U1331 (N_1331,N_1299,N_1213);
and U1332 (N_1332,N_1265,N_1236);
nand U1333 (N_1333,N_1278,N_1219);
or U1334 (N_1334,N_1289,N_1247);
and U1335 (N_1335,N_1214,N_1209);
or U1336 (N_1336,N_1215,N_1295);
and U1337 (N_1337,N_1208,N_1285);
and U1338 (N_1338,N_1254,N_1217);
or U1339 (N_1339,N_1266,N_1220);
nor U1340 (N_1340,N_1211,N_1224);
nor U1341 (N_1341,N_1223,N_1287);
or U1342 (N_1342,N_1234,N_1293);
or U1343 (N_1343,N_1202,N_1283);
nor U1344 (N_1344,N_1203,N_1248);
and U1345 (N_1345,N_1294,N_1238);
nand U1346 (N_1346,N_1267,N_1216);
nand U1347 (N_1347,N_1221,N_1280);
or U1348 (N_1348,N_1232,N_1241);
nand U1349 (N_1349,N_1233,N_1231);
and U1350 (N_1350,N_1262,N_1293);
nor U1351 (N_1351,N_1294,N_1224);
and U1352 (N_1352,N_1218,N_1294);
and U1353 (N_1353,N_1213,N_1233);
nand U1354 (N_1354,N_1229,N_1277);
nand U1355 (N_1355,N_1270,N_1227);
and U1356 (N_1356,N_1294,N_1229);
and U1357 (N_1357,N_1282,N_1254);
or U1358 (N_1358,N_1276,N_1209);
xor U1359 (N_1359,N_1256,N_1257);
nand U1360 (N_1360,N_1297,N_1209);
and U1361 (N_1361,N_1292,N_1290);
nand U1362 (N_1362,N_1268,N_1245);
or U1363 (N_1363,N_1287,N_1264);
and U1364 (N_1364,N_1278,N_1282);
nand U1365 (N_1365,N_1215,N_1272);
nand U1366 (N_1366,N_1242,N_1278);
and U1367 (N_1367,N_1207,N_1280);
or U1368 (N_1368,N_1224,N_1276);
or U1369 (N_1369,N_1205,N_1277);
and U1370 (N_1370,N_1224,N_1263);
nor U1371 (N_1371,N_1253,N_1286);
nor U1372 (N_1372,N_1240,N_1257);
nor U1373 (N_1373,N_1295,N_1270);
xor U1374 (N_1374,N_1293,N_1202);
and U1375 (N_1375,N_1260,N_1240);
nand U1376 (N_1376,N_1208,N_1262);
and U1377 (N_1377,N_1206,N_1292);
or U1378 (N_1378,N_1209,N_1222);
and U1379 (N_1379,N_1264,N_1220);
and U1380 (N_1380,N_1211,N_1213);
and U1381 (N_1381,N_1259,N_1209);
nand U1382 (N_1382,N_1206,N_1226);
xnor U1383 (N_1383,N_1252,N_1203);
nor U1384 (N_1384,N_1282,N_1248);
or U1385 (N_1385,N_1276,N_1218);
nor U1386 (N_1386,N_1291,N_1273);
or U1387 (N_1387,N_1283,N_1221);
nor U1388 (N_1388,N_1252,N_1209);
nor U1389 (N_1389,N_1246,N_1254);
or U1390 (N_1390,N_1247,N_1256);
and U1391 (N_1391,N_1270,N_1250);
nor U1392 (N_1392,N_1272,N_1210);
nand U1393 (N_1393,N_1231,N_1284);
and U1394 (N_1394,N_1206,N_1229);
nand U1395 (N_1395,N_1249,N_1287);
nand U1396 (N_1396,N_1249,N_1248);
nor U1397 (N_1397,N_1291,N_1293);
nand U1398 (N_1398,N_1200,N_1274);
nor U1399 (N_1399,N_1222,N_1298);
nand U1400 (N_1400,N_1307,N_1339);
or U1401 (N_1401,N_1364,N_1313);
nor U1402 (N_1402,N_1361,N_1365);
nor U1403 (N_1403,N_1399,N_1320);
nor U1404 (N_1404,N_1350,N_1373);
nand U1405 (N_1405,N_1341,N_1380);
or U1406 (N_1406,N_1393,N_1377);
nand U1407 (N_1407,N_1379,N_1310);
nor U1408 (N_1408,N_1346,N_1368);
or U1409 (N_1409,N_1372,N_1333);
or U1410 (N_1410,N_1383,N_1314);
nand U1411 (N_1411,N_1354,N_1392);
nand U1412 (N_1412,N_1323,N_1389);
nor U1413 (N_1413,N_1303,N_1300);
and U1414 (N_1414,N_1319,N_1388);
or U1415 (N_1415,N_1366,N_1357);
nand U1416 (N_1416,N_1334,N_1316);
or U1417 (N_1417,N_1344,N_1376);
nor U1418 (N_1418,N_1340,N_1332);
xor U1419 (N_1419,N_1387,N_1351);
or U1420 (N_1420,N_1391,N_1335);
xor U1421 (N_1421,N_1358,N_1378);
nor U1422 (N_1422,N_1347,N_1304);
nand U1423 (N_1423,N_1337,N_1356);
nor U1424 (N_1424,N_1311,N_1374);
nand U1425 (N_1425,N_1327,N_1382);
and U1426 (N_1426,N_1315,N_1331);
or U1427 (N_1427,N_1355,N_1363);
or U1428 (N_1428,N_1395,N_1398);
and U1429 (N_1429,N_1348,N_1396);
and U1430 (N_1430,N_1336,N_1367);
nand U1431 (N_1431,N_1390,N_1309);
or U1432 (N_1432,N_1308,N_1328);
nand U1433 (N_1433,N_1352,N_1329);
nand U1434 (N_1434,N_1369,N_1338);
nand U1435 (N_1435,N_1349,N_1359);
and U1436 (N_1436,N_1325,N_1330);
or U1437 (N_1437,N_1397,N_1345);
and U1438 (N_1438,N_1302,N_1384);
nor U1439 (N_1439,N_1371,N_1306);
or U1440 (N_1440,N_1301,N_1362);
and U1441 (N_1441,N_1370,N_1318);
and U1442 (N_1442,N_1324,N_1305);
and U1443 (N_1443,N_1322,N_1326);
nand U1444 (N_1444,N_1342,N_1375);
or U1445 (N_1445,N_1360,N_1386);
nand U1446 (N_1446,N_1312,N_1321);
or U1447 (N_1447,N_1317,N_1385);
nor U1448 (N_1448,N_1381,N_1343);
or U1449 (N_1449,N_1353,N_1394);
and U1450 (N_1450,N_1307,N_1326);
nand U1451 (N_1451,N_1323,N_1363);
nand U1452 (N_1452,N_1386,N_1347);
and U1453 (N_1453,N_1396,N_1315);
and U1454 (N_1454,N_1317,N_1321);
or U1455 (N_1455,N_1377,N_1340);
nor U1456 (N_1456,N_1344,N_1361);
and U1457 (N_1457,N_1332,N_1310);
or U1458 (N_1458,N_1357,N_1359);
or U1459 (N_1459,N_1384,N_1315);
nand U1460 (N_1460,N_1350,N_1342);
nor U1461 (N_1461,N_1388,N_1395);
nor U1462 (N_1462,N_1396,N_1372);
nand U1463 (N_1463,N_1328,N_1389);
xor U1464 (N_1464,N_1316,N_1399);
nor U1465 (N_1465,N_1344,N_1323);
or U1466 (N_1466,N_1303,N_1330);
nor U1467 (N_1467,N_1363,N_1366);
nor U1468 (N_1468,N_1327,N_1368);
or U1469 (N_1469,N_1347,N_1354);
nor U1470 (N_1470,N_1348,N_1311);
and U1471 (N_1471,N_1356,N_1323);
nand U1472 (N_1472,N_1321,N_1392);
nand U1473 (N_1473,N_1313,N_1328);
and U1474 (N_1474,N_1331,N_1329);
or U1475 (N_1475,N_1326,N_1343);
and U1476 (N_1476,N_1363,N_1332);
nand U1477 (N_1477,N_1393,N_1346);
nor U1478 (N_1478,N_1392,N_1381);
or U1479 (N_1479,N_1360,N_1329);
or U1480 (N_1480,N_1323,N_1377);
or U1481 (N_1481,N_1321,N_1391);
and U1482 (N_1482,N_1367,N_1355);
or U1483 (N_1483,N_1372,N_1300);
or U1484 (N_1484,N_1326,N_1352);
or U1485 (N_1485,N_1327,N_1339);
or U1486 (N_1486,N_1350,N_1361);
nor U1487 (N_1487,N_1332,N_1319);
and U1488 (N_1488,N_1392,N_1325);
nor U1489 (N_1489,N_1359,N_1333);
nand U1490 (N_1490,N_1311,N_1370);
nor U1491 (N_1491,N_1322,N_1369);
or U1492 (N_1492,N_1369,N_1312);
or U1493 (N_1493,N_1358,N_1391);
and U1494 (N_1494,N_1346,N_1314);
and U1495 (N_1495,N_1367,N_1354);
nand U1496 (N_1496,N_1387,N_1393);
nand U1497 (N_1497,N_1353,N_1319);
or U1498 (N_1498,N_1388,N_1314);
and U1499 (N_1499,N_1309,N_1330);
nor U1500 (N_1500,N_1475,N_1482);
or U1501 (N_1501,N_1462,N_1464);
nor U1502 (N_1502,N_1460,N_1467);
and U1503 (N_1503,N_1418,N_1401);
or U1504 (N_1504,N_1451,N_1453);
and U1505 (N_1505,N_1438,N_1425);
or U1506 (N_1506,N_1457,N_1428);
nor U1507 (N_1507,N_1446,N_1483);
or U1508 (N_1508,N_1441,N_1443);
nor U1509 (N_1509,N_1494,N_1432);
and U1510 (N_1510,N_1478,N_1450);
and U1511 (N_1511,N_1471,N_1442);
nand U1512 (N_1512,N_1436,N_1426);
and U1513 (N_1513,N_1496,N_1461);
and U1514 (N_1514,N_1434,N_1412);
nand U1515 (N_1515,N_1417,N_1497);
or U1516 (N_1516,N_1458,N_1491);
nand U1517 (N_1517,N_1484,N_1440);
or U1518 (N_1518,N_1449,N_1437);
or U1519 (N_1519,N_1452,N_1470);
and U1520 (N_1520,N_1403,N_1445);
and U1521 (N_1521,N_1455,N_1486);
nand U1522 (N_1522,N_1448,N_1459);
or U1523 (N_1523,N_1489,N_1492);
and U1524 (N_1524,N_1466,N_1490);
or U1525 (N_1525,N_1479,N_1414);
nor U1526 (N_1526,N_1487,N_1410);
nor U1527 (N_1527,N_1402,N_1473);
nand U1528 (N_1528,N_1439,N_1488);
or U1529 (N_1529,N_1495,N_1411);
or U1530 (N_1530,N_1400,N_1454);
nor U1531 (N_1531,N_1415,N_1477);
or U1532 (N_1532,N_1465,N_1406);
and U1533 (N_1533,N_1416,N_1420);
and U1534 (N_1534,N_1424,N_1493);
or U1535 (N_1535,N_1480,N_1481);
nand U1536 (N_1536,N_1456,N_1447);
nor U1537 (N_1537,N_1498,N_1430);
or U1538 (N_1538,N_1405,N_1472);
and U1539 (N_1539,N_1469,N_1422);
nand U1540 (N_1540,N_1433,N_1408);
nand U1541 (N_1541,N_1409,N_1419);
nand U1542 (N_1542,N_1499,N_1474);
and U1543 (N_1543,N_1468,N_1444);
and U1544 (N_1544,N_1485,N_1423);
or U1545 (N_1545,N_1429,N_1407);
or U1546 (N_1546,N_1421,N_1427);
nand U1547 (N_1547,N_1463,N_1476);
nor U1548 (N_1548,N_1431,N_1404);
nor U1549 (N_1549,N_1413,N_1435);
or U1550 (N_1550,N_1491,N_1475);
nand U1551 (N_1551,N_1450,N_1435);
nand U1552 (N_1552,N_1464,N_1417);
and U1553 (N_1553,N_1472,N_1487);
or U1554 (N_1554,N_1442,N_1437);
and U1555 (N_1555,N_1453,N_1418);
nand U1556 (N_1556,N_1412,N_1400);
nor U1557 (N_1557,N_1483,N_1447);
nand U1558 (N_1558,N_1403,N_1484);
nand U1559 (N_1559,N_1467,N_1472);
nand U1560 (N_1560,N_1455,N_1492);
nor U1561 (N_1561,N_1474,N_1400);
nor U1562 (N_1562,N_1427,N_1475);
and U1563 (N_1563,N_1424,N_1467);
and U1564 (N_1564,N_1484,N_1480);
and U1565 (N_1565,N_1400,N_1424);
and U1566 (N_1566,N_1488,N_1473);
nand U1567 (N_1567,N_1495,N_1478);
nand U1568 (N_1568,N_1479,N_1421);
nor U1569 (N_1569,N_1447,N_1485);
nand U1570 (N_1570,N_1467,N_1446);
or U1571 (N_1571,N_1413,N_1405);
or U1572 (N_1572,N_1416,N_1425);
nor U1573 (N_1573,N_1435,N_1462);
nand U1574 (N_1574,N_1409,N_1491);
or U1575 (N_1575,N_1420,N_1407);
and U1576 (N_1576,N_1413,N_1408);
nand U1577 (N_1577,N_1446,N_1499);
nand U1578 (N_1578,N_1441,N_1482);
nand U1579 (N_1579,N_1418,N_1464);
and U1580 (N_1580,N_1471,N_1448);
nor U1581 (N_1581,N_1442,N_1425);
or U1582 (N_1582,N_1440,N_1478);
xnor U1583 (N_1583,N_1459,N_1402);
and U1584 (N_1584,N_1415,N_1438);
nand U1585 (N_1585,N_1451,N_1403);
nand U1586 (N_1586,N_1464,N_1495);
nor U1587 (N_1587,N_1499,N_1415);
or U1588 (N_1588,N_1465,N_1467);
nand U1589 (N_1589,N_1474,N_1498);
xor U1590 (N_1590,N_1450,N_1485);
nand U1591 (N_1591,N_1488,N_1495);
or U1592 (N_1592,N_1402,N_1422);
or U1593 (N_1593,N_1427,N_1403);
nand U1594 (N_1594,N_1498,N_1465);
nand U1595 (N_1595,N_1457,N_1496);
nor U1596 (N_1596,N_1418,N_1454);
and U1597 (N_1597,N_1482,N_1403);
or U1598 (N_1598,N_1496,N_1479);
or U1599 (N_1599,N_1473,N_1432);
and U1600 (N_1600,N_1503,N_1523);
nor U1601 (N_1601,N_1539,N_1567);
xor U1602 (N_1602,N_1542,N_1596);
nor U1603 (N_1603,N_1590,N_1525);
nor U1604 (N_1604,N_1589,N_1517);
nor U1605 (N_1605,N_1592,N_1521);
nor U1606 (N_1606,N_1530,N_1549);
or U1607 (N_1607,N_1564,N_1540);
and U1608 (N_1608,N_1512,N_1568);
xor U1609 (N_1609,N_1509,N_1534);
nor U1610 (N_1610,N_1504,N_1576);
nor U1611 (N_1611,N_1599,N_1529);
nand U1612 (N_1612,N_1572,N_1513);
nor U1613 (N_1613,N_1581,N_1566);
and U1614 (N_1614,N_1526,N_1583);
and U1615 (N_1615,N_1577,N_1559);
and U1616 (N_1616,N_1531,N_1561);
nand U1617 (N_1617,N_1501,N_1519);
and U1618 (N_1618,N_1546,N_1598);
nand U1619 (N_1619,N_1533,N_1544);
or U1620 (N_1620,N_1570,N_1569);
nand U1621 (N_1621,N_1545,N_1541);
or U1622 (N_1622,N_1594,N_1505);
and U1623 (N_1623,N_1516,N_1555);
and U1624 (N_1624,N_1588,N_1571);
or U1625 (N_1625,N_1597,N_1547);
nor U1626 (N_1626,N_1508,N_1586);
nor U1627 (N_1627,N_1557,N_1595);
nand U1628 (N_1628,N_1579,N_1573);
nor U1629 (N_1629,N_1585,N_1538);
xnor U1630 (N_1630,N_1527,N_1500);
nor U1631 (N_1631,N_1580,N_1565);
nand U1632 (N_1632,N_1528,N_1591);
or U1633 (N_1633,N_1510,N_1562);
or U1634 (N_1634,N_1522,N_1537);
or U1635 (N_1635,N_1554,N_1553);
or U1636 (N_1636,N_1578,N_1593);
or U1637 (N_1637,N_1560,N_1575);
or U1638 (N_1638,N_1536,N_1524);
nand U1639 (N_1639,N_1520,N_1582);
nand U1640 (N_1640,N_1506,N_1518);
nand U1641 (N_1641,N_1502,N_1552);
and U1642 (N_1642,N_1543,N_1507);
nand U1643 (N_1643,N_1515,N_1587);
and U1644 (N_1644,N_1532,N_1551);
and U1645 (N_1645,N_1563,N_1511);
nor U1646 (N_1646,N_1558,N_1574);
or U1647 (N_1647,N_1550,N_1584);
and U1648 (N_1648,N_1514,N_1556);
and U1649 (N_1649,N_1548,N_1535);
and U1650 (N_1650,N_1528,N_1522);
or U1651 (N_1651,N_1593,N_1503);
or U1652 (N_1652,N_1501,N_1585);
nor U1653 (N_1653,N_1594,N_1537);
and U1654 (N_1654,N_1582,N_1598);
nand U1655 (N_1655,N_1501,N_1540);
nor U1656 (N_1656,N_1547,N_1546);
or U1657 (N_1657,N_1597,N_1578);
nor U1658 (N_1658,N_1515,N_1510);
nor U1659 (N_1659,N_1521,N_1572);
nand U1660 (N_1660,N_1591,N_1526);
nand U1661 (N_1661,N_1511,N_1578);
or U1662 (N_1662,N_1575,N_1543);
nand U1663 (N_1663,N_1509,N_1555);
nor U1664 (N_1664,N_1550,N_1578);
nor U1665 (N_1665,N_1522,N_1525);
and U1666 (N_1666,N_1513,N_1544);
nor U1667 (N_1667,N_1564,N_1568);
nor U1668 (N_1668,N_1518,N_1591);
and U1669 (N_1669,N_1579,N_1545);
or U1670 (N_1670,N_1550,N_1529);
and U1671 (N_1671,N_1526,N_1578);
nor U1672 (N_1672,N_1573,N_1596);
xor U1673 (N_1673,N_1513,N_1501);
nand U1674 (N_1674,N_1567,N_1503);
nor U1675 (N_1675,N_1551,N_1518);
nand U1676 (N_1676,N_1536,N_1521);
nand U1677 (N_1677,N_1552,N_1571);
or U1678 (N_1678,N_1503,N_1543);
or U1679 (N_1679,N_1539,N_1535);
and U1680 (N_1680,N_1587,N_1598);
or U1681 (N_1681,N_1541,N_1550);
nor U1682 (N_1682,N_1564,N_1504);
and U1683 (N_1683,N_1515,N_1585);
or U1684 (N_1684,N_1585,N_1539);
xnor U1685 (N_1685,N_1519,N_1583);
and U1686 (N_1686,N_1570,N_1595);
xnor U1687 (N_1687,N_1547,N_1551);
nand U1688 (N_1688,N_1519,N_1556);
nor U1689 (N_1689,N_1584,N_1572);
nand U1690 (N_1690,N_1524,N_1551);
nand U1691 (N_1691,N_1527,N_1542);
nand U1692 (N_1692,N_1515,N_1573);
nor U1693 (N_1693,N_1520,N_1505);
or U1694 (N_1694,N_1504,N_1537);
xor U1695 (N_1695,N_1519,N_1568);
nor U1696 (N_1696,N_1558,N_1519);
or U1697 (N_1697,N_1593,N_1544);
or U1698 (N_1698,N_1542,N_1590);
nor U1699 (N_1699,N_1536,N_1571);
nor U1700 (N_1700,N_1631,N_1676);
nand U1701 (N_1701,N_1681,N_1665);
nand U1702 (N_1702,N_1630,N_1680);
nand U1703 (N_1703,N_1610,N_1651);
nand U1704 (N_1704,N_1641,N_1618);
or U1705 (N_1705,N_1657,N_1656);
nor U1706 (N_1706,N_1604,N_1647);
xor U1707 (N_1707,N_1626,N_1697);
nor U1708 (N_1708,N_1632,N_1691);
or U1709 (N_1709,N_1690,N_1617);
and U1710 (N_1710,N_1698,N_1619);
nor U1711 (N_1711,N_1685,N_1668);
nand U1712 (N_1712,N_1674,N_1622);
nand U1713 (N_1713,N_1611,N_1609);
xor U1714 (N_1714,N_1603,N_1634);
nor U1715 (N_1715,N_1678,N_1649);
nand U1716 (N_1716,N_1629,N_1662);
xor U1717 (N_1717,N_1650,N_1688);
nor U1718 (N_1718,N_1648,N_1637);
or U1719 (N_1719,N_1639,N_1664);
xnor U1720 (N_1720,N_1640,N_1695);
nor U1721 (N_1721,N_1633,N_1661);
nor U1722 (N_1722,N_1699,N_1621);
or U1723 (N_1723,N_1686,N_1660);
nor U1724 (N_1724,N_1644,N_1623);
and U1725 (N_1725,N_1667,N_1605);
nand U1726 (N_1726,N_1670,N_1620);
nand U1727 (N_1727,N_1666,N_1694);
nand U1728 (N_1728,N_1607,N_1692);
nand U1729 (N_1729,N_1624,N_1642);
nor U1730 (N_1730,N_1677,N_1615);
nand U1731 (N_1731,N_1672,N_1693);
nand U1732 (N_1732,N_1646,N_1652);
or U1733 (N_1733,N_1663,N_1612);
nor U1734 (N_1734,N_1608,N_1671);
or U1735 (N_1735,N_1689,N_1601);
and U1736 (N_1736,N_1613,N_1654);
or U1737 (N_1737,N_1655,N_1658);
nand U1738 (N_1738,N_1627,N_1684);
or U1739 (N_1739,N_1600,N_1683);
nor U1740 (N_1740,N_1653,N_1643);
or U1741 (N_1741,N_1696,N_1659);
nand U1742 (N_1742,N_1673,N_1682);
and U1743 (N_1743,N_1635,N_1628);
nor U1744 (N_1744,N_1675,N_1614);
and U1745 (N_1745,N_1602,N_1625);
nor U1746 (N_1746,N_1669,N_1606);
nand U1747 (N_1747,N_1638,N_1687);
nand U1748 (N_1748,N_1636,N_1645);
and U1749 (N_1749,N_1616,N_1679);
and U1750 (N_1750,N_1671,N_1666);
nor U1751 (N_1751,N_1608,N_1685);
or U1752 (N_1752,N_1673,N_1695);
nor U1753 (N_1753,N_1622,N_1685);
or U1754 (N_1754,N_1673,N_1693);
nand U1755 (N_1755,N_1699,N_1679);
nor U1756 (N_1756,N_1641,N_1651);
or U1757 (N_1757,N_1685,N_1698);
nor U1758 (N_1758,N_1655,N_1678);
nand U1759 (N_1759,N_1612,N_1652);
and U1760 (N_1760,N_1652,N_1601);
nor U1761 (N_1761,N_1660,N_1611);
or U1762 (N_1762,N_1656,N_1643);
nand U1763 (N_1763,N_1613,N_1647);
and U1764 (N_1764,N_1671,N_1618);
and U1765 (N_1765,N_1662,N_1682);
nand U1766 (N_1766,N_1633,N_1622);
or U1767 (N_1767,N_1696,N_1688);
nor U1768 (N_1768,N_1675,N_1687);
or U1769 (N_1769,N_1620,N_1635);
and U1770 (N_1770,N_1643,N_1636);
nor U1771 (N_1771,N_1651,N_1693);
nor U1772 (N_1772,N_1673,N_1601);
and U1773 (N_1773,N_1649,N_1621);
or U1774 (N_1774,N_1653,N_1659);
nor U1775 (N_1775,N_1634,N_1620);
nor U1776 (N_1776,N_1672,N_1668);
or U1777 (N_1777,N_1682,N_1644);
or U1778 (N_1778,N_1615,N_1624);
and U1779 (N_1779,N_1698,N_1607);
and U1780 (N_1780,N_1678,N_1666);
and U1781 (N_1781,N_1645,N_1651);
nor U1782 (N_1782,N_1681,N_1615);
nand U1783 (N_1783,N_1617,N_1658);
or U1784 (N_1784,N_1678,N_1646);
or U1785 (N_1785,N_1653,N_1646);
or U1786 (N_1786,N_1630,N_1603);
nand U1787 (N_1787,N_1684,N_1613);
nand U1788 (N_1788,N_1672,N_1628);
or U1789 (N_1789,N_1611,N_1695);
or U1790 (N_1790,N_1627,N_1634);
or U1791 (N_1791,N_1662,N_1675);
nor U1792 (N_1792,N_1657,N_1678);
and U1793 (N_1793,N_1656,N_1644);
nor U1794 (N_1794,N_1663,N_1670);
nor U1795 (N_1795,N_1687,N_1612);
xnor U1796 (N_1796,N_1655,N_1614);
or U1797 (N_1797,N_1688,N_1606);
and U1798 (N_1798,N_1686,N_1695);
nor U1799 (N_1799,N_1685,N_1602);
nand U1800 (N_1800,N_1738,N_1722);
nand U1801 (N_1801,N_1744,N_1725);
or U1802 (N_1802,N_1792,N_1740);
and U1803 (N_1803,N_1774,N_1754);
or U1804 (N_1804,N_1776,N_1746);
nand U1805 (N_1805,N_1712,N_1717);
and U1806 (N_1806,N_1750,N_1724);
or U1807 (N_1807,N_1769,N_1735);
nand U1808 (N_1808,N_1796,N_1704);
and U1809 (N_1809,N_1785,N_1702);
nor U1810 (N_1810,N_1730,N_1718);
and U1811 (N_1811,N_1710,N_1731);
nand U1812 (N_1812,N_1760,N_1777);
and U1813 (N_1813,N_1737,N_1732);
xnor U1814 (N_1814,N_1736,N_1773);
and U1815 (N_1815,N_1742,N_1770);
nand U1816 (N_1816,N_1759,N_1720);
nor U1817 (N_1817,N_1709,N_1705);
nand U1818 (N_1818,N_1766,N_1745);
nor U1819 (N_1819,N_1701,N_1786);
nand U1820 (N_1820,N_1767,N_1751);
nand U1821 (N_1821,N_1711,N_1723);
nor U1822 (N_1822,N_1761,N_1753);
or U1823 (N_1823,N_1780,N_1763);
or U1824 (N_1824,N_1791,N_1755);
nor U1825 (N_1825,N_1716,N_1790);
nand U1826 (N_1826,N_1797,N_1721);
nand U1827 (N_1827,N_1788,N_1756);
and U1828 (N_1828,N_1719,N_1739);
nand U1829 (N_1829,N_1799,N_1743);
or U1830 (N_1830,N_1748,N_1728);
nand U1831 (N_1831,N_1714,N_1726);
nand U1832 (N_1832,N_1789,N_1729);
or U1833 (N_1833,N_1768,N_1783);
nand U1834 (N_1834,N_1794,N_1762);
nor U1835 (N_1835,N_1706,N_1781);
nand U1836 (N_1836,N_1703,N_1795);
and U1837 (N_1837,N_1787,N_1708);
and U1838 (N_1838,N_1741,N_1757);
and U1839 (N_1839,N_1715,N_1764);
nand U1840 (N_1840,N_1793,N_1772);
nand U1841 (N_1841,N_1778,N_1784);
or U1842 (N_1842,N_1758,N_1765);
nand U1843 (N_1843,N_1775,N_1707);
nor U1844 (N_1844,N_1734,N_1747);
nor U1845 (N_1845,N_1779,N_1713);
nor U1846 (N_1846,N_1752,N_1782);
and U1847 (N_1847,N_1727,N_1733);
nand U1848 (N_1848,N_1700,N_1798);
and U1849 (N_1849,N_1771,N_1749);
and U1850 (N_1850,N_1764,N_1790);
and U1851 (N_1851,N_1725,N_1763);
nand U1852 (N_1852,N_1739,N_1753);
nand U1853 (N_1853,N_1792,N_1723);
and U1854 (N_1854,N_1774,N_1712);
nor U1855 (N_1855,N_1772,N_1758);
and U1856 (N_1856,N_1741,N_1745);
or U1857 (N_1857,N_1744,N_1788);
or U1858 (N_1858,N_1737,N_1781);
and U1859 (N_1859,N_1739,N_1731);
nor U1860 (N_1860,N_1796,N_1726);
nand U1861 (N_1861,N_1771,N_1718);
nand U1862 (N_1862,N_1737,N_1766);
nand U1863 (N_1863,N_1709,N_1739);
nor U1864 (N_1864,N_1783,N_1717);
xor U1865 (N_1865,N_1767,N_1766);
or U1866 (N_1866,N_1734,N_1791);
or U1867 (N_1867,N_1749,N_1700);
or U1868 (N_1868,N_1730,N_1765);
nor U1869 (N_1869,N_1747,N_1760);
nand U1870 (N_1870,N_1797,N_1798);
or U1871 (N_1871,N_1738,N_1740);
nand U1872 (N_1872,N_1761,N_1776);
nor U1873 (N_1873,N_1751,N_1745);
or U1874 (N_1874,N_1742,N_1798);
and U1875 (N_1875,N_1737,N_1753);
nor U1876 (N_1876,N_1788,N_1718);
or U1877 (N_1877,N_1756,N_1732);
or U1878 (N_1878,N_1730,N_1781);
xnor U1879 (N_1879,N_1761,N_1715);
and U1880 (N_1880,N_1715,N_1719);
or U1881 (N_1881,N_1711,N_1728);
nand U1882 (N_1882,N_1764,N_1745);
and U1883 (N_1883,N_1725,N_1732);
nand U1884 (N_1884,N_1750,N_1718);
nand U1885 (N_1885,N_1782,N_1703);
or U1886 (N_1886,N_1711,N_1765);
nand U1887 (N_1887,N_1770,N_1703);
xnor U1888 (N_1888,N_1724,N_1700);
or U1889 (N_1889,N_1772,N_1712);
and U1890 (N_1890,N_1799,N_1705);
nand U1891 (N_1891,N_1783,N_1752);
nor U1892 (N_1892,N_1770,N_1733);
or U1893 (N_1893,N_1750,N_1737);
nor U1894 (N_1894,N_1752,N_1777);
xnor U1895 (N_1895,N_1784,N_1711);
or U1896 (N_1896,N_1796,N_1744);
or U1897 (N_1897,N_1799,N_1781);
nor U1898 (N_1898,N_1701,N_1704);
and U1899 (N_1899,N_1779,N_1794);
nand U1900 (N_1900,N_1812,N_1887);
nor U1901 (N_1901,N_1855,N_1876);
and U1902 (N_1902,N_1872,N_1871);
or U1903 (N_1903,N_1821,N_1844);
and U1904 (N_1904,N_1899,N_1827);
and U1905 (N_1905,N_1819,N_1836);
nand U1906 (N_1906,N_1817,N_1840);
nand U1907 (N_1907,N_1848,N_1842);
nor U1908 (N_1908,N_1815,N_1891);
nor U1909 (N_1909,N_1835,N_1801);
and U1910 (N_1910,N_1864,N_1890);
nor U1911 (N_1911,N_1893,N_1838);
or U1912 (N_1912,N_1843,N_1868);
and U1913 (N_1913,N_1892,N_1863);
nand U1914 (N_1914,N_1880,N_1830);
nor U1915 (N_1915,N_1878,N_1857);
nor U1916 (N_1916,N_1841,N_1802);
nand U1917 (N_1917,N_1822,N_1896);
and U1918 (N_1918,N_1833,N_1845);
nand U1919 (N_1919,N_1865,N_1824);
nand U1920 (N_1920,N_1806,N_1853);
xor U1921 (N_1921,N_1885,N_1861);
nand U1922 (N_1922,N_1866,N_1803);
or U1923 (N_1923,N_1847,N_1839);
and U1924 (N_1924,N_1886,N_1807);
nand U1925 (N_1925,N_1882,N_1895);
or U1926 (N_1926,N_1877,N_1849);
or U1927 (N_1927,N_1862,N_1820);
or U1928 (N_1928,N_1825,N_1883);
and U1929 (N_1929,N_1859,N_1816);
and U1930 (N_1930,N_1851,N_1884);
or U1931 (N_1931,N_1858,N_1846);
or U1932 (N_1932,N_1879,N_1852);
nor U1933 (N_1933,N_1814,N_1828);
xnor U1934 (N_1934,N_1829,N_1888);
nand U1935 (N_1935,N_1813,N_1897);
nand U1936 (N_1936,N_1837,N_1850);
nand U1937 (N_1937,N_1811,N_1874);
or U1938 (N_1938,N_1894,N_1867);
nor U1939 (N_1939,N_1869,N_1834);
nor U1940 (N_1940,N_1826,N_1808);
nand U1941 (N_1941,N_1804,N_1831);
and U1942 (N_1942,N_1860,N_1889);
or U1943 (N_1943,N_1805,N_1823);
or U1944 (N_1944,N_1809,N_1854);
nor U1945 (N_1945,N_1875,N_1800);
and U1946 (N_1946,N_1810,N_1818);
or U1947 (N_1947,N_1832,N_1881);
nor U1948 (N_1948,N_1873,N_1898);
nor U1949 (N_1949,N_1870,N_1856);
nand U1950 (N_1950,N_1826,N_1884);
nor U1951 (N_1951,N_1841,N_1811);
nor U1952 (N_1952,N_1896,N_1844);
and U1953 (N_1953,N_1897,N_1859);
or U1954 (N_1954,N_1848,N_1839);
nor U1955 (N_1955,N_1832,N_1823);
nand U1956 (N_1956,N_1895,N_1859);
or U1957 (N_1957,N_1858,N_1813);
nor U1958 (N_1958,N_1874,N_1838);
or U1959 (N_1959,N_1825,N_1882);
nand U1960 (N_1960,N_1899,N_1873);
or U1961 (N_1961,N_1836,N_1805);
nor U1962 (N_1962,N_1875,N_1823);
or U1963 (N_1963,N_1849,N_1863);
and U1964 (N_1964,N_1805,N_1897);
and U1965 (N_1965,N_1808,N_1859);
and U1966 (N_1966,N_1829,N_1819);
nand U1967 (N_1967,N_1846,N_1832);
nor U1968 (N_1968,N_1866,N_1808);
nor U1969 (N_1969,N_1812,N_1837);
and U1970 (N_1970,N_1838,N_1883);
and U1971 (N_1971,N_1878,N_1867);
and U1972 (N_1972,N_1881,N_1887);
nor U1973 (N_1973,N_1814,N_1893);
nor U1974 (N_1974,N_1862,N_1848);
and U1975 (N_1975,N_1895,N_1832);
nand U1976 (N_1976,N_1860,N_1812);
or U1977 (N_1977,N_1881,N_1826);
and U1978 (N_1978,N_1889,N_1814);
or U1979 (N_1979,N_1892,N_1896);
nand U1980 (N_1980,N_1835,N_1873);
or U1981 (N_1981,N_1868,N_1801);
and U1982 (N_1982,N_1872,N_1819);
or U1983 (N_1983,N_1863,N_1818);
and U1984 (N_1984,N_1801,N_1816);
nor U1985 (N_1985,N_1844,N_1845);
or U1986 (N_1986,N_1833,N_1890);
nor U1987 (N_1987,N_1891,N_1837);
and U1988 (N_1988,N_1870,N_1895);
nand U1989 (N_1989,N_1833,N_1851);
nor U1990 (N_1990,N_1801,N_1895);
xnor U1991 (N_1991,N_1896,N_1861);
or U1992 (N_1992,N_1857,N_1887);
nand U1993 (N_1993,N_1856,N_1844);
and U1994 (N_1994,N_1896,N_1863);
or U1995 (N_1995,N_1836,N_1850);
and U1996 (N_1996,N_1877,N_1895);
or U1997 (N_1997,N_1854,N_1869);
nand U1998 (N_1998,N_1864,N_1837);
or U1999 (N_1999,N_1819,N_1894);
nor U2000 (N_2000,N_1941,N_1960);
and U2001 (N_2001,N_1920,N_1999);
or U2002 (N_2002,N_1957,N_1973);
nand U2003 (N_2003,N_1932,N_1967);
nand U2004 (N_2004,N_1910,N_1905);
and U2005 (N_2005,N_1947,N_1938);
and U2006 (N_2006,N_1976,N_1968);
or U2007 (N_2007,N_1948,N_1979);
nor U2008 (N_2008,N_1923,N_1916);
nor U2009 (N_2009,N_1959,N_1915);
nor U2010 (N_2010,N_1961,N_1945);
or U2011 (N_2011,N_1940,N_1975);
and U2012 (N_2012,N_1949,N_1982);
nand U2013 (N_2013,N_1919,N_1954);
or U2014 (N_2014,N_1935,N_1912);
and U2015 (N_2015,N_1930,N_1917);
or U2016 (N_2016,N_1989,N_1969);
or U2017 (N_2017,N_1997,N_1925);
nor U2018 (N_2018,N_1987,N_1983);
nand U2019 (N_2019,N_1900,N_1981);
and U2020 (N_2020,N_1922,N_1931);
and U2021 (N_2021,N_1974,N_1965);
nand U2022 (N_2022,N_1956,N_1901);
nand U2023 (N_2023,N_1986,N_1977);
or U2024 (N_2024,N_1903,N_1924);
or U2025 (N_2025,N_1946,N_1936);
nor U2026 (N_2026,N_1902,N_1921);
and U2027 (N_2027,N_1958,N_1966);
and U2028 (N_2028,N_1951,N_1985);
and U2029 (N_2029,N_1927,N_1963);
and U2030 (N_2030,N_1971,N_1918);
or U2031 (N_2031,N_1970,N_1988);
nor U2032 (N_2032,N_1995,N_1913);
nor U2033 (N_2033,N_1937,N_1906);
and U2034 (N_2034,N_1907,N_1984);
nand U2035 (N_2035,N_1952,N_1994);
nor U2036 (N_2036,N_1962,N_1914);
and U2037 (N_2037,N_1904,N_1908);
xnor U2038 (N_2038,N_1942,N_1990);
or U2039 (N_2039,N_1953,N_1911);
nor U2040 (N_2040,N_1929,N_1978);
nand U2041 (N_2041,N_1950,N_1998);
and U2042 (N_2042,N_1928,N_1991);
xor U2043 (N_2043,N_1909,N_1934);
or U2044 (N_2044,N_1992,N_1964);
and U2045 (N_2045,N_1993,N_1926);
nand U2046 (N_2046,N_1939,N_1933);
and U2047 (N_2047,N_1980,N_1955);
nand U2048 (N_2048,N_1972,N_1996);
or U2049 (N_2049,N_1944,N_1943);
or U2050 (N_2050,N_1927,N_1984);
or U2051 (N_2051,N_1928,N_1960);
or U2052 (N_2052,N_1985,N_1964);
and U2053 (N_2053,N_1914,N_1957);
nor U2054 (N_2054,N_1901,N_1900);
nor U2055 (N_2055,N_1933,N_1923);
and U2056 (N_2056,N_1916,N_1915);
or U2057 (N_2057,N_1941,N_1982);
nor U2058 (N_2058,N_1940,N_1951);
nand U2059 (N_2059,N_1951,N_1924);
and U2060 (N_2060,N_1907,N_1937);
nand U2061 (N_2061,N_1979,N_1953);
or U2062 (N_2062,N_1975,N_1970);
or U2063 (N_2063,N_1943,N_1954);
and U2064 (N_2064,N_1934,N_1995);
nand U2065 (N_2065,N_1928,N_1957);
nor U2066 (N_2066,N_1909,N_1929);
nor U2067 (N_2067,N_1984,N_1915);
nand U2068 (N_2068,N_1920,N_1964);
nor U2069 (N_2069,N_1900,N_1998);
or U2070 (N_2070,N_1930,N_1997);
nor U2071 (N_2071,N_1993,N_1961);
nor U2072 (N_2072,N_1930,N_1969);
nand U2073 (N_2073,N_1950,N_1972);
nor U2074 (N_2074,N_1961,N_1982);
and U2075 (N_2075,N_1985,N_1935);
nor U2076 (N_2076,N_1945,N_1976);
nand U2077 (N_2077,N_1935,N_1967);
nor U2078 (N_2078,N_1901,N_1985);
or U2079 (N_2079,N_1924,N_1972);
nand U2080 (N_2080,N_1935,N_1913);
nor U2081 (N_2081,N_1972,N_1970);
nor U2082 (N_2082,N_1962,N_1937);
or U2083 (N_2083,N_1963,N_1904);
or U2084 (N_2084,N_1965,N_1975);
xor U2085 (N_2085,N_1955,N_1922);
nand U2086 (N_2086,N_1903,N_1927);
or U2087 (N_2087,N_1904,N_1927);
or U2088 (N_2088,N_1966,N_1975);
nand U2089 (N_2089,N_1968,N_1959);
xnor U2090 (N_2090,N_1908,N_1929);
and U2091 (N_2091,N_1972,N_1959);
nor U2092 (N_2092,N_1932,N_1915);
nor U2093 (N_2093,N_1978,N_1925);
or U2094 (N_2094,N_1965,N_1916);
or U2095 (N_2095,N_1926,N_1929);
and U2096 (N_2096,N_1923,N_1960);
nand U2097 (N_2097,N_1996,N_1984);
nand U2098 (N_2098,N_1924,N_1976);
or U2099 (N_2099,N_1929,N_1914);
or U2100 (N_2100,N_2055,N_2060);
or U2101 (N_2101,N_2038,N_2042);
or U2102 (N_2102,N_2002,N_2090);
and U2103 (N_2103,N_2019,N_2046);
nand U2104 (N_2104,N_2040,N_2009);
nand U2105 (N_2105,N_2097,N_2013);
or U2106 (N_2106,N_2054,N_2065);
nor U2107 (N_2107,N_2053,N_2078);
nand U2108 (N_2108,N_2056,N_2092);
and U2109 (N_2109,N_2045,N_2057);
nor U2110 (N_2110,N_2099,N_2016);
nor U2111 (N_2111,N_2072,N_2073);
nor U2112 (N_2112,N_2018,N_2077);
xnor U2113 (N_2113,N_2027,N_2021);
or U2114 (N_2114,N_2029,N_2037);
and U2115 (N_2115,N_2047,N_2082);
xor U2116 (N_2116,N_2030,N_2003);
nand U2117 (N_2117,N_2012,N_2049);
and U2118 (N_2118,N_2050,N_2080);
nand U2119 (N_2119,N_2096,N_2091);
nand U2120 (N_2120,N_2067,N_2095);
or U2121 (N_2121,N_2031,N_2089);
and U2122 (N_2122,N_2087,N_2081);
xor U2123 (N_2123,N_2017,N_2064);
and U2124 (N_2124,N_2084,N_2076);
or U2125 (N_2125,N_2032,N_2074);
or U2126 (N_2126,N_2005,N_2034);
nor U2127 (N_2127,N_2094,N_2025);
and U2128 (N_2128,N_2052,N_2071);
and U2129 (N_2129,N_2098,N_2028);
and U2130 (N_2130,N_2011,N_2085);
nand U2131 (N_2131,N_2039,N_2014);
nand U2132 (N_2132,N_2083,N_2059);
or U2133 (N_2133,N_2024,N_2066);
or U2134 (N_2134,N_2020,N_2075);
nand U2135 (N_2135,N_2007,N_2023);
and U2136 (N_2136,N_2086,N_2068);
nand U2137 (N_2137,N_2001,N_2048);
or U2138 (N_2138,N_2070,N_2000);
and U2139 (N_2139,N_2069,N_2033);
or U2140 (N_2140,N_2062,N_2010);
and U2141 (N_2141,N_2015,N_2022);
and U2142 (N_2142,N_2026,N_2004);
nand U2143 (N_2143,N_2044,N_2035);
nor U2144 (N_2144,N_2051,N_2093);
nand U2145 (N_2145,N_2088,N_2079);
nor U2146 (N_2146,N_2036,N_2008);
or U2147 (N_2147,N_2061,N_2058);
and U2148 (N_2148,N_2063,N_2043);
nand U2149 (N_2149,N_2006,N_2041);
nand U2150 (N_2150,N_2012,N_2051);
nand U2151 (N_2151,N_2033,N_2008);
and U2152 (N_2152,N_2045,N_2096);
nor U2153 (N_2153,N_2082,N_2071);
or U2154 (N_2154,N_2008,N_2045);
and U2155 (N_2155,N_2048,N_2052);
nand U2156 (N_2156,N_2078,N_2069);
nor U2157 (N_2157,N_2098,N_2030);
nand U2158 (N_2158,N_2000,N_2060);
and U2159 (N_2159,N_2004,N_2098);
or U2160 (N_2160,N_2062,N_2067);
and U2161 (N_2161,N_2027,N_2042);
nor U2162 (N_2162,N_2032,N_2004);
nor U2163 (N_2163,N_2079,N_2051);
xor U2164 (N_2164,N_2084,N_2071);
and U2165 (N_2165,N_2045,N_2067);
or U2166 (N_2166,N_2093,N_2064);
or U2167 (N_2167,N_2048,N_2065);
or U2168 (N_2168,N_2055,N_2002);
or U2169 (N_2169,N_2074,N_2050);
nand U2170 (N_2170,N_2005,N_2061);
nor U2171 (N_2171,N_2051,N_2098);
or U2172 (N_2172,N_2088,N_2016);
nor U2173 (N_2173,N_2023,N_2088);
or U2174 (N_2174,N_2093,N_2079);
nand U2175 (N_2175,N_2059,N_2065);
nand U2176 (N_2176,N_2056,N_2002);
nand U2177 (N_2177,N_2086,N_2050);
nor U2178 (N_2178,N_2071,N_2003);
or U2179 (N_2179,N_2007,N_2014);
nand U2180 (N_2180,N_2002,N_2088);
nand U2181 (N_2181,N_2025,N_2026);
and U2182 (N_2182,N_2087,N_2073);
and U2183 (N_2183,N_2091,N_2097);
nor U2184 (N_2184,N_2002,N_2085);
or U2185 (N_2185,N_2067,N_2054);
and U2186 (N_2186,N_2077,N_2022);
or U2187 (N_2187,N_2018,N_2080);
or U2188 (N_2188,N_2056,N_2069);
nand U2189 (N_2189,N_2040,N_2003);
nand U2190 (N_2190,N_2093,N_2095);
or U2191 (N_2191,N_2011,N_2078);
nand U2192 (N_2192,N_2063,N_2087);
nand U2193 (N_2193,N_2087,N_2037);
nor U2194 (N_2194,N_2069,N_2051);
or U2195 (N_2195,N_2068,N_2056);
nor U2196 (N_2196,N_2015,N_2010);
nor U2197 (N_2197,N_2050,N_2027);
and U2198 (N_2198,N_2076,N_2093);
nand U2199 (N_2199,N_2063,N_2015);
nor U2200 (N_2200,N_2187,N_2147);
nor U2201 (N_2201,N_2139,N_2149);
or U2202 (N_2202,N_2131,N_2121);
and U2203 (N_2203,N_2177,N_2146);
and U2204 (N_2204,N_2162,N_2199);
and U2205 (N_2205,N_2119,N_2148);
nand U2206 (N_2206,N_2120,N_2107);
nor U2207 (N_2207,N_2175,N_2114);
and U2208 (N_2208,N_2105,N_2143);
nand U2209 (N_2209,N_2125,N_2185);
nor U2210 (N_2210,N_2173,N_2118);
nand U2211 (N_2211,N_2158,N_2153);
nor U2212 (N_2212,N_2113,N_2128);
or U2213 (N_2213,N_2115,N_2197);
xnor U2214 (N_2214,N_2106,N_2111);
or U2215 (N_2215,N_2160,N_2135);
nand U2216 (N_2216,N_2117,N_2123);
xnor U2217 (N_2217,N_2150,N_2196);
nor U2218 (N_2218,N_2145,N_2133);
nand U2219 (N_2219,N_2180,N_2186);
nand U2220 (N_2220,N_2190,N_2193);
and U2221 (N_2221,N_2104,N_2109);
and U2222 (N_2222,N_2142,N_2168);
nor U2223 (N_2223,N_2138,N_2172);
or U2224 (N_2224,N_2194,N_2103);
or U2225 (N_2225,N_2176,N_2166);
nor U2226 (N_2226,N_2108,N_2179);
and U2227 (N_2227,N_2192,N_2191);
or U2228 (N_2228,N_2195,N_2183);
or U2229 (N_2229,N_2152,N_2124);
nor U2230 (N_2230,N_2112,N_2184);
or U2231 (N_2231,N_2169,N_2161);
nor U2232 (N_2232,N_2100,N_2141);
and U2233 (N_2233,N_2182,N_2136);
or U2234 (N_2234,N_2181,N_2126);
nor U2235 (N_2235,N_2132,N_2164);
xnor U2236 (N_2236,N_2157,N_2140);
nand U2237 (N_2237,N_2127,N_2188);
nor U2238 (N_2238,N_2110,N_2174);
nor U2239 (N_2239,N_2170,N_2171);
nand U2240 (N_2240,N_2163,N_2122);
and U2241 (N_2241,N_2165,N_2101);
and U2242 (N_2242,N_2178,N_2137);
nor U2243 (N_2243,N_2155,N_2159);
and U2244 (N_2244,N_2198,N_2154);
and U2245 (N_2245,N_2129,N_2156);
nor U2246 (N_2246,N_2151,N_2134);
or U2247 (N_2247,N_2116,N_2167);
or U2248 (N_2248,N_2102,N_2130);
nor U2249 (N_2249,N_2189,N_2144);
or U2250 (N_2250,N_2170,N_2184);
and U2251 (N_2251,N_2174,N_2108);
and U2252 (N_2252,N_2156,N_2196);
and U2253 (N_2253,N_2188,N_2169);
nor U2254 (N_2254,N_2135,N_2179);
or U2255 (N_2255,N_2131,N_2142);
xnor U2256 (N_2256,N_2124,N_2115);
nand U2257 (N_2257,N_2144,N_2116);
and U2258 (N_2258,N_2196,N_2173);
and U2259 (N_2259,N_2130,N_2145);
nor U2260 (N_2260,N_2156,N_2166);
or U2261 (N_2261,N_2136,N_2193);
nor U2262 (N_2262,N_2100,N_2197);
or U2263 (N_2263,N_2185,N_2142);
nand U2264 (N_2264,N_2198,N_2128);
or U2265 (N_2265,N_2170,N_2153);
nand U2266 (N_2266,N_2149,N_2181);
or U2267 (N_2267,N_2158,N_2167);
or U2268 (N_2268,N_2181,N_2154);
nand U2269 (N_2269,N_2130,N_2179);
or U2270 (N_2270,N_2109,N_2156);
or U2271 (N_2271,N_2124,N_2187);
and U2272 (N_2272,N_2150,N_2128);
or U2273 (N_2273,N_2103,N_2138);
and U2274 (N_2274,N_2147,N_2151);
nor U2275 (N_2275,N_2117,N_2124);
nor U2276 (N_2276,N_2194,N_2105);
nor U2277 (N_2277,N_2173,N_2113);
nor U2278 (N_2278,N_2158,N_2154);
and U2279 (N_2279,N_2101,N_2133);
nand U2280 (N_2280,N_2195,N_2130);
and U2281 (N_2281,N_2100,N_2165);
nand U2282 (N_2282,N_2113,N_2130);
nor U2283 (N_2283,N_2181,N_2121);
nand U2284 (N_2284,N_2160,N_2110);
nand U2285 (N_2285,N_2145,N_2104);
nor U2286 (N_2286,N_2180,N_2115);
nand U2287 (N_2287,N_2160,N_2133);
and U2288 (N_2288,N_2179,N_2189);
nand U2289 (N_2289,N_2144,N_2153);
or U2290 (N_2290,N_2197,N_2107);
or U2291 (N_2291,N_2187,N_2199);
and U2292 (N_2292,N_2151,N_2179);
nor U2293 (N_2293,N_2194,N_2190);
or U2294 (N_2294,N_2164,N_2140);
or U2295 (N_2295,N_2142,N_2151);
nor U2296 (N_2296,N_2180,N_2147);
or U2297 (N_2297,N_2182,N_2169);
and U2298 (N_2298,N_2161,N_2159);
nor U2299 (N_2299,N_2181,N_2124);
nand U2300 (N_2300,N_2248,N_2203);
or U2301 (N_2301,N_2263,N_2289);
or U2302 (N_2302,N_2286,N_2200);
nand U2303 (N_2303,N_2222,N_2245);
or U2304 (N_2304,N_2228,N_2214);
nor U2305 (N_2305,N_2215,N_2246);
and U2306 (N_2306,N_2235,N_2249);
nor U2307 (N_2307,N_2239,N_2251);
and U2308 (N_2308,N_2219,N_2208);
or U2309 (N_2309,N_2240,N_2210);
or U2310 (N_2310,N_2247,N_2252);
nor U2311 (N_2311,N_2216,N_2297);
or U2312 (N_2312,N_2271,N_2272);
nor U2313 (N_2313,N_2242,N_2296);
nand U2314 (N_2314,N_2298,N_2294);
nor U2315 (N_2315,N_2260,N_2233);
and U2316 (N_2316,N_2254,N_2264);
and U2317 (N_2317,N_2244,N_2268);
nor U2318 (N_2318,N_2241,N_2284);
nand U2319 (N_2319,N_2231,N_2281);
nor U2320 (N_2320,N_2236,N_2265);
nor U2321 (N_2321,N_2259,N_2274);
or U2322 (N_2322,N_2204,N_2270);
and U2323 (N_2323,N_2225,N_2266);
and U2324 (N_2324,N_2269,N_2217);
and U2325 (N_2325,N_2292,N_2211);
nor U2326 (N_2326,N_2232,N_2273);
or U2327 (N_2327,N_2221,N_2223);
and U2328 (N_2328,N_2220,N_2250);
or U2329 (N_2329,N_2288,N_2279);
nand U2330 (N_2330,N_2299,N_2229);
nand U2331 (N_2331,N_2291,N_2293);
nor U2332 (N_2332,N_2205,N_2257);
nand U2333 (N_2333,N_2290,N_2280);
or U2334 (N_2334,N_2243,N_2267);
or U2335 (N_2335,N_2237,N_2218);
or U2336 (N_2336,N_2230,N_2224);
nor U2337 (N_2337,N_2209,N_2253);
nor U2338 (N_2338,N_2277,N_2226);
nor U2339 (N_2339,N_2276,N_2212);
nor U2340 (N_2340,N_2201,N_2282);
xnor U2341 (N_2341,N_2207,N_2255);
nand U2342 (N_2342,N_2213,N_2295);
nor U2343 (N_2343,N_2285,N_2227);
nor U2344 (N_2344,N_2258,N_2275);
or U2345 (N_2345,N_2278,N_2262);
and U2346 (N_2346,N_2206,N_2261);
nand U2347 (N_2347,N_2283,N_2234);
or U2348 (N_2348,N_2256,N_2202);
nand U2349 (N_2349,N_2287,N_2238);
and U2350 (N_2350,N_2245,N_2242);
and U2351 (N_2351,N_2224,N_2231);
nand U2352 (N_2352,N_2225,N_2229);
and U2353 (N_2353,N_2253,N_2275);
or U2354 (N_2354,N_2273,N_2245);
nand U2355 (N_2355,N_2231,N_2284);
nor U2356 (N_2356,N_2209,N_2216);
nor U2357 (N_2357,N_2271,N_2207);
and U2358 (N_2358,N_2277,N_2234);
and U2359 (N_2359,N_2265,N_2212);
nor U2360 (N_2360,N_2228,N_2280);
or U2361 (N_2361,N_2230,N_2204);
or U2362 (N_2362,N_2230,N_2207);
and U2363 (N_2363,N_2274,N_2243);
nand U2364 (N_2364,N_2279,N_2217);
nor U2365 (N_2365,N_2228,N_2255);
nand U2366 (N_2366,N_2234,N_2266);
or U2367 (N_2367,N_2298,N_2284);
and U2368 (N_2368,N_2278,N_2223);
or U2369 (N_2369,N_2255,N_2284);
and U2370 (N_2370,N_2213,N_2203);
nor U2371 (N_2371,N_2213,N_2294);
nor U2372 (N_2372,N_2232,N_2276);
xnor U2373 (N_2373,N_2244,N_2260);
xor U2374 (N_2374,N_2247,N_2212);
or U2375 (N_2375,N_2241,N_2262);
nand U2376 (N_2376,N_2218,N_2288);
nor U2377 (N_2377,N_2222,N_2206);
or U2378 (N_2378,N_2203,N_2264);
and U2379 (N_2379,N_2249,N_2244);
nand U2380 (N_2380,N_2263,N_2246);
or U2381 (N_2381,N_2217,N_2253);
and U2382 (N_2382,N_2206,N_2202);
nand U2383 (N_2383,N_2207,N_2222);
nor U2384 (N_2384,N_2241,N_2268);
and U2385 (N_2385,N_2228,N_2237);
nand U2386 (N_2386,N_2242,N_2295);
nand U2387 (N_2387,N_2240,N_2218);
xnor U2388 (N_2388,N_2253,N_2258);
nor U2389 (N_2389,N_2271,N_2239);
nor U2390 (N_2390,N_2203,N_2216);
nand U2391 (N_2391,N_2245,N_2248);
nor U2392 (N_2392,N_2224,N_2259);
nor U2393 (N_2393,N_2271,N_2263);
nand U2394 (N_2394,N_2218,N_2287);
nand U2395 (N_2395,N_2262,N_2249);
or U2396 (N_2396,N_2244,N_2239);
or U2397 (N_2397,N_2286,N_2284);
nand U2398 (N_2398,N_2233,N_2220);
or U2399 (N_2399,N_2217,N_2263);
nor U2400 (N_2400,N_2304,N_2363);
nor U2401 (N_2401,N_2353,N_2336);
nand U2402 (N_2402,N_2306,N_2317);
nor U2403 (N_2403,N_2382,N_2378);
or U2404 (N_2404,N_2332,N_2364);
nand U2405 (N_2405,N_2349,N_2385);
or U2406 (N_2406,N_2322,N_2381);
nand U2407 (N_2407,N_2374,N_2320);
nor U2408 (N_2408,N_2330,N_2370);
nand U2409 (N_2409,N_2391,N_2362);
and U2410 (N_2410,N_2329,N_2326);
nand U2411 (N_2411,N_2371,N_2303);
nand U2412 (N_2412,N_2325,N_2309);
nand U2413 (N_2413,N_2394,N_2343);
nor U2414 (N_2414,N_2323,N_2331);
nand U2415 (N_2415,N_2384,N_2351);
or U2416 (N_2416,N_2339,N_2399);
or U2417 (N_2417,N_2380,N_2354);
nand U2418 (N_2418,N_2396,N_2307);
and U2419 (N_2419,N_2383,N_2379);
nor U2420 (N_2420,N_2376,N_2398);
or U2421 (N_2421,N_2366,N_2301);
or U2422 (N_2422,N_2367,N_2345);
and U2423 (N_2423,N_2348,N_2327);
nand U2424 (N_2424,N_2318,N_2324);
nor U2425 (N_2425,N_2352,N_2333);
or U2426 (N_2426,N_2355,N_2377);
and U2427 (N_2427,N_2337,N_2347);
and U2428 (N_2428,N_2365,N_2300);
nand U2429 (N_2429,N_2328,N_2321);
or U2430 (N_2430,N_2315,N_2341);
xor U2431 (N_2431,N_2360,N_2373);
nor U2432 (N_2432,N_2312,N_2397);
nand U2433 (N_2433,N_2392,N_2335);
and U2434 (N_2434,N_2314,N_2311);
nand U2435 (N_2435,N_2361,N_2358);
and U2436 (N_2436,N_2368,N_2344);
nor U2437 (N_2437,N_2308,N_2393);
or U2438 (N_2438,N_2319,N_2359);
nand U2439 (N_2439,N_2390,N_2387);
or U2440 (N_2440,N_2389,N_2356);
or U2441 (N_2441,N_2388,N_2375);
nand U2442 (N_2442,N_2338,N_2340);
nand U2443 (N_2443,N_2305,N_2386);
nor U2444 (N_2444,N_2369,N_2395);
nor U2445 (N_2445,N_2310,N_2372);
and U2446 (N_2446,N_2316,N_2302);
or U2447 (N_2447,N_2334,N_2357);
nor U2448 (N_2448,N_2350,N_2342);
nand U2449 (N_2449,N_2346,N_2313);
or U2450 (N_2450,N_2332,N_2350);
and U2451 (N_2451,N_2333,N_2335);
nand U2452 (N_2452,N_2324,N_2366);
and U2453 (N_2453,N_2363,N_2313);
or U2454 (N_2454,N_2362,N_2308);
or U2455 (N_2455,N_2384,N_2338);
or U2456 (N_2456,N_2378,N_2347);
or U2457 (N_2457,N_2334,N_2344);
and U2458 (N_2458,N_2307,N_2335);
nor U2459 (N_2459,N_2326,N_2302);
and U2460 (N_2460,N_2358,N_2300);
nand U2461 (N_2461,N_2384,N_2385);
and U2462 (N_2462,N_2358,N_2314);
nand U2463 (N_2463,N_2375,N_2378);
or U2464 (N_2464,N_2316,N_2340);
and U2465 (N_2465,N_2341,N_2330);
and U2466 (N_2466,N_2339,N_2366);
and U2467 (N_2467,N_2340,N_2355);
or U2468 (N_2468,N_2375,N_2353);
nand U2469 (N_2469,N_2311,N_2356);
and U2470 (N_2470,N_2306,N_2338);
or U2471 (N_2471,N_2301,N_2389);
or U2472 (N_2472,N_2316,N_2331);
nor U2473 (N_2473,N_2372,N_2343);
or U2474 (N_2474,N_2323,N_2301);
nand U2475 (N_2475,N_2373,N_2362);
nor U2476 (N_2476,N_2339,N_2392);
or U2477 (N_2477,N_2390,N_2348);
nand U2478 (N_2478,N_2374,N_2324);
and U2479 (N_2479,N_2350,N_2393);
nor U2480 (N_2480,N_2399,N_2324);
or U2481 (N_2481,N_2383,N_2359);
and U2482 (N_2482,N_2318,N_2308);
and U2483 (N_2483,N_2352,N_2390);
or U2484 (N_2484,N_2356,N_2303);
nand U2485 (N_2485,N_2330,N_2316);
and U2486 (N_2486,N_2303,N_2378);
nor U2487 (N_2487,N_2377,N_2374);
or U2488 (N_2488,N_2374,N_2332);
or U2489 (N_2489,N_2363,N_2355);
or U2490 (N_2490,N_2393,N_2362);
nor U2491 (N_2491,N_2340,N_2366);
nand U2492 (N_2492,N_2382,N_2366);
or U2493 (N_2493,N_2329,N_2382);
or U2494 (N_2494,N_2367,N_2346);
and U2495 (N_2495,N_2329,N_2387);
or U2496 (N_2496,N_2325,N_2320);
or U2497 (N_2497,N_2307,N_2333);
nor U2498 (N_2498,N_2366,N_2357);
nor U2499 (N_2499,N_2393,N_2383);
and U2500 (N_2500,N_2495,N_2486);
nand U2501 (N_2501,N_2444,N_2466);
nand U2502 (N_2502,N_2440,N_2457);
nand U2503 (N_2503,N_2409,N_2458);
and U2504 (N_2504,N_2428,N_2438);
and U2505 (N_2505,N_2482,N_2410);
and U2506 (N_2506,N_2418,N_2412);
or U2507 (N_2507,N_2445,N_2405);
nand U2508 (N_2508,N_2441,N_2452);
and U2509 (N_2509,N_2433,N_2450);
nor U2510 (N_2510,N_2416,N_2429);
nor U2511 (N_2511,N_2487,N_2456);
nand U2512 (N_2512,N_2406,N_2432);
or U2513 (N_2513,N_2446,N_2474);
nor U2514 (N_2514,N_2413,N_2415);
or U2515 (N_2515,N_2430,N_2496);
and U2516 (N_2516,N_2483,N_2431);
or U2517 (N_2517,N_2476,N_2451);
nor U2518 (N_2518,N_2453,N_2449);
nand U2519 (N_2519,N_2499,N_2434);
nand U2520 (N_2520,N_2493,N_2491);
nor U2521 (N_2521,N_2471,N_2464);
or U2522 (N_2522,N_2484,N_2439);
or U2523 (N_2523,N_2423,N_2421);
and U2524 (N_2524,N_2447,N_2494);
nand U2525 (N_2525,N_2463,N_2419);
nor U2526 (N_2526,N_2492,N_2498);
and U2527 (N_2527,N_2426,N_2477);
nor U2528 (N_2528,N_2489,N_2472);
nor U2529 (N_2529,N_2408,N_2459);
nor U2530 (N_2530,N_2437,N_2401);
nand U2531 (N_2531,N_2490,N_2465);
nor U2532 (N_2532,N_2481,N_2414);
nand U2533 (N_2533,N_2473,N_2425);
or U2534 (N_2534,N_2461,N_2455);
nor U2535 (N_2535,N_2448,N_2402);
and U2536 (N_2536,N_2467,N_2475);
and U2537 (N_2537,N_2443,N_2436);
and U2538 (N_2538,N_2403,N_2479);
nand U2539 (N_2539,N_2460,N_2400);
or U2540 (N_2540,N_2454,N_2485);
or U2541 (N_2541,N_2411,N_2497);
nand U2542 (N_2542,N_2427,N_2442);
nand U2543 (N_2543,N_2422,N_2424);
and U2544 (N_2544,N_2435,N_2462);
nand U2545 (N_2545,N_2478,N_2470);
nor U2546 (N_2546,N_2480,N_2404);
and U2547 (N_2547,N_2468,N_2420);
or U2548 (N_2548,N_2407,N_2469);
or U2549 (N_2549,N_2488,N_2417);
and U2550 (N_2550,N_2405,N_2418);
nor U2551 (N_2551,N_2463,N_2422);
nor U2552 (N_2552,N_2453,N_2409);
or U2553 (N_2553,N_2462,N_2469);
nand U2554 (N_2554,N_2409,N_2439);
or U2555 (N_2555,N_2434,N_2412);
or U2556 (N_2556,N_2495,N_2404);
and U2557 (N_2557,N_2410,N_2463);
and U2558 (N_2558,N_2496,N_2417);
nor U2559 (N_2559,N_2499,N_2475);
or U2560 (N_2560,N_2471,N_2479);
nor U2561 (N_2561,N_2423,N_2410);
nand U2562 (N_2562,N_2406,N_2495);
nor U2563 (N_2563,N_2499,N_2476);
nor U2564 (N_2564,N_2448,N_2452);
or U2565 (N_2565,N_2406,N_2422);
nor U2566 (N_2566,N_2434,N_2478);
and U2567 (N_2567,N_2441,N_2446);
nand U2568 (N_2568,N_2454,N_2406);
nor U2569 (N_2569,N_2465,N_2448);
or U2570 (N_2570,N_2419,N_2489);
nand U2571 (N_2571,N_2414,N_2480);
or U2572 (N_2572,N_2425,N_2464);
and U2573 (N_2573,N_2419,N_2475);
and U2574 (N_2574,N_2481,N_2428);
and U2575 (N_2575,N_2498,N_2479);
nand U2576 (N_2576,N_2470,N_2490);
and U2577 (N_2577,N_2455,N_2498);
nor U2578 (N_2578,N_2477,N_2425);
or U2579 (N_2579,N_2450,N_2465);
or U2580 (N_2580,N_2476,N_2459);
nand U2581 (N_2581,N_2418,N_2400);
or U2582 (N_2582,N_2474,N_2464);
xor U2583 (N_2583,N_2485,N_2472);
nor U2584 (N_2584,N_2495,N_2436);
nor U2585 (N_2585,N_2436,N_2418);
xnor U2586 (N_2586,N_2471,N_2465);
nand U2587 (N_2587,N_2413,N_2494);
or U2588 (N_2588,N_2473,N_2494);
and U2589 (N_2589,N_2462,N_2482);
nor U2590 (N_2590,N_2474,N_2444);
nor U2591 (N_2591,N_2484,N_2473);
nor U2592 (N_2592,N_2412,N_2405);
and U2593 (N_2593,N_2481,N_2467);
nand U2594 (N_2594,N_2418,N_2456);
and U2595 (N_2595,N_2458,N_2438);
nor U2596 (N_2596,N_2442,N_2485);
and U2597 (N_2597,N_2434,N_2449);
or U2598 (N_2598,N_2469,N_2484);
nand U2599 (N_2599,N_2413,N_2401);
nand U2600 (N_2600,N_2515,N_2512);
xnor U2601 (N_2601,N_2513,N_2564);
or U2602 (N_2602,N_2578,N_2541);
and U2603 (N_2603,N_2579,N_2577);
and U2604 (N_2604,N_2553,N_2544);
or U2605 (N_2605,N_2556,N_2500);
or U2606 (N_2606,N_2521,N_2599);
or U2607 (N_2607,N_2528,N_2571);
nor U2608 (N_2608,N_2555,N_2565);
nor U2609 (N_2609,N_2581,N_2584);
nor U2610 (N_2610,N_2530,N_2563);
nor U2611 (N_2611,N_2519,N_2551);
or U2612 (N_2612,N_2550,N_2595);
or U2613 (N_2613,N_2575,N_2524);
nor U2614 (N_2614,N_2545,N_2590);
nor U2615 (N_2615,N_2502,N_2529);
nand U2616 (N_2616,N_2503,N_2548);
or U2617 (N_2617,N_2535,N_2586);
and U2618 (N_2618,N_2570,N_2525);
and U2619 (N_2619,N_2508,N_2576);
nand U2620 (N_2620,N_2543,N_2574);
or U2621 (N_2621,N_2589,N_2592);
or U2622 (N_2622,N_2510,N_2533);
or U2623 (N_2623,N_2527,N_2585);
or U2624 (N_2624,N_2588,N_2557);
and U2625 (N_2625,N_2542,N_2504);
or U2626 (N_2626,N_2554,N_2507);
nor U2627 (N_2627,N_2559,N_2509);
or U2628 (N_2628,N_2552,N_2511);
or U2629 (N_2629,N_2567,N_2547);
nand U2630 (N_2630,N_2580,N_2520);
nand U2631 (N_2631,N_2568,N_2596);
nand U2632 (N_2632,N_2546,N_2566);
or U2633 (N_2633,N_2523,N_2549);
nand U2634 (N_2634,N_2598,N_2591);
and U2635 (N_2635,N_2593,N_2517);
or U2636 (N_2636,N_2572,N_2522);
or U2637 (N_2637,N_2561,N_2536);
nor U2638 (N_2638,N_2506,N_2532);
or U2639 (N_2639,N_2582,N_2538);
nand U2640 (N_2640,N_2594,N_2534);
nand U2641 (N_2641,N_2558,N_2573);
nor U2642 (N_2642,N_2540,N_2531);
nor U2643 (N_2643,N_2562,N_2518);
nor U2644 (N_2644,N_2583,N_2560);
and U2645 (N_2645,N_2505,N_2539);
nand U2646 (N_2646,N_2516,N_2587);
nand U2647 (N_2647,N_2537,N_2597);
nor U2648 (N_2648,N_2514,N_2526);
nor U2649 (N_2649,N_2569,N_2501);
and U2650 (N_2650,N_2512,N_2595);
nand U2651 (N_2651,N_2507,N_2510);
nand U2652 (N_2652,N_2572,N_2560);
nand U2653 (N_2653,N_2563,N_2595);
or U2654 (N_2654,N_2584,N_2544);
or U2655 (N_2655,N_2510,N_2535);
nand U2656 (N_2656,N_2581,N_2598);
nor U2657 (N_2657,N_2520,N_2524);
and U2658 (N_2658,N_2534,N_2585);
or U2659 (N_2659,N_2571,N_2529);
or U2660 (N_2660,N_2578,N_2527);
nor U2661 (N_2661,N_2554,N_2582);
nand U2662 (N_2662,N_2558,N_2512);
or U2663 (N_2663,N_2543,N_2568);
or U2664 (N_2664,N_2553,N_2532);
nand U2665 (N_2665,N_2589,N_2543);
xnor U2666 (N_2666,N_2592,N_2554);
xnor U2667 (N_2667,N_2521,N_2518);
xnor U2668 (N_2668,N_2564,N_2508);
nand U2669 (N_2669,N_2545,N_2530);
nor U2670 (N_2670,N_2572,N_2531);
or U2671 (N_2671,N_2581,N_2550);
and U2672 (N_2672,N_2510,N_2532);
or U2673 (N_2673,N_2545,N_2540);
and U2674 (N_2674,N_2536,N_2529);
and U2675 (N_2675,N_2593,N_2515);
or U2676 (N_2676,N_2539,N_2594);
and U2677 (N_2677,N_2545,N_2546);
nor U2678 (N_2678,N_2505,N_2524);
nor U2679 (N_2679,N_2553,N_2575);
or U2680 (N_2680,N_2519,N_2572);
or U2681 (N_2681,N_2566,N_2550);
or U2682 (N_2682,N_2507,N_2537);
nand U2683 (N_2683,N_2594,N_2592);
nand U2684 (N_2684,N_2553,N_2513);
nand U2685 (N_2685,N_2524,N_2541);
xor U2686 (N_2686,N_2549,N_2568);
and U2687 (N_2687,N_2563,N_2583);
nor U2688 (N_2688,N_2516,N_2566);
or U2689 (N_2689,N_2545,N_2567);
nand U2690 (N_2690,N_2539,N_2562);
nand U2691 (N_2691,N_2507,N_2559);
or U2692 (N_2692,N_2579,N_2530);
nand U2693 (N_2693,N_2597,N_2573);
xnor U2694 (N_2694,N_2594,N_2536);
or U2695 (N_2695,N_2543,N_2520);
or U2696 (N_2696,N_2508,N_2504);
nor U2697 (N_2697,N_2596,N_2580);
or U2698 (N_2698,N_2513,N_2518);
and U2699 (N_2699,N_2538,N_2573);
nand U2700 (N_2700,N_2670,N_2662);
nand U2701 (N_2701,N_2651,N_2608);
nor U2702 (N_2702,N_2673,N_2652);
nor U2703 (N_2703,N_2602,N_2618);
and U2704 (N_2704,N_2635,N_2684);
or U2705 (N_2705,N_2639,N_2656);
and U2706 (N_2706,N_2621,N_2630);
or U2707 (N_2707,N_2692,N_2629);
and U2708 (N_2708,N_2641,N_2697);
xnor U2709 (N_2709,N_2658,N_2623);
nand U2710 (N_2710,N_2661,N_2606);
nand U2711 (N_2711,N_2698,N_2681);
nor U2712 (N_2712,N_2647,N_2686);
or U2713 (N_2713,N_2677,N_2694);
nand U2714 (N_2714,N_2685,N_2678);
and U2715 (N_2715,N_2669,N_2616);
nand U2716 (N_2716,N_2613,N_2626);
or U2717 (N_2717,N_2695,N_2693);
xnor U2718 (N_2718,N_2633,N_2603);
nor U2719 (N_2719,N_2612,N_2675);
or U2720 (N_2720,N_2649,N_2696);
or U2721 (N_2721,N_2691,N_2659);
and U2722 (N_2722,N_2699,N_2674);
nand U2723 (N_2723,N_2620,N_2636);
or U2724 (N_2724,N_2624,N_2682);
or U2725 (N_2725,N_2655,N_2689);
or U2726 (N_2726,N_2680,N_2657);
nor U2727 (N_2727,N_2676,N_2634);
or U2728 (N_2728,N_2600,N_2642);
and U2729 (N_2729,N_2628,N_2671);
and U2730 (N_2730,N_2643,N_2645);
nor U2731 (N_2731,N_2663,N_2625);
or U2732 (N_2732,N_2605,N_2640);
nor U2733 (N_2733,N_2660,N_2638);
or U2734 (N_2734,N_2679,N_2666);
or U2735 (N_2735,N_2622,N_2607);
nor U2736 (N_2736,N_2611,N_2683);
or U2737 (N_2737,N_2672,N_2690);
nand U2738 (N_2738,N_2609,N_2664);
and U2739 (N_2739,N_2687,N_2601);
or U2740 (N_2740,N_2688,N_2615);
nand U2741 (N_2741,N_2627,N_2637);
and U2742 (N_2742,N_2610,N_2665);
nor U2743 (N_2743,N_2632,N_2650);
and U2744 (N_2744,N_2654,N_2646);
and U2745 (N_2745,N_2648,N_2644);
nor U2746 (N_2746,N_2668,N_2653);
nor U2747 (N_2747,N_2604,N_2619);
and U2748 (N_2748,N_2617,N_2667);
nand U2749 (N_2749,N_2631,N_2614);
or U2750 (N_2750,N_2682,N_2675);
or U2751 (N_2751,N_2681,N_2600);
and U2752 (N_2752,N_2671,N_2618);
xnor U2753 (N_2753,N_2629,N_2691);
nor U2754 (N_2754,N_2678,N_2638);
or U2755 (N_2755,N_2636,N_2642);
or U2756 (N_2756,N_2676,N_2609);
nor U2757 (N_2757,N_2679,N_2629);
nor U2758 (N_2758,N_2608,N_2611);
nand U2759 (N_2759,N_2619,N_2639);
and U2760 (N_2760,N_2655,N_2635);
nand U2761 (N_2761,N_2645,N_2693);
or U2762 (N_2762,N_2677,N_2697);
or U2763 (N_2763,N_2639,N_2666);
or U2764 (N_2764,N_2638,N_2665);
or U2765 (N_2765,N_2655,N_2673);
or U2766 (N_2766,N_2646,N_2601);
nand U2767 (N_2767,N_2652,N_2660);
and U2768 (N_2768,N_2692,N_2628);
nand U2769 (N_2769,N_2652,N_2650);
and U2770 (N_2770,N_2633,N_2661);
nand U2771 (N_2771,N_2611,N_2666);
xnor U2772 (N_2772,N_2662,N_2643);
nand U2773 (N_2773,N_2655,N_2615);
nor U2774 (N_2774,N_2698,N_2677);
and U2775 (N_2775,N_2646,N_2642);
nor U2776 (N_2776,N_2694,N_2650);
nand U2777 (N_2777,N_2697,N_2645);
or U2778 (N_2778,N_2604,N_2665);
nor U2779 (N_2779,N_2611,N_2638);
and U2780 (N_2780,N_2645,N_2675);
nor U2781 (N_2781,N_2641,N_2621);
nand U2782 (N_2782,N_2603,N_2608);
or U2783 (N_2783,N_2600,N_2643);
or U2784 (N_2784,N_2696,N_2634);
nand U2785 (N_2785,N_2630,N_2654);
nand U2786 (N_2786,N_2690,N_2640);
and U2787 (N_2787,N_2686,N_2622);
and U2788 (N_2788,N_2607,N_2631);
nand U2789 (N_2789,N_2679,N_2648);
nor U2790 (N_2790,N_2632,N_2672);
and U2791 (N_2791,N_2666,N_2654);
nor U2792 (N_2792,N_2644,N_2643);
nand U2793 (N_2793,N_2632,N_2615);
nand U2794 (N_2794,N_2613,N_2641);
or U2795 (N_2795,N_2660,N_2605);
nand U2796 (N_2796,N_2670,N_2600);
nor U2797 (N_2797,N_2643,N_2659);
or U2798 (N_2798,N_2610,N_2633);
or U2799 (N_2799,N_2614,N_2642);
nand U2800 (N_2800,N_2763,N_2744);
nor U2801 (N_2801,N_2700,N_2716);
xnor U2802 (N_2802,N_2720,N_2746);
nand U2803 (N_2803,N_2701,N_2710);
nand U2804 (N_2804,N_2783,N_2713);
nand U2805 (N_2805,N_2762,N_2768);
and U2806 (N_2806,N_2789,N_2704);
nand U2807 (N_2807,N_2711,N_2794);
nor U2808 (N_2808,N_2736,N_2776);
or U2809 (N_2809,N_2740,N_2772);
xor U2810 (N_2810,N_2766,N_2737);
nand U2811 (N_2811,N_2753,N_2721);
nor U2812 (N_2812,N_2738,N_2729);
nand U2813 (N_2813,N_2715,N_2791);
nand U2814 (N_2814,N_2760,N_2742);
or U2815 (N_2815,N_2725,N_2767);
nor U2816 (N_2816,N_2702,N_2795);
and U2817 (N_2817,N_2792,N_2788);
nand U2818 (N_2818,N_2796,N_2733);
or U2819 (N_2819,N_2761,N_2751);
and U2820 (N_2820,N_2784,N_2741);
xor U2821 (N_2821,N_2735,N_2775);
or U2822 (N_2822,N_2764,N_2756);
or U2823 (N_2823,N_2706,N_2727);
or U2824 (N_2824,N_2790,N_2745);
xnor U2825 (N_2825,N_2750,N_2730);
nor U2826 (N_2826,N_2748,N_2754);
or U2827 (N_2827,N_2728,N_2758);
nor U2828 (N_2828,N_2717,N_2726);
or U2829 (N_2829,N_2759,N_2797);
or U2830 (N_2830,N_2781,N_2707);
nand U2831 (N_2831,N_2774,N_2752);
and U2832 (N_2832,N_2749,N_2787);
and U2833 (N_2833,N_2769,N_2778);
and U2834 (N_2834,N_2793,N_2757);
and U2835 (N_2835,N_2718,N_2732);
nand U2836 (N_2836,N_2770,N_2722);
nor U2837 (N_2837,N_2786,N_2798);
nor U2838 (N_2838,N_2765,N_2782);
nor U2839 (N_2839,N_2712,N_2719);
and U2840 (N_2840,N_2771,N_2773);
and U2841 (N_2841,N_2743,N_2705);
or U2842 (N_2842,N_2714,N_2785);
and U2843 (N_2843,N_2780,N_2799);
nand U2844 (N_2844,N_2703,N_2739);
or U2845 (N_2845,N_2779,N_2709);
nor U2846 (N_2846,N_2731,N_2734);
nor U2847 (N_2847,N_2724,N_2747);
or U2848 (N_2848,N_2708,N_2723);
nand U2849 (N_2849,N_2755,N_2777);
and U2850 (N_2850,N_2737,N_2739);
or U2851 (N_2851,N_2788,N_2720);
nand U2852 (N_2852,N_2780,N_2786);
nand U2853 (N_2853,N_2722,N_2754);
nor U2854 (N_2854,N_2719,N_2771);
or U2855 (N_2855,N_2745,N_2721);
or U2856 (N_2856,N_2786,N_2793);
or U2857 (N_2857,N_2786,N_2706);
nor U2858 (N_2858,N_2715,N_2728);
and U2859 (N_2859,N_2760,N_2766);
nor U2860 (N_2860,N_2737,N_2758);
nor U2861 (N_2861,N_2701,N_2767);
nand U2862 (N_2862,N_2769,N_2739);
nor U2863 (N_2863,N_2719,N_2706);
or U2864 (N_2864,N_2700,N_2737);
nand U2865 (N_2865,N_2725,N_2746);
nand U2866 (N_2866,N_2751,N_2759);
and U2867 (N_2867,N_2743,N_2737);
nor U2868 (N_2868,N_2724,N_2745);
or U2869 (N_2869,N_2782,N_2713);
xnor U2870 (N_2870,N_2713,N_2760);
or U2871 (N_2871,N_2799,N_2741);
or U2872 (N_2872,N_2786,N_2783);
nor U2873 (N_2873,N_2707,N_2752);
and U2874 (N_2874,N_2725,N_2795);
and U2875 (N_2875,N_2797,N_2794);
or U2876 (N_2876,N_2705,N_2763);
nor U2877 (N_2877,N_2757,N_2753);
or U2878 (N_2878,N_2795,N_2751);
and U2879 (N_2879,N_2707,N_2782);
nand U2880 (N_2880,N_2782,N_2771);
nand U2881 (N_2881,N_2786,N_2792);
or U2882 (N_2882,N_2735,N_2728);
and U2883 (N_2883,N_2731,N_2740);
nand U2884 (N_2884,N_2796,N_2774);
nand U2885 (N_2885,N_2797,N_2755);
nand U2886 (N_2886,N_2778,N_2742);
nor U2887 (N_2887,N_2755,N_2769);
nand U2888 (N_2888,N_2709,N_2722);
nand U2889 (N_2889,N_2771,N_2774);
and U2890 (N_2890,N_2749,N_2750);
nor U2891 (N_2891,N_2780,N_2765);
nand U2892 (N_2892,N_2768,N_2713);
nand U2893 (N_2893,N_2764,N_2721);
nor U2894 (N_2894,N_2791,N_2723);
or U2895 (N_2895,N_2770,N_2788);
nor U2896 (N_2896,N_2725,N_2704);
nor U2897 (N_2897,N_2764,N_2793);
and U2898 (N_2898,N_2751,N_2756);
or U2899 (N_2899,N_2786,N_2733);
and U2900 (N_2900,N_2829,N_2885);
nor U2901 (N_2901,N_2865,N_2894);
and U2902 (N_2902,N_2826,N_2876);
nand U2903 (N_2903,N_2804,N_2847);
or U2904 (N_2904,N_2802,N_2891);
and U2905 (N_2905,N_2858,N_2848);
and U2906 (N_2906,N_2805,N_2837);
and U2907 (N_2907,N_2831,N_2857);
or U2908 (N_2908,N_2841,N_2806);
and U2909 (N_2909,N_2836,N_2861);
nand U2910 (N_2910,N_2842,N_2873);
nor U2911 (N_2911,N_2889,N_2877);
nand U2912 (N_2912,N_2834,N_2881);
or U2913 (N_2913,N_2807,N_2815);
nor U2914 (N_2914,N_2884,N_2833);
nand U2915 (N_2915,N_2882,N_2869);
nor U2916 (N_2916,N_2895,N_2803);
nor U2917 (N_2917,N_2886,N_2855);
xnor U2918 (N_2918,N_2880,N_2812);
nand U2919 (N_2919,N_2817,N_2823);
or U2920 (N_2920,N_2888,N_2813);
nand U2921 (N_2921,N_2890,N_2808);
or U2922 (N_2922,N_2820,N_2879);
and U2923 (N_2923,N_2859,N_2830);
nand U2924 (N_2924,N_2893,N_2868);
and U2925 (N_2925,N_2878,N_2821);
nand U2926 (N_2926,N_2846,N_2863);
or U2927 (N_2927,N_2883,N_2898);
nand U2928 (N_2928,N_2874,N_2853);
and U2929 (N_2929,N_2828,N_2892);
and U2930 (N_2930,N_2851,N_2896);
nand U2931 (N_2931,N_2819,N_2822);
and U2932 (N_2932,N_2816,N_2844);
nand U2933 (N_2933,N_2810,N_2860);
and U2934 (N_2934,N_2864,N_2856);
and U2935 (N_2935,N_2832,N_2897);
and U2936 (N_2936,N_2850,N_2866);
nor U2937 (N_2937,N_2870,N_2835);
nand U2938 (N_2938,N_2809,N_2843);
nand U2939 (N_2939,N_2872,N_2875);
and U2940 (N_2940,N_2840,N_2825);
nand U2941 (N_2941,N_2839,N_2818);
and U2942 (N_2942,N_2862,N_2827);
nand U2943 (N_2943,N_2871,N_2814);
or U2944 (N_2944,N_2849,N_2838);
and U2945 (N_2945,N_2824,N_2801);
and U2946 (N_2946,N_2867,N_2852);
nand U2947 (N_2947,N_2800,N_2811);
and U2948 (N_2948,N_2899,N_2854);
and U2949 (N_2949,N_2845,N_2887);
nand U2950 (N_2950,N_2866,N_2826);
nor U2951 (N_2951,N_2835,N_2894);
nand U2952 (N_2952,N_2840,N_2812);
xor U2953 (N_2953,N_2852,N_2825);
or U2954 (N_2954,N_2859,N_2807);
nand U2955 (N_2955,N_2858,N_2815);
and U2956 (N_2956,N_2887,N_2852);
nand U2957 (N_2957,N_2843,N_2859);
nand U2958 (N_2958,N_2873,N_2864);
and U2959 (N_2959,N_2854,N_2879);
and U2960 (N_2960,N_2800,N_2889);
and U2961 (N_2961,N_2841,N_2829);
nor U2962 (N_2962,N_2861,N_2808);
nor U2963 (N_2963,N_2800,N_2877);
nor U2964 (N_2964,N_2840,N_2853);
nor U2965 (N_2965,N_2895,N_2813);
nor U2966 (N_2966,N_2827,N_2888);
or U2967 (N_2967,N_2899,N_2871);
nand U2968 (N_2968,N_2865,N_2890);
nor U2969 (N_2969,N_2801,N_2888);
nor U2970 (N_2970,N_2867,N_2882);
or U2971 (N_2971,N_2888,N_2815);
nand U2972 (N_2972,N_2891,N_2872);
nand U2973 (N_2973,N_2800,N_2861);
or U2974 (N_2974,N_2845,N_2803);
and U2975 (N_2975,N_2870,N_2883);
nand U2976 (N_2976,N_2850,N_2899);
nor U2977 (N_2977,N_2888,N_2808);
nand U2978 (N_2978,N_2831,N_2892);
or U2979 (N_2979,N_2878,N_2839);
or U2980 (N_2980,N_2808,N_2822);
nand U2981 (N_2981,N_2810,N_2894);
and U2982 (N_2982,N_2802,N_2853);
and U2983 (N_2983,N_2842,N_2899);
and U2984 (N_2984,N_2879,N_2898);
nand U2985 (N_2985,N_2848,N_2886);
or U2986 (N_2986,N_2868,N_2886);
and U2987 (N_2987,N_2828,N_2877);
nor U2988 (N_2988,N_2814,N_2879);
and U2989 (N_2989,N_2880,N_2808);
and U2990 (N_2990,N_2856,N_2803);
and U2991 (N_2991,N_2824,N_2834);
nor U2992 (N_2992,N_2817,N_2809);
xor U2993 (N_2993,N_2871,N_2863);
or U2994 (N_2994,N_2855,N_2859);
or U2995 (N_2995,N_2881,N_2847);
and U2996 (N_2996,N_2855,N_2834);
nor U2997 (N_2997,N_2810,N_2870);
and U2998 (N_2998,N_2849,N_2821);
nand U2999 (N_2999,N_2805,N_2851);
and U3000 (N_3000,N_2912,N_2905);
nand U3001 (N_3001,N_2967,N_2970);
or U3002 (N_3002,N_2983,N_2925);
nand U3003 (N_3003,N_2942,N_2987);
nor U3004 (N_3004,N_2930,N_2989);
nand U3005 (N_3005,N_2922,N_2933);
nor U3006 (N_3006,N_2962,N_2928);
nand U3007 (N_3007,N_2906,N_2993);
and U3008 (N_3008,N_2901,N_2958);
or U3009 (N_3009,N_2900,N_2924);
and U3010 (N_3010,N_2915,N_2941);
and U3011 (N_3011,N_2994,N_2953);
or U3012 (N_3012,N_2917,N_2982);
nor U3013 (N_3013,N_2923,N_2939);
nand U3014 (N_3014,N_2964,N_2975);
or U3015 (N_3015,N_2911,N_2954);
nor U3016 (N_3016,N_2921,N_2995);
nand U3017 (N_3017,N_2974,N_2966);
and U3018 (N_3018,N_2937,N_2984);
or U3019 (N_3019,N_2902,N_2968);
nand U3020 (N_3020,N_2957,N_2944);
nand U3021 (N_3021,N_2961,N_2997);
nor U3022 (N_3022,N_2955,N_2907);
nand U3023 (N_3023,N_2980,N_2959);
and U3024 (N_3024,N_2965,N_2913);
nor U3025 (N_3025,N_2992,N_2914);
nand U3026 (N_3026,N_2998,N_2935);
and U3027 (N_3027,N_2952,N_2963);
nand U3028 (N_3028,N_2910,N_2948);
or U3029 (N_3029,N_2929,N_2971);
nor U3030 (N_3030,N_2931,N_2903);
xor U3031 (N_3031,N_2976,N_2950);
or U3032 (N_3032,N_2978,N_2909);
and U3033 (N_3033,N_2936,N_2926);
nand U3034 (N_3034,N_2990,N_2945);
or U3035 (N_3035,N_2949,N_2977);
xnor U3036 (N_3036,N_2985,N_2940);
nand U3037 (N_3037,N_2951,N_2934);
nand U3038 (N_3038,N_2988,N_2999);
nand U3039 (N_3039,N_2981,N_2916);
nor U3040 (N_3040,N_2938,N_2986);
nor U3041 (N_3041,N_2996,N_2947);
and U3042 (N_3042,N_2946,N_2908);
nor U3043 (N_3043,N_2956,N_2919);
nand U3044 (N_3044,N_2927,N_2943);
xor U3045 (N_3045,N_2932,N_2979);
and U3046 (N_3046,N_2991,N_2920);
nand U3047 (N_3047,N_2972,N_2904);
or U3048 (N_3048,N_2918,N_2960);
and U3049 (N_3049,N_2969,N_2973);
and U3050 (N_3050,N_2973,N_2923);
nand U3051 (N_3051,N_2902,N_2962);
or U3052 (N_3052,N_2907,N_2990);
nor U3053 (N_3053,N_2978,N_2904);
nor U3054 (N_3054,N_2939,N_2929);
nand U3055 (N_3055,N_2910,N_2972);
nand U3056 (N_3056,N_2951,N_2960);
nor U3057 (N_3057,N_2969,N_2959);
and U3058 (N_3058,N_2944,N_2940);
and U3059 (N_3059,N_2924,N_2915);
nand U3060 (N_3060,N_2990,N_2989);
or U3061 (N_3061,N_2948,N_2955);
or U3062 (N_3062,N_2998,N_2907);
and U3063 (N_3063,N_2985,N_2935);
or U3064 (N_3064,N_2926,N_2909);
and U3065 (N_3065,N_2917,N_2915);
and U3066 (N_3066,N_2935,N_2926);
and U3067 (N_3067,N_2968,N_2986);
nand U3068 (N_3068,N_2957,N_2960);
nand U3069 (N_3069,N_2907,N_2952);
nor U3070 (N_3070,N_2974,N_2944);
nand U3071 (N_3071,N_2975,N_2990);
nor U3072 (N_3072,N_2943,N_2963);
nand U3073 (N_3073,N_2952,N_2918);
and U3074 (N_3074,N_2947,N_2953);
and U3075 (N_3075,N_2956,N_2915);
nor U3076 (N_3076,N_2991,N_2960);
nand U3077 (N_3077,N_2911,N_2930);
nor U3078 (N_3078,N_2946,N_2923);
nor U3079 (N_3079,N_2922,N_2911);
nand U3080 (N_3080,N_2924,N_2941);
nor U3081 (N_3081,N_2968,N_2964);
or U3082 (N_3082,N_2956,N_2941);
nor U3083 (N_3083,N_2968,N_2965);
or U3084 (N_3084,N_2921,N_2934);
nand U3085 (N_3085,N_2948,N_2951);
and U3086 (N_3086,N_2965,N_2953);
nor U3087 (N_3087,N_2908,N_2961);
or U3088 (N_3088,N_2943,N_2978);
or U3089 (N_3089,N_2955,N_2995);
and U3090 (N_3090,N_2972,N_2995);
nor U3091 (N_3091,N_2977,N_2969);
or U3092 (N_3092,N_2938,N_2905);
and U3093 (N_3093,N_2918,N_2961);
or U3094 (N_3094,N_2910,N_2944);
or U3095 (N_3095,N_2945,N_2937);
or U3096 (N_3096,N_2994,N_2990);
or U3097 (N_3097,N_2914,N_2985);
and U3098 (N_3098,N_2993,N_2917);
or U3099 (N_3099,N_2995,N_2905);
nand U3100 (N_3100,N_3022,N_3099);
xnor U3101 (N_3101,N_3064,N_3066);
nand U3102 (N_3102,N_3015,N_3039);
xnor U3103 (N_3103,N_3044,N_3025);
or U3104 (N_3104,N_3002,N_3092);
nor U3105 (N_3105,N_3021,N_3003);
or U3106 (N_3106,N_3074,N_3070);
and U3107 (N_3107,N_3035,N_3068);
or U3108 (N_3108,N_3071,N_3030);
nand U3109 (N_3109,N_3041,N_3065);
nand U3110 (N_3110,N_3079,N_3058);
or U3111 (N_3111,N_3050,N_3098);
or U3112 (N_3112,N_3094,N_3009);
and U3113 (N_3113,N_3036,N_3052);
or U3114 (N_3114,N_3073,N_3067);
nand U3115 (N_3115,N_3096,N_3043);
and U3116 (N_3116,N_3091,N_3017);
xnor U3117 (N_3117,N_3000,N_3087);
nand U3118 (N_3118,N_3088,N_3019);
nor U3119 (N_3119,N_3006,N_3059);
or U3120 (N_3120,N_3080,N_3047);
nor U3121 (N_3121,N_3063,N_3014);
nand U3122 (N_3122,N_3008,N_3028);
or U3123 (N_3123,N_3013,N_3054);
or U3124 (N_3124,N_3027,N_3057);
nand U3125 (N_3125,N_3016,N_3075);
nor U3126 (N_3126,N_3062,N_3010);
nand U3127 (N_3127,N_3020,N_3093);
and U3128 (N_3128,N_3084,N_3069);
and U3129 (N_3129,N_3097,N_3023);
nand U3130 (N_3130,N_3082,N_3034);
nand U3131 (N_3131,N_3032,N_3033);
or U3132 (N_3132,N_3031,N_3060);
and U3133 (N_3133,N_3037,N_3053);
nor U3134 (N_3134,N_3077,N_3042);
nor U3135 (N_3135,N_3011,N_3083);
or U3136 (N_3136,N_3026,N_3051);
and U3137 (N_3137,N_3086,N_3045);
and U3138 (N_3138,N_3055,N_3095);
and U3139 (N_3139,N_3018,N_3001);
nor U3140 (N_3140,N_3040,N_3005);
and U3141 (N_3141,N_3090,N_3076);
nand U3142 (N_3142,N_3046,N_3078);
and U3143 (N_3143,N_3072,N_3056);
or U3144 (N_3144,N_3081,N_3029);
nand U3145 (N_3145,N_3012,N_3089);
nand U3146 (N_3146,N_3061,N_3085);
or U3147 (N_3147,N_3024,N_3038);
or U3148 (N_3148,N_3048,N_3007);
nor U3149 (N_3149,N_3049,N_3004);
and U3150 (N_3150,N_3053,N_3040);
nor U3151 (N_3151,N_3055,N_3042);
nand U3152 (N_3152,N_3027,N_3040);
or U3153 (N_3153,N_3082,N_3055);
nand U3154 (N_3154,N_3032,N_3079);
and U3155 (N_3155,N_3096,N_3058);
and U3156 (N_3156,N_3015,N_3037);
xnor U3157 (N_3157,N_3083,N_3045);
nor U3158 (N_3158,N_3003,N_3042);
nand U3159 (N_3159,N_3067,N_3095);
nand U3160 (N_3160,N_3060,N_3028);
nor U3161 (N_3161,N_3023,N_3062);
or U3162 (N_3162,N_3030,N_3057);
nor U3163 (N_3163,N_3003,N_3024);
and U3164 (N_3164,N_3032,N_3048);
or U3165 (N_3165,N_3069,N_3020);
nand U3166 (N_3166,N_3054,N_3081);
or U3167 (N_3167,N_3038,N_3096);
and U3168 (N_3168,N_3013,N_3003);
nor U3169 (N_3169,N_3041,N_3071);
nor U3170 (N_3170,N_3093,N_3045);
and U3171 (N_3171,N_3083,N_3056);
and U3172 (N_3172,N_3034,N_3072);
nand U3173 (N_3173,N_3064,N_3081);
or U3174 (N_3174,N_3026,N_3099);
or U3175 (N_3175,N_3055,N_3070);
xnor U3176 (N_3176,N_3081,N_3086);
or U3177 (N_3177,N_3097,N_3086);
nand U3178 (N_3178,N_3058,N_3052);
or U3179 (N_3179,N_3054,N_3089);
xnor U3180 (N_3180,N_3073,N_3027);
nand U3181 (N_3181,N_3001,N_3077);
or U3182 (N_3182,N_3070,N_3024);
or U3183 (N_3183,N_3045,N_3008);
nor U3184 (N_3184,N_3081,N_3090);
nor U3185 (N_3185,N_3041,N_3045);
nor U3186 (N_3186,N_3006,N_3045);
and U3187 (N_3187,N_3025,N_3008);
nand U3188 (N_3188,N_3000,N_3025);
and U3189 (N_3189,N_3059,N_3044);
or U3190 (N_3190,N_3091,N_3035);
and U3191 (N_3191,N_3003,N_3014);
and U3192 (N_3192,N_3014,N_3054);
nand U3193 (N_3193,N_3029,N_3078);
or U3194 (N_3194,N_3067,N_3069);
nand U3195 (N_3195,N_3033,N_3056);
and U3196 (N_3196,N_3035,N_3095);
or U3197 (N_3197,N_3068,N_3022);
and U3198 (N_3198,N_3020,N_3074);
nand U3199 (N_3199,N_3092,N_3050);
nand U3200 (N_3200,N_3139,N_3149);
and U3201 (N_3201,N_3135,N_3178);
or U3202 (N_3202,N_3114,N_3147);
and U3203 (N_3203,N_3143,N_3140);
and U3204 (N_3204,N_3126,N_3116);
nor U3205 (N_3205,N_3105,N_3101);
nand U3206 (N_3206,N_3193,N_3127);
nand U3207 (N_3207,N_3167,N_3190);
or U3208 (N_3208,N_3179,N_3118);
or U3209 (N_3209,N_3115,N_3123);
nand U3210 (N_3210,N_3148,N_3177);
or U3211 (N_3211,N_3121,N_3157);
nand U3212 (N_3212,N_3187,N_3119);
or U3213 (N_3213,N_3181,N_3124);
or U3214 (N_3214,N_3122,N_3166);
and U3215 (N_3215,N_3163,N_3182);
nor U3216 (N_3216,N_3175,N_3112);
nand U3217 (N_3217,N_3154,N_3168);
nor U3218 (N_3218,N_3192,N_3189);
nand U3219 (N_3219,N_3111,N_3131);
or U3220 (N_3220,N_3134,N_3165);
nor U3221 (N_3221,N_3174,N_3155);
nand U3222 (N_3222,N_3194,N_3162);
nand U3223 (N_3223,N_3150,N_3160);
or U3224 (N_3224,N_3146,N_3152);
xor U3225 (N_3225,N_3142,N_3137);
nor U3226 (N_3226,N_3185,N_3113);
nor U3227 (N_3227,N_3129,N_3156);
and U3228 (N_3228,N_3107,N_3159);
and U3229 (N_3229,N_3169,N_3144);
or U3230 (N_3230,N_3186,N_3153);
or U3231 (N_3231,N_3102,N_3100);
nand U3232 (N_3232,N_3138,N_3128);
nand U3233 (N_3233,N_3188,N_3180);
nand U3234 (N_3234,N_3106,N_3151);
and U3235 (N_3235,N_3164,N_3172);
or U3236 (N_3236,N_3108,N_3161);
nor U3237 (N_3237,N_3145,N_3170);
and U3238 (N_3238,N_3191,N_3199);
nand U3239 (N_3239,N_3120,N_3171);
and U3240 (N_3240,N_3196,N_3158);
nand U3241 (N_3241,N_3141,N_3110);
or U3242 (N_3242,N_3103,N_3197);
nand U3243 (N_3243,N_3125,N_3176);
nand U3244 (N_3244,N_3198,N_3173);
or U3245 (N_3245,N_3133,N_3109);
and U3246 (N_3246,N_3183,N_3184);
and U3247 (N_3247,N_3195,N_3130);
and U3248 (N_3248,N_3117,N_3136);
nand U3249 (N_3249,N_3132,N_3104);
or U3250 (N_3250,N_3128,N_3168);
nor U3251 (N_3251,N_3178,N_3191);
nor U3252 (N_3252,N_3105,N_3117);
or U3253 (N_3253,N_3101,N_3145);
nor U3254 (N_3254,N_3164,N_3142);
or U3255 (N_3255,N_3119,N_3114);
nor U3256 (N_3256,N_3157,N_3193);
nor U3257 (N_3257,N_3103,N_3183);
or U3258 (N_3258,N_3179,N_3195);
and U3259 (N_3259,N_3126,N_3112);
nand U3260 (N_3260,N_3126,N_3136);
and U3261 (N_3261,N_3150,N_3168);
and U3262 (N_3262,N_3109,N_3142);
nand U3263 (N_3263,N_3108,N_3127);
and U3264 (N_3264,N_3173,N_3113);
nand U3265 (N_3265,N_3187,N_3179);
and U3266 (N_3266,N_3127,N_3155);
and U3267 (N_3267,N_3147,N_3117);
or U3268 (N_3268,N_3103,N_3101);
nand U3269 (N_3269,N_3178,N_3138);
nand U3270 (N_3270,N_3164,N_3174);
nor U3271 (N_3271,N_3176,N_3196);
or U3272 (N_3272,N_3141,N_3114);
nor U3273 (N_3273,N_3173,N_3106);
nor U3274 (N_3274,N_3178,N_3158);
nand U3275 (N_3275,N_3182,N_3120);
and U3276 (N_3276,N_3104,N_3101);
or U3277 (N_3277,N_3165,N_3189);
nor U3278 (N_3278,N_3101,N_3131);
nand U3279 (N_3279,N_3192,N_3168);
or U3280 (N_3280,N_3110,N_3191);
nand U3281 (N_3281,N_3119,N_3172);
or U3282 (N_3282,N_3179,N_3142);
nor U3283 (N_3283,N_3104,N_3105);
nand U3284 (N_3284,N_3144,N_3177);
and U3285 (N_3285,N_3180,N_3187);
nor U3286 (N_3286,N_3105,N_3168);
nand U3287 (N_3287,N_3152,N_3130);
nand U3288 (N_3288,N_3136,N_3190);
and U3289 (N_3289,N_3144,N_3165);
nand U3290 (N_3290,N_3188,N_3178);
and U3291 (N_3291,N_3166,N_3135);
xnor U3292 (N_3292,N_3179,N_3103);
and U3293 (N_3293,N_3131,N_3124);
or U3294 (N_3294,N_3146,N_3160);
xor U3295 (N_3295,N_3169,N_3148);
nor U3296 (N_3296,N_3180,N_3189);
or U3297 (N_3297,N_3103,N_3188);
nand U3298 (N_3298,N_3191,N_3100);
nor U3299 (N_3299,N_3125,N_3159);
nor U3300 (N_3300,N_3283,N_3258);
nor U3301 (N_3301,N_3275,N_3291);
nand U3302 (N_3302,N_3210,N_3299);
or U3303 (N_3303,N_3220,N_3268);
nor U3304 (N_3304,N_3239,N_3229);
nand U3305 (N_3305,N_3213,N_3250);
or U3306 (N_3306,N_3221,N_3256);
or U3307 (N_3307,N_3204,N_3251);
and U3308 (N_3308,N_3223,N_3224);
nor U3309 (N_3309,N_3203,N_3267);
nor U3310 (N_3310,N_3284,N_3245);
nand U3311 (N_3311,N_3214,N_3294);
nor U3312 (N_3312,N_3247,N_3272);
and U3313 (N_3313,N_3263,N_3222);
or U3314 (N_3314,N_3237,N_3248);
or U3315 (N_3315,N_3232,N_3254);
nand U3316 (N_3316,N_3255,N_3234);
or U3317 (N_3317,N_3226,N_3262);
or U3318 (N_3318,N_3297,N_3277);
and U3319 (N_3319,N_3273,N_3261);
nand U3320 (N_3320,N_3270,N_3238);
and U3321 (N_3321,N_3208,N_3227);
nor U3322 (N_3322,N_3292,N_3233);
or U3323 (N_3323,N_3231,N_3280);
nor U3324 (N_3324,N_3235,N_3217);
or U3325 (N_3325,N_3271,N_3200);
nand U3326 (N_3326,N_3253,N_3274);
or U3327 (N_3327,N_3240,N_3230);
and U3328 (N_3328,N_3228,N_3285);
and U3329 (N_3329,N_3282,N_3241);
or U3330 (N_3330,N_3225,N_3246);
nand U3331 (N_3331,N_3236,N_3259);
and U3332 (N_3332,N_3281,N_3278);
nand U3333 (N_3333,N_3201,N_3289);
nor U3334 (N_3334,N_3269,N_3212);
and U3335 (N_3335,N_3252,N_3287);
and U3336 (N_3336,N_3216,N_3205);
nor U3337 (N_3337,N_3266,N_3215);
nand U3338 (N_3338,N_3249,N_3296);
or U3339 (N_3339,N_3265,N_3209);
or U3340 (N_3340,N_3244,N_3290);
and U3341 (N_3341,N_3279,N_3257);
and U3342 (N_3342,N_3264,N_3202);
nand U3343 (N_3343,N_3207,N_3242);
and U3344 (N_3344,N_3298,N_3293);
and U3345 (N_3345,N_3276,N_3243);
nor U3346 (N_3346,N_3219,N_3218);
nor U3347 (N_3347,N_3295,N_3286);
nor U3348 (N_3348,N_3211,N_3260);
nor U3349 (N_3349,N_3288,N_3206);
and U3350 (N_3350,N_3291,N_3221);
or U3351 (N_3351,N_3224,N_3211);
nor U3352 (N_3352,N_3213,N_3297);
and U3353 (N_3353,N_3219,N_3202);
nand U3354 (N_3354,N_3219,N_3293);
nor U3355 (N_3355,N_3238,N_3261);
nor U3356 (N_3356,N_3255,N_3281);
nand U3357 (N_3357,N_3248,N_3265);
nand U3358 (N_3358,N_3295,N_3204);
or U3359 (N_3359,N_3200,N_3243);
nor U3360 (N_3360,N_3205,N_3246);
nor U3361 (N_3361,N_3248,N_3291);
nand U3362 (N_3362,N_3269,N_3297);
nor U3363 (N_3363,N_3298,N_3252);
nor U3364 (N_3364,N_3295,N_3210);
nor U3365 (N_3365,N_3208,N_3297);
nor U3366 (N_3366,N_3227,N_3285);
and U3367 (N_3367,N_3232,N_3200);
nand U3368 (N_3368,N_3245,N_3242);
nand U3369 (N_3369,N_3266,N_3256);
nor U3370 (N_3370,N_3280,N_3263);
or U3371 (N_3371,N_3212,N_3286);
nand U3372 (N_3372,N_3242,N_3260);
and U3373 (N_3373,N_3240,N_3206);
and U3374 (N_3374,N_3227,N_3271);
or U3375 (N_3375,N_3299,N_3267);
and U3376 (N_3376,N_3220,N_3236);
or U3377 (N_3377,N_3237,N_3277);
nor U3378 (N_3378,N_3249,N_3270);
and U3379 (N_3379,N_3270,N_3281);
or U3380 (N_3380,N_3236,N_3242);
or U3381 (N_3381,N_3295,N_3203);
and U3382 (N_3382,N_3281,N_3266);
nor U3383 (N_3383,N_3246,N_3252);
nand U3384 (N_3384,N_3276,N_3279);
or U3385 (N_3385,N_3227,N_3269);
nand U3386 (N_3386,N_3259,N_3221);
or U3387 (N_3387,N_3299,N_3238);
or U3388 (N_3388,N_3226,N_3281);
nand U3389 (N_3389,N_3224,N_3299);
or U3390 (N_3390,N_3278,N_3227);
nor U3391 (N_3391,N_3221,N_3237);
nand U3392 (N_3392,N_3266,N_3283);
and U3393 (N_3393,N_3267,N_3258);
and U3394 (N_3394,N_3247,N_3218);
nor U3395 (N_3395,N_3293,N_3241);
or U3396 (N_3396,N_3243,N_3273);
or U3397 (N_3397,N_3249,N_3204);
or U3398 (N_3398,N_3207,N_3214);
or U3399 (N_3399,N_3246,N_3227);
nand U3400 (N_3400,N_3371,N_3305);
and U3401 (N_3401,N_3330,N_3300);
nand U3402 (N_3402,N_3393,N_3394);
or U3403 (N_3403,N_3398,N_3307);
nor U3404 (N_3404,N_3389,N_3347);
nor U3405 (N_3405,N_3359,N_3324);
xnor U3406 (N_3406,N_3362,N_3391);
nor U3407 (N_3407,N_3322,N_3318);
and U3408 (N_3408,N_3319,N_3352);
or U3409 (N_3409,N_3327,N_3355);
nor U3410 (N_3410,N_3311,N_3378);
nor U3411 (N_3411,N_3383,N_3396);
or U3412 (N_3412,N_3360,N_3346);
nor U3413 (N_3413,N_3341,N_3345);
nor U3414 (N_3414,N_3316,N_3310);
nand U3415 (N_3415,N_3301,N_3302);
nor U3416 (N_3416,N_3313,N_3353);
nand U3417 (N_3417,N_3397,N_3368);
or U3418 (N_3418,N_3376,N_3337);
or U3419 (N_3419,N_3384,N_3356);
nor U3420 (N_3420,N_3370,N_3367);
and U3421 (N_3421,N_3375,N_3329);
nand U3422 (N_3422,N_3320,N_3335);
nand U3423 (N_3423,N_3344,N_3385);
and U3424 (N_3424,N_3365,N_3323);
nor U3425 (N_3425,N_3336,N_3306);
or U3426 (N_3426,N_3340,N_3342);
xnor U3427 (N_3427,N_3374,N_3373);
xnor U3428 (N_3428,N_3326,N_3338);
nor U3429 (N_3429,N_3332,N_3382);
nor U3430 (N_3430,N_3357,N_3304);
or U3431 (N_3431,N_3364,N_3379);
or U3432 (N_3432,N_3387,N_3339);
nor U3433 (N_3433,N_3315,N_3361);
nand U3434 (N_3434,N_3363,N_3314);
nor U3435 (N_3435,N_3333,N_3308);
and U3436 (N_3436,N_3349,N_3348);
and U3437 (N_3437,N_3388,N_3366);
and U3438 (N_3438,N_3372,N_3312);
and U3439 (N_3439,N_3386,N_3321);
or U3440 (N_3440,N_3380,N_3334);
nand U3441 (N_3441,N_3351,N_3395);
nor U3442 (N_3442,N_3369,N_3390);
or U3443 (N_3443,N_3358,N_3392);
nor U3444 (N_3444,N_3377,N_3399);
and U3445 (N_3445,N_3317,N_3354);
and U3446 (N_3446,N_3343,N_3303);
xnor U3447 (N_3447,N_3309,N_3350);
nand U3448 (N_3448,N_3328,N_3325);
nand U3449 (N_3449,N_3381,N_3331);
and U3450 (N_3450,N_3338,N_3306);
and U3451 (N_3451,N_3349,N_3386);
or U3452 (N_3452,N_3364,N_3333);
nor U3453 (N_3453,N_3375,N_3361);
and U3454 (N_3454,N_3338,N_3318);
nand U3455 (N_3455,N_3362,N_3346);
or U3456 (N_3456,N_3384,N_3367);
nand U3457 (N_3457,N_3319,N_3316);
and U3458 (N_3458,N_3348,N_3366);
and U3459 (N_3459,N_3316,N_3357);
or U3460 (N_3460,N_3317,N_3384);
or U3461 (N_3461,N_3380,N_3340);
and U3462 (N_3462,N_3391,N_3333);
and U3463 (N_3463,N_3305,N_3342);
nand U3464 (N_3464,N_3346,N_3340);
nand U3465 (N_3465,N_3354,N_3337);
or U3466 (N_3466,N_3377,N_3302);
or U3467 (N_3467,N_3371,N_3359);
or U3468 (N_3468,N_3331,N_3384);
nand U3469 (N_3469,N_3368,N_3395);
nand U3470 (N_3470,N_3313,N_3367);
or U3471 (N_3471,N_3386,N_3309);
or U3472 (N_3472,N_3329,N_3300);
nor U3473 (N_3473,N_3337,N_3335);
nand U3474 (N_3474,N_3378,N_3321);
or U3475 (N_3475,N_3310,N_3335);
or U3476 (N_3476,N_3357,N_3354);
nor U3477 (N_3477,N_3317,N_3339);
and U3478 (N_3478,N_3371,N_3335);
and U3479 (N_3479,N_3383,N_3323);
nor U3480 (N_3480,N_3361,N_3388);
nand U3481 (N_3481,N_3385,N_3319);
nor U3482 (N_3482,N_3310,N_3386);
nand U3483 (N_3483,N_3348,N_3323);
and U3484 (N_3484,N_3389,N_3378);
nor U3485 (N_3485,N_3340,N_3357);
xnor U3486 (N_3486,N_3321,N_3344);
and U3487 (N_3487,N_3327,N_3309);
nor U3488 (N_3488,N_3377,N_3328);
nor U3489 (N_3489,N_3323,N_3349);
and U3490 (N_3490,N_3341,N_3377);
or U3491 (N_3491,N_3368,N_3380);
and U3492 (N_3492,N_3346,N_3359);
nor U3493 (N_3493,N_3338,N_3369);
and U3494 (N_3494,N_3346,N_3336);
nand U3495 (N_3495,N_3325,N_3371);
or U3496 (N_3496,N_3323,N_3381);
or U3497 (N_3497,N_3396,N_3317);
nor U3498 (N_3498,N_3334,N_3348);
or U3499 (N_3499,N_3389,N_3381);
and U3500 (N_3500,N_3448,N_3453);
nor U3501 (N_3501,N_3482,N_3458);
nor U3502 (N_3502,N_3480,N_3470);
or U3503 (N_3503,N_3429,N_3431);
or U3504 (N_3504,N_3493,N_3463);
or U3505 (N_3505,N_3414,N_3464);
and U3506 (N_3506,N_3485,N_3495);
nand U3507 (N_3507,N_3428,N_3455);
or U3508 (N_3508,N_3457,N_3424);
and U3509 (N_3509,N_3408,N_3417);
nor U3510 (N_3510,N_3427,N_3450);
and U3511 (N_3511,N_3479,N_3456);
nand U3512 (N_3512,N_3487,N_3468);
and U3513 (N_3513,N_3467,N_3425);
or U3514 (N_3514,N_3401,N_3440);
and U3515 (N_3515,N_3484,N_3496);
or U3516 (N_3516,N_3486,N_3462);
and U3517 (N_3517,N_3413,N_3412);
and U3518 (N_3518,N_3445,N_3419);
nor U3519 (N_3519,N_3476,N_3441);
nor U3520 (N_3520,N_3451,N_3471);
or U3521 (N_3521,N_3426,N_3400);
and U3522 (N_3522,N_3406,N_3472);
nand U3523 (N_3523,N_3442,N_3474);
nand U3524 (N_3524,N_3415,N_3443);
nand U3525 (N_3525,N_3483,N_3421);
nand U3526 (N_3526,N_3465,N_3498);
and U3527 (N_3527,N_3490,N_3488);
nand U3528 (N_3528,N_3418,N_3407);
nor U3529 (N_3529,N_3432,N_3435);
nand U3530 (N_3530,N_3404,N_3447);
nor U3531 (N_3531,N_3409,N_3439);
or U3532 (N_3532,N_3436,N_3449);
nor U3533 (N_3533,N_3405,N_3434);
or U3534 (N_3534,N_3423,N_3475);
nor U3535 (N_3535,N_3489,N_3491);
nor U3536 (N_3536,N_3420,N_3430);
or U3537 (N_3537,N_3469,N_3494);
or U3538 (N_3538,N_3416,N_3466);
or U3539 (N_3539,N_3452,N_3492);
and U3540 (N_3540,N_3497,N_3477);
nand U3541 (N_3541,N_3473,N_3403);
nand U3542 (N_3542,N_3481,N_3478);
nand U3543 (N_3543,N_3438,N_3454);
nor U3544 (N_3544,N_3444,N_3460);
and U3545 (N_3545,N_3422,N_3411);
nor U3546 (N_3546,N_3433,N_3499);
and U3547 (N_3547,N_3461,N_3459);
nor U3548 (N_3548,N_3437,N_3410);
nand U3549 (N_3549,N_3446,N_3402);
nor U3550 (N_3550,N_3425,N_3488);
nand U3551 (N_3551,N_3490,N_3420);
nor U3552 (N_3552,N_3460,N_3457);
nor U3553 (N_3553,N_3484,N_3495);
nor U3554 (N_3554,N_3474,N_3482);
or U3555 (N_3555,N_3408,N_3429);
nand U3556 (N_3556,N_3446,N_3440);
nor U3557 (N_3557,N_3459,N_3487);
nor U3558 (N_3558,N_3427,N_3446);
or U3559 (N_3559,N_3434,N_3467);
nand U3560 (N_3560,N_3486,N_3422);
nor U3561 (N_3561,N_3432,N_3434);
nand U3562 (N_3562,N_3428,N_3454);
and U3563 (N_3563,N_3485,N_3453);
nor U3564 (N_3564,N_3487,N_3485);
nor U3565 (N_3565,N_3434,N_3400);
nor U3566 (N_3566,N_3451,N_3443);
nor U3567 (N_3567,N_3423,N_3460);
nor U3568 (N_3568,N_3413,N_3443);
nor U3569 (N_3569,N_3489,N_3416);
nor U3570 (N_3570,N_3442,N_3409);
or U3571 (N_3571,N_3487,N_3450);
nor U3572 (N_3572,N_3464,N_3473);
nand U3573 (N_3573,N_3485,N_3407);
nor U3574 (N_3574,N_3407,N_3409);
and U3575 (N_3575,N_3466,N_3483);
and U3576 (N_3576,N_3463,N_3484);
nor U3577 (N_3577,N_3488,N_3437);
nand U3578 (N_3578,N_3410,N_3490);
or U3579 (N_3579,N_3495,N_3458);
or U3580 (N_3580,N_3436,N_3419);
nand U3581 (N_3581,N_3492,N_3475);
and U3582 (N_3582,N_3467,N_3429);
nor U3583 (N_3583,N_3421,N_3462);
nor U3584 (N_3584,N_3461,N_3492);
nand U3585 (N_3585,N_3475,N_3443);
nand U3586 (N_3586,N_3457,N_3422);
nor U3587 (N_3587,N_3402,N_3468);
and U3588 (N_3588,N_3494,N_3451);
nand U3589 (N_3589,N_3410,N_3419);
or U3590 (N_3590,N_3479,N_3448);
nor U3591 (N_3591,N_3408,N_3464);
and U3592 (N_3592,N_3453,N_3402);
nor U3593 (N_3593,N_3401,N_3455);
nand U3594 (N_3594,N_3447,N_3498);
and U3595 (N_3595,N_3405,N_3448);
nand U3596 (N_3596,N_3494,N_3466);
nand U3597 (N_3597,N_3470,N_3411);
or U3598 (N_3598,N_3412,N_3441);
and U3599 (N_3599,N_3417,N_3492);
or U3600 (N_3600,N_3541,N_3509);
or U3601 (N_3601,N_3577,N_3597);
or U3602 (N_3602,N_3518,N_3501);
and U3603 (N_3603,N_3590,N_3513);
nor U3604 (N_3604,N_3503,N_3540);
or U3605 (N_3605,N_3538,N_3592);
and U3606 (N_3606,N_3578,N_3524);
nand U3607 (N_3607,N_3552,N_3507);
nand U3608 (N_3608,N_3564,N_3531);
and U3609 (N_3609,N_3566,N_3594);
nand U3610 (N_3610,N_3582,N_3534);
or U3611 (N_3611,N_3567,N_3551);
nor U3612 (N_3612,N_3520,N_3599);
nor U3613 (N_3613,N_3543,N_3537);
nor U3614 (N_3614,N_3533,N_3526);
nor U3615 (N_3615,N_3598,N_3562);
or U3616 (N_3616,N_3559,N_3593);
and U3617 (N_3617,N_3587,N_3547);
and U3618 (N_3618,N_3536,N_3502);
nor U3619 (N_3619,N_3523,N_3532);
nor U3620 (N_3620,N_3546,N_3585);
xnor U3621 (N_3621,N_3595,N_3514);
nand U3622 (N_3622,N_3572,N_3563);
and U3623 (N_3623,N_3511,N_3504);
or U3624 (N_3624,N_3516,N_3557);
nor U3625 (N_3625,N_3568,N_3542);
nor U3626 (N_3626,N_3576,N_3522);
or U3627 (N_3627,N_3589,N_3556);
and U3628 (N_3628,N_3508,N_3580);
nand U3629 (N_3629,N_3570,N_3548);
or U3630 (N_3630,N_3530,N_3545);
or U3631 (N_3631,N_3591,N_3553);
nor U3632 (N_3632,N_3517,N_3588);
nand U3633 (N_3633,N_3573,N_3505);
or U3634 (N_3634,N_3519,N_3500);
nand U3635 (N_3635,N_3544,N_3506);
nor U3636 (N_3636,N_3569,N_3575);
xor U3637 (N_3637,N_3528,N_3574);
or U3638 (N_3638,N_3581,N_3558);
and U3639 (N_3639,N_3560,N_3521);
or U3640 (N_3640,N_3596,N_3565);
and U3641 (N_3641,N_3549,N_3554);
and U3642 (N_3642,N_3579,N_3586);
nand U3643 (N_3643,N_3561,N_3535);
and U3644 (N_3644,N_3525,N_3515);
or U3645 (N_3645,N_3527,N_3529);
or U3646 (N_3646,N_3539,N_3571);
nand U3647 (N_3647,N_3550,N_3512);
and U3648 (N_3648,N_3583,N_3555);
nand U3649 (N_3649,N_3584,N_3510);
or U3650 (N_3650,N_3564,N_3570);
and U3651 (N_3651,N_3572,N_3584);
nand U3652 (N_3652,N_3533,N_3542);
nand U3653 (N_3653,N_3587,N_3581);
nor U3654 (N_3654,N_3576,N_3567);
or U3655 (N_3655,N_3568,N_3510);
or U3656 (N_3656,N_3575,N_3591);
or U3657 (N_3657,N_3598,N_3559);
nor U3658 (N_3658,N_3522,N_3566);
nor U3659 (N_3659,N_3574,N_3535);
or U3660 (N_3660,N_3536,N_3576);
or U3661 (N_3661,N_3522,N_3581);
xor U3662 (N_3662,N_3558,N_3527);
and U3663 (N_3663,N_3554,N_3552);
nor U3664 (N_3664,N_3519,N_3518);
and U3665 (N_3665,N_3507,N_3544);
nor U3666 (N_3666,N_3587,N_3522);
or U3667 (N_3667,N_3590,N_3582);
or U3668 (N_3668,N_3527,N_3518);
nand U3669 (N_3669,N_3570,N_3559);
nand U3670 (N_3670,N_3535,N_3573);
or U3671 (N_3671,N_3590,N_3525);
or U3672 (N_3672,N_3578,N_3566);
nand U3673 (N_3673,N_3535,N_3572);
nand U3674 (N_3674,N_3513,N_3561);
and U3675 (N_3675,N_3506,N_3562);
and U3676 (N_3676,N_3533,N_3520);
or U3677 (N_3677,N_3572,N_3523);
or U3678 (N_3678,N_3519,N_3508);
nor U3679 (N_3679,N_3515,N_3540);
and U3680 (N_3680,N_3595,N_3565);
nand U3681 (N_3681,N_3534,N_3597);
or U3682 (N_3682,N_3547,N_3572);
nor U3683 (N_3683,N_3590,N_3540);
nand U3684 (N_3684,N_3586,N_3533);
and U3685 (N_3685,N_3555,N_3545);
and U3686 (N_3686,N_3504,N_3533);
nor U3687 (N_3687,N_3584,N_3544);
and U3688 (N_3688,N_3548,N_3564);
and U3689 (N_3689,N_3568,N_3563);
or U3690 (N_3690,N_3515,N_3508);
or U3691 (N_3691,N_3548,N_3505);
or U3692 (N_3692,N_3596,N_3559);
and U3693 (N_3693,N_3500,N_3570);
nor U3694 (N_3694,N_3552,N_3549);
and U3695 (N_3695,N_3558,N_3530);
and U3696 (N_3696,N_3550,N_3506);
nand U3697 (N_3697,N_3520,N_3572);
and U3698 (N_3698,N_3588,N_3537);
nand U3699 (N_3699,N_3591,N_3554);
nand U3700 (N_3700,N_3602,N_3693);
nor U3701 (N_3701,N_3649,N_3675);
xor U3702 (N_3702,N_3623,N_3603);
nor U3703 (N_3703,N_3629,N_3676);
and U3704 (N_3704,N_3685,N_3642);
nor U3705 (N_3705,N_3688,N_3660);
nand U3706 (N_3706,N_3671,N_3696);
or U3707 (N_3707,N_3614,N_3673);
or U3708 (N_3708,N_3665,N_3601);
nand U3709 (N_3709,N_3608,N_3641);
or U3710 (N_3710,N_3624,N_3638);
or U3711 (N_3711,N_3651,N_3692);
and U3712 (N_3712,N_3611,N_3618);
and U3713 (N_3713,N_3655,N_3643);
or U3714 (N_3714,N_3637,N_3644);
or U3715 (N_3715,N_3681,N_3636);
and U3716 (N_3716,N_3697,N_3625);
and U3717 (N_3717,N_3647,N_3633);
or U3718 (N_3718,N_3658,N_3699);
and U3719 (N_3719,N_3615,N_3659);
or U3720 (N_3720,N_3619,N_3683);
or U3721 (N_3721,N_3687,N_3656);
or U3722 (N_3722,N_3639,N_3664);
nor U3723 (N_3723,N_3600,N_3682);
and U3724 (N_3724,N_3621,N_3635);
and U3725 (N_3725,N_3630,N_3670);
nor U3726 (N_3726,N_3605,N_3640);
nor U3727 (N_3727,N_3652,N_3684);
nand U3728 (N_3728,N_3672,N_3694);
and U3729 (N_3729,N_3669,N_3654);
nand U3730 (N_3730,N_3607,N_3634);
nor U3731 (N_3731,N_3627,N_3691);
or U3732 (N_3732,N_3668,N_3690);
or U3733 (N_3733,N_3679,N_3622);
nor U3734 (N_3734,N_3689,N_3645);
nand U3735 (N_3735,N_3612,N_3613);
and U3736 (N_3736,N_3661,N_3663);
nand U3737 (N_3737,N_3626,N_3616);
nand U3738 (N_3738,N_3653,N_3610);
nor U3739 (N_3739,N_3609,N_3695);
and U3740 (N_3740,N_3617,N_3678);
nand U3741 (N_3741,N_3628,N_3662);
or U3742 (N_3742,N_3632,N_3666);
nand U3743 (N_3743,N_3698,N_3674);
nand U3744 (N_3744,N_3631,N_3646);
nand U3745 (N_3745,N_3667,N_3657);
or U3746 (N_3746,N_3606,N_3648);
nor U3747 (N_3747,N_3686,N_3677);
or U3748 (N_3748,N_3680,N_3604);
nor U3749 (N_3749,N_3650,N_3620);
nand U3750 (N_3750,N_3626,N_3607);
nand U3751 (N_3751,N_3693,N_3668);
nand U3752 (N_3752,N_3621,N_3617);
nor U3753 (N_3753,N_3683,N_3650);
and U3754 (N_3754,N_3652,N_3638);
nand U3755 (N_3755,N_3602,N_3624);
or U3756 (N_3756,N_3691,N_3637);
nand U3757 (N_3757,N_3638,N_3658);
nor U3758 (N_3758,N_3600,N_3602);
nor U3759 (N_3759,N_3614,N_3605);
nor U3760 (N_3760,N_3669,N_3670);
or U3761 (N_3761,N_3638,N_3683);
or U3762 (N_3762,N_3677,N_3674);
or U3763 (N_3763,N_3613,N_3610);
nand U3764 (N_3764,N_3606,N_3601);
and U3765 (N_3765,N_3643,N_3689);
nor U3766 (N_3766,N_3626,N_3611);
or U3767 (N_3767,N_3618,N_3683);
nand U3768 (N_3768,N_3663,N_3642);
nor U3769 (N_3769,N_3653,N_3678);
nor U3770 (N_3770,N_3674,N_3689);
and U3771 (N_3771,N_3608,N_3657);
or U3772 (N_3772,N_3618,N_3679);
nand U3773 (N_3773,N_3665,N_3643);
and U3774 (N_3774,N_3617,N_3600);
nand U3775 (N_3775,N_3661,N_3624);
nand U3776 (N_3776,N_3674,N_3675);
nand U3777 (N_3777,N_3670,N_3663);
nand U3778 (N_3778,N_3615,N_3683);
nand U3779 (N_3779,N_3634,N_3615);
nand U3780 (N_3780,N_3681,N_3655);
nand U3781 (N_3781,N_3677,N_3646);
nor U3782 (N_3782,N_3675,N_3641);
and U3783 (N_3783,N_3695,N_3621);
nand U3784 (N_3784,N_3647,N_3675);
or U3785 (N_3785,N_3624,N_3640);
xnor U3786 (N_3786,N_3694,N_3639);
or U3787 (N_3787,N_3610,N_3607);
or U3788 (N_3788,N_3640,N_3684);
nand U3789 (N_3789,N_3636,N_3677);
nand U3790 (N_3790,N_3640,N_3638);
and U3791 (N_3791,N_3612,N_3638);
or U3792 (N_3792,N_3670,N_3625);
or U3793 (N_3793,N_3669,N_3677);
nand U3794 (N_3794,N_3617,N_3685);
nand U3795 (N_3795,N_3632,N_3678);
and U3796 (N_3796,N_3617,N_3680);
or U3797 (N_3797,N_3623,N_3645);
and U3798 (N_3798,N_3635,N_3643);
or U3799 (N_3799,N_3650,N_3677);
or U3800 (N_3800,N_3705,N_3740);
nor U3801 (N_3801,N_3770,N_3747);
or U3802 (N_3802,N_3796,N_3783);
or U3803 (N_3803,N_3773,N_3780);
or U3804 (N_3804,N_3715,N_3721);
nor U3805 (N_3805,N_3711,N_3743);
nand U3806 (N_3806,N_3726,N_3703);
nand U3807 (N_3807,N_3720,N_3768);
or U3808 (N_3808,N_3708,N_3787);
nor U3809 (N_3809,N_3762,N_3707);
nand U3810 (N_3810,N_3792,N_3727);
nor U3811 (N_3811,N_3799,N_3746);
nand U3812 (N_3812,N_3774,N_3772);
xnor U3813 (N_3813,N_3785,N_3771);
or U3814 (N_3814,N_3712,N_3704);
and U3815 (N_3815,N_3791,N_3764);
nand U3816 (N_3816,N_3742,N_3753);
and U3817 (N_3817,N_3752,N_3744);
nand U3818 (N_3818,N_3793,N_3706);
and U3819 (N_3819,N_3700,N_3778);
nor U3820 (N_3820,N_3731,N_3710);
xnor U3821 (N_3821,N_3763,N_3790);
nor U3822 (N_3822,N_3737,N_3709);
or U3823 (N_3823,N_3769,N_3733);
and U3824 (N_3824,N_3748,N_3736);
or U3825 (N_3825,N_3776,N_3754);
and U3826 (N_3826,N_3716,N_3723);
nand U3827 (N_3827,N_3741,N_3789);
and U3828 (N_3828,N_3755,N_3781);
and U3829 (N_3829,N_3782,N_3725);
and U3830 (N_3830,N_3729,N_3775);
or U3831 (N_3831,N_3738,N_3797);
nand U3832 (N_3832,N_3761,N_3779);
or U3833 (N_3833,N_3794,N_3750);
xor U3834 (N_3834,N_3786,N_3722);
and U3835 (N_3835,N_3788,N_3735);
or U3836 (N_3836,N_3730,N_3795);
nand U3837 (N_3837,N_3767,N_3756);
or U3838 (N_3838,N_3732,N_3760);
xnor U3839 (N_3839,N_3713,N_3759);
nor U3840 (N_3840,N_3758,N_3749);
and U3841 (N_3841,N_3718,N_3739);
nor U3842 (N_3842,N_3784,N_3777);
or U3843 (N_3843,N_3757,N_3702);
nor U3844 (N_3844,N_3766,N_3701);
and U3845 (N_3845,N_3714,N_3745);
nor U3846 (N_3846,N_3717,N_3751);
xor U3847 (N_3847,N_3765,N_3798);
or U3848 (N_3848,N_3734,N_3724);
and U3849 (N_3849,N_3728,N_3719);
and U3850 (N_3850,N_3784,N_3756);
nor U3851 (N_3851,N_3705,N_3742);
and U3852 (N_3852,N_3771,N_3793);
xor U3853 (N_3853,N_3792,N_3769);
nand U3854 (N_3854,N_3750,N_3702);
or U3855 (N_3855,N_3722,N_3706);
nor U3856 (N_3856,N_3716,N_3746);
nor U3857 (N_3857,N_3777,N_3763);
nand U3858 (N_3858,N_3709,N_3792);
nor U3859 (N_3859,N_3747,N_3783);
nand U3860 (N_3860,N_3762,N_3726);
or U3861 (N_3861,N_3782,N_3706);
nand U3862 (N_3862,N_3708,N_3791);
and U3863 (N_3863,N_3723,N_3738);
nand U3864 (N_3864,N_3702,N_3785);
or U3865 (N_3865,N_3756,N_3728);
and U3866 (N_3866,N_3724,N_3736);
nand U3867 (N_3867,N_3755,N_3790);
and U3868 (N_3868,N_3720,N_3709);
nor U3869 (N_3869,N_3719,N_3795);
nand U3870 (N_3870,N_3747,N_3781);
or U3871 (N_3871,N_3753,N_3760);
or U3872 (N_3872,N_3734,N_3706);
nor U3873 (N_3873,N_3717,N_3755);
or U3874 (N_3874,N_3784,N_3794);
nand U3875 (N_3875,N_3734,N_3796);
nor U3876 (N_3876,N_3730,N_3786);
nor U3877 (N_3877,N_3756,N_3759);
nor U3878 (N_3878,N_3739,N_3759);
or U3879 (N_3879,N_3795,N_3708);
nand U3880 (N_3880,N_3781,N_3738);
nor U3881 (N_3881,N_3766,N_3712);
or U3882 (N_3882,N_3701,N_3706);
nand U3883 (N_3883,N_3705,N_3725);
or U3884 (N_3884,N_3746,N_3762);
xor U3885 (N_3885,N_3792,N_3762);
nor U3886 (N_3886,N_3718,N_3773);
xnor U3887 (N_3887,N_3756,N_3747);
nand U3888 (N_3888,N_3748,N_3764);
and U3889 (N_3889,N_3744,N_3721);
nor U3890 (N_3890,N_3762,N_3701);
nor U3891 (N_3891,N_3712,N_3741);
nand U3892 (N_3892,N_3704,N_3733);
and U3893 (N_3893,N_3789,N_3711);
or U3894 (N_3894,N_3724,N_3798);
xnor U3895 (N_3895,N_3721,N_3734);
and U3896 (N_3896,N_3744,N_3797);
xor U3897 (N_3897,N_3760,N_3745);
or U3898 (N_3898,N_3704,N_3799);
nor U3899 (N_3899,N_3757,N_3780);
nand U3900 (N_3900,N_3877,N_3805);
nor U3901 (N_3901,N_3839,N_3878);
and U3902 (N_3902,N_3825,N_3851);
nand U3903 (N_3903,N_3895,N_3870);
nor U3904 (N_3904,N_3844,N_3823);
nor U3905 (N_3905,N_3834,N_3821);
nand U3906 (N_3906,N_3810,N_3854);
xor U3907 (N_3907,N_3872,N_3848);
or U3908 (N_3908,N_3875,N_3861);
and U3909 (N_3909,N_3815,N_3824);
or U3910 (N_3910,N_3892,N_3853);
nor U3911 (N_3911,N_3890,N_3847);
nand U3912 (N_3912,N_3850,N_3829);
nand U3913 (N_3913,N_3894,N_3873);
nor U3914 (N_3914,N_3887,N_3889);
nor U3915 (N_3915,N_3886,N_3813);
nand U3916 (N_3916,N_3803,N_3862);
and U3917 (N_3917,N_3863,N_3860);
or U3918 (N_3918,N_3883,N_3896);
nor U3919 (N_3919,N_3801,N_3898);
nor U3920 (N_3920,N_3893,N_3846);
nor U3921 (N_3921,N_3806,N_3855);
nand U3922 (N_3922,N_3817,N_3897);
and U3923 (N_3923,N_3812,N_3831);
or U3924 (N_3924,N_3818,N_3868);
nor U3925 (N_3925,N_3884,N_3858);
nor U3926 (N_3926,N_3866,N_3835);
or U3927 (N_3927,N_3852,N_3876);
or U3928 (N_3928,N_3869,N_3811);
and U3929 (N_3929,N_3865,N_3856);
or U3930 (N_3930,N_3871,N_3822);
or U3931 (N_3931,N_3807,N_3864);
nand U3932 (N_3932,N_3842,N_3891);
or U3933 (N_3933,N_3840,N_3859);
xor U3934 (N_3934,N_3843,N_3899);
or U3935 (N_3935,N_3880,N_3814);
or U3936 (N_3936,N_3800,N_3830);
nor U3937 (N_3937,N_3836,N_3885);
nor U3938 (N_3938,N_3838,N_3820);
and U3939 (N_3939,N_3837,N_3849);
or U3940 (N_3940,N_3874,N_3826);
nand U3941 (N_3941,N_3857,N_3888);
xor U3942 (N_3942,N_3882,N_3832);
or U3943 (N_3943,N_3881,N_3845);
or U3944 (N_3944,N_3816,N_3828);
or U3945 (N_3945,N_3841,N_3802);
and U3946 (N_3946,N_3827,N_3819);
nand U3947 (N_3947,N_3808,N_3879);
or U3948 (N_3948,N_3804,N_3809);
or U3949 (N_3949,N_3867,N_3833);
or U3950 (N_3950,N_3861,N_3865);
nor U3951 (N_3951,N_3870,N_3832);
and U3952 (N_3952,N_3832,N_3876);
or U3953 (N_3953,N_3882,N_3814);
and U3954 (N_3954,N_3874,N_3823);
nor U3955 (N_3955,N_3874,N_3853);
and U3956 (N_3956,N_3898,N_3849);
and U3957 (N_3957,N_3817,N_3829);
nand U3958 (N_3958,N_3803,N_3834);
xnor U3959 (N_3959,N_3859,N_3814);
nand U3960 (N_3960,N_3831,N_3844);
or U3961 (N_3961,N_3838,N_3882);
or U3962 (N_3962,N_3817,N_3895);
nand U3963 (N_3963,N_3889,N_3802);
nand U3964 (N_3964,N_3851,N_3886);
or U3965 (N_3965,N_3820,N_3854);
and U3966 (N_3966,N_3882,N_3880);
nor U3967 (N_3967,N_3851,N_3870);
and U3968 (N_3968,N_3821,N_3828);
or U3969 (N_3969,N_3811,N_3824);
or U3970 (N_3970,N_3868,N_3886);
or U3971 (N_3971,N_3822,N_3827);
nor U3972 (N_3972,N_3829,N_3819);
nor U3973 (N_3973,N_3846,N_3895);
and U3974 (N_3974,N_3839,N_3837);
xnor U3975 (N_3975,N_3827,N_3866);
and U3976 (N_3976,N_3815,N_3892);
and U3977 (N_3977,N_3832,N_3808);
and U3978 (N_3978,N_3897,N_3829);
nand U3979 (N_3979,N_3822,N_3862);
nand U3980 (N_3980,N_3874,N_3850);
xnor U3981 (N_3981,N_3823,N_3855);
nor U3982 (N_3982,N_3805,N_3837);
nor U3983 (N_3983,N_3810,N_3813);
nor U3984 (N_3984,N_3829,N_3804);
and U3985 (N_3985,N_3876,N_3891);
nor U3986 (N_3986,N_3877,N_3804);
nor U3987 (N_3987,N_3812,N_3859);
nand U3988 (N_3988,N_3885,N_3853);
or U3989 (N_3989,N_3862,N_3850);
and U3990 (N_3990,N_3800,N_3820);
and U3991 (N_3991,N_3893,N_3866);
nand U3992 (N_3992,N_3872,N_3845);
nand U3993 (N_3993,N_3881,N_3870);
and U3994 (N_3994,N_3860,N_3879);
nand U3995 (N_3995,N_3800,N_3826);
and U3996 (N_3996,N_3883,N_3871);
nand U3997 (N_3997,N_3894,N_3846);
or U3998 (N_3998,N_3837,N_3871);
nor U3999 (N_3999,N_3885,N_3880);
or U4000 (N_4000,N_3954,N_3948);
or U4001 (N_4001,N_3907,N_3900);
nor U4002 (N_4002,N_3932,N_3978);
xor U4003 (N_4003,N_3987,N_3906);
and U4004 (N_4004,N_3999,N_3974);
nand U4005 (N_4005,N_3961,N_3905);
or U4006 (N_4006,N_3953,N_3980);
nand U4007 (N_4007,N_3911,N_3975);
nor U4008 (N_4008,N_3997,N_3977);
nor U4009 (N_4009,N_3935,N_3926);
and U4010 (N_4010,N_3910,N_3966);
nand U4011 (N_4011,N_3941,N_3996);
nand U4012 (N_4012,N_3918,N_3973);
and U4013 (N_4013,N_3925,N_3972);
and U4014 (N_4014,N_3934,N_3938);
nand U4015 (N_4015,N_3922,N_3928);
nand U4016 (N_4016,N_3957,N_3937);
or U4017 (N_4017,N_3908,N_3927);
nand U4018 (N_4018,N_3904,N_3981);
and U4019 (N_4019,N_3903,N_3990);
nor U4020 (N_4020,N_3991,N_3936);
xnor U4021 (N_4021,N_3982,N_3914);
nand U4022 (N_4022,N_3963,N_3946);
nor U4023 (N_4023,N_3947,N_3976);
or U4024 (N_4024,N_3939,N_3902);
nor U4025 (N_4025,N_3960,N_3979);
and U4026 (N_4026,N_3912,N_3913);
or U4027 (N_4027,N_3971,N_3952);
and U4028 (N_4028,N_3956,N_3945);
or U4029 (N_4029,N_3964,N_3915);
nor U4030 (N_4030,N_3959,N_3940);
nand U4031 (N_4031,N_3958,N_3909);
nand U4032 (N_4032,N_3920,N_3968);
nand U4033 (N_4033,N_3919,N_3992);
nor U4034 (N_4034,N_3970,N_3929);
and U4035 (N_4035,N_3988,N_3955);
and U4036 (N_4036,N_3994,N_3930);
nand U4037 (N_4037,N_3986,N_3983);
and U4038 (N_4038,N_3917,N_3950);
nor U4039 (N_4039,N_3965,N_3967);
or U4040 (N_4040,N_3944,N_3924);
xnor U4041 (N_4041,N_3949,N_3933);
nor U4042 (N_4042,N_3923,N_3984);
nand U4043 (N_4043,N_3989,N_3969);
nand U4044 (N_4044,N_3995,N_3985);
xnor U4045 (N_4045,N_3931,N_3916);
and U4046 (N_4046,N_3993,N_3901);
or U4047 (N_4047,N_3998,N_3943);
nor U4048 (N_4048,N_3942,N_3962);
and U4049 (N_4049,N_3921,N_3951);
and U4050 (N_4050,N_3964,N_3959);
or U4051 (N_4051,N_3993,N_3945);
or U4052 (N_4052,N_3913,N_3981);
or U4053 (N_4053,N_3981,N_3918);
xnor U4054 (N_4054,N_3906,N_3915);
nand U4055 (N_4055,N_3932,N_3997);
nor U4056 (N_4056,N_3985,N_3950);
nand U4057 (N_4057,N_3900,N_3986);
or U4058 (N_4058,N_3923,N_3951);
and U4059 (N_4059,N_3911,N_3901);
nand U4060 (N_4060,N_3936,N_3970);
xnor U4061 (N_4061,N_3961,N_3994);
nor U4062 (N_4062,N_3910,N_3938);
and U4063 (N_4063,N_3950,N_3921);
and U4064 (N_4064,N_3965,N_3901);
or U4065 (N_4065,N_3922,N_3979);
nand U4066 (N_4066,N_3951,N_3915);
and U4067 (N_4067,N_3920,N_3941);
or U4068 (N_4068,N_3922,N_3998);
and U4069 (N_4069,N_3901,N_3927);
and U4070 (N_4070,N_3917,N_3945);
or U4071 (N_4071,N_3985,N_3953);
or U4072 (N_4072,N_3962,N_3967);
nor U4073 (N_4073,N_3930,N_3989);
or U4074 (N_4074,N_3963,N_3932);
or U4075 (N_4075,N_3958,N_3915);
or U4076 (N_4076,N_3993,N_3934);
nor U4077 (N_4077,N_3918,N_3990);
nand U4078 (N_4078,N_3921,N_3997);
nand U4079 (N_4079,N_3998,N_3940);
nand U4080 (N_4080,N_3955,N_3903);
nand U4081 (N_4081,N_3949,N_3938);
nor U4082 (N_4082,N_3945,N_3933);
xnor U4083 (N_4083,N_3945,N_3963);
and U4084 (N_4084,N_3969,N_3977);
or U4085 (N_4085,N_3977,N_3938);
and U4086 (N_4086,N_3980,N_3922);
and U4087 (N_4087,N_3951,N_3969);
nand U4088 (N_4088,N_3949,N_3991);
and U4089 (N_4089,N_3903,N_3997);
or U4090 (N_4090,N_3925,N_3978);
and U4091 (N_4091,N_3975,N_3901);
or U4092 (N_4092,N_3997,N_3999);
or U4093 (N_4093,N_3980,N_3909);
nand U4094 (N_4094,N_3983,N_3908);
or U4095 (N_4095,N_3942,N_3956);
nor U4096 (N_4096,N_3946,N_3978);
nor U4097 (N_4097,N_3994,N_3959);
or U4098 (N_4098,N_3923,N_3982);
nor U4099 (N_4099,N_3982,N_3962);
or U4100 (N_4100,N_4002,N_4082);
nand U4101 (N_4101,N_4080,N_4064);
or U4102 (N_4102,N_4024,N_4046);
and U4103 (N_4103,N_4099,N_4015);
nor U4104 (N_4104,N_4007,N_4037);
and U4105 (N_4105,N_4068,N_4012);
and U4106 (N_4106,N_4045,N_4013);
and U4107 (N_4107,N_4021,N_4084);
and U4108 (N_4108,N_4086,N_4057);
and U4109 (N_4109,N_4066,N_4028);
and U4110 (N_4110,N_4033,N_4088);
nor U4111 (N_4111,N_4091,N_4003);
or U4112 (N_4112,N_4052,N_4025);
and U4113 (N_4113,N_4072,N_4078);
nor U4114 (N_4114,N_4041,N_4043);
nand U4115 (N_4115,N_4069,N_4048);
nand U4116 (N_4116,N_4085,N_4074);
nor U4117 (N_4117,N_4040,N_4060);
and U4118 (N_4118,N_4009,N_4026);
or U4119 (N_4119,N_4031,N_4093);
or U4120 (N_4120,N_4073,N_4008);
nor U4121 (N_4121,N_4010,N_4035);
or U4122 (N_4122,N_4044,N_4051);
and U4123 (N_4123,N_4098,N_4067);
nand U4124 (N_4124,N_4097,N_4022);
nand U4125 (N_4125,N_4090,N_4059);
or U4126 (N_4126,N_4020,N_4058);
or U4127 (N_4127,N_4063,N_4030);
nor U4128 (N_4128,N_4023,N_4038);
nor U4129 (N_4129,N_4083,N_4032);
and U4130 (N_4130,N_4065,N_4034);
nand U4131 (N_4131,N_4081,N_4001);
nor U4132 (N_4132,N_4053,N_4079);
nand U4133 (N_4133,N_4062,N_4094);
and U4134 (N_4134,N_4016,N_4070);
nand U4135 (N_4135,N_4006,N_4011);
nand U4136 (N_4136,N_4095,N_4089);
or U4137 (N_4137,N_4077,N_4027);
xor U4138 (N_4138,N_4014,N_4029);
nor U4139 (N_4139,N_4004,N_4096);
xnor U4140 (N_4140,N_4055,N_4076);
nor U4141 (N_4141,N_4087,N_4005);
nor U4142 (N_4142,N_4017,N_4042);
nand U4143 (N_4143,N_4047,N_4019);
nor U4144 (N_4144,N_4056,N_4049);
nor U4145 (N_4145,N_4039,N_4061);
nor U4146 (N_4146,N_4054,N_4092);
nand U4147 (N_4147,N_4071,N_4036);
nand U4148 (N_4148,N_4075,N_4050);
and U4149 (N_4149,N_4018,N_4000);
nand U4150 (N_4150,N_4002,N_4098);
or U4151 (N_4151,N_4061,N_4041);
nand U4152 (N_4152,N_4006,N_4026);
nand U4153 (N_4153,N_4055,N_4058);
and U4154 (N_4154,N_4065,N_4037);
and U4155 (N_4155,N_4058,N_4075);
nand U4156 (N_4156,N_4063,N_4038);
nor U4157 (N_4157,N_4074,N_4053);
nand U4158 (N_4158,N_4048,N_4099);
or U4159 (N_4159,N_4020,N_4055);
xnor U4160 (N_4160,N_4054,N_4095);
or U4161 (N_4161,N_4082,N_4025);
nor U4162 (N_4162,N_4035,N_4028);
nand U4163 (N_4163,N_4002,N_4008);
nor U4164 (N_4164,N_4040,N_4033);
and U4165 (N_4165,N_4009,N_4045);
nor U4166 (N_4166,N_4071,N_4057);
and U4167 (N_4167,N_4078,N_4032);
or U4168 (N_4168,N_4079,N_4072);
and U4169 (N_4169,N_4064,N_4015);
or U4170 (N_4170,N_4075,N_4064);
nand U4171 (N_4171,N_4022,N_4033);
nor U4172 (N_4172,N_4037,N_4010);
nor U4173 (N_4173,N_4080,N_4032);
nand U4174 (N_4174,N_4044,N_4062);
nor U4175 (N_4175,N_4061,N_4074);
nand U4176 (N_4176,N_4008,N_4054);
nand U4177 (N_4177,N_4031,N_4004);
and U4178 (N_4178,N_4009,N_4094);
nor U4179 (N_4179,N_4084,N_4056);
and U4180 (N_4180,N_4040,N_4026);
nor U4181 (N_4181,N_4035,N_4000);
and U4182 (N_4182,N_4027,N_4093);
or U4183 (N_4183,N_4006,N_4003);
nand U4184 (N_4184,N_4026,N_4050);
nand U4185 (N_4185,N_4078,N_4039);
nor U4186 (N_4186,N_4040,N_4074);
nor U4187 (N_4187,N_4068,N_4077);
nor U4188 (N_4188,N_4058,N_4085);
xnor U4189 (N_4189,N_4067,N_4004);
or U4190 (N_4190,N_4033,N_4069);
nand U4191 (N_4191,N_4092,N_4025);
nor U4192 (N_4192,N_4079,N_4011);
or U4193 (N_4193,N_4083,N_4026);
nor U4194 (N_4194,N_4060,N_4080);
and U4195 (N_4195,N_4071,N_4092);
or U4196 (N_4196,N_4012,N_4061);
or U4197 (N_4197,N_4048,N_4008);
or U4198 (N_4198,N_4060,N_4016);
nor U4199 (N_4199,N_4036,N_4092);
or U4200 (N_4200,N_4149,N_4156);
nand U4201 (N_4201,N_4150,N_4177);
and U4202 (N_4202,N_4142,N_4132);
nand U4203 (N_4203,N_4130,N_4193);
nand U4204 (N_4204,N_4106,N_4137);
nor U4205 (N_4205,N_4176,N_4166);
and U4206 (N_4206,N_4148,N_4109);
nor U4207 (N_4207,N_4157,N_4111);
and U4208 (N_4208,N_4160,N_4159);
and U4209 (N_4209,N_4141,N_4189);
and U4210 (N_4210,N_4154,N_4100);
nor U4211 (N_4211,N_4131,N_4153);
or U4212 (N_4212,N_4113,N_4195);
and U4213 (N_4213,N_4158,N_4163);
and U4214 (N_4214,N_4172,N_4114);
nor U4215 (N_4215,N_4125,N_4134);
nor U4216 (N_4216,N_4182,N_4191);
nand U4217 (N_4217,N_4138,N_4135);
nor U4218 (N_4218,N_4152,N_4161);
or U4219 (N_4219,N_4129,N_4143);
or U4220 (N_4220,N_4105,N_4115);
and U4221 (N_4221,N_4155,N_4169);
nand U4222 (N_4222,N_4104,N_4121);
or U4223 (N_4223,N_4127,N_4175);
and U4224 (N_4224,N_4194,N_4110);
and U4225 (N_4225,N_4184,N_4108);
nand U4226 (N_4226,N_4185,N_4116);
nand U4227 (N_4227,N_4174,N_4179);
nand U4228 (N_4228,N_4119,N_4186);
nor U4229 (N_4229,N_4196,N_4197);
and U4230 (N_4230,N_4162,N_4122);
nand U4231 (N_4231,N_4183,N_4165);
xnor U4232 (N_4232,N_4145,N_4128);
and U4233 (N_4233,N_4188,N_4139);
or U4234 (N_4234,N_4170,N_4126);
and U4235 (N_4235,N_4178,N_4123);
or U4236 (N_4236,N_4101,N_4151);
nor U4237 (N_4237,N_4198,N_4136);
and U4238 (N_4238,N_4180,N_4102);
nand U4239 (N_4239,N_4133,N_4167);
nand U4240 (N_4240,N_4171,N_4107);
and U4241 (N_4241,N_4168,N_4112);
or U4242 (N_4242,N_4190,N_4146);
nor U4243 (N_4243,N_4140,N_4164);
nand U4244 (N_4244,N_4124,N_4187);
and U4245 (N_4245,N_4117,N_4118);
or U4246 (N_4246,N_4144,N_4192);
nor U4247 (N_4247,N_4199,N_4173);
nand U4248 (N_4248,N_4147,N_4120);
or U4249 (N_4249,N_4103,N_4181);
nand U4250 (N_4250,N_4121,N_4142);
and U4251 (N_4251,N_4123,N_4127);
and U4252 (N_4252,N_4141,N_4144);
and U4253 (N_4253,N_4124,N_4101);
nor U4254 (N_4254,N_4170,N_4197);
nor U4255 (N_4255,N_4197,N_4147);
and U4256 (N_4256,N_4103,N_4198);
nand U4257 (N_4257,N_4172,N_4163);
or U4258 (N_4258,N_4156,N_4117);
or U4259 (N_4259,N_4175,N_4173);
nor U4260 (N_4260,N_4164,N_4165);
nor U4261 (N_4261,N_4146,N_4170);
or U4262 (N_4262,N_4167,N_4188);
nor U4263 (N_4263,N_4143,N_4134);
and U4264 (N_4264,N_4176,N_4196);
or U4265 (N_4265,N_4117,N_4150);
or U4266 (N_4266,N_4139,N_4122);
and U4267 (N_4267,N_4125,N_4121);
and U4268 (N_4268,N_4163,N_4146);
or U4269 (N_4269,N_4139,N_4106);
and U4270 (N_4270,N_4170,N_4171);
nand U4271 (N_4271,N_4114,N_4104);
and U4272 (N_4272,N_4128,N_4129);
and U4273 (N_4273,N_4128,N_4118);
and U4274 (N_4274,N_4132,N_4159);
nand U4275 (N_4275,N_4185,N_4129);
nand U4276 (N_4276,N_4112,N_4105);
and U4277 (N_4277,N_4150,N_4108);
nand U4278 (N_4278,N_4136,N_4156);
or U4279 (N_4279,N_4114,N_4180);
nor U4280 (N_4280,N_4130,N_4182);
or U4281 (N_4281,N_4142,N_4155);
nand U4282 (N_4282,N_4190,N_4186);
nor U4283 (N_4283,N_4162,N_4197);
and U4284 (N_4284,N_4198,N_4179);
nand U4285 (N_4285,N_4114,N_4194);
nor U4286 (N_4286,N_4189,N_4157);
or U4287 (N_4287,N_4189,N_4174);
or U4288 (N_4288,N_4156,N_4160);
or U4289 (N_4289,N_4149,N_4190);
or U4290 (N_4290,N_4116,N_4133);
xor U4291 (N_4291,N_4102,N_4153);
or U4292 (N_4292,N_4165,N_4110);
and U4293 (N_4293,N_4167,N_4172);
nand U4294 (N_4294,N_4113,N_4193);
nand U4295 (N_4295,N_4125,N_4190);
or U4296 (N_4296,N_4161,N_4147);
xnor U4297 (N_4297,N_4110,N_4133);
nor U4298 (N_4298,N_4144,N_4139);
or U4299 (N_4299,N_4184,N_4177);
or U4300 (N_4300,N_4237,N_4261);
nor U4301 (N_4301,N_4248,N_4269);
nand U4302 (N_4302,N_4254,N_4205);
or U4303 (N_4303,N_4262,N_4234);
nor U4304 (N_4304,N_4280,N_4223);
or U4305 (N_4305,N_4271,N_4226);
and U4306 (N_4306,N_4227,N_4284);
nand U4307 (N_4307,N_4244,N_4221);
nor U4308 (N_4308,N_4243,N_4279);
nor U4309 (N_4309,N_4275,N_4277);
nor U4310 (N_4310,N_4213,N_4242);
nor U4311 (N_4311,N_4260,N_4245);
nand U4312 (N_4312,N_4214,N_4217);
nand U4313 (N_4313,N_4209,N_4216);
or U4314 (N_4314,N_4203,N_4294);
or U4315 (N_4315,N_4208,N_4256);
and U4316 (N_4316,N_4225,N_4249);
nor U4317 (N_4317,N_4283,N_4289);
nor U4318 (N_4318,N_4235,N_4298);
and U4319 (N_4319,N_4230,N_4296);
and U4320 (N_4320,N_4270,N_4282);
and U4321 (N_4321,N_4274,N_4204);
and U4322 (N_4322,N_4247,N_4233);
and U4323 (N_4323,N_4295,N_4202);
or U4324 (N_4324,N_4287,N_4246);
nand U4325 (N_4325,N_4236,N_4240);
and U4326 (N_4326,N_4250,N_4281);
nor U4327 (N_4327,N_4253,N_4290);
nand U4328 (N_4328,N_4259,N_4278);
nor U4329 (N_4329,N_4229,N_4268);
or U4330 (N_4330,N_4286,N_4212);
and U4331 (N_4331,N_4276,N_4272);
or U4332 (N_4332,N_4215,N_4258);
and U4333 (N_4333,N_4228,N_4218);
or U4334 (N_4334,N_4273,N_4238);
and U4335 (N_4335,N_4222,N_4255);
and U4336 (N_4336,N_4231,N_4257);
and U4337 (N_4337,N_4292,N_4252);
nand U4338 (N_4338,N_4241,N_4264);
and U4339 (N_4339,N_4201,N_4293);
nand U4340 (N_4340,N_4207,N_4263);
and U4341 (N_4341,N_4285,N_4288);
or U4342 (N_4342,N_4239,N_4206);
nand U4343 (N_4343,N_4219,N_4299);
xor U4344 (N_4344,N_4251,N_4200);
or U4345 (N_4345,N_4224,N_4265);
nor U4346 (N_4346,N_4266,N_4210);
and U4347 (N_4347,N_4297,N_4220);
nor U4348 (N_4348,N_4267,N_4232);
nand U4349 (N_4349,N_4211,N_4291);
or U4350 (N_4350,N_4244,N_4209);
nor U4351 (N_4351,N_4230,N_4237);
or U4352 (N_4352,N_4239,N_4233);
or U4353 (N_4353,N_4267,N_4224);
and U4354 (N_4354,N_4254,N_4269);
and U4355 (N_4355,N_4258,N_4245);
and U4356 (N_4356,N_4237,N_4299);
or U4357 (N_4357,N_4248,N_4264);
or U4358 (N_4358,N_4282,N_4200);
nand U4359 (N_4359,N_4227,N_4251);
nand U4360 (N_4360,N_4282,N_4298);
or U4361 (N_4361,N_4209,N_4252);
or U4362 (N_4362,N_4218,N_4291);
nor U4363 (N_4363,N_4224,N_4217);
and U4364 (N_4364,N_4286,N_4261);
and U4365 (N_4365,N_4238,N_4276);
nor U4366 (N_4366,N_4203,N_4226);
and U4367 (N_4367,N_4226,N_4202);
nor U4368 (N_4368,N_4279,N_4289);
and U4369 (N_4369,N_4202,N_4243);
or U4370 (N_4370,N_4202,N_4208);
nand U4371 (N_4371,N_4260,N_4220);
and U4372 (N_4372,N_4262,N_4283);
nand U4373 (N_4373,N_4222,N_4274);
and U4374 (N_4374,N_4213,N_4215);
nand U4375 (N_4375,N_4253,N_4249);
nor U4376 (N_4376,N_4292,N_4229);
and U4377 (N_4377,N_4295,N_4275);
or U4378 (N_4378,N_4245,N_4241);
and U4379 (N_4379,N_4219,N_4294);
or U4380 (N_4380,N_4243,N_4263);
and U4381 (N_4381,N_4270,N_4267);
and U4382 (N_4382,N_4295,N_4268);
and U4383 (N_4383,N_4245,N_4248);
and U4384 (N_4384,N_4234,N_4255);
and U4385 (N_4385,N_4208,N_4222);
nor U4386 (N_4386,N_4219,N_4231);
nor U4387 (N_4387,N_4215,N_4238);
nor U4388 (N_4388,N_4297,N_4205);
and U4389 (N_4389,N_4209,N_4227);
and U4390 (N_4390,N_4276,N_4286);
and U4391 (N_4391,N_4293,N_4210);
and U4392 (N_4392,N_4219,N_4218);
and U4393 (N_4393,N_4265,N_4286);
and U4394 (N_4394,N_4275,N_4255);
nand U4395 (N_4395,N_4210,N_4262);
or U4396 (N_4396,N_4236,N_4262);
and U4397 (N_4397,N_4262,N_4243);
or U4398 (N_4398,N_4246,N_4278);
nand U4399 (N_4399,N_4287,N_4248);
and U4400 (N_4400,N_4344,N_4338);
nand U4401 (N_4401,N_4334,N_4372);
and U4402 (N_4402,N_4357,N_4306);
nand U4403 (N_4403,N_4399,N_4354);
nand U4404 (N_4404,N_4359,N_4349);
nor U4405 (N_4405,N_4319,N_4360);
and U4406 (N_4406,N_4337,N_4329);
or U4407 (N_4407,N_4331,N_4317);
and U4408 (N_4408,N_4336,N_4316);
nor U4409 (N_4409,N_4308,N_4352);
and U4410 (N_4410,N_4379,N_4304);
and U4411 (N_4411,N_4377,N_4366);
nand U4412 (N_4412,N_4341,N_4323);
or U4413 (N_4413,N_4368,N_4330);
nand U4414 (N_4414,N_4393,N_4335);
nand U4415 (N_4415,N_4356,N_4300);
or U4416 (N_4416,N_4396,N_4353);
nor U4417 (N_4417,N_4386,N_4376);
nand U4418 (N_4418,N_4333,N_4397);
or U4419 (N_4419,N_4387,N_4355);
nor U4420 (N_4420,N_4381,N_4362);
or U4421 (N_4421,N_4325,N_4358);
or U4422 (N_4422,N_4318,N_4378);
nand U4423 (N_4423,N_4347,N_4315);
or U4424 (N_4424,N_4348,N_4384);
or U4425 (N_4425,N_4391,N_4312);
or U4426 (N_4426,N_4320,N_4327);
nor U4427 (N_4427,N_4382,N_4324);
and U4428 (N_4428,N_4380,N_4350);
or U4429 (N_4429,N_4374,N_4388);
and U4430 (N_4430,N_4392,N_4390);
nor U4431 (N_4431,N_4307,N_4321);
and U4432 (N_4432,N_4371,N_4339);
xnor U4433 (N_4433,N_4309,N_4395);
xnor U4434 (N_4434,N_4332,N_4369);
nor U4435 (N_4435,N_4351,N_4367);
and U4436 (N_4436,N_4383,N_4373);
nand U4437 (N_4437,N_4328,N_4361);
and U4438 (N_4438,N_4340,N_4365);
nand U4439 (N_4439,N_4314,N_4311);
and U4440 (N_4440,N_4364,N_4303);
nor U4441 (N_4441,N_4363,N_4346);
and U4442 (N_4442,N_4389,N_4305);
nor U4443 (N_4443,N_4302,N_4345);
nor U4444 (N_4444,N_4343,N_4301);
or U4445 (N_4445,N_4313,N_4398);
or U4446 (N_4446,N_4375,N_4385);
and U4447 (N_4447,N_4394,N_4370);
and U4448 (N_4448,N_4326,N_4322);
nor U4449 (N_4449,N_4310,N_4342);
nand U4450 (N_4450,N_4353,N_4304);
and U4451 (N_4451,N_4333,N_4359);
nor U4452 (N_4452,N_4340,N_4319);
nor U4453 (N_4453,N_4373,N_4396);
or U4454 (N_4454,N_4354,N_4333);
and U4455 (N_4455,N_4398,N_4382);
or U4456 (N_4456,N_4309,N_4389);
and U4457 (N_4457,N_4364,N_4398);
or U4458 (N_4458,N_4301,N_4399);
and U4459 (N_4459,N_4339,N_4306);
nand U4460 (N_4460,N_4394,N_4337);
nor U4461 (N_4461,N_4348,N_4358);
or U4462 (N_4462,N_4349,N_4358);
nor U4463 (N_4463,N_4342,N_4346);
nor U4464 (N_4464,N_4308,N_4375);
or U4465 (N_4465,N_4350,N_4352);
nand U4466 (N_4466,N_4372,N_4307);
nor U4467 (N_4467,N_4327,N_4353);
nor U4468 (N_4468,N_4330,N_4361);
nor U4469 (N_4469,N_4391,N_4382);
or U4470 (N_4470,N_4309,N_4339);
and U4471 (N_4471,N_4378,N_4358);
nand U4472 (N_4472,N_4368,N_4301);
or U4473 (N_4473,N_4343,N_4381);
nor U4474 (N_4474,N_4359,N_4384);
nand U4475 (N_4475,N_4393,N_4317);
or U4476 (N_4476,N_4351,N_4352);
nand U4477 (N_4477,N_4305,N_4340);
or U4478 (N_4478,N_4389,N_4350);
nor U4479 (N_4479,N_4368,N_4399);
and U4480 (N_4480,N_4370,N_4378);
or U4481 (N_4481,N_4302,N_4369);
and U4482 (N_4482,N_4327,N_4347);
or U4483 (N_4483,N_4389,N_4399);
nand U4484 (N_4484,N_4342,N_4361);
and U4485 (N_4485,N_4302,N_4372);
nand U4486 (N_4486,N_4319,N_4369);
nor U4487 (N_4487,N_4332,N_4352);
nand U4488 (N_4488,N_4364,N_4310);
nand U4489 (N_4489,N_4351,N_4364);
and U4490 (N_4490,N_4390,N_4335);
xnor U4491 (N_4491,N_4390,N_4308);
nor U4492 (N_4492,N_4305,N_4325);
and U4493 (N_4493,N_4393,N_4302);
nor U4494 (N_4494,N_4335,N_4332);
xor U4495 (N_4495,N_4370,N_4338);
nor U4496 (N_4496,N_4327,N_4383);
and U4497 (N_4497,N_4365,N_4373);
or U4498 (N_4498,N_4395,N_4367);
nand U4499 (N_4499,N_4376,N_4306);
nand U4500 (N_4500,N_4476,N_4431);
or U4501 (N_4501,N_4425,N_4404);
and U4502 (N_4502,N_4468,N_4445);
nor U4503 (N_4503,N_4470,N_4459);
nor U4504 (N_4504,N_4441,N_4411);
and U4505 (N_4505,N_4475,N_4403);
or U4506 (N_4506,N_4478,N_4440);
nand U4507 (N_4507,N_4498,N_4472);
and U4508 (N_4508,N_4483,N_4439);
or U4509 (N_4509,N_4433,N_4462);
nand U4510 (N_4510,N_4435,N_4443);
or U4511 (N_4511,N_4499,N_4466);
and U4512 (N_4512,N_4492,N_4457);
or U4513 (N_4513,N_4451,N_4465);
nand U4514 (N_4514,N_4494,N_4495);
nand U4515 (N_4515,N_4408,N_4450);
nor U4516 (N_4516,N_4484,N_4497);
and U4517 (N_4517,N_4409,N_4458);
xor U4518 (N_4518,N_4456,N_4463);
nand U4519 (N_4519,N_4415,N_4416);
nor U4520 (N_4520,N_4452,N_4421);
or U4521 (N_4521,N_4434,N_4461);
nand U4522 (N_4522,N_4474,N_4471);
and U4523 (N_4523,N_4401,N_4413);
or U4524 (N_4524,N_4464,N_4430);
nor U4525 (N_4525,N_4428,N_4407);
or U4526 (N_4526,N_4487,N_4423);
nor U4527 (N_4527,N_4481,N_4454);
nor U4528 (N_4528,N_4410,N_4467);
xor U4529 (N_4529,N_4400,N_4460);
nor U4530 (N_4530,N_4426,N_4414);
nand U4531 (N_4531,N_4473,N_4489);
nor U4532 (N_4532,N_4479,N_4469);
xnor U4533 (N_4533,N_4448,N_4419);
nand U4534 (N_4534,N_4491,N_4482);
and U4535 (N_4535,N_4449,N_4488);
or U4536 (N_4536,N_4438,N_4442);
nand U4537 (N_4537,N_4446,N_4455);
and U4538 (N_4538,N_4485,N_4417);
nor U4539 (N_4539,N_4490,N_4496);
nand U4540 (N_4540,N_4432,N_4437);
nor U4541 (N_4541,N_4412,N_4418);
and U4542 (N_4542,N_4424,N_4406);
nand U4543 (N_4543,N_4477,N_4480);
nand U4544 (N_4544,N_4436,N_4420);
and U4545 (N_4545,N_4444,N_4493);
nand U4546 (N_4546,N_4422,N_4447);
nor U4547 (N_4547,N_4453,N_4429);
or U4548 (N_4548,N_4405,N_4402);
nand U4549 (N_4549,N_4427,N_4486);
and U4550 (N_4550,N_4418,N_4429);
and U4551 (N_4551,N_4433,N_4427);
nand U4552 (N_4552,N_4452,N_4442);
and U4553 (N_4553,N_4494,N_4405);
or U4554 (N_4554,N_4437,N_4450);
xor U4555 (N_4555,N_4431,N_4481);
nor U4556 (N_4556,N_4441,N_4446);
or U4557 (N_4557,N_4404,N_4457);
nor U4558 (N_4558,N_4475,N_4474);
nor U4559 (N_4559,N_4408,N_4411);
or U4560 (N_4560,N_4467,N_4448);
nand U4561 (N_4561,N_4488,N_4404);
nand U4562 (N_4562,N_4488,N_4455);
or U4563 (N_4563,N_4499,N_4487);
or U4564 (N_4564,N_4416,N_4453);
and U4565 (N_4565,N_4480,N_4470);
nand U4566 (N_4566,N_4472,N_4488);
nand U4567 (N_4567,N_4457,N_4476);
nand U4568 (N_4568,N_4434,N_4478);
nand U4569 (N_4569,N_4439,N_4478);
xnor U4570 (N_4570,N_4452,N_4448);
or U4571 (N_4571,N_4434,N_4419);
xor U4572 (N_4572,N_4499,N_4459);
and U4573 (N_4573,N_4469,N_4459);
and U4574 (N_4574,N_4428,N_4452);
nand U4575 (N_4575,N_4447,N_4431);
nand U4576 (N_4576,N_4493,N_4408);
and U4577 (N_4577,N_4404,N_4426);
nor U4578 (N_4578,N_4443,N_4449);
nor U4579 (N_4579,N_4443,N_4447);
nor U4580 (N_4580,N_4494,N_4498);
nand U4581 (N_4581,N_4428,N_4471);
nand U4582 (N_4582,N_4411,N_4473);
and U4583 (N_4583,N_4459,N_4416);
or U4584 (N_4584,N_4451,N_4455);
and U4585 (N_4585,N_4476,N_4488);
nand U4586 (N_4586,N_4462,N_4498);
and U4587 (N_4587,N_4437,N_4482);
or U4588 (N_4588,N_4417,N_4486);
nand U4589 (N_4589,N_4417,N_4456);
nand U4590 (N_4590,N_4400,N_4434);
and U4591 (N_4591,N_4427,N_4415);
and U4592 (N_4592,N_4421,N_4486);
or U4593 (N_4593,N_4430,N_4469);
or U4594 (N_4594,N_4467,N_4442);
and U4595 (N_4595,N_4491,N_4419);
and U4596 (N_4596,N_4494,N_4419);
or U4597 (N_4597,N_4484,N_4498);
or U4598 (N_4598,N_4407,N_4481);
and U4599 (N_4599,N_4413,N_4493);
nand U4600 (N_4600,N_4575,N_4517);
nand U4601 (N_4601,N_4587,N_4567);
nand U4602 (N_4602,N_4505,N_4535);
or U4603 (N_4603,N_4516,N_4553);
nor U4604 (N_4604,N_4566,N_4557);
nand U4605 (N_4605,N_4564,N_4511);
nand U4606 (N_4606,N_4509,N_4545);
and U4607 (N_4607,N_4506,N_4508);
nor U4608 (N_4608,N_4562,N_4594);
nand U4609 (N_4609,N_4599,N_4552);
or U4610 (N_4610,N_4561,N_4504);
and U4611 (N_4611,N_4558,N_4555);
xor U4612 (N_4612,N_4591,N_4588);
nor U4613 (N_4613,N_4534,N_4538);
nand U4614 (N_4614,N_4548,N_4597);
or U4615 (N_4615,N_4518,N_4572);
and U4616 (N_4616,N_4565,N_4581);
nor U4617 (N_4617,N_4573,N_4503);
nor U4618 (N_4618,N_4593,N_4524);
nand U4619 (N_4619,N_4579,N_4549);
and U4620 (N_4620,N_4531,N_4513);
or U4621 (N_4621,N_4570,N_4583);
nand U4622 (N_4622,N_4554,N_4560);
nand U4623 (N_4623,N_4590,N_4577);
nand U4624 (N_4624,N_4522,N_4574);
and U4625 (N_4625,N_4595,N_4532);
nor U4626 (N_4626,N_4585,N_4507);
nand U4627 (N_4627,N_4556,N_4541);
and U4628 (N_4628,N_4576,N_4542);
nor U4629 (N_4629,N_4521,N_4536);
and U4630 (N_4630,N_4596,N_4501);
nor U4631 (N_4631,N_4529,N_4500);
or U4632 (N_4632,N_4540,N_4519);
nand U4633 (N_4633,N_4528,N_4598);
nor U4634 (N_4634,N_4547,N_4515);
nor U4635 (N_4635,N_4520,N_4527);
nor U4636 (N_4636,N_4523,N_4546);
nand U4637 (N_4637,N_4582,N_4571);
nor U4638 (N_4638,N_4512,N_4569);
nand U4639 (N_4639,N_4563,N_4580);
or U4640 (N_4640,N_4551,N_4537);
and U4641 (N_4641,N_4530,N_4586);
nand U4642 (N_4642,N_4510,N_4592);
and U4643 (N_4643,N_4526,N_4543);
nand U4644 (N_4644,N_4550,N_4578);
or U4645 (N_4645,N_4539,N_4559);
nand U4646 (N_4646,N_4584,N_4525);
nor U4647 (N_4647,N_4502,N_4589);
nand U4648 (N_4648,N_4514,N_4533);
or U4649 (N_4649,N_4544,N_4568);
or U4650 (N_4650,N_4558,N_4503);
nor U4651 (N_4651,N_4594,N_4555);
nor U4652 (N_4652,N_4565,N_4523);
nand U4653 (N_4653,N_4562,N_4557);
nand U4654 (N_4654,N_4595,N_4517);
nor U4655 (N_4655,N_4538,N_4581);
nand U4656 (N_4656,N_4583,N_4543);
nor U4657 (N_4657,N_4513,N_4578);
and U4658 (N_4658,N_4573,N_4504);
and U4659 (N_4659,N_4505,N_4530);
and U4660 (N_4660,N_4587,N_4549);
and U4661 (N_4661,N_4570,N_4598);
and U4662 (N_4662,N_4585,N_4540);
or U4663 (N_4663,N_4595,N_4587);
nor U4664 (N_4664,N_4529,N_4599);
nor U4665 (N_4665,N_4509,N_4551);
or U4666 (N_4666,N_4587,N_4583);
and U4667 (N_4667,N_4598,N_4511);
nor U4668 (N_4668,N_4561,N_4521);
nand U4669 (N_4669,N_4598,N_4591);
nor U4670 (N_4670,N_4515,N_4542);
nand U4671 (N_4671,N_4563,N_4564);
nor U4672 (N_4672,N_4574,N_4554);
nand U4673 (N_4673,N_4546,N_4525);
nand U4674 (N_4674,N_4519,N_4528);
nand U4675 (N_4675,N_4566,N_4596);
and U4676 (N_4676,N_4539,N_4531);
nor U4677 (N_4677,N_4529,N_4574);
xor U4678 (N_4678,N_4502,N_4592);
and U4679 (N_4679,N_4510,N_4578);
nand U4680 (N_4680,N_4590,N_4547);
nor U4681 (N_4681,N_4510,N_4590);
nand U4682 (N_4682,N_4518,N_4579);
and U4683 (N_4683,N_4559,N_4517);
nand U4684 (N_4684,N_4561,N_4574);
nand U4685 (N_4685,N_4517,N_4585);
or U4686 (N_4686,N_4522,N_4513);
nand U4687 (N_4687,N_4540,N_4547);
and U4688 (N_4688,N_4599,N_4580);
or U4689 (N_4689,N_4577,N_4552);
or U4690 (N_4690,N_4513,N_4502);
nand U4691 (N_4691,N_4599,N_4568);
nand U4692 (N_4692,N_4521,N_4583);
nand U4693 (N_4693,N_4529,N_4580);
or U4694 (N_4694,N_4578,N_4568);
nor U4695 (N_4695,N_4583,N_4559);
xnor U4696 (N_4696,N_4583,N_4503);
nand U4697 (N_4697,N_4508,N_4571);
nand U4698 (N_4698,N_4504,N_4566);
nor U4699 (N_4699,N_4580,N_4557);
and U4700 (N_4700,N_4608,N_4618);
nor U4701 (N_4701,N_4627,N_4678);
or U4702 (N_4702,N_4665,N_4600);
and U4703 (N_4703,N_4664,N_4616);
and U4704 (N_4704,N_4699,N_4611);
nand U4705 (N_4705,N_4651,N_4612);
nand U4706 (N_4706,N_4692,N_4650);
nand U4707 (N_4707,N_4646,N_4657);
nand U4708 (N_4708,N_4666,N_4684);
xnor U4709 (N_4709,N_4621,N_4647);
nor U4710 (N_4710,N_4673,N_4663);
or U4711 (N_4711,N_4668,N_4652);
and U4712 (N_4712,N_4683,N_4636);
xor U4713 (N_4713,N_4698,N_4662);
nand U4714 (N_4714,N_4632,N_4686);
nor U4715 (N_4715,N_4640,N_4679);
nor U4716 (N_4716,N_4660,N_4639);
and U4717 (N_4717,N_4631,N_4688);
and U4718 (N_4718,N_4638,N_4603);
and U4719 (N_4719,N_4635,N_4623);
nor U4720 (N_4720,N_4643,N_4674);
nand U4721 (N_4721,N_4677,N_4671);
nor U4722 (N_4722,N_4625,N_4676);
nand U4723 (N_4723,N_4630,N_4667);
nor U4724 (N_4724,N_4648,N_4693);
nand U4725 (N_4725,N_4680,N_4637);
and U4726 (N_4726,N_4624,N_4644);
and U4727 (N_4727,N_4656,N_4687);
nor U4728 (N_4728,N_4685,N_4659);
nand U4729 (N_4729,N_4697,N_4669);
or U4730 (N_4730,N_4689,N_4670);
nor U4731 (N_4731,N_4610,N_4654);
nor U4732 (N_4732,N_4696,N_4620);
nand U4733 (N_4733,N_4642,N_4622);
nor U4734 (N_4734,N_4602,N_4691);
nor U4735 (N_4735,N_4653,N_4614);
or U4736 (N_4736,N_4649,N_4607);
nor U4737 (N_4737,N_4661,N_4655);
nand U4738 (N_4738,N_4601,N_4634);
and U4739 (N_4739,N_4645,N_4604);
nor U4740 (N_4740,N_4617,N_4641);
nand U4741 (N_4741,N_4633,N_4615);
nand U4742 (N_4742,N_4609,N_4694);
nor U4743 (N_4743,N_4605,N_4682);
nor U4744 (N_4744,N_4606,N_4629);
and U4745 (N_4745,N_4626,N_4681);
and U4746 (N_4746,N_4690,N_4619);
or U4747 (N_4747,N_4695,N_4628);
or U4748 (N_4748,N_4675,N_4672);
and U4749 (N_4749,N_4613,N_4658);
or U4750 (N_4750,N_4635,N_4649);
nand U4751 (N_4751,N_4616,N_4693);
nand U4752 (N_4752,N_4678,N_4661);
or U4753 (N_4753,N_4694,N_4652);
or U4754 (N_4754,N_4602,N_4641);
nand U4755 (N_4755,N_4642,N_4688);
nand U4756 (N_4756,N_4653,N_4609);
and U4757 (N_4757,N_4675,N_4609);
nand U4758 (N_4758,N_4643,N_4690);
or U4759 (N_4759,N_4611,N_4646);
and U4760 (N_4760,N_4623,N_4669);
and U4761 (N_4761,N_4662,N_4637);
nor U4762 (N_4762,N_4659,N_4646);
nand U4763 (N_4763,N_4654,N_4645);
nor U4764 (N_4764,N_4694,N_4628);
nor U4765 (N_4765,N_4673,N_4661);
or U4766 (N_4766,N_4671,N_4611);
or U4767 (N_4767,N_4613,N_4633);
or U4768 (N_4768,N_4626,N_4693);
nor U4769 (N_4769,N_4642,N_4637);
and U4770 (N_4770,N_4629,N_4655);
nand U4771 (N_4771,N_4625,N_4660);
nand U4772 (N_4772,N_4656,N_4664);
or U4773 (N_4773,N_4680,N_4602);
or U4774 (N_4774,N_4649,N_4652);
or U4775 (N_4775,N_4665,N_4697);
nor U4776 (N_4776,N_4657,N_4651);
and U4777 (N_4777,N_4697,N_4651);
or U4778 (N_4778,N_4651,N_4632);
nor U4779 (N_4779,N_4689,N_4684);
and U4780 (N_4780,N_4691,N_4614);
nand U4781 (N_4781,N_4628,N_4636);
or U4782 (N_4782,N_4627,N_4692);
nor U4783 (N_4783,N_4625,N_4658);
or U4784 (N_4784,N_4636,N_4612);
nor U4785 (N_4785,N_4684,N_4606);
and U4786 (N_4786,N_4607,N_4690);
or U4787 (N_4787,N_4608,N_4689);
and U4788 (N_4788,N_4663,N_4675);
nand U4789 (N_4789,N_4635,N_4678);
nand U4790 (N_4790,N_4672,N_4686);
and U4791 (N_4791,N_4692,N_4624);
and U4792 (N_4792,N_4606,N_4654);
nand U4793 (N_4793,N_4644,N_4619);
or U4794 (N_4794,N_4605,N_4648);
nor U4795 (N_4795,N_4602,N_4698);
and U4796 (N_4796,N_4629,N_4659);
or U4797 (N_4797,N_4633,N_4689);
nand U4798 (N_4798,N_4611,N_4686);
nor U4799 (N_4799,N_4677,N_4695);
and U4800 (N_4800,N_4770,N_4735);
nand U4801 (N_4801,N_4748,N_4754);
nand U4802 (N_4802,N_4739,N_4701);
and U4803 (N_4803,N_4796,N_4791);
nor U4804 (N_4804,N_4743,N_4798);
or U4805 (N_4805,N_4734,N_4787);
or U4806 (N_4806,N_4708,N_4780);
and U4807 (N_4807,N_4722,N_4745);
nor U4808 (N_4808,N_4714,N_4768);
or U4809 (N_4809,N_4730,N_4793);
or U4810 (N_4810,N_4725,N_4712);
or U4811 (N_4811,N_4774,N_4795);
nand U4812 (N_4812,N_4716,N_4727);
nor U4813 (N_4813,N_4707,N_4717);
and U4814 (N_4814,N_4729,N_4741);
nand U4815 (N_4815,N_4713,N_4749);
and U4816 (N_4816,N_4789,N_4711);
or U4817 (N_4817,N_4705,N_4794);
nor U4818 (N_4818,N_4723,N_4778);
or U4819 (N_4819,N_4760,N_4753);
and U4820 (N_4820,N_4732,N_4763);
and U4821 (N_4821,N_4757,N_4790);
nor U4822 (N_4822,N_4799,N_4766);
or U4823 (N_4823,N_4733,N_4724);
nor U4824 (N_4824,N_4736,N_4746);
or U4825 (N_4825,N_4744,N_4755);
and U4826 (N_4826,N_4776,N_4703);
nand U4827 (N_4827,N_4700,N_4775);
or U4828 (N_4828,N_4718,N_4773);
and U4829 (N_4829,N_4720,N_4737);
nand U4830 (N_4830,N_4704,N_4764);
nand U4831 (N_4831,N_4797,N_4792);
or U4832 (N_4832,N_4786,N_4756);
nor U4833 (N_4833,N_4769,N_4772);
or U4834 (N_4834,N_4750,N_4747);
nand U4835 (N_4835,N_4731,N_4715);
nand U4836 (N_4836,N_4765,N_4738);
nor U4837 (N_4837,N_4762,N_4709);
nor U4838 (N_4838,N_4719,N_4702);
nor U4839 (N_4839,N_4740,N_4761);
nand U4840 (N_4840,N_4710,N_4751);
and U4841 (N_4841,N_4783,N_4742);
and U4842 (N_4842,N_4779,N_4784);
or U4843 (N_4843,N_4726,N_4752);
or U4844 (N_4844,N_4706,N_4782);
nor U4845 (N_4845,N_4759,N_4728);
or U4846 (N_4846,N_4777,N_4767);
nor U4847 (N_4847,N_4758,N_4721);
and U4848 (N_4848,N_4781,N_4771);
nor U4849 (N_4849,N_4788,N_4785);
nand U4850 (N_4850,N_4737,N_4724);
or U4851 (N_4851,N_4707,N_4734);
and U4852 (N_4852,N_4794,N_4784);
nand U4853 (N_4853,N_4766,N_4753);
or U4854 (N_4854,N_4706,N_4775);
and U4855 (N_4855,N_4764,N_4774);
nor U4856 (N_4856,N_4795,N_4779);
nand U4857 (N_4857,N_4787,N_4784);
nand U4858 (N_4858,N_4771,N_4702);
nand U4859 (N_4859,N_4718,N_4755);
and U4860 (N_4860,N_4741,N_4786);
nor U4861 (N_4861,N_4789,N_4748);
nand U4862 (N_4862,N_4752,N_4769);
or U4863 (N_4863,N_4727,N_4753);
nor U4864 (N_4864,N_4754,N_4782);
nand U4865 (N_4865,N_4723,N_4751);
nand U4866 (N_4866,N_4793,N_4705);
nor U4867 (N_4867,N_4727,N_4751);
nand U4868 (N_4868,N_4768,N_4775);
or U4869 (N_4869,N_4768,N_4791);
nor U4870 (N_4870,N_4760,N_4769);
or U4871 (N_4871,N_4760,N_4740);
or U4872 (N_4872,N_4754,N_4729);
nor U4873 (N_4873,N_4743,N_4711);
nor U4874 (N_4874,N_4787,N_4796);
nor U4875 (N_4875,N_4706,N_4711);
xor U4876 (N_4876,N_4756,N_4703);
and U4877 (N_4877,N_4719,N_4764);
and U4878 (N_4878,N_4728,N_4729);
nand U4879 (N_4879,N_4799,N_4785);
nor U4880 (N_4880,N_4770,N_4739);
nand U4881 (N_4881,N_4796,N_4737);
nand U4882 (N_4882,N_4700,N_4749);
or U4883 (N_4883,N_4731,N_4733);
nor U4884 (N_4884,N_4792,N_4786);
nor U4885 (N_4885,N_4795,N_4728);
nand U4886 (N_4886,N_4727,N_4778);
nor U4887 (N_4887,N_4754,N_4749);
or U4888 (N_4888,N_4783,N_4789);
xor U4889 (N_4889,N_4777,N_4726);
xnor U4890 (N_4890,N_4759,N_4727);
and U4891 (N_4891,N_4748,N_4774);
nor U4892 (N_4892,N_4726,N_4766);
and U4893 (N_4893,N_4791,N_4771);
and U4894 (N_4894,N_4788,N_4750);
or U4895 (N_4895,N_4732,N_4724);
nand U4896 (N_4896,N_4727,N_4715);
nor U4897 (N_4897,N_4764,N_4743);
or U4898 (N_4898,N_4746,N_4759);
nor U4899 (N_4899,N_4798,N_4719);
xor U4900 (N_4900,N_4819,N_4859);
nor U4901 (N_4901,N_4850,N_4847);
nor U4902 (N_4902,N_4845,N_4866);
nor U4903 (N_4903,N_4855,N_4826);
or U4904 (N_4904,N_4827,N_4839);
nand U4905 (N_4905,N_4880,N_4864);
xnor U4906 (N_4906,N_4884,N_4806);
or U4907 (N_4907,N_4860,N_4846);
nand U4908 (N_4908,N_4882,N_4803);
nand U4909 (N_4909,N_4840,N_4804);
or U4910 (N_4910,N_4897,N_4878);
nor U4911 (N_4911,N_4816,N_4872);
nor U4912 (N_4912,N_4867,N_4874);
or U4913 (N_4913,N_4852,N_4899);
nand U4914 (N_4914,N_4853,N_4894);
nor U4915 (N_4915,N_4814,N_4865);
nand U4916 (N_4916,N_4858,N_4810);
nand U4917 (N_4917,N_4862,N_4818);
or U4918 (N_4918,N_4876,N_4832);
or U4919 (N_4919,N_4833,N_4849);
nand U4920 (N_4920,N_4811,N_4813);
nor U4921 (N_4921,N_4830,N_4815);
and U4922 (N_4922,N_4841,N_4886);
or U4923 (N_4923,N_4891,N_4892);
nand U4924 (N_4924,N_4896,N_4800);
or U4925 (N_4925,N_4883,N_4854);
nor U4926 (N_4926,N_4805,N_4885);
nand U4927 (N_4927,N_4857,N_4822);
or U4928 (N_4928,N_4837,N_4869);
and U4929 (N_4929,N_4817,N_4820);
or U4930 (N_4930,N_4823,N_4835);
or U4931 (N_4931,N_4873,N_4856);
and U4932 (N_4932,N_4890,N_4861);
and U4933 (N_4933,N_4848,N_4871);
or U4934 (N_4934,N_4895,N_4863);
or U4935 (N_4935,N_4879,N_4842);
nand U4936 (N_4936,N_4844,N_4831);
nor U4937 (N_4937,N_4825,N_4807);
and U4938 (N_4938,N_4893,N_4898);
nor U4939 (N_4939,N_4875,N_4838);
nand U4940 (N_4940,N_4843,N_4888);
nor U4941 (N_4941,N_4801,N_4868);
nand U4942 (N_4942,N_4821,N_4829);
or U4943 (N_4943,N_4828,N_4834);
and U4944 (N_4944,N_4877,N_4889);
and U4945 (N_4945,N_4809,N_4824);
nor U4946 (N_4946,N_4887,N_4802);
and U4947 (N_4947,N_4881,N_4836);
and U4948 (N_4948,N_4812,N_4851);
or U4949 (N_4949,N_4870,N_4808);
nor U4950 (N_4950,N_4899,N_4829);
nor U4951 (N_4951,N_4880,N_4847);
and U4952 (N_4952,N_4831,N_4810);
nor U4953 (N_4953,N_4850,N_4899);
or U4954 (N_4954,N_4867,N_4857);
nor U4955 (N_4955,N_4805,N_4837);
or U4956 (N_4956,N_4814,N_4850);
nand U4957 (N_4957,N_4898,N_4864);
nor U4958 (N_4958,N_4875,N_4820);
nor U4959 (N_4959,N_4866,N_4890);
and U4960 (N_4960,N_4822,N_4884);
and U4961 (N_4961,N_4805,N_4857);
nand U4962 (N_4962,N_4848,N_4868);
or U4963 (N_4963,N_4893,N_4859);
nand U4964 (N_4964,N_4876,N_4873);
nand U4965 (N_4965,N_4873,N_4853);
and U4966 (N_4966,N_4894,N_4812);
nor U4967 (N_4967,N_4821,N_4882);
or U4968 (N_4968,N_4810,N_4841);
and U4969 (N_4969,N_4896,N_4804);
nor U4970 (N_4970,N_4890,N_4809);
or U4971 (N_4971,N_4825,N_4869);
and U4972 (N_4972,N_4841,N_4848);
or U4973 (N_4973,N_4891,N_4841);
and U4974 (N_4974,N_4829,N_4867);
or U4975 (N_4975,N_4856,N_4880);
nand U4976 (N_4976,N_4802,N_4863);
nand U4977 (N_4977,N_4804,N_4806);
and U4978 (N_4978,N_4825,N_4803);
and U4979 (N_4979,N_4882,N_4852);
nor U4980 (N_4980,N_4807,N_4849);
xnor U4981 (N_4981,N_4829,N_4828);
nand U4982 (N_4982,N_4868,N_4812);
nand U4983 (N_4983,N_4876,N_4857);
nor U4984 (N_4984,N_4817,N_4831);
or U4985 (N_4985,N_4851,N_4884);
and U4986 (N_4986,N_4873,N_4813);
nor U4987 (N_4987,N_4877,N_4812);
and U4988 (N_4988,N_4803,N_4861);
and U4989 (N_4989,N_4874,N_4800);
nand U4990 (N_4990,N_4836,N_4865);
or U4991 (N_4991,N_4845,N_4813);
nor U4992 (N_4992,N_4872,N_4820);
nand U4993 (N_4993,N_4833,N_4898);
nand U4994 (N_4994,N_4877,N_4898);
or U4995 (N_4995,N_4876,N_4872);
nor U4996 (N_4996,N_4884,N_4824);
or U4997 (N_4997,N_4802,N_4866);
or U4998 (N_4998,N_4828,N_4803);
nand U4999 (N_4999,N_4876,N_4885);
and U5000 (N_5000,N_4941,N_4970);
nor U5001 (N_5001,N_4950,N_4919);
nor U5002 (N_5002,N_4914,N_4988);
and U5003 (N_5003,N_4904,N_4909);
and U5004 (N_5004,N_4974,N_4984);
nor U5005 (N_5005,N_4900,N_4963);
and U5006 (N_5006,N_4953,N_4976);
or U5007 (N_5007,N_4949,N_4918);
and U5008 (N_5008,N_4930,N_4969);
or U5009 (N_5009,N_4958,N_4986);
nand U5010 (N_5010,N_4975,N_4973);
nor U5011 (N_5011,N_4936,N_4981);
nand U5012 (N_5012,N_4994,N_4987);
nor U5013 (N_5013,N_4916,N_4947);
or U5014 (N_5014,N_4964,N_4942);
nand U5015 (N_5015,N_4907,N_4902);
or U5016 (N_5016,N_4935,N_4990);
and U5017 (N_5017,N_4960,N_4903);
nor U5018 (N_5018,N_4929,N_4989);
and U5019 (N_5019,N_4979,N_4998);
nor U5020 (N_5020,N_4971,N_4952);
nand U5021 (N_5021,N_4978,N_4925);
and U5022 (N_5022,N_4945,N_4999);
nand U5023 (N_5023,N_4993,N_4922);
nor U5024 (N_5024,N_4956,N_4906);
or U5025 (N_5025,N_4944,N_4997);
and U5026 (N_5026,N_4991,N_4980);
nand U5027 (N_5027,N_4995,N_4917);
or U5028 (N_5028,N_4911,N_4908);
nand U5029 (N_5029,N_4954,N_4966);
nor U5030 (N_5030,N_4901,N_4915);
or U5031 (N_5031,N_4968,N_4913);
xor U5032 (N_5032,N_4951,N_4962);
nand U5033 (N_5033,N_4939,N_4967);
or U5034 (N_5034,N_4961,N_4937);
nor U5035 (N_5035,N_4912,N_4957);
and U5036 (N_5036,N_4910,N_4983);
nand U5037 (N_5037,N_4934,N_4972);
and U5038 (N_5038,N_4946,N_4923);
nor U5039 (N_5039,N_4959,N_4927);
nand U5040 (N_5040,N_4926,N_4985);
or U5041 (N_5041,N_4996,N_4940);
or U5042 (N_5042,N_4965,N_4932);
nand U5043 (N_5043,N_4948,N_4982);
and U5044 (N_5044,N_4928,N_4933);
and U5045 (N_5045,N_4992,N_4921);
nor U5046 (N_5046,N_4955,N_4977);
and U5047 (N_5047,N_4931,N_4938);
nand U5048 (N_5048,N_4943,N_4924);
and U5049 (N_5049,N_4920,N_4905);
nand U5050 (N_5050,N_4952,N_4980);
and U5051 (N_5051,N_4903,N_4941);
or U5052 (N_5052,N_4940,N_4906);
nand U5053 (N_5053,N_4922,N_4916);
nand U5054 (N_5054,N_4991,N_4919);
nor U5055 (N_5055,N_4922,N_4949);
or U5056 (N_5056,N_4941,N_4957);
nand U5057 (N_5057,N_4929,N_4948);
or U5058 (N_5058,N_4916,N_4972);
and U5059 (N_5059,N_4971,N_4930);
or U5060 (N_5060,N_4985,N_4962);
nor U5061 (N_5061,N_4997,N_4959);
nand U5062 (N_5062,N_4949,N_4919);
or U5063 (N_5063,N_4980,N_4916);
xnor U5064 (N_5064,N_4928,N_4944);
nor U5065 (N_5065,N_4917,N_4969);
and U5066 (N_5066,N_4968,N_4905);
nor U5067 (N_5067,N_4984,N_4966);
and U5068 (N_5068,N_4945,N_4925);
or U5069 (N_5069,N_4979,N_4972);
nand U5070 (N_5070,N_4914,N_4909);
or U5071 (N_5071,N_4915,N_4932);
or U5072 (N_5072,N_4987,N_4955);
and U5073 (N_5073,N_4908,N_4909);
or U5074 (N_5074,N_4910,N_4990);
nand U5075 (N_5075,N_4924,N_4998);
nand U5076 (N_5076,N_4981,N_4932);
and U5077 (N_5077,N_4915,N_4960);
nand U5078 (N_5078,N_4959,N_4915);
nor U5079 (N_5079,N_4925,N_4993);
nand U5080 (N_5080,N_4930,N_4995);
nor U5081 (N_5081,N_4966,N_4998);
and U5082 (N_5082,N_4925,N_4916);
or U5083 (N_5083,N_4961,N_4958);
nand U5084 (N_5084,N_4969,N_4964);
or U5085 (N_5085,N_4939,N_4906);
nand U5086 (N_5086,N_4969,N_4910);
and U5087 (N_5087,N_4987,N_4907);
nand U5088 (N_5088,N_4920,N_4927);
nand U5089 (N_5089,N_4939,N_4932);
nand U5090 (N_5090,N_4920,N_4935);
and U5091 (N_5091,N_4923,N_4979);
or U5092 (N_5092,N_4992,N_4980);
nand U5093 (N_5093,N_4966,N_4938);
or U5094 (N_5094,N_4906,N_4944);
nor U5095 (N_5095,N_4908,N_4942);
and U5096 (N_5096,N_4973,N_4950);
and U5097 (N_5097,N_4986,N_4904);
and U5098 (N_5098,N_4955,N_4975);
or U5099 (N_5099,N_4968,N_4911);
and U5100 (N_5100,N_5001,N_5060);
nand U5101 (N_5101,N_5037,N_5050);
nor U5102 (N_5102,N_5020,N_5009);
or U5103 (N_5103,N_5099,N_5012);
or U5104 (N_5104,N_5072,N_5054);
nor U5105 (N_5105,N_5021,N_5045);
nand U5106 (N_5106,N_5029,N_5011);
or U5107 (N_5107,N_5059,N_5058);
and U5108 (N_5108,N_5008,N_5097);
nand U5109 (N_5109,N_5024,N_5081);
and U5110 (N_5110,N_5073,N_5052);
nor U5111 (N_5111,N_5022,N_5023);
and U5112 (N_5112,N_5006,N_5056);
and U5113 (N_5113,N_5025,N_5080);
or U5114 (N_5114,N_5064,N_5070);
or U5115 (N_5115,N_5031,N_5047);
nor U5116 (N_5116,N_5077,N_5066);
or U5117 (N_5117,N_5017,N_5068);
and U5118 (N_5118,N_5089,N_5033);
xnor U5119 (N_5119,N_5078,N_5004);
and U5120 (N_5120,N_5085,N_5091);
or U5121 (N_5121,N_5003,N_5087);
or U5122 (N_5122,N_5018,N_5075);
or U5123 (N_5123,N_5084,N_5076);
nand U5124 (N_5124,N_5096,N_5032);
and U5125 (N_5125,N_5007,N_5049);
and U5126 (N_5126,N_5014,N_5005);
nand U5127 (N_5127,N_5048,N_5069);
nor U5128 (N_5128,N_5026,N_5061);
or U5129 (N_5129,N_5013,N_5098);
or U5130 (N_5130,N_5036,N_5035);
and U5131 (N_5131,N_5079,N_5027);
or U5132 (N_5132,N_5088,N_5057);
or U5133 (N_5133,N_5090,N_5082);
nor U5134 (N_5134,N_5038,N_5044);
and U5135 (N_5135,N_5094,N_5000);
and U5136 (N_5136,N_5034,N_5065);
and U5137 (N_5137,N_5010,N_5086);
nor U5138 (N_5138,N_5053,N_5083);
nor U5139 (N_5139,N_5095,N_5063);
and U5140 (N_5140,N_5043,N_5051);
or U5141 (N_5141,N_5030,N_5002);
or U5142 (N_5142,N_5062,N_5092);
nand U5143 (N_5143,N_5019,N_5040);
nor U5144 (N_5144,N_5093,N_5067);
nand U5145 (N_5145,N_5042,N_5055);
and U5146 (N_5146,N_5074,N_5046);
and U5147 (N_5147,N_5041,N_5028);
and U5148 (N_5148,N_5015,N_5039);
nand U5149 (N_5149,N_5016,N_5071);
and U5150 (N_5150,N_5018,N_5086);
nand U5151 (N_5151,N_5095,N_5013);
nor U5152 (N_5152,N_5074,N_5086);
or U5153 (N_5153,N_5040,N_5060);
and U5154 (N_5154,N_5061,N_5040);
or U5155 (N_5155,N_5073,N_5077);
or U5156 (N_5156,N_5000,N_5040);
nand U5157 (N_5157,N_5004,N_5089);
or U5158 (N_5158,N_5042,N_5016);
nand U5159 (N_5159,N_5014,N_5070);
and U5160 (N_5160,N_5043,N_5056);
and U5161 (N_5161,N_5037,N_5096);
or U5162 (N_5162,N_5013,N_5056);
nor U5163 (N_5163,N_5066,N_5054);
nor U5164 (N_5164,N_5054,N_5076);
and U5165 (N_5165,N_5099,N_5098);
nor U5166 (N_5166,N_5024,N_5064);
and U5167 (N_5167,N_5049,N_5040);
nor U5168 (N_5168,N_5050,N_5047);
nor U5169 (N_5169,N_5043,N_5010);
or U5170 (N_5170,N_5040,N_5005);
nand U5171 (N_5171,N_5014,N_5098);
or U5172 (N_5172,N_5091,N_5071);
nor U5173 (N_5173,N_5007,N_5066);
or U5174 (N_5174,N_5091,N_5032);
xnor U5175 (N_5175,N_5001,N_5006);
nand U5176 (N_5176,N_5004,N_5015);
and U5177 (N_5177,N_5012,N_5013);
nand U5178 (N_5178,N_5052,N_5081);
xor U5179 (N_5179,N_5072,N_5065);
nand U5180 (N_5180,N_5023,N_5004);
nand U5181 (N_5181,N_5048,N_5022);
nor U5182 (N_5182,N_5027,N_5043);
nor U5183 (N_5183,N_5015,N_5093);
or U5184 (N_5184,N_5094,N_5018);
nand U5185 (N_5185,N_5005,N_5012);
nor U5186 (N_5186,N_5074,N_5060);
nand U5187 (N_5187,N_5022,N_5033);
xor U5188 (N_5188,N_5014,N_5052);
and U5189 (N_5189,N_5096,N_5030);
xor U5190 (N_5190,N_5056,N_5090);
nor U5191 (N_5191,N_5014,N_5038);
or U5192 (N_5192,N_5051,N_5048);
nand U5193 (N_5193,N_5055,N_5009);
nor U5194 (N_5194,N_5052,N_5077);
and U5195 (N_5195,N_5047,N_5091);
nor U5196 (N_5196,N_5078,N_5074);
or U5197 (N_5197,N_5024,N_5066);
or U5198 (N_5198,N_5053,N_5064);
nand U5199 (N_5199,N_5092,N_5049);
xor U5200 (N_5200,N_5116,N_5128);
or U5201 (N_5201,N_5132,N_5137);
and U5202 (N_5202,N_5143,N_5159);
nand U5203 (N_5203,N_5169,N_5190);
nand U5204 (N_5204,N_5112,N_5161);
nor U5205 (N_5205,N_5113,N_5176);
and U5206 (N_5206,N_5171,N_5181);
or U5207 (N_5207,N_5163,N_5199);
or U5208 (N_5208,N_5157,N_5115);
nor U5209 (N_5209,N_5136,N_5119);
nand U5210 (N_5210,N_5125,N_5168);
and U5211 (N_5211,N_5158,N_5123);
nand U5212 (N_5212,N_5167,N_5110);
nor U5213 (N_5213,N_5187,N_5105);
nand U5214 (N_5214,N_5146,N_5107);
xor U5215 (N_5215,N_5152,N_5197);
and U5216 (N_5216,N_5134,N_5172);
or U5217 (N_5217,N_5196,N_5193);
and U5218 (N_5218,N_5165,N_5102);
nand U5219 (N_5219,N_5108,N_5162);
nand U5220 (N_5220,N_5147,N_5164);
or U5221 (N_5221,N_5144,N_5114);
nand U5222 (N_5222,N_5149,N_5129);
or U5223 (N_5223,N_5179,N_5145);
nor U5224 (N_5224,N_5194,N_5142);
nor U5225 (N_5225,N_5118,N_5101);
or U5226 (N_5226,N_5153,N_5109);
or U5227 (N_5227,N_5170,N_5195);
and U5228 (N_5228,N_5173,N_5138);
and U5229 (N_5229,N_5198,N_5185);
nand U5230 (N_5230,N_5126,N_5184);
and U5231 (N_5231,N_5121,N_5127);
or U5232 (N_5232,N_5156,N_5140);
nor U5233 (N_5233,N_5192,N_5141);
nor U5234 (N_5234,N_5111,N_5103);
and U5235 (N_5235,N_5148,N_5117);
nand U5236 (N_5236,N_5160,N_5100);
or U5237 (N_5237,N_5154,N_5188);
nand U5238 (N_5238,N_5191,N_5166);
nor U5239 (N_5239,N_5120,N_5174);
nand U5240 (N_5240,N_5139,N_5189);
nand U5241 (N_5241,N_5104,N_5180);
nor U5242 (N_5242,N_5131,N_5155);
or U5243 (N_5243,N_5106,N_5186);
nand U5244 (N_5244,N_5175,N_5151);
nand U5245 (N_5245,N_5133,N_5178);
nor U5246 (N_5246,N_5183,N_5135);
nand U5247 (N_5247,N_5124,N_5122);
and U5248 (N_5248,N_5177,N_5150);
and U5249 (N_5249,N_5182,N_5130);
nor U5250 (N_5250,N_5114,N_5108);
or U5251 (N_5251,N_5174,N_5125);
xor U5252 (N_5252,N_5104,N_5133);
and U5253 (N_5253,N_5103,N_5167);
or U5254 (N_5254,N_5120,N_5122);
nand U5255 (N_5255,N_5101,N_5167);
xnor U5256 (N_5256,N_5108,N_5150);
nand U5257 (N_5257,N_5191,N_5131);
nor U5258 (N_5258,N_5152,N_5143);
and U5259 (N_5259,N_5145,N_5197);
nor U5260 (N_5260,N_5104,N_5186);
and U5261 (N_5261,N_5170,N_5175);
nor U5262 (N_5262,N_5185,N_5136);
or U5263 (N_5263,N_5177,N_5154);
nand U5264 (N_5264,N_5175,N_5190);
or U5265 (N_5265,N_5113,N_5122);
nor U5266 (N_5266,N_5168,N_5179);
and U5267 (N_5267,N_5184,N_5178);
xor U5268 (N_5268,N_5130,N_5174);
nand U5269 (N_5269,N_5100,N_5188);
xnor U5270 (N_5270,N_5113,N_5197);
and U5271 (N_5271,N_5148,N_5174);
or U5272 (N_5272,N_5172,N_5166);
and U5273 (N_5273,N_5125,N_5139);
or U5274 (N_5274,N_5165,N_5138);
xnor U5275 (N_5275,N_5130,N_5151);
nor U5276 (N_5276,N_5190,N_5187);
nand U5277 (N_5277,N_5183,N_5106);
nor U5278 (N_5278,N_5120,N_5144);
and U5279 (N_5279,N_5131,N_5197);
nand U5280 (N_5280,N_5197,N_5160);
nor U5281 (N_5281,N_5172,N_5178);
nand U5282 (N_5282,N_5104,N_5199);
or U5283 (N_5283,N_5103,N_5143);
nor U5284 (N_5284,N_5147,N_5137);
and U5285 (N_5285,N_5101,N_5176);
or U5286 (N_5286,N_5125,N_5198);
or U5287 (N_5287,N_5129,N_5178);
and U5288 (N_5288,N_5129,N_5117);
or U5289 (N_5289,N_5126,N_5132);
nor U5290 (N_5290,N_5153,N_5121);
nand U5291 (N_5291,N_5151,N_5155);
nor U5292 (N_5292,N_5175,N_5140);
nand U5293 (N_5293,N_5186,N_5100);
or U5294 (N_5294,N_5111,N_5187);
or U5295 (N_5295,N_5119,N_5164);
xor U5296 (N_5296,N_5152,N_5188);
nand U5297 (N_5297,N_5120,N_5166);
nand U5298 (N_5298,N_5137,N_5193);
and U5299 (N_5299,N_5108,N_5137);
nor U5300 (N_5300,N_5236,N_5295);
or U5301 (N_5301,N_5239,N_5290);
nor U5302 (N_5302,N_5207,N_5273);
and U5303 (N_5303,N_5294,N_5251);
and U5304 (N_5304,N_5259,N_5274);
or U5305 (N_5305,N_5254,N_5269);
xor U5306 (N_5306,N_5224,N_5219);
and U5307 (N_5307,N_5291,N_5240);
nand U5308 (N_5308,N_5272,N_5264);
nand U5309 (N_5309,N_5298,N_5256);
nand U5310 (N_5310,N_5226,N_5211);
nor U5311 (N_5311,N_5262,N_5267);
nor U5312 (N_5312,N_5214,N_5292);
nand U5313 (N_5313,N_5248,N_5299);
nand U5314 (N_5314,N_5209,N_5233);
and U5315 (N_5315,N_5281,N_5201);
or U5316 (N_5316,N_5263,N_5255);
nor U5317 (N_5317,N_5205,N_5223);
nand U5318 (N_5318,N_5275,N_5268);
nand U5319 (N_5319,N_5204,N_5238);
and U5320 (N_5320,N_5210,N_5222);
nand U5321 (N_5321,N_5242,N_5297);
and U5322 (N_5322,N_5244,N_5231);
nand U5323 (N_5323,N_5202,N_5283);
nand U5324 (N_5324,N_5227,N_5237);
nand U5325 (N_5325,N_5225,N_5229);
or U5326 (N_5326,N_5252,N_5208);
nand U5327 (N_5327,N_5250,N_5279);
nand U5328 (N_5328,N_5289,N_5288);
nand U5329 (N_5329,N_5213,N_5278);
or U5330 (N_5330,N_5266,N_5203);
and U5331 (N_5331,N_5277,N_5271);
nor U5332 (N_5332,N_5232,N_5260);
or U5333 (N_5333,N_5276,N_5215);
or U5334 (N_5334,N_5245,N_5284);
nor U5335 (N_5335,N_5287,N_5206);
or U5336 (N_5336,N_5230,N_5217);
or U5337 (N_5337,N_5234,N_5228);
xnor U5338 (N_5338,N_5247,N_5221);
nor U5339 (N_5339,N_5218,N_5235);
and U5340 (N_5340,N_5249,N_5270);
nand U5341 (N_5341,N_5200,N_5282);
xor U5342 (N_5342,N_5243,N_5293);
nor U5343 (N_5343,N_5253,N_5285);
nor U5344 (N_5344,N_5286,N_5216);
nor U5345 (N_5345,N_5212,N_5257);
nand U5346 (N_5346,N_5296,N_5258);
nand U5347 (N_5347,N_5241,N_5261);
or U5348 (N_5348,N_5280,N_5220);
nand U5349 (N_5349,N_5246,N_5265);
nor U5350 (N_5350,N_5295,N_5280);
nor U5351 (N_5351,N_5299,N_5214);
nor U5352 (N_5352,N_5238,N_5220);
nor U5353 (N_5353,N_5287,N_5283);
nand U5354 (N_5354,N_5241,N_5227);
or U5355 (N_5355,N_5209,N_5225);
or U5356 (N_5356,N_5257,N_5299);
or U5357 (N_5357,N_5218,N_5264);
xnor U5358 (N_5358,N_5260,N_5280);
or U5359 (N_5359,N_5229,N_5279);
nor U5360 (N_5360,N_5200,N_5230);
xnor U5361 (N_5361,N_5219,N_5206);
and U5362 (N_5362,N_5250,N_5214);
or U5363 (N_5363,N_5251,N_5264);
and U5364 (N_5364,N_5286,N_5289);
or U5365 (N_5365,N_5271,N_5219);
and U5366 (N_5366,N_5267,N_5217);
nand U5367 (N_5367,N_5277,N_5259);
or U5368 (N_5368,N_5229,N_5299);
nor U5369 (N_5369,N_5232,N_5207);
and U5370 (N_5370,N_5273,N_5264);
or U5371 (N_5371,N_5267,N_5200);
nand U5372 (N_5372,N_5227,N_5298);
and U5373 (N_5373,N_5264,N_5206);
nand U5374 (N_5374,N_5288,N_5219);
or U5375 (N_5375,N_5201,N_5229);
nand U5376 (N_5376,N_5219,N_5222);
nor U5377 (N_5377,N_5215,N_5232);
nand U5378 (N_5378,N_5215,N_5204);
or U5379 (N_5379,N_5225,N_5217);
nand U5380 (N_5380,N_5283,N_5257);
nand U5381 (N_5381,N_5227,N_5226);
and U5382 (N_5382,N_5272,N_5275);
nor U5383 (N_5383,N_5206,N_5200);
or U5384 (N_5384,N_5200,N_5264);
or U5385 (N_5385,N_5232,N_5269);
and U5386 (N_5386,N_5264,N_5290);
or U5387 (N_5387,N_5282,N_5255);
nand U5388 (N_5388,N_5274,N_5202);
nand U5389 (N_5389,N_5274,N_5252);
nand U5390 (N_5390,N_5233,N_5294);
or U5391 (N_5391,N_5237,N_5231);
nand U5392 (N_5392,N_5217,N_5280);
nor U5393 (N_5393,N_5294,N_5220);
or U5394 (N_5394,N_5225,N_5268);
nor U5395 (N_5395,N_5277,N_5278);
nand U5396 (N_5396,N_5233,N_5234);
and U5397 (N_5397,N_5279,N_5249);
nand U5398 (N_5398,N_5271,N_5236);
or U5399 (N_5399,N_5290,N_5296);
nor U5400 (N_5400,N_5315,N_5323);
nor U5401 (N_5401,N_5345,N_5343);
nor U5402 (N_5402,N_5378,N_5399);
nor U5403 (N_5403,N_5367,N_5336);
or U5404 (N_5404,N_5317,N_5354);
nand U5405 (N_5405,N_5351,N_5330);
or U5406 (N_5406,N_5321,N_5359);
nor U5407 (N_5407,N_5381,N_5316);
and U5408 (N_5408,N_5314,N_5393);
nand U5409 (N_5409,N_5370,N_5347);
nor U5410 (N_5410,N_5320,N_5371);
or U5411 (N_5411,N_5379,N_5350);
and U5412 (N_5412,N_5349,N_5365);
nor U5413 (N_5413,N_5335,N_5332);
nand U5414 (N_5414,N_5392,N_5303);
or U5415 (N_5415,N_5374,N_5326);
nand U5416 (N_5416,N_5307,N_5355);
and U5417 (N_5417,N_5356,N_5395);
and U5418 (N_5418,N_5388,N_5384);
and U5419 (N_5419,N_5376,N_5311);
nor U5420 (N_5420,N_5305,N_5346);
and U5421 (N_5421,N_5318,N_5360);
and U5422 (N_5422,N_5310,N_5300);
or U5423 (N_5423,N_5301,N_5382);
and U5424 (N_5424,N_5362,N_5369);
nand U5425 (N_5425,N_5322,N_5380);
nand U5426 (N_5426,N_5366,N_5333);
or U5427 (N_5427,N_5302,N_5327);
nand U5428 (N_5428,N_5334,N_5397);
or U5429 (N_5429,N_5389,N_5385);
nand U5430 (N_5430,N_5308,N_5312);
and U5431 (N_5431,N_5364,N_5372);
or U5432 (N_5432,N_5339,N_5325);
or U5433 (N_5433,N_5353,N_5344);
nor U5434 (N_5434,N_5337,N_5341);
and U5435 (N_5435,N_5329,N_5377);
or U5436 (N_5436,N_5340,N_5357);
or U5437 (N_5437,N_5304,N_5373);
and U5438 (N_5438,N_5352,N_5342);
or U5439 (N_5439,N_5361,N_5313);
and U5440 (N_5440,N_5328,N_5396);
and U5441 (N_5441,N_5319,N_5383);
or U5442 (N_5442,N_5375,N_5394);
nand U5443 (N_5443,N_5391,N_5331);
nor U5444 (N_5444,N_5386,N_5387);
and U5445 (N_5445,N_5338,N_5398);
or U5446 (N_5446,N_5363,N_5358);
nand U5447 (N_5447,N_5390,N_5324);
nand U5448 (N_5448,N_5368,N_5348);
or U5449 (N_5449,N_5306,N_5309);
and U5450 (N_5450,N_5358,N_5353);
nor U5451 (N_5451,N_5334,N_5391);
nor U5452 (N_5452,N_5306,N_5314);
nor U5453 (N_5453,N_5392,N_5325);
nor U5454 (N_5454,N_5385,N_5398);
or U5455 (N_5455,N_5379,N_5305);
or U5456 (N_5456,N_5395,N_5305);
nand U5457 (N_5457,N_5331,N_5388);
nor U5458 (N_5458,N_5349,N_5363);
nor U5459 (N_5459,N_5342,N_5349);
nand U5460 (N_5460,N_5306,N_5340);
nor U5461 (N_5461,N_5385,N_5395);
nand U5462 (N_5462,N_5336,N_5317);
nor U5463 (N_5463,N_5392,N_5360);
nand U5464 (N_5464,N_5330,N_5380);
or U5465 (N_5465,N_5366,N_5337);
or U5466 (N_5466,N_5318,N_5300);
and U5467 (N_5467,N_5389,N_5359);
nor U5468 (N_5468,N_5374,N_5378);
and U5469 (N_5469,N_5318,N_5398);
or U5470 (N_5470,N_5326,N_5333);
or U5471 (N_5471,N_5365,N_5317);
and U5472 (N_5472,N_5312,N_5329);
nor U5473 (N_5473,N_5314,N_5326);
or U5474 (N_5474,N_5365,N_5371);
nand U5475 (N_5475,N_5314,N_5397);
nand U5476 (N_5476,N_5355,N_5363);
nor U5477 (N_5477,N_5390,N_5386);
or U5478 (N_5478,N_5386,N_5385);
or U5479 (N_5479,N_5320,N_5336);
nor U5480 (N_5480,N_5394,N_5382);
or U5481 (N_5481,N_5371,N_5330);
or U5482 (N_5482,N_5394,N_5360);
nand U5483 (N_5483,N_5329,N_5379);
or U5484 (N_5484,N_5321,N_5312);
nand U5485 (N_5485,N_5391,N_5392);
xnor U5486 (N_5486,N_5384,N_5355);
and U5487 (N_5487,N_5316,N_5346);
nor U5488 (N_5488,N_5351,N_5321);
xnor U5489 (N_5489,N_5369,N_5392);
or U5490 (N_5490,N_5366,N_5365);
nor U5491 (N_5491,N_5319,N_5397);
nor U5492 (N_5492,N_5301,N_5302);
and U5493 (N_5493,N_5331,N_5393);
and U5494 (N_5494,N_5372,N_5354);
nor U5495 (N_5495,N_5311,N_5375);
nand U5496 (N_5496,N_5350,N_5399);
or U5497 (N_5497,N_5322,N_5393);
and U5498 (N_5498,N_5310,N_5350);
nand U5499 (N_5499,N_5311,N_5302);
or U5500 (N_5500,N_5431,N_5474);
nor U5501 (N_5501,N_5437,N_5412);
nand U5502 (N_5502,N_5470,N_5475);
nor U5503 (N_5503,N_5442,N_5404);
nand U5504 (N_5504,N_5494,N_5425);
nor U5505 (N_5505,N_5400,N_5443);
nand U5506 (N_5506,N_5430,N_5462);
nand U5507 (N_5507,N_5478,N_5498);
nand U5508 (N_5508,N_5420,N_5441);
nand U5509 (N_5509,N_5409,N_5427);
or U5510 (N_5510,N_5445,N_5461);
nand U5511 (N_5511,N_5432,N_5444);
xnor U5512 (N_5512,N_5477,N_5439);
nand U5513 (N_5513,N_5416,N_5495);
or U5514 (N_5514,N_5429,N_5402);
or U5515 (N_5515,N_5447,N_5467);
nand U5516 (N_5516,N_5491,N_5450);
nand U5517 (N_5517,N_5496,N_5436);
or U5518 (N_5518,N_5471,N_5446);
nand U5519 (N_5519,N_5406,N_5480);
nand U5520 (N_5520,N_5497,N_5405);
nand U5521 (N_5521,N_5403,N_5401);
and U5522 (N_5522,N_5454,N_5489);
nand U5523 (N_5523,N_5458,N_5426);
nand U5524 (N_5524,N_5449,N_5499);
nor U5525 (N_5525,N_5463,N_5479);
and U5526 (N_5526,N_5423,N_5493);
and U5527 (N_5527,N_5448,N_5459);
or U5528 (N_5528,N_5457,N_5440);
nand U5529 (N_5529,N_5490,N_5408);
nor U5530 (N_5530,N_5482,N_5464);
and U5531 (N_5531,N_5452,N_5419);
nand U5532 (N_5532,N_5418,N_5483);
nand U5533 (N_5533,N_5469,N_5456);
nor U5534 (N_5534,N_5428,N_5434);
nor U5535 (N_5535,N_5460,N_5473);
or U5536 (N_5536,N_5492,N_5433);
xnor U5537 (N_5537,N_5417,N_5424);
or U5538 (N_5538,N_5485,N_5410);
nor U5539 (N_5539,N_5411,N_5472);
and U5540 (N_5540,N_5487,N_5438);
nor U5541 (N_5541,N_5481,N_5466);
nor U5542 (N_5542,N_5407,N_5476);
nand U5543 (N_5543,N_5468,N_5413);
xor U5544 (N_5544,N_5421,N_5414);
or U5545 (N_5545,N_5435,N_5451);
nand U5546 (N_5546,N_5484,N_5455);
and U5547 (N_5547,N_5486,N_5415);
nor U5548 (N_5548,N_5422,N_5453);
nand U5549 (N_5549,N_5488,N_5465);
or U5550 (N_5550,N_5413,N_5483);
nand U5551 (N_5551,N_5475,N_5454);
nor U5552 (N_5552,N_5427,N_5431);
and U5553 (N_5553,N_5424,N_5468);
or U5554 (N_5554,N_5406,N_5481);
or U5555 (N_5555,N_5478,N_5447);
nand U5556 (N_5556,N_5493,N_5459);
and U5557 (N_5557,N_5456,N_5486);
nand U5558 (N_5558,N_5461,N_5430);
nor U5559 (N_5559,N_5419,N_5464);
and U5560 (N_5560,N_5498,N_5476);
and U5561 (N_5561,N_5439,N_5445);
and U5562 (N_5562,N_5431,N_5417);
nand U5563 (N_5563,N_5403,N_5488);
nor U5564 (N_5564,N_5411,N_5487);
and U5565 (N_5565,N_5401,N_5468);
nand U5566 (N_5566,N_5442,N_5441);
nor U5567 (N_5567,N_5442,N_5496);
nor U5568 (N_5568,N_5410,N_5439);
nor U5569 (N_5569,N_5443,N_5404);
and U5570 (N_5570,N_5424,N_5483);
nor U5571 (N_5571,N_5435,N_5470);
and U5572 (N_5572,N_5435,N_5439);
nand U5573 (N_5573,N_5483,N_5441);
or U5574 (N_5574,N_5415,N_5432);
and U5575 (N_5575,N_5479,N_5433);
and U5576 (N_5576,N_5400,N_5424);
or U5577 (N_5577,N_5420,N_5448);
nor U5578 (N_5578,N_5452,N_5475);
nor U5579 (N_5579,N_5473,N_5451);
nand U5580 (N_5580,N_5414,N_5426);
and U5581 (N_5581,N_5454,N_5468);
nor U5582 (N_5582,N_5436,N_5481);
nand U5583 (N_5583,N_5466,N_5475);
and U5584 (N_5584,N_5427,N_5484);
and U5585 (N_5585,N_5414,N_5441);
or U5586 (N_5586,N_5453,N_5477);
nand U5587 (N_5587,N_5411,N_5471);
nand U5588 (N_5588,N_5487,N_5473);
or U5589 (N_5589,N_5497,N_5496);
nand U5590 (N_5590,N_5483,N_5465);
nand U5591 (N_5591,N_5466,N_5449);
nand U5592 (N_5592,N_5463,N_5407);
nand U5593 (N_5593,N_5402,N_5477);
xor U5594 (N_5594,N_5479,N_5499);
nor U5595 (N_5595,N_5432,N_5439);
nor U5596 (N_5596,N_5492,N_5429);
xor U5597 (N_5597,N_5409,N_5465);
nor U5598 (N_5598,N_5451,N_5477);
nor U5599 (N_5599,N_5416,N_5438);
or U5600 (N_5600,N_5558,N_5577);
and U5601 (N_5601,N_5508,N_5580);
xnor U5602 (N_5602,N_5599,N_5517);
nand U5603 (N_5603,N_5583,N_5516);
nand U5604 (N_5604,N_5551,N_5555);
nor U5605 (N_5605,N_5571,N_5548);
nand U5606 (N_5606,N_5523,N_5528);
nand U5607 (N_5607,N_5588,N_5511);
and U5608 (N_5608,N_5538,N_5535);
or U5609 (N_5609,N_5586,N_5527);
or U5610 (N_5610,N_5579,N_5522);
or U5611 (N_5611,N_5503,N_5539);
or U5612 (N_5612,N_5585,N_5524);
and U5613 (N_5613,N_5594,N_5595);
nor U5614 (N_5614,N_5504,N_5512);
or U5615 (N_5615,N_5540,N_5542);
and U5616 (N_5616,N_5592,N_5500);
nand U5617 (N_5617,N_5509,N_5520);
xor U5618 (N_5618,N_5566,N_5559);
or U5619 (N_5619,N_5532,N_5572);
nor U5620 (N_5620,N_5531,N_5581);
nor U5621 (N_5621,N_5590,N_5530);
and U5622 (N_5622,N_5513,N_5563);
nor U5623 (N_5623,N_5591,N_5507);
or U5624 (N_5624,N_5596,N_5575);
or U5625 (N_5625,N_5501,N_5536);
nand U5626 (N_5626,N_5560,N_5545);
nand U5627 (N_5627,N_5506,N_5514);
and U5628 (N_5628,N_5549,N_5568);
xor U5629 (N_5629,N_5510,N_5552);
or U5630 (N_5630,N_5564,N_5598);
and U5631 (N_5631,N_5561,N_5574);
and U5632 (N_5632,N_5562,N_5544);
nor U5633 (N_5633,N_5505,N_5529);
or U5634 (N_5634,N_5593,N_5573);
or U5635 (N_5635,N_5533,N_5541);
nand U5636 (N_5636,N_5578,N_5547);
and U5637 (N_5637,N_5570,N_5521);
nor U5638 (N_5638,N_5569,N_5515);
nor U5639 (N_5639,N_5543,N_5537);
nand U5640 (N_5640,N_5597,N_5546);
nand U5641 (N_5641,N_5553,N_5565);
nor U5642 (N_5642,N_5576,N_5518);
nor U5643 (N_5643,N_5550,N_5519);
or U5644 (N_5644,N_5526,N_5589);
nor U5645 (N_5645,N_5587,N_5502);
nor U5646 (N_5646,N_5557,N_5584);
and U5647 (N_5647,N_5582,N_5525);
and U5648 (N_5648,N_5567,N_5556);
and U5649 (N_5649,N_5554,N_5534);
nor U5650 (N_5650,N_5539,N_5549);
nor U5651 (N_5651,N_5526,N_5573);
or U5652 (N_5652,N_5574,N_5546);
or U5653 (N_5653,N_5547,N_5567);
xor U5654 (N_5654,N_5508,N_5579);
nand U5655 (N_5655,N_5576,N_5566);
and U5656 (N_5656,N_5543,N_5560);
nor U5657 (N_5657,N_5538,N_5565);
nor U5658 (N_5658,N_5595,N_5569);
nand U5659 (N_5659,N_5561,N_5568);
nor U5660 (N_5660,N_5554,N_5587);
or U5661 (N_5661,N_5503,N_5512);
and U5662 (N_5662,N_5517,N_5561);
nor U5663 (N_5663,N_5521,N_5507);
or U5664 (N_5664,N_5515,N_5559);
or U5665 (N_5665,N_5547,N_5559);
and U5666 (N_5666,N_5513,N_5522);
and U5667 (N_5667,N_5550,N_5561);
or U5668 (N_5668,N_5555,N_5553);
and U5669 (N_5669,N_5507,N_5548);
and U5670 (N_5670,N_5560,N_5569);
nor U5671 (N_5671,N_5512,N_5508);
or U5672 (N_5672,N_5555,N_5587);
nor U5673 (N_5673,N_5589,N_5546);
and U5674 (N_5674,N_5511,N_5543);
nor U5675 (N_5675,N_5551,N_5517);
nand U5676 (N_5676,N_5550,N_5526);
and U5677 (N_5677,N_5501,N_5555);
nor U5678 (N_5678,N_5557,N_5505);
nand U5679 (N_5679,N_5557,N_5509);
or U5680 (N_5680,N_5538,N_5591);
or U5681 (N_5681,N_5553,N_5577);
nor U5682 (N_5682,N_5542,N_5593);
nor U5683 (N_5683,N_5584,N_5574);
nand U5684 (N_5684,N_5596,N_5524);
nand U5685 (N_5685,N_5526,N_5500);
and U5686 (N_5686,N_5541,N_5511);
and U5687 (N_5687,N_5585,N_5582);
or U5688 (N_5688,N_5562,N_5516);
nor U5689 (N_5689,N_5553,N_5530);
and U5690 (N_5690,N_5587,N_5535);
or U5691 (N_5691,N_5566,N_5518);
and U5692 (N_5692,N_5573,N_5566);
xor U5693 (N_5693,N_5524,N_5567);
nor U5694 (N_5694,N_5539,N_5573);
and U5695 (N_5695,N_5542,N_5551);
nand U5696 (N_5696,N_5550,N_5590);
and U5697 (N_5697,N_5504,N_5503);
or U5698 (N_5698,N_5506,N_5561);
nand U5699 (N_5699,N_5520,N_5591);
nand U5700 (N_5700,N_5608,N_5612);
and U5701 (N_5701,N_5620,N_5637);
and U5702 (N_5702,N_5640,N_5663);
nand U5703 (N_5703,N_5668,N_5661);
nor U5704 (N_5704,N_5665,N_5646);
nand U5705 (N_5705,N_5662,N_5628);
nor U5706 (N_5706,N_5695,N_5631);
nor U5707 (N_5707,N_5658,N_5685);
nor U5708 (N_5708,N_5644,N_5659);
and U5709 (N_5709,N_5666,N_5609);
nor U5710 (N_5710,N_5642,N_5635);
nand U5711 (N_5711,N_5690,N_5625);
nand U5712 (N_5712,N_5610,N_5672);
and U5713 (N_5713,N_5657,N_5688);
and U5714 (N_5714,N_5618,N_5617);
nor U5715 (N_5715,N_5601,N_5606);
nor U5716 (N_5716,N_5675,N_5670);
and U5717 (N_5717,N_5611,N_5650);
xnor U5718 (N_5718,N_5687,N_5679);
nor U5719 (N_5719,N_5616,N_5667);
or U5720 (N_5720,N_5613,N_5673);
and U5721 (N_5721,N_5671,N_5623);
or U5722 (N_5722,N_5634,N_5632);
or U5723 (N_5723,N_5604,N_5639);
or U5724 (N_5724,N_5699,N_5697);
and U5725 (N_5725,N_5653,N_5677);
or U5726 (N_5726,N_5689,N_5615);
and U5727 (N_5727,N_5624,N_5603);
nand U5728 (N_5728,N_5643,N_5645);
nor U5729 (N_5729,N_5651,N_5605);
or U5730 (N_5730,N_5621,N_5676);
nand U5731 (N_5731,N_5664,N_5681);
nor U5732 (N_5732,N_5693,N_5619);
and U5733 (N_5733,N_5649,N_5633);
and U5734 (N_5734,N_5614,N_5683);
nand U5735 (N_5735,N_5684,N_5641);
or U5736 (N_5736,N_5674,N_5622);
nor U5737 (N_5737,N_5638,N_5652);
or U5738 (N_5738,N_5648,N_5669);
nand U5739 (N_5739,N_5680,N_5655);
or U5740 (N_5740,N_5698,N_5636);
nand U5741 (N_5741,N_5656,N_5686);
nor U5742 (N_5742,N_5696,N_5682);
and U5743 (N_5743,N_5600,N_5647);
nand U5744 (N_5744,N_5607,N_5602);
and U5745 (N_5745,N_5694,N_5630);
and U5746 (N_5746,N_5627,N_5678);
nand U5747 (N_5747,N_5660,N_5691);
nor U5748 (N_5748,N_5654,N_5626);
or U5749 (N_5749,N_5692,N_5629);
or U5750 (N_5750,N_5690,N_5676);
nor U5751 (N_5751,N_5650,N_5669);
and U5752 (N_5752,N_5657,N_5676);
and U5753 (N_5753,N_5613,N_5678);
or U5754 (N_5754,N_5634,N_5670);
nand U5755 (N_5755,N_5643,N_5619);
and U5756 (N_5756,N_5610,N_5658);
nand U5757 (N_5757,N_5672,N_5637);
or U5758 (N_5758,N_5696,N_5625);
or U5759 (N_5759,N_5691,N_5631);
or U5760 (N_5760,N_5673,N_5683);
or U5761 (N_5761,N_5634,N_5699);
nand U5762 (N_5762,N_5607,N_5697);
and U5763 (N_5763,N_5679,N_5659);
and U5764 (N_5764,N_5628,N_5660);
and U5765 (N_5765,N_5643,N_5687);
nand U5766 (N_5766,N_5695,N_5697);
and U5767 (N_5767,N_5686,N_5637);
and U5768 (N_5768,N_5606,N_5658);
and U5769 (N_5769,N_5602,N_5687);
nand U5770 (N_5770,N_5611,N_5665);
nor U5771 (N_5771,N_5695,N_5679);
or U5772 (N_5772,N_5639,N_5626);
nor U5773 (N_5773,N_5602,N_5697);
nor U5774 (N_5774,N_5694,N_5659);
and U5775 (N_5775,N_5690,N_5615);
nor U5776 (N_5776,N_5651,N_5644);
and U5777 (N_5777,N_5669,N_5619);
and U5778 (N_5778,N_5674,N_5642);
nor U5779 (N_5779,N_5602,N_5612);
and U5780 (N_5780,N_5658,N_5624);
or U5781 (N_5781,N_5672,N_5649);
nor U5782 (N_5782,N_5614,N_5604);
and U5783 (N_5783,N_5682,N_5695);
xnor U5784 (N_5784,N_5675,N_5692);
or U5785 (N_5785,N_5690,N_5687);
nand U5786 (N_5786,N_5690,N_5694);
nor U5787 (N_5787,N_5639,N_5633);
nor U5788 (N_5788,N_5648,N_5607);
nand U5789 (N_5789,N_5671,N_5641);
nor U5790 (N_5790,N_5606,N_5648);
nor U5791 (N_5791,N_5611,N_5669);
and U5792 (N_5792,N_5669,N_5642);
nand U5793 (N_5793,N_5610,N_5686);
or U5794 (N_5794,N_5632,N_5649);
nor U5795 (N_5795,N_5639,N_5615);
or U5796 (N_5796,N_5613,N_5672);
nor U5797 (N_5797,N_5664,N_5629);
and U5798 (N_5798,N_5626,N_5610);
xnor U5799 (N_5799,N_5606,N_5696);
nand U5800 (N_5800,N_5739,N_5706);
nand U5801 (N_5801,N_5757,N_5788);
or U5802 (N_5802,N_5724,N_5720);
nor U5803 (N_5803,N_5742,N_5799);
nor U5804 (N_5804,N_5755,N_5730);
or U5805 (N_5805,N_5723,N_5786);
or U5806 (N_5806,N_5728,N_5767);
nand U5807 (N_5807,N_5719,N_5778);
and U5808 (N_5808,N_5796,N_5714);
and U5809 (N_5809,N_5744,N_5798);
xnor U5810 (N_5810,N_5797,N_5743);
nor U5811 (N_5811,N_5772,N_5701);
and U5812 (N_5812,N_5762,N_5780);
or U5813 (N_5813,N_5703,N_5737);
and U5814 (N_5814,N_5771,N_5764);
or U5815 (N_5815,N_5726,N_5754);
or U5816 (N_5816,N_5727,N_5787);
nand U5817 (N_5817,N_5745,N_5702);
nor U5818 (N_5818,N_5777,N_5781);
and U5819 (N_5819,N_5741,N_5748);
nor U5820 (N_5820,N_5717,N_5752);
or U5821 (N_5821,N_5746,N_5761);
and U5822 (N_5822,N_5700,N_5793);
or U5823 (N_5823,N_5710,N_5713);
and U5824 (N_5824,N_5722,N_5791);
xnor U5825 (N_5825,N_5756,N_5709);
nand U5826 (N_5826,N_5765,N_5733);
or U5827 (N_5827,N_5750,N_5763);
and U5828 (N_5828,N_5769,N_5734);
nor U5829 (N_5829,N_5735,N_5759);
or U5830 (N_5830,N_5758,N_5747);
and U5831 (N_5831,N_5712,N_5785);
or U5832 (N_5832,N_5768,N_5775);
nand U5833 (N_5833,N_5718,N_5716);
or U5834 (N_5834,N_5736,N_5732);
and U5835 (N_5835,N_5766,N_5770);
nand U5836 (N_5836,N_5725,N_5794);
and U5837 (N_5837,N_5740,N_5721);
and U5838 (N_5838,N_5749,N_5774);
nand U5839 (N_5839,N_5753,N_5715);
or U5840 (N_5840,N_5704,N_5792);
nand U5841 (N_5841,N_5711,N_5789);
or U5842 (N_5842,N_5708,N_5795);
or U5843 (N_5843,N_5784,N_5790);
and U5844 (N_5844,N_5760,N_5783);
or U5845 (N_5845,N_5738,N_5773);
nor U5846 (N_5846,N_5705,N_5782);
nor U5847 (N_5847,N_5731,N_5776);
nor U5848 (N_5848,N_5729,N_5779);
nand U5849 (N_5849,N_5707,N_5751);
nand U5850 (N_5850,N_5774,N_5771);
or U5851 (N_5851,N_5717,N_5730);
nand U5852 (N_5852,N_5720,N_5770);
nor U5853 (N_5853,N_5778,N_5716);
nor U5854 (N_5854,N_5765,N_5759);
and U5855 (N_5855,N_5712,N_5722);
nor U5856 (N_5856,N_5755,N_5795);
nand U5857 (N_5857,N_5717,N_5759);
or U5858 (N_5858,N_5791,N_5767);
or U5859 (N_5859,N_5783,N_5737);
nor U5860 (N_5860,N_5741,N_5753);
nand U5861 (N_5861,N_5741,N_5705);
and U5862 (N_5862,N_5787,N_5757);
or U5863 (N_5863,N_5706,N_5730);
nor U5864 (N_5864,N_5733,N_5704);
nor U5865 (N_5865,N_5787,N_5764);
nand U5866 (N_5866,N_5771,N_5790);
nand U5867 (N_5867,N_5706,N_5736);
nand U5868 (N_5868,N_5775,N_5725);
nor U5869 (N_5869,N_5731,N_5757);
or U5870 (N_5870,N_5732,N_5799);
and U5871 (N_5871,N_5767,N_5788);
or U5872 (N_5872,N_5722,N_5733);
nand U5873 (N_5873,N_5766,N_5729);
or U5874 (N_5874,N_5726,N_5744);
or U5875 (N_5875,N_5788,N_5730);
or U5876 (N_5876,N_5771,N_5778);
or U5877 (N_5877,N_5742,N_5781);
and U5878 (N_5878,N_5725,N_5781);
nand U5879 (N_5879,N_5798,N_5733);
or U5880 (N_5880,N_5767,N_5710);
xnor U5881 (N_5881,N_5710,N_5756);
and U5882 (N_5882,N_5732,N_5703);
nor U5883 (N_5883,N_5767,N_5784);
and U5884 (N_5884,N_5794,N_5769);
nor U5885 (N_5885,N_5726,N_5743);
or U5886 (N_5886,N_5725,N_5730);
nor U5887 (N_5887,N_5799,N_5712);
nor U5888 (N_5888,N_5794,N_5740);
nand U5889 (N_5889,N_5724,N_5730);
nor U5890 (N_5890,N_5753,N_5793);
or U5891 (N_5891,N_5722,N_5795);
nand U5892 (N_5892,N_5777,N_5715);
or U5893 (N_5893,N_5750,N_5745);
and U5894 (N_5894,N_5799,N_5714);
or U5895 (N_5895,N_5753,N_5795);
nand U5896 (N_5896,N_5763,N_5727);
nand U5897 (N_5897,N_5775,N_5746);
nand U5898 (N_5898,N_5739,N_5723);
nor U5899 (N_5899,N_5762,N_5753);
and U5900 (N_5900,N_5845,N_5888);
xor U5901 (N_5901,N_5898,N_5881);
or U5902 (N_5902,N_5844,N_5893);
or U5903 (N_5903,N_5841,N_5816);
and U5904 (N_5904,N_5859,N_5899);
or U5905 (N_5905,N_5891,N_5812);
nor U5906 (N_5906,N_5874,N_5871);
and U5907 (N_5907,N_5896,N_5823);
or U5908 (N_5908,N_5866,N_5892);
and U5909 (N_5909,N_5811,N_5853);
nand U5910 (N_5910,N_5843,N_5822);
and U5911 (N_5911,N_5840,N_5814);
and U5912 (N_5912,N_5856,N_5826);
nor U5913 (N_5913,N_5818,N_5804);
nand U5914 (N_5914,N_5854,N_5890);
or U5915 (N_5915,N_5828,N_5837);
or U5916 (N_5916,N_5894,N_5864);
nand U5917 (N_5917,N_5813,N_5803);
or U5918 (N_5918,N_5867,N_5834);
and U5919 (N_5919,N_5865,N_5862);
and U5920 (N_5920,N_5838,N_5879);
or U5921 (N_5921,N_5877,N_5817);
nor U5922 (N_5922,N_5806,N_5831);
nor U5923 (N_5923,N_5868,N_5850);
nor U5924 (N_5924,N_5809,N_5833);
nand U5925 (N_5925,N_5882,N_5897);
nor U5926 (N_5926,N_5855,N_5861);
nand U5927 (N_5927,N_5895,N_5849);
nor U5928 (N_5928,N_5886,N_5873);
and U5929 (N_5929,N_5857,N_5870);
nor U5930 (N_5930,N_5802,N_5836);
nand U5931 (N_5931,N_5889,N_5858);
or U5932 (N_5932,N_5825,N_5805);
or U5933 (N_5933,N_5846,N_5885);
or U5934 (N_5934,N_5887,N_5875);
nor U5935 (N_5935,N_5832,N_5883);
nand U5936 (N_5936,N_5847,N_5880);
nor U5937 (N_5937,N_5869,N_5815);
nand U5938 (N_5938,N_5819,N_5839);
and U5939 (N_5939,N_5835,N_5851);
nor U5940 (N_5940,N_5827,N_5872);
and U5941 (N_5941,N_5848,N_5878);
or U5942 (N_5942,N_5863,N_5860);
and U5943 (N_5943,N_5876,N_5808);
nand U5944 (N_5944,N_5810,N_5842);
or U5945 (N_5945,N_5824,N_5830);
or U5946 (N_5946,N_5800,N_5852);
nor U5947 (N_5947,N_5820,N_5821);
nand U5948 (N_5948,N_5829,N_5807);
nor U5949 (N_5949,N_5801,N_5884);
and U5950 (N_5950,N_5800,N_5882);
nor U5951 (N_5951,N_5861,N_5811);
nand U5952 (N_5952,N_5849,N_5896);
and U5953 (N_5953,N_5863,N_5890);
and U5954 (N_5954,N_5870,N_5873);
or U5955 (N_5955,N_5876,N_5857);
xor U5956 (N_5956,N_5850,N_5870);
nand U5957 (N_5957,N_5875,N_5826);
nand U5958 (N_5958,N_5837,N_5801);
nor U5959 (N_5959,N_5896,N_5891);
and U5960 (N_5960,N_5845,N_5846);
or U5961 (N_5961,N_5886,N_5824);
and U5962 (N_5962,N_5861,N_5876);
nand U5963 (N_5963,N_5859,N_5840);
nor U5964 (N_5964,N_5807,N_5806);
nand U5965 (N_5965,N_5804,N_5806);
xnor U5966 (N_5966,N_5878,N_5821);
nor U5967 (N_5967,N_5834,N_5882);
nand U5968 (N_5968,N_5896,N_5800);
nand U5969 (N_5969,N_5874,N_5825);
nor U5970 (N_5970,N_5840,N_5800);
nor U5971 (N_5971,N_5848,N_5874);
and U5972 (N_5972,N_5888,N_5806);
and U5973 (N_5973,N_5801,N_5895);
and U5974 (N_5974,N_5866,N_5851);
nor U5975 (N_5975,N_5813,N_5882);
and U5976 (N_5976,N_5858,N_5822);
and U5977 (N_5977,N_5824,N_5872);
nand U5978 (N_5978,N_5823,N_5868);
nand U5979 (N_5979,N_5886,N_5829);
nor U5980 (N_5980,N_5875,N_5871);
nand U5981 (N_5981,N_5869,N_5810);
nor U5982 (N_5982,N_5889,N_5888);
nor U5983 (N_5983,N_5803,N_5849);
nor U5984 (N_5984,N_5807,N_5832);
nand U5985 (N_5985,N_5890,N_5889);
or U5986 (N_5986,N_5850,N_5801);
nor U5987 (N_5987,N_5846,N_5820);
nor U5988 (N_5988,N_5843,N_5812);
nor U5989 (N_5989,N_5820,N_5831);
nand U5990 (N_5990,N_5889,N_5843);
and U5991 (N_5991,N_5842,N_5892);
and U5992 (N_5992,N_5820,N_5826);
nand U5993 (N_5993,N_5893,N_5858);
nand U5994 (N_5994,N_5897,N_5898);
or U5995 (N_5995,N_5828,N_5801);
nor U5996 (N_5996,N_5873,N_5833);
and U5997 (N_5997,N_5868,N_5858);
xnor U5998 (N_5998,N_5867,N_5888);
and U5999 (N_5999,N_5847,N_5853);
nor U6000 (N_6000,N_5903,N_5994);
or U6001 (N_6001,N_5939,N_5918);
nor U6002 (N_6002,N_5986,N_5914);
nor U6003 (N_6003,N_5917,N_5909);
and U6004 (N_6004,N_5983,N_5926);
xor U6005 (N_6005,N_5971,N_5992);
nor U6006 (N_6006,N_5933,N_5974);
nor U6007 (N_6007,N_5961,N_5979);
and U6008 (N_6008,N_5934,N_5982);
nor U6009 (N_6009,N_5993,N_5964);
nand U6010 (N_6010,N_5904,N_5955);
nor U6011 (N_6011,N_5946,N_5944);
or U6012 (N_6012,N_5967,N_5991);
and U6013 (N_6013,N_5916,N_5924);
and U6014 (N_6014,N_5948,N_5911);
nor U6015 (N_6015,N_5997,N_5966);
or U6016 (N_6016,N_5998,N_5927);
or U6017 (N_6017,N_5996,N_5938);
nand U6018 (N_6018,N_5954,N_5910);
nor U6019 (N_6019,N_5935,N_5922);
and U6020 (N_6020,N_5920,N_5989);
or U6021 (N_6021,N_5969,N_5973);
nand U6022 (N_6022,N_5958,N_5932);
nor U6023 (N_6023,N_5942,N_5928);
nand U6024 (N_6024,N_5900,N_5913);
and U6025 (N_6025,N_5929,N_5941);
nand U6026 (N_6026,N_5962,N_5949);
or U6027 (N_6027,N_5923,N_5912);
nor U6028 (N_6028,N_5930,N_5978);
or U6029 (N_6029,N_5953,N_5931);
or U6030 (N_6030,N_5943,N_5907);
and U6031 (N_6031,N_5999,N_5976);
and U6032 (N_6032,N_5959,N_5950);
nor U6033 (N_6033,N_5936,N_5902);
or U6034 (N_6034,N_5901,N_5977);
nand U6035 (N_6035,N_5908,N_5951);
xnor U6036 (N_6036,N_5952,N_5970);
nor U6037 (N_6037,N_5995,N_5972);
xnor U6038 (N_6038,N_5905,N_5906);
or U6039 (N_6039,N_5965,N_5990);
and U6040 (N_6040,N_5945,N_5947);
nor U6041 (N_6041,N_5915,N_5919);
nor U6042 (N_6042,N_5988,N_5921);
and U6043 (N_6043,N_5957,N_5984);
and U6044 (N_6044,N_5937,N_5985);
nor U6045 (N_6045,N_5925,N_5956);
nand U6046 (N_6046,N_5940,N_5963);
nor U6047 (N_6047,N_5981,N_5960);
nand U6048 (N_6048,N_5987,N_5975);
nand U6049 (N_6049,N_5980,N_5968);
nor U6050 (N_6050,N_5966,N_5972);
or U6051 (N_6051,N_5996,N_5975);
nand U6052 (N_6052,N_5958,N_5987);
nor U6053 (N_6053,N_5946,N_5921);
or U6054 (N_6054,N_5921,N_5904);
nand U6055 (N_6055,N_5969,N_5901);
nand U6056 (N_6056,N_5915,N_5965);
nand U6057 (N_6057,N_5970,N_5998);
nand U6058 (N_6058,N_5964,N_5944);
or U6059 (N_6059,N_5924,N_5944);
nand U6060 (N_6060,N_5942,N_5989);
nand U6061 (N_6061,N_5923,N_5915);
or U6062 (N_6062,N_5941,N_5924);
or U6063 (N_6063,N_5940,N_5989);
nand U6064 (N_6064,N_5932,N_5972);
nand U6065 (N_6065,N_5901,N_5948);
or U6066 (N_6066,N_5916,N_5954);
and U6067 (N_6067,N_5949,N_5932);
or U6068 (N_6068,N_5982,N_5974);
nand U6069 (N_6069,N_5936,N_5994);
or U6070 (N_6070,N_5953,N_5963);
nor U6071 (N_6071,N_5980,N_5951);
nand U6072 (N_6072,N_5908,N_5939);
and U6073 (N_6073,N_5996,N_5946);
and U6074 (N_6074,N_5956,N_5946);
and U6075 (N_6075,N_5974,N_5910);
or U6076 (N_6076,N_5927,N_5976);
and U6077 (N_6077,N_5961,N_5950);
or U6078 (N_6078,N_5971,N_5945);
or U6079 (N_6079,N_5948,N_5919);
and U6080 (N_6080,N_5989,N_5936);
or U6081 (N_6081,N_5912,N_5989);
nand U6082 (N_6082,N_5968,N_5904);
nand U6083 (N_6083,N_5938,N_5993);
and U6084 (N_6084,N_5912,N_5981);
or U6085 (N_6085,N_5938,N_5971);
and U6086 (N_6086,N_5941,N_5959);
nor U6087 (N_6087,N_5946,N_5967);
nor U6088 (N_6088,N_5945,N_5973);
and U6089 (N_6089,N_5931,N_5911);
nor U6090 (N_6090,N_5907,N_5920);
and U6091 (N_6091,N_5945,N_5910);
nand U6092 (N_6092,N_5984,N_5910);
nor U6093 (N_6093,N_5907,N_5965);
nand U6094 (N_6094,N_5902,N_5922);
or U6095 (N_6095,N_5980,N_5923);
nor U6096 (N_6096,N_5936,N_5964);
nand U6097 (N_6097,N_5941,N_5931);
and U6098 (N_6098,N_5997,N_5928);
nand U6099 (N_6099,N_5943,N_5991);
nand U6100 (N_6100,N_6007,N_6022);
or U6101 (N_6101,N_6043,N_6066);
xnor U6102 (N_6102,N_6069,N_6078);
nand U6103 (N_6103,N_6077,N_6020);
nand U6104 (N_6104,N_6091,N_6097);
nand U6105 (N_6105,N_6045,N_6070);
nand U6106 (N_6106,N_6041,N_6042);
and U6107 (N_6107,N_6075,N_6008);
or U6108 (N_6108,N_6094,N_6060);
nor U6109 (N_6109,N_6010,N_6006);
or U6110 (N_6110,N_6090,N_6074);
nand U6111 (N_6111,N_6039,N_6013);
or U6112 (N_6112,N_6011,N_6062);
nor U6113 (N_6113,N_6002,N_6044);
nor U6114 (N_6114,N_6084,N_6052);
xnor U6115 (N_6115,N_6033,N_6047);
nand U6116 (N_6116,N_6086,N_6004);
nor U6117 (N_6117,N_6058,N_6083);
and U6118 (N_6118,N_6037,N_6092);
and U6119 (N_6119,N_6009,N_6036);
or U6120 (N_6120,N_6017,N_6095);
nand U6121 (N_6121,N_6067,N_6025);
nand U6122 (N_6122,N_6080,N_6024);
and U6123 (N_6123,N_6064,N_6098);
nand U6124 (N_6124,N_6087,N_6054);
nand U6125 (N_6125,N_6046,N_6056);
nand U6126 (N_6126,N_6055,N_6057);
or U6127 (N_6127,N_6034,N_6026);
nand U6128 (N_6128,N_6019,N_6021);
or U6129 (N_6129,N_6031,N_6081);
and U6130 (N_6130,N_6088,N_6003);
or U6131 (N_6131,N_6016,N_6029);
or U6132 (N_6132,N_6012,N_6030);
nand U6133 (N_6133,N_6048,N_6050);
or U6134 (N_6134,N_6051,N_6023);
or U6135 (N_6135,N_6018,N_6065);
nor U6136 (N_6136,N_6079,N_6068);
and U6137 (N_6137,N_6073,N_6015);
nor U6138 (N_6138,N_6059,N_6005);
and U6139 (N_6139,N_6049,N_6014);
xnor U6140 (N_6140,N_6038,N_6085);
nor U6141 (N_6141,N_6076,N_6040);
nand U6142 (N_6142,N_6001,N_6071);
nand U6143 (N_6143,N_6028,N_6072);
or U6144 (N_6144,N_6063,N_6096);
or U6145 (N_6145,N_6082,N_6089);
nor U6146 (N_6146,N_6027,N_6053);
xor U6147 (N_6147,N_6000,N_6093);
xor U6148 (N_6148,N_6099,N_6032);
or U6149 (N_6149,N_6035,N_6061);
and U6150 (N_6150,N_6059,N_6061);
and U6151 (N_6151,N_6012,N_6061);
nand U6152 (N_6152,N_6039,N_6084);
nand U6153 (N_6153,N_6007,N_6020);
and U6154 (N_6154,N_6003,N_6089);
nor U6155 (N_6155,N_6038,N_6013);
or U6156 (N_6156,N_6021,N_6050);
and U6157 (N_6157,N_6037,N_6024);
nand U6158 (N_6158,N_6033,N_6081);
or U6159 (N_6159,N_6039,N_6014);
or U6160 (N_6160,N_6004,N_6030);
nand U6161 (N_6161,N_6064,N_6020);
nand U6162 (N_6162,N_6049,N_6002);
or U6163 (N_6163,N_6002,N_6000);
and U6164 (N_6164,N_6032,N_6090);
or U6165 (N_6165,N_6012,N_6087);
nand U6166 (N_6166,N_6043,N_6008);
and U6167 (N_6167,N_6069,N_6068);
and U6168 (N_6168,N_6031,N_6005);
or U6169 (N_6169,N_6001,N_6084);
nand U6170 (N_6170,N_6020,N_6092);
or U6171 (N_6171,N_6092,N_6094);
nor U6172 (N_6172,N_6000,N_6092);
nor U6173 (N_6173,N_6089,N_6049);
xnor U6174 (N_6174,N_6026,N_6064);
or U6175 (N_6175,N_6038,N_6077);
and U6176 (N_6176,N_6085,N_6058);
nand U6177 (N_6177,N_6011,N_6018);
and U6178 (N_6178,N_6099,N_6015);
and U6179 (N_6179,N_6027,N_6093);
nor U6180 (N_6180,N_6036,N_6063);
and U6181 (N_6181,N_6045,N_6065);
or U6182 (N_6182,N_6036,N_6028);
nand U6183 (N_6183,N_6005,N_6029);
nand U6184 (N_6184,N_6081,N_6052);
nand U6185 (N_6185,N_6002,N_6057);
and U6186 (N_6186,N_6074,N_6001);
and U6187 (N_6187,N_6064,N_6031);
or U6188 (N_6188,N_6084,N_6029);
nor U6189 (N_6189,N_6000,N_6099);
and U6190 (N_6190,N_6086,N_6033);
nand U6191 (N_6191,N_6081,N_6028);
or U6192 (N_6192,N_6089,N_6077);
nand U6193 (N_6193,N_6037,N_6021);
xor U6194 (N_6194,N_6064,N_6067);
nand U6195 (N_6195,N_6048,N_6006);
nor U6196 (N_6196,N_6037,N_6065);
nand U6197 (N_6197,N_6049,N_6053);
nor U6198 (N_6198,N_6072,N_6089);
nand U6199 (N_6199,N_6053,N_6088);
nor U6200 (N_6200,N_6156,N_6145);
or U6201 (N_6201,N_6170,N_6104);
or U6202 (N_6202,N_6108,N_6198);
and U6203 (N_6203,N_6119,N_6162);
nor U6204 (N_6204,N_6178,N_6180);
nor U6205 (N_6205,N_6112,N_6130);
and U6206 (N_6206,N_6103,N_6191);
nand U6207 (N_6207,N_6152,N_6172);
or U6208 (N_6208,N_6185,N_6102);
and U6209 (N_6209,N_6109,N_6171);
nand U6210 (N_6210,N_6174,N_6139);
xor U6211 (N_6211,N_6136,N_6132);
nor U6212 (N_6212,N_6131,N_6150);
and U6213 (N_6213,N_6193,N_6163);
nor U6214 (N_6214,N_6110,N_6154);
nand U6215 (N_6215,N_6168,N_6125);
or U6216 (N_6216,N_6179,N_6124);
nor U6217 (N_6217,N_6142,N_6157);
nand U6218 (N_6218,N_6187,N_6114);
nand U6219 (N_6219,N_6192,N_6167);
or U6220 (N_6220,N_6149,N_6160);
or U6221 (N_6221,N_6140,N_6166);
or U6222 (N_6222,N_6107,N_6158);
nor U6223 (N_6223,N_6137,N_6115);
and U6224 (N_6224,N_6186,N_6127);
and U6225 (N_6225,N_6197,N_6173);
nor U6226 (N_6226,N_6188,N_6196);
and U6227 (N_6227,N_6117,N_6113);
nor U6228 (N_6228,N_6146,N_6181);
nor U6229 (N_6229,N_6148,N_6116);
or U6230 (N_6230,N_6147,N_6123);
nor U6231 (N_6231,N_6101,N_6161);
nor U6232 (N_6232,N_6190,N_6183);
or U6233 (N_6233,N_6169,N_6155);
and U6234 (N_6234,N_6135,N_6120);
nor U6235 (N_6235,N_6126,N_6121);
or U6236 (N_6236,N_6151,N_6111);
nor U6237 (N_6237,N_6143,N_6176);
and U6238 (N_6238,N_6175,N_6106);
or U6239 (N_6239,N_6122,N_6105);
nor U6240 (N_6240,N_6189,N_6182);
xor U6241 (N_6241,N_6128,N_6134);
nand U6242 (N_6242,N_6138,N_6194);
or U6243 (N_6243,N_6141,N_6118);
nor U6244 (N_6244,N_6195,N_6129);
nor U6245 (N_6245,N_6100,N_6159);
nand U6246 (N_6246,N_6133,N_6153);
or U6247 (N_6247,N_6164,N_6144);
nand U6248 (N_6248,N_6177,N_6199);
nor U6249 (N_6249,N_6184,N_6165);
nor U6250 (N_6250,N_6111,N_6162);
and U6251 (N_6251,N_6142,N_6131);
nor U6252 (N_6252,N_6138,N_6137);
or U6253 (N_6253,N_6121,N_6119);
and U6254 (N_6254,N_6167,N_6116);
and U6255 (N_6255,N_6196,N_6170);
nand U6256 (N_6256,N_6128,N_6166);
nor U6257 (N_6257,N_6132,N_6106);
or U6258 (N_6258,N_6191,N_6188);
nand U6259 (N_6259,N_6153,N_6143);
nand U6260 (N_6260,N_6120,N_6101);
nor U6261 (N_6261,N_6119,N_6167);
or U6262 (N_6262,N_6135,N_6150);
nand U6263 (N_6263,N_6147,N_6125);
nor U6264 (N_6264,N_6105,N_6131);
nor U6265 (N_6265,N_6108,N_6170);
or U6266 (N_6266,N_6180,N_6137);
or U6267 (N_6267,N_6184,N_6190);
nand U6268 (N_6268,N_6169,N_6115);
nor U6269 (N_6269,N_6198,N_6199);
nand U6270 (N_6270,N_6133,N_6124);
and U6271 (N_6271,N_6185,N_6167);
nand U6272 (N_6272,N_6140,N_6165);
and U6273 (N_6273,N_6179,N_6153);
nand U6274 (N_6274,N_6164,N_6180);
nor U6275 (N_6275,N_6100,N_6136);
nor U6276 (N_6276,N_6162,N_6122);
nor U6277 (N_6277,N_6120,N_6138);
and U6278 (N_6278,N_6159,N_6174);
nor U6279 (N_6279,N_6199,N_6171);
and U6280 (N_6280,N_6189,N_6137);
nor U6281 (N_6281,N_6118,N_6115);
nor U6282 (N_6282,N_6113,N_6118);
nor U6283 (N_6283,N_6186,N_6145);
or U6284 (N_6284,N_6166,N_6118);
nor U6285 (N_6285,N_6115,N_6101);
or U6286 (N_6286,N_6109,N_6161);
nor U6287 (N_6287,N_6172,N_6131);
or U6288 (N_6288,N_6196,N_6105);
or U6289 (N_6289,N_6153,N_6110);
nor U6290 (N_6290,N_6135,N_6140);
nor U6291 (N_6291,N_6190,N_6125);
or U6292 (N_6292,N_6180,N_6159);
nor U6293 (N_6293,N_6130,N_6113);
nor U6294 (N_6294,N_6124,N_6105);
and U6295 (N_6295,N_6163,N_6142);
nor U6296 (N_6296,N_6157,N_6115);
nor U6297 (N_6297,N_6172,N_6166);
nand U6298 (N_6298,N_6121,N_6133);
or U6299 (N_6299,N_6155,N_6143);
and U6300 (N_6300,N_6202,N_6241);
and U6301 (N_6301,N_6283,N_6295);
and U6302 (N_6302,N_6211,N_6227);
nor U6303 (N_6303,N_6223,N_6234);
nor U6304 (N_6304,N_6264,N_6224);
nand U6305 (N_6305,N_6204,N_6250);
and U6306 (N_6306,N_6267,N_6210);
nand U6307 (N_6307,N_6226,N_6231);
or U6308 (N_6308,N_6201,N_6261);
nand U6309 (N_6309,N_6277,N_6289);
nand U6310 (N_6310,N_6280,N_6281);
or U6311 (N_6311,N_6265,N_6240);
or U6312 (N_6312,N_6215,N_6262);
nand U6313 (N_6313,N_6249,N_6273);
or U6314 (N_6314,N_6285,N_6279);
xnor U6315 (N_6315,N_6259,N_6270);
nand U6316 (N_6316,N_6209,N_6278);
or U6317 (N_6317,N_6220,N_6213);
nand U6318 (N_6318,N_6255,N_6271);
or U6319 (N_6319,N_6291,N_6237);
nand U6320 (N_6320,N_6219,N_6256);
or U6321 (N_6321,N_6214,N_6266);
nand U6322 (N_6322,N_6290,N_6206);
or U6323 (N_6323,N_6292,N_6257);
nor U6324 (N_6324,N_6221,N_6243);
and U6325 (N_6325,N_6272,N_6247);
and U6326 (N_6326,N_6207,N_6225);
and U6327 (N_6327,N_6205,N_6244);
nand U6328 (N_6328,N_6246,N_6268);
nor U6329 (N_6329,N_6288,N_6284);
and U6330 (N_6330,N_6239,N_6293);
or U6331 (N_6331,N_6218,N_6228);
or U6332 (N_6332,N_6248,N_6296);
nor U6333 (N_6333,N_6260,N_6251);
or U6334 (N_6334,N_6269,N_6263);
nor U6335 (N_6335,N_6253,N_6203);
nor U6336 (N_6336,N_6217,N_6282);
and U6337 (N_6337,N_6252,N_6287);
and U6338 (N_6338,N_6230,N_6254);
and U6339 (N_6339,N_6229,N_6238);
nor U6340 (N_6340,N_6236,N_6294);
nand U6341 (N_6341,N_6245,N_6222);
nor U6342 (N_6342,N_6258,N_6212);
nand U6343 (N_6343,N_6200,N_6276);
or U6344 (N_6344,N_6297,N_6208);
xnor U6345 (N_6345,N_6232,N_6233);
nor U6346 (N_6346,N_6298,N_6299);
nor U6347 (N_6347,N_6216,N_6275);
nand U6348 (N_6348,N_6235,N_6286);
or U6349 (N_6349,N_6242,N_6274);
nand U6350 (N_6350,N_6247,N_6212);
nand U6351 (N_6351,N_6285,N_6209);
nor U6352 (N_6352,N_6213,N_6253);
nand U6353 (N_6353,N_6215,N_6255);
and U6354 (N_6354,N_6200,N_6296);
or U6355 (N_6355,N_6240,N_6276);
or U6356 (N_6356,N_6260,N_6211);
nand U6357 (N_6357,N_6263,N_6280);
nor U6358 (N_6358,N_6236,N_6224);
or U6359 (N_6359,N_6291,N_6219);
nor U6360 (N_6360,N_6282,N_6256);
or U6361 (N_6361,N_6228,N_6240);
nor U6362 (N_6362,N_6216,N_6239);
nand U6363 (N_6363,N_6243,N_6291);
and U6364 (N_6364,N_6279,N_6272);
nand U6365 (N_6365,N_6272,N_6257);
nor U6366 (N_6366,N_6255,N_6282);
nor U6367 (N_6367,N_6261,N_6258);
and U6368 (N_6368,N_6242,N_6280);
nand U6369 (N_6369,N_6289,N_6214);
nor U6370 (N_6370,N_6234,N_6283);
and U6371 (N_6371,N_6259,N_6280);
and U6372 (N_6372,N_6200,N_6279);
nor U6373 (N_6373,N_6276,N_6298);
or U6374 (N_6374,N_6206,N_6299);
xor U6375 (N_6375,N_6235,N_6220);
nand U6376 (N_6376,N_6299,N_6244);
or U6377 (N_6377,N_6216,N_6220);
and U6378 (N_6378,N_6214,N_6231);
nor U6379 (N_6379,N_6228,N_6297);
or U6380 (N_6380,N_6225,N_6200);
or U6381 (N_6381,N_6283,N_6217);
nand U6382 (N_6382,N_6217,N_6228);
or U6383 (N_6383,N_6207,N_6210);
nor U6384 (N_6384,N_6235,N_6240);
and U6385 (N_6385,N_6287,N_6231);
nor U6386 (N_6386,N_6221,N_6251);
nand U6387 (N_6387,N_6212,N_6223);
and U6388 (N_6388,N_6265,N_6288);
nand U6389 (N_6389,N_6291,N_6245);
or U6390 (N_6390,N_6210,N_6245);
and U6391 (N_6391,N_6221,N_6203);
nand U6392 (N_6392,N_6248,N_6209);
nand U6393 (N_6393,N_6243,N_6244);
and U6394 (N_6394,N_6285,N_6208);
and U6395 (N_6395,N_6253,N_6200);
and U6396 (N_6396,N_6206,N_6289);
and U6397 (N_6397,N_6240,N_6263);
nand U6398 (N_6398,N_6254,N_6281);
nand U6399 (N_6399,N_6212,N_6201);
nand U6400 (N_6400,N_6304,N_6380);
nor U6401 (N_6401,N_6362,N_6321);
and U6402 (N_6402,N_6342,N_6381);
or U6403 (N_6403,N_6368,N_6327);
and U6404 (N_6404,N_6371,N_6383);
nor U6405 (N_6405,N_6394,N_6303);
and U6406 (N_6406,N_6322,N_6374);
nand U6407 (N_6407,N_6388,N_6318);
and U6408 (N_6408,N_6337,N_6348);
and U6409 (N_6409,N_6328,N_6398);
or U6410 (N_6410,N_6332,N_6306);
nor U6411 (N_6411,N_6351,N_6352);
nand U6412 (N_6412,N_6338,N_6384);
nor U6413 (N_6413,N_6360,N_6320);
and U6414 (N_6414,N_6354,N_6345);
nand U6415 (N_6415,N_6323,N_6344);
and U6416 (N_6416,N_6369,N_6331);
nor U6417 (N_6417,N_6363,N_6353);
nor U6418 (N_6418,N_6308,N_6376);
nor U6419 (N_6419,N_6329,N_6390);
nor U6420 (N_6420,N_6379,N_6311);
or U6421 (N_6421,N_6377,N_6382);
and U6422 (N_6422,N_6375,N_6310);
and U6423 (N_6423,N_6370,N_6386);
and U6424 (N_6424,N_6378,N_6366);
nand U6425 (N_6425,N_6317,N_6314);
or U6426 (N_6426,N_6347,N_6300);
xor U6427 (N_6427,N_6391,N_6350);
nand U6428 (N_6428,N_6389,N_6339);
and U6429 (N_6429,N_6324,N_6349);
or U6430 (N_6430,N_6367,N_6302);
or U6431 (N_6431,N_6316,N_6373);
xor U6432 (N_6432,N_6340,N_6365);
nor U6433 (N_6433,N_6326,N_6355);
xor U6434 (N_6434,N_6361,N_6358);
or U6435 (N_6435,N_6319,N_6346);
nor U6436 (N_6436,N_6364,N_6385);
or U6437 (N_6437,N_6334,N_6313);
or U6438 (N_6438,N_6396,N_6315);
and U6439 (N_6439,N_6341,N_6343);
nand U6440 (N_6440,N_6330,N_6372);
or U6441 (N_6441,N_6301,N_6305);
or U6442 (N_6442,N_6395,N_6357);
nor U6443 (N_6443,N_6335,N_6399);
nand U6444 (N_6444,N_6359,N_6333);
and U6445 (N_6445,N_6387,N_6356);
and U6446 (N_6446,N_6392,N_6312);
or U6447 (N_6447,N_6309,N_6393);
or U6448 (N_6448,N_6336,N_6325);
nand U6449 (N_6449,N_6307,N_6397);
and U6450 (N_6450,N_6396,N_6381);
nand U6451 (N_6451,N_6320,N_6311);
nor U6452 (N_6452,N_6371,N_6342);
and U6453 (N_6453,N_6395,N_6315);
or U6454 (N_6454,N_6390,N_6373);
or U6455 (N_6455,N_6300,N_6370);
and U6456 (N_6456,N_6386,N_6324);
and U6457 (N_6457,N_6306,N_6334);
nand U6458 (N_6458,N_6342,N_6309);
and U6459 (N_6459,N_6325,N_6396);
nand U6460 (N_6460,N_6367,N_6381);
nand U6461 (N_6461,N_6311,N_6315);
or U6462 (N_6462,N_6320,N_6303);
xor U6463 (N_6463,N_6330,N_6345);
and U6464 (N_6464,N_6392,N_6313);
nor U6465 (N_6465,N_6379,N_6371);
nor U6466 (N_6466,N_6314,N_6385);
nor U6467 (N_6467,N_6346,N_6379);
or U6468 (N_6468,N_6320,N_6352);
or U6469 (N_6469,N_6367,N_6322);
nor U6470 (N_6470,N_6346,N_6301);
nor U6471 (N_6471,N_6356,N_6353);
or U6472 (N_6472,N_6396,N_6314);
nand U6473 (N_6473,N_6328,N_6390);
nand U6474 (N_6474,N_6359,N_6301);
nand U6475 (N_6475,N_6332,N_6338);
nand U6476 (N_6476,N_6386,N_6333);
nand U6477 (N_6477,N_6378,N_6384);
or U6478 (N_6478,N_6318,N_6392);
nand U6479 (N_6479,N_6307,N_6367);
nor U6480 (N_6480,N_6383,N_6328);
nor U6481 (N_6481,N_6383,N_6363);
nand U6482 (N_6482,N_6308,N_6398);
or U6483 (N_6483,N_6399,N_6336);
and U6484 (N_6484,N_6374,N_6357);
nor U6485 (N_6485,N_6309,N_6375);
nand U6486 (N_6486,N_6333,N_6317);
and U6487 (N_6487,N_6333,N_6310);
and U6488 (N_6488,N_6301,N_6334);
and U6489 (N_6489,N_6357,N_6364);
or U6490 (N_6490,N_6342,N_6398);
nand U6491 (N_6491,N_6350,N_6313);
nor U6492 (N_6492,N_6313,N_6337);
or U6493 (N_6493,N_6390,N_6321);
nor U6494 (N_6494,N_6376,N_6329);
nor U6495 (N_6495,N_6318,N_6346);
xnor U6496 (N_6496,N_6320,N_6331);
nand U6497 (N_6497,N_6305,N_6334);
and U6498 (N_6498,N_6390,N_6342);
nand U6499 (N_6499,N_6340,N_6396);
or U6500 (N_6500,N_6447,N_6455);
or U6501 (N_6501,N_6476,N_6486);
and U6502 (N_6502,N_6487,N_6414);
nor U6503 (N_6503,N_6420,N_6452);
or U6504 (N_6504,N_6475,N_6460);
and U6505 (N_6505,N_6430,N_6490);
xnor U6506 (N_6506,N_6413,N_6496);
nor U6507 (N_6507,N_6407,N_6469);
or U6508 (N_6508,N_6462,N_6438);
or U6509 (N_6509,N_6454,N_6464);
and U6510 (N_6510,N_6432,N_6449);
nand U6511 (N_6511,N_6471,N_6443);
nor U6512 (N_6512,N_6493,N_6422);
and U6513 (N_6513,N_6494,N_6474);
or U6514 (N_6514,N_6448,N_6434);
and U6515 (N_6515,N_6461,N_6488);
nor U6516 (N_6516,N_6445,N_6491);
and U6517 (N_6517,N_6457,N_6467);
nand U6518 (N_6518,N_6408,N_6427);
or U6519 (N_6519,N_6444,N_6441);
and U6520 (N_6520,N_6406,N_6463);
or U6521 (N_6521,N_6426,N_6468);
and U6522 (N_6522,N_6465,N_6489);
xnor U6523 (N_6523,N_6401,N_6410);
and U6524 (N_6524,N_6405,N_6456);
nor U6525 (N_6525,N_6425,N_6421);
nor U6526 (N_6526,N_6495,N_6412);
nand U6527 (N_6527,N_6436,N_6442);
xnor U6528 (N_6528,N_6482,N_6417);
or U6529 (N_6529,N_6453,N_6418);
or U6530 (N_6530,N_6416,N_6402);
and U6531 (N_6531,N_6484,N_6411);
or U6532 (N_6532,N_6428,N_6497);
and U6533 (N_6533,N_6450,N_6403);
or U6534 (N_6534,N_6470,N_6437);
nand U6535 (N_6535,N_6423,N_6485);
or U6536 (N_6536,N_6431,N_6459);
or U6537 (N_6537,N_6478,N_6451);
or U6538 (N_6538,N_6458,N_6415);
and U6539 (N_6539,N_6446,N_6440);
nand U6540 (N_6540,N_6481,N_6473);
nand U6541 (N_6541,N_6498,N_6433);
and U6542 (N_6542,N_6483,N_6499);
nand U6543 (N_6543,N_6477,N_6472);
nor U6544 (N_6544,N_6492,N_6479);
and U6545 (N_6545,N_6466,N_6435);
or U6546 (N_6546,N_6404,N_6480);
nor U6547 (N_6547,N_6419,N_6424);
nor U6548 (N_6548,N_6429,N_6409);
and U6549 (N_6549,N_6439,N_6400);
xor U6550 (N_6550,N_6419,N_6407);
nand U6551 (N_6551,N_6471,N_6462);
nand U6552 (N_6552,N_6490,N_6493);
or U6553 (N_6553,N_6445,N_6412);
and U6554 (N_6554,N_6453,N_6408);
nand U6555 (N_6555,N_6427,N_6450);
nor U6556 (N_6556,N_6445,N_6455);
and U6557 (N_6557,N_6492,N_6429);
nand U6558 (N_6558,N_6499,N_6452);
nor U6559 (N_6559,N_6406,N_6449);
nor U6560 (N_6560,N_6448,N_6401);
nor U6561 (N_6561,N_6441,N_6498);
or U6562 (N_6562,N_6409,N_6478);
nand U6563 (N_6563,N_6416,N_6410);
nand U6564 (N_6564,N_6418,N_6484);
or U6565 (N_6565,N_6470,N_6495);
and U6566 (N_6566,N_6470,N_6405);
nor U6567 (N_6567,N_6458,N_6474);
nand U6568 (N_6568,N_6445,N_6415);
or U6569 (N_6569,N_6407,N_6429);
nand U6570 (N_6570,N_6425,N_6409);
and U6571 (N_6571,N_6451,N_6467);
nor U6572 (N_6572,N_6406,N_6402);
and U6573 (N_6573,N_6487,N_6489);
or U6574 (N_6574,N_6479,N_6433);
nor U6575 (N_6575,N_6442,N_6437);
nor U6576 (N_6576,N_6481,N_6451);
nor U6577 (N_6577,N_6461,N_6486);
xor U6578 (N_6578,N_6406,N_6461);
and U6579 (N_6579,N_6477,N_6418);
nor U6580 (N_6580,N_6463,N_6438);
nor U6581 (N_6581,N_6402,N_6477);
nor U6582 (N_6582,N_6442,N_6477);
and U6583 (N_6583,N_6439,N_6475);
and U6584 (N_6584,N_6473,N_6459);
and U6585 (N_6585,N_6457,N_6428);
and U6586 (N_6586,N_6474,N_6472);
or U6587 (N_6587,N_6413,N_6454);
and U6588 (N_6588,N_6433,N_6429);
xnor U6589 (N_6589,N_6467,N_6498);
and U6590 (N_6590,N_6407,N_6400);
and U6591 (N_6591,N_6401,N_6483);
or U6592 (N_6592,N_6472,N_6402);
and U6593 (N_6593,N_6492,N_6440);
and U6594 (N_6594,N_6456,N_6494);
nor U6595 (N_6595,N_6418,N_6479);
nor U6596 (N_6596,N_6484,N_6447);
nand U6597 (N_6597,N_6460,N_6430);
and U6598 (N_6598,N_6405,N_6426);
and U6599 (N_6599,N_6472,N_6425);
and U6600 (N_6600,N_6550,N_6554);
nor U6601 (N_6601,N_6524,N_6586);
nor U6602 (N_6602,N_6561,N_6510);
and U6603 (N_6603,N_6577,N_6517);
and U6604 (N_6604,N_6505,N_6562);
nand U6605 (N_6605,N_6543,N_6578);
and U6606 (N_6606,N_6521,N_6572);
nor U6607 (N_6607,N_6504,N_6541);
or U6608 (N_6608,N_6575,N_6515);
or U6609 (N_6609,N_6542,N_6568);
nand U6610 (N_6610,N_6549,N_6501);
nor U6611 (N_6611,N_6584,N_6538);
or U6612 (N_6612,N_6533,N_6571);
nand U6613 (N_6613,N_6532,N_6570);
or U6614 (N_6614,N_6514,N_6518);
nor U6615 (N_6615,N_6595,N_6511);
and U6616 (N_6616,N_6523,N_6580);
nor U6617 (N_6617,N_6579,N_6583);
nor U6618 (N_6618,N_6507,N_6573);
and U6619 (N_6619,N_6547,N_6530);
and U6620 (N_6620,N_6551,N_6536);
and U6621 (N_6621,N_6512,N_6563);
nand U6622 (N_6622,N_6594,N_6588);
or U6623 (N_6623,N_6581,N_6556);
and U6624 (N_6624,N_6544,N_6548);
and U6625 (N_6625,N_6593,N_6552);
and U6626 (N_6626,N_6557,N_6566);
nand U6627 (N_6627,N_6502,N_6589);
and U6628 (N_6628,N_6585,N_6503);
nor U6629 (N_6629,N_6531,N_6587);
nor U6630 (N_6630,N_6564,N_6520);
nand U6631 (N_6631,N_6537,N_6527);
or U6632 (N_6632,N_6535,N_6553);
or U6633 (N_6633,N_6596,N_6555);
or U6634 (N_6634,N_6598,N_6558);
or U6635 (N_6635,N_6540,N_6597);
and U6636 (N_6636,N_6582,N_6576);
nor U6637 (N_6637,N_6529,N_6500);
nand U6638 (N_6638,N_6574,N_6513);
nor U6639 (N_6639,N_6539,N_6546);
or U6640 (N_6640,N_6599,N_6506);
or U6641 (N_6641,N_6560,N_6525);
nor U6642 (N_6642,N_6592,N_6545);
and U6643 (N_6643,N_6591,N_6565);
nand U6644 (N_6644,N_6590,N_6509);
nor U6645 (N_6645,N_6559,N_6528);
and U6646 (N_6646,N_6526,N_6522);
nand U6647 (N_6647,N_6534,N_6519);
nand U6648 (N_6648,N_6516,N_6567);
or U6649 (N_6649,N_6569,N_6508);
nand U6650 (N_6650,N_6552,N_6524);
nand U6651 (N_6651,N_6586,N_6554);
nor U6652 (N_6652,N_6528,N_6503);
nor U6653 (N_6653,N_6576,N_6560);
or U6654 (N_6654,N_6531,N_6537);
nor U6655 (N_6655,N_6514,N_6596);
nand U6656 (N_6656,N_6596,N_6545);
nand U6657 (N_6657,N_6597,N_6501);
and U6658 (N_6658,N_6543,N_6564);
or U6659 (N_6659,N_6511,N_6567);
and U6660 (N_6660,N_6508,N_6510);
and U6661 (N_6661,N_6569,N_6507);
or U6662 (N_6662,N_6566,N_6507);
or U6663 (N_6663,N_6520,N_6503);
and U6664 (N_6664,N_6595,N_6551);
nand U6665 (N_6665,N_6571,N_6536);
nand U6666 (N_6666,N_6593,N_6583);
or U6667 (N_6667,N_6579,N_6542);
nor U6668 (N_6668,N_6573,N_6555);
and U6669 (N_6669,N_6551,N_6590);
nand U6670 (N_6670,N_6500,N_6509);
or U6671 (N_6671,N_6547,N_6517);
nor U6672 (N_6672,N_6577,N_6569);
nand U6673 (N_6673,N_6518,N_6537);
xnor U6674 (N_6674,N_6581,N_6597);
nor U6675 (N_6675,N_6554,N_6531);
nor U6676 (N_6676,N_6562,N_6569);
and U6677 (N_6677,N_6521,N_6529);
or U6678 (N_6678,N_6516,N_6540);
or U6679 (N_6679,N_6595,N_6580);
nor U6680 (N_6680,N_6565,N_6553);
and U6681 (N_6681,N_6506,N_6586);
xor U6682 (N_6682,N_6519,N_6598);
or U6683 (N_6683,N_6505,N_6580);
and U6684 (N_6684,N_6544,N_6565);
or U6685 (N_6685,N_6568,N_6545);
nand U6686 (N_6686,N_6572,N_6539);
xor U6687 (N_6687,N_6517,N_6562);
nand U6688 (N_6688,N_6577,N_6570);
and U6689 (N_6689,N_6509,N_6545);
nor U6690 (N_6690,N_6572,N_6523);
nand U6691 (N_6691,N_6522,N_6534);
and U6692 (N_6692,N_6532,N_6503);
nand U6693 (N_6693,N_6500,N_6566);
nand U6694 (N_6694,N_6524,N_6541);
nand U6695 (N_6695,N_6573,N_6583);
and U6696 (N_6696,N_6526,N_6569);
or U6697 (N_6697,N_6539,N_6589);
or U6698 (N_6698,N_6581,N_6594);
and U6699 (N_6699,N_6572,N_6520);
nand U6700 (N_6700,N_6650,N_6627);
and U6701 (N_6701,N_6643,N_6616);
nand U6702 (N_6702,N_6651,N_6662);
nand U6703 (N_6703,N_6615,N_6665);
xnor U6704 (N_6704,N_6631,N_6669);
nor U6705 (N_6705,N_6689,N_6682);
nor U6706 (N_6706,N_6619,N_6673);
and U6707 (N_6707,N_6601,N_6604);
nor U6708 (N_6708,N_6655,N_6680);
and U6709 (N_6709,N_6690,N_6644);
and U6710 (N_6710,N_6668,N_6613);
and U6711 (N_6711,N_6639,N_6638);
nand U6712 (N_6712,N_6600,N_6624);
or U6713 (N_6713,N_6633,N_6617);
and U6714 (N_6714,N_6664,N_6612);
or U6715 (N_6715,N_6646,N_6609);
nand U6716 (N_6716,N_6610,N_6687);
nor U6717 (N_6717,N_6675,N_6681);
nor U6718 (N_6718,N_6611,N_6648);
or U6719 (N_6719,N_6694,N_6686);
and U6720 (N_6720,N_6658,N_6623);
nor U6721 (N_6721,N_6636,N_6630);
nand U6722 (N_6722,N_6625,N_6659);
nand U6723 (N_6723,N_6663,N_6618);
nor U6724 (N_6724,N_6637,N_6641);
and U6725 (N_6725,N_6672,N_6670);
nor U6726 (N_6726,N_6674,N_6621);
nor U6727 (N_6727,N_6653,N_6602);
nor U6728 (N_6728,N_6628,N_6649);
nor U6729 (N_6729,N_6608,N_6677);
or U6730 (N_6730,N_6645,N_6695);
nor U6731 (N_6731,N_6642,N_6685);
nor U6732 (N_6732,N_6676,N_6699);
xor U6733 (N_6733,N_6647,N_6660);
nor U6734 (N_6734,N_6698,N_6693);
nor U6735 (N_6735,N_6684,N_6683);
or U6736 (N_6736,N_6688,N_6661);
and U6737 (N_6737,N_6657,N_6679);
and U6738 (N_6738,N_6696,N_6605);
xor U6739 (N_6739,N_6667,N_6671);
or U6740 (N_6740,N_6614,N_6697);
and U6741 (N_6741,N_6678,N_6629);
or U6742 (N_6742,N_6603,N_6632);
and U6743 (N_6743,N_6640,N_6634);
nor U6744 (N_6744,N_6622,N_6691);
and U6745 (N_6745,N_6607,N_6666);
nor U6746 (N_6746,N_6620,N_6654);
or U6747 (N_6747,N_6656,N_6635);
and U6748 (N_6748,N_6652,N_6606);
nand U6749 (N_6749,N_6692,N_6626);
nand U6750 (N_6750,N_6674,N_6664);
nand U6751 (N_6751,N_6656,N_6665);
nor U6752 (N_6752,N_6643,N_6665);
or U6753 (N_6753,N_6680,N_6684);
nor U6754 (N_6754,N_6677,N_6655);
nand U6755 (N_6755,N_6682,N_6652);
and U6756 (N_6756,N_6607,N_6684);
and U6757 (N_6757,N_6697,N_6628);
or U6758 (N_6758,N_6614,N_6619);
or U6759 (N_6759,N_6670,N_6659);
and U6760 (N_6760,N_6699,N_6615);
xor U6761 (N_6761,N_6659,N_6689);
or U6762 (N_6762,N_6623,N_6606);
or U6763 (N_6763,N_6634,N_6645);
or U6764 (N_6764,N_6664,N_6628);
nor U6765 (N_6765,N_6680,N_6600);
or U6766 (N_6766,N_6674,N_6660);
or U6767 (N_6767,N_6633,N_6634);
nor U6768 (N_6768,N_6677,N_6631);
nand U6769 (N_6769,N_6648,N_6601);
nand U6770 (N_6770,N_6604,N_6603);
nand U6771 (N_6771,N_6685,N_6657);
nor U6772 (N_6772,N_6636,N_6690);
and U6773 (N_6773,N_6617,N_6603);
or U6774 (N_6774,N_6601,N_6640);
xnor U6775 (N_6775,N_6673,N_6624);
and U6776 (N_6776,N_6626,N_6670);
nand U6777 (N_6777,N_6628,N_6652);
nor U6778 (N_6778,N_6665,N_6616);
nand U6779 (N_6779,N_6605,N_6692);
nor U6780 (N_6780,N_6677,N_6635);
nand U6781 (N_6781,N_6660,N_6685);
and U6782 (N_6782,N_6622,N_6610);
nor U6783 (N_6783,N_6627,N_6678);
nand U6784 (N_6784,N_6614,N_6652);
or U6785 (N_6785,N_6688,N_6600);
or U6786 (N_6786,N_6667,N_6668);
and U6787 (N_6787,N_6612,N_6682);
nor U6788 (N_6788,N_6655,N_6679);
nor U6789 (N_6789,N_6646,N_6656);
or U6790 (N_6790,N_6684,N_6687);
and U6791 (N_6791,N_6667,N_6646);
and U6792 (N_6792,N_6648,N_6636);
or U6793 (N_6793,N_6626,N_6646);
nand U6794 (N_6794,N_6616,N_6695);
and U6795 (N_6795,N_6694,N_6676);
and U6796 (N_6796,N_6657,N_6607);
and U6797 (N_6797,N_6628,N_6640);
nor U6798 (N_6798,N_6690,N_6616);
or U6799 (N_6799,N_6674,N_6676);
nor U6800 (N_6800,N_6724,N_6796);
nand U6801 (N_6801,N_6789,N_6766);
nor U6802 (N_6802,N_6786,N_6744);
nor U6803 (N_6803,N_6706,N_6708);
or U6804 (N_6804,N_6787,N_6751);
nand U6805 (N_6805,N_6714,N_6713);
and U6806 (N_6806,N_6700,N_6718);
nor U6807 (N_6807,N_6747,N_6758);
or U6808 (N_6808,N_6716,N_6755);
or U6809 (N_6809,N_6793,N_6749);
and U6810 (N_6810,N_6703,N_6738);
nor U6811 (N_6811,N_6710,N_6733);
xnor U6812 (N_6812,N_6788,N_6792);
or U6813 (N_6813,N_6798,N_6791);
or U6814 (N_6814,N_6702,N_6799);
and U6815 (N_6815,N_6748,N_6753);
and U6816 (N_6816,N_6754,N_6771);
nand U6817 (N_6817,N_6770,N_6774);
nand U6818 (N_6818,N_6775,N_6757);
nand U6819 (N_6819,N_6723,N_6720);
or U6820 (N_6820,N_6735,N_6722);
nor U6821 (N_6821,N_6780,N_6727);
xnor U6822 (N_6822,N_6704,N_6750);
nand U6823 (N_6823,N_6797,N_6762);
and U6824 (N_6824,N_6709,N_6705);
or U6825 (N_6825,N_6779,N_6730);
or U6826 (N_6826,N_6739,N_6728);
nor U6827 (N_6827,N_6778,N_6781);
nand U6828 (N_6828,N_6729,N_6701);
or U6829 (N_6829,N_6785,N_6794);
and U6830 (N_6830,N_6717,N_6736);
and U6831 (N_6831,N_6726,N_6712);
nand U6832 (N_6832,N_6719,N_6764);
or U6833 (N_6833,N_6740,N_6763);
or U6834 (N_6834,N_6795,N_6761);
nand U6835 (N_6835,N_6711,N_6743);
and U6836 (N_6836,N_6732,N_6741);
nor U6837 (N_6837,N_6777,N_6760);
xnor U6838 (N_6838,N_6725,N_6756);
nand U6839 (N_6839,N_6784,N_6742);
nand U6840 (N_6840,N_6768,N_6783);
or U6841 (N_6841,N_6759,N_6790);
nand U6842 (N_6842,N_6776,N_6737);
nand U6843 (N_6843,N_6731,N_6746);
nor U6844 (N_6844,N_6721,N_6782);
and U6845 (N_6845,N_6715,N_6765);
nor U6846 (N_6846,N_6769,N_6745);
or U6847 (N_6847,N_6773,N_6772);
nand U6848 (N_6848,N_6707,N_6734);
and U6849 (N_6849,N_6767,N_6752);
nand U6850 (N_6850,N_6753,N_6723);
nor U6851 (N_6851,N_6756,N_6783);
and U6852 (N_6852,N_6741,N_6761);
and U6853 (N_6853,N_6773,N_6797);
nand U6854 (N_6854,N_6760,N_6763);
nor U6855 (N_6855,N_6719,N_6726);
and U6856 (N_6856,N_6742,N_6704);
nand U6857 (N_6857,N_6780,N_6790);
nand U6858 (N_6858,N_6769,N_6792);
nand U6859 (N_6859,N_6784,N_6703);
and U6860 (N_6860,N_6704,N_6795);
nand U6861 (N_6861,N_6710,N_6712);
nor U6862 (N_6862,N_6726,N_6772);
nor U6863 (N_6863,N_6736,N_6787);
nand U6864 (N_6864,N_6742,N_6746);
nand U6865 (N_6865,N_6737,N_6775);
nand U6866 (N_6866,N_6709,N_6736);
nor U6867 (N_6867,N_6706,N_6758);
and U6868 (N_6868,N_6725,N_6787);
and U6869 (N_6869,N_6751,N_6718);
nand U6870 (N_6870,N_6795,N_6705);
xor U6871 (N_6871,N_6793,N_6781);
or U6872 (N_6872,N_6743,N_6727);
or U6873 (N_6873,N_6772,N_6756);
or U6874 (N_6874,N_6745,N_6743);
nor U6875 (N_6875,N_6707,N_6766);
nand U6876 (N_6876,N_6768,N_6754);
or U6877 (N_6877,N_6771,N_6746);
nor U6878 (N_6878,N_6726,N_6703);
nand U6879 (N_6879,N_6730,N_6764);
nand U6880 (N_6880,N_6740,N_6755);
nand U6881 (N_6881,N_6790,N_6729);
nor U6882 (N_6882,N_6710,N_6752);
nand U6883 (N_6883,N_6764,N_6775);
nand U6884 (N_6884,N_6740,N_6733);
nor U6885 (N_6885,N_6767,N_6797);
or U6886 (N_6886,N_6731,N_6762);
or U6887 (N_6887,N_6793,N_6731);
and U6888 (N_6888,N_6715,N_6793);
and U6889 (N_6889,N_6769,N_6710);
nand U6890 (N_6890,N_6737,N_6725);
nor U6891 (N_6891,N_6733,N_6707);
nor U6892 (N_6892,N_6727,N_6768);
and U6893 (N_6893,N_6738,N_6782);
nor U6894 (N_6894,N_6739,N_6704);
or U6895 (N_6895,N_6737,N_6793);
nor U6896 (N_6896,N_6707,N_6701);
and U6897 (N_6897,N_6787,N_6705);
nor U6898 (N_6898,N_6746,N_6758);
or U6899 (N_6899,N_6752,N_6782);
nor U6900 (N_6900,N_6854,N_6874);
or U6901 (N_6901,N_6897,N_6822);
or U6902 (N_6902,N_6823,N_6868);
and U6903 (N_6903,N_6809,N_6817);
nor U6904 (N_6904,N_6880,N_6812);
xor U6905 (N_6905,N_6820,N_6856);
and U6906 (N_6906,N_6850,N_6834);
or U6907 (N_6907,N_6845,N_6846);
nand U6908 (N_6908,N_6882,N_6804);
nand U6909 (N_6909,N_6848,N_6884);
or U6910 (N_6910,N_6832,N_6819);
nand U6911 (N_6911,N_6890,N_6801);
nor U6912 (N_6912,N_6835,N_6885);
and U6913 (N_6913,N_6878,N_6840);
nor U6914 (N_6914,N_6838,N_6826);
and U6915 (N_6915,N_6870,N_6827);
nor U6916 (N_6916,N_6810,N_6857);
nor U6917 (N_6917,N_6816,N_6841);
and U6918 (N_6918,N_6866,N_6876);
nand U6919 (N_6919,N_6807,N_6886);
nor U6920 (N_6920,N_6881,N_6844);
and U6921 (N_6921,N_6824,N_6864);
or U6922 (N_6922,N_6843,N_6862);
nand U6923 (N_6923,N_6806,N_6847);
and U6924 (N_6924,N_6836,N_6825);
and U6925 (N_6925,N_6828,N_6893);
nand U6926 (N_6926,N_6839,N_6800);
nor U6927 (N_6927,N_6851,N_6852);
and U6928 (N_6928,N_6860,N_6891);
nand U6929 (N_6929,N_6814,N_6802);
or U6930 (N_6930,N_6858,N_6899);
nand U6931 (N_6931,N_6811,N_6875);
nor U6932 (N_6932,N_6895,N_6829);
or U6933 (N_6933,N_6873,N_6813);
and U6934 (N_6934,N_6821,N_6888);
nand U6935 (N_6935,N_6805,N_6833);
nor U6936 (N_6936,N_6867,N_6892);
or U6937 (N_6937,N_6883,N_6898);
and U6938 (N_6938,N_6853,N_6877);
nor U6939 (N_6939,N_6879,N_6871);
nand U6940 (N_6940,N_6855,N_6894);
nand U6941 (N_6941,N_6872,N_6889);
and U6942 (N_6942,N_6803,N_6815);
nor U6943 (N_6943,N_6831,N_6837);
xor U6944 (N_6944,N_6865,N_6849);
or U6945 (N_6945,N_6863,N_6859);
nand U6946 (N_6946,N_6869,N_6896);
nand U6947 (N_6947,N_6830,N_6887);
and U6948 (N_6948,N_6861,N_6842);
and U6949 (N_6949,N_6818,N_6808);
or U6950 (N_6950,N_6849,N_6871);
nand U6951 (N_6951,N_6867,N_6881);
nor U6952 (N_6952,N_6839,N_6867);
and U6953 (N_6953,N_6872,N_6859);
nor U6954 (N_6954,N_6832,N_6867);
and U6955 (N_6955,N_6847,N_6864);
nor U6956 (N_6956,N_6836,N_6868);
and U6957 (N_6957,N_6864,N_6817);
or U6958 (N_6958,N_6815,N_6882);
and U6959 (N_6959,N_6801,N_6867);
or U6960 (N_6960,N_6845,N_6813);
xor U6961 (N_6961,N_6865,N_6853);
and U6962 (N_6962,N_6880,N_6848);
nand U6963 (N_6963,N_6894,N_6810);
and U6964 (N_6964,N_6852,N_6868);
and U6965 (N_6965,N_6892,N_6858);
and U6966 (N_6966,N_6891,N_6809);
nor U6967 (N_6967,N_6819,N_6891);
nand U6968 (N_6968,N_6898,N_6800);
or U6969 (N_6969,N_6875,N_6883);
and U6970 (N_6970,N_6852,N_6862);
nand U6971 (N_6971,N_6840,N_6830);
nor U6972 (N_6972,N_6836,N_6802);
or U6973 (N_6973,N_6871,N_6823);
or U6974 (N_6974,N_6829,N_6807);
nand U6975 (N_6975,N_6863,N_6896);
and U6976 (N_6976,N_6834,N_6831);
nand U6977 (N_6977,N_6875,N_6837);
nand U6978 (N_6978,N_6809,N_6842);
and U6979 (N_6979,N_6871,N_6858);
and U6980 (N_6980,N_6885,N_6800);
nor U6981 (N_6981,N_6869,N_6881);
nor U6982 (N_6982,N_6824,N_6871);
nor U6983 (N_6983,N_6859,N_6804);
or U6984 (N_6984,N_6801,N_6887);
nor U6985 (N_6985,N_6851,N_6801);
xor U6986 (N_6986,N_6855,N_6803);
nor U6987 (N_6987,N_6849,N_6840);
and U6988 (N_6988,N_6855,N_6887);
or U6989 (N_6989,N_6891,N_6864);
or U6990 (N_6990,N_6831,N_6892);
nor U6991 (N_6991,N_6827,N_6892);
or U6992 (N_6992,N_6803,N_6841);
and U6993 (N_6993,N_6848,N_6823);
or U6994 (N_6994,N_6831,N_6898);
or U6995 (N_6995,N_6836,N_6806);
nor U6996 (N_6996,N_6806,N_6834);
and U6997 (N_6997,N_6833,N_6886);
and U6998 (N_6998,N_6888,N_6898);
nor U6999 (N_6999,N_6856,N_6899);
and U7000 (N_7000,N_6941,N_6998);
nand U7001 (N_7001,N_6936,N_6937);
nand U7002 (N_7002,N_6984,N_6963);
or U7003 (N_7003,N_6950,N_6932);
nor U7004 (N_7004,N_6991,N_6913);
or U7005 (N_7005,N_6933,N_6988);
nand U7006 (N_7006,N_6951,N_6902);
or U7007 (N_7007,N_6931,N_6993);
nand U7008 (N_7008,N_6957,N_6904);
or U7009 (N_7009,N_6939,N_6920);
and U7010 (N_7010,N_6956,N_6995);
and U7011 (N_7011,N_6918,N_6960);
and U7012 (N_7012,N_6911,N_6949);
nor U7013 (N_7013,N_6938,N_6966);
nand U7014 (N_7014,N_6926,N_6952);
nor U7015 (N_7015,N_6935,N_6953);
and U7016 (N_7016,N_6983,N_6955);
or U7017 (N_7017,N_6934,N_6996);
and U7018 (N_7018,N_6948,N_6974);
nand U7019 (N_7019,N_6980,N_6946);
and U7020 (N_7020,N_6917,N_6973);
or U7021 (N_7021,N_6916,N_6962);
nor U7022 (N_7022,N_6999,N_6914);
nor U7023 (N_7023,N_6922,N_6985);
and U7024 (N_7024,N_6900,N_6987);
nand U7025 (N_7025,N_6901,N_6986);
nor U7026 (N_7026,N_6997,N_6942);
xor U7027 (N_7027,N_6964,N_6958);
xor U7028 (N_7028,N_6924,N_6903);
and U7029 (N_7029,N_6943,N_6954);
nor U7030 (N_7030,N_6940,N_6965);
nand U7031 (N_7031,N_6994,N_6947);
nor U7032 (N_7032,N_6977,N_6961);
and U7033 (N_7033,N_6989,N_6990);
or U7034 (N_7034,N_6908,N_6929);
nor U7035 (N_7035,N_6930,N_6928);
and U7036 (N_7036,N_6907,N_6915);
or U7037 (N_7037,N_6978,N_6981);
or U7038 (N_7038,N_6905,N_6910);
nor U7039 (N_7039,N_6982,N_6959);
nor U7040 (N_7040,N_6944,N_6923);
nand U7041 (N_7041,N_6979,N_6912);
or U7042 (N_7042,N_6975,N_6921);
and U7043 (N_7043,N_6992,N_6976);
and U7044 (N_7044,N_6909,N_6970);
nand U7045 (N_7045,N_6971,N_6972);
nor U7046 (N_7046,N_6927,N_6906);
nand U7047 (N_7047,N_6925,N_6945);
or U7048 (N_7048,N_6968,N_6969);
nand U7049 (N_7049,N_6919,N_6967);
nand U7050 (N_7050,N_6971,N_6941);
nand U7051 (N_7051,N_6968,N_6911);
nor U7052 (N_7052,N_6964,N_6944);
nand U7053 (N_7053,N_6969,N_6961);
and U7054 (N_7054,N_6904,N_6990);
nand U7055 (N_7055,N_6981,N_6996);
or U7056 (N_7056,N_6946,N_6935);
and U7057 (N_7057,N_6950,N_6997);
or U7058 (N_7058,N_6925,N_6908);
nand U7059 (N_7059,N_6965,N_6951);
xnor U7060 (N_7060,N_6992,N_6902);
or U7061 (N_7061,N_6969,N_6988);
nor U7062 (N_7062,N_6929,N_6981);
or U7063 (N_7063,N_6945,N_6982);
or U7064 (N_7064,N_6931,N_6917);
or U7065 (N_7065,N_6966,N_6942);
or U7066 (N_7066,N_6932,N_6955);
nand U7067 (N_7067,N_6977,N_6968);
nor U7068 (N_7068,N_6916,N_6910);
or U7069 (N_7069,N_6920,N_6999);
and U7070 (N_7070,N_6942,N_6958);
and U7071 (N_7071,N_6915,N_6974);
nand U7072 (N_7072,N_6951,N_6937);
nand U7073 (N_7073,N_6918,N_6927);
nor U7074 (N_7074,N_6945,N_6921);
and U7075 (N_7075,N_6976,N_6972);
or U7076 (N_7076,N_6914,N_6911);
nor U7077 (N_7077,N_6939,N_6906);
and U7078 (N_7078,N_6919,N_6954);
and U7079 (N_7079,N_6922,N_6977);
and U7080 (N_7080,N_6957,N_6926);
nor U7081 (N_7081,N_6992,N_6930);
nand U7082 (N_7082,N_6981,N_6907);
nor U7083 (N_7083,N_6939,N_6903);
or U7084 (N_7084,N_6979,N_6969);
nand U7085 (N_7085,N_6993,N_6988);
or U7086 (N_7086,N_6956,N_6902);
and U7087 (N_7087,N_6990,N_6902);
or U7088 (N_7088,N_6994,N_6997);
nand U7089 (N_7089,N_6940,N_6921);
and U7090 (N_7090,N_6960,N_6907);
nand U7091 (N_7091,N_6924,N_6905);
nand U7092 (N_7092,N_6913,N_6976);
or U7093 (N_7093,N_6985,N_6982);
or U7094 (N_7094,N_6971,N_6929);
or U7095 (N_7095,N_6948,N_6979);
or U7096 (N_7096,N_6916,N_6936);
nor U7097 (N_7097,N_6997,N_6944);
or U7098 (N_7098,N_6952,N_6966);
and U7099 (N_7099,N_6951,N_6921);
nor U7100 (N_7100,N_7023,N_7079);
nor U7101 (N_7101,N_7027,N_7063);
or U7102 (N_7102,N_7041,N_7059);
and U7103 (N_7103,N_7009,N_7095);
nor U7104 (N_7104,N_7008,N_7058);
and U7105 (N_7105,N_7048,N_7025);
or U7106 (N_7106,N_7033,N_7078);
and U7107 (N_7107,N_7034,N_7030);
and U7108 (N_7108,N_7050,N_7091);
nand U7109 (N_7109,N_7031,N_7022);
and U7110 (N_7110,N_7013,N_7011);
nor U7111 (N_7111,N_7044,N_7068);
nor U7112 (N_7112,N_7045,N_7056);
nand U7113 (N_7113,N_7037,N_7075);
nand U7114 (N_7114,N_7010,N_7081);
xnor U7115 (N_7115,N_7051,N_7060);
and U7116 (N_7116,N_7040,N_7019);
and U7117 (N_7117,N_7085,N_7087);
or U7118 (N_7118,N_7067,N_7001);
or U7119 (N_7119,N_7003,N_7089);
nand U7120 (N_7120,N_7053,N_7005);
nand U7121 (N_7121,N_7097,N_7086);
nor U7122 (N_7122,N_7052,N_7099);
nor U7123 (N_7123,N_7038,N_7055);
nand U7124 (N_7124,N_7083,N_7065);
nand U7125 (N_7125,N_7029,N_7049);
nor U7126 (N_7126,N_7096,N_7039);
nor U7127 (N_7127,N_7006,N_7054);
and U7128 (N_7128,N_7093,N_7046);
and U7129 (N_7129,N_7074,N_7021);
or U7130 (N_7130,N_7017,N_7026);
or U7131 (N_7131,N_7012,N_7072);
or U7132 (N_7132,N_7036,N_7077);
nand U7133 (N_7133,N_7062,N_7066);
nand U7134 (N_7134,N_7064,N_7002);
nor U7135 (N_7135,N_7080,N_7007);
or U7136 (N_7136,N_7047,N_7057);
nand U7137 (N_7137,N_7014,N_7042);
or U7138 (N_7138,N_7016,N_7032);
nor U7139 (N_7139,N_7018,N_7024);
and U7140 (N_7140,N_7071,N_7084);
nand U7141 (N_7141,N_7076,N_7094);
or U7142 (N_7142,N_7000,N_7043);
nor U7143 (N_7143,N_7020,N_7015);
and U7144 (N_7144,N_7090,N_7028);
or U7145 (N_7145,N_7070,N_7069);
and U7146 (N_7146,N_7004,N_7082);
nand U7147 (N_7147,N_7098,N_7035);
nand U7148 (N_7148,N_7073,N_7088);
nand U7149 (N_7149,N_7061,N_7092);
or U7150 (N_7150,N_7025,N_7076);
or U7151 (N_7151,N_7072,N_7013);
and U7152 (N_7152,N_7084,N_7072);
nand U7153 (N_7153,N_7080,N_7021);
nor U7154 (N_7154,N_7053,N_7031);
nand U7155 (N_7155,N_7037,N_7011);
nor U7156 (N_7156,N_7050,N_7066);
xor U7157 (N_7157,N_7016,N_7010);
or U7158 (N_7158,N_7095,N_7043);
and U7159 (N_7159,N_7095,N_7033);
and U7160 (N_7160,N_7077,N_7008);
and U7161 (N_7161,N_7077,N_7025);
or U7162 (N_7162,N_7027,N_7086);
nor U7163 (N_7163,N_7003,N_7070);
nand U7164 (N_7164,N_7059,N_7067);
or U7165 (N_7165,N_7085,N_7091);
and U7166 (N_7166,N_7070,N_7096);
nor U7167 (N_7167,N_7093,N_7073);
and U7168 (N_7168,N_7011,N_7090);
nor U7169 (N_7169,N_7089,N_7042);
and U7170 (N_7170,N_7082,N_7090);
and U7171 (N_7171,N_7023,N_7074);
and U7172 (N_7172,N_7071,N_7034);
or U7173 (N_7173,N_7017,N_7020);
nor U7174 (N_7174,N_7021,N_7055);
nand U7175 (N_7175,N_7064,N_7011);
and U7176 (N_7176,N_7034,N_7047);
xnor U7177 (N_7177,N_7057,N_7056);
nor U7178 (N_7178,N_7080,N_7020);
and U7179 (N_7179,N_7099,N_7089);
nor U7180 (N_7180,N_7084,N_7096);
nand U7181 (N_7181,N_7022,N_7070);
nor U7182 (N_7182,N_7034,N_7077);
or U7183 (N_7183,N_7065,N_7098);
nor U7184 (N_7184,N_7058,N_7057);
or U7185 (N_7185,N_7076,N_7056);
nand U7186 (N_7186,N_7062,N_7048);
and U7187 (N_7187,N_7093,N_7036);
and U7188 (N_7188,N_7056,N_7008);
and U7189 (N_7189,N_7080,N_7073);
nor U7190 (N_7190,N_7008,N_7085);
nor U7191 (N_7191,N_7056,N_7064);
and U7192 (N_7192,N_7020,N_7057);
or U7193 (N_7193,N_7032,N_7061);
nor U7194 (N_7194,N_7008,N_7054);
and U7195 (N_7195,N_7041,N_7080);
nor U7196 (N_7196,N_7092,N_7089);
nand U7197 (N_7197,N_7061,N_7008);
nor U7198 (N_7198,N_7085,N_7076);
and U7199 (N_7199,N_7073,N_7065);
and U7200 (N_7200,N_7136,N_7148);
nor U7201 (N_7201,N_7181,N_7170);
nor U7202 (N_7202,N_7116,N_7128);
or U7203 (N_7203,N_7168,N_7156);
nor U7204 (N_7204,N_7121,N_7154);
and U7205 (N_7205,N_7171,N_7146);
nand U7206 (N_7206,N_7125,N_7197);
or U7207 (N_7207,N_7142,N_7118);
or U7208 (N_7208,N_7175,N_7179);
nor U7209 (N_7209,N_7195,N_7133);
nand U7210 (N_7210,N_7132,N_7131);
or U7211 (N_7211,N_7180,N_7176);
and U7212 (N_7212,N_7111,N_7137);
or U7213 (N_7213,N_7196,N_7143);
and U7214 (N_7214,N_7126,N_7151);
or U7215 (N_7215,N_7110,N_7161);
nand U7216 (N_7216,N_7117,N_7124);
nand U7217 (N_7217,N_7188,N_7104);
nor U7218 (N_7218,N_7177,N_7193);
nor U7219 (N_7219,N_7192,N_7119);
or U7220 (N_7220,N_7178,N_7160);
nand U7221 (N_7221,N_7157,N_7108);
nor U7222 (N_7222,N_7144,N_7190);
and U7223 (N_7223,N_7138,N_7194);
nand U7224 (N_7224,N_7182,N_7165);
nor U7225 (N_7225,N_7127,N_7172);
or U7226 (N_7226,N_7198,N_7103);
nor U7227 (N_7227,N_7189,N_7149);
nor U7228 (N_7228,N_7139,N_7153);
or U7229 (N_7229,N_7134,N_7141);
and U7230 (N_7230,N_7164,N_7166);
or U7231 (N_7231,N_7129,N_7169);
or U7232 (N_7232,N_7167,N_7122);
or U7233 (N_7233,N_7107,N_7102);
and U7234 (N_7234,N_7163,N_7187);
or U7235 (N_7235,N_7174,N_7101);
nor U7236 (N_7236,N_7150,N_7186);
nor U7237 (N_7237,N_7109,N_7158);
nor U7238 (N_7238,N_7120,N_7113);
nand U7239 (N_7239,N_7115,N_7147);
and U7240 (N_7240,N_7191,N_7185);
or U7241 (N_7241,N_7105,N_7106);
nand U7242 (N_7242,N_7159,N_7183);
nand U7243 (N_7243,N_7135,N_7100);
or U7244 (N_7244,N_7140,N_7152);
and U7245 (N_7245,N_7199,N_7155);
and U7246 (N_7246,N_7173,N_7162);
and U7247 (N_7247,N_7145,N_7130);
nand U7248 (N_7248,N_7112,N_7114);
or U7249 (N_7249,N_7184,N_7123);
or U7250 (N_7250,N_7174,N_7162);
and U7251 (N_7251,N_7180,N_7103);
nor U7252 (N_7252,N_7136,N_7126);
nor U7253 (N_7253,N_7124,N_7145);
nor U7254 (N_7254,N_7118,N_7190);
nor U7255 (N_7255,N_7176,N_7110);
or U7256 (N_7256,N_7197,N_7168);
nor U7257 (N_7257,N_7165,N_7109);
nand U7258 (N_7258,N_7138,N_7173);
and U7259 (N_7259,N_7163,N_7128);
or U7260 (N_7260,N_7145,N_7151);
nor U7261 (N_7261,N_7134,N_7166);
nor U7262 (N_7262,N_7136,N_7101);
nor U7263 (N_7263,N_7144,N_7159);
nor U7264 (N_7264,N_7199,N_7141);
nor U7265 (N_7265,N_7191,N_7128);
or U7266 (N_7266,N_7192,N_7112);
and U7267 (N_7267,N_7129,N_7175);
xor U7268 (N_7268,N_7186,N_7195);
or U7269 (N_7269,N_7110,N_7111);
and U7270 (N_7270,N_7105,N_7169);
nor U7271 (N_7271,N_7107,N_7164);
nand U7272 (N_7272,N_7129,N_7184);
nand U7273 (N_7273,N_7183,N_7192);
nor U7274 (N_7274,N_7165,N_7128);
or U7275 (N_7275,N_7136,N_7172);
nor U7276 (N_7276,N_7168,N_7190);
or U7277 (N_7277,N_7129,N_7158);
and U7278 (N_7278,N_7149,N_7118);
nand U7279 (N_7279,N_7173,N_7109);
and U7280 (N_7280,N_7113,N_7161);
or U7281 (N_7281,N_7137,N_7166);
xor U7282 (N_7282,N_7199,N_7100);
nand U7283 (N_7283,N_7164,N_7199);
nor U7284 (N_7284,N_7183,N_7123);
or U7285 (N_7285,N_7108,N_7190);
and U7286 (N_7286,N_7117,N_7126);
nand U7287 (N_7287,N_7165,N_7169);
and U7288 (N_7288,N_7154,N_7149);
and U7289 (N_7289,N_7102,N_7105);
or U7290 (N_7290,N_7125,N_7104);
nor U7291 (N_7291,N_7149,N_7171);
or U7292 (N_7292,N_7179,N_7116);
and U7293 (N_7293,N_7104,N_7141);
or U7294 (N_7294,N_7136,N_7157);
and U7295 (N_7295,N_7143,N_7138);
and U7296 (N_7296,N_7109,N_7170);
xor U7297 (N_7297,N_7182,N_7104);
and U7298 (N_7298,N_7185,N_7140);
and U7299 (N_7299,N_7143,N_7105);
nand U7300 (N_7300,N_7256,N_7248);
or U7301 (N_7301,N_7290,N_7230);
nand U7302 (N_7302,N_7298,N_7215);
nand U7303 (N_7303,N_7260,N_7209);
or U7304 (N_7304,N_7272,N_7224);
nor U7305 (N_7305,N_7287,N_7271);
nor U7306 (N_7306,N_7258,N_7235);
xnor U7307 (N_7307,N_7255,N_7210);
nor U7308 (N_7308,N_7237,N_7242);
and U7309 (N_7309,N_7202,N_7220);
and U7310 (N_7310,N_7231,N_7219);
and U7311 (N_7311,N_7251,N_7232);
nand U7312 (N_7312,N_7234,N_7229);
and U7313 (N_7313,N_7236,N_7291);
nor U7314 (N_7314,N_7212,N_7216);
nor U7315 (N_7315,N_7223,N_7240);
nand U7316 (N_7316,N_7203,N_7250);
nor U7317 (N_7317,N_7285,N_7201);
nor U7318 (N_7318,N_7281,N_7275);
xor U7319 (N_7319,N_7208,N_7293);
nor U7320 (N_7320,N_7211,N_7283);
and U7321 (N_7321,N_7282,N_7217);
and U7322 (N_7322,N_7280,N_7245);
nand U7323 (N_7323,N_7213,N_7222);
or U7324 (N_7324,N_7253,N_7277);
nand U7325 (N_7325,N_7257,N_7269);
nor U7326 (N_7326,N_7259,N_7284);
and U7327 (N_7327,N_7205,N_7266);
nor U7328 (N_7328,N_7292,N_7296);
nor U7329 (N_7329,N_7226,N_7276);
or U7330 (N_7330,N_7244,N_7264);
nor U7331 (N_7331,N_7238,N_7214);
and U7332 (N_7332,N_7288,N_7261);
nand U7333 (N_7333,N_7206,N_7289);
nor U7334 (N_7334,N_7297,N_7274);
nand U7335 (N_7335,N_7286,N_7279);
and U7336 (N_7336,N_7204,N_7262);
or U7337 (N_7337,N_7241,N_7294);
nor U7338 (N_7338,N_7200,N_7239);
xor U7339 (N_7339,N_7273,N_7295);
nand U7340 (N_7340,N_7268,N_7265);
and U7341 (N_7341,N_7218,N_7247);
nand U7342 (N_7342,N_7233,N_7299);
nor U7343 (N_7343,N_7263,N_7267);
or U7344 (N_7344,N_7278,N_7227);
nand U7345 (N_7345,N_7249,N_7228);
and U7346 (N_7346,N_7246,N_7243);
nor U7347 (N_7347,N_7270,N_7221);
and U7348 (N_7348,N_7254,N_7207);
nor U7349 (N_7349,N_7225,N_7252);
and U7350 (N_7350,N_7246,N_7286);
nor U7351 (N_7351,N_7206,N_7287);
and U7352 (N_7352,N_7234,N_7295);
xor U7353 (N_7353,N_7263,N_7272);
nor U7354 (N_7354,N_7298,N_7201);
nor U7355 (N_7355,N_7200,N_7264);
and U7356 (N_7356,N_7204,N_7297);
nor U7357 (N_7357,N_7220,N_7245);
nand U7358 (N_7358,N_7218,N_7217);
and U7359 (N_7359,N_7218,N_7200);
nand U7360 (N_7360,N_7289,N_7281);
and U7361 (N_7361,N_7240,N_7262);
nor U7362 (N_7362,N_7234,N_7245);
or U7363 (N_7363,N_7220,N_7230);
xnor U7364 (N_7364,N_7205,N_7217);
xor U7365 (N_7365,N_7230,N_7226);
nand U7366 (N_7366,N_7233,N_7236);
nand U7367 (N_7367,N_7271,N_7262);
and U7368 (N_7368,N_7234,N_7232);
or U7369 (N_7369,N_7237,N_7212);
and U7370 (N_7370,N_7208,N_7277);
nor U7371 (N_7371,N_7215,N_7267);
or U7372 (N_7372,N_7202,N_7264);
and U7373 (N_7373,N_7206,N_7286);
nor U7374 (N_7374,N_7280,N_7253);
and U7375 (N_7375,N_7262,N_7265);
and U7376 (N_7376,N_7204,N_7263);
or U7377 (N_7377,N_7268,N_7295);
nor U7378 (N_7378,N_7285,N_7205);
and U7379 (N_7379,N_7208,N_7264);
or U7380 (N_7380,N_7257,N_7274);
nor U7381 (N_7381,N_7210,N_7226);
nor U7382 (N_7382,N_7286,N_7218);
nor U7383 (N_7383,N_7298,N_7251);
nor U7384 (N_7384,N_7299,N_7214);
or U7385 (N_7385,N_7206,N_7260);
nor U7386 (N_7386,N_7223,N_7281);
and U7387 (N_7387,N_7234,N_7217);
or U7388 (N_7388,N_7260,N_7283);
and U7389 (N_7389,N_7298,N_7211);
nor U7390 (N_7390,N_7281,N_7273);
nor U7391 (N_7391,N_7292,N_7250);
and U7392 (N_7392,N_7248,N_7271);
nor U7393 (N_7393,N_7215,N_7229);
or U7394 (N_7394,N_7241,N_7286);
nand U7395 (N_7395,N_7288,N_7249);
nand U7396 (N_7396,N_7271,N_7224);
and U7397 (N_7397,N_7238,N_7224);
and U7398 (N_7398,N_7209,N_7201);
nand U7399 (N_7399,N_7291,N_7208);
and U7400 (N_7400,N_7370,N_7309);
or U7401 (N_7401,N_7364,N_7352);
nor U7402 (N_7402,N_7382,N_7327);
and U7403 (N_7403,N_7312,N_7373);
nand U7404 (N_7404,N_7383,N_7391);
nor U7405 (N_7405,N_7399,N_7323);
nand U7406 (N_7406,N_7300,N_7339);
or U7407 (N_7407,N_7390,N_7308);
nand U7408 (N_7408,N_7392,N_7303);
nor U7409 (N_7409,N_7398,N_7318);
or U7410 (N_7410,N_7344,N_7397);
and U7411 (N_7411,N_7386,N_7395);
and U7412 (N_7412,N_7307,N_7359);
nand U7413 (N_7413,N_7372,N_7378);
nor U7414 (N_7414,N_7356,N_7369);
or U7415 (N_7415,N_7363,N_7351);
and U7416 (N_7416,N_7388,N_7320);
or U7417 (N_7417,N_7367,N_7336);
nor U7418 (N_7418,N_7314,N_7346);
xor U7419 (N_7419,N_7313,N_7380);
nand U7420 (N_7420,N_7304,N_7325);
nand U7421 (N_7421,N_7358,N_7368);
or U7422 (N_7422,N_7328,N_7357);
or U7423 (N_7423,N_7396,N_7324);
and U7424 (N_7424,N_7384,N_7353);
nor U7425 (N_7425,N_7393,N_7330);
or U7426 (N_7426,N_7377,N_7333);
and U7427 (N_7427,N_7354,N_7317);
and U7428 (N_7428,N_7301,N_7311);
xnor U7429 (N_7429,N_7387,N_7350);
or U7430 (N_7430,N_7326,N_7341);
or U7431 (N_7431,N_7376,N_7319);
nor U7432 (N_7432,N_7332,N_7322);
nor U7433 (N_7433,N_7316,N_7348);
or U7434 (N_7434,N_7305,N_7375);
nand U7435 (N_7435,N_7335,N_7343);
or U7436 (N_7436,N_7389,N_7349);
xor U7437 (N_7437,N_7362,N_7365);
nand U7438 (N_7438,N_7381,N_7315);
and U7439 (N_7439,N_7337,N_7385);
nand U7440 (N_7440,N_7329,N_7302);
nand U7441 (N_7441,N_7340,N_7334);
or U7442 (N_7442,N_7374,N_7338);
and U7443 (N_7443,N_7306,N_7321);
or U7444 (N_7444,N_7361,N_7355);
nor U7445 (N_7445,N_7394,N_7371);
nand U7446 (N_7446,N_7360,N_7345);
nor U7447 (N_7447,N_7342,N_7379);
or U7448 (N_7448,N_7310,N_7347);
nor U7449 (N_7449,N_7331,N_7366);
nor U7450 (N_7450,N_7392,N_7323);
nor U7451 (N_7451,N_7328,N_7396);
nor U7452 (N_7452,N_7378,N_7356);
and U7453 (N_7453,N_7395,N_7306);
or U7454 (N_7454,N_7302,N_7306);
or U7455 (N_7455,N_7376,N_7344);
or U7456 (N_7456,N_7327,N_7332);
or U7457 (N_7457,N_7331,N_7392);
and U7458 (N_7458,N_7346,N_7399);
nor U7459 (N_7459,N_7354,N_7342);
nand U7460 (N_7460,N_7350,N_7330);
or U7461 (N_7461,N_7339,N_7345);
nand U7462 (N_7462,N_7319,N_7373);
or U7463 (N_7463,N_7382,N_7307);
nor U7464 (N_7464,N_7320,N_7357);
nand U7465 (N_7465,N_7325,N_7374);
nand U7466 (N_7466,N_7322,N_7323);
and U7467 (N_7467,N_7334,N_7380);
or U7468 (N_7468,N_7376,N_7304);
nand U7469 (N_7469,N_7300,N_7326);
nor U7470 (N_7470,N_7397,N_7307);
nor U7471 (N_7471,N_7323,N_7356);
nand U7472 (N_7472,N_7385,N_7391);
nor U7473 (N_7473,N_7351,N_7374);
nand U7474 (N_7474,N_7369,N_7377);
or U7475 (N_7475,N_7370,N_7349);
nand U7476 (N_7476,N_7385,N_7327);
and U7477 (N_7477,N_7377,N_7316);
nor U7478 (N_7478,N_7390,N_7338);
and U7479 (N_7479,N_7328,N_7391);
nor U7480 (N_7480,N_7366,N_7354);
nand U7481 (N_7481,N_7340,N_7369);
or U7482 (N_7482,N_7333,N_7371);
and U7483 (N_7483,N_7342,N_7333);
nand U7484 (N_7484,N_7331,N_7319);
and U7485 (N_7485,N_7348,N_7392);
and U7486 (N_7486,N_7392,N_7334);
nor U7487 (N_7487,N_7374,N_7352);
and U7488 (N_7488,N_7313,N_7309);
or U7489 (N_7489,N_7389,N_7370);
nand U7490 (N_7490,N_7332,N_7376);
nor U7491 (N_7491,N_7324,N_7368);
or U7492 (N_7492,N_7389,N_7367);
and U7493 (N_7493,N_7361,N_7388);
and U7494 (N_7494,N_7344,N_7335);
nand U7495 (N_7495,N_7320,N_7374);
or U7496 (N_7496,N_7371,N_7349);
and U7497 (N_7497,N_7300,N_7384);
nor U7498 (N_7498,N_7338,N_7384);
nor U7499 (N_7499,N_7380,N_7316);
and U7500 (N_7500,N_7454,N_7449);
nand U7501 (N_7501,N_7417,N_7444);
or U7502 (N_7502,N_7463,N_7441);
or U7503 (N_7503,N_7496,N_7411);
nor U7504 (N_7504,N_7421,N_7495);
nand U7505 (N_7505,N_7403,N_7446);
nand U7506 (N_7506,N_7480,N_7431);
and U7507 (N_7507,N_7475,N_7465);
and U7508 (N_7508,N_7445,N_7426);
nor U7509 (N_7509,N_7456,N_7453);
nor U7510 (N_7510,N_7455,N_7481);
nor U7511 (N_7511,N_7405,N_7418);
nor U7512 (N_7512,N_7439,N_7408);
or U7513 (N_7513,N_7435,N_7482);
nor U7514 (N_7514,N_7400,N_7416);
and U7515 (N_7515,N_7451,N_7477);
or U7516 (N_7516,N_7459,N_7457);
nor U7517 (N_7517,N_7499,N_7448);
or U7518 (N_7518,N_7437,N_7409);
nor U7519 (N_7519,N_7497,N_7429);
xnor U7520 (N_7520,N_7420,N_7461);
or U7521 (N_7521,N_7402,N_7489);
or U7522 (N_7522,N_7438,N_7413);
nand U7523 (N_7523,N_7494,N_7423);
nand U7524 (N_7524,N_7466,N_7460);
and U7525 (N_7525,N_7412,N_7490);
nor U7526 (N_7526,N_7478,N_7406);
or U7527 (N_7527,N_7487,N_7471);
nor U7528 (N_7528,N_7458,N_7474);
or U7529 (N_7529,N_7440,N_7469);
and U7530 (N_7530,N_7419,N_7436);
and U7531 (N_7531,N_7468,N_7433);
nand U7532 (N_7532,N_7410,N_7467);
or U7533 (N_7533,N_7483,N_7486);
and U7534 (N_7534,N_7424,N_7452);
nand U7535 (N_7535,N_7447,N_7414);
and U7536 (N_7536,N_7491,N_7427);
xnor U7537 (N_7537,N_7462,N_7498);
nand U7538 (N_7538,N_7428,N_7479);
or U7539 (N_7539,N_7432,N_7443);
nand U7540 (N_7540,N_7473,N_7464);
nand U7541 (N_7541,N_7434,N_7430);
nor U7542 (N_7542,N_7415,N_7422);
and U7543 (N_7543,N_7485,N_7476);
nand U7544 (N_7544,N_7442,N_7401);
nand U7545 (N_7545,N_7492,N_7493);
nor U7546 (N_7546,N_7450,N_7404);
and U7547 (N_7547,N_7484,N_7488);
nor U7548 (N_7548,N_7470,N_7407);
or U7549 (N_7549,N_7472,N_7425);
nand U7550 (N_7550,N_7455,N_7441);
and U7551 (N_7551,N_7402,N_7405);
nor U7552 (N_7552,N_7417,N_7411);
or U7553 (N_7553,N_7445,N_7496);
nand U7554 (N_7554,N_7481,N_7488);
and U7555 (N_7555,N_7468,N_7467);
nand U7556 (N_7556,N_7432,N_7404);
nand U7557 (N_7557,N_7479,N_7419);
and U7558 (N_7558,N_7456,N_7488);
or U7559 (N_7559,N_7461,N_7428);
or U7560 (N_7560,N_7415,N_7405);
or U7561 (N_7561,N_7436,N_7463);
or U7562 (N_7562,N_7408,N_7467);
xnor U7563 (N_7563,N_7463,N_7415);
xnor U7564 (N_7564,N_7499,N_7438);
and U7565 (N_7565,N_7474,N_7416);
or U7566 (N_7566,N_7401,N_7460);
or U7567 (N_7567,N_7494,N_7438);
nand U7568 (N_7568,N_7499,N_7429);
nor U7569 (N_7569,N_7478,N_7405);
nand U7570 (N_7570,N_7488,N_7434);
and U7571 (N_7571,N_7406,N_7494);
and U7572 (N_7572,N_7469,N_7413);
or U7573 (N_7573,N_7452,N_7402);
nand U7574 (N_7574,N_7465,N_7408);
nor U7575 (N_7575,N_7441,N_7451);
or U7576 (N_7576,N_7405,N_7449);
nor U7577 (N_7577,N_7466,N_7441);
and U7578 (N_7578,N_7406,N_7499);
or U7579 (N_7579,N_7439,N_7443);
or U7580 (N_7580,N_7474,N_7432);
and U7581 (N_7581,N_7441,N_7495);
and U7582 (N_7582,N_7446,N_7479);
and U7583 (N_7583,N_7459,N_7497);
and U7584 (N_7584,N_7439,N_7488);
and U7585 (N_7585,N_7400,N_7479);
or U7586 (N_7586,N_7467,N_7401);
nand U7587 (N_7587,N_7432,N_7400);
and U7588 (N_7588,N_7438,N_7485);
and U7589 (N_7589,N_7413,N_7489);
and U7590 (N_7590,N_7426,N_7474);
nor U7591 (N_7591,N_7447,N_7488);
or U7592 (N_7592,N_7493,N_7445);
nor U7593 (N_7593,N_7417,N_7434);
and U7594 (N_7594,N_7490,N_7457);
or U7595 (N_7595,N_7468,N_7409);
and U7596 (N_7596,N_7411,N_7463);
or U7597 (N_7597,N_7480,N_7495);
and U7598 (N_7598,N_7454,N_7411);
or U7599 (N_7599,N_7484,N_7424);
nand U7600 (N_7600,N_7555,N_7590);
xnor U7601 (N_7601,N_7575,N_7554);
and U7602 (N_7602,N_7568,N_7581);
and U7603 (N_7603,N_7599,N_7551);
nor U7604 (N_7604,N_7566,N_7538);
and U7605 (N_7605,N_7597,N_7531);
xor U7606 (N_7606,N_7539,N_7580);
or U7607 (N_7607,N_7571,N_7572);
and U7608 (N_7608,N_7574,N_7549);
and U7609 (N_7609,N_7537,N_7507);
and U7610 (N_7610,N_7548,N_7529);
nor U7611 (N_7611,N_7552,N_7545);
nand U7612 (N_7612,N_7559,N_7542);
nor U7613 (N_7613,N_7594,N_7584);
nor U7614 (N_7614,N_7520,N_7522);
nand U7615 (N_7615,N_7585,N_7513);
and U7616 (N_7616,N_7583,N_7596);
nor U7617 (N_7617,N_7514,N_7503);
nor U7618 (N_7618,N_7533,N_7563);
and U7619 (N_7619,N_7587,N_7561);
and U7620 (N_7620,N_7527,N_7576);
nand U7621 (N_7621,N_7534,N_7540);
or U7622 (N_7622,N_7504,N_7565);
and U7623 (N_7623,N_7501,N_7598);
nand U7624 (N_7624,N_7591,N_7567);
nand U7625 (N_7625,N_7579,N_7578);
or U7626 (N_7626,N_7560,N_7500);
nand U7627 (N_7627,N_7506,N_7556);
xor U7628 (N_7628,N_7516,N_7511);
or U7629 (N_7629,N_7586,N_7592);
and U7630 (N_7630,N_7508,N_7577);
nor U7631 (N_7631,N_7562,N_7593);
nor U7632 (N_7632,N_7564,N_7570);
and U7633 (N_7633,N_7558,N_7589);
or U7634 (N_7634,N_7523,N_7582);
and U7635 (N_7635,N_7510,N_7536);
and U7636 (N_7636,N_7546,N_7550);
nand U7637 (N_7637,N_7569,N_7518);
nand U7638 (N_7638,N_7573,N_7521);
nand U7639 (N_7639,N_7532,N_7588);
nor U7640 (N_7640,N_7595,N_7544);
or U7641 (N_7641,N_7530,N_7517);
nor U7642 (N_7642,N_7509,N_7553);
nand U7643 (N_7643,N_7515,N_7543);
and U7644 (N_7644,N_7541,N_7505);
and U7645 (N_7645,N_7512,N_7524);
nor U7646 (N_7646,N_7519,N_7535);
or U7647 (N_7647,N_7525,N_7526);
and U7648 (N_7648,N_7502,N_7557);
nand U7649 (N_7649,N_7528,N_7547);
and U7650 (N_7650,N_7572,N_7525);
nand U7651 (N_7651,N_7533,N_7578);
nand U7652 (N_7652,N_7508,N_7559);
or U7653 (N_7653,N_7556,N_7542);
nand U7654 (N_7654,N_7507,N_7571);
and U7655 (N_7655,N_7582,N_7507);
nand U7656 (N_7656,N_7552,N_7535);
or U7657 (N_7657,N_7571,N_7519);
or U7658 (N_7658,N_7539,N_7583);
nand U7659 (N_7659,N_7558,N_7521);
and U7660 (N_7660,N_7523,N_7567);
and U7661 (N_7661,N_7565,N_7560);
or U7662 (N_7662,N_7549,N_7540);
xor U7663 (N_7663,N_7540,N_7584);
and U7664 (N_7664,N_7507,N_7520);
or U7665 (N_7665,N_7531,N_7510);
nand U7666 (N_7666,N_7525,N_7522);
or U7667 (N_7667,N_7505,N_7512);
nor U7668 (N_7668,N_7552,N_7558);
and U7669 (N_7669,N_7513,N_7576);
xnor U7670 (N_7670,N_7507,N_7517);
nand U7671 (N_7671,N_7561,N_7504);
or U7672 (N_7672,N_7573,N_7502);
nor U7673 (N_7673,N_7506,N_7588);
or U7674 (N_7674,N_7565,N_7507);
and U7675 (N_7675,N_7587,N_7595);
nor U7676 (N_7676,N_7533,N_7501);
and U7677 (N_7677,N_7566,N_7536);
and U7678 (N_7678,N_7583,N_7570);
or U7679 (N_7679,N_7530,N_7519);
or U7680 (N_7680,N_7567,N_7559);
nand U7681 (N_7681,N_7598,N_7525);
and U7682 (N_7682,N_7510,N_7503);
nor U7683 (N_7683,N_7572,N_7595);
nand U7684 (N_7684,N_7509,N_7542);
or U7685 (N_7685,N_7544,N_7555);
nand U7686 (N_7686,N_7596,N_7511);
nand U7687 (N_7687,N_7534,N_7589);
nor U7688 (N_7688,N_7564,N_7550);
or U7689 (N_7689,N_7528,N_7503);
nand U7690 (N_7690,N_7576,N_7580);
nor U7691 (N_7691,N_7504,N_7508);
nand U7692 (N_7692,N_7547,N_7511);
and U7693 (N_7693,N_7574,N_7569);
and U7694 (N_7694,N_7567,N_7589);
nor U7695 (N_7695,N_7595,N_7511);
and U7696 (N_7696,N_7517,N_7585);
or U7697 (N_7697,N_7534,N_7570);
nand U7698 (N_7698,N_7520,N_7550);
and U7699 (N_7699,N_7578,N_7513);
xor U7700 (N_7700,N_7698,N_7617);
nand U7701 (N_7701,N_7647,N_7613);
nor U7702 (N_7702,N_7662,N_7699);
nand U7703 (N_7703,N_7656,N_7689);
or U7704 (N_7704,N_7653,N_7674);
and U7705 (N_7705,N_7646,N_7667);
and U7706 (N_7706,N_7641,N_7692);
or U7707 (N_7707,N_7635,N_7649);
and U7708 (N_7708,N_7658,N_7680);
nand U7709 (N_7709,N_7648,N_7611);
nor U7710 (N_7710,N_7672,N_7614);
nor U7711 (N_7711,N_7675,N_7664);
nand U7712 (N_7712,N_7620,N_7661);
or U7713 (N_7713,N_7626,N_7612);
and U7714 (N_7714,N_7631,N_7695);
and U7715 (N_7715,N_7687,N_7696);
or U7716 (N_7716,N_7655,N_7616);
nor U7717 (N_7717,N_7642,N_7634);
nor U7718 (N_7718,N_7679,N_7624);
and U7719 (N_7719,N_7683,N_7666);
nor U7720 (N_7720,N_7619,N_7629);
nand U7721 (N_7721,N_7607,N_7645);
or U7722 (N_7722,N_7632,N_7684);
and U7723 (N_7723,N_7618,N_7682);
nand U7724 (N_7724,N_7676,N_7660);
and U7725 (N_7725,N_7638,N_7671);
nor U7726 (N_7726,N_7633,N_7650);
nand U7727 (N_7727,N_7690,N_7665);
or U7728 (N_7728,N_7673,N_7615);
and U7729 (N_7729,N_7601,N_7693);
xor U7730 (N_7730,N_7640,N_7694);
and U7731 (N_7731,N_7621,N_7605);
nor U7732 (N_7732,N_7670,N_7677);
nor U7733 (N_7733,N_7681,N_7657);
or U7734 (N_7734,N_7669,N_7609);
nand U7735 (N_7735,N_7623,N_7636);
and U7736 (N_7736,N_7685,N_7688);
nand U7737 (N_7737,N_7608,N_7686);
and U7738 (N_7738,N_7622,N_7600);
nand U7739 (N_7739,N_7625,N_7630);
nor U7740 (N_7740,N_7643,N_7652);
and U7741 (N_7741,N_7668,N_7637);
xnor U7742 (N_7742,N_7663,N_7678);
and U7743 (N_7743,N_7603,N_7697);
nand U7744 (N_7744,N_7659,N_7654);
nand U7745 (N_7745,N_7610,N_7627);
or U7746 (N_7746,N_7628,N_7644);
or U7747 (N_7747,N_7651,N_7606);
nor U7748 (N_7748,N_7602,N_7604);
and U7749 (N_7749,N_7691,N_7639);
nand U7750 (N_7750,N_7628,N_7665);
and U7751 (N_7751,N_7607,N_7697);
nor U7752 (N_7752,N_7617,N_7691);
and U7753 (N_7753,N_7648,N_7616);
nand U7754 (N_7754,N_7614,N_7698);
or U7755 (N_7755,N_7647,N_7621);
nor U7756 (N_7756,N_7627,N_7681);
and U7757 (N_7757,N_7675,N_7698);
or U7758 (N_7758,N_7698,N_7664);
or U7759 (N_7759,N_7605,N_7641);
or U7760 (N_7760,N_7615,N_7641);
or U7761 (N_7761,N_7656,N_7670);
nor U7762 (N_7762,N_7614,N_7601);
or U7763 (N_7763,N_7699,N_7694);
nor U7764 (N_7764,N_7605,N_7603);
or U7765 (N_7765,N_7699,N_7693);
and U7766 (N_7766,N_7699,N_7603);
nor U7767 (N_7767,N_7619,N_7657);
or U7768 (N_7768,N_7667,N_7660);
nor U7769 (N_7769,N_7606,N_7655);
nand U7770 (N_7770,N_7673,N_7632);
and U7771 (N_7771,N_7625,N_7652);
nor U7772 (N_7772,N_7693,N_7692);
and U7773 (N_7773,N_7686,N_7602);
or U7774 (N_7774,N_7673,N_7676);
and U7775 (N_7775,N_7646,N_7664);
or U7776 (N_7776,N_7669,N_7687);
and U7777 (N_7777,N_7631,N_7664);
nand U7778 (N_7778,N_7601,N_7641);
nor U7779 (N_7779,N_7653,N_7663);
nand U7780 (N_7780,N_7670,N_7642);
and U7781 (N_7781,N_7645,N_7606);
and U7782 (N_7782,N_7601,N_7624);
nor U7783 (N_7783,N_7674,N_7610);
nor U7784 (N_7784,N_7698,N_7687);
nor U7785 (N_7785,N_7628,N_7690);
or U7786 (N_7786,N_7673,N_7695);
nor U7787 (N_7787,N_7634,N_7631);
or U7788 (N_7788,N_7657,N_7617);
or U7789 (N_7789,N_7649,N_7609);
nand U7790 (N_7790,N_7625,N_7646);
nor U7791 (N_7791,N_7642,N_7690);
or U7792 (N_7792,N_7642,N_7672);
nor U7793 (N_7793,N_7643,N_7695);
and U7794 (N_7794,N_7672,N_7626);
nor U7795 (N_7795,N_7698,N_7620);
nand U7796 (N_7796,N_7692,N_7670);
or U7797 (N_7797,N_7658,N_7678);
nor U7798 (N_7798,N_7644,N_7607);
or U7799 (N_7799,N_7691,N_7671);
nor U7800 (N_7800,N_7796,N_7748);
nor U7801 (N_7801,N_7769,N_7758);
xor U7802 (N_7802,N_7750,N_7798);
xnor U7803 (N_7803,N_7751,N_7741);
nor U7804 (N_7804,N_7727,N_7712);
nand U7805 (N_7805,N_7760,N_7706);
xor U7806 (N_7806,N_7725,N_7749);
nor U7807 (N_7807,N_7742,N_7777);
and U7808 (N_7808,N_7782,N_7700);
nor U7809 (N_7809,N_7763,N_7746);
nand U7810 (N_7810,N_7759,N_7754);
nand U7811 (N_7811,N_7778,N_7784);
nor U7812 (N_7812,N_7715,N_7774);
nor U7813 (N_7813,N_7775,N_7762);
or U7814 (N_7814,N_7795,N_7710);
or U7815 (N_7815,N_7770,N_7717);
or U7816 (N_7816,N_7730,N_7729);
and U7817 (N_7817,N_7757,N_7786);
and U7818 (N_7818,N_7735,N_7740);
or U7819 (N_7819,N_7747,N_7716);
and U7820 (N_7820,N_7714,N_7731);
nand U7821 (N_7821,N_7745,N_7726);
and U7822 (N_7822,N_7783,N_7734);
nor U7823 (N_7823,N_7765,N_7788);
nand U7824 (N_7824,N_7709,N_7772);
and U7825 (N_7825,N_7722,N_7752);
nor U7826 (N_7826,N_7711,N_7732);
and U7827 (N_7827,N_7720,N_7728);
nor U7828 (N_7828,N_7793,N_7785);
nor U7829 (N_7829,N_7733,N_7773);
nor U7830 (N_7830,N_7781,N_7713);
nand U7831 (N_7831,N_7780,N_7724);
nor U7832 (N_7832,N_7767,N_7753);
or U7833 (N_7833,N_7776,N_7768);
and U7834 (N_7834,N_7703,N_7721);
nor U7835 (N_7835,N_7761,N_7764);
and U7836 (N_7836,N_7736,N_7704);
or U7837 (N_7837,N_7779,N_7799);
or U7838 (N_7838,N_7789,N_7797);
or U7839 (N_7839,N_7771,N_7723);
or U7840 (N_7840,N_7719,N_7705);
nand U7841 (N_7841,N_7791,N_7743);
nand U7842 (N_7842,N_7707,N_7737);
or U7843 (N_7843,N_7792,N_7756);
nor U7844 (N_7844,N_7790,N_7794);
or U7845 (N_7845,N_7738,N_7787);
and U7846 (N_7846,N_7701,N_7708);
nand U7847 (N_7847,N_7744,N_7766);
nor U7848 (N_7848,N_7702,N_7755);
nor U7849 (N_7849,N_7739,N_7718);
or U7850 (N_7850,N_7791,N_7748);
and U7851 (N_7851,N_7788,N_7744);
or U7852 (N_7852,N_7702,N_7781);
xor U7853 (N_7853,N_7736,N_7718);
or U7854 (N_7854,N_7744,N_7785);
nor U7855 (N_7855,N_7707,N_7726);
or U7856 (N_7856,N_7714,N_7728);
nand U7857 (N_7857,N_7739,N_7754);
and U7858 (N_7858,N_7764,N_7720);
and U7859 (N_7859,N_7778,N_7779);
nor U7860 (N_7860,N_7733,N_7711);
or U7861 (N_7861,N_7725,N_7794);
nand U7862 (N_7862,N_7708,N_7760);
or U7863 (N_7863,N_7739,N_7740);
and U7864 (N_7864,N_7733,N_7762);
and U7865 (N_7865,N_7758,N_7790);
or U7866 (N_7866,N_7774,N_7700);
nor U7867 (N_7867,N_7760,N_7721);
or U7868 (N_7868,N_7764,N_7757);
nand U7869 (N_7869,N_7774,N_7725);
nand U7870 (N_7870,N_7746,N_7700);
and U7871 (N_7871,N_7751,N_7754);
nor U7872 (N_7872,N_7799,N_7730);
nand U7873 (N_7873,N_7731,N_7761);
or U7874 (N_7874,N_7722,N_7771);
and U7875 (N_7875,N_7787,N_7797);
and U7876 (N_7876,N_7789,N_7760);
nand U7877 (N_7877,N_7793,N_7740);
nand U7878 (N_7878,N_7716,N_7709);
nand U7879 (N_7879,N_7722,N_7739);
or U7880 (N_7880,N_7727,N_7762);
nor U7881 (N_7881,N_7729,N_7741);
nand U7882 (N_7882,N_7739,N_7702);
nor U7883 (N_7883,N_7780,N_7717);
and U7884 (N_7884,N_7710,N_7702);
and U7885 (N_7885,N_7759,N_7788);
nor U7886 (N_7886,N_7748,N_7797);
xnor U7887 (N_7887,N_7712,N_7761);
nor U7888 (N_7888,N_7703,N_7765);
or U7889 (N_7889,N_7745,N_7773);
nand U7890 (N_7890,N_7753,N_7780);
or U7891 (N_7891,N_7736,N_7752);
or U7892 (N_7892,N_7780,N_7798);
nand U7893 (N_7893,N_7766,N_7759);
or U7894 (N_7894,N_7723,N_7735);
and U7895 (N_7895,N_7789,N_7715);
and U7896 (N_7896,N_7750,N_7776);
or U7897 (N_7897,N_7773,N_7775);
nand U7898 (N_7898,N_7777,N_7797);
nor U7899 (N_7899,N_7777,N_7705);
nand U7900 (N_7900,N_7800,N_7852);
nand U7901 (N_7901,N_7876,N_7875);
nor U7902 (N_7902,N_7807,N_7815);
and U7903 (N_7903,N_7871,N_7805);
or U7904 (N_7904,N_7828,N_7836);
nand U7905 (N_7905,N_7850,N_7853);
or U7906 (N_7906,N_7808,N_7880);
or U7907 (N_7907,N_7830,N_7892);
nor U7908 (N_7908,N_7893,N_7867);
and U7909 (N_7909,N_7868,N_7841);
nor U7910 (N_7910,N_7861,N_7846);
nand U7911 (N_7911,N_7898,N_7821);
and U7912 (N_7912,N_7844,N_7822);
nor U7913 (N_7913,N_7810,N_7825);
or U7914 (N_7914,N_7865,N_7854);
nand U7915 (N_7915,N_7813,N_7820);
and U7916 (N_7916,N_7848,N_7862);
nand U7917 (N_7917,N_7863,N_7802);
nor U7918 (N_7918,N_7882,N_7885);
nor U7919 (N_7919,N_7877,N_7809);
nand U7920 (N_7920,N_7895,N_7842);
nand U7921 (N_7921,N_7827,N_7896);
and U7922 (N_7922,N_7849,N_7832);
and U7923 (N_7923,N_7824,N_7811);
and U7924 (N_7924,N_7856,N_7845);
and U7925 (N_7925,N_7831,N_7866);
nor U7926 (N_7926,N_7881,N_7818);
nand U7927 (N_7927,N_7886,N_7860);
nand U7928 (N_7928,N_7847,N_7838);
or U7929 (N_7929,N_7884,N_7874);
and U7930 (N_7930,N_7872,N_7823);
nor U7931 (N_7931,N_7814,N_7869);
nand U7932 (N_7932,N_7855,N_7834);
and U7933 (N_7933,N_7888,N_7839);
nand U7934 (N_7934,N_7803,N_7859);
nand U7935 (N_7935,N_7816,N_7840);
nand U7936 (N_7936,N_7806,N_7817);
nor U7937 (N_7937,N_7878,N_7887);
or U7938 (N_7938,N_7890,N_7857);
nand U7939 (N_7939,N_7835,N_7891);
or U7940 (N_7940,N_7829,N_7879);
and U7941 (N_7941,N_7837,N_7889);
nor U7942 (N_7942,N_7851,N_7812);
or U7943 (N_7943,N_7899,N_7864);
and U7944 (N_7944,N_7858,N_7801);
nor U7945 (N_7945,N_7833,N_7897);
nor U7946 (N_7946,N_7873,N_7883);
nand U7947 (N_7947,N_7843,N_7826);
or U7948 (N_7948,N_7804,N_7819);
nand U7949 (N_7949,N_7870,N_7894);
nand U7950 (N_7950,N_7815,N_7811);
nand U7951 (N_7951,N_7852,N_7813);
and U7952 (N_7952,N_7865,N_7878);
and U7953 (N_7953,N_7886,N_7840);
and U7954 (N_7954,N_7872,N_7857);
or U7955 (N_7955,N_7840,N_7898);
nor U7956 (N_7956,N_7898,N_7839);
nor U7957 (N_7957,N_7835,N_7839);
or U7958 (N_7958,N_7829,N_7881);
and U7959 (N_7959,N_7807,N_7823);
and U7960 (N_7960,N_7861,N_7822);
or U7961 (N_7961,N_7869,N_7807);
and U7962 (N_7962,N_7869,N_7810);
or U7963 (N_7963,N_7887,N_7880);
or U7964 (N_7964,N_7805,N_7821);
or U7965 (N_7965,N_7810,N_7837);
nor U7966 (N_7966,N_7875,N_7865);
nand U7967 (N_7967,N_7869,N_7892);
nor U7968 (N_7968,N_7855,N_7874);
nor U7969 (N_7969,N_7855,N_7812);
and U7970 (N_7970,N_7875,N_7874);
nor U7971 (N_7971,N_7891,N_7805);
nand U7972 (N_7972,N_7852,N_7858);
or U7973 (N_7973,N_7802,N_7897);
nor U7974 (N_7974,N_7882,N_7867);
nand U7975 (N_7975,N_7851,N_7870);
or U7976 (N_7976,N_7865,N_7800);
and U7977 (N_7977,N_7829,N_7823);
nand U7978 (N_7978,N_7812,N_7815);
nor U7979 (N_7979,N_7813,N_7855);
or U7980 (N_7980,N_7850,N_7805);
nor U7981 (N_7981,N_7842,N_7855);
or U7982 (N_7982,N_7842,N_7827);
nor U7983 (N_7983,N_7892,N_7800);
nand U7984 (N_7984,N_7822,N_7887);
or U7985 (N_7985,N_7898,N_7860);
and U7986 (N_7986,N_7819,N_7842);
or U7987 (N_7987,N_7870,N_7863);
or U7988 (N_7988,N_7824,N_7807);
and U7989 (N_7989,N_7825,N_7860);
or U7990 (N_7990,N_7831,N_7898);
nor U7991 (N_7991,N_7859,N_7888);
nand U7992 (N_7992,N_7862,N_7860);
and U7993 (N_7993,N_7871,N_7833);
and U7994 (N_7994,N_7827,N_7825);
and U7995 (N_7995,N_7876,N_7817);
nand U7996 (N_7996,N_7803,N_7845);
or U7997 (N_7997,N_7864,N_7851);
or U7998 (N_7998,N_7877,N_7803);
or U7999 (N_7999,N_7842,N_7836);
and U8000 (N_8000,N_7904,N_7933);
or U8001 (N_8001,N_7972,N_7968);
and U8002 (N_8002,N_7994,N_7932);
and U8003 (N_8003,N_7910,N_7909);
and U8004 (N_8004,N_7934,N_7961);
or U8005 (N_8005,N_7905,N_7917);
nand U8006 (N_8006,N_7952,N_7946);
nor U8007 (N_8007,N_7983,N_7986);
nor U8008 (N_8008,N_7997,N_7935);
nand U8009 (N_8009,N_7954,N_7988);
and U8010 (N_8010,N_7945,N_7930);
or U8011 (N_8011,N_7918,N_7973);
nor U8012 (N_8012,N_7940,N_7995);
or U8013 (N_8013,N_7967,N_7998);
or U8014 (N_8014,N_7941,N_7914);
nor U8015 (N_8015,N_7912,N_7959);
nor U8016 (N_8016,N_7903,N_7916);
xnor U8017 (N_8017,N_7943,N_7979);
or U8018 (N_8018,N_7956,N_7987);
and U8019 (N_8019,N_7915,N_7901);
xor U8020 (N_8020,N_7942,N_7978);
nand U8021 (N_8021,N_7911,N_7964);
nand U8022 (N_8022,N_7924,N_7960);
xor U8023 (N_8023,N_7970,N_7923);
and U8024 (N_8024,N_7939,N_7929);
and U8025 (N_8025,N_7928,N_7955);
or U8026 (N_8026,N_7953,N_7982);
nand U8027 (N_8027,N_7969,N_7984);
nor U8028 (N_8028,N_7949,N_7963);
nand U8029 (N_8029,N_7927,N_7947);
or U8030 (N_8030,N_7966,N_7907);
and U8031 (N_8031,N_7957,N_7980);
nor U8032 (N_8032,N_7999,N_7958);
and U8033 (N_8033,N_7992,N_7906);
or U8034 (N_8034,N_7937,N_7926);
and U8035 (N_8035,N_7991,N_7908);
or U8036 (N_8036,N_7981,N_7962);
nand U8037 (N_8037,N_7902,N_7944);
nand U8038 (N_8038,N_7922,N_7993);
or U8039 (N_8039,N_7925,N_7974);
nand U8040 (N_8040,N_7913,N_7919);
nor U8041 (N_8041,N_7965,N_7948);
or U8042 (N_8042,N_7975,N_7900);
or U8043 (N_8043,N_7950,N_7971);
nor U8044 (N_8044,N_7990,N_7938);
or U8045 (N_8045,N_7921,N_7985);
xor U8046 (N_8046,N_7976,N_7989);
and U8047 (N_8047,N_7996,N_7931);
nand U8048 (N_8048,N_7936,N_7920);
nor U8049 (N_8049,N_7951,N_7977);
nand U8050 (N_8050,N_7941,N_7943);
nor U8051 (N_8051,N_7976,N_7958);
nand U8052 (N_8052,N_7924,N_7941);
and U8053 (N_8053,N_7975,N_7953);
nor U8054 (N_8054,N_7962,N_7916);
or U8055 (N_8055,N_7983,N_7971);
and U8056 (N_8056,N_7915,N_7923);
or U8057 (N_8057,N_7991,N_7903);
nor U8058 (N_8058,N_7911,N_7980);
nand U8059 (N_8059,N_7919,N_7912);
and U8060 (N_8060,N_7949,N_7966);
nand U8061 (N_8061,N_7939,N_7961);
and U8062 (N_8062,N_7991,N_7935);
and U8063 (N_8063,N_7941,N_7908);
and U8064 (N_8064,N_7961,N_7950);
nand U8065 (N_8065,N_7940,N_7998);
nand U8066 (N_8066,N_7959,N_7983);
and U8067 (N_8067,N_7962,N_7979);
nand U8068 (N_8068,N_7976,N_7953);
and U8069 (N_8069,N_7988,N_7947);
nor U8070 (N_8070,N_7953,N_7902);
nor U8071 (N_8071,N_7928,N_7984);
xnor U8072 (N_8072,N_7980,N_7963);
nand U8073 (N_8073,N_7957,N_7944);
or U8074 (N_8074,N_7976,N_7912);
nor U8075 (N_8075,N_7908,N_7917);
nor U8076 (N_8076,N_7920,N_7962);
or U8077 (N_8077,N_7991,N_7956);
and U8078 (N_8078,N_7973,N_7989);
xnor U8079 (N_8079,N_7920,N_7994);
nor U8080 (N_8080,N_7913,N_7994);
nand U8081 (N_8081,N_7924,N_7933);
nor U8082 (N_8082,N_7927,N_7990);
nor U8083 (N_8083,N_7945,N_7927);
and U8084 (N_8084,N_7946,N_7930);
or U8085 (N_8085,N_7950,N_7926);
and U8086 (N_8086,N_7977,N_7907);
nor U8087 (N_8087,N_7996,N_7956);
or U8088 (N_8088,N_7958,N_7989);
and U8089 (N_8089,N_7950,N_7912);
or U8090 (N_8090,N_7985,N_7930);
nand U8091 (N_8091,N_7970,N_7953);
nor U8092 (N_8092,N_7978,N_7992);
or U8093 (N_8093,N_7988,N_7901);
nor U8094 (N_8094,N_7955,N_7908);
nand U8095 (N_8095,N_7901,N_7922);
and U8096 (N_8096,N_7907,N_7923);
nand U8097 (N_8097,N_7926,N_7974);
nand U8098 (N_8098,N_7991,N_7923);
or U8099 (N_8099,N_7980,N_7993);
nand U8100 (N_8100,N_8068,N_8088);
nand U8101 (N_8101,N_8056,N_8054);
or U8102 (N_8102,N_8052,N_8080);
nor U8103 (N_8103,N_8086,N_8034);
nor U8104 (N_8104,N_8030,N_8074);
nor U8105 (N_8105,N_8071,N_8072);
nor U8106 (N_8106,N_8003,N_8009);
or U8107 (N_8107,N_8013,N_8002);
nand U8108 (N_8108,N_8055,N_8098);
or U8109 (N_8109,N_8087,N_8060);
and U8110 (N_8110,N_8090,N_8062);
or U8111 (N_8111,N_8059,N_8029);
nand U8112 (N_8112,N_8026,N_8097);
nand U8113 (N_8113,N_8015,N_8005);
nand U8114 (N_8114,N_8017,N_8046);
or U8115 (N_8115,N_8092,N_8010);
and U8116 (N_8116,N_8039,N_8020);
or U8117 (N_8117,N_8000,N_8045);
nand U8118 (N_8118,N_8011,N_8022);
nor U8119 (N_8119,N_8091,N_8069);
nand U8120 (N_8120,N_8031,N_8082);
nor U8121 (N_8121,N_8024,N_8028);
and U8122 (N_8122,N_8021,N_8075);
and U8123 (N_8123,N_8096,N_8037);
or U8124 (N_8124,N_8050,N_8099);
nand U8125 (N_8125,N_8077,N_8057);
and U8126 (N_8126,N_8008,N_8004);
and U8127 (N_8127,N_8065,N_8063);
nand U8128 (N_8128,N_8093,N_8027);
or U8129 (N_8129,N_8083,N_8044);
or U8130 (N_8130,N_8070,N_8051);
nor U8131 (N_8131,N_8095,N_8035);
or U8132 (N_8132,N_8040,N_8081);
and U8133 (N_8133,N_8043,N_8025);
nand U8134 (N_8134,N_8007,N_8067);
nand U8135 (N_8135,N_8064,N_8061);
and U8136 (N_8136,N_8012,N_8079);
or U8137 (N_8137,N_8073,N_8023);
nand U8138 (N_8138,N_8006,N_8048);
or U8139 (N_8139,N_8089,N_8018);
and U8140 (N_8140,N_8049,N_8085);
and U8141 (N_8141,N_8041,N_8084);
and U8142 (N_8142,N_8014,N_8032);
and U8143 (N_8143,N_8019,N_8001);
nand U8144 (N_8144,N_8033,N_8094);
nand U8145 (N_8145,N_8076,N_8078);
or U8146 (N_8146,N_8042,N_8016);
nand U8147 (N_8147,N_8066,N_8038);
xor U8148 (N_8148,N_8036,N_8047);
nand U8149 (N_8149,N_8058,N_8053);
nor U8150 (N_8150,N_8087,N_8005);
nand U8151 (N_8151,N_8046,N_8098);
or U8152 (N_8152,N_8086,N_8051);
nand U8153 (N_8153,N_8094,N_8077);
or U8154 (N_8154,N_8061,N_8078);
nor U8155 (N_8155,N_8080,N_8032);
and U8156 (N_8156,N_8084,N_8063);
or U8157 (N_8157,N_8081,N_8085);
nand U8158 (N_8158,N_8002,N_8087);
nand U8159 (N_8159,N_8085,N_8074);
or U8160 (N_8160,N_8015,N_8006);
or U8161 (N_8161,N_8072,N_8008);
or U8162 (N_8162,N_8091,N_8042);
xnor U8163 (N_8163,N_8037,N_8009);
nand U8164 (N_8164,N_8001,N_8034);
or U8165 (N_8165,N_8015,N_8043);
and U8166 (N_8166,N_8077,N_8086);
nor U8167 (N_8167,N_8007,N_8045);
nand U8168 (N_8168,N_8000,N_8085);
nor U8169 (N_8169,N_8065,N_8013);
nand U8170 (N_8170,N_8083,N_8029);
nand U8171 (N_8171,N_8046,N_8023);
or U8172 (N_8172,N_8052,N_8013);
or U8173 (N_8173,N_8032,N_8058);
or U8174 (N_8174,N_8055,N_8009);
and U8175 (N_8175,N_8055,N_8035);
nand U8176 (N_8176,N_8043,N_8094);
nand U8177 (N_8177,N_8063,N_8086);
and U8178 (N_8178,N_8046,N_8037);
nand U8179 (N_8179,N_8080,N_8031);
and U8180 (N_8180,N_8055,N_8058);
nand U8181 (N_8181,N_8067,N_8071);
or U8182 (N_8182,N_8020,N_8071);
nand U8183 (N_8183,N_8079,N_8099);
or U8184 (N_8184,N_8049,N_8034);
nand U8185 (N_8185,N_8034,N_8037);
nand U8186 (N_8186,N_8046,N_8082);
or U8187 (N_8187,N_8079,N_8091);
and U8188 (N_8188,N_8058,N_8090);
and U8189 (N_8189,N_8078,N_8081);
and U8190 (N_8190,N_8041,N_8032);
or U8191 (N_8191,N_8030,N_8098);
and U8192 (N_8192,N_8005,N_8080);
and U8193 (N_8193,N_8056,N_8089);
nor U8194 (N_8194,N_8070,N_8039);
or U8195 (N_8195,N_8084,N_8011);
nor U8196 (N_8196,N_8004,N_8035);
nand U8197 (N_8197,N_8054,N_8052);
nor U8198 (N_8198,N_8005,N_8023);
and U8199 (N_8199,N_8075,N_8008);
nor U8200 (N_8200,N_8136,N_8153);
or U8201 (N_8201,N_8154,N_8165);
nand U8202 (N_8202,N_8191,N_8109);
and U8203 (N_8203,N_8117,N_8103);
and U8204 (N_8204,N_8143,N_8172);
nand U8205 (N_8205,N_8183,N_8173);
xnor U8206 (N_8206,N_8113,N_8171);
or U8207 (N_8207,N_8149,N_8186);
nor U8208 (N_8208,N_8124,N_8176);
nor U8209 (N_8209,N_8137,N_8174);
and U8210 (N_8210,N_8129,N_8192);
nor U8211 (N_8211,N_8170,N_8115);
nand U8212 (N_8212,N_8161,N_8121);
or U8213 (N_8213,N_8105,N_8159);
nand U8214 (N_8214,N_8158,N_8152);
xor U8215 (N_8215,N_8193,N_8151);
and U8216 (N_8216,N_8156,N_8155);
nor U8217 (N_8217,N_8185,N_8106);
nand U8218 (N_8218,N_8187,N_8189);
and U8219 (N_8219,N_8147,N_8125);
nor U8220 (N_8220,N_8112,N_8101);
and U8221 (N_8221,N_8180,N_8169);
nand U8222 (N_8222,N_8182,N_8190);
nand U8223 (N_8223,N_8140,N_8122);
or U8224 (N_8224,N_8199,N_8118);
or U8225 (N_8225,N_8168,N_8135);
nand U8226 (N_8226,N_8107,N_8134);
or U8227 (N_8227,N_8157,N_8138);
nor U8228 (N_8228,N_8131,N_8177);
nor U8229 (N_8229,N_8181,N_8163);
and U8230 (N_8230,N_8188,N_8148);
xnor U8231 (N_8231,N_8197,N_8166);
xor U8232 (N_8232,N_8195,N_8104);
and U8233 (N_8233,N_8108,N_8123);
nor U8234 (N_8234,N_8175,N_8102);
or U8235 (N_8235,N_8164,N_8179);
nor U8236 (N_8236,N_8130,N_8167);
nand U8237 (N_8237,N_8142,N_8100);
nand U8238 (N_8238,N_8145,N_8146);
xor U8239 (N_8239,N_8132,N_8110);
and U8240 (N_8240,N_8120,N_8141);
and U8241 (N_8241,N_8178,N_8198);
and U8242 (N_8242,N_8133,N_8196);
and U8243 (N_8243,N_8116,N_8162);
nand U8244 (N_8244,N_8126,N_8144);
nor U8245 (N_8245,N_8127,N_8150);
nor U8246 (N_8246,N_8128,N_8111);
or U8247 (N_8247,N_8139,N_8114);
nand U8248 (N_8248,N_8160,N_8119);
and U8249 (N_8249,N_8184,N_8194);
and U8250 (N_8250,N_8104,N_8162);
and U8251 (N_8251,N_8142,N_8143);
nor U8252 (N_8252,N_8176,N_8199);
xor U8253 (N_8253,N_8166,N_8110);
nand U8254 (N_8254,N_8199,N_8162);
and U8255 (N_8255,N_8171,N_8105);
nand U8256 (N_8256,N_8178,N_8173);
xnor U8257 (N_8257,N_8187,N_8169);
nor U8258 (N_8258,N_8139,N_8136);
nor U8259 (N_8259,N_8134,N_8165);
nand U8260 (N_8260,N_8176,N_8186);
and U8261 (N_8261,N_8130,N_8136);
nand U8262 (N_8262,N_8188,N_8145);
and U8263 (N_8263,N_8140,N_8155);
and U8264 (N_8264,N_8153,N_8135);
nand U8265 (N_8265,N_8128,N_8163);
nor U8266 (N_8266,N_8123,N_8147);
and U8267 (N_8267,N_8135,N_8126);
and U8268 (N_8268,N_8195,N_8127);
nor U8269 (N_8269,N_8196,N_8162);
and U8270 (N_8270,N_8129,N_8197);
or U8271 (N_8271,N_8146,N_8105);
and U8272 (N_8272,N_8182,N_8136);
nand U8273 (N_8273,N_8177,N_8168);
and U8274 (N_8274,N_8197,N_8160);
nor U8275 (N_8275,N_8189,N_8175);
nor U8276 (N_8276,N_8184,N_8104);
nand U8277 (N_8277,N_8180,N_8114);
nor U8278 (N_8278,N_8172,N_8138);
xor U8279 (N_8279,N_8187,N_8153);
nor U8280 (N_8280,N_8102,N_8122);
or U8281 (N_8281,N_8190,N_8139);
nand U8282 (N_8282,N_8122,N_8157);
and U8283 (N_8283,N_8185,N_8160);
and U8284 (N_8284,N_8101,N_8158);
nand U8285 (N_8285,N_8187,N_8168);
nand U8286 (N_8286,N_8105,N_8184);
nand U8287 (N_8287,N_8153,N_8163);
and U8288 (N_8288,N_8101,N_8173);
nor U8289 (N_8289,N_8146,N_8155);
nand U8290 (N_8290,N_8176,N_8175);
and U8291 (N_8291,N_8162,N_8108);
nand U8292 (N_8292,N_8173,N_8152);
nor U8293 (N_8293,N_8146,N_8154);
nand U8294 (N_8294,N_8141,N_8176);
nor U8295 (N_8295,N_8123,N_8180);
nand U8296 (N_8296,N_8189,N_8172);
or U8297 (N_8297,N_8149,N_8128);
nand U8298 (N_8298,N_8120,N_8156);
or U8299 (N_8299,N_8127,N_8138);
or U8300 (N_8300,N_8299,N_8265);
and U8301 (N_8301,N_8226,N_8241);
and U8302 (N_8302,N_8207,N_8200);
and U8303 (N_8303,N_8252,N_8220);
or U8304 (N_8304,N_8229,N_8204);
or U8305 (N_8305,N_8257,N_8264);
or U8306 (N_8306,N_8276,N_8287);
nor U8307 (N_8307,N_8279,N_8277);
or U8308 (N_8308,N_8254,N_8281);
and U8309 (N_8309,N_8209,N_8272);
nor U8310 (N_8310,N_8240,N_8271);
nor U8311 (N_8311,N_8213,N_8235);
nor U8312 (N_8312,N_8206,N_8224);
nor U8313 (N_8313,N_8263,N_8208);
nor U8314 (N_8314,N_8251,N_8225);
nor U8315 (N_8315,N_8256,N_8295);
nand U8316 (N_8316,N_8219,N_8223);
and U8317 (N_8317,N_8232,N_8227);
and U8318 (N_8318,N_8212,N_8261);
and U8319 (N_8319,N_8230,N_8296);
nor U8320 (N_8320,N_8245,N_8236);
or U8321 (N_8321,N_8250,N_8273);
nand U8322 (N_8322,N_8228,N_8266);
or U8323 (N_8323,N_8290,N_8249);
nor U8324 (N_8324,N_8258,N_8255);
nor U8325 (N_8325,N_8205,N_8292);
nor U8326 (N_8326,N_8274,N_8280);
and U8327 (N_8327,N_8222,N_8260);
nand U8328 (N_8328,N_8286,N_8262);
nand U8329 (N_8329,N_8270,N_8210);
nand U8330 (N_8330,N_8243,N_8246);
or U8331 (N_8331,N_8248,N_8239);
and U8332 (N_8332,N_8201,N_8217);
and U8333 (N_8333,N_8291,N_8214);
nor U8334 (N_8334,N_8294,N_8268);
or U8335 (N_8335,N_8233,N_8288);
nand U8336 (N_8336,N_8298,N_8203);
and U8337 (N_8337,N_8259,N_8202);
or U8338 (N_8338,N_8237,N_8238);
nand U8339 (N_8339,N_8253,N_8285);
or U8340 (N_8340,N_8215,N_8231);
nor U8341 (N_8341,N_8242,N_8216);
or U8342 (N_8342,N_8289,N_8234);
nor U8343 (N_8343,N_8269,N_8293);
nand U8344 (N_8344,N_8283,N_8221);
or U8345 (N_8345,N_8297,N_8278);
nand U8346 (N_8346,N_8284,N_8275);
and U8347 (N_8347,N_8282,N_8247);
nand U8348 (N_8348,N_8244,N_8267);
nand U8349 (N_8349,N_8211,N_8218);
nand U8350 (N_8350,N_8264,N_8282);
or U8351 (N_8351,N_8280,N_8269);
nor U8352 (N_8352,N_8235,N_8208);
and U8353 (N_8353,N_8237,N_8243);
and U8354 (N_8354,N_8279,N_8214);
and U8355 (N_8355,N_8271,N_8224);
xor U8356 (N_8356,N_8295,N_8272);
xor U8357 (N_8357,N_8293,N_8287);
xnor U8358 (N_8358,N_8264,N_8204);
and U8359 (N_8359,N_8244,N_8286);
and U8360 (N_8360,N_8221,N_8265);
nor U8361 (N_8361,N_8224,N_8232);
nand U8362 (N_8362,N_8268,N_8288);
nor U8363 (N_8363,N_8278,N_8291);
and U8364 (N_8364,N_8205,N_8290);
or U8365 (N_8365,N_8299,N_8201);
nor U8366 (N_8366,N_8274,N_8233);
nand U8367 (N_8367,N_8237,N_8293);
or U8368 (N_8368,N_8215,N_8243);
or U8369 (N_8369,N_8203,N_8235);
nand U8370 (N_8370,N_8219,N_8256);
or U8371 (N_8371,N_8236,N_8204);
nand U8372 (N_8372,N_8225,N_8236);
nor U8373 (N_8373,N_8273,N_8243);
nor U8374 (N_8374,N_8204,N_8245);
nand U8375 (N_8375,N_8210,N_8246);
or U8376 (N_8376,N_8246,N_8211);
nor U8377 (N_8377,N_8205,N_8202);
nand U8378 (N_8378,N_8265,N_8204);
or U8379 (N_8379,N_8274,N_8221);
nand U8380 (N_8380,N_8221,N_8264);
nor U8381 (N_8381,N_8252,N_8236);
nor U8382 (N_8382,N_8280,N_8228);
nor U8383 (N_8383,N_8264,N_8244);
or U8384 (N_8384,N_8287,N_8252);
nand U8385 (N_8385,N_8218,N_8207);
nor U8386 (N_8386,N_8263,N_8255);
and U8387 (N_8387,N_8278,N_8262);
nand U8388 (N_8388,N_8264,N_8201);
and U8389 (N_8389,N_8243,N_8297);
and U8390 (N_8390,N_8276,N_8255);
nand U8391 (N_8391,N_8250,N_8290);
and U8392 (N_8392,N_8210,N_8236);
nor U8393 (N_8393,N_8200,N_8265);
or U8394 (N_8394,N_8246,N_8242);
and U8395 (N_8395,N_8274,N_8282);
nand U8396 (N_8396,N_8288,N_8264);
and U8397 (N_8397,N_8266,N_8227);
or U8398 (N_8398,N_8288,N_8241);
or U8399 (N_8399,N_8237,N_8201);
or U8400 (N_8400,N_8368,N_8304);
and U8401 (N_8401,N_8388,N_8385);
nand U8402 (N_8402,N_8313,N_8371);
and U8403 (N_8403,N_8395,N_8341);
or U8404 (N_8404,N_8366,N_8315);
nand U8405 (N_8405,N_8327,N_8397);
or U8406 (N_8406,N_8342,N_8344);
or U8407 (N_8407,N_8346,N_8323);
and U8408 (N_8408,N_8307,N_8390);
or U8409 (N_8409,N_8314,N_8391);
and U8410 (N_8410,N_8343,N_8347);
or U8411 (N_8411,N_8357,N_8382);
nand U8412 (N_8412,N_8328,N_8372);
and U8413 (N_8413,N_8399,N_8378);
nand U8414 (N_8414,N_8369,N_8386);
and U8415 (N_8415,N_8305,N_8380);
or U8416 (N_8416,N_8396,N_8302);
nor U8417 (N_8417,N_8303,N_8345);
nor U8418 (N_8418,N_8330,N_8300);
nor U8419 (N_8419,N_8350,N_8316);
nor U8420 (N_8420,N_8312,N_8373);
or U8421 (N_8421,N_8338,N_8348);
nor U8422 (N_8422,N_8301,N_8360);
and U8423 (N_8423,N_8326,N_8365);
nor U8424 (N_8424,N_8393,N_8394);
and U8425 (N_8425,N_8392,N_8337);
or U8426 (N_8426,N_8318,N_8362);
or U8427 (N_8427,N_8356,N_8379);
xor U8428 (N_8428,N_8376,N_8364);
and U8429 (N_8429,N_8325,N_8354);
nand U8430 (N_8430,N_8321,N_8398);
or U8431 (N_8431,N_8331,N_8367);
or U8432 (N_8432,N_8377,N_8374);
nand U8433 (N_8433,N_8361,N_8359);
nand U8434 (N_8434,N_8387,N_8322);
or U8435 (N_8435,N_8339,N_8319);
or U8436 (N_8436,N_8329,N_8381);
nand U8437 (N_8437,N_8355,N_8317);
or U8438 (N_8438,N_8383,N_8363);
or U8439 (N_8439,N_8335,N_8333);
nor U8440 (N_8440,N_8334,N_8336);
and U8441 (N_8441,N_8384,N_8352);
or U8442 (N_8442,N_8324,N_8311);
xor U8443 (N_8443,N_8353,N_8320);
and U8444 (N_8444,N_8370,N_8375);
and U8445 (N_8445,N_8340,N_8306);
nor U8446 (N_8446,N_8351,N_8308);
nor U8447 (N_8447,N_8332,N_8310);
nand U8448 (N_8448,N_8349,N_8358);
nor U8449 (N_8449,N_8389,N_8309);
or U8450 (N_8450,N_8339,N_8325);
or U8451 (N_8451,N_8343,N_8388);
or U8452 (N_8452,N_8347,N_8328);
or U8453 (N_8453,N_8307,N_8366);
nor U8454 (N_8454,N_8396,N_8397);
or U8455 (N_8455,N_8331,N_8311);
or U8456 (N_8456,N_8322,N_8341);
or U8457 (N_8457,N_8303,N_8353);
nor U8458 (N_8458,N_8333,N_8377);
nor U8459 (N_8459,N_8393,N_8337);
nor U8460 (N_8460,N_8370,N_8338);
nor U8461 (N_8461,N_8343,N_8305);
and U8462 (N_8462,N_8336,N_8386);
nor U8463 (N_8463,N_8395,N_8372);
or U8464 (N_8464,N_8326,N_8303);
or U8465 (N_8465,N_8341,N_8360);
nor U8466 (N_8466,N_8330,N_8310);
and U8467 (N_8467,N_8394,N_8314);
and U8468 (N_8468,N_8378,N_8349);
nand U8469 (N_8469,N_8383,N_8376);
or U8470 (N_8470,N_8372,N_8300);
nor U8471 (N_8471,N_8389,N_8331);
or U8472 (N_8472,N_8307,N_8305);
or U8473 (N_8473,N_8373,N_8392);
nor U8474 (N_8474,N_8397,N_8391);
or U8475 (N_8475,N_8347,N_8383);
or U8476 (N_8476,N_8394,N_8337);
and U8477 (N_8477,N_8345,N_8396);
or U8478 (N_8478,N_8348,N_8395);
nand U8479 (N_8479,N_8357,N_8365);
or U8480 (N_8480,N_8341,N_8334);
nor U8481 (N_8481,N_8304,N_8302);
and U8482 (N_8482,N_8347,N_8332);
nor U8483 (N_8483,N_8377,N_8335);
or U8484 (N_8484,N_8325,N_8359);
or U8485 (N_8485,N_8377,N_8353);
and U8486 (N_8486,N_8338,N_8354);
nor U8487 (N_8487,N_8309,N_8384);
xnor U8488 (N_8488,N_8337,N_8331);
and U8489 (N_8489,N_8317,N_8334);
nand U8490 (N_8490,N_8358,N_8388);
or U8491 (N_8491,N_8358,N_8377);
nor U8492 (N_8492,N_8315,N_8376);
or U8493 (N_8493,N_8388,N_8350);
nand U8494 (N_8494,N_8378,N_8334);
and U8495 (N_8495,N_8355,N_8368);
nand U8496 (N_8496,N_8353,N_8384);
nor U8497 (N_8497,N_8300,N_8375);
nand U8498 (N_8498,N_8310,N_8321);
xnor U8499 (N_8499,N_8382,N_8348);
or U8500 (N_8500,N_8416,N_8443);
or U8501 (N_8501,N_8467,N_8439);
nand U8502 (N_8502,N_8453,N_8424);
or U8503 (N_8503,N_8410,N_8454);
xor U8504 (N_8504,N_8427,N_8426);
nor U8505 (N_8505,N_8421,N_8469);
and U8506 (N_8506,N_8489,N_8475);
or U8507 (N_8507,N_8472,N_8493);
or U8508 (N_8508,N_8411,N_8418);
or U8509 (N_8509,N_8490,N_8466);
nand U8510 (N_8510,N_8409,N_8423);
nand U8511 (N_8511,N_8414,N_8407);
and U8512 (N_8512,N_8496,N_8444);
or U8513 (N_8513,N_8406,N_8457);
nand U8514 (N_8514,N_8481,N_8437);
or U8515 (N_8515,N_8495,N_8491);
and U8516 (N_8516,N_8446,N_8420);
or U8517 (N_8517,N_8450,N_8499);
nor U8518 (N_8518,N_8452,N_8468);
nand U8519 (N_8519,N_8474,N_8478);
and U8520 (N_8520,N_8488,N_8436);
nand U8521 (N_8521,N_8403,N_8408);
and U8522 (N_8522,N_8431,N_8432);
nand U8523 (N_8523,N_8405,N_8415);
nand U8524 (N_8524,N_8498,N_8479);
or U8525 (N_8525,N_8476,N_8462);
nand U8526 (N_8526,N_8465,N_8486);
and U8527 (N_8527,N_8463,N_8487);
or U8528 (N_8528,N_8483,N_8460);
and U8529 (N_8529,N_8419,N_8494);
nor U8530 (N_8530,N_8445,N_8417);
xnor U8531 (N_8531,N_8404,N_8485);
or U8532 (N_8532,N_8430,N_8412);
nor U8533 (N_8533,N_8497,N_8400);
or U8534 (N_8534,N_8433,N_8425);
nand U8535 (N_8535,N_8461,N_8458);
or U8536 (N_8536,N_8438,N_8413);
and U8537 (N_8537,N_8471,N_8428);
or U8538 (N_8538,N_8484,N_8464);
and U8539 (N_8539,N_8470,N_8492);
and U8540 (N_8540,N_8473,N_8455);
nand U8541 (N_8541,N_8442,N_8440);
nor U8542 (N_8542,N_8456,N_8422);
and U8543 (N_8543,N_8451,N_8449);
and U8544 (N_8544,N_8447,N_8448);
or U8545 (N_8545,N_8459,N_8435);
or U8546 (N_8546,N_8480,N_8401);
nor U8547 (N_8547,N_8441,N_8477);
nand U8548 (N_8548,N_8429,N_8402);
or U8549 (N_8549,N_8482,N_8434);
xor U8550 (N_8550,N_8415,N_8445);
nand U8551 (N_8551,N_8430,N_8497);
nand U8552 (N_8552,N_8497,N_8423);
nor U8553 (N_8553,N_8424,N_8443);
or U8554 (N_8554,N_8439,N_8441);
nand U8555 (N_8555,N_8407,N_8408);
and U8556 (N_8556,N_8412,N_8440);
or U8557 (N_8557,N_8439,N_8429);
xor U8558 (N_8558,N_8442,N_8451);
and U8559 (N_8559,N_8416,N_8447);
and U8560 (N_8560,N_8475,N_8455);
and U8561 (N_8561,N_8405,N_8401);
and U8562 (N_8562,N_8454,N_8476);
or U8563 (N_8563,N_8410,N_8497);
nor U8564 (N_8564,N_8464,N_8492);
and U8565 (N_8565,N_8474,N_8410);
nand U8566 (N_8566,N_8429,N_8407);
or U8567 (N_8567,N_8454,N_8425);
or U8568 (N_8568,N_8428,N_8456);
or U8569 (N_8569,N_8434,N_8438);
and U8570 (N_8570,N_8406,N_8446);
nor U8571 (N_8571,N_8471,N_8427);
nand U8572 (N_8572,N_8423,N_8474);
nor U8573 (N_8573,N_8433,N_8401);
or U8574 (N_8574,N_8414,N_8475);
and U8575 (N_8575,N_8423,N_8485);
nor U8576 (N_8576,N_8446,N_8407);
nand U8577 (N_8577,N_8430,N_8450);
and U8578 (N_8578,N_8438,N_8486);
nor U8579 (N_8579,N_8481,N_8469);
or U8580 (N_8580,N_8458,N_8483);
nor U8581 (N_8581,N_8410,N_8459);
nand U8582 (N_8582,N_8489,N_8462);
nand U8583 (N_8583,N_8461,N_8491);
nor U8584 (N_8584,N_8451,N_8476);
nand U8585 (N_8585,N_8439,N_8405);
or U8586 (N_8586,N_8436,N_8463);
nor U8587 (N_8587,N_8434,N_8410);
and U8588 (N_8588,N_8403,N_8452);
nor U8589 (N_8589,N_8492,N_8413);
and U8590 (N_8590,N_8432,N_8440);
nand U8591 (N_8591,N_8450,N_8418);
or U8592 (N_8592,N_8429,N_8419);
nor U8593 (N_8593,N_8462,N_8470);
and U8594 (N_8594,N_8487,N_8438);
or U8595 (N_8595,N_8475,N_8439);
nand U8596 (N_8596,N_8444,N_8451);
xnor U8597 (N_8597,N_8441,N_8491);
nor U8598 (N_8598,N_8460,N_8438);
and U8599 (N_8599,N_8415,N_8488);
and U8600 (N_8600,N_8560,N_8590);
nand U8601 (N_8601,N_8593,N_8556);
nor U8602 (N_8602,N_8558,N_8575);
and U8603 (N_8603,N_8540,N_8578);
nor U8604 (N_8604,N_8567,N_8520);
nand U8605 (N_8605,N_8597,N_8529);
nand U8606 (N_8606,N_8534,N_8552);
nor U8607 (N_8607,N_8503,N_8500);
nor U8608 (N_8608,N_8538,N_8588);
nand U8609 (N_8609,N_8587,N_8525);
nor U8610 (N_8610,N_8562,N_8507);
nor U8611 (N_8611,N_8523,N_8584);
and U8612 (N_8612,N_8533,N_8595);
nand U8613 (N_8613,N_8596,N_8573);
nand U8614 (N_8614,N_8536,N_8524);
and U8615 (N_8615,N_8554,N_8566);
nand U8616 (N_8616,N_8547,N_8516);
and U8617 (N_8617,N_8557,N_8545);
nor U8618 (N_8618,N_8504,N_8592);
nor U8619 (N_8619,N_8506,N_8543);
and U8620 (N_8620,N_8565,N_8585);
nand U8621 (N_8621,N_8577,N_8555);
or U8622 (N_8622,N_8549,N_8550);
nor U8623 (N_8623,N_8531,N_8517);
nand U8624 (N_8624,N_8576,N_8564);
or U8625 (N_8625,N_8586,N_8509);
and U8626 (N_8626,N_8508,N_8580);
nor U8627 (N_8627,N_8527,N_8522);
nand U8628 (N_8628,N_8544,N_8502);
and U8629 (N_8629,N_8528,N_8511);
or U8630 (N_8630,N_8513,N_8583);
nand U8631 (N_8631,N_8582,N_8537);
nor U8632 (N_8632,N_8553,N_8568);
nand U8633 (N_8633,N_8542,N_8515);
or U8634 (N_8634,N_8572,N_8591);
or U8635 (N_8635,N_8559,N_8546);
nor U8636 (N_8636,N_8535,N_8518);
nor U8637 (N_8637,N_8521,N_8598);
and U8638 (N_8638,N_8589,N_8530);
nand U8639 (N_8639,N_8594,N_8581);
nand U8640 (N_8640,N_8526,N_8548);
nor U8641 (N_8641,N_8561,N_8512);
nand U8642 (N_8642,N_8563,N_8532);
xnor U8643 (N_8643,N_8599,N_8539);
or U8644 (N_8644,N_8571,N_8569);
nand U8645 (N_8645,N_8501,N_8519);
nand U8646 (N_8646,N_8579,N_8510);
or U8647 (N_8647,N_8570,N_8514);
nor U8648 (N_8648,N_8541,N_8505);
nand U8649 (N_8649,N_8551,N_8574);
or U8650 (N_8650,N_8559,N_8529);
nand U8651 (N_8651,N_8551,N_8599);
xor U8652 (N_8652,N_8555,N_8521);
or U8653 (N_8653,N_8550,N_8553);
and U8654 (N_8654,N_8566,N_8545);
nor U8655 (N_8655,N_8505,N_8500);
nand U8656 (N_8656,N_8594,N_8535);
nor U8657 (N_8657,N_8520,N_8509);
and U8658 (N_8658,N_8544,N_8593);
and U8659 (N_8659,N_8577,N_8550);
or U8660 (N_8660,N_8529,N_8526);
or U8661 (N_8661,N_8571,N_8590);
or U8662 (N_8662,N_8594,N_8572);
or U8663 (N_8663,N_8575,N_8550);
and U8664 (N_8664,N_8525,N_8562);
nand U8665 (N_8665,N_8519,N_8520);
or U8666 (N_8666,N_8534,N_8532);
or U8667 (N_8667,N_8523,N_8503);
nand U8668 (N_8668,N_8550,N_8565);
nand U8669 (N_8669,N_8533,N_8504);
or U8670 (N_8670,N_8574,N_8521);
nand U8671 (N_8671,N_8590,N_8551);
or U8672 (N_8672,N_8552,N_8589);
nand U8673 (N_8673,N_8582,N_8571);
or U8674 (N_8674,N_8555,N_8559);
and U8675 (N_8675,N_8568,N_8598);
nor U8676 (N_8676,N_8578,N_8521);
or U8677 (N_8677,N_8501,N_8532);
nor U8678 (N_8678,N_8506,N_8594);
nand U8679 (N_8679,N_8516,N_8551);
and U8680 (N_8680,N_8589,N_8545);
nand U8681 (N_8681,N_8536,N_8570);
and U8682 (N_8682,N_8513,N_8557);
and U8683 (N_8683,N_8521,N_8516);
or U8684 (N_8684,N_8589,N_8551);
or U8685 (N_8685,N_8539,N_8557);
nor U8686 (N_8686,N_8591,N_8587);
and U8687 (N_8687,N_8578,N_8509);
nor U8688 (N_8688,N_8527,N_8582);
nor U8689 (N_8689,N_8518,N_8514);
nand U8690 (N_8690,N_8542,N_8592);
xor U8691 (N_8691,N_8517,N_8558);
nand U8692 (N_8692,N_8571,N_8536);
and U8693 (N_8693,N_8580,N_8573);
and U8694 (N_8694,N_8571,N_8501);
and U8695 (N_8695,N_8562,N_8578);
nor U8696 (N_8696,N_8574,N_8595);
or U8697 (N_8697,N_8550,N_8595);
nor U8698 (N_8698,N_8563,N_8514);
nor U8699 (N_8699,N_8573,N_8501);
and U8700 (N_8700,N_8690,N_8610);
nand U8701 (N_8701,N_8615,N_8608);
nand U8702 (N_8702,N_8694,N_8698);
xnor U8703 (N_8703,N_8679,N_8631);
nor U8704 (N_8704,N_8637,N_8685);
nand U8705 (N_8705,N_8645,N_8624);
nand U8706 (N_8706,N_8693,N_8646);
or U8707 (N_8707,N_8620,N_8648);
nor U8708 (N_8708,N_8614,N_8670);
and U8709 (N_8709,N_8621,N_8687);
and U8710 (N_8710,N_8697,N_8618);
or U8711 (N_8711,N_8630,N_8665);
and U8712 (N_8712,N_8611,N_8692);
nor U8713 (N_8713,N_8688,N_8644);
and U8714 (N_8714,N_8617,N_8663);
and U8715 (N_8715,N_8673,N_8683);
and U8716 (N_8716,N_8638,N_8639);
or U8717 (N_8717,N_8666,N_8628);
and U8718 (N_8718,N_8669,N_8604);
and U8719 (N_8719,N_8600,N_8672);
or U8720 (N_8720,N_8625,N_8619);
nand U8721 (N_8721,N_8671,N_8699);
nor U8722 (N_8722,N_8664,N_8634);
or U8723 (N_8723,N_8650,N_8613);
nand U8724 (N_8724,N_8656,N_8653);
nand U8725 (N_8725,N_8636,N_8658);
and U8726 (N_8726,N_8632,N_8643);
and U8727 (N_8727,N_8605,N_8678);
nand U8728 (N_8728,N_8668,N_8675);
or U8729 (N_8729,N_8680,N_8684);
nand U8730 (N_8730,N_8640,N_8662);
and U8731 (N_8731,N_8616,N_8695);
and U8732 (N_8732,N_8626,N_8682);
nand U8733 (N_8733,N_8603,N_8681);
or U8734 (N_8734,N_8623,N_8609);
nand U8735 (N_8735,N_8602,N_8696);
or U8736 (N_8736,N_8660,N_8654);
nor U8737 (N_8737,N_8661,N_8659);
or U8738 (N_8738,N_8633,N_8607);
and U8739 (N_8739,N_8622,N_8635);
or U8740 (N_8740,N_8691,N_8647);
nand U8741 (N_8741,N_8686,N_8627);
nor U8742 (N_8742,N_8655,N_8657);
or U8743 (N_8743,N_8677,N_8674);
or U8744 (N_8744,N_8689,N_8667);
and U8745 (N_8745,N_8642,N_8606);
and U8746 (N_8746,N_8652,N_8641);
and U8747 (N_8747,N_8629,N_8649);
nor U8748 (N_8748,N_8676,N_8612);
or U8749 (N_8749,N_8651,N_8601);
nor U8750 (N_8750,N_8617,N_8606);
and U8751 (N_8751,N_8633,N_8649);
nor U8752 (N_8752,N_8658,N_8681);
nor U8753 (N_8753,N_8698,N_8622);
and U8754 (N_8754,N_8665,N_8642);
nor U8755 (N_8755,N_8662,N_8652);
and U8756 (N_8756,N_8635,N_8676);
or U8757 (N_8757,N_8644,N_8675);
and U8758 (N_8758,N_8610,N_8628);
nor U8759 (N_8759,N_8689,N_8690);
xnor U8760 (N_8760,N_8659,N_8656);
or U8761 (N_8761,N_8684,N_8652);
or U8762 (N_8762,N_8649,N_8662);
or U8763 (N_8763,N_8657,N_8685);
nand U8764 (N_8764,N_8613,N_8609);
nand U8765 (N_8765,N_8684,N_8687);
nor U8766 (N_8766,N_8698,N_8666);
nand U8767 (N_8767,N_8629,N_8662);
or U8768 (N_8768,N_8641,N_8688);
xor U8769 (N_8769,N_8612,N_8602);
xnor U8770 (N_8770,N_8656,N_8687);
or U8771 (N_8771,N_8694,N_8693);
nor U8772 (N_8772,N_8620,N_8689);
and U8773 (N_8773,N_8680,N_8613);
or U8774 (N_8774,N_8690,N_8682);
nand U8775 (N_8775,N_8624,N_8633);
nand U8776 (N_8776,N_8682,N_8638);
and U8777 (N_8777,N_8690,N_8637);
xnor U8778 (N_8778,N_8637,N_8617);
or U8779 (N_8779,N_8678,N_8619);
and U8780 (N_8780,N_8627,N_8687);
nor U8781 (N_8781,N_8685,N_8610);
and U8782 (N_8782,N_8668,N_8643);
or U8783 (N_8783,N_8688,N_8621);
nor U8784 (N_8784,N_8680,N_8673);
or U8785 (N_8785,N_8672,N_8635);
and U8786 (N_8786,N_8642,N_8650);
nor U8787 (N_8787,N_8613,N_8632);
and U8788 (N_8788,N_8694,N_8697);
and U8789 (N_8789,N_8699,N_8625);
nand U8790 (N_8790,N_8676,N_8641);
and U8791 (N_8791,N_8625,N_8648);
nor U8792 (N_8792,N_8650,N_8637);
nand U8793 (N_8793,N_8616,N_8673);
and U8794 (N_8794,N_8609,N_8691);
nand U8795 (N_8795,N_8698,N_8612);
and U8796 (N_8796,N_8659,N_8681);
xor U8797 (N_8797,N_8639,N_8601);
or U8798 (N_8798,N_8602,N_8673);
or U8799 (N_8799,N_8658,N_8614);
and U8800 (N_8800,N_8784,N_8736);
and U8801 (N_8801,N_8775,N_8789);
or U8802 (N_8802,N_8707,N_8730);
nand U8803 (N_8803,N_8710,N_8734);
nor U8804 (N_8804,N_8791,N_8798);
or U8805 (N_8805,N_8754,N_8708);
and U8806 (N_8806,N_8751,N_8711);
nand U8807 (N_8807,N_8735,N_8753);
nor U8808 (N_8808,N_8780,N_8704);
or U8809 (N_8809,N_8700,N_8769);
or U8810 (N_8810,N_8746,N_8726);
xnor U8811 (N_8811,N_8758,N_8783);
or U8812 (N_8812,N_8721,N_8712);
or U8813 (N_8813,N_8778,N_8706);
or U8814 (N_8814,N_8703,N_8781);
nor U8815 (N_8815,N_8755,N_8748);
and U8816 (N_8816,N_8779,N_8722);
nand U8817 (N_8817,N_8796,N_8720);
and U8818 (N_8818,N_8770,N_8794);
nand U8819 (N_8819,N_8756,N_8714);
and U8820 (N_8820,N_8709,N_8719);
and U8821 (N_8821,N_8749,N_8725);
and U8822 (N_8822,N_8795,N_8782);
or U8823 (N_8823,N_8718,N_8763);
or U8824 (N_8824,N_8760,N_8792);
or U8825 (N_8825,N_8768,N_8728);
nor U8826 (N_8826,N_8771,N_8793);
xor U8827 (N_8827,N_8765,N_8799);
or U8828 (N_8828,N_8797,N_8786);
and U8829 (N_8829,N_8713,N_8729);
nor U8830 (N_8830,N_8705,N_8752);
and U8831 (N_8831,N_8739,N_8731);
or U8832 (N_8832,N_8742,N_8750);
or U8833 (N_8833,N_8774,N_8741);
nand U8834 (N_8834,N_8716,N_8740);
and U8835 (N_8835,N_8747,N_8788);
nor U8836 (N_8836,N_8787,N_8764);
and U8837 (N_8837,N_8724,N_8702);
and U8838 (N_8838,N_8772,N_8727);
and U8839 (N_8839,N_8759,N_8776);
nand U8840 (N_8840,N_8701,N_8732);
nand U8841 (N_8841,N_8785,N_8767);
nand U8842 (N_8842,N_8790,N_8757);
nor U8843 (N_8843,N_8766,N_8762);
nor U8844 (N_8844,N_8744,N_8723);
nand U8845 (N_8845,N_8733,N_8715);
and U8846 (N_8846,N_8761,N_8717);
or U8847 (N_8847,N_8738,N_8773);
or U8848 (N_8848,N_8745,N_8777);
and U8849 (N_8849,N_8737,N_8743);
nand U8850 (N_8850,N_8742,N_8710);
nor U8851 (N_8851,N_8773,N_8755);
or U8852 (N_8852,N_8728,N_8749);
or U8853 (N_8853,N_8717,N_8769);
nor U8854 (N_8854,N_8729,N_8719);
or U8855 (N_8855,N_8727,N_8766);
nor U8856 (N_8856,N_8767,N_8729);
and U8857 (N_8857,N_8775,N_8784);
nand U8858 (N_8858,N_8794,N_8717);
nand U8859 (N_8859,N_8767,N_8704);
nand U8860 (N_8860,N_8767,N_8757);
or U8861 (N_8861,N_8728,N_8706);
or U8862 (N_8862,N_8771,N_8715);
xor U8863 (N_8863,N_8788,N_8728);
or U8864 (N_8864,N_8777,N_8778);
nor U8865 (N_8865,N_8798,N_8706);
nor U8866 (N_8866,N_8707,N_8728);
nor U8867 (N_8867,N_8786,N_8749);
and U8868 (N_8868,N_8782,N_8764);
nand U8869 (N_8869,N_8765,N_8775);
or U8870 (N_8870,N_8741,N_8710);
nand U8871 (N_8871,N_8776,N_8741);
or U8872 (N_8872,N_8726,N_8776);
or U8873 (N_8873,N_8720,N_8763);
and U8874 (N_8874,N_8720,N_8759);
or U8875 (N_8875,N_8783,N_8731);
or U8876 (N_8876,N_8734,N_8790);
nor U8877 (N_8877,N_8793,N_8720);
nor U8878 (N_8878,N_8789,N_8778);
or U8879 (N_8879,N_8737,N_8751);
and U8880 (N_8880,N_8731,N_8732);
nor U8881 (N_8881,N_8774,N_8739);
and U8882 (N_8882,N_8780,N_8795);
and U8883 (N_8883,N_8722,N_8720);
nor U8884 (N_8884,N_8746,N_8778);
or U8885 (N_8885,N_8720,N_8771);
nor U8886 (N_8886,N_8707,N_8788);
xor U8887 (N_8887,N_8795,N_8770);
or U8888 (N_8888,N_8785,N_8792);
or U8889 (N_8889,N_8770,N_8720);
or U8890 (N_8890,N_8757,N_8717);
or U8891 (N_8891,N_8772,N_8751);
nand U8892 (N_8892,N_8716,N_8783);
and U8893 (N_8893,N_8700,N_8701);
nand U8894 (N_8894,N_8720,N_8749);
and U8895 (N_8895,N_8739,N_8782);
nor U8896 (N_8896,N_8775,N_8774);
or U8897 (N_8897,N_8773,N_8705);
nand U8898 (N_8898,N_8708,N_8780);
nand U8899 (N_8899,N_8734,N_8760);
nor U8900 (N_8900,N_8856,N_8853);
nand U8901 (N_8901,N_8817,N_8868);
or U8902 (N_8902,N_8863,N_8801);
and U8903 (N_8903,N_8880,N_8804);
or U8904 (N_8904,N_8811,N_8845);
or U8905 (N_8905,N_8821,N_8806);
and U8906 (N_8906,N_8892,N_8897);
and U8907 (N_8907,N_8859,N_8814);
nand U8908 (N_8908,N_8866,N_8839);
nor U8909 (N_8909,N_8864,N_8881);
or U8910 (N_8910,N_8875,N_8871);
nor U8911 (N_8911,N_8837,N_8883);
nand U8912 (N_8912,N_8832,N_8886);
nor U8913 (N_8913,N_8885,N_8812);
nand U8914 (N_8914,N_8869,N_8838);
nand U8915 (N_8915,N_8895,N_8808);
and U8916 (N_8916,N_8825,N_8860);
xnor U8917 (N_8917,N_8867,N_8873);
or U8918 (N_8918,N_8848,N_8815);
nand U8919 (N_8919,N_8849,N_8876);
or U8920 (N_8920,N_8861,N_8822);
nand U8921 (N_8921,N_8857,N_8833);
or U8922 (N_8922,N_8851,N_8888);
and U8923 (N_8923,N_8800,N_8810);
and U8924 (N_8924,N_8835,N_8834);
nor U8925 (N_8925,N_8803,N_8844);
and U8926 (N_8926,N_8893,N_8846);
nor U8927 (N_8927,N_8840,N_8874);
or U8928 (N_8928,N_8850,N_8865);
or U8929 (N_8929,N_8802,N_8836);
nand U8930 (N_8930,N_8805,N_8898);
nand U8931 (N_8931,N_8824,N_8855);
xor U8932 (N_8932,N_8852,N_8819);
or U8933 (N_8933,N_8807,N_8843);
or U8934 (N_8934,N_8847,N_8884);
and U8935 (N_8935,N_8870,N_8896);
and U8936 (N_8936,N_8809,N_8887);
xor U8937 (N_8937,N_8889,N_8854);
xor U8938 (N_8938,N_8826,N_8899);
nor U8939 (N_8939,N_8842,N_8894);
nor U8940 (N_8940,N_8828,N_8877);
nand U8941 (N_8941,N_8818,N_8872);
and U8942 (N_8942,N_8827,N_8813);
nor U8943 (N_8943,N_8820,N_8831);
nand U8944 (N_8944,N_8882,N_8879);
nand U8945 (N_8945,N_8862,N_8878);
or U8946 (N_8946,N_8858,N_8830);
nand U8947 (N_8947,N_8829,N_8841);
and U8948 (N_8948,N_8890,N_8816);
nor U8949 (N_8949,N_8823,N_8891);
or U8950 (N_8950,N_8825,N_8887);
nand U8951 (N_8951,N_8832,N_8867);
nor U8952 (N_8952,N_8875,N_8884);
or U8953 (N_8953,N_8860,N_8861);
nor U8954 (N_8954,N_8892,N_8832);
xnor U8955 (N_8955,N_8896,N_8808);
xor U8956 (N_8956,N_8843,N_8887);
or U8957 (N_8957,N_8817,N_8810);
or U8958 (N_8958,N_8897,N_8873);
nor U8959 (N_8959,N_8884,N_8881);
nand U8960 (N_8960,N_8886,N_8838);
nand U8961 (N_8961,N_8840,N_8847);
or U8962 (N_8962,N_8886,N_8808);
or U8963 (N_8963,N_8811,N_8816);
and U8964 (N_8964,N_8890,N_8833);
or U8965 (N_8965,N_8842,N_8833);
nor U8966 (N_8966,N_8866,N_8850);
or U8967 (N_8967,N_8861,N_8812);
nand U8968 (N_8968,N_8816,N_8858);
nor U8969 (N_8969,N_8860,N_8898);
nand U8970 (N_8970,N_8852,N_8823);
nand U8971 (N_8971,N_8894,N_8841);
and U8972 (N_8972,N_8887,N_8842);
and U8973 (N_8973,N_8883,N_8811);
nand U8974 (N_8974,N_8847,N_8898);
and U8975 (N_8975,N_8833,N_8883);
nand U8976 (N_8976,N_8835,N_8878);
nand U8977 (N_8977,N_8838,N_8896);
and U8978 (N_8978,N_8828,N_8829);
nor U8979 (N_8979,N_8822,N_8827);
or U8980 (N_8980,N_8817,N_8842);
or U8981 (N_8981,N_8801,N_8800);
or U8982 (N_8982,N_8852,N_8836);
xor U8983 (N_8983,N_8872,N_8809);
nand U8984 (N_8984,N_8841,N_8879);
and U8985 (N_8985,N_8802,N_8814);
nand U8986 (N_8986,N_8818,N_8823);
and U8987 (N_8987,N_8810,N_8869);
nor U8988 (N_8988,N_8828,N_8823);
or U8989 (N_8989,N_8818,N_8897);
and U8990 (N_8990,N_8857,N_8866);
nand U8991 (N_8991,N_8897,N_8864);
nand U8992 (N_8992,N_8862,N_8853);
nand U8993 (N_8993,N_8869,N_8855);
nor U8994 (N_8994,N_8879,N_8885);
nand U8995 (N_8995,N_8888,N_8821);
or U8996 (N_8996,N_8870,N_8814);
nor U8997 (N_8997,N_8885,N_8810);
and U8998 (N_8998,N_8829,N_8827);
and U8999 (N_8999,N_8876,N_8861);
or U9000 (N_9000,N_8969,N_8981);
nor U9001 (N_9001,N_8960,N_8950);
or U9002 (N_9002,N_8921,N_8966);
nand U9003 (N_9003,N_8935,N_8991);
nand U9004 (N_9004,N_8961,N_8962);
or U9005 (N_9005,N_8920,N_8913);
and U9006 (N_9006,N_8941,N_8959);
nor U9007 (N_9007,N_8994,N_8933);
and U9008 (N_9008,N_8971,N_8903);
and U9009 (N_9009,N_8942,N_8964);
or U9010 (N_9010,N_8987,N_8939);
nand U9011 (N_9011,N_8990,N_8974);
nand U9012 (N_9012,N_8914,N_8984);
and U9013 (N_9013,N_8926,N_8992);
or U9014 (N_9014,N_8937,N_8980);
or U9015 (N_9015,N_8965,N_8997);
and U9016 (N_9016,N_8955,N_8931);
and U9017 (N_9017,N_8949,N_8934);
or U9018 (N_9018,N_8976,N_8917);
and U9019 (N_9019,N_8975,N_8911);
nor U9020 (N_9020,N_8948,N_8982);
nand U9021 (N_9021,N_8954,N_8916);
and U9022 (N_9022,N_8938,N_8958);
nor U9023 (N_9023,N_8918,N_8972);
or U9024 (N_9024,N_8929,N_8944);
or U9025 (N_9025,N_8977,N_8996);
nor U9026 (N_9026,N_8907,N_8956);
nor U9027 (N_9027,N_8973,N_8932);
nand U9028 (N_9028,N_8989,N_8923);
or U9029 (N_9029,N_8922,N_8925);
or U9030 (N_9030,N_8995,N_8908);
or U9031 (N_9031,N_8909,N_8983);
nand U9032 (N_9032,N_8986,N_8985);
nor U9033 (N_9033,N_8936,N_8940);
and U9034 (N_9034,N_8912,N_8953);
nand U9035 (N_9035,N_8915,N_8901);
or U9036 (N_9036,N_8945,N_8963);
nand U9037 (N_9037,N_8970,N_8947);
nor U9038 (N_9038,N_8930,N_8967);
nand U9039 (N_9039,N_8946,N_8999);
xnor U9040 (N_9040,N_8943,N_8904);
nor U9041 (N_9041,N_8951,N_8902);
nor U9042 (N_9042,N_8906,N_8900);
nand U9043 (N_9043,N_8952,N_8927);
nand U9044 (N_9044,N_8905,N_8910);
nand U9045 (N_9045,N_8919,N_8924);
nand U9046 (N_9046,N_8957,N_8998);
and U9047 (N_9047,N_8993,N_8928);
or U9048 (N_9048,N_8978,N_8979);
or U9049 (N_9049,N_8968,N_8988);
nand U9050 (N_9050,N_8986,N_8961);
and U9051 (N_9051,N_8966,N_8960);
or U9052 (N_9052,N_8955,N_8942);
nand U9053 (N_9053,N_8957,N_8936);
and U9054 (N_9054,N_8984,N_8982);
and U9055 (N_9055,N_8990,N_8925);
nand U9056 (N_9056,N_8981,N_8948);
and U9057 (N_9057,N_8912,N_8924);
nand U9058 (N_9058,N_8904,N_8969);
nor U9059 (N_9059,N_8960,N_8935);
nand U9060 (N_9060,N_8957,N_8953);
nor U9061 (N_9061,N_8995,N_8952);
nand U9062 (N_9062,N_8971,N_8946);
and U9063 (N_9063,N_8917,N_8911);
and U9064 (N_9064,N_8916,N_8926);
and U9065 (N_9065,N_8938,N_8937);
or U9066 (N_9066,N_8983,N_8961);
nand U9067 (N_9067,N_8935,N_8921);
nand U9068 (N_9068,N_8925,N_8933);
nor U9069 (N_9069,N_8973,N_8903);
or U9070 (N_9070,N_8904,N_8926);
nand U9071 (N_9071,N_8919,N_8934);
or U9072 (N_9072,N_8960,N_8951);
and U9073 (N_9073,N_8908,N_8948);
and U9074 (N_9074,N_8991,N_8979);
xor U9075 (N_9075,N_8911,N_8945);
nor U9076 (N_9076,N_8946,N_8987);
nor U9077 (N_9077,N_8916,N_8935);
nor U9078 (N_9078,N_8967,N_8943);
or U9079 (N_9079,N_8928,N_8910);
or U9080 (N_9080,N_8981,N_8980);
and U9081 (N_9081,N_8929,N_8994);
and U9082 (N_9082,N_8954,N_8902);
nor U9083 (N_9083,N_8974,N_8978);
or U9084 (N_9084,N_8972,N_8935);
nand U9085 (N_9085,N_8911,N_8920);
and U9086 (N_9086,N_8957,N_8952);
or U9087 (N_9087,N_8966,N_8986);
and U9088 (N_9088,N_8910,N_8975);
nor U9089 (N_9089,N_8917,N_8910);
or U9090 (N_9090,N_8914,N_8910);
and U9091 (N_9091,N_8948,N_8985);
nor U9092 (N_9092,N_8960,N_8990);
and U9093 (N_9093,N_8965,N_8995);
or U9094 (N_9094,N_8920,N_8914);
nor U9095 (N_9095,N_8911,N_8924);
or U9096 (N_9096,N_8925,N_8978);
nor U9097 (N_9097,N_8997,N_8964);
or U9098 (N_9098,N_8913,N_8953);
nor U9099 (N_9099,N_8990,N_8955);
nor U9100 (N_9100,N_9090,N_9087);
nor U9101 (N_9101,N_9064,N_9020);
or U9102 (N_9102,N_9081,N_9018);
or U9103 (N_9103,N_9010,N_9000);
nand U9104 (N_9104,N_9097,N_9037);
nand U9105 (N_9105,N_9013,N_9095);
nand U9106 (N_9106,N_9016,N_9041);
nor U9107 (N_9107,N_9091,N_9039);
nor U9108 (N_9108,N_9014,N_9038);
or U9109 (N_9109,N_9035,N_9077);
nand U9110 (N_9110,N_9063,N_9099);
or U9111 (N_9111,N_9061,N_9034);
or U9112 (N_9112,N_9055,N_9056);
or U9113 (N_9113,N_9044,N_9006);
xor U9114 (N_9114,N_9030,N_9031);
and U9115 (N_9115,N_9001,N_9052);
or U9116 (N_9116,N_9096,N_9040);
nor U9117 (N_9117,N_9043,N_9008);
nand U9118 (N_9118,N_9088,N_9015);
nand U9119 (N_9119,N_9082,N_9066);
nor U9120 (N_9120,N_9046,N_9042);
or U9121 (N_9121,N_9032,N_9069);
nand U9122 (N_9122,N_9024,N_9048);
nor U9123 (N_9123,N_9050,N_9002);
or U9124 (N_9124,N_9026,N_9054);
nor U9125 (N_9125,N_9084,N_9049);
or U9126 (N_9126,N_9098,N_9004);
or U9127 (N_9127,N_9071,N_9047);
nand U9128 (N_9128,N_9027,N_9058);
and U9129 (N_9129,N_9089,N_9073);
or U9130 (N_9130,N_9068,N_9005);
or U9131 (N_9131,N_9060,N_9028);
and U9132 (N_9132,N_9075,N_9009);
or U9133 (N_9133,N_9007,N_9080);
nor U9134 (N_9134,N_9053,N_9059);
and U9135 (N_9135,N_9093,N_9057);
nor U9136 (N_9136,N_9094,N_9012);
or U9137 (N_9137,N_9074,N_9062);
and U9138 (N_9138,N_9036,N_9083);
nor U9139 (N_9139,N_9011,N_9086);
nor U9140 (N_9140,N_9065,N_9070);
nor U9141 (N_9141,N_9025,N_9019);
nand U9142 (N_9142,N_9085,N_9045);
nor U9143 (N_9143,N_9022,N_9072);
or U9144 (N_9144,N_9051,N_9003);
nand U9145 (N_9145,N_9033,N_9023);
and U9146 (N_9146,N_9078,N_9067);
and U9147 (N_9147,N_9092,N_9079);
and U9148 (N_9148,N_9029,N_9017);
nand U9149 (N_9149,N_9076,N_9021);
or U9150 (N_9150,N_9036,N_9060);
and U9151 (N_9151,N_9002,N_9044);
nand U9152 (N_9152,N_9026,N_9041);
and U9153 (N_9153,N_9007,N_9084);
or U9154 (N_9154,N_9098,N_9070);
and U9155 (N_9155,N_9020,N_9067);
nor U9156 (N_9156,N_9014,N_9003);
and U9157 (N_9157,N_9093,N_9023);
or U9158 (N_9158,N_9006,N_9075);
or U9159 (N_9159,N_9096,N_9086);
xor U9160 (N_9160,N_9019,N_9099);
or U9161 (N_9161,N_9034,N_9060);
and U9162 (N_9162,N_9062,N_9050);
nor U9163 (N_9163,N_9030,N_9083);
xnor U9164 (N_9164,N_9010,N_9015);
nand U9165 (N_9165,N_9072,N_9045);
nor U9166 (N_9166,N_9041,N_9029);
nand U9167 (N_9167,N_9098,N_9036);
and U9168 (N_9168,N_9032,N_9018);
and U9169 (N_9169,N_9091,N_9005);
and U9170 (N_9170,N_9009,N_9014);
nor U9171 (N_9171,N_9053,N_9010);
or U9172 (N_9172,N_9053,N_9028);
or U9173 (N_9173,N_9077,N_9088);
and U9174 (N_9174,N_9061,N_9052);
nor U9175 (N_9175,N_9012,N_9029);
or U9176 (N_9176,N_9091,N_9027);
nor U9177 (N_9177,N_9084,N_9025);
and U9178 (N_9178,N_9024,N_9056);
and U9179 (N_9179,N_9031,N_9042);
or U9180 (N_9180,N_9097,N_9015);
nand U9181 (N_9181,N_9080,N_9069);
and U9182 (N_9182,N_9010,N_9038);
or U9183 (N_9183,N_9038,N_9081);
or U9184 (N_9184,N_9067,N_9099);
nor U9185 (N_9185,N_9072,N_9083);
nor U9186 (N_9186,N_9044,N_9068);
and U9187 (N_9187,N_9026,N_9015);
nand U9188 (N_9188,N_9091,N_9094);
and U9189 (N_9189,N_9030,N_9029);
nand U9190 (N_9190,N_9095,N_9019);
or U9191 (N_9191,N_9075,N_9011);
or U9192 (N_9192,N_9085,N_9094);
nand U9193 (N_9193,N_9037,N_9035);
or U9194 (N_9194,N_9065,N_9003);
and U9195 (N_9195,N_9065,N_9082);
nand U9196 (N_9196,N_9004,N_9093);
nand U9197 (N_9197,N_9065,N_9013);
or U9198 (N_9198,N_9075,N_9039);
xnor U9199 (N_9199,N_9052,N_9042);
or U9200 (N_9200,N_9142,N_9138);
nand U9201 (N_9201,N_9106,N_9197);
or U9202 (N_9202,N_9193,N_9195);
nand U9203 (N_9203,N_9181,N_9169);
or U9204 (N_9204,N_9135,N_9100);
or U9205 (N_9205,N_9148,N_9118);
and U9206 (N_9206,N_9149,N_9122);
nor U9207 (N_9207,N_9176,N_9133);
nand U9208 (N_9208,N_9196,N_9105);
nor U9209 (N_9209,N_9199,N_9154);
nand U9210 (N_9210,N_9109,N_9175);
nor U9211 (N_9211,N_9143,N_9136);
nand U9212 (N_9212,N_9180,N_9139);
and U9213 (N_9213,N_9185,N_9117);
nand U9214 (N_9214,N_9187,N_9165);
xnor U9215 (N_9215,N_9146,N_9152);
nor U9216 (N_9216,N_9194,N_9102);
or U9217 (N_9217,N_9128,N_9107);
nand U9218 (N_9218,N_9191,N_9160);
nand U9219 (N_9219,N_9127,N_9171);
nor U9220 (N_9220,N_9140,N_9132);
nand U9221 (N_9221,N_9120,N_9111);
nand U9222 (N_9222,N_9147,N_9151);
xor U9223 (N_9223,N_9115,N_9108);
nand U9224 (N_9224,N_9110,N_9178);
nor U9225 (N_9225,N_9101,N_9119);
nor U9226 (N_9226,N_9144,N_9159);
or U9227 (N_9227,N_9153,N_9186);
nor U9228 (N_9228,N_9188,N_9131);
or U9229 (N_9229,N_9156,N_9112);
nor U9230 (N_9230,N_9182,N_9150);
nor U9231 (N_9231,N_9104,N_9123);
or U9232 (N_9232,N_9141,N_9189);
and U9233 (N_9233,N_9164,N_9125);
or U9234 (N_9234,N_9179,N_9158);
and U9235 (N_9235,N_9163,N_9137);
or U9236 (N_9236,N_9198,N_9130);
or U9237 (N_9237,N_9121,N_9103);
nor U9238 (N_9238,N_9190,N_9177);
nor U9239 (N_9239,N_9172,N_9174);
nand U9240 (N_9240,N_9173,N_9116);
nand U9241 (N_9241,N_9157,N_9162);
nand U9242 (N_9242,N_9168,N_9126);
and U9243 (N_9243,N_9124,N_9134);
and U9244 (N_9244,N_9167,N_9155);
nor U9245 (N_9245,N_9170,N_9183);
nand U9246 (N_9246,N_9161,N_9192);
xnor U9247 (N_9247,N_9145,N_9113);
nor U9248 (N_9248,N_9166,N_9184);
nor U9249 (N_9249,N_9114,N_9129);
and U9250 (N_9250,N_9135,N_9164);
nor U9251 (N_9251,N_9167,N_9151);
and U9252 (N_9252,N_9176,N_9165);
and U9253 (N_9253,N_9104,N_9147);
nand U9254 (N_9254,N_9175,N_9121);
nor U9255 (N_9255,N_9120,N_9130);
and U9256 (N_9256,N_9150,N_9165);
nor U9257 (N_9257,N_9150,N_9121);
nor U9258 (N_9258,N_9176,N_9127);
and U9259 (N_9259,N_9149,N_9151);
nor U9260 (N_9260,N_9183,N_9102);
nand U9261 (N_9261,N_9127,N_9157);
nand U9262 (N_9262,N_9172,N_9104);
nor U9263 (N_9263,N_9104,N_9134);
nand U9264 (N_9264,N_9172,N_9134);
nand U9265 (N_9265,N_9184,N_9104);
and U9266 (N_9266,N_9192,N_9196);
nand U9267 (N_9267,N_9125,N_9177);
nand U9268 (N_9268,N_9189,N_9195);
nand U9269 (N_9269,N_9128,N_9122);
or U9270 (N_9270,N_9130,N_9167);
and U9271 (N_9271,N_9162,N_9132);
and U9272 (N_9272,N_9114,N_9123);
and U9273 (N_9273,N_9192,N_9199);
and U9274 (N_9274,N_9144,N_9119);
nand U9275 (N_9275,N_9197,N_9125);
or U9276 (N_9276,N_9107,N_9163);
or U9277 (N_9277,N_9138,N_9102);
or U9278 (N_9278,N_9140,N_9136);
nand U9279 (N_9279,N_9111,N_9161);
nand U9280 (N_9280,N_9185,N_9193);
and U9281 (N_9281,N_9195,N_9106);
and U9282 (N_9282,N_9186,N_9108);
or U9283 (N_9283,N_9159,N_9197);
and U9284 (N_9284,N_9174,N_9183);
nor U9285 (N_9285,N_9118,N_9157);
or U9286 (N_9286,N_9162,N_9116);
or U9287 (N_9287,N_9175,N_9179);
nand U9288 (N_9288,N_9153,N_9136);
nor U9289 (N_9289,N_9176,N_9153);
nand U9290 (N_9290,N_9174,N_9140);
nand U9291 (N_9291,N_9113,N_9143);
nand U9292 (N_9292,N_9119,N_9135);
nand U9293 (N_9293,N_9122,N_9167);
nor U9294 (N_9294,N_9132,N_9198);
nand U9295 (N_9295,N_9145,N_9148);
or U9296 (N_9296,N_9152,N_9185);
nor U9297 (N_9297,N_9160,N_9131);
nor U9298 (N_9298,N_9133,N_9166);
nor U9299 (N_9299,N_9148,N_9199);
nand U9300 (N_9300,N_9239,N_9286);
nor U9301 (N_9301,N_9292,N_9223);
or U9302 (N_9302,N_9285,N_9244);
nand U9303 (N_9303,N_9284,N_9289);
and U9304 (N_9304,N_9237,N_9235);
and U9305 (N_9305,N_9218,N_9249);
and U9306 (N_9306,N_9280,N_9236);
or U9307 (N_9307,N_9206,N_9202);
or U9308 (N_9308,N_9271,N_9219);
nand U9309 (N_9309,N_9291,N_9261);
or U9310 (N_9310,N_9293,N_9201);
or U9311 (N_9311,N_9262,N_9257);
and U9312 (N_9312,N_9273,N_9264);
nor U9313 (N_9313,N_9252,N_9298);
nor U9314 (N_9314,N_9258,N_9242);
and U9315 (N_9315,N_9296,N_9200);
and U9316 (N_9316,N_9234,N_9294);
nand U9317 (N_9317,N_9255,N_9259);
and U9318 (N_9318,N_9208,N_9212);
nor U9319 (N_9319,N_9213,N_9220);
and U9320 (N_9320,N_9299,N_9278);
xnor U9321 (N_9321,N_9229,N_9226);
or U9322 (N_9322,N_9251,N_9211);
nand U9323 (N_9323,N_9222,N_9221);
xnor U9324 (N_9324,N_9279,N_9297);
and U9325 (N_9325,N_9287,N_9240);
nor U9326 (N_9326,N_9267,N_9241);
or U9327 (N_9327,N_9243,N_9276);
nor U9328 (N_9328,N_9204,N_9225);
nor U9329 (N_9329,N_9248,N_9283);
and U9330 (N_9330,N_9269,N_9270);
nand U9331 (N_9331,N_9214,N_9233);
or U9332 (N_9332,N_9231,N_9209);
and U9333 (N_9333,N_9228,N_9247);
nor U9334 (N_9334,N_9272,N_9246);
and U9335 (N_9335,N_9203,N_9230);
and U9336 (N_9336,N_9224,N_9205);
nand U9337 (N_9337,N_9245,N_9282);
and U9338 (N_9338,N_9265,N_9215);
nand U9339 (N_9339,N_9295,N_9217);
nand U9340 (N_9340,N_9281,N_9275);
and U9341 (N_9341,N_9266,N_9274);
nand U9342 (N_9342,N_9210,N_9227);
nor U9343 (N_9343,N_9256,N_9216);
or U9344 (N_9344,N_9268,N_9250);
nand U9345 (N_9345,N_9238,N_9263);
nand U9346 (N_9346,N_9253,N_9288);
or U9347 (N_9347,N_9290,N_9254);
or U9348 (N_9348,N_9260,N_9207);
nand U9349 (N_9349,N_9277,N_9232);
nor U9350 (N_9350,N_9253,N_9216);
nor U9351 (N_9351,N_9202,N_9264);
or U9352 (N_9352,N_9293,N_9256);
nor U9353 (N_9353,N_9233,N_9267);
nand U9354 (N_9354,N_9299,N_9231);
and U9355 (N_9355,N_9230,N_9265);
nand U9356 (N_9356,N_9247,N_9218);
and U9357 (N_9357,N_9248,N_9208);
nor U9358 (N_9358,N_9204,N_9208);
nor U9359 (N_9359,N_9233,N_9282);
nor U9360 (N_9360,N_9214,N_9262);
or U9361 (N_9361,N_9247,N_9293);
nor U9362 (N_9362,N_9215,N_9289);
and U9363 (N_9363,N_9293,N_9271);
and U9364 (N_9364,N_9288,N_9238);
nor U9365 (N_9365,N_9235,N_9251);
or U9366 (N_9366,N_9295,N_9297);
nor U9367 (N_9367,N_9290,N_9253);
or U9368 (N_9368,N_9256,N_9229);
xnor U9369 (N_9369,N_9298,N_9218);
and U9370 (N_9370,N_9278,N_9254);
and U9371 (N_9371,N_9238,N_9229);
xor U9372 (N_9372,N_9248,N_9211);
and U9373 (N_9373,N_9275,N_9254);
or U9374 (N_9374,N_9287,N_9246);
nor U9375 (N_9375,N_9237,N_9222);
nor U9376 (N_9376,N_9219,N_9229);
or U9377 (N_9377,N_9267,N_9290);
nand U9378 (N_9378,N_9278,N_9234);
nor U9379 (N_9379,N_9297,N_9294);
nand U9380 (N_9380,N_9294,N_9265);
and U9381 (N_9381,N_9202,N_9242);
and U9382 (N_9382,N_9202,N_9217);
and U9383 (N_9383,N_9279,N_9214);
or U9384 (N_9384,N_9273,N_9275);
or U9385 (N_9385,N_9291,N_9218);
or U9386 (N_9386,N_9295,N_9220);
nor U9387 (N_9387,N_9227,N_9257);
nand U9388 (N_9388,N_9290,N_9235);
or U9389 (N_9389,N_9285,N_9253);
or U9390 (N_9390,N_9257,N_9237);
and U9391 (N_9391,N_9282,N_9239);
and U9392 (N_9392,N_9223,N_9258);
and U9393 (N_9393,N_9224,N_9272);
or U9394 (N_9394,N_9213,N_9223);
or U9395 (N_9395,N_9203,N_9202);
or U9396 (N_9396,N_9265,N_9220);
or U9397 (N_9397,N_9271,N_9261);
nor U9398 (N_9398,N_9231,N_9234);
and U9399 (N_9399,N_9210,N_9209);
nand U9400 (N_9400,N_9318,N_9386);
or U9401 (N_9401,N_9304,N_9305);
or U9402 (N_9402,N_9359,N_9343);
or U9403 (N_9403,N_9350,N_9302);
nor U9404 (N_9404,N_9332,N_9349);
nand U9405 (N_9405,N_9338,N_9375);
and U9406 (N_9406,N_9394,N_9361);
or U9407 (N_9407,N_9309,N_9320);
nand U9408 (N_9408,N_9388,N_9310);
or U9409 (N_9409,N_9357,N_9348);
nand U9410 (N_9410,N_9328,N_9396);
nor U9411 (N_9411,N_9319,N_9389);
and U9412 (N_9412,N_9303,N_9353);
and U9413 (N_9413,N_9397,N_9365);
nand U9414 (N_9414,N_9399,N_9323);
nand U9415 (N_9415,N_9300,N_9367);
nor U9416 (N_9416,N_9387,N_9314);
nand U9417 (N_9417,N_9313,N_9381);
and U9418 (N_9418,N_9382,N_9390);
nand U9419 (N_9419,N_9373,N_9371);
nor U9420 (N_9420,N_9383,N_9356);
or U9421 (N_9421,N_9307,N_9311);
and U9422 (N_9422,N_9393,N_9329);
and U9423 (N_9423,N_9391,N_9360);
or U9424 (N_9424,N_9363,N_9384);
nor U9425 (N_9425,N_9306,N_9308);
nor U9426 (N_9426,N_9342,N_9326);
and U9427 (N_9427,N_9379,N_9377);
or U9428 (N_9428,N_9370,N_9337);
and U9429 (N_9429,N_9344,N_9358);
and U9430 (N_9430,N_9347,N_9364);
and U9431 (N_9431,N_9336,N_9333);
or U9432 (N_9432,N_9385,N_9335);
or U9433 (N_9433,N_9327,N_9374);
nand U9434 (N_9434,N_9317,N_9315);
nor U9435 (N_9435,N_9378,N_9372);
nand U9436 (N_9436,N_9324,N_9345);
xnor U9437 (N_9437,N_9351,N_9398);
nand U9438 (N_9438,N_9321,N_9352);
or U9439 (N_9439,N_9316,N_9341);
nor U9440 (N_9440,N_9368,N_9301);
or U9441 (N_9441,N_9331,N_9380);
nand U9442 (N_9442,N_9330,N_9339);
or U9443 (N_9443,N_9312,N_9366);
and U9444 (N_9444,N_9376,N_9392);
or U9445 (N_9445,N_9325,N_9346);
xor U9446 (N_9446,N_9322,N_9362);
nor U9447 (N_9447,N_9369,N_9354);
and U9448 (N_9448,N_9340,N_9395);
or U9449 (N_9449,N_9334,N_9355);
and U9450 (N_9450,N_9378,N_9361);
and U9451 (N_9451,N_9348,N_9375);
and U9452 (N_9452,N_9358,N_9327);
nand U9453 (N_9453,N_9300,N_9385);
and U9454 (N_9454,N_9337,N_9357);
or U9455 (N_9455,N_9398,N_9389);
and U9456 (N_9456,N_9306,N_9389);
nand U9457 (N_9457,N_9387,N_9303);
nand U9458 (N_9458,N_9357,N_9352);
nand U9459 (N_9459,N_9383,N_9346);
and U9460 (N_9460,N_9309,N_9354);
or U9461 (N_9461,N_9368,N_9379);
and U9462 (N_9462,N_9381,N_9346);
nor U9463 (N_9463,N_9346,N_9335);
nor U9464 (N_9464,N_9310,N_9306);
nor U9465 (N_9465,N_9335,N_9338);
and U9466 (N_9466,N_9313,N_9314);
nand U9467 (N_9467,N_9389,N_9394);
and U9468 (N_9468,N_9318,N_9335);
xnor U9469 (N_9469,N_9326,N_9314);
and U9470 (N_9470,N_9305,N_9347);
or U9471 (N_9471,N_9319,N_9384);
nand U9472 (N_9472,N_9380,N_9308);
or U9473 (N_9473,N_9386,N_9395);
nor U9474 (N_9474,N_9352,N_9371);
nor U9475 (N_9475,N_9360,N_9384);
nor U9476 (N_9476,N_9349,N_9314);
nand U9477 (N_9477,N_9343,N_9399);
nand U9478 (N_9478,N_9392,N_9355);
and U9479 (N_9479,N_9371,N_9326);
nand U9480 (N_9480,N_9328,N_9321);
or U9481 (N_9481,N_9395,N_9300);
or U9482 (N_9482,N_9393,N_9370);
and U9483 (N_9483,N_9342,N_9358);
nor U9484 (N_9484,N_9342,N_9336);
nor U9485 (N_9485,N_9342,N_9370);
or U9486 (N_9486,N_9381,N_9387);
nand U9487 (N_9487,N_9312,N_9303);
and U9488 (N_9488,N_9318,N_9383);
nand U9489 (N_9489,N_9382,N_9335);
nor U9490 (N_9490,N_9359,N_9350);
and U9491 (N_9491,N_9337,N_9343);
nand U9492 (N_9492,N_9345,N_9333);
nand U9493 (N_9493,N_9344,N_9330);
nor U9494 (N_9494,N_9321,N_9300);
and U9495 (N_9495,N_9335,N_9309);
or U9496 (N_9496,N_9376,N_9358);
and U9497 (N_9497,N_9372,N_9308);
and U9498 (N_9498,N_9356,N_9329);
nor U9499 (N_9499,N_9323,N_9361);
nand U9500 (N_9500,N_9465,N_9483);
nor U9501 (N_9501,N_9494,N_9481);
or U9502 (N_9502,N_9422,N_9408);
or U9503 (N_9503,N_9480,N_9445);
or U9504 (N_9504,N_9491,N_9479);
nand U9505 (N_9505,N_9403,N_9469);
or U9506 (N_9506,N_9471,N_9426);
nor U9507 (N_9507,N_9489,N_9490);
and U9508 (N_9508,N_9427,N_9405);
nand U9509 (N_9509,N_9435,N_9438);
and U9510 (N_9510,N_9410,N_9452);
and U9511 (N_9511,N_9417,N_9448);
nand U9512 (N_9512,N_9460,N_9472);
or U9513 (N_9513,N_9484,N_9461);
or U9514 (N_9514,N_9488,N_9402);
or U9515 (N_9515,N_9433,N_9455);
or U9516 (N_9516,N_9470,N_9486);
xnor U9517 (N_9517,N_9434,N_9428);
or U9518 (N_9518,N_9497,N_9451);
nand U9519 (N_9519,N_9493,N_9464);
nor U9520 (N_9520,N_9456,N_9459);
nand U9521 (N_9521,N_9423,N_9476);
nor U9522 (N_9522,N_9409,N_9412);
nand U9523 (N_9523,N_9466,N_9425);
and U9524 (N_9524,N_9457,N_9413);
nor U9525 (N_9525,N_9404,N_9499);
and U9526 (N_9526,N_9444,N_9416);
nor U9527 (N_9527,N_9496,N_9478);
and U9528 (N_9528,N_9424,N_9421);
or U9529 (N_9529,N_9442,N_9418);
or U9530 (N_9530,N_9437,N_9429);
or U9531 (N_9531,N_9432,N_9482);
xnor U9532 (N_9532,N_9449,N_9458);
and U9533 (N_9533,N_9419,N_9407);
nand U9534 (N_9534,N_9401,N_9411);
nor U9535 (N_9535,N_9443,N_9446);
nor U9536 (N_9536,N_9498,N_9474);
and U9537 (N_9537,N_9431,N_9475);
nand U9538 (N_9538,N_9467,N_9492);
nand U9539 (N_9539,N_9414,N_9454);
or U9540 (N_9540,N_9415,N_9485);
nand U9541 (N_9541,N_9462,N_9447);
and U9542 (N_9542,N_9473,N_9468);
nor U9543 (N_9543,N_9477,N_9420);
and U9544 (N_9544,N_9400,N_9450);
nand U9545 (N_9545,N_9439,N_9453);
nor U9546 (N_9546,N_9436,N_9463);
nand U9547 (N_9547,N_9495,N_9406);
and U9548 (N_9548,N_9440,N_9430);
or U9549 (N_9549,N_9441,N_9487);
nor U9550 (N_9550,N_9455,N_9468);
or U9551 (N_9551,N_9473,N_9417);
or U9552 (N_9552,N_9424,N_9418);
nand U9553 (N_9553,N_9476,N_9420);
nor U9554 (N_9554,N_9437,N_9402);
xor U9555 (N_9555,N_9412,N_9428);
nand U9556 (N_9556,N_9465,N_9485);
nand U9557 (N_9557,N_9462,N_9408);
nand U9558 (N_9558,N_9469,N_9497);
and U9559 (N_9559,N_9433,N_9428);
nand U9560 (N_9560,N_9406,N_9476);
nand U9561 (N_9561,N_9453,N_9458);
or U9562 (N_9562,N_9471,N_9467);
nor U9563 (N_9563,N_9474,N_9438);
and U9564 (N_9564,N_9408,N_9496);
nand U9565 (N_9565,N_9447,N_9451);
and U9566 (N_9566,N_9474,N_9450);
nand U9567 (N_9567,N_9450,N_9478);
nand U9568 (N_9568,N_9420,N_9444);
nor U9569 (N_9569,N_9482,N_9415);
nand U9570 (N_9570,N_9448,N_9461);
nor U9571 (N_9571,N_9477,N_9473);
and U9572 (N_9572,N_9486,N_9477);
or U9573 (N_9573,N_9471,N_9479);
nand U9574 (N_9574,N_9433,N_9426);
or U9575 (N_9575,N_9467,N_9469);
or U9576 (N_9576,N_9418,N_9423);
and U9577 (N_9577,N_9416,N_9439);
and U9578 (N_9578,N_9406,N_9451);
xnor U9579 (N_9579,N_9438,N_9448);
and U9580 (N_9580,N_9452,N_9443);
and U9581 (N_9581,N_9421,N_9478);
and U9582 (N_9582,N_9456,N_9401);
nand U9583 (N_9583,N_9490,N_9406);
nor U9584 (N_9584,N_9431,N_9464);
and U9585 (N_9585,N_9458,N_9491);
nand U9586 (N_9586,N_9431,N_9400);
and U9587 (N_9587,N_9497,N_9459);
nor U9588 (N_9588,N_9421,N_9475);
nor U9589 (N_9589,N_9419,N_9473);
and U9590 (N_9590,N_9460,N_9499);
or U9591 (N_9591,N_9416,N_9426);
and U9592 (N_9592,N_9465,N_9442);
or U9593 (N_9593,N_9412,N_9481);
nand U9594 (N_9594,N_9407,N_9484);
and U9595 (N_9595,N_9439,N_9489);
and U9596 (N_9596,N_9415,N_9466);
nor U9597 (N_9597,N_9401,N_9433);
nand U9598 (N_9598,N_9452,N_9465);
or U9599 (N_9599,N_9402,N_9470);
and U9600 (N_9600,N_9555,N_9557);
or U9601 (N_9601,N_9548,N_9561);
xnor U9602 (N_9602,N_9515,N_9542);
nand U9603 (N_9603,N_9524,N_9559);
or U9604 (N_9604,N_9569,N_9594);
or U9605 (N_9605,N_9523,N_9549);
nand U9606 (N_9606,N_9573,N_9541);
nor U9607 (N_9607,N_9592,N_9575);
or U9608 (N_9608,N_9572,N_9582);
or U9609 (N_9609,N_9584,N_9506);
or U9610 (N_9610,N_9577,N_9505);
nor U9611 (N_9611,N_9564,N_9534);
and U9612 (N_9612,N_9558,N_9586);
nor U9613 (N_9613,N_9585,N_9518);
or U9614 (N_9614,N_9591,N_9512);
xor U9615 (N_9615,N_9526,N_9571);
and U9616 (N_9616,N_9517,N_9508);
nand U9617 (N_9617,N_9513,N_9560);
and U9618 (N_9618,N_9578,N_9597);
or U9619 (N_9619,N_9538,N_9514);
or U9620 (N_9620,N_9570,N_9544);
nand U9621 (N_9621,N_9530,N_9507);
nand U9622 (N_9622,N_9547,N_9503);
or U9623 (N_9623,N_9554,N_9589);
nor U9624 (N_9624,N_9536,N_9567);
nor U9625 (N_9625,N_9562,N_9537);
nor U9626 (N_9626,N_9576,N_9553);
and U9627 (N_9627,N_9504,N_9520);
nand U9628 (N_9628,N_9556,N_9583);
and U9629 (N_9629,N_9516,N_9535);
nand U9630 (N_9630,N_9566,N_9529);
or U9631 (N_9631,N_9579,N_9552);
and U9632 (N_9632,N_9593,N_9580);
or U9633 (N_9633,N_9521,N_9533);
nor U9634 (N_9634,N_9511,N_9590);
and U9635 (N_9635,N_9563,N_9595);
and U9636 (N_9636,N_9598,N_9545);
nand U9637 (N_9637,N_9550,N_9596);
nor U9638 (N_9638,N_9546,N_9588);
and U9639 (N_9639,N_9540,N_9599);
nor U9640 (N_9640,N_9574,N_9587);
and U9641 (N_9641,N_9568,N_9581);
or U9642 (N_9642,N_9543,N_9551);
nand U9643 (N_9643,N_9500,N_9527);
nor U9644 (N_9644,N_9528,N_9519);
nor U9645 (N_9645,N_9532,N_9510);
nand U9646 (N_9646,N_9531,N_9525);
nand U9647 (N_9647,N_9509,N_9565);
and U9648 (N_9648,N_9502,N_9501);
or U9649 (N_9649,N_9539,N_9522);
nand U9650 (N_9650,N_9524,N_9541);
nor U9651 (N_9651,N_9516,N_9545);
and U9652 (N_9652,N_9575,N_9517);
nand U9653 (N_9653,N_9579,N_9594);
xor U9654 (N_9654,N_9578,N_9538);
and U9655 (N_9655,N_9540,N_9532);
nor U9656 (N_9656,N_9516,N_9544);
nor U9657 (N_9657,N_9551,N_9589);
and U9658 (N_9658,N_9557,N_9595);
nor U9659 (N_9659,N_9575,N_9528);
and U9660 (N_9660,N_9589,N_9549);
nor U9661 (N_9661,N_9572,N_9504);
or U9662 (N_9662,N_9562,N_9574);
or U9663 (N_9663,N_9585,N_9510);
and U9664 (N_9664,N_9517,N_9507);
nor U9665 (N_9665,N_9505,N_9525);
or U9666 (N_9666,N_9585,N_9575);
and U9667 (N_9667,N_9542,N_9513);
nand U9668 (N_9668,N_9548,N_9515);
nor U9669 (N_9669,N_9533,N_9508);
nand U9670 (N_9670,N_9594,N_9552);
or U9671 (N_9671,N_9592,N_9524);
and U9672 (N_9672,N_9565,N_9582);
and U9673 (N_9673,N_9500,N_9544);
or U9674 (N_9674,N_9528,N_9591);
and U9675 (N_9675,N_9598,N_9527);
and U9676 (N_9676,N_9576,N_9570);
or U9677 (N_9677,N_9534,N_9546);
nand U9678 (N_9678,N_9506,N_9591);
and U9679 (N_9679,N_9547,N_9533);
and U9680 (N_9680,N_9578,N_9572);
or U9681 (N_9681,N_9581,N_9533);
xnor U9682 (N_9682,N_9539,N_9541);
and U9683 (N_9683,N_9509,N_9553);
nor U9684 (N_9684,N_9527,N_9549);
nor U9685 (N_9685,N_9569,N_9500);
and U9686 (N_9686,N_9534,N_9533);
nand U9687 (N_9687,N_9510,N_9583);
or U9688 (N_9688,N_9548,N_9514);
or U9689 (N_9689,N_9512,N_9572);
or U9690 (N_9690,N_9571,N_9517);
nand U9691 (N_9691,N_9578,N_9599);
or U9692 (N_9692,N_9542,N_9571);
and U9693 (N_9693,N_9570,N_9561);
nor U9694 (N_9694,N_9510,N_9542);
and U9695 (N_9695,N_9556,N_9590);
and U9696 (N_9696,N_9516,N_9527);
and U9697 (N_9697,N_9585,N_9541);
nor U9698 (N_9698,N_9501,N_9526);
and U9699 (N_9699,N_9576,N_9589);
nand U9700 (N_9700,N_9659,N_9621);
nor U9701 (N_9701,N_9687,N_9605);
or U9702 (N_9702,N_9661,N_9693);
and U9703 (N_9703,N_9674,N_9651);
nor U9704 (N_9704,N_9609,N_9640);
nand U9705 (N_9705,N_9678,N_9649);
nor U9706 (N_9706,N_9614,N_9671);
or U9707 (N_9707,N_9630,N_9601);
and U9708 (N_9708,N_9684,N_9648);
or U9709 (N_9709,N_9642,N_9673);
or U9710 (N_9710,N_9619,N_9698);
and U9711 (N_9711,N_9663,N_9675);
nand U9712 (N_9712,N_9699,N_9672);
and U9713 (N_9713,N_9688,N_9634);
nand U9714 (N_9714,N_9669,N_9655);
or U9715 (N_9715,N_9626,N_9611);
nor U9716 (N_9716,N_9652,N_9633);
xnor U9717 (N_9717,N_9682,N_9676);
nor U9718 (N_9718,N_9691,N_9620);
nand U9719 (N_9719,N_9666,N_9679);
nand U9720 (N_9720,N_9606,N_9697);
nand U9721 (N_9721,N_9692,N_9604);
and U9722 (N_9722,N_9664,N_9646);
or U9723 (N_9723,N_9623,N_9656);
xor U9724 (N_9724,N_9685,N_9628);
and U9725 (N_9725,N_9647,N_9668);
nor U9726 (N_9726,N_9635,N_9681);
nor U9727 (N_9727,N_9662,N_9677);
or U9728 (N_9728,N_9667,N_9641);
and U9729 (N_9729,N_9644,N_9638);
and U9730 (N_9730,N_9643,N_9689);
xor U9731 (N_9731,N_9615,N_9610);
nand U9732 (N_9732,N_9665,N_9658);
or U9733 (N_9733,N_9618,N_9603);
nand U9734 (N_9734,N_9650,N_9612);
nand U9735 (N_9735,N_9627,N_9690);
or U9736 (N_9736,N_9654,N_9680);
nor U9737 (N_9737,N_9629,N_9653);
nand U9738 (N_9738,N_9645,N_9636);
or U9739 (N_9739,N_9608,N_9660);
or U9740 (N_9740,N_9657,N_9602);
nand U9741 (N_9741,N_9617,N_9639);
nor U9742 (N_9742,N_9607,N_9686);
nor U9743 (N_9743,N_9624,N_9696);
xnor U9744 (N_9744,N_9600,N_9694);
nand U9745 (N_9745,N_9637,N_9670);
or U9746 (N_9746,N_9616,N_9683);
or U9747 (N_9747,N_9632,N_9613);
and U9748 (N_9748,N_9695,N_9622);
and U9749 (N_9749,N_9631,N_9625);
nand U9750 (N_9750,N_9672,N_9674);
nand U9751 (N_9751,N_9662,N_9665);
nand U9752 (N_9752,N_9659,N_9624);
and U9753 (N_9753,N_9652,N_9650);
and U9754 (N_9754,N_9601,N_9672);
and U9755 (N_9755,N_9638,N_9696);
nand U9756 (N_9756,N_9657,N_9604);
nand U9757 (N_9757,N_9698,N_9641);
and U9758 (N_9758,N_9654,N_9690);
or U9759 (N_9759,N_9628,N_9639);
nor U9760 (N_9760,N_9665,N_9681);
or U9761 (N_9761,N_9603,N_9654);
and U9762 (N_9762,N_9696,N_9684);
nand U9763 (N_9763,N_9652,N_9685);
xnor U9764 (N_9764,N_9687,N_9682);
and U9765 (N_9765,N_9646,N_9612);
and U9766 (N_9766,N_9635,N_9671);
and U9767 (N_9767,N_9688,N_9629);
nand U9768 (N_9768,N_9647,N_9675);
and U9769 (N_9769,N_9665,N_9634);
and U9770 (N_9770,N_9690,N_9618);
and U9771 (N_9771,N_9673,N_9682);
nor U9772 (N_9772,N_9649,N_9671);
nand U9773 (N_9773,N_9643,N_9695);
and U9774 (N_9774,N_9682,N_9631);
nor U9775 (N_9775,N_9681,N_9631);
and U9776 (N_9776,N_9666,N_9626);
nor U9777 (N_9777,N_9669,N_9639);
or U9778 (N_9778,N_9659,N_9613);
or U9779 (N_9779,N_9600,N_9682);
nor U9780 (N_9780,N_9637,N_9621);
and U9781 (N_9781,N_9664,N_9629);
or U9782 (N_9782,N_9617,N_9638);
nand U9783 (N_9783,N_9600,N_9631);
nand U9784 (N_9784,N_9656,N_9699);
nor U9785 (N_9785,N_9611,N_9660);
nand U9786 (N_9786,N_9637,N_9684);
nor U9787 (N_9787,N_9607,N_9694);
nand U9788 (N_9788,N_9660,N_9668);
and U9789 (N_9789,N_9673,N_9609);
nor U9790 (N_9790,N_9618,N_9614);
nand U9791 (N_9791,N_9621,N_9656);
or U9792 (N_9792,N_9680,N_9678);
xor U9793 (N_9793,N_9698,N_9650);
nor U9794 (N_9794,N_9671,N_9645);
or U9795 (N_9795,N_9631,N_9692);
nor U9796 (N_9796,N_9642,N_9685);
or U9797 (N_9797,N_9603,N_9652);
and U9798 (N_9798,N_9633,N_9639);
and U9799 (N_9799,N_9673,N_9643);
and U9800 (N_9800,N_9779,N_9720);
and U9801 (N_9801,N_9746,N_9769);
nor U9802 (N_9802,N_9767,N_9776);
nor U9803 (N_9803,N_9717,N_9713);
or U9804 (N_9804,N_9701,N_9735);
nand U9805 (N_9805,N_9722,N_9754);
nor U9806 (N_9806,N_9721,N_9723);
nor U9807 (N_9807,N_9773,N_9743);
or U9808 (N_9808,N_9711,N_9732);
nor U9809 (N_9809,N_9738,N_9733);
and U9810 (N_9810,N_9751,N_9762);
nand U9811 (N_9811,N_9799,N_9755);
and U9812 (N_9812,N_9729,N_9787);
nor U9813 (N_9813,N_9750,N_9777);
nor U9814 (N_9814,N_9763,N_9758);
xor U9815 (N_9815,N_9781,N_9736);
nand U9816 (N_9816,N_9794,N_9700);
nor U9817 (N_9817,N_9745,N_9796);
and U9818 (N_9818,N_9749,N_9795);
or U9819 (N_9819,N_9719,N_9739);
nand U9820 (N_9820,N_9706,N_9757);
nand U9821 (N_9821,N_9766,N_9791);
nor U9822 (N_9822,N_9759,N_9785);
nand U9823 (N_9823,N_9790,N_9734);
nor U9824 (N_9824,N_9764,N_9712);
or U9825 (N_9825,N_9715,N_9770);
nor U9826 (N_9826,N_9768,N_9782);
nand U9827 (N_9827,N_9772,N_9707);
and U9828 (N_9828,N_9793,N_9748);
or U9829 (N_9829,N_9747,N_9741);
nand U9830 (N_9830,N_9774,N_9783);
or U9831 (N_9831,N_9744,N_9731);
or U9832 (N_9832,N_9752,N_9765);
nor U9833 (N_9833,N_9716,N_9709);
nand U9834 (N_9834,N_9771,N_9740);
or U9835 (N_9835,N_9761,N_9704);
nor U9836 (N_9836,N_9718,N_9784);
nor U9837 (N_9837,N_9725,N_9705);
nor U9838 (N_9838,N_9742,N_9798);
nor U9839 (N_9839,N_9760,N_9780);
and U9840 (N_9840,N_9703,N_9792);
or U9841 (N_9841,N_9724,N_9756);
nand U9842 (N_9842,N_9788,N_9778);
nor U9843 (N_9843,N_9797,N_9714);
or U9844 (N_9844,N_9737,N_9702);
and U9845 (N_9845,N_9730,N_9789);
nand U9846 (N_9846,N_9708,N_9753);
nor U9847 (N_9847,N_9710,N_9727);
nand U9848 (N_9848,N_9786,N_9728);
or U9849 (N_9849,N_9775,N_9726);
nor U9850 (N_9850,N_9785,N_9732);
nand U9851 (N_9851,N_9755,N_9766);
or U9852 (N_9852,N_9793,N_9780);
or U9853 (N_9853,N_9703,N_9787);
nor U9854 (N_9854,N_9717,N_9766);
or U9855 (N_9855,N_9784,N_9748);
nand U9856 (N_9856,N_9793,N_9713);
and U9857 (N_9857,N_9786,N_9712);
nand U9858 (N_9858,N_9703,N_9764);
or U9859 (N_9859,N_9769,N_9739);
or U9860 (N_9860,N_9754,N_9743);
nand U9861 (N_9861,N_9705,N_9741);
nor U9862 (N_9862,N_9795,N_9777);
nand U9863 (N_9863,N_9729,N_9763);
and U9864 (N_9864,N_9775,N_9741);
or U9865 (N_9865,N_9780,N_9787);
nor U9866 (N_9866,N_9789,N_9780);
and U9867 (N_9867,N_9789,N_9791);
nand U9868 (N_9868,N_9765,N_9758);
nand U9869 (N_9869,N_9734,N_9779);
nand U9870 (N_9870,N_9731,N_9749);
and U9871 (N_9871,N_9708,N_9701);
nor U9872 (N_9872,N_9739,N_9767);
nor U9873 (N_9873,N_9748,N_9714);
nor U9874 (N_9874,N_9704,N_9734);
and U9875 (N_9875,N_9753,N_9772);
nand U9876 (N_9876,N_9776,N_9756);
or U9877 (N_9877,N_9728,N_9788);
nor U9878 (N_9878,N_9715,N_9742);
and U9879 (N_9879,N_9733,N_9741);
and U9880 (N_9880,N_9708,N_9723);
nor U9881 (N_9881,N_9747,N_9748);
or U9882 (N_9882,N_9781,N_9732);
nor U9883 (N_9883,N_9732,N_9747);
or U9884 (N_9884,N_9758,N_9762);
and U9885 (N_9885,N_9751,N_9745);
and U9886 (N_9886,N_9746,N_9794);
and U9887 (N_9887,N_9767,N_9775);
and U9888 (N_9888,N_9731,N_9739);
nor U9889 (N_9889,N_9718,N_9773);
and U9890 (N_9890,N_9757,N_9787);
nor U9891 (N_9891,N_9723,N_9742);
and U9892 (N_9892,N_9701,N_9709);
nor U9893 (N_9893,N_9701,N_9746);
and U9894 (N_9894,N_9716,N_9771);
and U9895 (N_9895,N_9705,N_9782);
nor U9896 (N_9896,N_9731,N_9784);
and U9897 (N_9897,N_9727,N_9774);
nor U9898 (N_9898,N_9772,N_9727);
nor U9899 (N_9899,N_9730,N_9725);
and U9900 (N_9900,N_9871,N_9820);
nor U9901 (N_9901,N_9868,N_9889);
nor U9902 (N_9902,N_9809,N_9838);
or U9903 (N_9903,N_9874,N_9823);
or U9904 (N_9904,N_9898,N_9841);
nand U9905 (N_9905,N_9855,N_9846);
or U9906 (N_9906,N_9859,N_9863);
nand U9907 (N_9907,N_9864,N_9826);
nor U9908 (N_9908,N_9881,N_9870);
nand U9909 (N_9909,N_9814,N_9811);
and U9910 (N_9910,N_9839,N_9892);
nor U9911 (N_9911,N_9876,N_9819);
nand U9912 (N_9912,N_9850,N_9890);
or U9913 (N_9913,N_9843,N_9808);
and U9914 (N_9914,N_9817,N_9840);
and U9915 (N_9915,N_9802,N_9815);
or U9916 (N_9916,N_9877,N_9861);
or U9917 (N_9917,N_9872,N_9879);
and U9918 (N_9918,N_9832,N_9806);
nand U9919 (N_9919,N_9807,N_9849);
nand U9920 (N_9920,N_9828,N_9842);
or U9921 (N_9921,N_9836,N_9845);
and U9922 (N_9922,N_9812,N_9804);
nand U9923 (N_9923,N_9867,N_9880);
nor U9924 (N_9924,N_9818,N_9800);
and U9925 (N_9925,N_9831,N_9873);
nor U9926 (N_9926,N_9894,N_9805);
or U9927 (N_9927,N_9899,N_9816);
nor U9928 (N_9928,N_9810,N_9875);
and U9929 (N_9929,N_9886,N_9852);
or U9930 (N_9930,N_9869,N_9822);
and U9931 (N_9931,N_9866,N_9865);
and U9932 (N_9932,N_9882,N_9895);
or U9933 (N_9933,N_9885,N_9837);
or U9934 (N_9934,N_9801,N_9835);
or U9935 (N_9935,N_9813,N_9860);
or U9936 (N_9936,N_9858,N_9856);
and U9937 (N_9937,N_9853,N_9829);
and U9938 (N_9938,N_9833,N_9884);
or U9939 (N_9939,N_9887,N_9803);
nor U9940 (N_9940,N_9825,N_9888);
nand U9941 (N_9941,N_9848,N_9862);
nand U9942 (N_9942,N_9883,N_9827);
nor U9943 (N_9943,N_9844,N_9893);
and U9944 (N_9944,N_9896,N_9857);
nand U9945 (N_9945,N_9824,N_9821);
nor U9946 (N_9946,N_9830,N_9897);
and U9947 (N_9947,N_9854,N_9834);
nor U9948 (N_9948,N_9847,N_9851);
and U9949 (N_9949,N_9878,N_9891);
and U9950 (N_9950,N_9812,N_9845);
nor U9951 (N_9951,N_9801,N_9857);
or U9952 (N_9952,N_9873,N_9839);
nor U9953 (N_9953,N_9888,N_9814);
nand U9954 (N_9954,N_9837,N_9883);
nand U9955 (N_9955,N_9857,N_9800);
nor U9956 (N_9956,N_9861,N_9883);
and U9957 (N_9957,N_9836,N_9806);
and U9958 (N_9958,N_9830,N_9887);
nand U9959 (N_9959,N_9811,N_9855);
or U9960 (N_9960,N_9895,N_9860);
nor U9961 (N_9961,N_9842,N_9899);
or U9962 (N_9962,N_9857,N_9855);
and U9963 (N_9963,N_9886,N_9893);
and U9964 (N_9964,N_9805,N_9895);
nor U9965 (N_9965,N_9841,N_9884);
nor U9966 (N_9966,N_9898,N_9821);
nor U9967 (N_9967,N_9878,N_9864);
and U9968 (N_9968,N_9852,N_9872);
xor U9969 (N_9969,N_9832,N_9825);
or U9970 (N_9970,N_9868,N_9815);
or U9971 (N_9971,N_9886,N_9884);
nand U9972 (N_9972,N_9897,N_9816);
and U9973 (N_9973,N_9862,N_9830);
nor U9974 (N_9974,N_9866,N_9883);
and U9975 (N_9975,N_9887,N_9834);
or U9976 (N_9976,N_9842,N_9814);
nor U9977 (N_9977,N_9836,N_9871);
nor U9978 (N_9978,N_9832,N_9856);
and U9979 (N_9979,N_9822,N_9877);
nand U9980 (N_9980,N_9802,N_9801);
nor U9981 (N_9981,N_9844,N_9859);
nand U9982 (N_9982,N_9890,N_9809);
or U9983 (N_9983,N_9864,N_9883);
nor U9984 (N_9984,N_9876,N_9829);
nand U9985 (N_9985,N_9899,N_9838);
or U9986 (N_9986,N_9807,N_9873);
and U9987 (N_9987,N_9860,N_9890);
nor U9988 (N_9988,N_9840,N_9899);
and U9989 (N_9989,N_9802,N_9851);
nand U9990 (N_9990,N_9813,N_9887);
or U9991 (N_9991,N_9856,N_9881);
nand U9992 (N_9992,N_9869,N_9820);
and U9993 (N_9993,N_9801,N_9859);
nor U9994 (N_9994,N_9874,N_9897);
nor U9995 (N_9995,N_9832,N_9861);
and U9996 (N_9996,N_9847,N_9829);
nand U9997 (N_9997,N_9848,N_9869);
and U9998 (N_9998,N_9820,N_9882);
and U9999 (N_9999,N_9881,N_9822);
or UO_0 (O_0,N_9963,N_9930);
or UO_1 (O_1,N_9960,N_9915);
nand UO_2 (O_2,N_9909,N_9958);
nand UO_3 (O_3,N_9953,N_9990);
nor UO_4 (O_4,N_9956,N_9902);
nor UO_5 (O_5,N_9946,N_9987);
nand UO_6 (O_6,N_9967,N_9905);
and UO_7 (O_7,N_9941,N_9959);
or UO_8 (O_8,N_9901,N_9932);
nor UO_9 (O_9,N_9926,N_9961);
nor UO_10 (O_10,N_9934,N_9995);
or UO_11 (O_11,N_9970,N_9923);
or UO_12 (O_12,N_9936,N_9993);
nor UO_13 (O_13,N_9954,N_9984);
nor UO_14 (O_14,N_9935,N_9997);
and UO_15 (O_15,N_9974,N_9989);
or UO_16 (O_16,N_9910,N_9999);
nor UO_17 (O_17,N_9957,N_9916);
nand UO_18 (O_18,N_9913,N_9933);
nor UO_19 (O_19,N_9918,N_9942);
and UO_20 (O_20,N_9951,N_9948);
xor UO_21 (O_21,N_9996,N_9912);
xnor UO_22 (O_22,N_9925,N_9991);
nand UO_23 (O_23,N_9929,N_9920);
nand UO_24 (O_24,N_9911,N_9928);
nand UO_25 (O_25,N_9971,N_9917);
or UO_26 (O_26,N_9903,N_9973);
and UO_27 (O_27,N_9994,N_9919);
or UO_28 (O_28,N_9975,N_9980);
nor UO_29 (O_29,N_9906,N_9921);
and UO_30 (O_30,N_9983,N_9907);
or UO_31 (O_31,N_9943,N_9950);
nand UO_32 (O_32,N_9978,N_9955);
nand UO_33 (O_33,N_9972,N_9947);
or UO_34 (O_34,N_9939,N_9968);
and UO_35 (O_35,N_9908,N_9986);
nand UO_36 (O_36,N_9940,N_9979);
nor UO_37 (O_37,N_9900,N_9922);
nand UO_38 (O_38,N_9965,N_9969);
nand UO_39 (O_39,N_9985,N_9931);
nor UO_40 (O_40,N_9976,N_9952);
nor UO_41 (O_41,N_9914,N_9962);
nand UO_42 (O_42,N_9964,N_9981);
nor UO_43 (O_43,N_9924,N_9992);
nor UO_44 (O_44,N_9949,N_9982);
xor UO_45 (O_45,N_9927,N_9977);
nand UO_46 (O_46,N_9938,N_9945);
or UO_47 (O_47,N_9998,N_9944);
or UO_48 (O_48,N_9904,N_9988);
and UO_49 (O_49,N_9966,N_9937);
nand UO_50 (O_50,N_9996,N_9919);
or UO_51 (O_51,N_9931,N_9997);
nor UO_52 (O_52,N_9938,N_9920);
nor UO_53 (O_53,N_9982,N_9927);
xor UO_54 (O_54,N_9959,N_9994);
and UO_55 (O_55,N_9950,N_9998);
nor UO_56 (O_56,N_9997,N_9995);
and UO_57 (O_57,N_9901,N_9941);
and UO_58 (O_58,N_9952,N_9919);
xor UO_59 (O_59,N_9912,N_9946);
and UO_60 (O_60,N_9987,N_9943);
nand UO_61 (O_61,N_9930,N_9999);
nand UO_62 (O_62,N_9908,N_9935);
or UO_63 (O_63,N_9942,N_9955);
or UO_64 (O_64,N_9918,N_9929);
nand UO_65 (O_65,N_9959,N_9914);
and UO_66 (O_66,N_9992,N_9980);
or UO_67 (O_67,N_9988,N_9971);
nand UO_68 (O_68,N_9967,N_9941);
nor UO_69 (O_69,N_9976,N_9956);
nor UO_70 (O_70,N_9940,N_9969);
nor UO_71 (O_71,N_9965,N_9982);
nor UO_72 (O_72,N_9925,N_9953);
nand UO_73 (O_73,N_9928,N_9939);
nand UO_74 (O_74,N_9920,N_9975);
or UO_75 (O_75,N_9926,N_9920);
and UO_76 (O_76,N_9905,N_9985);
nand UO_77 (O_77,N_9993,N_9986);
nand UO_78 (O_78,N_9921,N_9919);
and UO_79 (O_79,N_9947,N_9936);
or UO_80 (O_80,N_9956,N_9931);
and UO_81 (O_81,N_9919,N_9986);
nor UO_82 (O_82,N_9960,N_9916);
nand UO_83 (O_83,N_9903,N_9927);
nor UO_84 (O_84,N_9929,N_9982);
and UO_85 (O_85,N_9976,N_9908);
or UO_86 (O_86,N_9926,N_9924);
and UO_87 (O_87,N_9994,N_9939);
nor UO_88 (O_88,N_9929,N_9914);
nor UO_89 (O_89,N_9988,N_9975);
or UO_90 (O_90,N_9967,N_9955);
and UO_91 (O_91,N_9952,N_9914);
and UO_92 (O_92,N_9940,N_9932);
and UO_93 (O_93,N_9962,N_9980);
or UO_94 (O_94,N_9945,N_9954);
xnor UO_95 (O_95,N_9991,N_9932);
and UO_96 (O_96,N_9983,N_9972);
or UO_97 (O_97,N_9970,N_9920);
nand UO_98 (O_98,N_9952,N_9986);
and UO_99 (O_99,N_9994,N_9968);
nor UO_100 (O_100,N_9942,N_9984);
nor UO_101 (O_101,N_9964,N_9932);
nand UO_102 (O_102,N_9959,N_9979);
nor UO_103 (O_103,N_9930,N_9982);
and UO_104 (O_104,N_9939,N_9904);
or UO_105 (O_105,N_9915,N_9901);
and UO_106 (O_106,N_9995,N_9974);
and UO_107 (O_107,N_9918,N_9936);
and UO_108 (O_108,N_9946,N_9921);
and UO_109 (O_109,N_9949,N_9956);
or UO_110 (O_110,N_9908,N_9990);
nand UO_111 (O_111,N_9923,N_9936);
nor UO_112 (O_112,N_9981,N_9968);
and UO_113 (O_113,N_9924,N_9935);
and UO_114 (O_114,N_9986,N_9944);
nor UO_115 (O_115,N_9997,N_9919);
nand UO_116 (O_116,N_9945,N_9950);
or UO_117 (O_117,N_9919,N_9933);
nor UO_118 (O_118,N_9969,N_9951);
nor UO_119 (O_119,N_9960,N_9963);
and UO_120 (O_120,N_9977,N_9937);
and UO_121 (O_121,N_9982,N_9912);
nor UO_122 (O_122,N_9992,N_9957);
nor UO_123 (O_123,N_9976,N_9995);
or UO_124 (O_124,N_9989,N_9939);
and UO_125 (O_125,N_9921,N_9962);
or UO_126 (O_126,N_9941,N_9993);
and UO_127 (O_127,N_9934,N_9955);
nand UO_128 (O_128,N_9987,N_9994);
nand UO_129 (O_129,N_9955,N_9997);
nand UO_130 (O_130,N_9962,N_9955);
or UO_131 (O_131,N_9962,N_9900);
nand UO_132 (O_132,N_9927,N_9922);
nand UO_133 (O_133,N_9961,N_9948);
or UO_134 (O_134,N_9974,N_9976);
or UO_135 (O_135,N_9946,N_9936);
nand UO_136 (O_136,N_9963,N_9990);
nor UO_137 (O_137,N_9914,N_9966);
nand UO_138 (O_138,N_9996,N_9949);
xnor UO_139 (O_139,N_9985,N_9953);
and UO_140 (O_140,N_9987,N_9904);
xor UO_141 (O_141,N_9992,N_9996);
nor UO_142 (O_142,N_9925,N_9926);
and UO_143 (O_143,N_9956,N_9986);
or UO_144 (O_144,N_9994,N_9989);
nand UO_145 (O_145,N_9977,N_9904);
xor UO_146 (O_146,N_9951,N_9925);
and UO_147 (O_147,N_9927,N_9962);
nand UO_148 (O_148,N_9972,N_9933);
and UO_149 (O_149,N_9977,N_9988);
and UO_150 (O_150,N_9994,N_9990);
nand UO_151 (O_151,N_9943,N_9908);
and UO_152 (O_152,N_9971,N_9987);
nand UO_153 (O_153,N_9966,N_9985);
or UO_154 (O_154,N_9962,N_9984);
or UO_155 (O_155,N_9903,N_9991);
nor UO_156 (O_156,N_9906,N_9931);
nand UO_157 (O_157,N_9918,N_9952);
and UO_158 (O_158,N_9914,N_9981);
or UO_159 (O_159,N_9935,N_9919);
nand UO_160 (O_160,N_9955,N_9904);
nand UO_161 (O_161,N_9931,N_9975);
nand UO_162 (O_162,N_9917,N_9981);
or UO_163 (O_163,N_9924,N_9995);
and UO_164 (O_164,N_9990,N_9980);
xnor UO_165 (O_165,N_9952,N_9926);
and UO_166 (O_166,N_9914,N_9969);
nand UO_167 (O_167,N_9907,N_9926);
or UO_168 (O_168,N_9914,N_9970);
and UO_169 (O_169,N_9922,N_9957);
and UO_170 (O_170,N_9928,N_9929);
nand UO_171 (O_171,N_9916,N_9920);
and UO_172 (O_172,N_9959,N_9968);
and UO_173 (O_173,N_9998,N_9993);
or UO_174 (O_174,N_9907,N_9911);
nor UO_175 (O_175,N_9935,N_9907);
nor UO_176 (O_176,N_9990,N_9937);
or UO_177 (O_177,N_9960,N_9956);
and UO_178 (O_178,N_9956,N_9989);
nor UO_179 (O_179,N_9904,N_9954);
nor UO_180 (O_180,N_9943,N_9977);
or UO_181 (O_181,N_9997,N_9913);
nand UO_182 (O_182,N_9945,N_9946);
nand UO_183 (O_183,N_9980,N_9974);
and UO_184 (O_184,N_9944,N_9997);
and UO_185 (O_185,N_9989,N_9914);
nand UO_186 (O_186,N_9926,N_9998);
nor UO_187 (O_187,N_9908,N_9945);
nor UO_188 (O_188,N_9928,N_9925);
and UO_189 (O_189,N_9930,N_9933);
nand UO_190 (O_190,N_9984,N_9932);
and UO_191 (O_191,N_9963,N_9996);
or UO_192 (O_192,N_9902,N_9944);
nand UO_193 (O_193,N_9908,N_9956);
or UO_194 (O_194,N_9935,N_9939);
and UO_195 (O_195,N_9962,N_9906);
nor UO_196 (O_196,N_9949,N_9943);
nand UO_197 (O_197,N_9918,N_9950);
and UO_198 (O_198,N_9929,N_9910);
nand UO_199 (O_199,N_9913,N_9990);
nand UO_200 (O_200,N_9956,N_9903);
and UO_201 (O_201,N_9932,N_9954);
and UO_202 (O_202,N_9980,N_9987);
nor UO_203 (O_203,N_9982,N_9924);
and UO_204 (O_204,N_9964,N_9913);
nor UO_205 (O_205,N_9917,N_9961);
nand UO_206 (O_206,N_9936,N_9987);
nand UO_207 (O_207,N_9977,N_9901);
nand UO_208 (O_208,N_9958,N_9965);
nand UO_209 (O_209,N_9906,N_9974);
or UO_210 (O_210,N_9971,N_9999);
nor UO_211 (O_211,N_9979,N_9904);
nor UO_212 (O_212,N_9963,N_9953);
and UO_213 (O_213,N_9954,N_9918);
and UO_214 (O_214,N_9950,N_9986);
or UO_215 (O_215,N_9930,N_9977);
nand UO_216 (O_216,N_9944,N_9981);
nor UO_217 (O_217,N_9909,N_9997);
and UO_218 (O_218,N_9904,N_9943);
and UO_219 (O_219,N_9901,N_9970);
or UO_220 (O_220,N_9992,N_9935);
or UO_221 (O_221,N_9912,N_9936);
nand UO_222 (O_222,N_9903,N_9965);
and UO_223 (O_223,N_9905,N_9998);
nor UO_224 (O_224,N_9980,N_9909);
or UO_225 (O_225,N_9916,N_9935);
and UO_226 (O_226,N_9963,N_9944);
and UO_227 (O_227,N_9957,N_9988);
or UO_228 (O_228,N_9911,N_9964);
or UO_229 (O_229,N_9989,N_9909);
and UO_230 (O_230,N_9972,N_9936);
or UO_231 (O_231,N_9948,N_9935);
nand UO_232 (O_232,N_9988,N_9911);
nand UO_233 (O_233,N_9991,N_9947);
nand UO_234 (O_234,N_9914,N_9961);
or UO_235 (O_235,N_9940,N_9957);
nor UO_236 (O_236,N_9971,N_9940);
and UO_237 (O_237,N_9975,N_9904);
or UO_238 (O_238,N_9936,N_9970);
nand UO_239 (O_239,N_9949,N_9998);
nor UO_240 (O_240,N_9975,N_9962);
and UO_241 (O_241,N_9993,N_9924);
nand UO_242 (O_242,N_9937,N_9971);
nor UO_243 (O_243,N_9993,N_9954);
nor UO_244 (O_244,N_9949,N_9924);
nor UO_245 (O_245,N_9936,N_9950);
and UO_246 (O_246,N_9956,N_9963);
or UO_247 (O_247,N_9914,N_9947);
or UO_248 (O_248,N_9945,N_9926);
and UO_249 (O_249,N_9977,N_9934);
nor UO_250 (O_250,N_9982,N_9914);
or UO_251 (O_251,N_9918,N_9976);
and UO_252 (O_252,N_9917,N_9944);
nand UO_253 (O_253,N_9986,N_9997);
nand UO_254 (O_254,N_9992,N_9911);
nand UO_255 (O_255,N_9942,N_9986);
or UO_256 (O_256,N_9966,N_9943);
nand UO_257 (O_257,N_9977,N_9918);
or UO_258 (O_258,N_9982,N_9953);
nand UO_259 (O_259,N_9960,N_9955);
nor UO_260 (O_260,N_9973,N_9989);
nand UO_261 (O_261,N_9940,N_9959);
nand UO_262 (O_262,N_9911,N_9982);
nor UO_263 (O_263,N_9921,N_9977);
nor UO_264 (O_264,N_9919,N_9957);
xnor UO_265 (O_265,N_9982,N_9985);
or UO_266 (O_266,N_9967,N_9909);
or UO_267 (O_267,N_9952,N_9971);
and UO_268 (O_268,N_9915,N_9955);
nor UO_269 (O_269,N_9957,N_9904);
xnor UO_270 (O_270,N_9975,N_9945);
nand UO_271 (O_271,N_9981,N_9961);
nand UO_272 (O_272,N_9905,N_9930);
and UO_273 (O_273,N_9999,N_9962);
and UO_274 (O_274,N_9913,N_9908);
nor UO_275 (O_275,N_9994,N_9943);
and UO_276 (O_276,N_9906,N_9960);
or UO_277 (O_277,N_9921,N_9918);
and UO_278 (O_278,N_9980,N_9994);
and UO_279 (O_279,N_9975,N_9916);
and UO_280 (O_280,N_9959,N_9986);
or UO_281 (O_281,N_9955,N_9988);
and UO_282 (O_282,N_9959,N_9935);
or UO_283 (O_283,N_9924,N_9980);
or UO_284 (O_284,N_9917,N_9966);
and UO_285 (O_285,N_9924,N_9936);
nand UO_286 (O_286,N_9912,N_9976);
or UO_287 (O_287,N_9908,N_9949);
or UO_288 (O_288,N_9934,N_9956);
or UO_289 (O_289,N_9941,N_9955);
and UO_290 (O_290,N_9947,N_9978);
nor UO_291 (O_291,N_9906,N_9964);
or UO_292 (O_292,N_9933,N_9922);
nand UO_293 (O_293,N_9921,N_9975);
nor UO_294 (O_294,N_9953,N_9914);
xnor UO_295 (O_295,N_9976,N_9937);
nor UO_296 (O_296,N_9965,N_9957);
and UO_297 (O_297,N_9955,N_9900);
nor UO_298 (O_298,N_9909,N_9940);
and UO_299 (O_299,N_9977,N_9999);
or UO_300 (O_300,N_9923,N_9945);
nor UO_301 (O_301,N_9993,N_9930);
and UO_302 (O_302,N_9999,N_9950);
nand UO_303 (O_303,N_9921,N_9955);
nor UO_304 (O_304,N_9971,N_9908);
nand UO_305 (O_305,N_9964,N_9958);
or UO_306 (O_306,N_9952,N_9945);
nor UO_307 (O_307,N_9984,N_9972);
nand UO_308 (O_308,N_9907,N_9970);
nand UO_309 (O_309,N_9934,N_9965);
nor UO_310 (O_310,N_9990,N_9902);
nor UO_311 (O_311,N_9912,N_9924);
or UO_312 (O_312,N_9998,N_9907);
xor UO_313 (O_313,N_9933,N_9909);
nor UO_314 (O_314,N_9973,N_9953);
and UO_315 (O_315,N_9998,N_9996);
xor UO_316 (O_316,N_9930,N_9954);
nand UO_317 (O_317,N_9953,N_9927);
and UO_318 (O_318,N_9951,N_9934);
xor UO_319 (O_319,N_9984,N_9944);
nand UO_320 (O_320,N_9957,N_9911);
nor UO_321 (O_321,N_9988,N_9908);
and UO_322 (O_322,N_9947,N_9950);
and UO_323 (O_323,N_9966,N_9934);
nor UO_324 (O_324,N_9991,N_9909);
nor UO_325 (O_325,N_9972,N_9944);
and UO_326 (O_326,N_9990,N_9946);
nor UO_327 (O_327,N_9985,N_9904);
or UO_328 (O_328,N_9935,N_9928);
nor UO_329 (O_329,N_9908,N_9992);
and UO_330 (O_330,N_9991,N_9963);
nor UO_331 (O_331,N_9960,N_9980);
nor UO_332 (O_332,N_9949,N_9987);
or UO_333 (O_333,N_9915,N_9996);
or UO_334 (O_334,N_9957,N_9945);
and UO_335 (O_335,N_9983,N_9902);
nor UO_336 (O_336,N_9954,N_9959);
xnor UO_337 (O_337,N_9997,N_9992);
nand UO_338 (O_338,N_9992,N_9960);
nand UO_339 (O_339,N_9907,N_9993);
nor UO_340 (O_340,N_9977,N_9978);
or UO_341 (O_341,N_9967,N_9944);
or UO_342 (O_342,N_9934,N_9940);
or UO_343 (O_343,N_9912,N_9979);
and UO_344 (O_344,N_9914,N_9964);
xor UO_345 (O_345,N_9937,N_9968);
and UO_346 (O_346,N_9992,N_9918);
nor UO_347 (O_347,N_9908,N_9969);
nor UO_348 (O_348,N_9916,N_9906);
nand UO_349 (O_349,N_9924,N_9966);
nor UO_350 (O_350,N_9945,N_9998);
or UO_351 (O_351,N_9955,N_9998);
xor UO_352 (O_352,N_9915,N_9971);
and UO_353 (O_353,N_9928,N_9941);
nor UO_354 (O_354,N_9925,N_9992);
nand UO_355 (O_355,N_9951,N_9961);
nand UO_356 (O_356,N_9915,N_9974);
xnor UO_357 (O_357,N_9944,N_9966);
nor UO_358 (O_358,N_9901,N_9938);
nor UO_359 (O_359,N_9902,N_9947);
nand UO_360 (O_360,N_9906,N_9943);
nand UO_361 (O_361,N_9989,N_9969);
and UO_362 (O_362,N_9928,N_9981);
nor UO_363 (O_363,N_9943,N_9972);
or UO_364 (O_364,N_9927,N_9914);
nor UO_365 (O_365,N_9919,N_9906);
nor UO_366 (O_366,N_9942,N_9909);
nand UO_367 (O_367,N_9949,N_9930);
nor UO_368 (O_368,N_9910,N_9981);
nor UO_369 (O_369,N_9959,N_9900);
or UO_370 (O_370,N_9940,N_9960);
xor UO_371 (O_371,N_9907,N_9999);
nor UO_372 (O_372,N_9928,N_9900);
and UO_373 (O_373,N_9958,N_9902);
nand UO_374 (O_374,N_9904,N_9964);
nand UO_375 (O_375,N_9926,N_9955);
and UO_376 (O_376,N_9942,N_9945);
or UO_377 (O_377,N_9959,N_9908);
and UO_378 (O_378,N_9933,N_9996);
nand UO_379 (O_379,N_9964,N_9945);
nand UO_380 (O_380,N_9921,N_9964);
or UO_381 (O_381,N_9934,N_9919);
nor UO_382 (O_382,N_9997,N_9918);
or UO_383 (O_383,N_9928,N_9947);
or UO_384 (O_384,N_9990,N_9976);
xnor UO_385 (O_385,N_9933,N_9916);
and UO_386 (O_386,N_9929,N_9990);
nor UO_387 (O_387,N_9903,N_9937);
nand UO_388 (O_388,N_9945,N_9902);
or UO_389 (O_389,N_9963,N_9903);
and UO_390 (O_390,N_9967,N_9911);
and UO_391 (O_391,N_9910,N_9987);
nand UO_392 (O_392,N_9987,N_9970);
and UO_393 (O_393,N_9995,N_9905);
nand UO_394 (O_394,N_9938,N_9979);
nand UO_395 (O_395,N_9985,N_9933);
xnor UO_396 (O_396,N_9989,N_9988);
and UO_397 (O_397,N_9901,N_9980);
or UO_398 (O_398,N_9955,N_9950);
or UO_399 (O_399,N_9918,N_9998);
nand UO_400 (O_400,N_9919,N_9961);
and UO_401 (O_401,N_9929,N_9931);
and UO_402 (O_402,N_9980,N_9907);
and UO_403 (O_403,N_9980,N_9922);
nand UO_404 (O_404,N_9906,N_9985);
or UO_405 (O_405,N_9977,N_9900);
nand UO_406 (O_406,N_9942,N_9967);
and UO_407 (O_407,N_9974,N_9997);
nand UO_408 (O_408,N_9935,N_9933);
nor UO_409 (O_409,N_9931,N_9903);
nor UO_410 (O_410,N_9916,N_9972);
and UO_411 (O_411,N_9915,N_9958);
and UO_412 (O_412,N_9973,N_9960);
or UO_413 (O_413,N_9973,N_9993);
nor UO_414 (O_414,N_9963,N_9919);
or UO_415 (O_415,N_9941,N_9990);
nor UO_416 (O_416,N_9969,N_9939);
or UO_417 (O_417,N_9905,N_9945);
nand UO_418 (O_418,N_9911,N_9981);
or UO_419 (O_419,N_9986,N_9923);
and UO_420 (O_420,N_9934,N_9946);
or UO_421 (O_421,N_9953,N_9918);
and UO_422 (O_422,N_9903,N_9953);
nor UO_423 (O_423,N_9962,N_9982);
xnor UO_424 (O_424,N_9921,N_9983);
nor UO_425 (O_425,N_9958,N_9926);
nand UO_426 (O_426,N_9982,N_9900);
or UO_427 (O_427,N_9926,N_9904);
and UO_428 (O_428,N_9917,N_9945);
nor UO_429 (O_429,N_9952,N_9934);
nand UO_430 (O_430,N_9967,N_9925);
or UO_431 (O_431,N_9930,N_9921);
nand UO_432 (O_432,N_9906,N_9928);
or UO_433 (O_433,N_9966,N_9946);
nor UO_434 (O_434,N_9964,N_9915);
or UO_435 (O_435,N_9995,N_9972);
nor UO_436 (O_436,N_9986,N_9985);
nand UO_437 (O_437,N_9900,N_9997);
nor UO_438 (O_438,N_9958,N_9942);
nand UO_439 (O_439,N_9974,N_9959);
nand UO_440 (O_440,N_9916,N_9977);
and UO_441 (O_441,N_9914,N_9991);
or UO_442 (O_442,N_9983,N_9989);
nor UO_443 (O_443,N_9911,N_9925);
or UO_444 (O_444,N_9986,N_9939);
nor UO_445 (O_445,N_9952,N_9994);
nor UO_446 (O_446,N_9924,N_9909);
or UO_447 (O_447,N_9947,N_9923);
or UO_448 (O_448,N_9959,N_9963);
and UO_449 (O_449,N_9935,N_9977);
and UO_450 (O_450,N_9999,N_9946);
nand UO_451 (O_451,N_9932,N_9931);
or UO_452 (O_452,N_9975,N_9908);
nor UO_453 (O_453,N_9952,N_9911);
nor UO_454 (O_454,N_9927,N_9915);
nand UO_455 (O_455,N_9920,N_9951);
nor UO_456 (O_456,N_9950,N_9907);
and UO_457 (O_457,N_9913,N_9931);
and UO_458 (O_458,N_9936,N_9909);
nor UO_459 (O_459,N_9997,N_9938);
and UO_460 (O_460,N_9941,N_9995);
nor UO_461 (O_461,N_9916,N_9999);
and UO_462 (O_462,N_9911,N_9932);
or UO_463 (O_463,N_9925,N_9993);
and UO_464 (O_464,N_9983,N_9966);
or UO_465 (O_465,N_9918,N_9928);
or UO_466 (O_466,N_9959,N_9985);
nor UO_467 (O_467,N_9981,N_9947);
nand UO_468 (O_468,N_9901,N_9995);
and UO_469 (O_469,N_9927,N_9902);
or UO_470 (O_470,N_9930,N_9901);
and UO_471 (O_471,N_9940,N_9946);
nor UO_472 (O_472,N_9933,N_9920);
nor UO_473 (O_473,N_9959,N_9993);
nor UO_474 (O_474,N_9904,N_9958);
nand UO_475 (O_475,N_9965,N_9976);
or UO_476 (O_476,N_9929,N_9915);
or UO_477 (O_477,N_9939,N_9995);
nand UO_478 (O_478,N_9938,N_9910);
or UO_479 (O_479,N_9904,N_9928);
or UO_480 (O_480,N_9934,N_9957);
nand UO_481 (O_481,N_9983,N_9970);
and UO_482 (O_482,N_9903,N_9943);
and UO_483 (O_483,N_9911,N_9945);
nor UO_484 (O_484,N_9953,N_9961);
nor UO_485 (O_485,N_9973,N_9963);
nand UO_486 (O_486,N_9981,N_9905);
and UO_487 (O_487,N_9950,N_9977);
nor UO_488 (O_488,N_9987,N_9976);
or UO_489 (O_489,N_9991,N_9989);
nand UO_490 (O_490,N_9952,N_9915);
or UO_491 (O_491,N_9924,N_9946);
and UO_492 (O_492,N_9919,N_9916);
nand UO_493 (O_493,N_9972,N_9932);
nand UO_494 (O_494,N_9938,N_9908);
nor UO_495 (O_495,N_9975,N_9978);
nand UO_496 (O_496,N_9975,N_9970);
nand UO_497 (O_497,N_9942,N_9976);
and UO_498 (O_498,N_9963,N_9966);
or UO_499 (O_499,N_9956,N_9994);
nand UO_500 (O_500,N_9928,N_9969);
nand UO_501 (O_501,N_9957,N_9973);
nor UO_502 (O_502,N_9939,N_9900);
or UO_503 (O_503,N_9934,N_9915);
nor UO_504 (O_504,N_9902,N_9980);
or UO_505 (O_505,N_9909,N_9910);
nand UO_506 (O_506,N_9959,N_9939);
nor UO_507 (O_507,N_9946,N_9995);
nand UO_508 (O_508,N_9967,N_9983);
and UO_509 (O_509,N_9969,N_9944);
nand UO_510 (O_510,N_9931,N_9983);
nor UO_511 (O_511,N_9962,N_9992);
nor UO_512 (O_512,N_9905,N_9971);
and UO_513 (O_513,N_9955,N_9958);
or UO_514 (O_514,N_9988,N_9960);
and UO_515 (O_515,N_9966,N_9938);
and UO_516 (O_516,N_9998,N_9983);
nand UO_517 (O_517,N_9965,N_9999);
nor UO_518 (O_518,N_9913,N_9996);
or UO_519 (O_519,N_9999,N_9964);
or UO_520 (O_520,N_9930,N_9953);
nor UO_521 (O_521,N_9978,N_9998);
and UO_522 (O_522,N_9985,N_9945);
nor UO_523 (O_523,N_9948,N_9915);
or UO_524 (O_524,N_9967,N_9973);
xor UO_525 (O_525,N_9967,N_9965);
nor UO_526 (O_526,N_9931,N_9974);
and UO_527 (O_527,N_9948,N_9949);
nand UO_528 (O_528,N_9925,N_9932);
and UO_529 (O_529,N_9947,N_9973);
or UO_530 (O_530,N_9932,N_9945);
and UO_531 (O_531,N_9944,N_9935);
or UO_532 (O_532,N_9924,N_9947);
or UO_533 (O_533,N_9971,N_9907);
nor UO_534 (O_534,N_9983,N_9929);
nand UO_535 (O_535,N_9900,N_9905);
nand UO_536 (O_536,N_9950,N_9984);
nor UO_537 (O_537,N_9992,N_9953);
nand UO_538 (O_538,N_9923,N_9979);
nor UO_539 (O_539,N_9920,N_9981);
nor UO_540 (O_540,N_9996,N_9982);
nor UO_541 (O_541,N_9993,N_9970);
or UO_542 (O_542,N_9961,N_9987);
and UO_543 (O_543,N_9928,N_9930);
nand UO_544 (O_544,N_9960,N_9964);
nand UO_545 (O_545,N_9949,N_9936);
nand UO_546 (O_546,N_9900,N_9952);
and UO_547 (O_547,N_9941,N_9906);
and UO_548 (O_548,N_9911,N_9914);
nand UO_549 (O_549,N_9938,N_9955);
nand UO_550 (O_550,N_9998,N_9935);
or UO_551 (O_551,N_9915,N_9963);
nor UO_552 (O_552,N_9957,N_9963);
and UO_553 (O_553,N_9971,N_9973);
or UO_554 (O_554,N_9936,N_9965);
nor UO_555 (O_555,N_9926,N_9919);
and UO_556 (O_556,N_9928,N_9961);
and UO_557 (O_557,N_9910,N_9951);
nand UO_558 (O_558,N_9956,N_9914);
nand UO_559 (O_559,N_9993,N_9995);
nor UO_560 (O_560,N_9911,N_9937);
and UO_561 (O_561,N_9999,N_9903);
and UO_562 (O_562,N_9949,N_9961);
or UO_563 (O_563,N_9900,N_9919);
or UO_564 (O_564,N_9920,N_9974);
and UO_565 (O_565,N_9953,N_9922);
nand UO_566 (O_566,N_9961,N_9970);
and UO_567 (O_567,N_9974,N_9911);
nor UO_568 (O_568,N_9972,N_9928);
or UO_569 (O_569,N_9960,N_9951);
or UO_570 (O_570,N_9933,N_9902);
nand UO_571 (O_571,N_9964,N_9947);
xor UO_572 (O_572,N_9928,N_9974);
or UO_573 (O_573,N_9987,N_9951);
and UO_574 (O_574,N_9995,N_9921);
xor UO_575 (O_575,N_9904,N_9982);
nor UO_576 (O_576,N_9971,N_9929);
or UO_577 (O_577,N_9925,N_9984);
and UO_578 (O_578,N_9918,N_9979);
or UO_579 (O_579,N_9951,N_9973);
or UO_580 (O_580,N_9991,N_9964);
nand UO_581 (O_581,N_9989,N_9903);
nor UO_582 (O_582,N_9996,N_9931);
xnor UO_583 (O_583,N_9991,N_9917);
nor UO_584 (O_584,N_9957,N_9978);
or UO_585 (O_585,N_9992,N_9916);
xor UO_586 (O_586,N_9978,N_9958);
nand UO_587 (O_587,N_9920,N_9989);
nand UO_588 (O_588,N_9960,N_9974);
xnor UO_589 (O_589,N_9958,N_9992);
or UO_590 (O_590,N_9948,N_9911);
nor UO_591 (O_591,N_9928,N_9954);
nor UO_592 (O_592,N_9950,N_9913);
nand UO_593 (O_593,N_9929,N_9939);
or UO_594 (O_594,N_9912,N_9945);
nor UO_595 (O_595,N_9950,N_9971);
nand UO_596 (O_596,N_9936,N_9901);
nand UO_597 (O_597,N_9984,N_9977);
xor UO_598 (O_598,N_9911,N_9975);
and UO_599 (O_599,N_9961,N_9916);
nand UO_600 (O_600,N_9991,N_9922);
nor UO_601 (O_601,N_9970,N_9990);
nand UO_602 (O_602,N_9978,N_9976);
or UO_603 (O_603,N_9911,N_9921);
or UO_604 (O_604,N_9946,N_9969);
nor UO_605 (O_605,N_9984,N_9905);
and UO_606 (O_606,N_9965,N_9983);
or UO_607 (O_607,N_9947,N_9975);
and UO_608 (O_608,N_9962,N_9969);
nor UO_609 (O_609,N_9987,N_9947);
nor UO_610 (O_610,N_9956,N_9965);
or UO_611 (O_611,N_9929,N_9923);
and UO_612 (O_612,N_9979,N_9977);
nand UO_613 (O_613,N_9948,N_9908);
nand UO_614 (O_614,N_9906,N_9914);
nor UO_615 (O_615,N_9958,N_9966);
or UO_616 (O_616,N_9968,N_9920);
nand UO_617 (O_617,N_9973,N_9913);
and UO_618 (O_618,N_9909,N_9999);
nor UO_619 (O_619,N_9943,N_9973);
and UO_620 (O_620,N_9974,N_9996);
nand UO_621 (O_621,N_9960,N_9996);
and UO_622 (O_622,N_9900,N_9995);
nand UO_623 (O_623,N_9913,N_9928);
nand UO_624 (O_624,N_9941,N_9976);
and UO_625 (O_625,N_9943,N_9952);
nand UO_626 (O_626,N_9956,N_9980);
or UO_627 (O_627,N_9958,N_9940);
nand UO_628 (O_628,N_9911,N_9995);
nor UO_629 (O_629,N_9925,N_9980);
and UO_630 (O_630,N_9986,N_9934);
nor UO_631 (O_631,N_9975,N_9917);
nand UO_632 (O_632,N_9984,N_9952);
nand UO_633 (O_633,N_9901,N_9959);
nand UO_634 (O_634,N_9910,N_9989);
and UO_635 (O_635,N_9942,N_9938);
or UO_636 (O_636,N_9948,N_9906);
or UO_637 (O_637,N_9948,N_9904);
or UO_638 (O_638,N_9974,N_9916);
and UO_639 (O_639,N_9943,N_9938);
and UO_640 (O_640,N_9919,N_9984);
nand UO_641 (O_641,N_9933,N_9989);
and UO_642 (O_642,N_9920,N_9904);
nand UO_643 (O_643,N_9923,N_9901);
nor UO_644 (O_644,N_9942,N_9914);
and UO_645 (O_645,N_9924,N_9986);
nor UO_646 (O_646,N_9947,N_9934);
or UO_647 (O_647,N_9919,N_9941);
nand UO_648 (O_648,N_9967,N_9906);
nand UO_649 (O_649,N_9954,N_9927);
nand UO_650 (O_650,N_9902,N_9922);
nand UO_651 (O_651,N_9942,N_9959);
nor UO_652 (O_652,N_9905,N_9987);
or UO_653 (O_653,N_9917,N_9942);
nand UO_654 (O_654,N_9998,N_9900);
and UO_655 (O_655,N_9943,N_9962);
nor UO_656 (O_656,N_9988,N_9982);
nor UO_657 (O_657,N_9972,N_9963);
nor UO_658 (O_658,N_9903,N_9917);
or UO_659 (O_659,N_9914,N_9941);
nor UO_660 (O_660,N_9962,N_9977);
and UO_661 (O_661,N_9991,N_9996);
or UO_662 (O_662,N_9942,N_9975);
or UO_663 (O_663,N_9907,N_9989);
nor UO_664 (O_664,N_9980,N_9965);
xor UO_665 (O_665,N_9975,N_9954);
nand UO_666 (O_666,N_9963,N_9922);
or UO_667 (O_667,N_9901,N_9997);
nor UO_668 (O_668,N_9927,N_9978);
and UO_669 (O_669,N_9991,N_9900);
nor UO_670 (O_670,N_9962,N_9945);
nand UO_671 (O_671,N_9972,N_9985);
or UO_672 (O_672,N_9983,N_9925);
and UO_673 (O_673,N_9923,N_9937);
and UO_674 (O_674,N_9926,N_9997);
nand UO_675 (O_675,N_9997,N_9999);
and UO_676 (O_676,N_9992,N_9921);
and UO_677 (O_677,N_9939,N_9945);
and UO_678 (O_678,N_9956,N_9961);
and UO_679 (O_679,N_9935,N_9987);
or UO_680 (O_680,N_9918,N_9958);
nand UO_681 (O_681,N_9940,N_9995);
nor UO_682 (O_682,N_9948,N_9947);
and UO_683 (O_683,N_9988,N_9965);
nor UO_684 (O_684,N_9901,N_9909);
nor UO_685 (O_685,N_9977,N_9915);
nor UO_686 (O_686,N_9905,N_9978);
xor UO_687 (O_687,N_9917,N_9962);
nor UO_688 (O_688,N_9920,N_9908);
or UO_689 (O_689,N_9909,N_9986);
and UO_690 (O_690,N_9965,N_9927);
and UO_691 (O_691,N_9984,N_9947);
nand UO_692 (O_692,N_9986,N_9918);
or UO_693 (O_693,N_9917,N_9915);
and UO_694 (O_694,N_9928,N_9952);
and UO_695 (O_695,N_9962,N_9908);
nand UO_696 (O_696,N_9912,N_9988);
nor UO_697 (O_697,N_9914,N_9967);
nand UO_698 (O_698,N_9928,N_9965);
nand UO_699 (O_699,N_9984,N_9913);
nand UO_700 (O_700,N_9968,N_9999);
and UO_701 (O_701,N_9971,N_9910);
nand UO_702 (O_702,N_9911,N_9941);
and UO_703 (O_703,N_9937,N_9955);
nand UO_704 (O_704,N_9965,N_9915);
or UO_705 (O_705,N_9998,N_9984);
nand UO_706 (O_706,N_9982,N_9983);
nor UO_707 (O_707,N_9920,N_9941);
nor UO_708 (O_708,N_9945,N_9987);
or UO_709 (O_709,N_9950,N_9974);
and UO_710 (O_710,N_9944,N_9936);
and UO_711 (O_711,N_9947,N_9968);
or UO_712 (O_712,N_9998,N_9931);
or UO_713 (O_713,N_9998,N_9975);
or UO_714 (O_714,N_9955,N_9961);
nand UO_715 (O_715,N_9930,N_9908);
and UO_716 (O_716,N_9979,N_9933);
nand UO_717 (O_717,N_9982,N_9964);
and UO_718 (O_718,N_9901,N_9974);
nand UO_719 (O_719,N_9996,N_9923);
nand UO_720 (O_720,N_9902,N_9929);
nand UO_721 (O_721,N_9971,N_9995);
nor UO_722 (O_722,N_9947,N_9912);
or UO_723 (O_723,N_9991,N_9950);
nand UO_724 (O_724,N_9928,N_9946);
nand UO_725 (O_725,N_9991,N_9977);
or UO_726 (O_726,N_9961,N_9974);
nand UO_727 (O_727,N_9968,N_9990);
nand UO_728 (O_728,N_9930,N_9927);
and UO_729 (O_729,N_9967,N_9991);
and UO_730 (O_730,N_9979,N_9925);
or UO_731 (O_731,N_9911,N_9976);
nor UO_732 (O_732,N_9987,N_9963);
or UO_733 (O_733,N_9996,N_9964);
and UO_734 (O_734,N_9918,N_9911);
or UO_735 (O_735,N_9983,N_9977);
nor UO_736 (O_736,N_9998,N_9929);
nand UO_737 (O_737,N_9906,N_9946);
or UO_738 (O_738,N_9970,N_9957);
nor UO_739 (O_739,N_9964,N_9986);
xor UO_740 (O_740,N_9938,N_9972);
nor UO_741 (O_741,N_9982,N_9998);
xor UO_742 (O_742,N_9957,N_9983);
and UO_743 (O_743,N_9992,N_9995);
or UO_744 (O_744,N_9922,N_9935);
or UO_745 (O_745,N_9914,N_9943);
or UO_746 (O_746,N_9921,N_9910);
nor UO_747 (O_747,N_9980,N_9903);
xor UO_748 (O_748,N_9954,N_9972);
or UO_749 (O_749,N_9959,N_9966);
or UO_750 (O_750,N_9990,N_9921);
nor UO_751 (O_751,N_9913,N_9935);
or UO_752 (O_752,N_9945,N_9934);
or UO_753 (O_753,N_9903,N_9913);
or UO_754 (O_754,N_9923,N_9969);
or UO_755 (O_755,N_9932,N_9934);
nand UO_756 (O_756,N_9983,N_9918);
nor UO_757 (O_757,N_9962,N_9911);
and UO_758 (O_758,N_9918,N_9927);
nand UO_759 (O_759,N_9911,N_9991);
and UO_760 (O_760,N_9979,N_9951);
nor UO_761 (O_761,N_9981,N_9966);
or UO_762 (O_762,N_9959,N_9927);
and UO_763 (O_763,N_9930,N_9936);
nor UO_764 (O_764,N_9994,N_9966);
nor UO_765 (O_765,N_9978,N_9993);
and UO_766 (O_766,N_9959,N_9995);
nor UO_767 (O_767,N_9998,N_9954);
nand UO_768 (O_768,N_9948,N_9962);
and UO_769 (O_769,N_9987,N_9978);
nor UO_770 (O_770,N_9907,N_9904);
nand UO_771 (O_771,N_9932,N_9922);
or UO_772 (O_772,N_9933,N_9980);
and UO_773 (O_773,N_9923,N_9998);
and UO_774 (O_774,N_9986,N_9987);
and UO_775 (O_775,N_9910,N_9928);
xor UO_776 (O_776,N_9994,N_9930);
and UO_777 (O_777,N_9926,N_9983);
or UO_778 (O_778,N_9998,N_9990);
nand UO_779 (O_779,N_9995,N_9960);
nand UO_780 (O_780,N_9960,N_9927);
and UO_781 (O_781,N_9943,N_9909);
nand UO_782 (O_782,N_9917,N_9937);
nor UO_783 (O_783,N_9960,N_9926);
nand UO_784 (O_784,N_9998,N_9969);
and UO_785 (O_785,N_9907,N_9910);
nand UO_786 (O_786,N_9973,N_9969);
nand UO_787 (O_787,N_9987,N_9998);
or UO_788 (O_788,N_9914,N_9954);
or UO_789 (O_789,N_9989,N_9952);
nand UO_790 (O_790,N_9939,N_9967);
and UO_791 (O_791,N_9934,N_9993);
nor UO_792 (O_792,N_9964,N_9916);
or UO_793 (O_793,N_9938,N_9958);
nor UO_794 (O_794,N_9977,N_9941);
or UO_795 (O_795,N_9937,N_9964);
and UO_796 (O_796,N_9935,N_9912);
nor UO_797 (O_797,N_9998,N_9994);
and UO_798 (O_798,N_9957,N_9986);
nor UO_799 (O_799,N_9981,N_9904);
nor UO_800 (O_800,N_9969,N_9995);
and UO_801 (O_801,N_9967,N_9985);
nor UO_802 (O_802,N_9988,N_9970);
nor UO_803 (O_803,N_9950,N_9957);
nand UO_804 (O_804,N_9963,N_9917);
nand UO_805 (O_805,N_9949,N_9977);
and UO_806 (O_806,N_9936,N_9941);
nor UO_807 (O_807,N_9927,N_9931);
nand UO_808 (O_808,N_9950,N_9988);
nand UO_809 (O_809,N_9976,N_9900);
nand UO_810 (O_810,N_9945,N_9978);
nand UO_811 (O_811,N_9967,N_9924);
nand UO_812 (O_812,N_9929,N_9906);
nand UO_813 (O_813,N_9944,N_9920);
and UO_814 (O_814,N_9913,N_9957);
nor UO_815 (O_815,N_9934,N_9922);
nor UO_816 (O_816,N_9994,N_9903);
and UO_817 (O_817,N_9921,N_9928);
nand UO_818 (O_818,N_9920,N_9985);
xnor UO_819 (O_819,N_9994,N_9986);
nor UO_820 (O_820,N_9921,N_9994);
or UO_821 (O_821,N_9915,N_9979);
nor UO_822 (O_822,N_9939,N_9954);
or UO_823 (O_823,N_9976,N_9930);
and UO_824 (O_824,N_9926,N_9914);
or UO_825 (O_825,N_9918,N_9917);
nor UO_826 (O_826,N_9950,N_9930);
and UO_827 (O_827,N_9911,N_9930);
nor UO_828 (O_828,N_9954,N_9900);
and UO_829 (O_829,N_9962,N_9960);
nand UO_830 (O_830,N_9916,N_9982);
and UO_831 (O_831,N_9963,N_9921);
or UO_832 (O_832,N_9925,N_9900);
nor UO_833 (O_833,N_9927,N_9942);
nor UO_834 (O_834,N_9928,N_9989);
nand UO_835 (O_835,N_9917,N_9994);
xnor UO_836 (O_836,N_9949,N_9939);
or UO_837 (O_837,N_9908,N_9989);
and UO_838 (O_838,N_9935,N_9927);
nand UO_839 (O_839,N_9923,N_9978);
nor UO_840 (O_840,N_9957,N_9908);
nor UO_841 (O_841,N_9971,N_9956);
nand UO_842 (O_842,N_9963,N_9967);
nor UO_843 (O_843,N_9943,N_9945);
nor UO_844 (O_844,N_9915,N_9968);
or UO_845 (O_845,N_9953,N_9926);
and UO_846 (O_846,N_9995,N_9904);
nor UO_847 (O_847,N_9901,N_9910);
and UO_848 (O_848,N_9959,N_9921);
nor UO_849 (O_849,N_9974,N_9972);
and UO_850 (O_850,N_9980,N_9912);
and UO_851 (O_851,N_9950,N_9963);
nand UO_852 (O_852,N_9944,N_9996);
and UO_853 (O_853,N_9919,N_9932);
nor UO_854 (O_854,N_9977,N_9959);
or UO_855 (O_855,N_9936,N_9940);
nand UO_856 (O_856,N_9945,N_9948);
and UO_857 (O_857,N_9905,N_9918);
nor UO_858 (O_858,N_9996,N_9948);
nand UO_859 (O_859,N_9923,N_9999);
or UO_860 (O_860,N_9945,N_9953);
and UO_861 (O_861,N_9961,N_9950);
nand UO_862 (O_862,N_9973,N_9917);
nor UO_863 (O_863,N_9996,N_9985);
nor UO_864 (O_864,N_9905,N_9956);
or UO_865 (O_865,N_9932,N_9907);
nand UO_866 (O_866,N_9968,N_9946);
and UO_867 (O_867,N_9960,N_9921);
nor UO_868 (O_868,N_9935,N_9969);
nor UO_869 (O_869,N_9932,N_9985);
nor UO_870 (O_870,N_9931,N_9916);
and UO_871 (O_871,N_9906,N_9995);
nor UO_872 (O_872,N_9909,N_9919);
or UO_873 (O_873,N_9916,N_9971);
nor UO_874 (O_874,N_9939,N_9948);
nor UO_875 (O_875,N_9953,N_9994);
and UO_876 (O_876,N_9982,N_9967);
nand UO_877 (O_877,N_9956,N_9991);
or UO_878 (O_878,N_9916,N_9983);
nand UO_879 (O_879,N_9991,N_9986);
nand UO_880 (O_880,N_9974,N_9939);
or UO_881 (O_881,N_9998,N_9970);
nand UO_882 (O_882,N_9970,N_9922);
or UO_883 (O_883,N_9951,N_9903);
and UO_884 (O_884,N_9911,N_9958);
nand UO_885 (O_885,N_9966,N_9910);
nand UO_886 (O_886,N_9943,N_9907);
nor UO_887 (O_887,N_9957,N_9974);
and UO_888 (O_888,N_9949,N_9965);
or UO_889 (O_889,N_9961,N_9925);
and UO_890 (O_890,N_9900,N_9936);
nand UO_891 (O_891,N_9906,N_9927);
nand UO_892 (O_892,N_9994,N_9957);
nand UO_893 (O_893,N_9974,N_9968);
nand UO_894 (O_894,N_9925,N_9916);
and UO_895 (O_895,N_9954,N_9996);
nand UO_896 (O_896,N_9961,N_9936);
or UO_897 (O_897,N_9926,N_9922);
or UO_898 (O_898,N_9941,N_9963);
nor UO_899 (O_899,N_9913,N_9971);
xnor UO_900 (O_900,N_9939,N_9947);
and UO_901 (O_901,N_9989,N_9949);
or UO_902 (O_902,N_9991,N_9984);
or UO_903 (O_903,N_9951,N_9946);
or UO_904 (O_904,N_9981,N_9998);
and UO_905 (O_905,N_9909,N_9900);
nor UO_906 (O_906,N_9925,N_9946);
nand UO_907 (O_907,N_9926,N_9973);
and UO_908 (O_908,N_9917,N_9957);
or UO_909 (O_909,N_9964,N_9938);
and UO_910 (O_910,N_9948,N_9952);
and UO_911 (O_911,N_9915,N_9916);
nor UO_912 (O_912,N_9995,N_9973);
nor UO_913 (O_913,N_9947,N_9906);
nand UO_914 (O_914,N_9905,N_9946);
and UO_915 (O_915,N_9949,N_9980);
nand UO_916 (O_916,N_9906,N_9977);
nand UO_917 (O_917,N_9979,N_9988);
or UO_918 (O_918,N_9960,N_9908);
and UO_919 (O_919,N_9917,N_9986);
and UO_920 (O_920,N_9931,N_9900);
nand UO_921 (O_921,N_9953,N_9901);
nand UO_922 (O_922,N_9923,N_9930);
and UO_923 (O_923,N_9919,N_9924);
nand UO_924 (O_924,N_9936,N_9935);
and UO_925 (O_925,N_9987,N_9996);
xnor UO_926 (O_926,N_9967,N_9977);
nor UO_927 (O_927,N_9963,N_9984);
nand UO_928 (O_928,N_9925,N_9960);
xor UO_929 (O_929,N_9974,N_9907);
or UO_930 (O_930,N_9937,N_9908);
xnor UO_931 (O_931,N_9945,N_9986);
and UO_932 (O_932,N_9927,N_9964);
nor UO_933 (O_933,N_9932,N_9951);
nor UO_934 (O_934,N_9950,N_9919);
and UO_935 (O_935,N_9981,N_9946);
and UO_936 (O_936,N_9990,N_9956);
nor UO_937 (O_937,N_9937,N_9934);
nor UO_938 (O_938,N_9905,N_9951);
nor UO_939 (O_939,N_9909,N_9908);
or UO_940 (O_940,N_9947,N_9963);
nand UO_941 (O_941,N_9984,N_9921);
nand UO_942 (O_942,N_9919,N_9912);
nand UO_943 (O_943,N_9924,N_9943);
nand UO_944 (O_944,N_9932,N_9942);
xor UO_945 (O_945,N_9933,N_9974);
and UO_946 (O_946,N_9970,N_9973);
or UO_947 (O_947,N_9929,N_9994);
and UO_948 (O_948,N_9935,N_9945);
and UO_949 (O_949,N_9907,N_9954);
nor UO_950 (O_950,N_9937,N_9993);
or UO_951 (O_951,N_9913,N_9952);
nand UO_952 (O_952,N_9946,N_9988);
and UO_953 (O_953,N_9911,N_9917);
nor UO_954 (O_954,N_9911,N_9951);
nand UO_955 (O_955,N_9970,N_9940);
nor UO_956 (O_956,N_9920,N_9946);
nand UO_957 (O_957,N_9929,N_9953);
and UO_958 (O_958,N_9965,N_9912);
nor UO_959 (O_959,N_9900,N_9937);
nor UO_960 (O_960,N_9925,N_9968);
and UO_961 (O_961,N_9958,N_9977);
nand UO_962 (O_962,N_9935,N_9983);
nor UO_963 (O_963,N_9981,N_9941);
nor UO_964 (O_964,N_9959,N_9929);
or UO_965 (O_965,N_9905,N_9911);
or UO_966 (O_966,N_9930,N_9919);
and UO_967 (O_967,N_9968,N_9998);
or UO_968 (O_968,N_9951,N_9963);
nor UO_969 (O_969,N_9961,N_9920);
xnor UO_970 (O_970,N_9951,N_9939);
and UO_971 (O_971,N_9927,N_9996);
nand UO_972 (O_972,N_9900,N_9986);
nor UO_973 (O_973,N_9988,N_9917);
or UO_974 (O_974,N_9982,N_9942);
xor UO_975 (O_975,N_9914,N_9971);
or UO_976 (O_976,N_9967,N_9989);
and UO_977 (O_977,N_9984,N_9935);
or UO_978 (O_978,N_9984,N_9975);
or UO_979 (O_979,N_9991,N_9961);
and UO_980 (O_980,N_9970,N_9954);
and UO_981 (O_981,N_9961,N_9959);
or UO_982 (O_982,N_9927,N_9941);
nor UO_983 (O_983,N_9943,N_9936);
nor UO_984 (O_984,N_9933,N_9999);
nand UO_985 (O_985,N_9943,N_9930);
and UO_986 (O_986,N_9959,N_9911);
and UO_987 (O_987,N_9951,N_9942);
and UO_988 (O_988,N_9976,N_9971);
or UO_989 (O_989,N_9967,N_9956);
nor UO_990 (O_990,N_9925,N_9918);
nand UO_991 (O_991,N_9937,N_9974);
and UO_992 (O_992,N_9954,N_9935);
and UO_993 (O_993,N_9980,N_9955);
nor UO_994 (O_994,N_9950,N_9942);
and UO_995 (O_995,N_9918,N_9962);
nor UO_996 (O_996,N_9939,N_9996);
or UO_997 (O_997,N_9939,N_9922);
or UO_998 (O_998,N_9941,N_9940);
or UO_999 (O_999,N_9993,N_9906);
and UO_1000 (O_1000,N_9950,N_9912);
nand UO_1001 (O_1001,N_9954,N_9967);
or UO_1002 (O_1002,N_9962,N_9994);
nand UO_1003 (O_1003,N_9947,N_9982);
or UO_1004 (O_1004,N_9978,N_9952);
or UO_1005 (O_1005,N_9963,N_9981);
and UO_1006 (O_1006,N_9923,N_9906);
or UO_1007 (O_1007,N_9973,N_9997);
or UO_1008 (O_1008,N_9910,N_9978);
and UO_1009 (O_1009,N_9929,N_9900);
or UO_1010 (O_1010,N_9923,N_9908);
nor UO_1011 (O_1011,N_9935,N_9964);
nand UO_1012 (O_1012,N_9969,N_9983);
or UO_1013 (O_1013,N_9998,N_9976);
nor UO_1014 (O_1014,N_9924,N_9921);
and UO_1015 (O_1015,N_9968,N_9917);
nor UO_1016 (O_1016,N_9969,N_9948);
or UO_1017 (O_1017,N_9917,N_9954);
nand UO_1018 (O_1018,N_9937,N_9984);
nor UO_1019 (O_1019,N_9973,N_9956);
xnor UO_1020 (O_1020,N_9948,N_9938);
xor UO_1021 (O_1021,N_9952,N_9975);
nand UO_1022 (O_1022,N_9966,N_9901);
nand UO_1023 (O_1023,N_9992,N_9985);
and UO_1024 (O_1024,N_9947,N_9931);
xnor UO_1025 (O_1025,N_9968,N_9955);
or UO_1026 (O_1026,N_9969,N_9960);
and UO_1027 (O_1027,N_9994,N_9951);
nand UO_1028 (O_1028,N_9912,N_9916);
or UO_1029 (O_1029,N_9954,N_9955);
nand UO_1030 (O_1030,N_9919,N_9991);
and UO_1031 (O_1031,N_9989,N_9922);
and UO_1032 (O_1032,N_9953,N_9936);
and UO_1033 (O_1033,N_9915,N_9946);
and UO_1034 (O_1034,N_9973,N_9920);
and UO_1035 (O_1035,N_9973,N_9979);
nor UO_1036 (O_1036,N_9909,N_9982);
nand UO_1037 (O_1037,N_9990,N_9935);
or UO_1038 (O_1038,N_9923,N_9985);
and UO_1039 (O_1039,N_9969,N_9947);
nand UO_1040 (O_1040,N_9928,N_9966);
nor UO_1041 (O_1041,N_9997,N_9949);
or UO_1042 (O_1042,N_9904,N_9956);
or UO_1043 (O_1043,N_9992,N_9967);
and UO_1044 (O_1044,N_9989,N_9917);
or UO_1045 (O_1045,N_9913,N_9940);
or UO_1046 (O_1046,N_9955,N_9966);
or UO_1047 (O_1047,N_9970,N_9935);
and UO_1048 (O_1048,N_9965,N_9933);
or UO_1049 (O_1049,N_9948,N_9980);
nor UO_1050 (O_1050,N_9901,N_9905);
nor UO_1051 (O_1051,N_9920,N_9965);
or UO_1052 (O_1052,N_9926,N_9944);
or UO_1053 (O_1053,N_9979,N_9958);
nand UO_1054 (O_1054,N_9917,N_9902);
nor UO_1055 (O_1055,N_9984,N_9978);
or UO_1056 (O_1056,N_9902,N_9960);
or UO_1057 (O_1057,N_9950,N_9962);
or UO_1058 (O_1058,N_9903,N_9997);
nand UO_1059 (O_1059,N_9925,N_9959);
or UO_1060 (O_1060,N_9926,N_9937);
nor UO_1061 (O_1061,N_9918,N_9930);
nand UO_1062 (O_1062,N_9955,N_9979);
nor UO_1063 (O_1063,N_9999,N_9959);
nor UO_1064 (O_1064,N_9907,N_9925);
nand UO_1065 (O_1065,N_9919,N_9977);
or UO_1066 (O_1066,N_9975,N_9993);
or UO_1067 (O_1067,N_9971,N_9949);
nor UO_1068 (O_1068,N_9949,N_9934);
and UO_1069 (O_1069,N_9909,N_9952);
or UO_1070 (O_1070,N_9939,N_9942);
or UO_1071 (O_1071,N_9980,N_9939);
or UO_1072 (O_1072,N_9923,N_9907);
xnor UO_1073 (O_1073,N_9902,N_9992);
nand UO_1074 (O_1074,N_9939,N_9924);
or UO_1075 (O_1075,N_9944,N_9907);
or UO_1076 (O_1076,N_9965,N_9985);
or UO_1077 (O_1077,N_9926,N_9978);
or UO_1078 (O_1078,N_9948,N_9981);
nand UO_1079 (O_1079,N_9993,N_9915);
nand UO_1080 (O_1080,N_9941,N_9935);
or UO_1081 (O_1081,N_9906,N_9978);
and UO_1082 (O_1082,N_9954,N_9934);
nor UO_1083 (O_1083,N_9918,N_9903);
nand UO_1084 (O_1084,N_9938,N_9973);
or UO_1085 (O_1085,N_9965,N_9942);
nand UO_1086 (O_1086,N_9971,N_9946);
nand UO_1087 (O_1087,N_9986,N_9963);
or UO_1088 (O_1088,N_9957,N_9912);
nand UO_1089 (O_1089,N_9972,N_9927);
nor UO_1090 (O_1090,N_9985,N_9946);
or UO_1091 (O_1091,N_9900,N_9934);
or UO_1092 (O_1092,N_9972,N_9964);
nor UO_1093 (O_1093,N_9960,N_9949);
or UO_1094 (O_1094,N_9994,N_9938);
nor UO_1095 (O_1095,N_9911,N_9996);
and UO_1096 (O_1096,N_9908,N_9922);
nand UO_1097 (O_1097,N_9969,N_9942);
and UO_1098 (O_1098,N_9992,N_9912);
nor UO_1099 (O_1099,N_9941,N_9945);
and UO_1100 (O_1100,N_9998,N_9928);
or UO_1101 (O_1101,N_9996,N_9968);
nor UO_1102 (O_1102,N_9900,N_9945);
nand UO_1103 (O_1103,N_9935,N_9986);
or UO_1104 (O_1104,N_9990,N_9993);
nor UO_1105 (O_1105,N_9937,N_9904);
nor UO_1106 (O_1106,N_9930,N_9945);
or UO_1107 (O_1107,N_9911,N_9987);
and UO_1108 (O_1108,N_9916,N_9955);
or UO_1109 (O_1109,N_9966,N_9962);
and UO_1110 (O_1110,N_9984,N_9904);
or UO_1111 (O_1111,N_9981,N_9992);
or UO_1112 (O_1112,N_9925,N_9903);
or UO_1113 (O_1113,N_9937,N_9938);
nor UO_1114 (O_1114,N_9947,N_9994);
nand UO_1115 (O_1115,N_9972,N_9970);
and UO_1116 (O_1116,N_9982,N_9923);
and UO_1117 (O_1117,N_9900,N_9901);
or UO_1118 (O_1118,N_9943,N_9916);
nand UO_1119 (O_1119,N_9965,N_9975);
nand UO_1120 (O_1120,N_9956,N_9959);
or UO_1121 (O_1121,N_9929,N_9973);
nor UO_1122 (O_1122,N_9977,N_9954);
nand UO_1123 (O_1123,N_9929,N_9938);
nand UO_1124 (O_1124,N_9912,N_9934);
or UO_1125 (O_1125,N_9910,N_9919);
nor UO_1126 (O_1126,N_9908,N_9925);
or UO_1127 (O_1127,N_9935,N_9955);
nand UO_1128 (O_1128,N_9992,N_9987);
nor UO_1129 (O_1129,N_9984,N_9901);
nand UO_1130 (O_1130,N_9965,N_9906);
and UO_1131 (O_1131,N_9926,N_9918);
or UO_1132 (O_1132,N_9932,N_9938);
and UO_1133 (O_1133,N_9934,N_9960);
and UO_1134 (O_1134,N_9986,N_9947);
and UO_1135 (O_1135,N_9925,N_9901);
nand UO_1136 (O_1136,N_9942,N_9906);
xnor UO_1137 (O_1137,N_9998,N_9933);
nor UO_1138 (O_1138,N_9987,N_9931);
nand UO_1139 (O_1139,N_9920,N_9978);
nand UO_1140 (O_1140,N_9933,N_9906);
nand UO_1141 (O_1141,N_9985,N_9902);
nand UO_1142 (O_1142,N_9934,N_9910);
and UO_1143 (O_1143,N_9989,N_9921);
nand UO_1144 (O_1144,N_9930,N_9920);
nor UO_1145 (O_1145,N_9936,N_9981);
and UO_1146 (O_1146,N_9951,N_9970);
nor UO_1147 (O_1147,N_9937,N_9946);
nand UO_1148 (O_1148,N_9903,N_9981);
or UO_1149 (O_1149,N_9934,N_9918);
nand UO_1150 (O_1150,N_9932,N_9941);
nand UO_1151 (O_1151,N_9908,N_9952);
nor UO_1152 (O_1152,N_9938,N_9949);
and UO_1153 (O_1153,N_9909,N_9911);
nor UO_1154 (O_1154,N_9902,N_9984);
or UO_1155 (O_1155,N_9995,N_9903);
nor UO_1156 (O_1156,N_9986,N_9904);
and UO_1157 (O_1157,N_9941,N_9992);
or UO_1158 (O_1158,N_9999,N_9958);
nand UO_1159 (O_1159,N_9965,N_9931);
or UO_1160 (O_1160,N_9906,N_9944);
or UO_1161 (O_1161,N_9918,N_9993);
and UO_1162 (O_1162,N_9902,N_9997);
and UO_1163 (O_1163,N_9968,N_9989);
nor UO_1164 (O_1164,N_9962,N_9931);
and UO_1165 (O_1165,N_9934,N_9999);
nor UO_1166 (O_1166,N_9918,N_9955);
nand UO_1167 (O_1167,N_9963,N_9934);
or UO_1168 (O_1168,N_9938,N_9998);
and UO_1169 (O_1169,N_9912,N_9968);
nand UO_1170 (O_1170,N_9941,N_9988);
nor UO_1171 (O_1171,N_9919,N_9983);
or UO_1172 (O_1172,N_9969,N_9924);
and UO_1173 (O_1173,N_9923,N_9989);
nor UO_1174 (O_1174,N_9914,N_9975);
or UO_1175 (O_1175,N_9908,N_9963);
or UO_1176 (O_1176,N_9972,N_9967);
nor UO_1177 (O_1177,N_9905,N_9907);
and UO_1178 (O_1178,N_9948,N_9959);
nand UO_1179 (O_1179,N_9918,N_9940);
nor UO_1180 (O_1180,N_9933,N_9995);
and UO_1181 (O_1181,N_9947,N_9995);
xor UO_1182 (O_1182,N_9932,N_9977);
and UO_1183 (O_1183,N_9915,N_9981);
and UO_1184 (O_1184,N_9959,N_9945);
or UO_1185 (O_1185,N_9959,N_9917);
and UO_1186 (O_1186,N_9941,N_9934);
or UO_1187 (O_1187,N_9939,N_9921);
and UO_1188 (O_1188,N_9954,N_9938);
nor UO_1189 (O_1189,N_9982,N_9976);
and UO_1190 (O_1190,N_9992,N_9970);
nand UO_1191 (O_1191,N_9920,N_9935);
or UO_1192 (O_1192,N_9923,N_9926);
or UO_1193 (O_1193,N_9944,N_9968);
nand UO_1194 (O_1194,N_9915,N_9953);
nor UO_1195 (O_1195,N_9945,N_9996);
and UO_1196 (O_1196,N_9944,N_9948);
nor UO_1197 (O_1197,N_9970,N_9919);
nand UO_1198 (O_1198,N_9970,N_9900);
nand UO_1199 (O_1199,N_9933,N_9992);
and UO_1200 (O_1200,N_9981,N_9957);
or UO_1201 (O_1201,N_9991,N_9927);
nor UO_1202 (O_1202,N_9947,N_9921);
and UO_1203 (O_1203,N_9951,N_9927);
or UO_1204 (O_1204,N_9926,N_9956);
nand UO_1205 (O_1205,N_9928,N_9923);
or UO_1206 (O_1206,N_9903,N_9915);
nand UO_1207 (O_1207,N_9951,N_9918);
and UO_1208 (O_1208,N_9941,N_9982);
nor UO_1209 (O_1209,N_9960,N_9933);
or UO_1210 (O_1210,N_9975,N_9935);
or UO_1211 (O_1211,N_9965,N_9971);
nor UO_1212 (O_1212,N_9943,N_9944);
and UO_1213 (O_1213,N_9993,N_9944);
and UO_1214 (O_1214,N_9985,N_9918);
nor UO_1215 (O_1215,N_9974,N_9919);
nor UO_1216 (O_1216,N_9998,N_9956);
and UO_1217 (O_1217,N_9988,N_9934);
or UO_1218 (O_1218,N_9950,N_9954);
or UO_1219 (O_1219,N_9939,N_9927);
or UO_1220 (O_1220,N_9996,N_9990);
nor UO_1221 (O_1221,N_9931,N_9992);
and UO_1222 (O_1222,N_9904,N_9971);
nand UO_1223 (O_1223,N_9902,N_9946);
nand UO_1224 (O_1224,N_9958,N_9967);
nor UO_1225 (O_1225,N_9970,N_9921);
nor UO_1226 (O_1226,N_9931,N_9989);
nand UO_1227 (O_1227,N_9919,N_9931);
and UO_1228 (O_1228,N_9918,N_9920);
or UO_1229 (O_1229,N_9908,N_9954);
or UO_1230 (O_1230,N_9966,N_9987);
and UO_1231 (O_1231,N_9968,N_9919);
nor UO_1232 (O_1232,N_9962,N_9920);
nand UO_1233 (O_1233,N_9986,N_9932);
nor UO_1234 (O_1234,N_9973,N_9981);
and UO_1235 (O_1235,N_9946,N_9963);
or UO_1236 (O_1236,N_9919,N_9903);
nor UO_1237 (O_1237,N_9951,N_9937);
nor UO_1238 (O_1238,N_9960,N_9943);
or UO_1239 (O_1239,N_9976,N_9992);
and UO_1240 (O_1240,N_9969,N_9915);
nor UO_1241 (O_1241,N_9995,N_9991);
nor UO_1242 (O_1242,N_9906,N_9938);
nor UO_1243 (O_1243,N_9909,N_9972);
nand UO_1244 (O_1244,N_9927,N_9948);
and UO_1245 (O_1245,N_9941,N_9916);
or UO_1246 (O_1246,N_9927,N_9925);
or UO_1247 (O_1247,N_9946,N_9970);
nand UO_1248 (O_1248,N_9903,N_9941);
nand UO_1249 (O_1249,N_9909,N_9947);
nand UO_1250 (O_1250,N_9946,N_9908);
and UO_1251 (O_1251,N_9933,N_9969);
or UO_1252 (O_1252,N_9906,N_9971);
nand UO_1253 (O_1253,N_9929,N_9950);
nor UO_1254 (O_1254,N_9954,N_9973);
nor UO_1255 (O_1255,N_9906,N_9910);
and UO_1256 (O_1256,N_9927,N_9997);
or UO_1257 (O_1257,N_9900,N_9987);
nand UO_1258 (O_1258,N_9965,N_9914);
or UO_1259 (O_1259,N_9981,N_9984);
nor UO_1260 (O_1260,N_9939,N_9975);
and UO_1261 (O_1261,N_9988,N_9925);
xnor UO_1262 (O_1262,N_9901,N_9973);
nor UO_1263 (O_1263,N_9918,N_9919);
nor UO_1264 (O_1264,N_9972,N_9957);
nor UO_1265 (O_1265,N_9922,N_9960);
or UO_1266 (O_1266,N_9983,N_9973);
and UO_1267 (O_1267,N_9954,N_9966);
nand UO_1268 (O_1268,N_9994,N_9923);
and UO_1269 (O_1269,N_9908,N_9901);
and UO_1270 (O_1270,N_9937,N_9914);
nand UO_1271 (O_1271,N_9994,N_9996);
nand UO_1272 (O_1272,N_9964,N_9983);
and UO_1273 (O_1273,N_9988,N_9997);
nand UO_1274 (O_1274,N_9996,N_9953);
or UO_1275 (O_1275,N_9949,N_9942);
and UO_1276 (O_1276,N_9930,N_9912);
and UO_1277 (O_1277,N_9969,N_9941);
nor UO_1278 (O_1278,N_9975,N_9958);
nand UO_1279 (O_1279,N_9904,N_9931);
nand UO_1280 (O_1280,N_9914,N_9908);
nand UO_1281 (O_1281,N_9900,N_9973);
and UO_1282 (O_1282,N_9917,N_9999);
nor UO_1283 (O_1283,N_9954,N_9925);
nor UO_1284 (O_1284,N_9912,N_9944);
and UO_1285 (O_1285,N_9950,N_9927);
nand UO_1286 (O_1286,N_9918,N_9937);
and UO_1287 (O_1287,N_9914,N_9994);
nor UO_1288 (O_1288,N_9903,N_9978);
or UO_1289 (O_1289,N_9914,N_9997);
nand UO_1290 (O_1290,N_9915,N_9956);
or UO_1291 (O_1291,N_9906,N_9992);
and UO_1292 (O_1292,N_9909,N_9917);
or UO_1293 (O_1293,N_9955,N_9953);
nand UO_1294 (O_1294,N_9971,N_9919);
or UO_1295 (O_1295,N_9915,N_9984);
and UO_1296 (O_1296,N_9980,N_9919);
nand UO_1297 (O_1297,N_9991,N_9957);
nand UO_1298 (O_1298,N_9978,N_9922);
nor UO_1299 (O_1299,N_9910,N_9900);
nor UO_1300 (O_1300,N_9991,N_9904);
nand UO_1301 (O_1301,N_9916,N_9910);
or UO_1302 (O_1302,N_9902,N_9939);
nor UO_1303 (O_1303,N_9951,N_9907);
nor UO_1304 (O_1304,N_9962,N_9934);
nand UO_1305 (O_1305,N_9997,N_9972);
or UO_1306 (O_1306,N_9939,N_9976);
nor UO_1307 (O_1307,N_9970,N_9944);
or UO_1308 (O_1308,N_9937,N_9980);
nand UO_1309 (O_1309,N_9977,N_9966);
or UO_1310 (O_1310,N_9970,N_9977);
nand UO_1311 (O_1311,N_9979,N_9971);
nor UO_1312 (O_1312,N_9981,N_9945);
or UO_1313 (O_1313,N_9913,N_9917);
or UO_1314 (O_1314,N_9904,N_9969);
or UO_1315 (O_1315,N_9904,N_9951);
nor UO_1316 (O_1316,N_9996,N_9980);
or UO_1317 (O_1317,N_9917,N_9985);
nor UO_1318 (O_1318,N_9983,N_9995);
and UO_1319 (O_1319,N_9936,N_9916);
and UO_1320 (O_1320,N_9910,N_9955);
and UO_1321 (O_1321,N_9941,N_9971);
and UO_1322 (O_1322,N_9985,N_9936);
nor UO_1323 (O_1323,N_9916,N_9917);
nor UO_1324 (O_1324,N_9961,N_9909);
and UO_1325 (O_1325,N_9919,N_9958);
nand UO_1326 (O_1326,N_9943,N_9959);
nand UO_1327 (O_1327,N_9942,N_9940);
or UO_1328 (O_1328,N_9964,N_9953);
or UO_1329 (O_1329,N_9951,N_9976);
or UO_1330 (O_1330,N_9919,N_9955);
nand UO_1331 (O_1331,N_9954,N_9911);
nor UO_1332 (O_1332,N_9945,N_9909);
and UO_1333 (O_1333,N_9936,N_9914);
nor UO_1334 (O_1334,N_9922,N_9918);
or UO_1335 (O_1335,N_9962,N_9951);
nor UO_1336 (O_1336,N_9942,N_9954);
and UO_1337 (O_1337,N_9936,N_9967);
or UO_1338 (O_1338,N_9941,N_9926);
or UO_1339 (O_1339,N_9903,N_9962);
nand UO_1340 (O_1340,N_9934,N_9909);
nand UO_1341 (O_1341,N_9992,N_9913);
xnor UO_1342 (O_1342,N_9966,N_9903);
nor UO_1343 (O_1343,N_9990,N_9971);
nand UO_1344 (O_1344,N_9976,N_9931);
nand UO_1345 (O_1345,N_9977,N_9939);
and UO_1346 (O_1346,N_9950,N_9975);
and UO_1347 (O_1347,N_9971,N_9970);
or UO_1348 (O_1348,N_9929,N_9989);
and UO_1349 (O_1349,N_9989,N_9926);
and UO_1350 (O_1350,N_9915,N_9904);
nand UO_1351 (O_1351,N_9903,N_9958);
or UO_1352 (O_1352,N_9902,N_9948);
nand UO_1353 (O_1353,N_9926,N_9948);
and UO_1354 (O_1354,N_9935,N_9915);
and UO_1355 (O_1355,N_9995,N_9982);
nor UO_1356 (O_1356,N_9965,N_9997);
or UO_1357 (O_1357,N_9938,N_9970);
and UO_1358 (O_1358,N_9997,N_9987);
and UO_1359 (O_1359,N_9934,N_9970);
nor UO_1360 (O_1360,N_9959,N_9910);
or UO_1361 (O_1361,N_9957,N_9924);
and UO_1362 (O_1362,N_9978,N_9959);
and UO_1363 (O_1363,N_9927,N_9985);
nand UO_1364 (O_1364,N_9989,N_9913);
nand UO_1365 (O_1365,N_9907,N_9939);
nor UO_1366 (O_1366,N_9934,N_9983);
nor UO_1367 (O_1367,N_9985,N_9988);
or UO_1368 (O_1368,N_9955,N_9949);
or UO_1369 (O_1369,N_9935,N_9972);
nor UO_1370 (O_1370,N_9902,N_9974);
nor UO_1371 (O_1371,N_9935,N_9991);
nand UO_1372 (O_1372,N_9949,N_9957);
nor UO_1373 (O_1373,N_9976,N_9950);
and UO_1374 (O_1374,N_9993,N_9916);
and UO_1375 (O_1375,N_9966,N_9929);
nand UO_1376 (O_1376,N_9977,N_9948);
nor UO_1377 (O_1377,N_9915,N_9908);
nand UO_1378 (O_1378,N_9970,N_9930);
or UO_1379 (O_1379,N_9997,N_9960);
and UO_1380 (O_1380,N_9924,N_9962);
or UO_1381 (O_1381,N_9988,N_9922);
nand UO_1382 (O_1382,N_9982,N_9935);
and UO_1383 (O_1383,N_9984,N_9949);
or UO_1384 (O_1384,N_9921,N_9956);
or UO_1385 (O_1385,N_9965,N_9905);
nand UO_1386 (O_1386,N_9933,N_9918);
nand UO_1387 (O_1387,N_9928,N_9956);
nor UO_1388 (O_1388,N_9902,N_9999);
or UO_1389 (O_1389,N_9990,N_9960);
nor UO_1390 (O_1390,N_9900,N_9921);
or UO_1391 (O_1391,N_9995,N_9931);
nand UO_1392 (O_1392,N_9983,N_9909);
or UO_1393 (O_1393,N_9940,N_9991);
nor UO_1394 (O_1394,N_9960,N_9920);
and UO_1395 (O_1395,N_9944,N_9913);
nand UO_1396 (O_1396,N_9930,N_9981);
xor UO_1397 (O_1397,N_9974,N_9998);
nand UO_1398 (O_1398,N_9958,N_9972);
nor UO_1399 (O_1399,N_9946,N_9983);
and UO_1400 (O_1400,N_9980,N_9917);
xnor UO_1401 (O_1401,N_9921,N_9941);
xor UO_1402 (O_1402,N_9927,N_9983);
or UO_1403 (O_1403,N_9923,N_9976);
or UO_1404 (O_1404,N_9941,N_9964);
nand UO_1405 (O_1405,N_9935,N_9965);
nand UO_1406 (O_1406,N_9944,N_9957);
xor UO_1407 (O_1407,N_9991,N_9933);
or UO_1408 (O_1408,N_9948,N_9970);
nor UO_1409 (O_1409,N_9967,N_9910);
nor UO_1410 (O_1410,N_9953,N_9951);
and UO_1411 (O_1411,N_9985,N_9980);
nand UO_1412 (O_1412,N_9900,N_9956);
and UO_1413 (O_1413,N_9907,N_9946);
nand UO_1414 (O_1414,N_9964,N_9939);
nor UO_1415 (O_1415,N_9979,N_9946);
and UO_1416 (O_1416,N_9965,N_9901);
nor UO_1417 (O_1417,N_9972,N_9903);
and UO_1418 (O_1418,N_9973,N_9988);
or UO_1419 (O_1419,N_9936,N_9964);
nor UO_1420 (O_1420,N_9902,N_9949);
or UO_1421 (O_1421,N_9939,N_9957);
and UO_1422 (O_1422,N_9938,N_9993);
and UO_1423 (O_1423,N_9996,N_9958);
or UO_1424 (O_1424,N_9975,N_9995);
nand UO_1425 (O_1425,N_9988,N_9916);
nor UO_1426 (O_1426,N_9904,N_9966);
and UO_1427 (O_1427,N_9968,N_9945);
and UO_1428 (O_1428,N_9980,N_9929);
nor UO_1429 (O_1429,N_9937,N_9948);
nand UO_1430 (O_1430,N_9948,N_9967);
nor UO_1431 (O_1431,N_9971,N_9953);
xnor UO_1432 (O_1432,N_9941,N_9975);
nand UO_1433 (O_1433,N_9954,N_9916);
nand UO_1434 (O_1434,N_9961,N_9918);
and UO_1435 (O_1435,N_9918,N_9989);
nand UO_1436 (O_1436,N_9952,N_9962);
nor UO_1437 (O_1437,N_9929,N_9965);
nand UO_1438 (O_1438,N_9960,N_9910);
or UO_1439 (O_1439,N_9996,N_9961);
or UO_1440 (O_1440,N_9979,N_9948);
and UO_1441 (O_1441,N_9943,N_9925);
xnor UO_1442 (O_1442,N_9967,N_9976);
nor UO_1443 (O_1443,N_9983,N_9920);
and UO_1444 (O_1444,N_9969,N_9911);
nand UO_1445 (O_1445,N_9912,N_9973);
or UO_1446 (O_1446,N_9917,N_9935);
nor UO_1447 (O_1447,N_9963,N_9904);
and UO_1448 (O_1448,N_9927,N_9936);
nand UO_1449 (O_1449,N_9991,N_9998);
and UO_1450 (O_1450,N_9971,N_9931);
nor UO_1451 (O_1451,N_9915,N_9936);
nor UO_1452 (O_1452,N_9941,N_9938);
nand UO_1453 (O_1453,N_9900,N_9971);
or UO_1454 (O_1454,N_9922,N_9920);
nand UO_1455 (O_1455,N_9928,N_9919);
and UO_1456 (O_1456,N_9935,N_9974);
or UO_1457 (O_1457,N_9996,N_9906);
nand UO_1458 (O_1458,N_9915,N_9933);
or UO_1459 (O_1459,N_9964,N_9902);
or UO_1460 (O_1460,N_9999,N_9972);
and UO_1461 (O_1461,N_9975,N_9903);
or UO_1462 (O_1462,N_9903,N_9992);
and UO_1463 (O_1463,N_9900,N_9943);
nor UO_1464 (O_1464,N_9966,N_9969);
nor UO_1465 (O_1465,N_9917,N_9904);
nor UO_1466 (O_1466,N_9925,N_9976);
nor UO_1467 (O_1467,N_9958,N_9982);
nor UO_1468 (O_1468,N_9919,N_9964);
nand UO_1469 (O_1469,N_9904,N_9900);
and UO_1470 (O_1470,N_9964,N_9980);
nor UO_1471 (O_1471,N_9922,N_9995);
nor UO_1472 (O_1472,N_9987,N_9958);
nand UO_1473 (O_1473,N_9944,N_9947);
nand UO_1474 (O_1474,N_9985,N_9943);
nand UO_1475 (O_1475,N_9995,N_9989);
or UO_1476 (O_1476,N_9968,N_9962);
and UO_1477 (O_1477,N_9949,N_9953);
and UO_1478 (O_1478,N_9917,N_9901);
nor UO_1479 (O_1479,N_9962,N_9993);
nand UO_1480 (O_1480,N_9910,N_9948);
and UO_1481 (O_1481,N_9952,N_9931);
and UO_1482 (O_1482,N_9977,N_9986);
or UO_1483 (O_1483,N_9958,N_9929);
or UO_1484 (O_1484,N_9928,N_9938);
nor UO_1485 (O_1485,N_9964,N_9926);
nor UO_1486 (O_1486,N_9904,N_9927);
nand UO_1487 (O_1487,N_9907,N_9917);
and UO_1488 (O_1488,N_9974,N_9947);
or UO_1489 (O_1489,N_9946,N_9972);
nor UO_1490 (O_1490,N_9910,N_9949);
nand UO_1491 (O_1491,N_9998,N_9979);
nand UO_1492 (O_1492,N_9913,N_9929);
and UO_1493 (O_1493,N_9994,N_9911);
and UO_1494 (O_1494,N_9911,N_9985);
xor UO_1495 (O_1495,N_9988,N_9949);
nor UO_1496 (O_1496,N_9902,N_9903);
or UO_1497 (O_1497,N_9942,N_9963);
or UO_1498 (O_1498,N_9988,N_9959);
or UO_1499 (O_1499,N_9965,N_9968);
endmodule