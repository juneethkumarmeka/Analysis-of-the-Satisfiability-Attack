module basic_2500_25000_3000_8_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_1626,In_486);
or U1 (N_1,In_810,In_1951);
nand U2 (N_2,In_11,In_475);
nor U3 (N_3,In_1400,In_1660);
xor U4 (N_4,In_194,In_78);
nor U5 (N_5,In_2260,In_1827);
or U6 (N_6,In_1601,In_1316);
nor U7 (N_7,In_647,In_714);
nand U8 (N_8,In_2460,In_2335);
nor U9 (N_9,In_1539,In_2011);
and U10 (N_10,In_1063,In_1489);
nand U11 (N_11,In_1867,In_291);
or U12 (N_12,In_914,In_1932);
or U13 (N_13,In_1862,In_808);
nand U14 (N_14,In_1227,In_2114);
nor U15 (N_15,In_1040,In_1217);
nor U16 (N_16,In_1977,In_1282);
and U17 (N_17,In_772,In_1308);
nand U18 (N_18,In_180,In_1831);
nor U19 (N_19,In_1385,In_695);
or U20 (N_20,In_2322,In_1826);
xor U21 (N_21,In_1098,In_1651);
or U22 (N_22,In_1224,In_2004);
nand U23 (N_23,In_2222,In_826);
nand U24 (N_24,In_251,In_1243);
and U25 (N_25,In_940,In_1418);
or U26 (N_26,In_1212,In_690);
or U27 (N_27,In_2394,In_173);
nor U28 (N_28,In_598,In_2443);
and U29 (N_29,In_2051,In_1680);
or U30 (N_30,In_101,In_1136);
xnor U31 (N_31,In_2223,In_2248);
xor U32 (N_32,In_2361,In_2093);
nand U33 (N_33,In_1646,In_1863);
and U34 (N_34,In_1786,In_75);
nor U35 (N_35,In_1958,In_1600);
nand U36 (N_36,In_245,In_1065);
or U37 (N_37,In_1384,In_89);
and U38 (N_38,In_1182,In_2070);
nor U39 (N_39,In_287,In_1046);
nand U40 (N_40,In_1256,In_374);
nand U41 (N_41,In_611,In_165);
or U42 (N_42,In_1787,In_2404);
nand U43 (N_43,In_2221,In_1604);
nor U44 (N_44,In_579,In_1440);
or U45 (N_45,In_2364,In_1568);
nor U46 (N_46,In_599,In_1861);
nand U47 (N_47,In_1115,In_2353);
or U48 (N_48,In_448,In_1934);
or U49 (N_49,In_2284,In_151);
and U50 (N_50,In_566,In_2005);
or U51 (N_51,In_83,In_1128);
or U52 (N_52,In_921,In_1573);
nor U53 (N_53,In_2037,In_2031);
nor U54 (N_54,In_136,In_1696);
nand U55 (N_55,In_1535,In_924);
or U56 (N_56,In_945,In_2342);
nor U57 (N_57,In_458,In_2239);
nand U58 (N_58,In_1043,In_237);
or U59 (N_59,In_60,In_390);
nor U60 (N_60,In_1843,In_1733);
nor U61 (N_61,In_986,In_2432);
and U62 (N_62,In_3,In_1691);
nor U63 (N_63,In_1850,In_1255);
or U64 (N_64,In_167,In_2403);
nor U65 (N_65,In_2198,In_295);
xnor U66 (N_66,In_1774,In_466);
nor U67 (N_67,In_126,In_1642);
xnor U68 (N_68,In_510,In_1302);
nand U69 (N_69,In_1513,In_322);
or U70 (N_70,In_1470,In_2344);
xnor U71 (N_71,In_1178,In_1961);
or U72 (N_72,In_660,In_65);
and U73 (N_73,In_158,In_1355);
nand U74 (N_74,In_1454,In_2481);
nand U75 (N_75,In_1715,In_2163);
nor U76 (N_76,In_1703,In_20);
xor U77 (N_77,In_32,In_987);
xnor U78 (N_78,In_1526,In_1238);
or U79 (N_79,In_2339,In_112);
nand U80 (N_80,In_1198,In_1174);
nand U81 (N_81,In_2234,In_2467);
xor U82 (N_82,In_2013,In_204);
xnor U83 (N_83,In_1929,In_2428);
nand U84 (N_84,In_1710,In_1779);
xnor U85 (N_85,In_1578,In_2391);
nand U86 (N_86,In_590,In_329);
and U87 (N_87,In_567,In_2319);
nand U88 (N_88,In_1666,In_2263);
or U89 (N_89,In_28,In_2162);
and U90 (N_90,In_903,In_854);
and U91 (N_91,In_1148,In_2369);
xor U92 (N_92,In_885,In_1986);
or U93 (N_93,In_845,In_2139);
or U94 (N_94,In_1373,In_1744);
or U95 (N_95,In_1451,In_668);
nand U96 (N_96,In_1589,In_82);
nand U97 (N_97,In_201,In_1156);
and U98 (N_98,In_1001,In_493);
or U99 (N_99,In_164,In_271);
or U100 (N_100,In_902,In_1802);
nand U101 (N_101,In_424,In_310);
nor U102 (N_102,In_444,In_827);
xor U103 (N_103,In_163,In_2420);
nand U104 (N_104,In_2079,In_1821);
nor U105 (N_105,In_1806,In_168);
nor U106 (N_106,In_1270,In_587);
and U107 (N_107,In_1448,In_554);
or U108 (N_108,In_775,In_1197);
xor U109 (N_109,In_1165,In_621);
nor U110 (N_110,In_953,In_104);
or U111 (N_111,In_831,In_898);
nor U112 (N_112,In_111,In_482);
or U113 (N_113,In_169,In_1189);
and U114 (N_114,In_942,In_1177);
and U115 (N_115,In_1566,In_879);
or U116 (N_116,In_1588,In_2053);
nor U117 (N_117,In_1816,In_2459);
nand U118 (N_118,In_1887,In_1413);
nand U119 (N_119,In_1899,In_1619);
nand U120 (N_120,In_1858,In_1202);
nor U121 (N_121,In_1902,In_2132);
and U122 (N_122,In_264,In_2461);
nand U123 (N_123,In_1503,In_1621);
nor U124 (N_124,In_1324,In_402);
nor U125 (N_125,In_634,In_742);
or U126 (N_126,In_1488,In_248);
xnor U127 (N_127,In_1277,In_1290);
or U128 (N_128,In_1331,In_1580);
nor U129 (N_129,In_1123,In_1127);
and U130 (N_130,In_1879,In_1328);
or U131 (N_131,In_1403,In_55);
or U132 (N_132,In_425,In_2110);
or U133 (N_133,In_629,In_2279);
and U134 (N_134,In_2450,In_882);
or U135 (N_135,In_891,In_1995);
nand U136 (N_136,In_1339,In_662);
nand U137 (N_137,In_1714,In_1145);
nand U138 (N_138,In_1649,In_584);
and U139 (N_139,In_1504,In_819);
and U140 (N_140,In_2097,In_132);
nand U141 (N_141,In_128,In_1812);
nand U142 (N_142,In_1734,In_330);
or U143 (N_143,In_2276,In_1069);
nand U144 (N_144,In_354,In_821);
or U145 (N_145,In_1250,In_1124);
nand U146 (N_146,In_2499,In_2156);
nor U147 (N_147,In_594,In_1447);
or U148 (N_148,In_376,In_571);
nand U149 (N_149,In_619,In_883);
nand U150 (N_150,In_706,In_575);
nand U151 (N_151,In_1967,In_964);
nor U152 (N_152,In_24,In_2010);
nand U153 (N_153,In_2111,In_2167);
nand U154 (N_154,In_130,In_2495);
nor U155 (N_155,In_347,In_2323);
nand U156 (N_156,In_997,In_754);
nand U157 (N_157,In_67,In_2257);
nor U158 (N_158,In_1976,In_266);
nand U159 (N_159,In_1367,In_2253);
or U160 (N_160,In_2038,In_1882);
or U161 (N_161,In_1775,In_1880);
or U162 (N_162,In_377,In_1438);
and U163 (N_163,In_1778,In_865);
or U164 (N_164,In_428,In_367);
xnor U165 (N_165,In_544,In_1999);
nor U166 (N_166,In_1397,In_622);
nand U167 (N_167,In_1251,In_728);
nor U168 (N_168,In_363,In_490);
or U169 (N_169,In_72,In_1372);
or U170 (N_170,In_1591,In_1970);
and U171 (N_171,In_263,In_1293);
nand U172 (N_172,In_1519,In_1275);
nor U173 (N_173,In_2451,In_1630);
or U174 (N_174,In_679,In_336);
or U175 (N_175,In_733,In_1204);
nand U176 (N_176,In_92,In_2085);
and U177 (N_177,In_2392,In_1664);
and U178 (N_178,In_944,In_1991);
and U179 (N_179,In_119,In_1450);
and U180 (N_180,In_1638,In_1603);
or U181 (N_181,In_1670,In_1808);
nor U182 (N_182,In_228,In_1186);
or U183 (N_183,In_1602,In_1482);
nor U184 (N_184,In_2042,In_1942);
and U185 (N_185,In_2147,In_325);
or U186 (N_186,In_37,In_149);
nor U187 (N_187,In_1110,In_643);
or U188 (N_188,In_2272,In_497);
nand U189 (N_189,In_1349,In_1449);
nor U190 (N_190,In_1966,In_1752);
nor U191 (N_191,In_227,In_1644);
nor U192 (N_192,In_743,In_721);
nor U193 (N_193,In_121,In_957);
xnor U194 (N_194,In_2425,In_698);
nand U195 (N_195,In_1549,In_1835);
nor U196 (N_196,In_1908,In_2023);
and U197 (N_197,In_703,In_923);
nor U198 (N_198,In_2411,In_423);
nand U199 (N_199,In_1502,In_303);
or U200 (N_200,In_793,In_1878);
nand U201 (N_201,In_1868,In_1654);
xor U202 (N_202,In_1254,In_2164);
nor U203 (N_203,In_2422,In_2048);
nand U204 (N_204,In_1841,In_1709);
nor U205 (N_205,In_820,In_371);
nand U206 (N_206,In_2380,In_514);
or U207 (N_207,In_1429,In_937);
and U208 (N_208,In_1390,In_1337);
nor U209 (N_209,In_1239,In_326);
and U210 (N_210,In_528,In_2088);
nand U211 (N_211,In_176,In_816);
nand U212 (N_212,In_2265,In_1102);
and U213 (N_213,In_1490,In_480);
and U214 (N_214,In_404,In_2205);
nand U215 (N_215,In_1894,In_2103);
xor U216 (N_216,In_1772,In_1719);
and U217 (N_217,In_2485,In_782);
or U218 (N_218,In_1939,In_1129);
or U219 (N_219,In_2184,In_40);
nand U220 (N_220,In_632,In_747);
nand U221 (N_221,In_2145,In_655);
xor U222 (N_222,In_2402,In_186);
nor U223 (N_223,In_463,In_1980);
nor U224 (N_224,In_2343,In_1329);
and U225 (N_225,In_676,In_935);
and U226 (N_226,In_368,In_2328);
nor U227 (N_227,In_2213,In_1469);
nand U228 (N_228,In_1954,In_1739);
xnor U229 (N_229,In_2295,In_1071);
nor U230 (N_230,In_351,In_2362);
nand U231 (N_231,In_1528,In_2413);
xnor U232 (N_232,In_539,In_1419);
xnor U233 (N_233,In_1045,In_1062);
or U234 (N_234,In_392,In_1788);
nand U235 (N_235,In_1996,In_1678);
or U236 (N_236,In_1311,In_2439);
and U237 (N_237,In_94,In_2405);
nand U238 (N_238,In_77,In_389);
and U239 (N_239,In_2182,In_829);
nor U240 (N_240,In_1221,In_1640);
or U241 (N_241,In_1381,In_114);
and U242 (N_242,In_1893,In_1789);
xnor U243 (N_243,In_1699,In_289);
and U244 (N_244,In_850,In_2129);
and U245 (N_245,In_2141,In_732);
or U246 (N_246,In_2293,In_456);
xnor U247 (N_247,In_1753,In_265);
and U248 (N_248,In_499,In_5);
or U249 (N_249,In_1889,In_10);
xor U250 (N_250,In_1936,In_1938);
nor U251 (N_251,In_2017,In_2027);
or U252 (N_252,In_370,In_1697);
nand U253 (N_253,In_1134,In_537);
nor U254 (N_254,In_438,In_515);
and U255 (N_255,In_779,In_17);
nand U256 (N_256,In_2202,In_177);
xor U257 (N_257,In_1348,In_1014);
xor U258 (N_258,In_1416,In_1633);
and U259 (N_259,In_1498,In_727);
nand U260 (N_260,In_1013,In_859);
xnor U261 (N_261,In_1499,In_1560);
nand U262 (N_262,In_1915,In_27);
nor U263 (N_263,In_2055,In_316);
or U264 (N_264,In_1721,In_578);
and U265 (N_265,In_1012,In_1183);
nor U266 (N_266,In_2130,In_185);
and U267 (N_267,In_2122,In_1582);
and U268 (N_268,In_2312,In_449);
nor U269 (N_269,In_2421,In_625);
and U270 (N_270,In_946,In_1673);
and U271 (N_271,In_1532,In_1520);
or U272 (N_272,In_1229,In_1852);
and U273 (N_273,In_443,In_1022);
or U274 (N_274,In_976,In_1953);
nor U275 (N_275,In_644,In_2483);
xor U276 (N_276,In_519,In_453);
and U277 (N_277,In_56,In_993);
nand U278 (N_278,In_1473,In_563);
and U279 (N_279,In_1848,In_858);
or U280 (N_280,In_1314,In_1810);
xor U281 (N_281,In_877,In_474);
nand U282 (N_282,In_2188,In_2146);
and U283 (N_283,In_2271,In_1394);
nor U284 (N_284,In_1048,In_1446);
xnor U285 (N_285,In_1836,In_551);
or U286 (N_286,In_321,In_1360);
nand U287 (N_287,In_2030,In_572);
or U288 (N_288,In_1614,In_1162);
nor U289 (N_289,In_64,In_1661);
nor U290 (N_290,In_699,In_2259);
nor U291 (N_291,In_426,In_835);
nand U292 (N_292,In_2197,In_1656);
nor U293 (N_293,In_1587,In_451);
nand U294 (N_294,In_1109,In_2326);
nor U295 (N_295,In_791,In_1326);
nor U296 (N_296,In_1682,In_1155);
and U297 (N_297,In_1572,In_596);
and U298 (N_298,In_1800,In_1032);
or U299 (N_299,In_1437,In_530);
nor U300 (N_300,In_229,In_1292);
nor U301 (N_301,In_1087,In_1305);
and U302 (N_302,In_508,In_211);
nand U303 (N_303,In_281,In_1598);
and U304 (N_304,In_2333,In_1782);
and U305 (N_305,In_150,In_1785);
or U306 (N_306,In_1401,In_70);
nor U307 (N_307,In_124,In_1100);
nand U308 (N_308,In_117,In_2406);
xor U309 (N_309,In_837,In_1439);
and U310 (N_310,In_760,In_1428);
and U311 (N_311,In_43,In_592);
or U312 (N_312,In_2207,In_863);
or U313 (N_313,In_200,In_1791);
nand U314 (N_314,In_2061,In_1702);
and U315 (N_315,In_171,In_1933);
or U316 (N_316,In_2099,In_758);
xor U317 (N_317,In_535,In_1625);
xor U318 (N_318,In_1635,In_191);
xor U319 (N_319,In_2477,In_777);
nor U320 (N_320,In_756,In_1610);
and U321 (N_321,In_2454,In_454);
nor U322 (N_322,In_1571,In_1956);
nor U323 (N_323,In_80,In_1295);
xor U324 (N_324,In_69,In_1839);
or U325 (N_325,In_7,In_255);
nand U326 (N_326,In_958,In_642);
xnor U327 (N_327,In_1613,In_306);
nor U328 (N_328,In_763,In_2287);
and U329 (N_329,In_31,In_1998);
nand U330 (N_330,In_118,In_250);
nor U331 (N_331,In_1284,In_851);
nor U332 (N_332,In_2250,In_682);
nor U333 (N_333,In_1180,In_2009);
nand U334 (N_334,In_1125,In_1257);
nand U335 (N_335,In_973,In_933);
nand U336 (N_336,In_9,In_2166);
nor U337 (N_337,In_492,In_1840);
nor U338 (N_338,In_1622,In_1727);
and U339 (N_339,In_1259,In_2315);
and U340 (N_340,In_2270,In_627);
and U341 (N_341,In_1246,In_1725);
nand U342 (N_342,In_403,In_350);
and U343 (N_343,In_1442,In_1232);
and U344 (N_344,In_1693,In_1236);
nor U345 (N_345,In_2463,In_1010);
nand U346 (N_346,In_678,In_1283);
xor U347 (N_347,In_154,In_8);
xor U348 (N_348,In_109,In_794);
nor U349 (N_349,In_1056,In_1493);
or U350 (N_350,In_2302,In_523);
nand U351 (N_351,In_418,In_187);
nor U352 (N_352,In_860,In_1960);
or U353 (N_353,In_39,In_2064);
and U354 (N_354,In_1459,In_538);
or U355 (N_355,In_1631,In_2006);
nand U356 (N_356,In_1496,In_215);
xnor U357 (N_357,In_1456,In_225);
or U358 (N_358,In_1741,In_138);
or U359 (N_359,In_2080,In_1139);
nand U360 (N_360,In_2448,In_34);
nand U361 (N_361,In_529,In_1859);
and U362 (N_362,In_704,In_1216);
and U363 (N_363,In_1007,In_233);
nand U364 (N_364,In_1694,In_1971);
or U365 (N_365,In_2498,In_1481);
nor U366 (N_366,In_1167,In_911);
nand U367 (N_367,In_1805,In_1468);
nor U368 (N_368,In_1088,In_1815);
and U369 (N_369,In_1120,In_1423);
nand U370 (N_370,In_2034,In_527);
nand U371 (N_371,In_1756,In_2497);
nor U372 (N_372,In_445,In_195);
nor U373 (N_373,In_765,In_894);
xnor U374 (N_374,In_1769,In_1405);
and U375 (N_375,In_897,In_844);
and U376 (N_376,In_1888,In_1313);
and U377 (N_377,In_1837,In_2220);
nor U378 (N_378,In_716,In_1132);
or U379 (N_379,In_1946,In_1793);
nor U380 (N_380,In_1795,In_343);
and U381 (N_381,In_996,In_2346);
nor U382 (N_382,In_362,In_2252);
xor U383 (N_383,In_2212,In_1406);
nor U384 (N_384,In_1105,In_333);
and U385 (N_385,In_1924,In_297);
and U386 (N_386,In_963,In_48);
nor U387 (N_387,In_2058,In_1854);
and U388 (N_388,In_518,In_434);
nand U389 (N_389,In_1285,In_1595);
nand U390 (N_390,In_1819,In_2219);
nand U391 (N_391,In_948,In_809);
xnor U392 (N_392,In_905,In_436);
xnor U393 (N_393,In_2415,In_90);
nand U394 (N_394,In_875,In_2142);
and U395 (N_395,In_1914,In_188);
and U396 (N_396,In_1818,In_1424);
or U397 (N_397,In_2032,In_1975);
or U398 (N_398,In_240,In_2424);
nand U399 (N_399,In_505,In_670);
nor U400 (N_400,In_1479,In_1191);
nand U401 (N_401,In_597,In_46);
or U402 (N_402,In_1463,In_1411);
nor U403 (N_403,In_696,In_2381);
xnor U404 (N_404,In_1435,In_1506);
nand U405 (N_405,In_2452,In_2359);
nor U406 (N_406,In_1597,In_1478);
nand U407 (N_407,In_2230,In_1092);
or U408 (N_408,In_1336,In_974);
nand U409 (N_409,In_926,In_134);
and U410 (N_410,In_414,In_2201);
or U411 (N_411,In_712,In_144);
nand U412 (N_412,In_677,In_1611);
nand U413 (N_413,In_1949,In_2441);
nand U414 (N_414,In_1193,In_58);
or U415 (N_415,In_774,In_2087);
and U416 (N_416,In_410,In_1296);
or U417 (N_417,In_1781,In_1555);
and U418 (N_418,In_719,In_1567);
and U419 (N_419,In_1742,In_1138);
nor U420 (N_420,In_1935,In_205);
and U421 (N_421,In_1833,In_1306);
xnor U422 (N_422,In_99,In_666);
xor U423 (N_423,In_998,In_2444);
or U424 (N_424,In_1323,In_1672);
nand U425 (N_425,In_1577,In_1195);
nand U426 (N_426,In_2178,In_113);
or U427 (N_427,In_2083,In_1135);
and U428 (N_428,In_62,In_284);
or U429 (N_429,In_1090,In_1652);
or U430 (N_430,In_2476,In_1210);
or U431 (N_431,In_904,In_2008);
and U432 (N_432,In_1223,In_2455);
nand U433 (N_433,In_1414,In_839);
and U434 (N_434,In_628,In_1757);
nor U435 (N_435,In_2482,In_1073);
nand U436 (N_436,In_2280,In_1300);
xor U437 (N_437,In_2352,In_586);
nand U438 (N_438,In_2154,In_697);
nor U439 (N_439,In_1031,In_2149);
and U440 (N_440,In_618,In_1466);
nor U441 (N_441,In_318,In_522);
nor U442 (N_442,In_1546,In_1807);
xnor U443 (N_443,In_36,In_559);
xnor U444 (N_444,In_1562,In_496);
and U445 (N_445,In_1759,In_657);
nor U446 (N_446,In_1773,In_561);
or U447 (N_447,In_41,In_1157);
nand U448 (N_448,In_2187,In_2417);
xnor U449 (N_449,In_715,In_100);
nor U450 (N_450,In_853,In_2261);
xnor U451 (N_451,In_2041,In_1000);
or U452 (N_452,In_680,In_1609);
nand U453 (N_453,In_1718,In_2321);
and U454 (N_454,In_388,In_1226);
nand U455 (N_455,In_219,In_665);
nand U456 (N_456,In_304,In_1495);
nand U457 (N_457,In_593,In_1052);
xor U458 (N_458,In_1559,In_954);
nand U459 (N_459,In_2233,In_710);
nand U460 (N_460,In_842,In_534);
and U461 (N_461,In_1901,In_1025);
and U462 (N_462,In_1099,In_604);
or U463 (N_463,In_1126,In_2474);
or U464 (N_464,In_2128,In_2063);
or U465 (N_465,In_2116,In_1443);
nor U466 (N_466,In_2269,In_1972);
nor U467 (N_467,In_2372,In_1273);
nor U468 (N_468,In_1093,In_2398);
and U469 (N_469,In_1671,In_2283);
or U470 (N_470,In_2386,In_2310);
xnor U471 (N_471,In_1851,In_2356);
or U472 (N_472,In_1679,In_383);
or U473 (N_473,In_524,In_739);
xnor U474 (N_474,In_1172,In_895);
nand U475 (N_475,In_2365,In_1377);
xor U476 (N_476,In_541,In_871);
or U477 (N_477,In_1334,In_1445);
nor U478 (N_478,In_762,In_701);
xnor U479 (N_479,In_833,In_1017);
and U480 (N_480,In_1564,In_1768);
nor U481 (N_481,In_900,In_2077);
and U482 (N_482,In_1783,In_1036);
nor U483 (N_483,In_2375,In_956);
nand U484 (N_484,In_1338,In_276);
and U485 (N_485,In_718,In_1813);
or U486 (N_486,In_1199,In_1750);
nor U487 (N_487,In_2399,In_568);
nand U488 (N_488,In_1291,In_1077);
nand U489 (N_489,In_1639,In_2376);
nor U490 (N_490,In_2371,In_674);
xor U491 (N_491,In_830,In_2026);
nand U492 (N_492,In_1985,In_2236);
or U493 (N_493,In_920,In_348);
xor U494 (N_494,In_2100,In_1379);
and U495 (N_495,In_405,In_750);
nand U496 (N_496,In_1235,In_1276);
nand U497 (N_497,In_941,In_2277);
nand U498 (N_498,In_1507,In_884);
or U499 (N_499,In_1085,In_1517);
or U500 (N_500,In_1267,In_148);
nor U501 (N_501,In_189,In_1857);
or U502 (N_502,In_51,In_2330);
or U503 (N_503,In_2062,In_1776);
and U504 (N_504,In_1369,In_1231);
nor U505 (N_505,In_759,In_1095);
and U506 (N_506,In_320,In_936);
xor U507 (N_507,In_548,In_1289);
xor U508 (N_508,In_1215,In_873);
or U509 (N_509,In_487,In_110);
nand U510 (N_510,In_1278,In_2374);
or U511 (N_511,In_2021,In_1133);
or U512 (N_512,In_1108,In_1537);
nor U513 (N_513,In_1796,In_2494);
xnor U514 (N_514,In_2307,In_127);
or U515 (N_515,In_1245,In_1408);
nor U516 (N_516,In_2232,In_108);
or U517 (N_517,In_2126,In_441);
nand U518 (N_518,In_1847,In_197);
and U519 (N_519,In_2473,In_2349);
nor U520 (N_520,In_2320,In_260);
and U521 (N_521,In_1327,In_1016);
nand U522 (N_522,In_1253,In_1542);
nand U523 (N_523,In_1067,In_1814);
nand U524 (N_524,In_971,In_683);
and U525 (N_525,In_1681,In_1160);
nor U526 (N_526,In_2290,In_938);
nand U527 (N_527,In_1911,In_2408);
nor U528 (N_528,In_640,In_1616);
or U529 (N_529,In_723,In_477);
nor U530 (N_530,In_283,In_671);
or U531 (N_531,In_2466,In_707);
nand U532 (N_532,In_1990,In_1515);
or U533 (N_533,In_2479,In_1989);
or U534 (N_534,In_1486,In_2227);
and U535 (N_535,In_840,In_531);
or U536 (N_536,In_1317,In_275);
nand U537 (N_537,In_437,In_342);
and U538 (N_538,In_2057,In_23);
or U539 (N_539,In_355,In_253);
xnor U540 (N_540,In_1342,In_272);
nand U541 (N_541,In_1075,In_912);
nand U542 (N_542,In_93,In_771);
and U543 (N_543,In_2350,In_74);
nor U544 (N_544,In_328,In_1545);
and U545 (N_545,In_1955,In_1002);
xnor U546 (N_546,In_2183,In_1551);
nor U547 (N_547,In_1467,In_408);
xor U548 (N_548,In_872,In_980);
nand U549 (N_549,In_981,In_335);
nor U550 (N_550,In_2496,In_1386);
nor U551 (N_551,In_966,In_653);
nor U552 (N_552,In_314,In_1747);
nor U553 (N_553,In_1175,In_1866);
nand U554 (N_554,In_14,In_1082);
xnor U555 (N_555,In_1540,In_1398);
or U556 (N_556,In_2228,In_1387);
nor U557 (N_557,In_1608,In_992);
or U558 (N_558,In_1920,In_79);
and U559 (N_559,In_382,In_613);
xnor U560 (N_560,In_1474,In_896);
or U561 (N_561,In_2436,In_207);
and U562 (N_562,In_2311,In_1286);
or U563 (N_563,In_778,In_1460);
and U564 (N_564,In_364,In_2136);
nand U565 (N_565,In_595,In_1049);
nor U566 (N_566,In_481,In_1181);
nor U567 (N_567,In_1143,In_1883);
nor U568 (N_568,In_1892,In_1068);
and U569 (N_569,In_1751,In_1505);
nor U570 (N_570,In_1820,In_692);
and U571 (N_571,In_360,In_1720);
nand U572 (N_572,In_746,In_462);
nor U573 (N_573,In_417,In_413);
xor U574 (N_574,In_2324,In_1089);
nor U575 (N_575,In_1230,In_1834);
nand U576 (N_576,In_558,In_856);
or U577 (N_577,In_2303,In_1556);
and U578 (N_578,In_1122,In_838);
and U579 (N_579,In_1310,In_874);
or U580 (N_580,In_2363,In_736);
xor U581 (N_581,In_800,In_2095);
nor U582 (N_582,In_279,In_2433);
nand U583 (N_583,In_1205,In_1033);
or U584 (N_584,In_852,In_421);
or U585 (N_585,In_1350,In_1228);
xor U586 (N_586,In_1207,In_789);
nor U587 (N_587,In_502,In_2275);
xor U588 (N_588,In_889,In_790);
xor U589 (N_589,In_2189,In_2148);
nand U590 (N_590,In_1558,In_2066);
nand U591 (N_591,In_560,In_1570);
and U592 (N_592,In_1365,In_1575);
and U593 (N_593,In_582,In_1957);
nand U594 (N_594,In_120,In_1020);
nor U595 (N_595,In_1299,In_1728);
or U596 (N_596,In_583,In_103);
nor U597 (N_597,In_145,In_274);
and U598 (N_598,In_292,In_533);
xnor U599 (N_599,In_1797,In_1615);
xor U600 (N_600,In_2193,In_2067);
nor U601 (N_601,In_507,In_1058);
or U602 (N_602,In_2355,In_2262);
nand U603 (N_603,In_1173,In_691);
nor U604 (N_604,In_967,In_133);
nand U605 (N_605,In_1521,In_479);
and U606 (N_606,In_549,In_131);
or U607 (N_607,In_241,In_1897);
xor U608 (N_608,In_1149,In_1599);
or U609 (N_609,In_234,In_1116);
nor U610 (N_610,In_218,In_13);
nor U611 (N_611,In_1344,In_300);
and U612 (N_612,In_345,In_1382);
or U613 (N_613,In_553,In_147);
or U614 (N_614,In_1484,In_44);
or U615 (N_615,In_630,In_2133);
nand U616 (N_616,In_2285,In_1978);
xor U617 (N_617,In_2449,In_929);
nand U618 (N_618,In_526,In_1525);
or U619 (N_619,In_1804,In_1341);
and U620 (N_620,In_2426,In_669);
or U621 (N_621,In_2069,In_1919);
nand U622 (N_622,In_722,In_447);
and U623 (N_623,In_1366,In_1121);
nor U624 (N_624,In_521,In_246);
nor U625 (N_625,In_1973,In_262);
or U626 (N_626,In_1131,In_1891);
nand U627 (N_627,In_489,In_861);
nor U628 (N_628,In_1988,In_1677);
xnor U629 (N_629,In_1817,In_1898);
xor U630 (N_630,In_532,In_2416);
nand U631 (N_631,In_2074,In_2181);
nor U632 (N_632,In_908,In_71);
nand U633 (N_633,In_1926,In_1005);
or U634 (N_634,In_1119,In_278);
nor U635 (N_635,In_1554,In_547);
or U636 (N_636,In_495,In_1737);
xor U637 (N_637,In_162,In_1716);
nand U638 (N_638,In_1396,In_1111);
xor U639 (N_639,In_1628,In_1322);
and U640 (N_640,In_1606,In_2059);
and U641 (N_641,In_542,In_857);
and U642 (N_642,In_472,In_751);
and U643 (N_643,In_214,In_2469);
nor U644 (N_644,In_1233,In_1021);
xnor U645 (N_645,In_1931,In_473);
and U646 (N_646,In_2264,In_764);
nor U647 (N_647,In_1307,In_641);
nor U648 (N_648,In_1059,In_1070);
nor U649 (N_649,In_91,In_491);
or U650 (N_650,In_419,In_427);
nand U651 (N_651,In_2089,In_2336);
nor U652 (N_652,In_1907,In_232);
xor U653 (N_653,In_2470,In_672);
xnor U654 (N_654,In_1219,In_1304);
nand U655 (N_655,In_626,In_1590);
nor U656 (N_656,In_749,In_452);
and U657 (N_657,In_2268,In_268);
nor U658 (N_658,In_57,In_2243);
nor U659 (N_659,In_1508,In_769);
or U660 (N_660,In_525,In_429);
and U661 (N_661,In_901,In_1359);
nor U662 (N_662,In_29,In_1501);
and U663 (N_663,In_757,In_1708);
and U664 (N_664,In_298,In_729);
or U665 (N_665,In_1809,In_254);
nand U666 (N_666,In_2423,In_1864);
xor U667 (N_667,In_2211,In_1712);
xor U668 (N_668,In_2194,In_6);
nor U669 (N_669,In_2165,In_317);
and U670 (N_670,In_1393,In_994);
nor U671 (N_671,In_708,In_440);
or U672 (N_672,In_16,In_880);
or U673 (N_673,In_1910,In_2401);
or U674 (N_674,In_1909,In_2119);
nor U675 (N_675,In_1683,In_2192);
nand U676 (N_676,In_509,In_1363);
and U677 (N_677,In_1011,In_1828);
xnor U678 (N_678,In_1055,In_422);
or U679 (N_679,In_2082,In_646);
nor U680 (N_680,In_238,In_2106);
xnor U681 (N_681,In_498,In_1345);
and U682 (N_682,In_2414,In_962);
and U683 (N_683,In_1147,In_1745);
nand U684 (N_684,In_309,In_61);
nand U685 (N_685,In_2191,In_1700);
xnor U686 (N_686,In_1927,In_890);
xor U687 (N_687,In_1655,In_652);
and U688 (N_688,In_1096,In_1748);
nor U689 (N_689,In_1192,In_1890);
or U690 (N_690,In_288,In_2073);
nor U691 (N_691,In_1144,In_2292);
nor U692 (N_692,In_2155,In_1767);
nand U693 (N_693,In_927,In_192);
nor U694 (N_694,In_2171,In_286);
and U695 (N_695,In_2431,In_307);
or U696 (N_696,In_931,In_1689);
nor U697 (N_697,In_1168,In_2159);
or U698 (N_698,In_1066,In_1035);
nand U699 (N_699,In_988,In_1112);
or U700 (N_700,In_2033,In_734);
or U701 (N_701,In_1364,In_357);
xnor U702 (N_702,In_97,In_784);
nand U703 (N_703,In_836,In_506);
and U704 (N_704,In_658,In_2313);
nor U705 (N_705,In_483,In_88);
nand U706 (N_706,In_745,In_1190);
nand U707 (N_707,In_45,In_1354);
or U708 (N_708,In_2289,In_1531);
nor U709 (N_709,In_1981,In_589);
nor U710 (N_710,In_1770,In_1303);
and U711 (N_711,In_1320,In_2172);
and U712 (N_712,In_577,In_143);
xor U713 (N_713,In_2338,In_1028);
and U714 (N_714,In_261,In_797);
nor U715 (N_715,In_2384,In_2049);
nor U716 (N_716,In_792,In_157);
and U717 (N_717,In_925,In_600);
xnor U718 (N_718,In_1853,In_802);
nand U719 (N_719,In_893,In_869);
nor U720 (N_720,In_435,In_1433);
nand U721 (N_721,In_1262,In_1579);
and U722 (N_722,In_1563,In_2435);
and U723 (N_723,In_359,In_1476);
and U724 (N_724,In_2304,In_1086);
nor U725 (N_725,In_324,In_807);
nor U726 (N_726,In_142,In_1220);
nor U727 (N_727,In_1659,In_624);
nand U728 (N_728,In_244,In_2102);
xnor U729 (N_729,In_1674,In_1030);
nor U730 (N_730,In_959,In_2170);
or U731 (N_731,In_620,In_1754);
or U732 (N_732,In_1494,In_2409);
or U733 (N_733,In_1461,In_1550);
and U734 (N_734,In_2267,In_1856);
and U735 (N_735,In_2241,In_1301);
nand U736 (N_736,In_461,In_1798);
or U737 (N_737,In_977,In_1916);
or U738 (N_738,In_955,In_87);
xnor U739 (N_739,In_1399,In_2115);
nor U740 (N_740,In_1176,In_2478);
nor U741 (N_741,In_1885,In_720);
xor U742 (N_742,In_0,In_2112);
and U743 (N_743,In_1346,In_1184);
nor U744 (N_744,In_1024,In_35);
and U745 (N_745,In_932,In_2072);
nor U746 (N_746,In_2332,In_834);
nor U747 (N_747,In_2429,In_947);
nand U748 (N_748,In_2462,In_338);
or U749 (N_749,In_1979,In_478);
or U750 (N_750,In_2229,In_96);
nand U751 (N_751,In_1876,In_406);
or U752 (N_752,In_2160,In_1676);
nor U753 (N_753,In_2291,In_323);
or U754 (N_754,In_565,In_19);
and U755 (N_755,In_2412,In_25);
nor U756 (N_756,In_805,In_803);
and U757 (N_757,In_781,In_2316);
or U758 (N_758,In_770,In_580);
and U759 (N_759,In_290,In_385);
nand U760 (N_760,In_270,In_1441);
or U761 (N_761,In_832,In_2340);
nor U762 (N_762,In_569,In_950);
or U763 (N_763,In_258,In_1650);
nor U764 (N_764,In_2081,In_1794);
and U765 (N_765,In_2168,In_2296);
or U766 (N_766,In_1458,In_785);
or U767 (N_767,In_213,In_381);
nor U768 (N_768,In_1380,In_555);
nor U769 (N_769,In_2493,In_1081);
or U770 (N_770,In_106,In_450);
and U771 (N_771,In_934,In_1258);
or U772 (N_772,In_1574,In_726);
nand U773 (N_773,In_1006,In_433);
or U774 (N_774,In_2124,In_1019);
nor U775 (N_775,In_1612,In_2484);
nor U776 (N_776,In_1872,In_1203);
and U777 (N_777,In_1675,In_2242);
and U778 (N_778,In_603,In_1886);
or U779 (N_779,In_1480,In_768);
or U780 (N_780,In_1298,In_2176);
or U781 (N_781,In_196,In_681);
or U782 (N_782,In_1263,In_1008);
and U783 (N_783,In_183,In_1895);
nand U784 (N_784,In_2367,In_512);
nand U785 (N_785,In_1266,In_1658);
nor U786 (N_786,In_965,In_892);
or U787 (N_787,In_398,In_1596);
or U788 (N_788,In_649,In_54);
nor U789 (N_789,In_1483,In_741);
nand U790 (N_790,In_631,In_1663);
or U791 (N_791,In_1717,In_2107);
and U792 (N_792,In_1705,In_1351);
or U793 (N_793,In_42,In_235);
and U794 (N_794,In_1607,In_1758);
xor U795 (N_795,In_285,In_1994);
nand U796 (N_796,In_1777,In_282);
nor U797 (N_797,In_1050,In_2);
xnor U798 (N_798,In_1417,In_1179);
and U799 (N_799,In_2442,In_1803);
nand U800 (N_800,In_471,In_312);
nand U801 (N_801,In_1874,In_2209);
nor U802 (N_802,In_1018,In_2468);
nor U803 (N_803,In_1208,In_787);
nor U804 (N_804,In_753,In_1247);
xor U805 (N_805,In_1527,In_991);
nand U806 (N_806,In_1151,In_1761);
nor U807 (N_807,In_504,In_2254);
xor U808 (N_808,In_1309,In_1343);
or U809 (N_809,In_1690,In_239);
or U810 (N_810,In_1206,In_344);
nand U811 (N_811,In_2123,In_1865);
or U812 (N_812,In_1335,In_2086);
nand U813 (N_813,In_1623,In_2022);
nand U814 (N_814,In_95,In_86);
or U815 (N_815,In_53,In_1244);
nand U816 (N_816,In_1565,In_230);
and U817 (N_817,In_2224,In_928);
and U818 (N_818,In_899,In_1287);
nand U819 (N_819,In_2179,In_1544);
nand U820 (N_820,In_66,In_1378);
nor U821 (N_821,In_411,In_2177);
nor U822 (N_822,In_2487,In_617);
or U823 (N_823,In_1,In_1740);
or U824 (N_824,In_1104,In_4);
nand U825 (N_825,In_2308,In_2354);
or U826 (N_826,In_2091,In_340);
and U827 (N_827,In_702,In_2245);
and U828 (N_828,In_2266,In_1462);
nor U829 (N_829,In_2127,In_146);
xnor U830 (N_830,In_2020,In_1618);
nor U831 (N_831,In_1557,In_1352);
nor U832 (N_832,In_2153,In_1707);
xor U833 (N_833,In_1509,In_1464);
nand U834 (N_834,In_1457,In_1041);
nor U835 (N_835,In_2306,In_585);
or U836 (N_836,In_1605,In_1332);
nand U837 (N_837,In_1315,In_748);
xnor U838 (N_838,In_713,In_876);
and U839 (N_839,In_724,In_814);
nand U840 (N_840,In_1425,In_21);
and U841 (N_841,In_1743,In_574);
and U842 (N_842,In_581,In_1940);
nand U843 (N_843,In_744,In_2370);
nand U844 (N_844,In_1749,In_1917);
and U845 (N_845,In_1844,In_294);
or U846 (N_846,In_1510,In_1047);
or U847 (N_847,In_651,In_795);
and U848 (N_848,In_1079,In_1569);
and U849 (N_849,In_2288,In_1518);
nand U850 (N_850,In_2383,In_1665);
and U851 (N_851,In_1669,In_125);
and U852 (N_852,In_212,In_552);
or U853 (N_853,In_484,In_1042);
nor U854 (N_854,In_2134,In_2373);
and U855 (N_855,In_1729,In_786);
nor U856 (N_856,In_1097,In_494);
nor U857 (N_857,In_2419,In_1799);
or U858 (N_858,In_2471,In_1142);
nor U859 (N_859,In_960,In_2445);
and U860 (N_860,In_280,In_1522);
or U861 (N_861,In_137,In_1617);
or U862 (N_862,In_105,In_610);
nand U863 (N_863,In_2090,In_1392);
nand U864 (N_864,In_1222,In_2195);
and U865 (N_865,In_1294,In_2393);
xnor U866 (N_866,In_684,In_1407);
and U867 (N_867,In_1492,In_469);
nand U868 (N_868,In_1792,In_2458);
nand U869 (N_869,In_1213,In_1074);
nor U870 (N_870,In_982,In_667);
nand U871 (N_871,In_2175,In_783);
nor U872 (N_872,In_301,In_731);
xor U873 (N_873,In_788,In_1388);
nand U874 (N_874,In_1117,In_315);
and U875 (N_875,In_906,In_415);
nor U876 (N_876,In_2121,In_1297);
nor U877 (N_877,In_711,In_1003);
or U878 (N_878,In_50,In_1027);
nand U879 (N_879,In_1593,In_601);
and U880 (N_880,In_2186,In_2035);
or U881 (N_881,In_2056,In_1163);
or U882 (N_882,In_267,In_1692);
or U883 (N_883,In_216,In_2185);
nand U884 (N_884,In_2040,In_256);
nand U885 (N_885,In_1913,In_2237);
or U886 (N_886,In_208,In_1060);
nand U887 (N_887,In_2273,In_47);
nand U888 (N_888,In_2137,In_868);
or U889 (N_889,In_22,In_650);
nor U890 (N_890,In_2475,In_1430);
and U891 (N_891,In_1698,In_2050);
and U892 (N_892,In_1592,In_717);
nor U893 (N_893,In_1512,In_1629);
nand U894 (N_894,In_878,In_1543);
nand U895 (N_895,In_339,In_1514);
nor U896 (N_896,In_2001,In_160);
xnor U897 (N_897,In_1584,In_1169);
xor U898 (N_898,In_1533,In_1091);
nand U899 (N_899,In_379,In_1771);
or U900 (N_900,In_1516,In_576);
or U901 (N_901,In_52,In_1524);
or U902 (N_902,In_612,In_179);
nor U903 (N_903,In_1695,In_2357);
or U904 (N_904,In_38,In_15);
or U905 (N_905,In_685,In_141);
or U906 (N_906,In_1362,In_659);
or U907 (N_907,In_2140,In_1984);
or U908 (N_908,In_1668,In_1319);
and U909 (N_909,In_1838,In_1585);
and U910 (N_910,In_709,In_773);
or U911 (N_911,In_116,In_516);
nand U912 (N_912,In_2440,In_49);
and U913 (N_913,In_1632,In_855);
nand U914 (N_914,In_231,In_2347);
and U915 (N_915,In_1268,In_1903);
nand U916 (N_916,In_358,In_2000);
nor U917 (N_917,In_1209,In_1053);
nor U918 (N_918,In_1150,In_605);
nand U919 (N_919,In_1657,In_886);
and U920 (N_920,In_488,In_1937);
and U921 (N_921,In_2203,In_1358);
nor U922 (N_922,In_1965,In_2225);
or U923 (N_923,In_346,In_1823);
nor U924 (N_924,In_2084,In_319);
or U925 (N_925,In_2235,In_968);
or U926 (N_926,In_1912,In_909);
or U927 (N_927,In_2138,In_846);
and U928 (N_928,In_1645,In_1722);
or U929 (N_929,In_536,In_1318);
or U930 (N_930,In_2204,In_166);
nand U931 (N_931,In_970,In_550);
nor U932 (N_932,In_983,In_1870);
and U933 (N_933,In_366,In_1784);
nand U934 (N_934,In_2206,In_2387);
nor U935 (N_935,In_545,In_217);
nand U936 (N_936,In_430,In_2314);
nor U937 (N_937,In_1738,In_2318);
nor U938 (N_938,In_2488,In_327);
or U939 (N_939,In_2199,In_961);
nor U940 (N_940,In_2258,In_222);
or U941 (N_941,In_2385,In_1845);
nand U942 (N_942,In_1038,In_2039);
nor U943 (N_943,In_1340,In_2157);
and U944 (N_944,In_1391,In_209);
or U945 (N_945,In_705,In_1875);
or U946 (N_946,In_378,In_1552);
nor U947 (N_947,In_1860,In_170);
and U948 (N_948,In_1421,In_1755);
nor U949 (N_949,In_2071,In_139);
or U950 (N_950,In_332,In_1992);
nand U951 (N_951,In_2047,In_1404);
nor U952 (N_952,In_656,In_1643);
nor U953 (N_953,In_199,In_2325);
xor U954 (N_954,In_693,In_2052);
xor U955 (N_955,In_1968,In_1790);
or U956 (N_956,In_766,In_175);
or U957 (N_957,In_334,In_1548);
nand U958 (N_958,In_159,In_439);
and U959 (N_959,In_1248,In_637);
and U960 (N_960,In_1171,In_1561);
nand U961 (N_961,In_1662,In_259);
nand U962 (N_962,In_76,In_1553);
nand U963 (N_963,In_386,In_1061);
nand U964 (N_964,In_2214,In_811);
or U965 (N_965,In_1944,In_978);
or U966 (N_966,In_817,In_156);
nor U967 (N_967,In_1974,In_387);
and U968 (N_968,In_476,In_1685);
or U969 (N_969,In_68,In_365);
nand U970 (N_970,In_588,In_349);
or U971 (N_971,In_2317,In_26);
and U972 (N_972,In_1529,In_123);
nor U973 (N_973,In_2446,In_1201);
and U974 (N_974,In_2341,In_2075);
nor U975 (N_975,In_2068,In_918);
xnor U976 (N_976,In_2465,In_907);
and U977 (N_977,In_638,In_1904);
nand U978 (N_978,In_1918,In_688);
and U979 (N_979,In_1166,In_616);
nand U980 (N_980,In_1420,In_1103);
nor U981 (N_981,In_1321,In_12);
or U982 (N_982,In_1993,In_85);
or U983 (N_983,In_1004,In_2045);
and U984 (N_984,In_1824,In_341);
and U985 (N_985,In_1375,In_556);
nand U986 (N_986,In_1241,In_972);
nand U987 (N_987,In_2348,In_2247);
or U988 (N_988,In_1962,In_1653);
nor U989 (N_989,In_1057,In_949);
or U990 (N_990,In_1465,In_84);
nand U991 (N_991,In_1374,In_1724);
nand U992 (N_992,In_1667,In_1780);
or U993 (N_993,In_393,In_226);
nand U994 (N_994,In_2378,In_752);
or U995 (N_995,In_848,In_252);
nor U996 (N_996,In_636,In_210);
nor U997 (N_997,In_2231,In_2218);
nor U998 (N_998,In_501,In_661);
nand U999 (N_999,In_1274,In_2131);
nand U1000 (N_1000,In_2101,In_203);
nor U1001 (N_1001,In_818,In_1583);
or U1002 (N_1002,In_1930,In_416);
and U1003 (N_1003,In_513,In_1842);
nand U1004 (N_1004,In_2249,In_1370);
xnor U1005 (N_1005,In_1905,In_2397);
and U1006 (N_1006,In_236,In_1987);
and U1007 (N_1007,In_193,In_645);
or U1008 (N_1008,In_1855,In_1218);
or U1009 (N_1009,In_2104,In_2366);
nor U1010 (N_1010,In_2274,In_2438);
or U1011 (N_1011,In_1538,In_1731);
nor U1012 (N_1012,In_412,In_2390);
nand U1013 (N_1013,In_2215,In_2360);
nor U1014 (N_1014,In_1849,In_155);
xor U1015 (N_1015,In_2044,In_1023);
and U1016 (N_1016,In_1044,In_407);
and U1017 (N_1017,In_864,In_485);
or U1018 (N_1018,In_887,In_570);
nand U1019 (N_1019,In_409,In_825);
nor U1020 (N_1020,In_799,In_2161);
or U1021 (N_1021,In_1648,In_2297);
nand U1022 (N_1022,In_804,In_2331);
nand U1023 (N_1023,In_939,In_63);
or U1024 (N_1024,In_2018,In_1211);
and U1025 (N_1025,In_2173,In_648);
nor U1026 (N_1026,In_384,In_1948);
or U1027 (N_1027,In_1452,In_1594);
nor U1028 (N_1028,In_1906,In_822);
nand U1029 (N_1029,In_59,In_2377);
and U1030 (N_1030,In_1325,In_161);
and U1031 (N_1031,In_353,In_1536);
and U1032 (N_1032,In_1107,In_2169);
and U1033 (N_1033,In_391,In_1982);
nor U1034 (N_1034,In_1873,In_1586);
and U1035 (N_1035,In_1735,In_1356);
nor U1036 (N_1036,In_1726,In_1801);
or U1037 (N_1037,In_801,In_1746);
or U1038 (N_1038,In_1240,In_2196);
and U1039 (N_1039,In_361,In_152);
nand U1040 (N_1040,In_1265,In_761);
and U1041 (N_1041,In_2351,In_1196);
or U1042 (N_1042,In_2113,In_1969);
nand U1043 (N_1043,In_2388,In_1158);
nand U1044 (N_1044,In_2135,In_2109);
nand U1045 (N_1045,In_951,In_455);
or U1046 (N_1046,In_1281,In_2430);
or U1047 (N_1047,In_1764,In_432);
or U1048 (N_1048,In_2491,In_1264);
xor U1049 (N_1049,In_1900,In_2256);
and U1050 (N_1050,In_2309,In_174);
nor U1051 (N_1051,In_1361,In_1947);
nand U1052 (N_1052,In_2208,In_178);
nand U1053 (N_1053,In_2210,In_1687);
xnor U1054 (N_1054,In_1922,In_181);
nand U1055 (N_1055,In_2012,In_2024);
nand U1056 (N_1056,In_1477,In_888);
nor U1057 (N_1057,In_823,In_915);
xor U1058 (N_1058,In_2240,In_623);
nand U1059 (N_1059,In_140,In_394);
xor U1060 (N_1060,In_500,In_2015);
xor U1061 (N_1061,In_1252,In_459);
or U1062 (N_1062,In_1130,In_1072);
and U1063 (N_1063,In_1376,In_373);
xor U1064 (N_1064,In_1711,In_806);
xor U1065 (N_1065,In_1637,In_687);
nand U1066 (N_1066,In_2151,In_910);
nor U1067 (N_1067,In_243,In_1846);
and U1068 (N_1068,In_98,In_1280);
xnor U1069 (N_1069,In_2143,In_1701);
and U1070 (N_1070,In_305,In_2327);
nand U1071 (N_1071,In_464,In_18);
and U1072 (N_1072,In_975,In_930);
nor U1073 (N_1073,In_457,In_562);
or U1074 (N_1074,In_730,In_1261);
or U1075 (N_1075,In_2286,In_609);
nand U1076 (N_1076,In_2251,In_2036);
nand U1077 (N_1077,In_1080,In_2472);
xor U1078 (N_1078,In_1534,In_557);
nor U1079 (N_1079,In_2028,In_2294);
and U1080 (N_1080,In_1923,In_798);
nand U1081 (N_1081,In_460,In_1730);
nand U1082 (N_1082,In_922,In_654);
nor U1083 (N_1083,In_2118,In_1620);
and U1084 (N_1084,In_608,In_1732);
nor U1085 (N_1085,In_2334,In_1704);
or U1086 (N_1086,In_1713,In_1170);
or U1087 (N_1087,In_81,In_2002);
and U1088 (N_1088,In_2246,In_664);
nand U1089 (N_1089,In_1581,In_520);
nand U1090 (N_1090,In_984,In_546);
nor U1091 (N_1091,In_2108,In_380);
xor U1092 (N_1092,In_1234,In_401);
nand U1093 (N_1093,In_2019,In_129);
and U1094 (N_1094,In_812,In_1636);
or U1095 (N_1095,In_919,In_755);
nand U1096 (N_1096,In_862,In_1627);
and U1097 (N_1097,In_1487,In_1896);
nor U1098 (N_1098,In_313,In_1547);
or U1099 (N_1099,In_1830,In_2046);
or U1100 (N_1100,In_1472,In_2410);
xnor U1101 (N_1101,In_1039,In_375);
or U1102 (N_1102,In_2396,In_1634);
xor U1103 (N_1103,In_2299,In_824);
nand U1104 (N_1104,In_1541,In_2457);
nor U1105 (N_1105,In_1763,In_2329);
nor U1106 (N_1106,In_299,In_517);
and U1107 (N_1107,In_221,In_1964);
and U1108 (N_1108,In_1164,In_1641);
nor U1109 (N_1109,In_1511,In_2486);
xor U1110 (N_1110,In_331,In_269);
nand U1111 (N_1111,In_995,In_1009);
or U1112 (N_1112,In_2174,In_2368);
and U1113 (N_1113,In_1415,In_352);
and U1114 (N_1114,In_1271,In_2065);
nor U1115 (N_1115,In_780,In_2226);
and U1116 (N_1116,In_2278,In_1925);
or U1117 (N_1117,In_725,In_866);
nand U1118 (N_1118,In_663,In_2337);
nor U1119 (N_1119,In_615,In_2282);
or U1120 (N_1120,In_1444,In_1260);
or U1121 (N_1121,In_2054,In_249);
and U1122 (N_1122,In_1943,In_431);
or U1123 (N_1123,In_614,In_979);
xor U1124 (N_1124,In_1455,In_2043);
or U1125 (N_1125,In_1146,In_73);
nor U1126 (N_1126,In_1491,In_673);
xnor U1127 (N_1127,In_1434,In_1983);
nand U1128 (N_1128,In_182,In_2281);
and U1129 (N_1129,In_2407,In_969);
and U1130 (N_1130,In_738,In_503);
nand U1131 (N_1131,In_999,In_1485);
and U1132 (N_1132,In_442,In_1871);
or U1133 (N_1133,In_2076,In_107);
xnor U1134 (N_1134,In_2395,In_2158);
nand U1135 (N_1135,In_573,In_257);
xor U1136 (N_1136,In_591,In_1884);
or U1137 (N_1137,In_2117,In_1412);
nor U1138 (N_1138,In_2217,In_395);
nor U1139 (N_1139,In_1500,In_372);
nor U1140 (N_1140,In_635,In_172);
nand U1141 (N_1141,In_1333,In_2489);
and U1142 (N_1142,In_1686,In_135);
xor U1143 (N_1143,In_1706,In_916);
or U1144 (N_1144,In_2125,In_815);
or U1145 (N_1145,In_1140,In_1141);
or U1146 (N_1146,In_1153,In_1249);
or U1147 (N_1147,In_985,In_1152);
nor U1148 (N_1148,In_694,In_735);
xnor U1149 (N_1149,In_700,In_847);
and U1150 (N_1150,In_1054,In_1279);
nand U1151 (N_1151,In_356,In_2007);
xnor U1152 (N_1152,In_1353,In_1436);
nand U1153 (N_1153,In_2490,In_2437);
nand U1154 (N_1154,In_1945,In_399);
and U1155 (N_1155,In_913,In_2098);
nand U1156 (N_1156,In_1034,In_1766);
and U1157 (N_1157,In_776,In_468);
nand U1158 (N_1158,In_2120,In_1431);
nor U1159 (N_1159,In_1427,In_1078);
nor U1160 (N_1160,In_1101,In_917);
nor U1161 (N_1161,In_1051,In_607);
nor U1162 (N_1162,In_1383,In_867);
and U1163 (N_1163,In_153,In_2060);
xnor U1164 (N_1164,In_1576,In_2298);
and U1165 (N_1165,In_689,In_843);
or U1166 (N_1166,In_302,In_1410);
nand U1167 (N_1167,In_1684,In_990);
or U1168 (N_1168,In_273,In_1688);
or U1169 (N_1169,In_2200,In_293);
nor U1170 (N_1170,In_2358,In_2216);
and U1171 (N_1171,In_400,In_813);
or U1172 (N_1172,In_1952,In_1225);
nand U1173 (N_1173,In_190,In_1368);
nor U1174 (N_1174,In_2456,In_1137);
xor U1175 (N_1175,In_223,In_2152);
and U1176 (N_1176,In_1214,In_1015);
or U1177 (N_1177,In_1200,In_1288);
nor U1178 (N_1178,In_2492,In_1811);
nor U1179 (N_1179,In_1762,In_102);
nand U1180 (N_1180,In_2150,In_1187);
or U1181 (N_1181,In_184,In_1312);
nor U1182 (N_1182,In_467,In_1094);
nor U1183 (N_1183,In_369,In_1409);
and U1184 (N_1184,In_2014,In_639);
xnor U1185 (N_1185,In_30,In_1921);
nand U1186 (N_1186,In_2029,In_2105);
nor U1187 (N_1187,In_1432,In_1832);
or U1188 (N_1188,In_1765,In_1026);
or U1189 (N_1189,In_2244,In_1269);
or U1190 (N_1190,In_2300,In_828);
or U1191 (N_1191,In_737,In_1475);
and U1192 (N_1192,In_397,In_1402);
and U1193 (N_1193,In_202,In_2400);
or U1194 (N_1194,In_543,In_2078);
xor U1195 (N_1195,In_767,In_2305);
nand U1196 (N_1196,In_247,In_2464);
and U1197 (N_1197,In_2096,In_2255);
or U1198 (N_1198,In_1159,In_2092);
or U1199 (N_1199,In_33,In_1647);
and U1200 (N_1200,In_2389,In_242);
nand U1201 (N_1201,In_2190,In_220);
nand U1202 (N_1202,In_1877,In_1869);
or U1203 (N_1203,In_1453,In_1188);
nor U1204 (N_1204,In_1242,In_2238);
and U1205 (N_1205,In_1497,In_952);
nor U1206 (N_1206,In_943,In_2480);
nand U1207 (N_1207,In_2301,In_881);
and U1208 (N_1208,In_796,In_602);
or U1209 (N_1209,In_2418,In_1076);
or U1210 (N_1210,In_841,In_1118);
nand U1211 (N_1211,In_2447,In_311);
nor U1212 (N_1212,In_989,In_2434);
nand U1213 (N_1213,In_1389,In_1959);
nor U1214 (N_1214,In_2003,In_1064);
nand U1215 (N_1215,In_2382,In_1330);
nor U1216 (N_1216,In_1357,In_1194);
or U1217 (N_1217,In_870,In_633);
nor U1218 (N_1218,In_1083,In_686);
nor U1219 (N_1219,In_420,In_1084);
and U1220 (N_1220,In_540,In_2094);
or U1221 (N_1221,In_1471,In_1272);
and U1222 (N_1222,In_1822,In_1530);
and U1223 (N_1223,In_740,In_1347);
or U1224 (N_1224,In_308,In_1963);
nand U1225 (N_1225,In_1161,In_277);
and U1226 (N_1226,In_2180,In_1825);
and U1227 (N_1227,In_396,In_564);
or U1228 (N_1228,In_2016,In_1523);
and U1229 (N_1229,In_1950,In_1881);
nor U1230 (N_1230,In_1723,In_1185);
and U1231 (N_1231,In_296,In_198);
or U1232 (N_1232,In_1237,In_849);
and U1233 (N_1233,In_115,In_1760);
or U1234 (N_1234,In_2025,In_1736);
nor U1235 (N_1235,In_1154,In_1624);
nor U1236 (N_1236,In_1829,In_1941);
and U1237 (N_1237,In_2345,In_446);
or U1238 (N_1238,In_224,In_675);
nor U1239 (N_1239,In_1395,In_122);
or U1240 (N_1240,In_1037,In_1997);
xnor U1241 (N_1241,In_2453,In_1422);
xnor U1242 (N_1242,In_465,In_1114);
nor U1243 (N_1243,In_1113,In_606);
xnor U1244 (N_1244,In_206,In_1371);
nand U1245 (N_1245,In_1029,In_511);
nand U1246 (N_1246,In_2144,In_2427);
nand U1247 (N_1247,In_1426,In_470);
nand U1248 (N_1248,In_1106,In_337);
and U1249 (N_1249,In_2379,In_1928);
and U1250 (N_1250,In_1141,In_1786);
nand U1251 (N_1251,In_630,In_2472);
or U1252 (N_1252,In_1973,In_1116);
and U1253 (N_1253,In_453,In_120);
nand U1254 (N_1254,In_286,In_1354);
or U1255 (N_1255,In_68,In_645);
xor U1256 (N_1256,In_1206,In_1591);
xnor U1257 (N_1257,In_687,In_2338);
and U1258 (N_1258,In_2036,In_2102);
nand U1259 (N_1259,In_1533,In_1631);
nor U1260 (N_1260,In_2000,In_1433);
xnor U1261 (N_1261,In_711,In_1629);
nand U1262 (N_1262,In_999,In_951);
and U1263 (N_1263,In_731,In_1953);
nor U1264 (N_1264,In_1439,In_222);
or U1265 (N_1265,In_2051,In_1796);
or U1266 (N_1266,In_390,In_380);
xor U1267 (N_1267,In_1041,In_1447);
and U1268 (N_1268,In_1876,In_456);
and U1269 (N_1269,In_992,In_1572);
nand U1270 (N_1270,In_487,In_1356);
nor U1271 (N_1271,In_2356,In_644);
and U1272 (N_1272,In_1296,In_2134);
or U1273 (N_1273,In_27,In_1927);
nor U1274 (N_1274,In_1023,In_871);
nor U1275 (N_1275,In_1159,In_975);
nor U1276 (N_1276,In_751,In_384);
nor U1277 (N_1277,In_1859,In_1254);
and U1278 (N_1278,In_2104,In_1326);
or U1279 (N_1279,In_991,In_2060);
or U1280 (N_1280,In_162,In_117);
nor U1281 (N_1281,In_638,In_697);
nor U1282 (N_1282,In_891,In_1496);
nor U1283 (N_1283,In_1298,In_857);
and U1284 (N_1284,In_2352,In_1441);
nand U1285 (N_1285,In_2068,In_2477);
xor U1286 (N_1286,In_2035,In_179);
nand U1287 (N_1287,In_1092,In_1315);
nand U1288 (N_1288,In_943,In_1098);
and U1289 (N_1289,In_628,In_1115);
xor U1290 (N_1290,In_852,In_2090);
nand U1291 (N_1291,In_661,In_743);
and U1292 (N_1292,In_774,In_1046);
nor U1293 (N_1293,In_2120,In_1890);
nor U1294 (N_1294,In_1930,In_152);
and U1295 (N_1295,In_1795,In_1999);
nor U1296 (N_1296,In_554,In_951);
and U1297 (N_1297,In_2149,In_2490);
nor U1298 (N_1298,In_147,In_521);
or U1299 (N_1299,In_1724,In_703);
or U1300 (N_1300,In_1306,In_584);
and U1301 (N_1301,In_2421,In_1817);
or U1302 (N_1302,In_2211,In_1189);
nor U1303 (N_1303,In_1489,In_2172);
nand U1304 (N_1304,In_176,In_2099);
nand U1305 (N_1305,In_749,In_577);
nor U1306 (N_1306,In_1594,In_1058);
or U1307 (N_1307,In_2474,In_664);
nor U1308 (N_1308,In_204,In_2293);
nand U1309 (N_1309,In_46,In_482);
or U1310 (N_1310,In_213,In_1483);
nor U1311 (N_1311,In_1072,In_8);
nand U1312 (N_1312,In_1622,In_469);
and U1313 (N_1313,In_2447,In_1246);
nand U1314 (N_1314,In_2429,In_2170);
nand U1315 (N_1315,In_1057,In_173);
and U1316 (N_1316,In_2059,In_788);
or U1317 (N_1317,In_1479,In_241);
nand U1318 (N_1318,In_612,In_1196);
nand U1319 (N_1319,In_2256,In_1405);
and U1320 (N_1320,In_1294,In_113);
and U1321 (N_1321,In_2465,In_1236);
or U1322 (N_1322,In_57,In_1127);
nor U1323 (N_1323,In_2294,In_524);
nand U1324 (N_1324,In_1328,In_1399);
or U1325 (N_1325,In_1854,In_1544);
nor U1326 (N_1326,In_598,In_1540);
or U1327 (N_1327,In_1658,In_1265);
nor U1328 (N_1328,In_956,In_1657);
nand U1329 (N_1329,In_2165,In_1147);
nor U1330 (N_1330,In_2208,In_960);
nand U1331 (N_1331,In_2384,In_60);
nor U1332 (N_1332,In_2012,In_337);
nor U1333 (N_1333,In_849,In_689);
nand U1334 (N_1334,In_2305,In_734);
and U1335 (N_1335,In_1681,In_1213);
nor U1336 (N_1336,In_1611,In_298);
and U1337 (N_1337,In_504,In_2483);
nand U1338 (N_1338,In_2207,In_1887);
and U1339 (N_1339,In_1148,In_1398);
and U1340 (N_1340,In_865,In_256);
and U1341 (N_1341,In_2102,In_1328);
xnor U1342 (N_1342,In_223,In_150);
or U1343 (N_1343,In_1325,In_1733);
nand U1344 (N_1344,In_856,In_49);
and U1345 (N_1345,In_1614,In_176);
or U1346 (N_1346,In_520,In_583);
or U1347 (N_1347,In_472,In_936);
nand U1348 (N_1348,In_2302,In_624);
xor U1349 (N_1349,In_1804,In_2127);
nand U1350 (N_1350,In_2378,In_2302);
nor U1351 (N_1351,In_1093,In_245);
nor U1352 (N_1352,In_668,In_2447);
nor U1353 (N_1353,In_944,In_251);
or U1354 (N_1354,In_728,In_1856);
nand U1355 (N_1355,In_594,In_1784);
nor U1356 (N_1356,In_1664,In_977);
nand U1357 (N_1357,In_921,In_1753);
nand U1358 (N_1358,In_1262,In_1342);
or U1359 (N_1359,In_0,In_837);
and U1360 (N_1360,In_284,In_493);
nor U1361 (N_1361,In_2045,In_1428);
nor U1362 (N_1362,In_1321,In_1402);
and U1363 (N_1363,In_332,In_1792);
nor U1364 (N_1364,In_1604,In_1431);
nor U1365 (N_1365,In_1257,In_1943);
nor U1366 (N_1366,In_2013,In_100);
xor U1367 (N_1367,In_392,In_2068);
or U1368 (N_1368,In_662,In_2262);
nor U1369 (N_1369,In_1799,In_2241);
nor U1370 (N_1370,In_1510,In_2334);
and U1371 (N_1371,In_1004,In_1737);
and U1372 (N_1372,In_1759,In_1825);
nand U1373 (N_1373,In_2433,In_1261);
or U1374 (N_1374,In_657,In_532);
or U1375 (N_1375,In_898,In_2017);
and U1376 (N_1376,In_1849,In_796);
or U1377 (N_1377,In_1522,In_1440);
or U1378 (N_1378,In_2199,In_780);
and U1379 (N_1379,In_2467,In_2430);
xnor U1380 (N_1380,In_1520,In_971);
nor U1381 (N_1381,In_1763,In_566);
and U1382 (N_1382,In_754,In_1777);
and U1383 (N_1383,In_1823,In_775);
nor U1384 (N_1384,In_2368,In_227);
nand U1385 (N_1385,In_1982,In_1203);
and U1386 (N_1386,In_665,In_417);
nand U1387 (N_1387,In_1569,In_158);
or U1388 (N_1388,In_1990,In_448);
and U1389 (N_1389,In_798,In_78);
or U1390 (N_1390,In_1080,In_1588);
and U1391 (N_1391,In_1765,In_406);
xnor U1392 (N_1392,In_1565,In_2289);
and U1393 (N_1393,In_50,In_2123);
xnor U1394 (N_1394,In_1087,In_2344);
nor U1395 (N_1395,In_2253,In_2061);
and U1396 (N_1396,In_426,In_2);
xnor U1397 (N_1397,In_2203,In_1193);
or U1398 (N_1398,In_1118,In_111);
and U1399 (N_1399,In_581,In_1749);
nand U1400 (N_1400,In_259,In_445);
or U1401 (N_1401,In_126,In_1450);
or U1402 (N_1402,In_1432,In_531);
nor U1403 (N_1403,In_121,In_316);
xnor U1404 (N_1404,In_912,In_1084);
nor U1405 (N_1405,In_1727,In_638);
or U1406 (N_1406,In_1901,In_506);
nand U1407 (N_1407,In_1630,In_248);
nor U1408 (N_1408,In_947,In_208);
or U1409 (N_1409,In_1787,In_1208);
or U1410 (N_1410,In_1449,In_1656);
xnor U1411 (N_1411,In_53,In_2020);
nor U1412 (N_1412,In_2336,In_1666);
xnor U1413 (N_1413,In_1699,In_371);
nand U1414 (N_1414,In_2316,In_1762);
and U1415 (N_1415,In_1171,In_1651);
and U1416 (N_1416,In_2192,In_1200);
nor U1417 (N_1417,In_643,In_1272);
nand U1418 (N_1418,In_2131,In_314);
nand U1419 (N_1419,In_522,In_769);
nand U1420 (N_1420,In_685,In_2421);
xnor U1421 (N_1421,In_1337,In_2112);
or U1422 (N_1422,In_825,In_768);
nand U1423 (N_1423,In_93,In_896);
xor U1424 (N_1424,In_1933,In_1009);
nor U1425 (N_1425,In_1394,In_81);
nor U1426 (N_1426,In_849,In_29);
nor U1427 (N_1427,In_1139,In_2215);
and U1428 (N_1428,In_16,In_1529);
and U1429 (N_1429,In_1068,In_2493);
nor U1430 (N_1430,In_1313,In_1456);
and U1431 (N_1431,In_1787,In_1041);
nor U1432 (N_1432,In_1831,In_964);
and U1433 (N_1433,In_909,In_2248);
nor U1434 (N_1434,In_1208,In_647);
nand U1435 (N_1435,In_2428,In_79);
or U1436 (N_1436,In_1526,In_2333);
or U1437 (N_1437,In_2341,In_2066);
nor U1438 (N_1438,In_2137,In_1351);
nor U1439 (N_1439,In_1523,In_945);
and U1440 (N_1440,In_2373,In_2085);
nand U1441 (N_1441,In_6,In_1147);
or U1442 (N_1442,In_168,In_1088);
nor U1443 (N_1443,In_104,In_1985);
nor U1444 (N_1444,In_326,In_179);
nand U1445 (N_1445,In_1377,In_1832);
or U1446 (N_1446,In_992,In_2243);
or U1447 (N_1447,In_363,In_694);
or U1448 (N_1448,In_1792,In_2406);
nor U1449 (N_1449,In_1466,In_54);
xor U1450 (N_1450,In_217,In_2062);
nand U1451 (N_1451,In_320,In_1748);
nand U1452 (N_1452,In_353,In_510);
or U1453 (N_1453,In_1009,In_1306);
or U1454 (N_1454,In_2342,In_1782);
or U1455 (N_1455,In_1962,In_1419);
nor U1456 (N_1456,In_864,In_2230);
and U1457 (N_1457,In_1464,In_1666);
or U1458 (N_1458,In_1887,In_234);
xor U1459 (N_1459,In_590,In_734);
or U1460 (N_1460,In_2386,In_480);
and U1461 (N_1461,In_2182,In_553);
nor U1462 (N_1462,In_1906,In_2126);
nor U1463 (N_1463,In_1712,In_2017);
xor U1464 (N_1464,In_294,In_2259);
and U1465 (N_1465,In_1213,In_1789);
or U1466 (N_1466,In_185,In_2458);
and U1467 (N_1467,In_1411,In_999);
or U1468 (N_1468,In_1980,In_1087);
nand U1469 (N_1469,In_326,In_855);
or U1470 (N_1470,In_627,In_2351);
or U1471 (N_1471,In_2375,In_604);
nor U1472 (N_1472,In_727,In_1865);
nand U1473 (N_1473,In_421,In_1727);
xnor U1474 (N_1474,In_1364,In_813);
or U1475 (N_1475,In_681,In_2262);
nor U1476 (N_1476,In_1456,In_1690);
xor U1477 (N_1477,In_2206,In_735);
and U1478 (N_1478,In_2090,In_2372);
nor U1479 (N_1479,In_358,In_925);
or U1480 (N_1480,In_818,In_1527);
or U1481 (N_1481,In_1954,In_231);
and U1482 (N_1482,In_572,In_54);
and U1483 (N_1483,In_619,In_537);
nor U1484 (N_1484,In_2293,In_919);
or U1485 (N_1485,In_1630,In_1192);
and U1486 (N_1486,In_951,In_1129);
nor U1487 (N_1487,In_2232,In_378);
and U1488 (N_1488,In_454,In_927);
nor U1489 (N_1489,In_1950,In_2165);
xnor U1490 (N_1490,In_650,In_915);
or U1491 (N_1491,In_1469,In_954);
nand U1492 (N_1492,In_525,In_490);
nor U1493 (N_1493,In_1534,In_964);
or U1494 (N_1494,In_686,In_1983);
nand U1495 (N_1495,In_142,In_877);
or U1496 (N_1496,In_1316,In_288);
or U1497 (N_1497,In_1180,In_2305);
nor U1498 (N_1498,In_257,In_1056);
xor U1499 (N_1499,In_2004,In_507);
nor U1500 (N_1500,In_101,In_1929);
nor U1501 (N_1501,In_1239,In_747);
nand U1502 (N_1502,In_2110,In_2227);
and U1503 (N_1503,In_1103,In_131);
nor U1504 (N_1504,In_697,In_806);
or U1505 (N_1505,In_1415,In_2237);
nand U1506 (N_1506,In_800,In_1501);
nor U1507 (N_1507,In_2343,In_1816);
or U1508 (N_1508,In_2489,In_682);
or U1509 (N_1509,In_1812,In_449);
nor U1510 (N_1510,In_1316,In_1084);
nand U1511 (N_1511,In_1886,In_1035);
or U1512 (N_1512,In_693,In_286);
or U1513 (N_1513,In_541,In_1629);
nor U1514 (N_1514,In_250,In_1932);
nand U1515 (N_1515,In_2188,In_130);
nand U1516 (N_1516,In_49,In_298);
nand U1517 (N_1517,In_52,In_2343);
nor U1518 (N_1518,In_2004,In_548);
and U1519 (N_1519,In_1024,In_2496);
nor U1520 (N_1520,In_1587,In_2195);
nand U1521 (N_1521,In_1868,In_853);
nor U1522 (N_1522,In_1713,In_2178);
and U1523 (N_1523,In_453,In_257);
or U1524 (N_1524,In_61,In_1861);
or U1525 (N_1525,In_2422,In_1969);
xor U1526 (N_1526,In_2392,In_1498);
or U1527 (N_1527,In_412,In_910);
and U1528 (N_1528,In_460,In_1939);
and U1529 (N_1529,In_39,In_1095);
or U1530 (N_1530,In_512,In_1701);
nor U1531 (N_1531,In_937,In_2291);
nand U1532 (N_1532,In_994,In_1964);
or U1533 (N_1533,In_2324,In_341);
and U1534 (N_1534,In_1229,In_1498);
and U1535 (N_1535,In_282,In_1452);
and U1536 (N_1536,In_1435,In_1794);
nor U1537 (N_1537,In_666,In_484);
and U1538 (N_1538,In_2385,In_2271);
or U1539 (N_1539,In_1870,In_219);
and U1540 (N_1540,In_1767,In_2300);
or U1541 (N_1541,In_1297,In_2264);
nor U1542 (N_1542,In_1876,In_761);
nand U1543 (N_1543,In_330,In_2144);
xor U1544 (N_1544,In_826,In_959);
or U1545 (N_1545,In_2320,In_2433);
nand U1546 (N_1546,In_2169,In_51);
nand U1547 (N_1547,In_694,In_2318);
nor U1548 (N_1548,In_1121,In_1139);
and U1549 (N_1549,In_1327,In_1187);
and U1550 (N_1550,In_1828,In_2381);
or U1551 (N_1551,In_834,In_1902);
or U1552 (N_1552,In_1147,In_1338);
or U1553 (N_1553,In_1802,In_578);
or U1554 (N_1554,In_1184,In_1447);
or U1555 (N_1555,In_2035,In_1188);
nor U1556 (N_1556,In_1091,In_957);
or U1557 (N_1557,In_1426,In_1634);
nand U1558 (N_1558,In_26,In_2360);
and U1559 (N_1559,In_21,In_1892);
nor U1560 (N_1560,In_939,In_859);
nand U1561 (N_1561,In_2260,In_832);
and U1562 (N_1562,In_1097,In_425);
nor U1563 (N_1563,In_1577,In_1002);
and U1564 (N_1564,In_1517,In_1295);
xor U1565 (N_1565,In_32,In_483);
xnor U1566 (N_1566,In_1301,In_34);
nor U1567 (N_1567,In_1540,In_2317);
nand U1568 (N_1568,In_2317,In_619);
nor U1569 (N_1569,In_2063,In_1488);
or U1570 (N_1570,In_1814,In_898);
nand U1571 (N_1571,In_1351,In_1962);
and U1572 (N_1572,In_2173,In_1118);
nand U1573 (N_1573,In_1678,In_725);
nand U1574 (N_1574,In_338,In_1947);
nand U1575 (N_1575,In_1594,In_1714);
and U1576 (N_1576,In_597,In_2318);
and U1577 (N_1577,In_152,In_118);
or U1578 (N_1578,In_1867,In_1669);
or U1579 (N_1579,In_1888,In_2424);
nand U1580 (N_1580,In_1189,In_1516);
nand U1581 (N_1581,In_1684,In_1359);
or U1582 (N_1582,In_1633,In_157);
and U1583 (N_1583,In_2247,In_2249);
and U1584 (N_1584,In_615,In_1470);
nor U1585 (N_1585,In_2049,In_1709);
nand U1586 (N_1586,In_1678,In_900);
or U1587 (N_1587,In_780,In_1421);
nor U1588 (N_1588,In_254,In_1952);
and U1589 (N_1589,In_2051,In_2295);
nor U1590 (N_1590,In_982,In_241);
nor U1591 (N_1591,In_905,In_1960);
xor U1592 (N_1592,In_2145,In_1588);
or U1593 (N_1593,In_863,In_1784);
nand U1594 (N_1594,In_603,In_1079);
or U1595 (N_1595,In_2342,In_386);
or U1596 (N_1596,In_1739,In_2381);
or U1597 (N_1597,In_596,In_440);
and U1598 (N_1598,In_172,In_247);
nor U1599 (N_1599,In_735,In_1852);
nand U1600 (N_1600,In_1307,In_1333);
and U1601 (N_1601,In_571,In_693);
nand U1602 (N_1602,In_362,In_2);
nand U1603 (N_1603,In_2232,In_1683);
nor U1604 (N_1604,In_1784,In_389);
xnor U1605 (N_1605,In_2464,In_640);
nor U1606 (N_1606,In_1707,In_1919);
nor U1607 (N_1607,In_408,In_2176);
or U1608 (N_1608,In_1622,In_568);
nand U1609 (N_1609,In_2114,In_40);
or U1610 (N_1610,In_1743,In_1111);
or U1611 (N_1611,In_1968,In_639);
and U1612 (N_1612,In_598,In_182);
and U1613 (N_1613,In_202,In_1443);
and U1614 (N_1614,In_1624,In_1508);
nand U1615 (N_1615,In_229,In_192);
nor U1616 (N_1616,In_1911,In_1208);
or U1617 (N_1617,In_2331,In_2064);
or U1618 (N_1618,In_919,In_1977);
nor U1619 (N_1619,In_1841,In_1371);
nand U1620 (N_1620,In_286,In_94);
nor U1621 (N_1621,In_1537,In_725);
nor U1622 (N_1622,In_1656,In_2411);
or U1623 (N_1623,In_2190,In_1422);
and U1624 (N_1624,In_2214,In_1797);
and U1625 (N_1625,In_410,In_2249);
or U1626 (N_1626,In_1838,In_1828);
nand U1627 (N_1627,In_2240,In_1175);
and U1628 (N_1628,In_1547,In_878);
nand U1629 (N_1629,In_1371,In_1067);
or U1630 (N_1630,In_204,In_492);
nor U1631 (N_1631,In_948,In_172);
nand U1632 (N_1632,In_2212,In_2249);
nor U1633 (N_1633,In_1871,In_506);
nor U1634 (N_1634,In_2299,In_18);
nor U1635 (N_1635,In_146,In_899);
nor U1636 (N_1636,In_1389,In_1589);
nor U1637 (N_1637,In_686,In_1653);
and U1638 (N_1638,In_1682,In_127);
xnor U1639 (N_1639,In_526,In_1887);
and U1640 (N_1640,In_905,In_223);
xnor U1641 (N_1641,In_1025,In_786);
or U1642 (N_1642,In_547,In_2416);
nand U1643 (N_1643,In_971,In_829);
and U1644 (N_1644,In_1599,In_382);
nor U1645 (N_1645,In_1563,In_197);
nor U1646 (N_1646,In_1317,In_955);
nand U1647 (N_1647,In_722,In_563);
xor U1648 (N_1648,In_435,In_2113);
xnor U1649 (N_1649,In_1882,In_1724);
and U1650 (N_1650,In_1229,In_1915);
nand U1651 (N_1651,In_2012,In_2232);
nand U1652 (N_1652,In_677,In_271);
nor U1653 (N_1653,In_1262,In_2221);
or U1654 (N_1654,In_1588,In_299);
nand U1655 (N_1655,In_2201,In_2468);
nand U1656 (N_1656,In_743,In_40);
xnor U1657 (N_1657,In_1092,In_1739);
and U1658 (N_1658,In_1930,In_2010);
and U1659 (N_1659,In_580,In_1940);
nor U1660 (N_1660,In_2152,In_1521);
and U1661 (N_1661,In_1126,In_140);
nor U1662 (N_1662,In_1667,In_1790);
or U1663 (N_1663,In_1504,In_1502);
nand U1664 (N_1664,In_321,In_1190);
and U1665 (N_1665,In_2100,In_1035);
nand U1666 (N_1666,In_1039,In_829);
and U1667 (N_1667,In_717,In_2484);
or U1668 (N_1668,In_2447,In_1686);
and U1669 (N_1669,In_2353,In_1240);
nand U1670 (N_1670,In_1065,In_1726);
nand U1671 (N_1671,In_2018,In_250);
or U1672 (N_1672,In_609,In_1626);
and U1673 (N_1673,In_14,In_445);
nand U1674 (N_1674,In_1855,In_1538);
nand U1675 (N_1675,In_536,In_146);
nor U1676 (N_1676,In_537,In_2333);
nor U1677 (N_1677,In_1249,In_65);
or U1678 (N_1678,In_1777,In_790);
or U1679 (N_1679,In_1596,In_587);
and U1680 (N_1680,In_139,In_1531);
and U1681 (N_1681,In_80,In_1885);
nor U1682 (N_1682,In_2103,In_1010);
nor U1683 (N_1683,In_989,In_2014);
xnor U1684 (N_1684,In_2375,In_1107);
nor U1685 (N_1685,In_1959,In_926);
or U1686 (N_1686,In_290,In_1161);
and U1687 (N_1687,In_2448,In_1098);
or U1688 (N_1688,In_1294,In_1055);
or U1689 (N_1689,In_610,In_2135);
or U1690 (N_1690,In_1903,In_1981);
xor U1691 (N_1691,In_2466,In_928);
nor U1692 (N_1692,In_1095,In_2047);
and U1693 (N_1693,In_2147,In_771);
nand U1694 (N_1694,In_2478,In_1861);
nand U1695 (N_1695,In_1266,In_545);
and U1696 (N_1696,In_2149,In_246);
nor U1697 (N_1697,In_1690,In_1524);
nor U1698 (N_1698,In_1559,In_2484);
nor U1699 (N_1699,In_2133,In_682);
or U1700 (N_1700,In_1205,In_1560);
and U1701 (N_1701,In_2295,In_195);
nand U1702 (N_1702,In_1080,In_2299);
nor U1703 (N_1703,In_184,In_1478);
nand U1704 (N_1704,In_769,In_1751);
and U1705 (N_1705,In_1848,In_1262);
nor U1706 (N_1706,In_616,In_2285);
nand U1707 (N_1707,In_1765,In_1784);
xnor U1708 (N_1708,In_1246,In_1302);
nand U1709 (N_1709,In_1998,In_15);
and U1710 (N_1710,In_1640,In_2441);
nor U1711 (N_1711,In_1959,In_2047);
and U1712 (N_1712,In_2037,In_523);
and U1713 (N_1713,In_2152,In_879);
xnor U1714 (N_1714,In_1088,In_1236);
and U1715 (N_1715,In_757,In_2483);
nand U1716 (N_1716,In_1108,In_553);
and U1717 (N_1717,In_2287,In_1934);
nor U1718 (N_1718,In_993,In_31);
or U1719 (N_1719,In_281,In_1632);
xor U1720 (N_1720,In_1356,In_322);
nor U1721 (N_1721,In_1053,In_349);
or U1722 (N_1722,In_1601,In_1242);
nor U1723 (N_1723,In_1595,In_1874);
or U1724 (N_1724,In_255,In_138);
nor U1725 (N_1725,In_2063,In_810);
or U1726 (N_1726,In_949,In_680);
nor U1727 (N_1727,In_1592,In_1699);
nand U1728 (N_1728,In_982,In_23);
nand U1729 (N_1729,In_696,In_503);
nand U1730 (N_1730,In_2307,In_803);
nor U1731 (N_1731,In_445,In_397);
and U1732 (N_1732,In_1159,In_1944);
xor U1733 (N_1733,In_1644,In_2402);
nor U1734 (N_1734,In_1648,In_1415);
xnor U1735 (N_1735,In_1678,In_1135);
nand U1736 (N_1736,In_287,In_162);
nand U1737 (N_1737,In_1088,In_626);
nor U1738 (N_1738,In_1461,In_957);
or U1739 (N_1739,In_174,In_1896);
xnor U1740 (N_1740,In_993,In_298);
nand U1741 (N_1741,In_1934,In_2084);
xnor U1742 (N_1742,In_2426,In_713);
nand U1743 (N_1743,In_1629,In_1318);
nor U1744 (N_1744,In_1608,In_1932);
or U1745 (N_1745,In_157,In_1246);
nor U1746 (N_1746,In_1681,In_434);
nand U1747 (N_1747,In_1820,In_1483);
nor U1748 (N_1748,In_1415,In_1219);
or U1749 (N_1749,In_155,In_1413);
nand U1750 (N_1750,In_582,In_2483);
and U1751 (N_1751,In_1831,In_1006);
or U1752 (N_1752,In_286,In_1915);
or U1753 (N_1753,In_1611,In_1561);
or U1754 (N_1754,In_2156,In_2031);
and U1755 (N_1755,In_2238,In_1799);
nand U1756 (N_1756,In_1286,In_1427);
nor U1757 (N_1757,In_1310,In_2405);
or U1758 (N_1758,In_2368,In_16);
nand U1759 (N_1759,In_1988,In_1388);
and U1760 (N_1760,In_2345,In_1335);
and U1761 (N_1761,In_114,In_2268);
or U1762 (N_1762,In_2481,In_13);
xor U1763 (N_1763,In_61,In_1019);
and U1764 (N_1764,In_1925,In_500);
and U1765 (N_1765,In_986,In_741);
and U1766 (N_1766,In_2455,In_14);
nor U1767 (N_1767,In_850,In_2186);
and U1768 (N_1768,In_775,In_1904);
nor U1769 (N_1769,In_155,In_645);
and U1770 (N_1770,In_2117,In_1118);
or U1771 (N_1771,In_1908,In_1726);
and U1772 (N_1772,In_30,In_300);
or U1773 (N_1773,In_1400,In_906);
xor U1774 (N_1774,In_1885,In_226);
nor U1775 (N_1775,In_208,In_1295);
and U1776 (N_1776,In_294,In_2256);
nand U1777 (N_1777,In_2024,In_1777);
xor U1778 (N_1778,In_2213,In_1825);
nor U1779 (N_1779,In_726,In_1199);
and U1780 (N_1780,In_2420,In_2466);
nand U1781 (N_1781,In_2268,In_29);
nand U1782 (N_1782,In_1446,In_1268);
nand U1783 (N_1783,In_367,In_477);
xor U1784 (N_1784,In_424,In_2280);
nor U1785 (N_1785,In_2479,In_2323);
nand U1786 (N_1786,In_844,In_2230);
nor U1787 (N_1787,In_1528,In_947);
nand U1788 (N_1788,In_1258,In_2241);
or U1789 (N_1789,In_659,In_1202);
nor U1790 (N_1790,In_1407,In_713);
nor U1791 (N_1791,In_2199,In_838);
nand U1792 (N_1792,In_1483,In_883);
or U1793 (N_1793,In_2082,In_1341);
and U1794 (N_1794,In_822,In_799);
and U1795 (N_1795,In_2072,In_309);
and U1796 (N_1796,In_2064,In_1369);
nor U1797 (N_1797,In_1711,In_1350);
and U1798 (N_1798,In_869,In_1267);
nor U1799 (N_1799,In_1708,In_626);
and U1800 (N_1800,In_1017,In_1236);
and U1801 (N_1801,In_652,In_110);
and U1802 (N_1802,In_334,In_1090);
and U1803 (N_1803,In_310,In_1549);
xor U1804 (N_1804,In_687,In_429);
and U1805 (N_1805,In_1380,In_1952);
nand U1806 (N_1806,In_1259,In_1938);
nand U1807 (N_1807,In_479,In_2040);
nand U1808 (N_1808,In_2207,In_230);
nand U1809 (N_1809,In_1445,In_537);
nor U1810 (N_1810,In_1343,In_1984);
nand U1811 (N_1811,In_234,In_1584);
and U1812 (N_1812,In_391,In_1036);
nor U1813 (N_1813,In_1369,In_1577);
nor U1814 (N_1814,In_120,In_988);
and U1815 (N_1815,In_125,In_2399);
and U1816 (N_1816,In_1320,In_345);
nand U1817 (N_1817,In_802,In_1771);
and U1818 (N_1818,In_426,In_1991);
or U1819 (N_1819,In_2387,In_95);
nor U1820 (N_1820,In_890,In_1779);
nor U1821 (N_1821,In_1846,In_1162);
or U1822 (N_1822,In_1231,In_1952);
and U1823 (N_1823,In_1562,In_340);
nand U1824 (N_1824,In_381,In_51);
nor U1825 (N_1825,In_167,In_2413);
nor U1826 (N_1826,In_875,In_2258);
nor U1827 (N_1827,In_710,In_1052);
or U1828 (N_1828,In_1596,In_2098);
xnor U1829 (N_1829,In_40,In_2014);
or U1830 (N_1830,In_144,In_1786);
nor U1831 (N_1831,In_508,In_813);
and U1832 (N_1832,In_1727,In_1069);
xor U1833 (N_1833,In_1406,In_239);
nor U1834 (N_1834,In_2339,In_945);
nor U1835 (N_1835,In_165,In_431);
nand U1836 (N_1836,In_2150,In_1997);
nor U1837 (N_1837,In_1521,In_221);
or U1838 (N_1838,In_139,In_2083);
or U1839 (N_1839,In_1955,In_2391);
nor U1840 (N_1840,In_251,In_930);
xnor U1841 (N_1841,In_871,In_349);
xor U1842 (N_1842,In_2058,In_462);
and U1843 (N_1843,In_1376,In_1496);
or U1844 (N_1844,In_1949,In_1308);
nand U1845 (N_1845,In_915,In_1519);
nor U1846 (N_1846,In_2072,In_2484);
or U1847 (N_1847,In_2334,In_212);
and U1848 (N_1848,In_1242,In_664);
nand U1849 (N_1849,In_1273,In_2223);
nor U1850 (N_1850,In_2473,In_1445);
and U1851 (N_1851,In_1263,In_2454);
and U1852 (N_1852,In_2211,In_2235);
or U1853 (N_1853,In_362,In_90);
nand U1854 (N_1854,In_1866,In_13);
and U1855 (N_1855,In_274,In_2085);
xnor U1856 (N_1856,In_889,In_583);
and U1857 (N_1857,In_1111,In_369);
and U1858 (N_1858,In_2364,In_547);
nand U1859 (N_1859,In_257,In_2077);
nand U1860 (N_1860,In_681,In_2285);
and U1861 (N_1861,In_1034,In_1251);
or U1862 (N_1862,In_983,In_2034);
or U1863 (N_1863,In_2393,In_1485);
nor U1864 (N_1864,In_2402,In_828);
xor U1865 (N_1865,In_2372,In_1760);
or U1866 (N_1866,In_1614,In_1109);
nor U1867 (N_1867,In_857,In_1365);
and U1868 (N_1868,In_588,In_492);
nand U1869 (N_1869,In_1806,In_488);
xor U1870 (N_1870,In_2464,In_948);
nand U1871 (N_1871,In_1184,In_1967);
and U1872 (N_1872,In_1559,In_1396);
and U1873 (N_1873,In_1168,In_362);
and U1874 (N_1874,In_2435,In_1139);
or U1875 (N_1875,In_1155,In_670);
nor U1876 (N_1876,In_1650,In_1439);
xnor U1877 (N_1877,In_2485,In_203);
nand U1878 (N_1878,In_556,In_786);
nand U1879 (N_1879,In_200,In_891);
nor U1880 (N_1880,In_394,In_1779);
nor U1881 (N_1881,In_835,In_1426);
and U1882 (N_1882,In_333,In_1297);
nor U1883 (N_1883,In_673,In_351);
nor U1884 (N_1884,In_1279,In_70);
nand U1885 (N_1885,In_454,In_1164);
and U1886 (N_1886,In_853,In_2418);
nand U1887 (N_1887,In_2164,In_1336);
nor U1888 (N_1888,In_2442,In_1613);
nand U1889 (N_1889,In_2243,In_233);
xnor U1890 (N_1890,In_1533,In_1112);
xor U1891 (N_1891,In_1378,In_1878);
or U1892 (N_1892,In_2471,In_2273);
nor U1893 (N_1893,In_336,In_760);
or U1894 (N_1894,In_2497,In_433);
or U1895 (N_1895,In_148,In_1916);
nor U1896 (N_1896,In_695,In_2431);
or U1897 (N_1897,In_755,In_504);
xor U1898 (N_1898,In_1996,In_1523);
nor U1899 (N_1899,In_590,In_1357);
nor U1900 (N_1900,In_123,In_1940);
nor U1901 (N_1901,In_969,In_636);
or U1902 (N_1902,In_245,In_1949);
and U1903 (N_1903,In_655,In_2040);
nand U1904 (N_1904,In_1344,In_1822);
or U1905 (N_1905,In_2174,In_2276);
and U1906 (N_1906,In_252,In_754);
and U1907 (N_1907,In_2373,In_2039);
nand U1908 (N_1908,In_594,In_352);
and U1909 (N_1909,In_331,In_1678);
or U1910 (N_1910,In_943,In_1022);
nand U1911 (N_1911,In_1363,In_1466);
nor U1912 (N_1912,In_2276,In_1754);
and U1913 (N_1913,In_1171,In_764);
or U1914 (N_1914,In_1739,In_1655);
and U1915 (N_1915,In_1079,In_403);
nand U1916 (N_1916,In_2377,In_191);
or U1917 (N_1917,In_557,In_1819);
or U1918 (N_1918,In_860,In_1654);
or U1919 (N_1919,In_675,In_38);
and U1920 (N_1920,In_2188,In_1474);
and U1921 (N_1921,In_1576,In_596);
xnor U1922 (N_1922,In_1990,In_346);
xnor U1923 (N_1923,In_850,In_480);
or U1924 (N_1924,In_2018,In_1574);
and U1925 (N_1925,In_141,In_2334);
nand U1926 (N_1926,In_1188,In_1796);
nand U1927 (N_1927,In_1967,In_1979);
nand U1928 (N_1928,In_2343,In_477);
nor U1929 (N_1929,In_2381,In_1862);
nand U1930 (N_1930,In_1618,In_1307);
nor U1931 (N_1931,In_1184,In_1950);
or U1932 (N_1932,In_1788,In_569);
or U1933 (N_1933,In_977,In_2464);
nand U1934 (N_1934,In_2405,In_1965);
nand U1935 (N_1935,In_1042,In_848);
and U1936 (N_1936,In_1681,In_2218);
and U1937 (N_1937,In_60,In_2119);
nand U1938 (N_1938,In_1574,In_815);
and U1939 (N_1939,In_324,In_2096);
nor U1940 (N_1940,In_1432,In_1010);
and U1941 (N_1941,In_2319,In_1763);
nor U1942 (N_1942,In_2079,In_1929);
nor U1943 (N_1943,In_158,In_597);
nand U1944 (N_1944,In_2477,In_1213);
and U1945 (N_1945,In_752,In_1940);
nor U1946 (N_1946,In_248,In_1921);
and U1947 (N_1947,In_827,In_1352);
nand U1948 (N_1948,In_121,In_1368);
or U1949 (N_1949,In_682,In_1673);
nand U1950 (N_1950,In_1231,In_1782);
or U1951 (N_1951,In_1686,In_2113);
or U1952 (N_1952,In_531,In_1649);
xnor U1953 (N_1953,In_2235,In_21);
and U1954 (N_1954,In_2105,In_456);
and U1955 (N_1955,In_2497,In_1781);
and U1956 (N_1956,In_2359,In_1862);
or U1957 (N_1957,In_16,In_2340);
nor U1958 (N_1958,In_1449,In_571);
nor U1959 (N_1959,In_1796,In_1374);
nand U1960 (N_1960,In_747,In_1448);
nor U1961 (N_1961,In_362,In_1988);
and U1962 (N_1962,In_474,In_984);
and U1963 (N_1963,In_1815,In_471);
or U1964 (N_1964,In_440,In_1748);
nand U1965 (N_1965,In_1207,In_1448);
nor U1966 (N_1966,In_1980,In_761);
nor U1967 (N_1967,In_1044,In_640);
nand U1968 (N_1968,In_2251,In_2247);
and U1969 (N_1969,In_397,In_1617);
and U1970 (N_1970,In_725,In_1463);
nand U1971 (N_1971,In_426,In_1741);
or U1972 (N_1972,In_1752,In_1083);
and U1973 (N_1973,In_369,In_1663);
or U1974 (N_1974,In_1107,In_239);
nand U1975 (N_1975,In_2279,In_1204);
nor U1976 (N_1976,In_1687,In_564);
xor U1977 (N_1977,In_2469,In_297);
xnor U1978 (N_1978,In_114,In_1687);
and U1979 (N_1979,In_708,In_1841);
nor U1980 (N_1980,In_1855,In_65);
and U1981 (N_1981,In_1005,In_1354);
or U1982 (N_1982,In_1715,In_2244);
or U1983 (N_1983,In_109,In_2222);
and U1984 (N_1984,In_907,In_2009);
xnor U1985 (N_1985,In_973,In_715);
nor U1986 (N_1986,In_1735,In_1619);
nand U1987 (N_1987,In_1387,In_1553);
nor U1988 (N_1988,In_791,In_1016);
and U1989 (N_1989,In_1322,In_86);
and U1990 (N_1990,In_1592,In_2188);
nor U1991 (N_1991,In_2311,In_1481);
nor U1992 (N_1992,In_2146,In_2227);
or U1993 (N_1993,In_220,In_1593);
nor U1994 (N_1994,In_120,In_513);
nor U1995 (N_1995,In_2071,In_2436);
and U1996 (N_1996,In_1949,In_1126);
or U1997 (N_1997,In_2265,In_1206);
and U1998 (N_1998,In_942,In_82);
nor U1999 (N_1999,In_57,In_2444);
nor U2000 (N_2000,In_1563,In_737);
nand U2001 (N_2001,In_671,In_1109);
nor U2002 (N_2002,In_1327,In_1559);
and U2003 (N_2003,In_2442,In_2411);
nor U2004 (N_2004,In_1386,In_1930);
nand U2005 (N_2005,In_258,In_369);
nor U2006 (N_2006,In_2437,In_1365);
nand U2007 (N_2007,In_1607,In_31);
nor U2008 (N_2008,In_1351,In_1247);
and U2009 (N_2009,In_880,In_2392);
or U2010 (N_2010,In_841,In_932);
nand U2011 (N_2011,In_1907,In_1364);
nor U2012 (N_2012,In_1239,In_614);
nor U2013 (N_2013,In_829,In_1289);
and U2014 (N_2014,In_228,In_1653);
nor U2015 (N_2015,In_1162,In_1076);
or U2016 (N_2016,In_1845,In_1786);
or U2017 (N_2017,In_1820,In_1743);
or U2018 (N_2018,In_1321,In_231);
nand U2019 (N_2019,In_218,In_2293);
or U2020 (N_2020,In_181,In_1335);
and U2021 (N_2021,In_2281,In_682);
xnor U2022 (N_2022,In_592,In_1583);
nand U2023 (N_2023,In_1111,In_1805);
nor U2024 (N_2024,In_2460,In_632);
or U2025 (N_2025,In_177,In_1873);
xnor U2026 (N_2026,In_1029,In_1368);
or U2027 (N_2027,In_1599,In_2264);
and U2028 (N_2028,In_1320,In_2441);
or U2029 (N_2029,In_2452,In_2038);
and U2030 (N_2030,In_154,In_1405);
nand U2031 (N_2031,In_1224,In_643);
or U2032 (N_2032,In_1570,In_1821);
nor U2033 (N_2033,In_521,In_1525);
nand U2034 (N_2034,In_1135,In_1133);
and U2035 (N_2035,In_2424,In_994);
nor U2036 (N_2036,In_2052,In_938);
or U2037 (N_2037,In_2234,In_1889);
or U2038 (N_2038,In_1337,In_1720);
and U2039 (N_2039,In_1313,In_1324);
and U2040 (N_2040,In_1540,In_1920);
or U2041 (N_2041,In_2000,In_1030);
or U2042 (N_2042,In_931,In_1537);
or U2043 (N_2043,In_398,In_2170);
and U2044 (N_2044,In_2390,In_314);
nand U2045 (N_2045,In_1816,In_2310);
and U2046 (N_2046,In_1155,In_98);
or U2047 (N_2047,In_155,In_2443);
nor U2048 (N_2048,In_1746,In_1074);
and U2049 (N_2049,In_1887,In_2241);
nand U2050 (N_2050,In_995,In_1218);
xor U2051 (N_2051,In_713,In_368);
or U2052 (N_2052,In_901,In_1706);
nor U2053 (N_2053,In_1945,In_1389);
or U2054 (N_2054,In_1865,In_2246);
and U2055 (N_2055,In_792,In_2023);
and U2056 (N_2056,In_1354,In_888);
and U2057 (N_2057,In_1262,In_890);
nand U2058 (N_2058,In_1184,In_1027);
nand U2059 (N_2059,In_1790,In_1825);
or U2060 (N_2060,In_2302,In_812);
or U2061 (N_2061,In_922,In_2110);
nor U2062 (N_2062,In_1393,In_191);
nor U2063 (N_2063,In_1934,In_493);
nor U2064 (N_2064,In_764,In_1018);
nand U2065 (N_2065,In_388,In_201);
xor U2066 (N_2066,In_224,In_2001);
nor U2067 (N_2067,In_436,In_45);
nor U2068 (N_2068,In_729,In_476);
and U2069 (N_2069,In_1611,In_1039);
and U2070 (N_2070,In_849,In_1577);
xor U2071 (N_2071,In_2424,In_438);
or U2072 (N_2072,In_1408,In_2307);
xnor U2073 (N_2073,In_920,In_2057);
and U2074 (N_2074,In_2155,In_1776);
nor U2075 (N_2075,In_2453,In_670);
nor U2076 (N_2076,In_393,In_1643);
and U2077 (N_2077,In_1678,In_1547);
and U2078 (N_2078,In_1177,In_244);
nand U2079 (N_2079,In_1869,In_1965);
nand U2080 (N_2080,In_1084,In_1208);
and U2081 (N_2081,In_699,In_621);
and U2082 (N_2082,In_1417,In_2213);
or U2083 (N_2083,In_1044,In_1437);
nor U2084 (N_2084,In_1787,In_1195);
nand U2085 (N_2085,In_394,In_1871);
or U2086 (N_2086,In_772,In_1066);
or U2087 (N_2087,In_1277,In_591);
nor U2088 (N_2088,In_206,In_399);
or U2089 (N_2089,In_1932,In_691);
nand U2090 (N_2090,In_792,In_1888);
nand U2091 (N_2091,In_1037,In_686);
or U2092 (N_2092,In_1082,In_1472);
or U2093 (N_2093,In_1546,In_362);
nor U2094 (N_2094,In_474,In_1515);
xor U2095 (N_2095,In_1982,In_823);
or U2096 (N_2096,In_2141,In_2328);
nor U2097 (N_2097,In_2264,In_2307);
or U2098 (N_2098,In_606,In_474);
and U2099 (N_2099,In_238,In_2090);
nand U2100 (N_2100,In_1869,In_619);
nand U2101 (N_2101,In_501,In_513);
and U2102 (N_2102,In_235,In_2424);
or U2103 (N_2103,In_2429,In_2105);
nor U2104 (N_2104,In_1872,In_1051);
and U2105 (N_2105,In_1812,In_817);
nor U2106 (N_2106,In_1424,In_408);
nand U2107 (N_2107,In_74,In_1048);
nand U2108 (N_2108,In_1576,In_2427);
or U2109 (N_2109,In_1025,In_2053);
and U2110 (N_2110,In_1250,In_1454);
nor U2111 (N_2111,In_603,In_463);
nand U2112 (N_2112,In_1101,In_848);
or U2113 (N_2113,In_74,In_1851);
or U2114 (N_2114,In_452,In_2445);
nor U2115 (N_2115,In_1329,In_1907);
xor U2116 (N_2116,In_453,In_816);
nand U2117 (N_2117,In_2474,In_695);
nor U2118 (N_2118,In_562,In_17);
and U2119 (N_2119,In_946,In_1332);
nor U2120 (N_2120,In_1774,In_1228);
and U2121 (N_2121,In_135,In_1620);
nor U2122 (N_2122,In_1255,In_214);
nor U2123 (N_2123,In_1750,In_2106);
and U2124 (N_2124,In_2235,In_2389);
and U2125 (N_2125,In_53,In_1213);
nand U2126 (N_2126,In_1924,In_1032);
or U2127 (N_2127,In_1623,In_1895);
and U2128 (N_2128,In_2164,In_2227);
or U2129 (N_2129,In_1005,In_1495);
nor U2130 (N_2130,In_1808,In_118);
nor U2131 (N_2131,In_2315,In_342);
and U2132 (N_2132,In_1074,In_1702);
and U2133 (N_2133,In_180,In_172);
nand U2134 (N_2134,In_2353,In_607);
nor U2135 (N_2135,In_2318,In_1992);
nand U2136 (N_2136,In_1004,In_1165);
or U2137 (N_2137,In_501,In_2250);
nor U2138 (N_2138,In_1127,In_64);
nor U2139 (N_2139,In_1707,In_1559);
and U2140 (N_2140,In_582,In_2246);
or U2141 (N_2141,In_795,In_1135);
nand U2142 (N_2142,In_2068,In_65);
nand U2143 (N_2143,In_2023,In_944);
xor U2144 (N_2144,In_2464,In_1480);
nor U2145 (N_2145,In_659,In_1725);
nand U2146 (N_2146,In_1909,In_1112);
or U2147 (N_2147,In_1534,In_948);
nand U2148 (N_2148,In_872,In_887);
and U2149 (N_2149,In_2038,In_236);
or U2150 (N_2150,In_888,In_125);
xor U2151 (N_2151,In_2292,In_1527);
nor U2152 (N_2152,In_929,In_863);
and U2153 (N_2153,In_1658,In_1173);
nand U2154 (N_2154,In_811,In_1180);
or U2155 (N_2155,In_2173,In_218);
or U2156 (N_2156,In_2117,In_1831);
or U2157 (N_2157,In_1430,In_2159);
nor U2158 (N_2158,In_763,In_432);
and U2159 (N_2159,In_1223,In_1119);
or U2160 (N_2160,In_675,In_944);
or U2161 (N_2161,In_1010,In_361);
or U2162 (N_2162,In_1228,In_1710);
nand U2163 (N_2163,In_1350,In_620);
nor U2164 (N_2164,In_1617,In_480);
and U2165 (N_2165,In_676,In_932);
and U2166 (N_2166,In_1116,In_489);
and U2167 (N_2167,In_1796,In_2254);
or U2168 (N_2168,In_121,In_1642);
and U2169 (N_2169,In_1424,In_2146);
and U2170 (N_2170,In_890,In_2010);
nand U2171 (N_2171,In_796,In_257);
or U2172 (N_2172,In_2243,In_1529);
or U2173 (N_2173,In_64,In_752);
and U2174 (N_2174,In_1480,In_1732);
or U2175 (N_2175,In_72,In_984);
nor U2176 (N_2176,In_1571,In_1324);
or U2177 (N_2177,In_621,In_2398);
nand U2178 (N_2178,In_2177,In_91);
nand U2179 (N_2179,In_1507,In_600);
nand U2180 (N_2180,In_2095,In_1805);
or U2181 (N_2181,In_341,In_2368);
xor U2182 (N_2182,In_1790,In_111);
and U2183 (N_2183,In_1643,In_239);
or U2184 (N_2184,In_38,In_1513);
nand U2185 (N_2185,In_1311,In_2247);
nor U2186 (N_2186,In_2375,In_2435);
and U2187 (N_2187,In_1083,In_783);
and U2188 (N_2188,In_493,In_1649);
nor U2189 (N_2189,In_1533,In_2374);
nor U2190 (N_2190,In_2111,In_187);
xnor U2191 (N_2191,In_1951,In_626);
xnor U2192 (N_2192,In_1496,In_654);
nand U2193 (N_2193,In_319,In_2314);
nor U2194 (N_2194,In_747,In_2046);
and U2195 (N_2195,In_1668,In_989);
nor U2196 (N_2196,In_246,In_1705);
and U2197 (N_2197,In_2481,In_1233);
and U2198 (N_2198,In_622,In_948);
nor U2199 (N_2199,In_623,In_2047);
or U2200 (N_2200,In_1541,In_1020);
and U2201 (N_2201,In_1339,In_93);
and U2202 (N_2202,In_1480,In_1343);
or U2203 (N_2203,In_2492,In_376);
nand U2204 (N_2204,In_759,In_1740);
nand U2205 (N_2205,In_1364,In_983);
nor U2206 (N_2206,In_1067,In_2482);
and U2207 (N_2207,In_172,In_1352);
nor U2208 (N_2208,In_65,In_335);
and U2209 (N_2209,In_662,In_810);
or U2210 (N_2210,In_732,In_1753);
nand U2211 (N_2211,In_1354,In_1924);
nor U2212 (N_2212,In_1770,In_1315);
or U2213 (N_2213,In_1258,In_168);
or U2214 (N_2214,In_855,In_1434);
nor U2215 (N_2215,In_2471,In_1174);
nor U2216 (N_2216,In_608,In_42);
nor U2217 (N_2217,In_1287,In_428);
and U2218 (N_2218,In_707,In_277);
nor U2219 (N_2219,In_612,In_166);
nor U2220 (N_2220,In_1710,In_635);
nand U2221 (N_2221,In_311,In_865);
nand U2222 (N_2222,In_1840,In_1459);
or U2223 (N_2223,In_1933,In_766);
nor U2224 (N_2224,In_1324,In_1783);
or U2225 (N_2225,In_429,In_656);
nand U2226 (N_2226,In_285,In_989);
and U2227 (N_2227,In_2390,In_1061);
nor U2228 (N_2228,In_1914,In_424);
or U2229 (N_2229,In_1608,In_183);
nand U2230 (N_2230,In_194,In_1890);
nor U2231 (N_2231,In_154,In_2244);
or U2232 (N_2232,In_1021,In_1721);
nand U2233 (N_2233,In_2072,In_1939);
and U2234 (N_2234,In_1311,In_1811);
or U2235 (N_2235,In_2427,In_2477);
nand U2236 (N_2236,In_2300,In_1904);
xor U2237 (N_2237,In_986,In_327);
and U2238 (N_2238,In_1527,In_2073);
and U2239 (N_2239,In_1171,In_938);
nand U2240 (N_2240,In_1029,In_2022);
and U2241 (N_2241,In_725,In_1907);
nor U2242 (N_2242,In_2476,In_53);
nand U2243 (N_2243,In_2304,In_1339);
nor U2244 (N_2244,In_2180,In_2429);
nand U2245 (N_2245,In_521,In_1812);
and U2246 (N_2246,In_2339,In_37);
or U2247 (N_2247,In_1657,In_454);
nor U2248 (N_2248,In_96,In_360);
nand U2249 (N_2249,In_942,In_2442);
and U2250 (N_2250,In_405,In_571);
or U2251 (N_2251,In_1338,In_106);
nor U2252 (N_2252,In_37,In_2112);
or U2253 (N_2253,In_283,In_1490);
nand U2254 (N_2254,In_1802,In_1574);
nor U2255 (N_2255,In_1313,In_1157);
xnor U2256 (N_2256,In_318,In_817);
nand U2257 (N_2257,In_1391,In_1679);
nand U2258 (N_2258,In_573,In_841);
and U2259 (N_2259,In_1786,In_2212);
xnor U2260 (N_2260,In_808,In_2034);
xnor U2261 (N_2261,In_2228,In_173);
nor U2262 (N_2262,In_790,In_2084);
nand U2263 (N_2263,In_2267,In_571);
xor U2264 (N_2264,In_692,In_380);
nor U2265 (N_2265,In_1338,In_2341);
nand U2266 (N_2266,In_1477,In_1685);
or U2267 (N_2267,In_1930,In_122);
nor U2268 (N_2268,In_1756,In_2216);
nor U2269 (N_2269,In_1478,In_196);
or U2270 (N_2270,In_1508,In_622);
and U2271 (N_2271,In_1155,In_2187);
nand U2272 (N_2272,In_1268,In_1383);
xor U2273 (N_2273,In_1027,In_2342);
and U2274 (N_2274,In_214,In_2001);
or U2275 (N_2275,In_560,In_796);
and U2276 (N_2276,In_1514,In_1169);
nor U2277 (N_2277,In_2305,In_2382);
or U2278 (N_2278,In_753,In_667);
nor U2279 (N_2279,In_2280,In_1711);
and U2280 (N_2280,In_645,In_1507);
and U2281 (N_2281,In_1554,In_579);
nand U2282 (N_2282,In_1467,In_1996);
or U2283 (N_2283,In_1211,In_1837);
xor U2284 (N_2284,In_86,In_2312);
and U2285 (N_2285,In_2310,In_2345);
and U2286 (N_2286,In_742,In_1542);
or U2287 (N_2287,In_1738,In_1310);
xnor U2288 (N_2288,In_2242,In_652);
or U2289 (N_2289,In_2082,In_2466);
nand U2290 (N_2290,In_1691,In_842);
or U2291 (N_2291,In_1679,In_959);
or U2292 (N_2292,In_1601,In_2045);
nand U2293 (N_2293,In_729,In_1691);
or U2294 (N_2294,In_1064,In_1167);
or U2295 (N_2295,In_1213,In_21);
or U2296 (N_2296,In_941,In_2268);
xnor U2297 (N_2297,In_1666,In_1907);
nand U2298 (N_2298,In_881,In_661);
and U2299 (N_2299,In_622,In_2409);
nand U2300 (N_2300,In_847,In_552);
nor U2301 (N_2301,In_1380,In_835);
nand U2302 (N_2302,In_2402,In_1706);
nand U2303 (N_2303,In_2126,In_2499);
nor U2304 (N_2304,In_262,In_2112);
xnor U2305 (N_2305,In_1577,In_1039);
nor U2306 (N_2306,In_719,In_1250);
and U2307 (N_2307,In_1479,In_1281);
xor U2308 (N_2308,In_1488,In_2022);
or U2309 (N_2309,In_2312,In_119);
nand U2310 (N_2310,In_699,In_2473);
xnor U2311 (N_2311,In_509,In_726);
xor U2312 (N_2312,In_1989,In_886);
nor U2313 (N_2313,In_818,In_1839);
nand U2314 (N_2314,In_53,In_208);
and U2315 (N_2315,In_738,In_529);
nand U2316 (N_2316,In_414,In_1827);
nand U2317 (N_2317,In_3,In_1612);
and U2318 (N_2318,In_807,In_208);
nand U2319 (N_2319,In_184,In_1392);
or U2320 (N_2320,In_2256,In_441);
nor U2321 (N_2321,In_250,In_1144);
nand U2322 (N_2322,In_2140,In_706);
nor U2323 (N_2323,In_566,In_1693);
or U2324 (N_2324,In_14,In_1945);
and U2325 (N_2325,In_906,In_717);
nor U2326 (N_2326,In_2116,In_2358);
or U2327 (N_2327,In_751,In_1537);
xor U2328 (N_2328,In_2365,In_1456);
nor U2329 (N_2329,In_1924,In_2466);
xnor U2330 (N_2330,In_2173,In_1878);
or U2331 (N_2331,In_1292,In_2249);
and U2332 (N_2332,In_1626,In_745);
or U2333 (N_2333,In_1283,In_774);
nor U2334 (N_2334,In_440,In_657);
nor U2335 (N_2335,In_1142,In_881);
nand U2336 (N_2336,In_2067,In_125);
or U2337 (N_2337,In_368,In_21);
and U2338 (N_2338,In_32,In_2109);
nor U2339 (N_2339,In_90,In_11);
and U2340 (N_2340,In_152,In_2318);
nor U2341 (N_2341,In_1268,In_2068);
or U2342 (N_2342,In_1717,In_1829);
nand U2343 (N_2343,In_2165,In_289);
nand U2344 (N_2344,In_692,In_989);
or U2345 (N_2345,In_1607,In_1964);
or U2346 (N_2346,In_525,In_2011);
nand U2347 (N_2347,In_811,In_995);
nor U2348 (N_2348,In_1643,In_1670);
xnor U2349 (N_2349,In_2369,In_2163);
nand U2350 (N_2350,In_1660,In_521);
and U2351 (N_2351,In_1876,In_2263);
or U2352 (N_2352,In_2470,In_1515);
xnor U2353 (N_2353,In_948,In_2306);
nand U2354 (N_2354,In_2308,In_895);
nor U2355 (N_2355,In_2351,In_2374);
nor U2356 (N_2356,In_436,In_633);
and U2357 (N_2357,In_747,In_1975);
xnor U2358 (N_2358,In_1694,In_919);
nor U2359 (N_2359,In_1336,In_786);
xor U2360 (N_2360,In_1552,In_1462);
or U2361 (N_2361,In_2245,In_1022);
nand U2362 (N_2362,In_168,In_442);
or U2363 (N_2363,In_182,In_547);
xnor U2364 (N_2364,In_106,In_2305);
or U2365 (N_2365,In_1818,In_591);
or U2366 (N_2366,In_2196,In_1831);
nand U2367 (N_2367,In_1999,In_66);
nand U2368 (N_2368,In_1999,In_2321);
or U2369 (N_2369,In_1467,In_2256);
or U2370 (N_2370,In_955,In_2464);
nor U2371 (N_2371,In_673,In_775);
xor U2372 (N_2372,In_563,In_2065);
or U2373 (N_2373,In_842,In_1140);
or U2374 (N_2374,In_827,In_2457);
or U2375 (N_2375,In_264,In_1286);
or U2376 (N_2376,In_2001,In_1836);
or U2377 (N_2377,In_260,In_2111);
or U2378 (N_2378,In_2316,In_1104);
xnor U2379 (N_2379,In_1258,In_2385);
and U2380 (N_2380,In_2058,In_2209);
and U2381 (N_2381,In_2477,In_1793);
nor U2382 (N_2382,In_673,In_2273);
or U2383 (N_2383,In_1019,In_1586);
or U2384 (N_2384,In_1357,In_1245);
xnor U2385 (N_2385,In_944,In_40);
nand U2386 (N_2386,In_193,In_2087);
and U2387 (N_2387,In_2300,In_733);
nand U2388 (N_2388,In_2161,In_794);
nor U2389 (N_2389,In_1012,In_1235);
nand U2390 (N_2390,In_2470,In_1668);
and U2391 (N_2391,In_2271,In_1863);
nand U2392 (N_2392,In_685,In_1413);
nor U2393 (N_2393,In_1671,In_655);
nand U2394 (N_2394,In_1389,In_361);
nor U2395 (N_2395,In_0,In_2055);
nand U2396 (N_2396,In_512,In_1742);
and U2397 (N_2397,In_338,In_1984);
nor U2398 (N_2398,In_2144,In_290);
and U2399 (N_2399,In_1768,In_394);
xnor U2400 (N_2400,In_1562,In_740);
or U2401 (N_2401,In_1156,In_1732);
xor U2402 (N_2402,In_2409,In_520);
nand U2403 (N_2403,In_1923,In_2094);
and U2404 (N_2404,In_1462,In_1770);
xor U2405 (N_2405,In_1316,In_439);
nand U2406 (N_2406,In_517,In_2156);
nand U2407 (N_2407,In_1999,In_154);
nand U2408 (N_2408,In_718,In_1720);
and U2409 (N_2409,In_846,In_1381);
or U2410 (N_2410,In_1312,In_1604);
and U2411 (N_2411,In_1377,In_675);
or U2412 (N_2412,In_658,In_1655);
nor U2413 (N_2413,In_105,In_317);
or U2414 (N_2414,In_1187,In_2311);
and U2415 (N_2415,In_2293,In_1503);
nand U2416 (N_2416,In_315,In_1911);
xor U2417 (N_2417,In_552,In_928);
nor U2418 (N_2418,In_28,In_1630);
nand U2419 (N_2419,In_2037,In_934);
nor U2420 (N_2420,In_1021,In_908);
xnor U2421 (N_2421,In_2290,In_1473);
nand U2422 (N_2422,In_2371,In_1402);
and U2423 (N_2423,In_617,In_2090);
or U2424 (N_2424,In_2494,In_445);
xnor U2425 (N_2425,In_1798,In_2216);
or U2426 (N_2426,In_552,In_1023);
or U2427 (N_2427,In_26,In_1472);
or U2428 (N_2428,In_834,In_1503);
and U2429 (N_2429,In_60,In_1775);
nor U2430 (N_2430,In_1359,In_768);
nor U2431 (N_2431,In_2428,In_1886);
nor U2432 (N_2432,In_616,In_1707);
nor U2433 (N_2433,In_1703,In_1282);
and U2434 (N_2434,In_543,In_1338);
nor U2435 (N_2435,In_273,In_806);
nand U2436 (N_2436,In_40,In_1848);
and U2437 (N_2437,In_2337,In_1022);
or U2438 (N_2438,In_2106,In_1948);
or U2439 (N_2439,In_2445,In_1820);
and U2440 (N_2440,In_1276,In_1375);
nand U2441 (N_2441,In_445,In_6);
nor U2442 (N_2442,In_1489,In_2356);
xor U2443 (N_2443,In_2442,In_203);
or U2444 (N_2444,In_628,In_1696);
and U2445 (N_2445,In_2496,In_396);
and U2446 (N_2446,In_203,In_883);
or U2447 (N_2447,In_2120,In_1279);
nor U2448 (N_2448,In_826,In_1543);
nand U2449 (N_2449,In_1443,In_551);
nor U2450 (N_2450,In_664,In_1917);
or U2451 (N_2451,In_1989,In_1158);
nor U2452 (N_2452,In_1806,In_2148);
or U2453 (N_2453,In_1416,In_1420);
and U2454 (N_2454,In_2024,In_945);
nand U2455 (N_2455,In_71,In_1275);
or U2456 (N_2456,In_1187,In_968);
or U2457 (N_2457,In_2135,In_796);
nor U2458 (N_2458,In_1317,In_280);
nand U2459 (N_2459,In_2141,In_266);
or U2460 (N_2460,In_1299,In_298);
and U2461 (N_2461,In_2059,In_753);
xor U2462 (N_2462,In_427,In_868);
or U2463 (N_2463,In_920,In_246);
nor U2464 (N_2464,In_2348,In_395);
nand U2465 (N_2465,In_2427,In_428);
nor U2466 (N_2466,In_253,In_35);
or U2467 (N_2467,In_309,In_909);
nor U2468 (N_2468,In_123,In_817);
nor U2469 (N_2469,In_1415,In_545);
and U2470 (N_2470,In_801,In_1273);
and U2471 (N_2471,In_1064,In_1105);
or U2472 (N_2472,In_54,In_1490);
nand U2473 (N_2473,In_2312,In_343);
xnor U2474 (N_2474,In_1322,In_2480);
or U2475 (N_2475,In_1158,In_333);
nand U2476 (N_2476,In_109,In_288);
xor U2477 (N_2477,In_138,In_1999);
xor U2478 (N_2478,In_1003,In_2322);
nand U2479 (N_2479,In_402,In_989);
and U2480 (N_2480,In_334,In_2138);
xnor U2481 (N_2481,In_972,In_1700);
xnor U2482 (N_2482,In_2379,In_162);
or U2483 (N_2483,In_2128,In_2058);
nor U2484 (N_2484,In_1611,In_1610);
nand U2485 (N_2485,In_2115,In_96);
and U2486 (N_2486,In_835,In_661);
xor U2487 (N_2487,In_1329,In_2300);
and U2488 (N_2488,In_329,In_63);
or U2489 (N_2489,In_1648,In_2454);
or U2490 (N_2490,In_2063,In_1437);
and U2491 (N_2491,In_571,In_1852);
or U2492 (N_2492,In_805,In_290);
and U2493 (N_2493,In_25,In_1610);
nor U2494 (N_2494,In_1381,In_1279);
nor U2495 (N_2495,In_202,In_1353);
nand U2496 (N_2496,In_117,In_1603);
xor U2497 (N_2497,In_394,In_1652);
and U2498 (N_2498,In_629,In_116);
nor U2499 (N_2499,In_1007,In_279);
nor U2500 (N_2500,In_1455,In_52);
and U2501 (N_2501,In_266,In_1923);
nor U2502 (N_2502,In_2135,In_481);
nand U2503 (N_2503,In_2236,In_1079);
nand U2504 (N_2504,In_2153,In_414);
nor U2505 (N_2505,In_2007,In_2265);
xor U2506 (N_2506,In_1939,In_2116);
and U2507 (N_2507,In_522,In_221);
nand U2508 (N_2508,In_675,In_2046);
or U2509 (N_2509,In_2118,In_2165);
nor U2510 (N_2510,In_2353,In_1802);
nor U2511 (N_2511,In_1960,In_480);
and U2512 (N_2512,In_1260,In_1215);
nand U2513 (N_2513,In_1187,In_1764);
and U2514 (N_2514,In_1273,In_394);
nand U2515 (N_2515,In_2485,In_1630);
and U2516 (N_2516,In_1908,In_516);
nand U2517 (N_2517,In_79,In_2480);
or U2518 (N_2518,In_1555,In_153);
and U2519 (N_2519,In_497,In_1495);
and U2520 (N_2520,In_1260,In_842);
nor U2521 (N_2521,In_789,In_1262);
nor U2522 (N_2522,In_300,In_2269);
and U2523 (N_2523,In_2189,In_922);
nand U2524 (N_2524,In_885,In_1875);
nand U2525 (N_2525,In_1741,In_1190);
or U2526 (N_2526,In_1979,In_325);
nor U2527 (N_2527,In_343,In_461);
xor U2528 (N_2528,In_1320,In_14);
or U2529 (N_2529,In_1548,In_513);
and U2530 (N_2530,In_461,In_133);
and U2531 (N_2531,In_2064,In_2369);
or U2532 (N_2532,In_1601,In_367);
nand U2533 (N_2533,In_2332,In_1919);
or U2534 (N_2534,In_538,In_1064);
or U2535 (N_2535,In_1118,In_252);
nand U2536 (N_2536,In_844,In_1276);
and U2537 (N_2537,In_570,In_1989);
or U2538 (N_2538,In_2295,In_118);
nand U2539 (N_2539,In_2483,In_2496);
nor U2540 (N_2540,In_1846,In_2260);
nand U2541 (N_2541,In_1867,In_2170);
xor U2542 (N_2542,In_658,In_950);
and U2543 (N_2543,In_301,In_250);
or U2544 (N_2544,In_571,In_1357);
and U2545 (N_2545,In_1087,In_907);
or U2546 (N_2546,In_842,In_2111);
and U2547 (N_2547,In_137,In_1861);
nand U2548 (N_2548,In_1453,In_1898);
nand U2549 (N_2549,In_2005,In_1400);
nand U2550 (N_2550,In_1393,In_1620);
or U2551 (N_2551,In_285,In_2251);
or U2552 (N_2552,In_859,In_730);
and U2553 (N_2553,In_2466,In_2165);
xnor U2554 (N_2554,In_1075,In_232);
nand U2555 (N_2555,In_2395,In_1691);
nand U2556 (N_2556,In_554,In_114);
and U2557 (N_2557,In_1587,In_1331);
nor U2558 (N_2558,In_1715,In_415);
nand U2559 (N_2559,In_84,In_237);
nor U2560 (N_2560,In_2479,In_264);
or U2561 (N_2561,In_2316,In_262);
xnor U2562 (N_2562,In_2362,In_7);
nor U2563 (N_2563,In_27,In_488);
and U2564 (N_2564,In_2032,In_1041);
nor U2565 (N_2565,In_2076,In_225);
nand U2566 (N_2566,In_1539,In_1308);
nand U2567 (N_2567,In_1680,In_1135);
and U2568 (N_2568,In_777,In_1165);
and U2569 (N_2569,In_2120,In_350);
and U2570 (N_2570,In_1557,In_1966);
and U2571 (N_2571,In_1413,In_1843);
and U2572 (N_2572,In_1214,In_598);
nand U2573 (N_2573,In_1380,In_572);
nand U2574 (N_2574,In_1567,In_385);
and U2575 (N_2575,In_1427,In_2392);
and U2576 (N_2576,In_2144,In_1662);
nor U2577 (N_2577,In_34,In_879);
or U2578 (N_2578,In_765,In_1591);
xor U2579 (N_2579,In_488,In_996);
xnor U2580 (N_2580,In_1822,In_2218);
nor U2581 (N_2581,In_1309,In_1303);
or U2582 (N_2582,In_1955,In_981);
and U2583 (N_2583,In_1725,In_2063);
nand U2584 (N_2584,In_1396,In_668);
or U2585 (N_2585,In_130,In_1266);
or U2586 (N_2586,In_317,In_2115);
nand U2587 (N_2587,In_1177,In_676);
and U2588 (N_2588,In_484,In_1119);
or U2589 (N_2589,In_343,In_2405);
nand U2590 (N_2590,In_1957,In_293);
nand U2591 (N_2591,In_271,In_707);
and U2592 (N_2592,In_2042,In_2351);
nand U2593 (N_2593,In_1726,In_1683);
nor U2594 (N_2594,In_496,In_1803);
and U2595 (N_2595,In_2052,In_156);
nand U2596 (N_2596,In_160,In_2365);
or U2597 (N_2597,In_989,In_2309);
nor U2598 (N_2598,In_1539,In_1230);
and U2599 (N_2599,In_1160,In_1671);
or U2600 (N_2600,In_343,In_2016);
nand U2601 (N_2601,In_1621,In_530);
nor U2602 (N_2602,In_799,In_1055);
nor U2603 (N_2603,In_1176,In_1865);
and U2604 (N_2604,In_1922,In_2393);
nand U2605 (N_2605,In_1227,In_1496);
or U2606 (N_2606,In_2167,In_2107);
nor U2607 (N_2607,In_976,In_271);
xnor U2608 (N_2608,In_1096,In_588);
and U2609 (N_2609,In_1093,In_1738);
xor U2610 (N_2610,In_1956,In_2472);
nor U2611 (N_2611,In_679,In_1391);
and U2612 (N_2612,In_1141,In_533);
xor U2613 (N_2613,In_28,In_454);
nor U2614 (N_2614,In_1299,In_1009);
and U2615 (N_2615,In_1805,In_2497);
and U2616 (N_2616,In_2125,In_2467);
and U2617 (N_2617,In_2090,In_2176);
nor U2618 (N_2618,In_118,In_165);
xor U2619 (N_2619,In_2395,In_1332);
nor U2620 (N_2620,In_90,In_969);
nand U2621 (N_2621,In_1210,In_1939);
and U2622 (N_2622,In_2216,In_1994);
or U2623 (N_2623,In_2231,In_1265);
or U2624 (N_2624,In_1616,In_731);
or U2625 (N_2625,In_1431,In_1720);
or U2626 (N_2626,In_1728,In_1462);
nor U2627 (N_2627,In_53,In_2033);
nand U2628 (N_2628,In_2481,In_2470);
and U2629 (N_2629,In_604,In_1618);
or U2630 (N_2630,In_715,In_2049);
nor U2631 (N_2631,In_1255,In_2385);
nor U2632 (N_2632,In_654,In_1495);
nor U2633 (N_2633,In_2067,In_2017);
and U2634 (N_2634,In_26,In_822);
nand U2635 (N_2635,In_1647,In_970);
nand U2636 (N_2636,In_632,In_90);
nor U2637 (N_2637,In_2372,In_2026);
nand U2638 (N_2638,In_1262,In_2108);
and U2639 (N_2639,In_124,In_1392);
nand U2640 (N_2640,In_2402,In_1176);
nand U2641 (N_2641,In_1233,In_26);
xor U2642 (N_2642,In_25,In_2059);
xor U2643 (N_2643,In_2037,In_1343);
nand U2644 (N_2644,In_1827,In_202);
nand U2645 (N_2645,In_2130,In_585);
nand U2646 (N_2646,In_115,In_199);
nor U2647 (N_2647,In_1741,In_1018);
nor U2648 (N_2648,In_1371,In_361);
nand U2649 (N_2649,In_1546,In_1588);
xor U2650 (N_2650,In_1791,In_941);
and U2651 (N_2651,In_960,In_893);
xor U2652 (N_2652,In_1546,In_9);
nand U2653 (N_2653,In_1320,In_1928);
and U2654 (N_2654,In_492,In_1988);
nor U2655 (N_2655,In_201,In_1439);
and U2656 (N_2656,In_2026,In_2051);
and U2657 (N_2657,In_805,In_263);
and U2658 (N_2658,In_206,In_487);
nand U2659 (N_2659,In_1687,In_1629);
or U2660 (N_2660,In_2049,In_635);
nor U2661 (N_2661,In_1282,In_1482);
nor U2662 (N_2662,In_2166,In_1873);
nand U2663 (N_2663,In_2120,In_1715);
or U2664 (N_2664,In_190,In_113);
or U2665 (N_2665,In_227,In_28);
nor U2666 (N_2666,In_1987,In_896);
or U2667 (N_2667,In_736,In_314);
or U2668 (N_2668,In_1920,In_1126);
or U2669 (N_2669,In_1372,In_677);
or U2670 (N_2670,In_522,In_155);
and U2671 (N_2671,In_588,In_1807);
nand U2672 (N_2672,In_1601,In_308);
or U2673 (N_2673,In_1691,In_2417);
nor U2674 (N_2674,In_2326,In_1794);
and U2675 (N_2675,In_2293,In_424);
or U2676 (N_2676,In_425,In_473);
and U2677 (N_2677,In_1647,In_1318);
or U2678 (N_2678,In_949,In_669);
or U2679 (N_2679,In_1346,In_2003);
nand U2680 (N_2680,In_1000,In_648);
or U2681 (N_2681,In_318,In_2133);
and U2682 (N_2682,In_604,In_243);
xnor U2683 (N_2683,In_1677,In_1811);
nand U2684 (N_2684,In_223,In_895);
nor U2685 (N_2685,In_656,In_1368);
and U2686 (N_2686,In_895,In_2092);
and U2687 (N_2687,In_194,In_837);
nor U2688 (N_2688,In_2102,In_894);
and U2689 (N_2689,In_532,In_497);
xnor U2690 (N_2690,In_324,In_887);
nor U2691 (N_2691,In_1524,In_110);
nor U2692 (N_2692,In_997,In_2002);
and U2693 (N_2693,In_1673,In_2304);
nor U2694 (N_2694,In_746,In_2437);
or U2695 (N_2695,In_194,In_1220);
nand U2696 (N_2696,In_2396,In_2195);
and U2697 (N_2697,In_1560,In_1196);
or U2698 (N_2698,In_1623,In_892);
or U2699 (N_2699,In_2227,In_58);
and U2700 (N_2700,In_160,In_1937);
or U2701 (N_2701,In_1667,In_516);
or U2702 (N_2702,In_2281,In_2098);
xnor U2703 (N_2703,In_682,In_2482);
or U2704 (N_2704,In_1928,In_2023);
or U2705 (N_2705,In_247,In_984);
nand U2706 (N_2706,In_1669,In_1685);
and U2707 (N_2707,In_1712,In_1186);
xor U2708 (N_2708,In_38,In_1638);
nor U2709 (N_2709,In_2469,In_311);
nand U2710 (N_2710,In_2110,In_2358);
or U2711 (N_2711,In_978,In_1071);
or U2712 (N_2712,In_590,In_2459);
nor U2713 (N_2713,In_580,In_461);
xor U2714 (N_2714,In_581,In_143);
nor U2715 (N_2715,In_1739,In_330);
or U2716 (N_2716,In_1148,In_1502);
nand U2717 (N_2717,In_670,In_2469);
xor U2718 (N_2718,In_1027,In_2364);
nor U2719 (N_2719,In_1369,In_2383);
nor U2720 (N_2720,In_279,In_612);
nand U2721 (N_2721,In_1473,In_1318);
or U2722 (N_2722,In_927,In_174);
nand U2723 (N_2723,In_1483,In_428);
or U2724 (N_2724,In_271,In_1007);
xor U2725 (N_2725,In_925,In_1392);
and U2726 (N_2726,In_212,In_2064);
and U2727 (N_2727,In_821,In_2101);
or U2728 (N_2728,In_2036,In_2401);
or U2729 (N_2729,In_156,In_809);
nand U2730 (N_2730,In_545,In_2196);
xnor U2731 (N_2731,In_1272,In_34);
and U2732 (N_2732,In_1809,In_1504);
xnor U2733 (N_2733,In_80,In_1653);
or U2734 (N_2734,In_1833,In_1065);
nor U2735 (N_2735,In_289,In_976);
nor U2736 (N_2736,In_1836,In_1979);
and U2737 (N_2737,In_2197,In_1231);
nand U2738 (N_2738,In_1320,In_1084);
or U2739 (N_2739,In_1984,In_1149);
nor U2740 (N_2740,In_1278,In_1901);
nor U2741 (N_2741,In_301,In_1030);
nor U2742 (N_2742,In_1492,In_1793);
nand U2743 (N_2743,In_936,In_1493);
xnor U2744 (N_2744,In_1744,In_1110);
xor U2745 (N_2745,In_2356,In_99);
nor U2746 (N_2746,In_1532,In_2494);
xnor U2747 (N_2747,In_319,In_1084);
or U2748 (N_2748,In_1690,In_1472);
nand U2749 (N_2749,In_0,In_86);
and U2750 (N_2750,In_52,In_312);
nand U2751 (N_2751,In_2028,In_1660);
nand U2752 (N_2752,In_1944,In_2388);
and U2753 (N_2753,In_1444,In_1440);
nand U2754 (N_2754,In_1566,In_599);
or U2755 (N_2755,In_143,In_283);
or U2756 (N_2756,In_203,In_606);
xnor U2757 (N_2757,In_528,In_2450);
xor U2758 (N_2758,In_1507,In_1049);
or U2759 (N_2759,In_1912,In_321);
or U2760 (N_2760,In_983,In_1690);
nand U2761 (N_2761,In_614,In_1517);
nand U2762 (N_2762,In_933,In_1732);
nor U2763 (N_2763,In_513,In_2363);
and U2764 (N_2764,In_2121,In_1582);
nor U2765 (N_2765,In_1382,In_1820);
or U2766 (N_2766,In_2089,In_1150);
and U2767 (N_2767,In_1457,In_2383);
and U2768 (N_2768,In_448,In_1611);
nand U2769 (N_2769,In_739,In_2084);
xor U2770 (N_2770,In_1950,In_296);
nand U2771 (N_2771,In_2261,In_1366);
or U2772 (N_2772,In_1612,In_1788);
nor U2773 (N_2773,In_159,In_1366);
nor U2774 (N_2774,In_1980,In_987);
and U2775 (N_2775,In_2035,In_2074);
and U2776 (N_2776,In_301,In_385);
nand U2777 (N_2777,In_2190,In_1829);
nand U2778 (N_2778,In_534,In_1805);
or U2779 (N_2779,In_584,In_139);
or U2780 (N_2780,In_2170,In_1737);
and U2781 (N_2781,In_1820,In_1578);
nor U2782 (N_2782,In_1636,In_1975);
nor U2783 (N_2783,In_211,In_1795);
nor U2784 (N_2784,In_15,In_897);
xor U2785 (N_2785,In_961,In_2265);
nor U2786 (N_2786,In_126,In_197);
or U2787 (N_2787,In_2465,In_2386);
nor U2788 (N_2788,In_419,In_671);
or U2789 (N_2789,In_590,In_65);
nand U2790 (N_2790,In_612,In_365);
nor U2791 (N_2791,In_559,In_1787);
or U2792 (N_2792,In_1175,In_445);
and U2793 (N_2793,In_2044,In_741);
nand U2794 (N_2794,In_881,In_2025);
nand U2795 (N_2795,In_2142,In_508);
or U2796 (N_2796,In_708,In_1198);
or U2797 (N_2797,In_1366,In_358);
nor U2798 (N_2798,In_180,In_1031);
nor U2799 (N_2799,In_1722,In_408);
nor U2800 (N_2800,In_2097,In_983);
nor U2801 (N_2801,In_2187,In_9);
or U2802 (N_2802,In_169,In_793);
nand U2803 (N_2803,In_2011,In_2397);
or U2804 (N_2804,In_199,In_263);
nand U2805 (N_2805,In_961,In_595);
nand U2806 (N_2806,In_2278,In_1546);
nand U2807 (N_2807,In_1897,In_643);
and U2808 (N_2808,In_1803,In_2221);
nor U2809 (N_2809,In_198,In_1114);
and U2810 (N_2810,In_166,In_2247);
or U2811 (N_2811,In_1212,In_301);
nor U2812 (N_2812,In_1378,In_117);
nand U2813 (N_2813,In_644,In_2405);
xnor U2814 (N_2814,In_656,In_396);
nand U2815 (N_2815,In_669,In_1630);
and U2816 (N_2816,In_1976,In_2077);
nor U2817 (N_2817,In_235,In_1320);
and U2818 (N_2818,In_467,In_1490);
or U2819 (N_2819,In_892,In_2284);
xnor U2820 (N_2820,In_2276,In_1852);
and U2821 (N_2821,In_612,In_2087);
nor U2822 (N_2822,In_1286,In_1751);
and U2823 (N_2823,In_1799,In_601);
nor U2824 (N_2824,In_7,In_89);
or U2825 (N_2825,In_2482,In_796);
and U2826 (N_2826,In_1348,In_1373);
and U2827 (N_2827,In_1534,In_334);
nand U2828 (N_2828,In_1543,In_415);
and U2829 (N_2829,In_618,In_532);
and U2830 (N_2830,In_2442,In_677);
nand U2831 (N_2831,In_396,In_649);
or U2832 (N_2832,In_1298,In_1802);
nor U2833 (N_2833,In_320,In_2253);
or U2834 (N_2834,In_2031,In_1509);
xor U2835 (N_2835,In_1854,In_33);
and U2836 (N_2836,In_41,In_581);
nand U2837 (N_2837,In_530,In_596);
and U2838 (N_2838,In_642,In_1843);
and U2839 (N_2839,In_2047,In_1347);
xnor U2840 (N_2840,In_1920,In_2461);
or U2841 (N_2841,In_1614,In_1521);
nand U2842 (N_2842,In_652,In_2405);
nor U2843 (N_2843,In_2284,In_834);
or U2844 (N_2844,In_672,In_821);
or U2845 (N_2845,In_2078,In_575);
and U2846 (N_2846,In_972,In_1399);
and U2847 (N_2847,In_540,In_1874);
or U2848 (N_2848,In_2079,In_984);
nor U2849 (N_2849,In_782,In_1575);
nor U2850 (N_2850,In_665,In_461);
or U2851 (N_2851,In_234,In_1172);
or U2852 (N_2852,In_1104,In_1519);
nor U2853 (N_2853,In_1397,In_361);
nand U2854 (N_2854,In_2166,In_1875);
nor U2855 (N_2855,In_787,In_213);
nor U2856 (N_2856,In_146,In_1736);
or U2857 (N_2857,In_1980,In_1541);
or U2858 (N_2858,In_1927,In_510);
nand U2859 (N_2859,In_2476,In_1494);
or U2860 (N_2860,In_684,In_403);
or U2861 (N_2861,In_1786,In_2375);
nor U2862 (N_2862,In_2361,In_309);
nand U2863 (N_2863,In_1635,In_1358);
xnor U2864 (N_2864,In_360,In_1265);
and U2865 (N_2865,In_2302,In_1339);
nand U2866 (N_2866,In_1520,In_1693);
or U2867 (N_2867,In_1687,In_1893);
nand U2868 (N_2868,In_110,In_1548);
and U2869 (N_2869,In_2098,In_1283);
or U2870 (N_2870,In_989,In_2024);
nor U2871 (N_2871,In_111,In_1225);
xor U2872 (N_2872,In_771,In_384);
nand U2873 (N_2873,In_799,In_1403);
or U2874 (N_2874,In_2165,In_576);
nand U2875 (N_2875,In_898,In_1531);
and U2876 (N_2876,In_1727,In_221);
nor U2877 (N_2877,In_1578,In_969);
or U2878 (N_2878,In_940,In_1998);
nor U2879 (N_2879,In_496,In_969);
nand U2880 (N_2880,In_2235,In_282);
or U2881 (N_2881,In_2324,In_2316);
nor U2882 (N_2882,In_66,In_1982);
and U2883 (N_2883,In_1242,In_2210);
and U2884 (N_2884,In_2009,In_845);
nor U2885 (N_2885,In_1948,In_1108);
nor U2886 (N_2886,In_2305,In_1869);
and U2887 (N_2887,In_1070,In_478);
and U2888 (N_2888,In_2283,In_100);
and U2889 (N_2889,In_2172,In_1956);
and U2890 (N_2890,In_1039,In_2259);
nand U2891 (N_2891,In_806,In_1213);
xnor U2892 (N_2892,In_649,In_11);
or U2893 (N_2893,In_1315,In_1254);
or U2894 (N_2894,In_1759,In_1981);
nand U2895 (N_2895,In_1847,In_2095);
nor U2896 (N_2896,In_285,In_1282);
nor U2897 (N_2897,In_279,In_375);
and U2898 (N_2898,In_1847,In_1532);
and U2899 (N_2899,In_1243,In_2200);
nand U2900 (N_2900,In_1615,In_2190);
nand U2901 (N_2901,In_1778,In_135);
xor U2902 (N_2902,In_1586,In_720);
and U2903 (N_2903,In_1584,In_929);
or U2904 (N_2904,In_833,In_1300);
nor U2905 (N_2905,In_2282,In_110);
nor U2906 (N_2906,In_1661,In_1123);
and U2907 (N_2907,In_1061,In_1446);
and U2908 (N_2908,In_2454,In_1984);
nand U2909 (N_2909,In_1000,In_796);
or U2910 (N_2910,In_748,In_477);
nand U2911 (N_2911,In_1345,In_841);
nor U2912 (N_2912,In_601,In_2465);
and U2913 (N_2913,In_1699,In_1356);
nor U2914 (N_2914,In_2344,In_1624);
and U2915 (N_2915,In_241,In_70);
nor U2916 (N_2916,In_1838,In_1128);
xor U2917 (N_2917,In_932,In_757);
nand U2918 (N_2918,In_2470,In_997);
nor U2919 (N_2919,In_1669,In_2435);
or U2920 (N_2920,In_2372,In_1650);
nor U2921 (N_2921,In_2168,In_1855);
nand U2922 (N_2922,In_2069,In_254);
or U2923 (N_2923,In_592,In_188);
or U2924 (N_2924,In_1859,In_1909);
nor U2925 (N_2925,In_1186,In_2054);
nor U2926 (N_2926,In_2303,In_2112);
and U2927 (N_2927,In_545,In_1375);
nor U2928 (N_2928,In_99,In_2251);
nor U2929 (N_2929,In_996,In_990);
and U2930 (N_2930,In_1614,In_113);
nor U2931 (N_2931,In_2444,In_764);
or U2932 (N_2932,In_1776,In_415);
or U2933 (N_2933,In_1083,In_1654);
or U2934 (N_2934,In_43,In_1537);
nor U2935 (N_2935,In_1929,In_1478);
and U2936 (N_2936,In_1197,In_29);
nor U2937 (N_2937,In_1111,In_2316);
or U2938 (N_2938,In_2053,In_1714);
or U2939 (N_2939,In_1169,In_1773);
nand U2940 (N_2940,In_2256,In_930);
and U2941 (N_2941,In_2285,In_289);
or U2942 (N_2942,In_1508,In_7);
xor U2943 (N_2943,In_23,In_2385);
nand U2944 (N_2944,In_782,In_2359);
or U2945 (N_2945,In_32,In_2014);
nand U2946 (N_2946,In_800,In_2340);
nand U2947 (N_2947,In_248,In_1130);
nor U2948 (N_2948,In_2143,In_940);
nand U2949 (N_2949,In_2379,In_1743);
or U2950 (N_2950,In_880,In_959);
and U2951 (N_2951,In_1652,In_757);
or U2952 (N_2952,In_2341,In_322);
nand U2953 (N_2953,In_1849,In_2366);
nor U2954 (N_2954,In_1911,In_384);
nand U2955 (N_2955,In_346,In_1049);
nor U2956 (N_2956,In_1808,In_2103);
nand U2957 (N_2957,In_395,In_1687);
or U2958 (N_2958,In_1951,In_713);
and U2959 (N_2959,In_50,In_86);
nand U2960 (N_2960,In_546,In_798);
or U2961 (N_2961,In_2019,In_236);
or U2962 (N_2962,In_861,In_995);
nand U2963 (N_2963,In_863,In_1626);
nor U2964 (N_2964,In_2470,In_1181);
nor U2965 (N_2965,In_1163,In_155);
nand U2966 (N_2966,In_2248,In_1926);
and U2967 (N_2967,In_2253,In_1786);
or U2968 (N_2968,In_856,In_2159);
xnor U2969 (N_2969,In_1591,In_779);
and U2970 (N_2970,In_439,In_1475);
or U2971 (N_2971,In_874,In_1922);
xnor U2972 (N_2972,In_812,In_518);
and U2973 (N_2973,In_1576,In_1658);
nand U2974 (N_2974,In_2295,In_2425);
xor U2975 (N_2975,In_2327,In_1072);
or U2976 (N_2976,In_902,In_2236);
or U2977 (N_2977,In_907,In_338);
nand U2978 (N_2978,In_2063,In_101);
or U2979 (N_2979,In_1642,In_613);
nand U2980 (N_2980,In_1491,In_461);
xnor U2981 (N_2981,In_2137,In_1180);
or U2982 (N_2982,In_347,In_2127);
and U2983 (N_2983,In_649,In_1827);
and U2984 (N_2984,In_1814,In_935);
nand U2985 (N_2985,In_908,In_1009);
or U2986 (N_2986,In_2490,In_2281);
nor U2987 (N_2987,In_1244,In_1317);
nand U2988 (N_2988,In_1844,In_2239);
nand U2989 (N_2989,In_909,In_1687);
nor U2990 (N_2990,In_336,In_1381);
nand U2991 (N_2991,In_1208,In_949);
or U2992 (N_2992,In_776,In_479);
nand U2993 (N_2993,In_381,In_342);
or U2994 (N_2994,In_1377,In_935);
xnor U2995 (N_2995,In_399,In_1071);
nand U2996 (N_2996,In_1362,In_1348);
and U2997 (N_2997,In_1440,In_349);
xor U2998 (N_2998,In_694,In_1843);
xor U2999 (N_2999,In_675,In_2386);
nand U3000 (N_3000,In_922,In_1377);
nor U3001 (N_3001,In_1225,In_890);
nand U3002 (N_3002,In_1329,In_1372);
nor U3003 (N_3003,In_1387,In_580);
nand U3004 (N_3004,In_747,In_2207);
xor U3005 (N_3005,In_1661,In_630);
nand U3006 (N_3006,In_678,In_248);
or U3007 (N_3007,In_16,In_860);
nand U3008 (N_3008,In_1344,In_574);
nand U3009 (N_3009,In_2023,In_688);
nand U3010 (N_3010,In_520,In_277);
nand U3011 (N_3011,In_283,In_125);
or U3012 (N_3012,In_941,In_493);
nor U3013 (N_3013,In_1138,In_1814);
nand U3014 (N_3014,In_1871,In_2172);
and U3015 (N_3015,In_238,In_1636);
nand U3016 (N_3016,In_2313,In_236);
and U3017 (N_3017,In_678,In_401);
nor U3018 (N_3018,In_854,In_2112);
nor U3019 (N_3019,In_1594,In_1839);
and U3020 (N_3020,In_1757,In_2144);
and U3021 (N_3021,In_2381,In_1682);
nand U3022 (N_3022,In_303,In_915);
and U3023 (N_3023,In_963,In_1382);
xnor U3024 (N_3024,In_549,In_528);
and U3025 (N_3025,In_1443,In_2190);
nand U3026 (N_3026,In_1446,In_310);
and U3027 (N_3027,In_407,In_18);
or U3028 (N_3028,In_282,In_770);
or U3029 (N_3029,In_2447,In_1788);
nand U3030 (N_3030,In_739,In_1358);
xor U3031 (N_3031,In_934,In_276);
and U3032 (N_3032,In_739,In_669);
xnor U3033 (N_3033,In_828,In_1913);
or U3034 (N_3034,In_1802,In_1785);
or U3035 (N_3035,In_904,In_262);
nand U3036 (N_3036,In_1585,In_1413);
or U3037 (N_3037,In_2186,In_2342);
or U3038 (N_3038,In_547,In_1526);
nor U3039 (N_3039,In_735,In_1609);
and U3040 (N_3040,In_1530,In_771);
nand U3041 (N_3041,In_2116,In_1898);
nor U3042 (N_3042,In_1631,In_2134);
and U3043 (N_3043,In_2409,In_1052);
nand U3044 (N_3044,In_161,In_270);
and U3045 (N_3045,In_1267,In_47);
nor U3046 (N_3046,In_1885,In_2192);
nand U3047 (N_3047,In_1897,In_2045);
nor U3048 (N_3048,In_675,In_734);
and U3049 (N_3049,In_522,In_1127);
xor U3050 (N_3050,In_2116,In_475);
and U3051 (N_3051,In_515,In_828);
and U3052 (N_3052,In_1818,In_425);
nand U3053 (N_3053,In_1263,In_2025);
nand U3054 (N_3054,In_2425,In_2135);
nor U3055 (N_3055,In_88,In_807);
and U3056 (N_3056,In_1511,In_1701);
nor U3057 (N_3057,In_1050,In_1260);
nor U3058 (N_3058,In_1200,In_906);
and U3059 (N_3059,In_234,In_1400);
and U3060 (N_3060,In_1802,In_2176);
nand U3061 (N_3061,In_452,In_1812);
or U3062 (N_3062,In_1000,In_1034);
and U3063 (N_3063,In_2286,In_167);
and U3064 (N_3064,In_2118,In_294);
nand U3065 (N_3065,In_212,In_1683);
xnor U3066 (N_3066,In_616,In_627);
and U3067 (N_3067,In_704,In_2323);
nor U3068 (N_3068,In_2306,In_1237);
xnor U3069 (N_3069,In_1545,In_342);
nor U3070 (N_3070,In_1794,In_1357);
and U3071 (N_3071,In_794,In_1421);
nor U3072 (N_3072,In_302,In_737);
nor U3073 (N_3073,In_1913,In_1557);
nor U3074 (N_3074,In_1739,In_208);
nand U3075 (N_3075,In_1884,In_667);
nor U3076 (N_3076,In_287,In_1207);
and U3077 (N_3077,In_2070,In_2430);
and U3078 (N_3078,In_1836,In_1472);
or U3079 (N_3079,In_2456,In_2074);
nand U3080 (N_3080,In_1513,In_2288);
and U3081 (N_3081,In_252,In_1851);
nand U3082 (N_3082,In_566,In_1392);
or U3083 (N_3083,In_1319,In_2286);
xor U3084 (N_3084,In_2364,In_2423);
nor U3085 (N_3085,In_1789,In_2445);
or U3086 (N_3086,In_197,In_855);
or U3087 (N_3087,In_2375,In_2428);
and U3088 (N_3088,In_1681,In_575);
and U3089 (N_3089,In_1781,In_1584);
or U3090 (N_3090,In_1250,In_94);
nand U3091 (N_3091,In_1221,In_2250);
nand U3092 (N_3092,In_1817,In_136);
and U3093 (N_3093,In_1480,In_558);
or U3094 (N_3094,In_650,In_709);
and U3095 (N_3095,In_1639,In_831);
or U3096 (N_3096,In_779,In_2423);
nor U3097 (N_3097,In_1689,In_1152);
xor U3098 (N_3098,In_534,In_2331);
nand U3099 (N_3099,In_148,In_1346);
nor U3100 (N_3100,In_1705,In_2087);
or U3101 (N_3101,In_2019,In_914);
nor U3102 (N_3102,In_1800,In_390);
nand U3103 (N_3103,In_1322,In_2210);
nor U3104 (N_3104,In_413,In_2446);
nor U3105 (N_3105,In_1743,In_481);
xnor U3106 (N_3106,In_211,In_1975);
or U3107 (N_3107,In_1589,In_1402);
xor U3108 (N_3108,In_1901,In_2291);
or U3109 (N_3109,In_299,In_195);
or U3110 (N_3110,In_666,In_538);
and U3111 (N_3111,In_1519,In_992);
nor U3112 (N_3112,In_1878,In_1766);
xor U3113 (N_3113,In_124,In_1863);
nor U3114 (N_3114,In_2273,In_2093);
xnor U3115 (N_3115,In_24,In_2027);
and U3116 (N_3116,In_2446,In_1439);
xor U3117 (N_3117,In_2156,In_1164);
nand U3118 (N_3118,In_1535,In_1723);
nand U3119 (N_3119,In_1480,In_2390);
nor U3120 (N_3120,In_856,In_682);
xnor U3121 (N_3121,In_2313,In_2124);
nand U3122 (N_3122,In_1340,In_1664);
nor U3123 (N_3123,In_1125,In_2168);
nor U3124 (N_3124,In_1629,In_1048);
or U3125 (N_3125,N_2202,N_1998);
nor U3126 (N_3126,N_1036,N_3014);
and U3127 (N_3127,N_1699,N_1035);
and U3128 (N_3128,N_2141,N_2538);
nand U3129 (N_3129,N_1774,N_648);
nor U3130 (N_3130,N_782,N_987);
nand U3131 (N_3131,N_109,N_142);
nor U3132 (N_3132,N_3048,N_1877);
nor U3133 (N_3133,N_870,N_2783);
and U3134 (N_3134,N_1918,N_1298);
nor U3135 (N_3135,N_264,N_1082);
or U3136 (N_3136,N_1529,N_2086);
nand U3137 (N_3137,N_163,N_1907);
or U3138 (N_3138,N_2999,N_2558);
and U3139 (N_3139,N_2012,N_1491);
nand U3140 (N_3140,N_2786,N_675);
and U3141 (N_3141,N_619,N_2873);
and U3142 (N_3142,N_271,N_1812);
xor U3143 (N_3143,N_2603,N_2859);
nand U3144 (N_3144,N_510,N_2038);
nor U3145 (N_3145,N_2888,N_2456);
or U3146 (N_3146,N_465,N_1126);
nand U3147 (N_3147,N_2741,N_371);
nand U3148 (N_3148,N_1144,N_2486);
and U3149 (N_3149,N_2687,N_18);
and U3150 (N_3150,N_1233,N_2890);
or U3151 (N_3151,N_35,N_2542);
nor U3152 (N_3152,N_1198,N_550);
and U3153 (N_3153,N_96,N_1706);
or U3154 (N_3154,N_2454,N_2482);
nor U3155 (N_3155,N_1408,N_962);
nor U3156 (N_3156,N_2507,N_2588);
nor U3157 (N_3157,N_165,N_2501);
xnor U3158 (N_3158,N_1927,N_1091);
and U3159 (N_3159,N_1637,N_3111);
nand U3160 (N_3160,N_356,N_1281);
nor U3161 (N_3161,N_1440,N_765);
and U3162 (N_3162,N_1331,N_429);
and U3163 (N_3163,N_71,N_800);
nor U3164 (N_3164,N_2157,N_663);
nand U3165 (N_3165,N_2282,N_2685);
or U3166 (N_3166,N_3033,N_1345);
or U3167 (N_3167,N_1869,N_2830);
or U3168 (N_3168,N_1382,N_1761);
nor U3169 (N_3169,N_1027,N_585);
nor U3170 (N_3170,N_1279,N_1465);
and U3171 (N_3171,N_2137,N_1937);
nor U3172 (N_3172,N_923,N_353);
or U3173 (N_3173,N_2314,N_2630);
or U3174 (N_3174,N_769,N_87);
nor U3175 (N_3175,N_3116,N_2054);
and U3176 (N_3176,N_2793,N_1575);
nand U3177 (N_3177,N_416,N_1950);
nor U3178 (N_3178,N_2616,N_1643);
nor U3179 (N_3179,N_1501,N_1486);
nand U3180 (N_3180,N_1583,N_1219);
and U3181 (N_3181,N_1939,N_1202);
nand U3182 (N_3182,N_2697,N_967);
nor U3183 (N_3183,N_2495,N_1217);
nor U3184 (N_3184,N_976,N_2342);
or U3185 (N_3185,N_583,N_2122);
nand U3186 (N_3186,N_334,N_2695);
nor U3187 (N_3187,N_1289,N_1482);
nand U3188 (N_3188,N_1243,N_2908);
xor U3189 (N_3189,N_3057,N_2654);
nor U3190 (N_3190,N_1825,N_956);
nor U3191 (N_3191,N_827,N_1444);
xor U3192 (N_3192,N_986,N_887);
nand U3193 (N_3193,N_1152,N_3124);
nor U3194 (N_3194,N_1291,N_843);
or U3195 (N_3195,N_674,N_1053);
and U3196 (N_3196,N_1627,N_2100);
xnor U3197 (N_3197,N_2795,N_2307);
or U3198 (N_3198,N_403,N_983);
nand U3199 (N_3199,N_1320,N_2528);
nand U3200 (N_3200,N_2945,N_667);
or U3201 (N_3201,N_588,N_1962);
xor U3202 (N_3202,N_2647,N_2133);
nor U3203 (N_3203,N_2306,N_32);
nand U3204 (N_3204,N_1128,N_1958);
or U3205 (N_3205,N_640,N_662);
and U3206 (N_3206,N_367,N_1665);
nand U3207 (N_3207,N_422,N_305);
or U3208 (N_3208,N_1608,N_941);
and U3209 (N_3209,N_512,N_1725);
nand U3210 (N_3210,N_1018,N_2714);
or U3211 (N_3211,N_1957,N_1159);
and U3212 (N_3212,N_826,N_2977);
and U3213 (N_3213,N_2920,N_2554);
and U3214 (N_3214,N_2042,N_735);
or U3215 (N_3215,N_2485,N_1125);
or U3216 (N_3216,N_485,N_3021);
nand U3217 (N_3217,N_2595,N_424);
and U3218 (N_3218,N_393,N_2023);
nand U3219 (N_3219,N_2121,N_131);
and U3220 (N_3220,N_2621,N_1337);
xnor U3221 (N_3221,N_2994,N_20);
and U3222 (N_3222,N_2826,N_2511);
or U3223 (N_3223,N_379,N_1271);
nor U3224 (N_3224,N_212,N_1141);
nor U3225 (N_3225,N_2798,N_1696);
xnor U3226 (N_3226,N_2426,N_2164);
nor U3227 (N_3227,N_2268,N_281);
nand U3228 (N_3228,N_2709,N_2794);
and U3229 (N_3229,N_2104,N_1364);
nor U3230 (N_3230,N_534,N_2912);
or U3231 (N_3231,N_920,N_1876);
and U3232 (N_3232,N_1682,N_338);
and U3233 (N_3233,N_1068,N_1329);
nor U3234 (N_3234,N_1565,N_196);
or U3235 (N_3235,N_2313,N_3080);
xor U3236 (N_3236,N_1509,N_2563);
nand U3237 (N_3237,N_1742,N_721);
nor U3238 (N_3238,N_1312,N_1722);
nor U3239 (N_3239,N_2990,N_2686);
or U3240 (N_3240,N_1392,N_1859);
nor U3241 (N_3241,N_1799,N_1296);
and U3242 (N_3242,N_2645,N_1433);
xor U3243 (N_3243,N_2058,N_1878);
nand U3244 (N_3244,N_2158,N_3056);
or U3245 (N_3245,N_2875,N_2403);
or U3246 (N_3246,N_1506,N_2636);
nor U3247 (N_3247,N_1210,N_2612);
and U3248 (N_3248,N_1779,N_405);
or U3249 (N_3249,N_1387,N_756);
and U3250 (N_3250,N_1758,N_1083);
and U3251 (N_3251,N_780,N_3004);
nor U3252 (N_3252,N_2478,N_489);
or U3253 (N_3253,N_3105,N_2672);
and U3254 (N_3254,N_1545,N_637);
nor U3255 (N_3255,N_3018,N_797);
nand U3256 (N_3256,N_1819,N_2127);
or U3257 (N_3257,N_3019,N_838);
xor U3258 (N_3258,N_844,N_1528);
nand U3259 (N_3259,N_2767,N_1460);
nor U3260 (N_3260,N_666,N_939);
and U3261 (N_3261,N_1169,N_208);
nand U3262 (N_3262,N_2573,N_2441);
or U3263 (N_3263,N_1882,N_308);
nor U3264 (N_3264,N_566,N_1335);
and U3265 (N_3265,N_1822,N_2919);
and U3266 (N_3266,N_355,N_1395);
nand U3267 (N_3267,N_1349,N_387);
nor U3268 (N_3268,N_1838,N_2224);
nand U3269 (N_3269,N_1259,N_1639);
or U3270 (N_3270,N_2231,N_238);
or U3271 (N_3271,N_350,N_2862);
xor U3272 (N_3272,N_1375,N_612);
or U3273 (N_3273,N_850,N_2723);
or U3274 (N_3274,N_1749,N_524);
or U3275 (N_3275,N_600,N_2349);
or U3276 (N_3276,N_85,N_1928);
and U3277 (N_3277,N_1798,N_712);
nand U3278 (N_3278,N_460,N_2229);
and U3279 (N_3279,N_2463,N_2174);
nand U3280 (N_3280,N_1192,N_2619);
nor U3281 (N_3281,N_310,N_636);
and U3282 (N_3282,N_2173,N_1393);
and U3283 (N_3283,N_2740,N_177);
nand U3284 (N_3284,N_15,N_1979);
and U3285 (N_3285,N_645,N_412);
xor U3286 (N_3286,N_300,N_2059);
or U3287 (N_3287,N_2763,N_2145);
and U3288 (N_3288,N_660,N_895);
nor U3289 (N_3289,N_1225,N_1666);
or U3290 (N_3290,N_1771,N_1974);
and U3291 (N_3291,N_1427,N_1121);
nor U3292 (N_3292,N_2123,N_346);
nand U3293 (N_3293,N_1969,N_1114);
nand U3294 (N_3294,N_1929,N_2604);
nand U3295 (N_3295,N_810,N_622);
nand U3296 (N_3296,N_579,N_4);
or U3297 (N_3297,N_1865,N_3071);
xnor U3298 (N_3298,N_2351,N_1924);
or U3299 (N_3299,N_761,N_2188);
or U3300 (N_3300,N_14,N_876);
xnor U3301 (N_3301,N_2562,N_2390);
xor U3302 (N_3302,N_1112,N_2101);
nand U3303 (N_3303,N_269,N_78);
nor U3304 (N_3304,N_2671,N_1542);
nand U3305 (N_3305,N_625,N_2730);
and U3306 (N_3306,N_2379,N_2570);
and U3307 (N_3307,N_2545,N_2503);
and U3308 (N_3308,N_1785,N_2263);
nor U3309 (N_3309,N_917,N_2816);
and U3310 (N_3310,N_807,N_542);
nor U3311 (N_3311,N_2972,N_1881);
and U3312 (N_3312,N_2978,N_318);
or U3313 (N_3313,N_2075,N_2450);
or U3314 (N_3314,N_1885,N_2009);
or U3315 (N_3315,N_2957,N_1668);
and U3316 (N_3316,N_2874,N_999);
and U3317 (N_3317,N_2365,N_1959);
nand U3318 (N_3318,N_2013,N_1441);
nor U3319 (N_3319,N_2240,N_938);
nand U3320 (N_3320,N_1490,N_1373);
nor U3321 (N_3321,N_1805,N_746);
or U3322 (N_3322,N_2370,N_997);
nand U3323 (N_3323,N_1580,N_651);
nand U3324 (N_3324,N_1138,N_2460);
nor U3325 (N_3325,N_1989,N_2722);
and U3326 (N_3326,N_53,N_124);
xnor U3327 (N_3327,N_3054,N_49);
nand U3328 (N_3328,N_587,N_2696);
or U3329 (N_3329,N_207,N_2850);
nand U3330 (N_3330,N_908,N_955);
and U3331 (N_3331,N_2219,N_1710);
nor U3332 (N_3332,N_482,N_1793);
and U3333 (N_3333,N_842,N_785);
or U3334 (N_3334,N_2377,N_2284);
nor U3335 (N_3335,N_573,N_869);
or U3336 (N_3336,N_2489,N_1512);
nand U3337 (N_3337,N_2781,N_1504);
or U3338 (N_3338,N_2475,N_2768);
and U3339 (N_3339,N_339,N_507);
nand U3340 (N_3340,N_753,N_1860);
nand U3341 (N_3341,N_247,N_2677);
xnor U3342 (N_3342,N_2857,N_2796);
and U3343 (N_3343,N_900,N_252);
or U3344 (N_3344,N_476,N_1892);
nor U3345 (N_3345,N_2238,N_3015);
and U3346 (N_3346,N_720,N_751);
nor U3347 (N_3347,N_2962,N_179);
or U3348 (N_3348,N_816,N_11);
nor U3349 (N_3349,N_1731,N_243);
nand U3350 (N_3350,N_1237,N_224);
and U3351 (N_3351,N_186,N_303);
and U3352 (N_3352,N_855,N_1644);
and U3353 (N_3353,N_457,N_1658);
and U3354 (N_3354,N_2119,N_2464);
and U3355 (N_3355,N_3008,N_1535);
or U3356 (N_3356,N_1116,N_1341);
nand U3357 (N_3357,N_220,N_3087);
nand U3358 (N_3358,N_945,N_2405);
or U3359 (N_3359,N_1350,N_1980);
xor U3360 (N_3360,N_2431,N_2543);
and U3361 (N_3361,N_1708,N_2419);
nor U3362 (N_3362,N_2439,N_2466);
or U3363 (N_3363,N_1617,N_1283);
and U3364 (N_3364,N_3108,N_2887);
or U3365 (N_3365,N_2402,N_1046);
or U3366 (N_3366,N_661,N_453);
or U3367 (N_3367,N_1163,N_1479);
nand U3368 (N_3368,N_584,N_1244);
and U3369 (N_3369,N_2675,N_2948);
nor U3370 (N_3370,N_1469,N_1503);
and U3371 (N_3371,N_1613,N_787);
or U3372 (N_3372,N_2773,N_1661);
or U3373 (N_3373,N_1925,N_2869);
or U3374 (N_3374,N_2320,N_1518);
nand U3375 (N_3375,N_894,N_2928);
nand U3376 (N_3376,N_2183,N_2579);
or U3377 (N_3377,N_123,N_912);
xor U3378 (N_3378,N_1883,N_2981);
and U3379 (N_3379,N_1587,N_503);
nand U3380 (N_3380,N_2970,N_1931);
nand U3381 (N_3381,N_2148,N_1737);
and U3382 (N_3382,N_319,N_3032);
and U3383 (N_3383,N_1578,N_312);
and U3384 (N_3384,N_2032,N_691);
and U3385 (N_3385,N_2373,N_1673);
or U3386 (N_3386,N_1450,N_169);
xnor U3387 (N_3387,N_2331,N_969);
and U3388 (N_3388,N_2517,N_2924);
nand U3389 (N_3389,N_2611,N_69);
nor U3390 (N_3390,N_1589,N_1972);
nand U3391 (N_3391,N_255,N_569);
nor U3392 (N_3392,N_2641,N_182);
nor U3393 (N_3393,N_1239,N_815);
nor U3394 (N_3394,N_2291,N_2536);
and U3395 (N_3395,N_62,N_1407);
and U3396 (N_3396,N_157,N_809);
and U3397 (N_3397,N_597,N_1261);
nand U3398 (N_3398,N_2213,N_1327);
or U3399 (N_3399,N_1355,N_1852);
nor U3400 (N_3400,N_135,N_9);
nor U3401 (N_3401,N_398,N_2323);
or U3402 (N_3402,N_2532,N_1769);
nand U3403 (N_3403,N_1703,N_1054);
or U3404 (N_3404,N_2077,N_2876);
nand U3405 (N_3405,N_1520,N_1476);
nor U3406 (N_3406,N_358,N_1858);
xnor U3407 (N_3407,N_3079,N_369);
nand U3408 (N_3408,N_729,N_802);
nand U3409 (N_3409,N_1926,N_1412);
nand U3410 (N_3410,N_1532,N_2860);
nor U3411 (N_3411,N_1790,N_642);
nor U3412 (N_3412,N_91,N_1338);
nor U3413 (N_3413,N_877,N_1629);
and U3414 (N_3414,N_1674,N_3012);
or U3415 (N_3415,N_1898,N_1357);
or U3416 (N_3416,N_1896,N_1763);
or U3417 (N_3417,N_2849,N_154);
or U3418 (N_3418,N_977,N_3102);
and U3419 (N_3419,N_345,N_927);
nand U3420 (N_3420,N_251,N_2176);
nand U3421 (N_3421,N_392,N_909);
nor U3422 (N_3422,N_994,N_490);
nand U3423 (N_3423,N_1832,N_3044);
or U3424 (N_3424,N_933,N_187);
nand U3425 (N_3425,N_1249,N_1577);
nand U3426 (N_3426,N_3119,N_794);
nand U3427 (N_3427,N_1568,N_1816);
nor U3428 (N_3428,N_2983,N_391);
nor U3429 (N_3429,N_30,N_2084);
xor U3430 (N_3430,N_530,N_1889);
nor U3431 (N_3431,N_513,N_1086);
nor U3432 (N_3432,N_2249,N_960);
xor U3433 (N_3433,N_134,N_1754);
and U3434 (N_3434,N_2694,N_2670);
nand U3435 (N_3435,N_2982,N_684);
xor U3436 (N_3436,N_1492,N_2046);
nand U3437 (N_3437,N_1258,N_2693);
or U3438 (N_3438,N_624,N_296);
nor U3439 (N_3439,N_3059,N_589);
nor U3440 (N_3440,N_2893,N_2234);
and U3441 (N_3441,N_2170,N_620);
and U3442 (N_3442,N_1455,N_1093);
nor U3443 (N_3443,N_285,N_1628);
and U3444 (N_3444,N_2810,N_1085);
or U3445 (N_3445,N_2348,N_1826);
nor U3446 (N_3446,N_2292,N_1765);
or U3447 (N_3447,N_253,N_1488);
and U3448 (N_3448,N_790,N_162);
nor U3449 (N_3449,N_357,N_1140);
or U3450 (N_3450,N_2669,N_2867);
nor U3451 (N_3451,N_1034,N_435);
and U3452 (N_3452,N_3035,N_3020);
nor U3453 (N_3453,N_1630,N_2060);
and U3454 (N_3454,N_3022,N_2625);
nor U3455 (N_3455,N_2879,N_420);
nand U3456 (N_3456,N_2580,N_2410);
xor U3457 (N_3457,N_1307,N_1599);
or U3458 (N_3458,N_570,N_2905);
nand U3459 (N_3459,N_1257,N_2550);
xnor U3460 (N_3460,N_1415,N_2939);
or U3461 (N_3461,N_284,N_1318);
nor U3462 (N_3462,N_1794,N_1031);
nand U3463 (N_3463,N_3074,N_2040);
or U3464 (N_3464,N_2846,N_1756);
nor U3465 (N_3465,N_1836,N_1485);
nor U3466 (N_3466,N_190,N_2615);
or U3467 (N_3467,N_2502,N_993);
nor U3468 (N_3468,N_2295,N_2169);
nor U3469 (N_3469,N_953,N_1453);
nor U3470 (N_3470,N_348,N_2780);
xor U3471 (N_3471,N_1134,N_2836);
xnor U3472 (N_3472,N_2565,N_1097);
nor U3473 (N_3473,N_1181,N_1348);
nand U3474 (N_3474,N_828,N_385);
nand U3475 (N_3475,N_258,N_1514);
and U3476 (N_3476,N_498,N_957);
nor U3477 (N_3477,N_652,N_1536);
and U3478 (N_3478,N_892,N_884);
nand U3479 (N_3479,N_1078,N_1207);
and U3480 (N_3480,N_916,N_1151);
nand U3481 (N_3481,N_647,N_1796);
nor U3482 (N_3482,N_2056,N_2681);
and U3483 (N_3483,N_2590,N_153);
xor U3484 (N_3484,N_1426,N_2117);
and U3485 (N_3485,N_493,N_1378);
nand U3486 (N_3486,N_329,N_2290);
nand U3487 (N_3487,N_383,N_2082);
nand U3488 (N_3488,N_2979,N_1124);
nor U3489 (N_3489,N_2750,N_1901);
and U3490 (N_3490,N_919,N_825);
and U3491 (N_3491,N_1588,N_1362);
nor U3492 (N_3492,N_742,N_270);
nor U3493 (N_3493,N_2500,N_140);
xnor U3494 (N_3494,N_1561,N_1061);
nor U3495 (N_3495,N_1922,N_1439);
and U3496 (N_3496,N_1005,N_2333);
nand U3497 (N_3497,N_2966,N_38);
nor U3498 (N_3498,N_1315,N_1548);
and U3499 (N_3499,N_2746,N_1938);
or U3500 (N_3500,N_2943,N_1397);
nand U3501 (N_3501,N_2281,N_2334);
and U3502 (N_3502,N_1640,N_1325);
nor U3503 (N_3503,N_2775,N_2468);
nor U3504 (N_3504,N_1302,N_536);
and U3505 (N_3505,N_591,N_1970);
nand U3506 (N_3506,N_664,N_2253);
and U3507 (N_3507,N_1176,N_1303);
nand U3508 (N_3508,N_2518,N_781);
or U3509 (N_3509,N_1420,N_226);
nand U3510 (N_3510,N_128,N_1968);
nand U3511 (N_3511,N_560,N_2574);
and U3512 (N_3512,N_671,N_1986);
nor U3513 (N_3513,N_322,N_822);
and U3514 (N_3514,N_829,N_1321);
or U3515 (N_3515,N_1234,N_132);
nor U3516 (N_3516,N_1723,N_839);
and U3517 (N_3517,N_2657,N_2577);
xnor U3518 (N_3518,N_2318,N_295);
nand U3519 (N_3519,N_1023,N_1619);
nor U3520 (N_3520,N_1156,N_2041);
nand U3521 (N_3521,N_514,N_861);
or U3522 (N_3522,N_1508,N_1157);
nor U3523 (N_3523,N_963,N_1032);
nor U3524 (N_3524,N_791,N_2124);
nor U3525 (N_3525,N_479,N_321);
nand U3526 (N_3526,N_95,N_3122);
or U3527 (N_3527,N_3112,N_1543);
or U3528 (N_3528,N_679,N_1359);
or U3529 (N_3529,N_1811,N_2302);
or U3530 (N_3530,N_1983,N_1055);
or U3531 (N_3531,N_2713,N_227);
and U3532 (N_3532,N_2438,N_2043);
nor U3533 (N_3533,N_2265,N_1960);
nand U3534 (N_3534,N_408,N_2343);
and U3535 (N_3535,N_2092,N_1458);
or U3536 (N_3536,N_1778,N_2522);
nor U3537 (N_3537,N_2700,N_1119);
or U3538 (N_3538,N_2422,N_101);
nand U3539 (N_3539,N_1245,N_2338);
nand U3540 (N_3540,N_2347,N_2413);
xnor U3541 (N_3541,N_1523,N_946);
nand U3542 (N_3542,N_2428,N_1484);
nand U3543 (N_3543,N_1719,N_120);
nand U3544 (N_3544,N_2147,N_2594);
nor U3545 (N_3545,N_1007,N_37);
and U3546 (N_3546,N_1709,N_1946);
nand U3547 (N_3547,N_2510,N_1065);
xnor U3548 (N_3548,N_2701,N_2653);
and U3549 (N_3549,N_2764,N_1012);
xor U3550 (N_3550,N_1704,N_1224);
nor U3551 (N_3551,N_508,N_1902);
nand U3552 (N_3552,N_635,N_1319);
nor U3553 (N_3553,N_2725,N_1419);
or U3554 (N_3554,N_2684,N_1870);
and U3555 (N_3555,N_3070,N_351);
nor U3556 (N_3556,N_174,N_2787);
or U3557 (N_3557,N_747,N_696);
nand U3558 (N_3558,N_2223,N_978);
nand U3559 (N_3559,N_1166,N_421);
nand U3560 (N_3560,N_1042,N_856);
nand U3561 (N_3561,N_1810,N_1801);
xnor U3562 (N_3562,N_2633,N_404);
nor U3563 (N_3563,N_914,N_3093);
nor U3564 (N_3564,N_1004,N_2132);
nor U3565 (N_3565,N_2901,N_2804);
or U3566 (N_3566,N_2973,N_1846);
nand U3567 (N_3567,N_1391,N_2896);
xor U3568 (N_3568,N_817,N_849);
xnor U3569 (N_3569,N_2418,N_488);
nor U3570 (N_3570,N_2656,N_2311);
or U3571 (N_3571,N_2028,N_2726);
and U3572 (N_3572,N_2854,N_3043);
xnor U3573 (N_3573,N_2553,N_107);
xor U3574 (N_3574,N_3072,N_288);
or U3575 (N_3575,N_2790,N_1275);
xnor U3576 (N_3576,N_2584,N_67);
nand U3577 (N_3577,N_2776,N_80);
nor U3578 (N_3578,N_328,N_2534);
or U3579 (N_3579,N_763,N_1873);
and U3580 (N_3580,N_2716,N_559);
or U3581 (N_3581,N_122,N_2880);
and U3582 (N_3582,N_905,N_1449);
or U3583 (N_3583,N_36,N_26);
or U3584 (N_3584,N_1084,N_409);
and U3585 (N_3585,N_2165,N_1788);
and U3586 (N_3586,N_3101,N_362);
or U3587 (N_3587,N_678,N_2476);
and U3588 (N_3588,N_2704,N_236);
and U3589 (N_3589,N_2254,N_1573);
xnor U3590 (N_3590,N_2541,N_518);
and U3591 (N_3591,N_2585,N_2600);
and U3592 (N_3592,N_3016,N_1333);
and U3593 (N_3593,N_924,N_854);
and U3594 (N_3594,N_244,N_2239);
or U3595 (N_3595,N_1604,N_1747);
or U3596 (N_3596,N_3065,N_868);
nor U3597 (N_3597,N_1659,N_1818);
xor U3598 (N_3598,N_1416,N_948);
and U3599 (N_3599,N_2627,N_1999);
or U3600 (N_3600,N_2710,N_2527);
nor U3601 (N_3601,N_1975,N_1728);
or U3602 (N_3602,N_741,N_1300);
nor U3603 (N_3603,N_2797,N_1933);
nor U3604 (N_3604,N_1821,N_616);
nand U3605 (N_3605,N_1934,N_673);
nand U3606 (N_3606,N_1967,N_1530);
nor U3607 (N_3607,N_2088,N_1429);
and U3608 (N_3608,N_2420,N_164);
or U3609 (N_3609,N_384,N_882);
and U3610 (N_3610,N_256,N_755);
nor U3611 (N_3611,N_525,N_52);
nand U3612 (N_3612,N_2734,N_1286);
and U3613 (N_3613,N_2415,N_1605);
or U3614 (N_3614,N_3040,N_2113);
nand U3615 (N_3615,N_158,N_1853);
xnor U3616 (N_3616,N_2705,N_118);
or U3617 (N_3617,N_2206,N_1063);
and U3618 (N_3618,N_1526,N_6);
and U3619 (N_3619,N_2991,N_2564);
or U3620 (N_3620,N_1009,N_1517);
and U3621 (N_3621,N_221,N_1274);
nand U3622 (N_3622,N_2679,N_3064);
nor U3623 (N_3623,N_2557,N_970);
xnor U3624 (N_3624,N_2451,N_21);
xor U3625 (N_3625,N_2001,N_237);
nand U3626 (N_3626,N_2017,N_1230);
or U3627 (N_3627,N_1278,N_2965);
and U3628 (N_3628,N_3,N_2276);
xnor U3629 (N_3629,N_239,N_2895);
or U3630 (N_3630,N_3005,N_659);
and U3631 (N_3631,N_1358,N_2822);
or U3632 (N_3632,N_1657,N_1712);
and U3633 (N_3633,N_2863,N_2483);
or U3634 (N_3634,N_442,N_930);
nand U3635 (N_3635,N_672,N_1209);
nand U3636 (N_3636,N_793,N_1477);
xor U3637 (N_3637,N_1354,N_1011);
nor U3638 (N_3638,N_2256,N_2014);
or U3639 (N_3639,N_297,N_293);
nand U3640 (N_3640,N_2387,N_2073);
or U3641 (N_3641,N_366,N_1591);
or U3642 (N_3642,N_2057,N_1648);
and U3643 (N_3643,N_2886,N_2555);
and U3644 (N_3644,N_1687,N_299);
or U3645 (N_3645,N_497,N_1863);
and U3646 (N_3646,N_744,N_495);
nor U3647 (N_3647,N_125,N_337);
and U3648 (N_3648,N_3029,N_115);
and U3649 (N_3649,N_904,N_1172);
and U3650 (N_3650,N_148,N_2091);
nor U3651 (N_3651,N_1976,N_2252);
and U3652 (N_3652,N_455,N_835);
nand U3653 (N_3653,N_1229,N_3025);
nor U3654 (N_3654,N_878,N_1050);
nand U3655 (N_3655,N_2280,N_733);
nor U3656 (N_3656,N_1273,N_2751);
or U3657 (N_3657,N_499,N_2242);
nand U3658 (N_3658,N_436,N_2884);
and U3659 (N_3659,N_1150,N_935);
or U3660 (N_3660,N_2984,N_2194);
xnor U3661 (N_3661,N_1301,N_1100);
nor U3662 (N_3662,N_1381,N_81);
nor U3663 (N_3663,N_2138,N_394);
and U3664 (N_3664,N_1498,N_1655);
or U3665 (N_3665,N_2275,N_1475);
or U3666 (N_3666,N_2356,N_1363);
or U3667 (N_3667,N_2397,N_417);
or U3668 (N_3668,N_160,N_2539);
nor U3669 (N_3669,N_267,N_1705);
nor U3670 (N_3670,N_2868,N_972);
and U3671 (N_3671,N_658,N_2791);
or U3672 (N_3672,N_1505,N_988);
nor U3673 (N_3673,N_1947,N_275);
and U3674 (N_3674,N_194,N_491);
and U3675 (N_3675,N_565,N_2903);
and U3676 (N_3676,N_3117,N_2599);
or U3677 (N_3677,N_1594,N_159);
nor U3678 (N_3678,N_2181,N_2809);
xnor U3679 (N_3679,N_2332,N_76);
nand U3680 (N_3680,N_2159,N_803);
or U3681 (N_3681,N_400,N_1624);
and U3682 (N_3682,N_1507,N_2782);
and U3683 (N_3683,N_981,N_1132);
and U3684 (N_3684,N_1955,N_1917);
nor U3685 (N_3685,N_758,N_2907);
xnor U3686 (N_3686,N_1915,N_554);
and U3687 (N_3687,N_738,N_1784);
and U3688 (N_3688,N_1267,N_2506);
xnor U3689 (N_3689,N_2108,N_851);
xor U3690 (N_3690,N_2769,N_2922);
nor U3691 (N_3691,N_2412,N_496);
nor U3692 (N_3692,N_2462,N_2733);
nand U3693 (N_3693,N_2208,N_764);
nand U3694 (N_3694,N_2407,N_2182);
nand U3695 (N_3695,N_2095,N_1135);
nor U3696 (N_3696,N_246,N_217);
or U3697 (N_3697,N_2301,N_2525);
or U3698 (N_3698,N_2904,N_2537);
nor U3699 (N_3699,N_1493,N_1480);
or U3700 (N_3700,N_1732,N_2029);
and U3701 (N_3701,N_2358,N_180);
nor U3702 (N_3702,N_832,N_2891);
or U3703 (N_3703,N_2271,N_2247);
xor U3704 (N_3704,N_1956,N_191);
or U3705 (N_3705,N_1070,N_1746);
xor U3706 (N_3706,N_1435,N_2861);
nor U3707 (N_3707,N_423,N_1149);
or U3708 (N_3708,N_438,N_2617);
and U3709 (N_3709,N_215,N_64);
xor U3710 (N_3710,N_1410,N_2216);
or U3711 (N_3711,N_344,N_1843);
or U3712 (N_3712,N_1603,N_759);
and U3713 (N_3713,N_1139,N_860);
nand U3714 (N_3714,N_1894,N_79);
nor U3715 (N_3715,N_188,N_1936);
nand U3716 (N_3716,N_2967,N_2380);
nor U3717 (N_3717,N_2207,N_2597);
or U3718 (N_3718,N_1932,N_43);
and U3719 (N_3719,N_2309,N_2021);
nor U3720 (N_3720,N_1193,N_2404);
nand U3721 (N_3721,N_2424,N_2640);
nor U3722 (N_3722,N_991,N_2909);
xnor U3723 (N_3723,N_2792,N_2218);
nor U3724 (N_3724,N_964,N_961);
xor U3725 (N_3725,N_2067,N_902);
nand U3726 (N_3726,N_1802,N_2136);
xor U3727 (N_3727,N_2228,N_2166);
nand U3728 (N_3728,N_2107,N_1040);
or U3729 (N_3729,N_2666,N_2414);
and U3730 (N_3730,N_519,N_760);
or U3731 (N_3731,N_1823,N_452);
or U3732 (N_3732,N_707,N_33);
nand U3733 (N_3733,N_1871,N_1422);
or U3734 (N_3734,N_1459,N_1595);
or U3735 (N_3735,N_1308,N_2639);
nand U3736 (N_3736,N_2526,N_562);
xor U3737 (N_3737,N_543,N_1766);
xnor U3738 (N_3738,N_1146,N_10);
and U3739 (N_3739,N_2858,N_748);
and U3740 (N_3740,N_1344,N_1949);
or U3741 (N_3741,N_3046,N_1733);
nor U3742 (N_3742,N_1328,N_2447);
and U3743 (N_3743,N_2085,N_1494);
nand U3744 (N_3744,N_1633,N_229);
or U3745 (N_3745,N_1201,N_2568);
or U3746 (N_3746,N_2698,N_1777);
nand U3747 (N_3747,N_506,N_1768);
nand U3748 (N_3748,N_2139,N_2593);
or U3749 (N_3749,N_50,N_548);
and U3750 (N_3750,N_1092,N_1284);
xor U3751 (N_3751,N_2448,N_1531);
nand U3752 (N_3752,N_2820,N_2774);
nor U3753 (N_3753,N_1045,N_2772);
or U3754 (N_3754,N_2759,N_2423);
and U3755 (N_3755,N_509,N_897);
or U3756 (N_3756,N_1880,N_2878);
or U3757 (N_3757,N_1681,N_2551);
and U3758 (N_3758,N_55,N_1569);
nor U3759 (N_3759,N_697,N_2575);
nor U3760 (N_3760,N_555,N_1194);
nor U3761 (N_3761,N_1370,N_1017);
and U3762 (N_3762,N_596,N_2490);
and U3763 (N_3763,N_2461,N_541);
nand U3764 (N_3764,N_349,N_2864);
nand U3765 (N_3765,N_2718,N_1642);
xnor U3766 (N_3766,N_1596,N_156);
and U3767 (N_3767,N_286,N_151);
nor U3768 (N_3768,N_680,N_74);
nor U3769 (N_3769,N_200,N_1002);
xnor U3770 (N_3770,N_1781,N_2329);
nand U3771 (N_3771,N_2834,N_1848);
or U3772 (N_3772,N_413,N_257);
or U3773 (N_3773,N_688,N_1203);
or U3774 (N_3774,N_1096,N_2156);
nand U3775 (N_3775,N_1891,N_204);
and U3776 (N_3776,N_2788,N_921);
and U3777 (N_3777,N_396,N_2492);
and U3778 (N_3778,N_1432,N_2071);
and U3779 (N_3779,N_695,N_2923);
or U3780 (N_3780,N_1671,N_677);
and U3781 (N_3781,N_1714,N_2634);
xnor U3782 (N_3782,N_1844,N_2189);
nand U3783 (N_3783,N_2708,N_599);
and U3784 (N_3784,N_1824,N_805);
xnor U3785 (N_3785,N_2484,N_2736);
or U3786 (N_3786,N_633,N_419);
nor U3787 (N_3787,N_3083,N_336);
nand U3788 (N_3788,N_2559,N_3118);
or U3789 (N_3789,N_657,N_1621);
nand U3790 (N_3790,N_2739,N_2312);
nand U3791 (N_3791,N_2472,N_539);
or U3792 (N_3792,N_487,N_136);
nand U3793 (N_3793,N_189,N_1102);
or U3794 (N_3794,N_1767,N_1043);
nor U3795 (N_3795,N_1782,N_98);
or U3796 (N_3796,N_397,N_399);
nor U3797 (N_3797,N_511,N_2011);
nor U3798 (N_3798,N_515,N_470);
xor U3799 (N_3799,N_54,N_3024);
nand U3800 (N_3800,N_1456,N_365);
xnor U3801 (N_3801,N_1553,N_1951);
or U3802 (N_3802,N_1692,N_1840);
or U3803 (N_3803,N_359,N_2264);
nor U3804 (N_3804,N_3096,N_2098);
nand U3805 (N_3805,N_434,N_3013);
and U3806 (N_3806,N_99,N_84);
nand U3807 (N_3807,N_2996,N_3042);
xnor U3808 (N_3808,N_2246,N_1987);
or U3809 (N_3809,N_1606,N_1470);
or U3810 (N_3810,N_1616,N_2146);
and U3811 (N_3811,N_494,N_2063);
nor U3812 (N_3812,N_990,N_1813);
xor U3813 (N_3813,N_965,N_1697);
or U3814 (N_3814,N_335,N_1544);
and U3815 (N_3815,N_57,N_72);
and U3816 (N_3816,N_1248,N_1047);
nand U3817 (N_3817,N_1973,N_911);
and U3818 (N_3818,N_2480,N_2659);
xnor U3819 (N_3819,N_2497,N_1849);
or U3820 (N_3820,N_610,N_2355);
nand U3821 (N_3821,N_481,N_47);
nand U3822 (N_3822,N_181,N_2933);
or U3823 (N_3823,N_1253,N_1690);
nand U3824 (N_3824,N_708,N_1294);
nand U3825 (N_3825,N_1037,N_1421);
and U3826 (N_3826,N_75,N_2993);
nor U3827 (N_3827,N_343,N_1576);
nand U3828 (N_3828,N_3121,N_1414);
nand U3829 (N_3829,N_852,N_1966);
nor U3830 (N_3830,N_2825,N_2549);
nor U3831 (N_3831,N_1991,N_263);
and U3832 (N_3832,N_2843,N_1164);
and U3833 (N_3833,N_628,N_2524);
nand U3834 (N_3834,N_1436,N_2350);
nor U3835 (N_3835,N_2221,N_1762);
nor U3836 (N_3836,N_1607,N_725);
nor U3837 (N_3837,N_3090,N_2523);
xor U3838 (N_3838,N_240,N_2727);
nor U3839 (N_3839,N_1527,N_51);
or U3840 (N_3840,N_324,N_2203);
nor U3841 (N_3841,N_1402,N_1855);
nor U3842 (N_3842,N_1610,N_3114);
xnor U3843 (N_3843,N_1347,N_1067);
nor U3844 (N_3844,N_2703,N_608);
nor U3845 (N_3845,N_598,N_2015);
nand U3846 (N_3846,N_2031,N_433);
and U3847 (N_3847,N_1446,N_896);
and U3848 (N_3848,N_12,N_2328);
nand U3849 (N_3849,N_595,N_2187);
xnor U3850 (N_3850,N_1242,N_646);
nor U3851 (N_3851,N_527,N_2737);
nand U3852 (N_3852,N_390,N_311);
nor U3853 (N_3853,N_2959,N_2711);
nand U3854 (N_3854,N_232,N_1772);
or U3855 (N_3855,N_1272,N_1374);
xnor U3856 (N_3856,N_291,N_2465);
or U3857 (N_3857,N_1467,N_2);
or U3858 (N_3858,N_2479,N_1222);
xnor U3859 (N_3859,N_3027,N_858);
nor U3860 (N_3860,N_2024,N_883);
nand U3861 (N_3861,N_2632,N_1651);
nand U3862 (N_3862,N_1481,N_2198);
or U3863 (N_3863,N_537,N_2571);
xnor U3864 (N_3864,N_1797,N_2745);
nor U3865 (N_3865,N_639,N_1304);
nand U3866 (N_3866,N_1874,N_1635);
nor U3867 (N_3867,N_1443,N_1541);
or U3868 (N_3868,N_3058,N_2493);
nor U3869 (N_3869,N_2748,N_458);
and U3870 (N_3870,N_1071,N_1994);
xnor U3871 (N_3871,N_3094,N_2942);
nor U3872 (N_3872,N_1142,N_2251);
nor U3873 (N_3873,N_893,N_985);
nor U3874 (N_3874,N_669,N_1089);
nor U3875 (N_3875,N_656,N_42);
nand U3876 (N_3876,N_1650,N_443);
nand U3877 (N_3877,N_611,N_2287);
or U3878 (N_3878,N_1914,N_1155);
and U3879 (N_3879,N_1748,N_1646);
xnor U3880 (N_3880,N_2964,N_1632);
nor U3881 (N_3881,N_17,N_1191);
and U3882 (N_3882,N_2304,N_1741);
xor U3883 (N_3883,N_2112,N_103);
xor U3884 (N_3884,N_2921,N_1827);
and U3885 (N_3885,N_2385,N_2020);
or U3886 (N_3886,N_2494,N_2065);
and U3887 (N_3887,N_2406,N_475);
nand U3888 (N_3888,N_501,N_2191);
and U3889 (N_3889,N_1263,N_3063);
xor U3890 (N_3890,N_2205,N_1299);
nand U3891 (N_3891,N_2300,N_2988);
nor U3892 (N_3892,N_1814,N_2259);
and U3893 (N_3893,N_576,N_1079);
nand U3894 (N_3894,N_944,N_2898);
or U3895 (N_3895,N_931,N_2150);
nor U3896 (N_3896,N_1352,N_1212);
nand U3897 (N_3897,N_13,N_557);
xor U3898 (N_3898,N_1806,N_2118);
or U3899 (N_3899,N_2039,N_2399);
xnor U3900 (N_3900,N_389,N_1270);
xnor U3901 (N_3901,N_795,N_2089);
nor U3902 (N_3902,N_1120,N_1069);
nor U3903 (N_3903,N_471,N_290);
nor U3904 (N_3904,N_178,N_1988);
nand U3905 (N_3905,N_1954,N_2660);
nand U3906 (N_3906,N_2197,N_2544);
nand U3907 (N_3907,N_750,N_1385);
or U3908 (N_3908,N_615,N_1609);
nand U3909 (N_3909,N_2394,N_2662);
or U3910 (N_3910,N_2400,N_830);
and U3911 (N_3911,N_520,N_377);
and U3912 (N_3912,N_1995,N_1753);
nand U3913 (N_3913,N_2613,N_2352);
xor U3914 (N_3914,N_2061,N_1196);
or U3915 (N_3915,N_282,N_1162);
nor U3916 (N_3916,N_363,N_638);
and U3917 (N_3917,N_2135,N_1293);
nand U3918 (N_3918,N_1638,N_1792);
and U3919 (N_3919,N_2211,N_1019);
xor U3920 (N_3920,N_1900,N_980);
nand U3921 (N_3921,N_380,N_2958);
and U3922 (N_3922,N_469,N_28);
or U3923 (N_3923,N_1399,N_1689);
and U3924 (N_3924,N_2818,N_1062);
nand U3925 (N_3925,N_2496,N_2828);
or U3926 (N_3926,N_937,N_2285);
nand U3927 (N_3927,N_447,N_1833);
or U3928 (N_3928,N_1552,N_1388);
or U3929 (N_3929,N_2185,N_3099);
nand U3930 (N_3930,N_2210,N_1567);
nand U3931 (N_3931,N_1941,N_2760);
or U3932 (N_3932,N_354,N_621);
nand U3933 (N_3933,N_2602,N_1534);
and U3934 (N_3934,N_1560,N_670);
nand U3935 (N_3935,N_820,N_2471);
and U3936 (N_3936,N_601,N_1310);
or U3937 (N_3937,N_467,N_2004);
or U3938 (N_3938,N_2902,N_1489);
nand U3939 (N_3939,N_1593,N_1691);
and U3940 (N_3940,N_2560,N_1309);
or U3941 (N_3941,N_105,N_2430);
and U3942 (N_3942,N_2360,N_2944);
or U3943 (N_3943,N_3031,N_2815);
or U3944 (N_3944,N_2578,N_464);
nor U3945 (N_3945,N_1964,N_586);
or U3946 (N_3946,N_1437,N_568);
nor U3947 (N_3947,N_492,N_262);
or U3948 (N_3948,N_114,N_2363);
or U3949 (N_3949,N_777,N_121);
nand U3950 (N_3950,N_2116,N_703);
and U3951 (N_3951,N_376,N_2250);
xor U3952 (N_3952,N_1857,N_694);
xor U3953 (N_3953,N_2248,N_727);
nor U3954 (N_3954,N_3103,N_873);
or U3955 (N_3955,N_2802,N_698);
nand U3956 (N_3956,N_1540,N_1376);
nor U3957 (N_3957,N_1795,N_1786);
and U3958 (N_3958,N_2643,N_864);
and U3959 (N_3959,N_2777,N_1652);
nor U3960 (N_3960,N_943,N_1764);
nor U3961 (N_3961,N_1899,N_1886);
and U3962 (N_3962,N_2076,N_929);
xor U3963 (N_3963,N_228,N_1487);
nor U3964 (N_3964,N_2744,N_2837);
and U3965 (N_3965,N_77,N_2591);
nor U3966 (N_3966,N_44,N_2025);
or U3967 (N_3967,N_2372,N_342);
nand U3968 (N_3968,N_971,N_1893);
and U3969 (N_3969,N_1519,N_1736);
nor U3970 (N_3970,N_1667,N_942);
xnor U3971 (N_3971,N_1056,N_910);
and U3972 (N_3972,N_1872,N_309);
and U3973 (N_3973,N_325,N_3097);
and U3974 (N_3974,N_2892,N_2624);
xor U3975 (N_3975,N_108,N_1525);
nor U3976 (N_3976,N_719,N_147);
nor U3977 (N_3977,N_655,N_1451);
xnor U3978 (N_3978,N_1165,N_898);
or U3979 (N_3979,N_2227,N_2010);
nor U3980 (N_3980,N_484,N_1180);
nand U3981 (N_3981,N_2319,N_3069);
or U3982 (N_3982,N_1170,N_1117);
nor U3983 (N_3983,N_2049,N_2852);
nand U3984 (N_3984,N_0,N_3055);
nor U3985 (N_3985,N_1216,N_2199);
xnor U3986 (N_3986,N_1750,N_2120);
nor U3987 (N_3987,N_395,N_431);
nand U3988 (N_3988,N_1041,N_1064);
or U3989 (N_3989,N_1539,N_1339);
nand U3990 (N_3990,N_274,N_2446);
and U3991 (N_3991,N_581,N_444);
xor U3992 (N_3992,N_840,N_155);
or U3993 (N_3993,N_316,N_2987);
nand U3994 (N_3994,N_1817,N_100);
or U3995 (N_3995,N_1572,N_1048);
xor U3996 (N_3996,N_602,N_2561);
and U3997 (N_3997,N_1590,N_283);
nor U3998 (N_3998,N_333,N_767);
and U3999 (N_3999,N_1636,N_451);
and U4000 (N_4000,N_2566,N_1049);
xnor U4001 (N_4001,N_1185,N_1516);
nor U4002 (N_4002,N_3100,N_1424);
or U4003 (N_4003,N_1631,N_1713);
nand U4004 (N_4004,N_2832,N_1022);
nor U4005 (N_4005,N_2421,N_745);
nor U4006 (N_4006,N_1729,N_614);
nor U4007 (N_4007,N_1438,N_175);
nor U4008 (N_4008,N_1118,N_2396);
or U4009 (N_4009,N_1250,N_113);
or U4010 (N_4010,N_2477,N_1074);
nor U4011 (N_4011,N_2976,N_323);
nor U4012 (N_4012,N_1252,N_259);
nand U4013 (N_4013,N_768,N_1463);
nor U4014 (N_4014,N_544,N_2074);
and U4015 (N_4015,N_1502,N_2911);
or U4016 (N_4016,N_1625,N_2963);
nand U4017 (N_4017,N_23,N_2831);
or U4018 (N_4018,N_728,N_1236);
nor U4019 (N_4019,N_2353,N_2894);
and U4020 (N_4020,N_2184,N_925);
nand U4021 (N_4021,N_2109,N_2614);
and U4022 (N_4022,N_2960,N_2220);
nor U4023 (N_4023,N_1276,N_516);
and U4024 (N_4024,N_1204,N_580);
and U4025 (N_4025,N_1195,N_3113);
xor U4026 (N_4026,N_2652,N_1683);
and U4027 (N_4027,N_1990,N_572);
and U4028 (N_4028,N_2648,N_2378);
nand U4029 (N_4029,N_2212,N_1213);
nand U4030 (N_4030,N_968,N_1727);
nand U4031 (N_4031,N_1978,N_574);
xor U4032 (N_4032,N_2111,N_950);
or U4033 (N_4033,N_1654,N_2225);
or U4034 (N_4034,N_2362,N_736);
xor U4035 (N_4035,N_1919,N_1716);
or U4036 (N_4036,N_1842,N_1850);
nand U4037 (N_4037,N_644,N_808);
nor U4038 (N_4038,N_1533,N_2072);
nand U4039 (N_4039,N_214,N_34);
nor U4040 (N_4040,N_1660,N_2779);
or U4041 (N_4041,N_340,N_119);
and U4042 (N_4042,N_1324,N_1809);
nor U4043 (N_4043,N_699,N_41);
nand U4044 (N_4044,N_2401,N_1051);
nor U4045 (N_4045,N_623,N_1611);
xnor U4046 (N_4046,N_2689,N_1123);
xnor U4047 (N_4047,N_831,N_2064);
or U4048 (N_4048,N_111,N_48);
nand U4049 (N_4049,N_2261,N_2785);
and U4050 (N_4050,N_1875,N_1400);
nor U4051 (N_4051,N_1107,N_1111);
and U4052 (N_4052,N_1653,N_2842);
nand U4053 (N_4053,N_1911,N_468);
nor U4054 (N_4054,N_104,N_1904);
or U4055 (N_4055,N_1417,N_2721);
and U4056 (N_4056,N_2006,N_2277);
and U4057 (N_4057,N_3115,N_1431);
nand U4058 (N_4058,N_3010,N_1807);
and U4059 (N_4059,N_1678,N_341);
or U4060 (N_4060,N_1413,N_1168);
nor U4061 (N_4061,N_2161,N_783);
nor U4062 (N_4062,N_2899,N_3068);
and U4063 (N_4063,N_3092,N_2270);
and U4064 (N_4064,N_173,N_2429);
and U4065 (N_4065,N_749,N_774);
nor U4066 (N_4066,N_426,N_2932);
and U4067 (N_4067,N_1129,N_3000);
nand U4068 (N_4068,N_966,N_2154);
and U4069 (N_4069,N_1343,N_2762);
nor U4070 (N_4070,N_1029,N_2151);
and U4071 (N_4071,N_428,N_210);
nor U4072 (N_4072,N_230,N_1044);
and U4073 (N_4073,N_254,N_2037);
and U4074 (N_4074,N_1199,N_718);
or U4075 (N_4075,N_1251,N_2357);
or U4076 (N_4076,N_2556,N_1052);
and U4077 (N_4077,N_701,N_88);
nand U4078 (N_4078,N_1686,N_1379);
nor U4079 (N_4079,N_2702,N_1744);
nand U4080 (N_4080,N_1695,N_2644);
and U4081 (N_4081,N_3075,N_2367);
and U4082 (N_4082,N_1038,N_1028);
nor U4083 (N_4083,N_2638,N_2055);
and U4084 (N_4084,N_3051,N_2392);
nor U4085 (N_4085,N_427,N_213);
nand U4086 (N_4086,N_304,N_804);
or U4087 (N_4087,N_1647,N_1693);
nand U4088 (N_4088,N_1179,N_2093);
and U4089 (N_4089,N_1394,N_3039);
or U4090 (N_4090,N_1346,N_857);
nand U4091 (N_4091,N_2848,N_1211);
or U4092 (N_4092,N_2715,N_1615);
and U4093 (N_4093,N_2217,N_185);
or U4094 (N_4094,N_801,N_193);
nor U4095 (N_4095,N_1598,N_2626);
or U4096 (N_4096,N_245,N_650);
nor U4097 (N_4097,N_975,N_2881);
and U4098 (N_4098,N_1330,N_1189);
nor U4099 (N_4099,N_1072,N_2168);
xor U4100 (N_4100,N_1025,N_1663);
and U4101 (N_4101,N_2838,N_1513);
nor U4102 (N_4102,N_2340,N_278);
nor U4103 (N_4103,N_2814,N_641);
nand U4104 (N_4104,N_1679,N_1205);
xnor U4105 (N_4105,N_989,N_73);
xor U4106 (N_4106,N_1965,N_3078);
nor U4107 (N_4107,N_1288,N_2680);
nor U4108 (N_4108,N_2985,N_1232);
or U4109 (N_4109,N_2883,N_880);
and U4110 (N_4110,N_1854,N_250);
and U4111 (N_4111,N_2844,N_2870);
or U4112 (N_4112,N_1547,N_86);
nand U4113 (N_4113,N_2961,N_83);
or U4114 (N_4114,N_2341,N_1262);
nand U4115 (N_4115,N_1014,N_2459);
or U4116 (N_4116,N_1145,N_2235);
nand U4117 (N_4117,N_1292,N_378);
xor U4118 (N_4118,N_1622,N_268);
nor U4119 (N_4119,N_685,N_1775);
xor U4120 (N_4120,N_693,N_3076);
nand U4121 (N_4121,N_531,N_2099);
nand U4122 (N_4122,N_901,N_936);
or U4123 (N_4123,N_2327,N_2260);
nand U4124 (N_4124,N_1351,N_1649);
or U4125 (N_4125,N_1510,N_1890);
nor U4126 (N_4126,N_2152,N_2467);
or U4127 (N_4127,N_2738,N_2036);
nor U4128 (N_4128,N_1751,N_2178);
and U4129 (N_4129,N_3061,N_1582);
nand U4130 (N_4130,N_456,N_2193);
nand U4131 (N_4131,N_1109,N_93);
nand U4132 (N_4132,N_2569,N_2416);
nand U4133 (N_4133,N_1447,N_2533);
nand U4134 (N_4134,N_307,N_448);
and U4135 (N_4135,N_2007,N_1039);
or U4136 (N_4136,N_3120,N_3037);
or U4137 (N_4137,N_364,N_31);
nand U4138 (N_4138,N_2384,N_2391);
and U4139 (N_4139,N_1188,N_1108);
or U4140 (N_4140,N_2233,N_388);
xor U4141 (N_4141,N_1471,N_1174);
nand U4142 (N_4142,N_2018,N_289);
or U4143 (N_4143,N_2255,N_2131);
and U4144 (N_4144,N_2369,N_2293);
or U4145 (N_4145,N_1106,N_301);
or U4146 (N_4146,N_1137,N_2209);
xnor U4147 (N_4147,N_1099,N_3086);
and U4148 (N_4148,N_1088,N_2930);
nand U4149 (N_4149,N_1555,N_906);
and U4150 (N_4150,N_2589,N_1755);
and U4151 (N_4151,N_1935,N_2955);
nand U4152 (N_4152,N_97,N_743);
nand U4153 (N_4153,N_1473,N_881);
xnor U4154 (N_4154,N_1945,N_2552);
or U4155 (N_4155,N_2567,N_2033);
or U4156 (N_4156,N_2022,N_954);
or U4157 (N_4157,N_2126,N_2529);
nor U4158 (N_4158,N_2513,N_1380);
or U4159 (N_4159,N_1265,N_1090);
nand U4160 (N_4160,N_1058,N_2925);
and U4161 (N_4161,N_2499,N_410);
or U4162 (N_4162,N_370,N_7);
nor U4163 (N_4163,N_913,N_2325);
and U4164 (N_4164,N_706,N_241);
nand U4165 (N_4165,N_2044,N_330);
nor U4166 (N_4166,N_702,N_1367);
xnor U4167 (N_4167,N_3007,N_740);
or U4168 (N_4168,N_1094,N_294);
nand U4169 (N_4169,N_1996,N_2019);
and U4170 (N_4170,N_1462,N_3104);
or U4171 (N_4171,N_2766,N_1579);
nor U4172 (N_4172,N_847,N_1981);
nor U4173 (N_4173,N_1511,N_871);
nand U4174 (N_4174,N_3041,N_1147);
xnor U4175 (N_4175,N_1306,N_1601);
or U4176 (N_4176,N_2789,N_1581);
and U4177 (N_4177,N_1418,N_2050);
or U4178 (N_4178,N_766,N_1562);
nand U4179 (N_4179,N_2310,N_1101);
nand U4180 (N_4180,N_1521,N_1241);
or U4181 (N_4181,N_1154,N_1143);
nor U4182 (N_4182,N_3089,N_430);
or U4183 (N_4183,N_627,N_3050);
nor U4184 (N_4184,N_3036,N_2330);
or U4185 (N_4185,N_558,N_1522);
nor U4186 (N_4186,N_1675,N_1497);
nand U4187 (N_4187,N_2204,N_223);
and U4188 (N_4188,N_2160,N_2676);
nor U4189 (N_4189,N_2605,N_700);
nor U4190 (N_4190,N_775,N_1098);
nor U4191 (N_4191,N_1184,N_1743);
nor U4192 (N_4192,N_2374,N_2882);
and U4193 (N_4193,N_2243,N_2003);
and U4194 (N_4194,N_2457,N_1235);
nand U4195 (N_4195,N_617,N_197);
xor U4196 (N_4196,N_1556,N_152);
nor U4197 (N_4197,N_1672,N_2047);
nor U4198 (N_4198,N_2812,N_1197);
or U4199 (N_4199,N_563,N_1760);
or U4200 (N_4200,N_1847,N_2444);
and U4201 (N_4201,N_2440,N_2433);
nand U4202 (N_4202,N_1944,N_1206);
or U4203 (N_4203,N_82,N_2368);
and U4204 (N_4204,N_2747,N_1131);
nand U4205 (N_4205,N_996,N_1669);
nand U4206 (N_4206,N_2583,N_2947);
xnor U4207 (N_4207,N_2607,N_551);
and U4208 (N_4208,N_1214,N_461);
nand U4209 (N_4209,N_737,N_1254);
or U4210 (N_4210,N_1474,N_3011);
nor U4211 (N_4211,N_710,N_1340);
and U4212 (N_4212,N_1887,N_2682);
or U4213 (N_4213,N_19,N_129);
or U4214 (N_4214,N_46,N_166);
nand U4215 (N_4215,N_242,N_2937);
nor U4216 (N_4216,N_2201,N_1428);
and U4217 (N_4217,N_1496,N_89);
xnor U4218 (N_4218,N_1365,N_754);
nor U4219 (N_4219,N_1323,N_2336);
nand U4220 (N_4220,N_2540,N_1551);
or U4221 (N_4221,N_1903,N_102);
nor U4222 (N_4222,N_1676,N_1313);
nand U4223 (N_4223,N_1557,N_2906);
xnor U4224 (N_4224,N_3034,N_789);
and U4225 (N_4225,N_505,N_1620);
nor U4226 (N_4226,N_2974,N_1656);
and U4227 (N_4227,N_533,N_1717);
nor U4228 (N_4228,N_1515,N_1977);
nand U4229 (N_4229,N_1829,N_2980);
xor U4230 (N_4230,N_2002,N_1026);
or U4231 (N_4231,N_2877,N_2140);
or U4232 (N_4232,N_3066,N_402);
and U4233 (N_4233,N_1317,N_811);
and U4234 (N_4234,N_1920,N_1483);
nand U4235 (N_4235,N_314,N_2936);
nand U4236 (N_4236,N_686,N_1834);
nand U4237 (N_4237,N_903,N_630);
xnor U4238 (N_4238,N_2324,N_2841);
or U4239 (N_4239,N_483,N_517);
and U4240 (N_4240,N_2469,N_211);
and U4241 (N_4241,N_2801,N_2519);
nand U4242 (N_4242,N_462,N_315);
xor U4243 (N_4243,N_1680,N_2296);
nor U4244 (N_4244,N_872,N_2729);
xnor U4245 (N_4245,N_2623,N_3026);
nand U4246 (N_4246,N_2754,N_618);
xnor U4247 (N_4247,N_1571,N_361);
nand U4248 (N_4248,N_2452,N_2752);
or U4249 (N_4249,N_1208,N_1905);
or U4250 (N_4250,N_726,N_1546);
or U4251 (N_4251,N_2083,N_2470);
and U4252 (N_4252,N_2665,N_1558);
or U4253 (N_4253,N_1670,N_1715);
or U4254 (N_4254,N_2395,N_1942);
nor U4255 (N_4255,N_1030,N_2655);
or U4256 (N_4256,N_1720,N_604);
xor U4257 (N_4257,N_2968,N_1623);
and U4258 (N_4258,N_1984,N_2866);
xnor U4259 (N_4259,N_2586,N_1148);
nand U4260 (N_4260,N_2756,N_161);
nor U4261 (N_4261,N_899,N_445);
nor U4262 (N_4262,N_1861,N_2800);
and U4263 (N_4263,N_218,N_368);
xor U4264 (N_4264,N_836,N_2215);
and U4265 (N_4265,N_2230,N_1361);
nor U4266 (N_4266,N_372,N_814);
or U4267 (N_4267,N_1158,N_2941);
nor U4268 (N_4268,N_2853,N_1711);
nand U4269 (N_4269,N_2629,N_979);
nor U4270 (N_4270,N_149,N_773);
and U4271 (N_4271,N_690,N_2839);
xor U4272 (N_4272,N_480,N_446);
nand U4273 (N_4273,N_2821,N_1182);
or U4274 (N_4274,N_676,N_2582);
or U4275 (N_4275,N_2153,N_819);
nand U4276 (N_4276,N_2531,N_2971);
and U4277 (N_4277,N_683,N_1495);
nand U4278 (N_4278,N_2989,N_2609);
or U4279 (N_4279,N_1862,N_757);
nor U4280 (N_4280,N_203,N_2398);
nor U4281 (N_4281,N_2386,N_225);
nand U4282 (N_4282,N_1851,N_2547);
nor U4283 (N_4283,N_1311,N_1076);
nor U4284 (N_4284,N_1390,N_2455);
or U4285 (N_4285,N_1122,N_643);
nand U4286 (N_4286,N_653,N_1554);
nand U4287 (N_4287,N_2900,N_1830);
or U4288 (N_4288,N_846,N_2732);
or U4289 (N_4289,N_439,N_266);
nor U4290 (N_4290,N_1759,N_2515);
and U4291 (N_4291,N_2425,N_486);
or U4292 (N_4292,N_1445,N_2761);
or U4293 (N_4293,N_922,N_45);
xnor U4294 (N_4294,N_3091,N_1780);
nand U4295 (N_4295,N_959,N_116);
nand U4296 (N_4296,N_634,N_2929);
and U4297 (N_4297,N_1177,N_331);
xor U4298 (N_4298,N_2226,N_974);
or U4299 (N_4299,N_1738,N_375);
and U4300 (N_4300,N_1403,N_771);
nor U4301 (N_4301,N_1161,N_848);
nor U4302 (N_4302,N_332,N_2053);
xnor U4303 (N_4303,N_1752,N_571);
xnor U4304 (N_4304,N_2449,N_2946);
nand U4305 (N_4305,N_2504,N_401);
and U4306 (N_4306,N_1389,N_2222);
or U4307 (N_4307,N_2833,N_1226);
and U4308 (N_4308,N_1586,N_2474);
and U4309 (N_4309,N_1081,N_2339);
xor U4310 (N_4310,N_2453,N_2079);
nor U4311 (N_4311,N_61,N_2090);
and U4312 (N_4312,N_1600,N_2717);
xnor U4313 (N_4313,N_2175,N_837);
nor U4314 (N_4314,N_2576,N_705);
and U4315 (N_4315,N_1316,N_2262);
and U4316 (N_4316,N_1524,N_592);
xor U4317 (N_4317,N_195,N_1322);
and U4318 (N_4318,N_2646,N_2997);
nor U4319 (N_4319,N_2487,N_1008);
nand U4320 (N_4320,N_2847,N_575);
or U4321 (N_4321,N_277,N_1740);
and U4322 (N_4322,N_1287,N_126);
or U4323 (N_4323,N_890,N_63);
and U4324 (N_4324,N_723,N_29);
nand U4325 (N_4325,N_273,N_1815);
and U4326 (N_4326,N_1369,N_549);
and U4327 (N_4327,N_235,N_1910);
and U4328 (N_4328,N_2337,N_689);
and U4329 (N_4329,N_2016,N_2817);
or U4330 (N_4330,N_1953,N_2735);
nor U4331 (N_4331,N_2115,N_2316);
nand U4332 (N_4332,N_2106,N_734);
or U4333 (N_4333,N_2317,N_2706);
nand U4334 (N_4334,N_1000,N_16);
or U4335 (N_4335,N_606,N_1948);
or U4336 (N_4336,N_567,N_1866);
and U4337 (N_4337,N_249,N_2992);
nor U4338 (N_4338,N_326,N_875);
and U4339 (N_4339,N_1884,N_2366);
and U4340 (N_4340,N_1773,N_472);
nor U4341 (N_4341,N_532,N_5);
nor U4342 (N_4342,N_1831,N_772);
and U4343 (N_4343,N_1130,N_1297);
and U4344 (N_4344,N_327,N_1057);
and U4345 (N_4345,N_139,N_2516);
nor U4346 (N_4346,N_2720,N_2381);
nor U4347 (N_4347,N_1730,N_2637);
nand U4348 (N_4348,N_3053,N_1662);
nor U4349 (N_4349,N_1707,N_845);
or U4350 (N_4350,N_1803,N_885);
or U4351 (N_4351,N_137,N_25);
nor U4352 (N_4352,N_2096,N_1867);
and U4353 (N_4353,N_1377,N_2142);
nand U4354 (N_4354,N_2297,N_2375);
xor U4355 (N_4355,N_500,N_2956);
or U4356 (N_4356,N_2712,N_2346);
nand U4357 (N_4357,N_1645,N_1285);
or U4358 (N_4358,N_1405,N_199);
and U4359 (N_4359,N_2177,N_2635);
nor U4360 (N_4360,N_1500,N_1066);
nor U4361 (N_4361,N_1001,N_1461);
nor U4362 (N_4362,N_1425,N_2505);
nand U4363 (N_4363,N_2155,N_891);
xor U4364 (N_4364,N_2622,N_2130);
and U4365 (N_4365,N_2432,N_2473);
and U4366 (N_4366,N_952,N_2661);
nor U4367 (N_4367,N_2027,N_2163);
or U4368 (N_4368,N_1783,N_2286);
xnor U4369 (N_4369,N_607,N_2409);
nand U4370 (N_4370,N_1916,N_1115);
and U4371 (N_4371,N_2608,N_2587);
nand U4372 (N_4372,N_287,N_1326);
nand U4373 (N_4373,N_547,N_2845);
and U4374 (N_4374,N_951,N_866);
and U4375 (N_4375,N_2856,N_2940);
nand U4376 (N_4376,N_2026,N_823);
nor U4377 (N_4377,N_2799,N_865);
or U4378 (N_4378,N_320,N_2442);
and U4379 (N_4379,N_1103,N_958);
nor U4380 (N_4380,N_2232,N_1721);
and U4381 (N_4381,N_947,N_414);
nor U4382 (N_4382,N_3095,N_812);
nand U4383 (N_4383,N_1835,N_2437);
and U4384 (N_4384,N_1059,N_127);
or U4385 (N_4385,N_704,N_1684);
nor U4386 (N_4386,N_915,N_2171);
and U4387 (N_4387,N_205,N_2935);
xnor U4388 (N_4388,N_1845,N_59);
nand U4389 (N_4389,N_2975,N_2771);
nand U4390 (N_4390,N_22,N_1077);
nand U4391 (N_4391,N_1366,N_1295);
nand U4392 (N_4392,N_171,N_779);
nand U4393 (N_4393,N_1856,N_58);
or U4394 (N_4394,N_3109,N_1167);
or U4395 (N_4395,N_613,N_1087);
or U4396 (N_4396,N_2683,N_2274);
nor U4397 (N_4397,N_1614,N_1280);
or U4398 (N_4398,N_2667,N_2278);
and U4399 (N_4399,N_521,N_2322);
nor U4400 (N_4400,N_632,N_1221);
nor U4401 (N_4401,N_603,N_784);
or U4402 (N_4402,N_731,N_1406);
nor U4403 (N_4403,N_1075,N_1789);
nand U4404 (N_4404,N_3030,N_1227);
nand U4405 (N_4405,N_3047,N_1776);
nand U4406 (N_4406,N_1701,N_2508);
nor U4407 (N_4407,N_1739,N_1183);
and U4408 (N_4408,N_1602,N_1360);
nor U4409 (N_4409,N_1175,N_2481);
and U4410 (N_4410,N_90,N_172);
nor U4411 (N_4411,N_1597,N_940);
nor U4412 (N_4412,N_112,N_577);
nor U4413 (N_4413,N_56,N_2008);
and U4414 (N_4414,N_2417,N_687);
nand U4415 (N_4415,N_1386,N_886);
or U4416 (N_4416,N_1912,N_3107);
and U4417 (N_4417,N_2688,N_415);
nor U4418 (N_4418,N_1260,N_2530);
nand U4419 (N_4419,N_432,N_2272);
or U4420 (N_4420,N_1398,N_1003);
nor U4421 (N_4421,N_1698,N_2952);
and U4422 (N_4422,N_1404,N_2364);
or U4423 (N_4423,N_2125,N_2094);
nor U4424 (N_4424,N_2954,N_1200);
nor U4425 (N_4425,N_1010,N_130);
nand U4426 (N_4426,N_27,N_879);
nor U4427 (N_4427,N_1013,N_143);
nand U4428 (N_4428,N_1448,N_1409);
and U4429 (N_4429,N_1264,N_1879);
or U4430 (N_4430,N_3045,N_2509);
nor U4431 (N_4431,N_2910,N_8);
or U4432 (N_4432,N_582,N_2144);
nand U4433 (N_4433,N_2535,N_2102);
nand U4434 (N_4434,N_692,N_141);
and U4435 (N_4435,N_374,N_66);
nand U4436 (N_4436,N_1268,N_3088);
or U4437 (N_4437,N_1228,N_2658);
and U4438 (N_4438,N_1231,N_1105);
xor U4439 (N_4439,N_110,N_2258);
and U4440 (N_4440,N_474,N_2949);
or U4441 (N_4441,N_1016,N_786);
nand U4442 (N_4442,N_862,N_1353);
nand U4443 (N_4443,N_2434,N_2885);
xnor U4444 (N_4444,N_1641,N_545);
xor U4445 (N_4445,N_546,N_1864);
nand U4446 (N_4446,N_715,N_3085);
and U4447 (N_4447,N_2068,N_2443);
or U4448 (N_4448,N_1411,N_2934);
nor U4449 (N_4449,N_2663,N_874);
nand U4450 (N_4450,N_2195,N_631);
nor U4451 (N_4451,N_770,N_2257);
or U4452 (N_4452,N_1401,N_2048);
nor U4453 (N_4453,N_92,N_2097);
nor U4454 (N_4454,N_535,N_540);
or U4455 (N_4455,N_3098,N_2897);
and U4456 (N_4456,N_1734,N_2000);
and U4457 (N_4457,N_2514,N_2427);
and U4458 (N_4458,N_1985,N_2294);
and U4459 (N_4459,N_824,N_219);
nor U4460 (N_4460,N_556,N_3110);
or U4461 (N_4461,N_1220,N_411);
or U4462 (N_4462,N_2692,N_1178);
and U4463 (N_4463,N_382,N_2805);
xor U4464 (N_4464,N_2865,N_1943);
nor U4465 (N_4465,N_2757,N_2062);
nor U4466 (N_4466,N_1888,N_2236);
nand U4467 (N_4467,N_1574,N_2719);
nand U4468 (N_4468,N_2628,N_2592);
nor U4469 (N_4469,N_347,N_280);
and U4470 (N_4470,N_788,N_716);
and U4471 (N_4471,N_1837,N_2435);
nor U4472 (N_4472,N_1452,N_992);
nand U4473 (N_4473,N_2596,N_2642);
and U4474 (N_4474,N_198,N_593);
or U4475 (N_4475,N_2651,N_792);
nor U4476 (N_4476,N_298,N_1992);
nor U4477 (N_4477,N_1828,N_117);
nor U4478 (N_4478,N_1282,N_2134);
nand U4479 (N_4479,N_1770,N_24);
or U4480 (N_4480,N_2196,N_2520);
and U4481 (N_4481,N_2214,N_2758);
and U4482 (N_4482,N_2926,N_1136);
nand U4483 (N_4483,N_2305,N_1186);
and U4484 (N_4484,N_776,N_2066);
or U4485 (N_4485,N_1442,N_2299);
nand U4486 (N_4486,N_1464,N_2190);
and U4487 (N_4487,N_2051,N_778);
nand U4488 (N_4488,N_2445,N_2913);
nand U4489 (N_4489,N_907,N_1702);
nand U4490 (N_4490,N_68,N_265);
nor U4491 (N_4491,N_2273,N_3023);
or U4492 (N_4492,N_2035,N_2045);
or U4493 (N_4493,N_1993,N_2070);
and U4494 (N_4494,N_437,N_3081);
nor U4495 (N_4495,N_553,N_2488);
and U4496 (N_4496,N_798,N_2393);
and U4497 (N_4497,N_2388,N_1173);
xnor U4498 (N_4498,N_1127,N_2143);
and U4499 (N_4499,N_2951,N_381);
nand U4500 (N_4500,N_2668,N_2321);
and U4501 (N_4501,N_2650,N_1564);
and U4502 (N_4502,N_1095,N_3067);
and U4503 (N_4503,N_1808,N_2200);
nand U4504 (N_4504,N_1332,N_1314);
nand U4505 (N_4505,N_1745,N_1724);
and U4506 (N_4506,N_552,N_949);
or U4507 (N_4507,N_450,N_1897);
nor U4508 (N_4508,N_1190,N_2411);
nor U4509 (N_4509,N_1906,N_594);
nand U4510 (N_4510,N_360,N_522);
nor U4511 (N_4511,N_1694,N_1499);
nand U4512 (N_4512,N_233,N_1021);
and U4513 (N_4513,N_2087,N_386);
nor U4514 (N_4514,N_1277,N_1371);
nor U4515 (N_4515,N_2382,N_2699);
nor U4516 (N_4516,N_2512,N_352);
or U4517 (N_4517,N_1466,N_813);
nand U4518 (N_4518,N_1356,N_473);
nand U4519 (N_4519,N_528,N_1559);
and U4520 (N_4520,N_2927,N_2808);
nor U4521 (N_4521,N_106,N_995);
nand U4522 (N_4522,N_2618,N_40);
or U4523 (N_4523,N_3077,N_578);
nand U4524 (N_4524,N_2753,N_292);
xnor U4525 (N_4525,N_2835,N_564);
or U4526 (N_4526,N_3017,N_1685);
and U4527 (N_4527,N_2180,N_1);
or U4528 (N_4528,N_1584,N_1384);
and U4529 (N_4529,N_2673,N_1634);
nor U4530 (N_4530,N_504,N_1971);
nand U4531 (N_4531,N_2829,N_60);
nor U4532 (N_4532,N_1290,N_1570);
xor U4533 (N_4533,N_833,N_682);
xor U4534 (N_4534,N_526,N_2765);
xor U4535 (N_4535,N_440,N_2344);
and U4536 (N_4536,N_306,N_834);
xnor U4537 (N_4537,N_821,N_2601);
or U4538 (N_4538,N_2241,N_1726);
nand U4539 (N_4539,N_407,N_2664);
and U4540 (N_4540,N_3106,N_146);
nor U4541 (N_4541,N_2998,N_2267);
nor U4542 (N_4542,N_2674,N_2731);
nor U4543 (N_4543,N_713,N_1952);
and U4544 (N_4544,N_714,N_681);
and U4545 (N_4545,N_1113,N_2823);
nand U4546 (N_4546,N_762,N_2827);
or U4547 (N_4547,N_867,N_629);
or U4548 (N_4548,N_609,N_1430);
xor U4549 (N_4549,N_1187,N_1396);
nand U4550 (N_4550,N_1538,N_3062);
nand U4551 (N_4551,N_1269,N_1372);
nor U4552 (N_4552,N_2167,N_2889);
xnor U4553 (N_4553,N_2871,N_1841);
nor U4554 (N_4554,N_1478,N_1895);
or U4555 (N_4555,N_144,N_928);
or U4556 (N_4556,N_302,N_94);
nor U4557 (N_4557,N_2755,N_313);
nor U4558 (N_4558,N_1073,N_841);
nand U4559 (N_4559,N_2244,N_2546);
nand U4560 (N_4560,N_260,N_2081);
or U4561 (N_4561,N_2807,N_206);
and U4562 (N_4562,N_231,N_1664);
nor U4563 (N_4563,N_2855,N_3009);
or U4564 (N_4564,N_317,N_1677);
and U4565 (N_4565,N_2631,N_2376);
xor U4566 (N_4566,N_2819,N_2572);
xor U4567 (N_4567,N_1133,N_2359);
or U4568 (N_4568,N_796,N_138);
nor U4569 (N_4569,N_2289,N_1820);
nand U4570 (N_4570,N_3001,N_449);
or U4571 (N_4571,N_932,N_2080);
xor U4572 (N_4572,N_654,N_3028);
xor U4573 (N_4573,N_1153,N_1982);
nand U4574 (N_4574,N_1256,N_2548);
and U4575 (N_4575,N_2770,N_1434);
xor U4576 (N_4576,N_2598,N_1688);
or U4577 (N_4577,N_2436,N_590);
nand U4578 (N_4578,N_2690,N_466);
and U4579 (N_4579,N_2162,N_406);
nand U4580 (N_4580,N_2813,N_2969);
xnor U4581 (N_4581,N_184,N_717);
and U4582 (N_4582,N_1171,N_2052);
nand U4583 (N_4583,N_3003,N_934);
nor U4584 (N_4584,N_2078,N_39);
and U4585 (N_4585,N_1033,N_1080);
nor U4586 (N_4586,N_2371,N_209);
xnor U4587 (N_4587,N_463,N_216);
or U4588 (N_4588,N_853,N_1215);
and U4589 (N_4589,N_192,N_2806);
nor U4590 (N_4590,N_1468,N_2498);
nand U4591 (N_4591,N_2269,N_272);
nor U4592 (N_4592,N_2649,N_1757);
and U4593 (N_4593,N_1700,N_709);
xnor U4594 (N_4594,N_477,N_2938);
nand U4595 (N_4595,N_2128,N_1908);
or U4596 (N_4596,N_1006,N_168);
and U4597 (N_4597,N_1909,N_1549);
or U4598 (N_4598,N_1383,N_1255);
or U4599 (N_4599,N_276,N_1218);
nor U4600 (N_4600,N_2707,N_1839);
and U4601 (N_4601,N_2172,N_1368);
nor U4602 (N_4602,N_722,N_1804);
or U4603 (N_4603,N_1472,N_1585);
nor U4604 (N_4604,N_441,N_1618);
nor U4605 (N_4605,N_3006,N_806);
nor U4606 (N_4606,N_1923,N_1334);
nand U4607 (N_4607,N_1454,N_523);
and U4608 (N_4608,N_1305,N_2069);
nor U4609 (N_4609,N_2872,N_2914);
nand U4610 (N_4610,N_2005,N_183);
or U4611 (N_4611,N_888,N_2931);
nand U4612 (N_4612,N_2491,N_2237);
or U4613 (N_4613,N_170,N_1800);
nand U4614 (N_4614,N_863,N_2192);
and U4615 (N_4615,N_799,N_2918);
nand U4616 (N_4616,N_1718,N_2458);
nand U4617 (N_4617,N_1336,N_2110);
nor U4618 (N_4618,N_3123,N_2521);
nor U4619 (N_4619,N_3038,N_1566);
nor U4620 (N_4620,N_2103,N_668);
xnor U4621 (N_4621,N_3049,N_752);
or U4622 (N_4622,N_1913,N_2851);
nand U4623 (N_4623,N_1160,N_373);
nor U4624 (N_4624,N_70,N_150);
xnor U4625 (N_4625,N_1024,N_145);
nor U4626 (N_4626,N_1997,N_2742);
nand U4627 (N_4627,N_2824,N_261);
nand U4628 (N_4628,N_2724,N_1423);
and U4629 (N_4629,N_2916,N_1238);
nand U4630 (N_4630,N_2678,N_3052);
nor U4631 (N_4631,N_1921,N_1110);
and U4632 (N_4632,N_2389,N_1735);
and U4633 (N_4633,N_998,N_2728);
nand U4634 (N_4634,N_724,N_3073);
and U4635 (N_4635,N_1537,N_2288);
and U4636 (N_4636,N_2840,N_454);
xnor U4637 (N_4637,N_3060,N_3084);
and U4638 (N_4638,N_133,N_973);
or U4639 (N_4639,N_1626,N_818);
or U4640 (N_4640,N_2995,N_918);
and U4641 (N_4641,N_279,N_1247);
or U4642 (N_4642,N_889,N_2034);
or U4643 (N_4643,N_984,N_167);
xor U4644 (N_4644,N_1550,N_605);
or U4645 (N_4645,N_2186,N_730);
or U4646 (N_4646,N_1342,N_2129);
or U4647 (N_4647,N_1963,N_2335);
nand U4648 (N_4648,N_478,N_425);
or U4649 (N_4649,N_2778,N_201);
nor U4650 (N_4650,N_3082,N_2749);
and U4651 (N_4651,N_502,N_459);
nand U4652 (N_4652,N_2915,N_1961);
or U4653 (N_4653,N_1930,N_418);
nor U4654 (N_4654,N_2308,N_2179);
nand U4655 (N_4655,N_2606,N_2950);
or U4656 (N_4656,N_248,N_2691);
and U4657 (N_4657,N_2803,N_2784);
or U4658 (N_4658,N_1060,N_711);
nand U4659 (N_4659,N_665,N_2917);
and U4660 (N_4660,N_1612,N_2620);
nand U4661 (N_4661,N_1223,N_739);
or U4662 (N_4662,N_2811,N_234);
nor U4663 (N_4663,N_1104,N_2361);
nand U4664 (N_4664,N_1868,N_2114);
nand U4665 (N_4665,N_1015,N_649);
nor U4666 (N_4666,N_529,N_2581);
and U4667 (N_4667,N_2986,N_176);
nor U4668 (N_4668,N_1020,N_2743);
nand U4669 (N_4669,N_1563,N_222);
and U4670 (N_4670,N_2245,N_2266);
or U4671 (N_4671,N_2408,N_1246);
or U4672 (N_4672,N_561,N_2610);
nor U4673 (N_4673,N_2279,N_1592);
nand U4674 (N_4674,N_2345,N_202);
nor U4675 (N_4675,N_2105,N_1266);
nand U4676 (N_4676,N_926,N_3002);
nand U4677 (N_4677,N_1940,N_2030);
or U4678 (N_4678,N_982,N_2315);
nor U4679 (N_4679,N_2149,N_2354);
nor U4680 (N_4680,N_2326,N_859);
nand U4681 (N_4681,N_626,N_1457);
or U4682 (N_4682,N_538,N_2283);
or U4683 (N_4683,N_65,N_2383);
nand U4684 (N_4684,N_732,N_1787);
nor U4685 (N_4685,N_1240,N_2298);
nand U4686 (N_4686,N_2303,N_1791);
or U4687 (N_4687,N_2953,N_906);
nand U4688 (N_4688,N_3022,N_3092);
nand U4689 (N_4689,N_1306,N_1980);
xor U4690 (N_4690,N_808,N_1185);
nor U4691 (N_4691,N_3068,N_756);
nor U4692 (N_4692,N_2320,N_645);
xor U4693 (N_4693,N_1265,N_198);
xnor U4694 (N_4694,N_2000,N_1027);
and U4695 (N_4695,N_2995,N_2727);
nand U4696 (N_4696,N_602,N_3022);
nor U4697 (N_4697,N_1025,N_1258);
nor U4698 (N_4698,N_2657,N_1631);
or U4699 (N_4699,N_1762,N_1121);
or U4700 (N_4700,N_403,N_1610);
and U4701 (N_4701,N_2788,N_1293);
and U4702 (N_4702,N_1321,N_1032);
xor U4703 (N_4703,N_643,N_2095);
or U4704 (N_4704,N_599,N_834);
nand U4705 (N_4705,N_465,N_226);
or U4706 (N_4706,N_2902,N_974);
nand U4707 (N_4707,N_2354,N_2361);
and U4708 (N_4708,N_2906,N_2323);
nand U4709 (N_4709,N_1084,N_868);
xor U4710 (N_4710,N_516,N_2646);
nor U4711 (N_4711,N_1301,N_211);
or U4712 (N_4712,N_97,N_33);
nor U4713 (N_4713,N_1723,N_357);
nor U4714 (N_4714,N_246,N_2935);
nand U4715 (N_4715,N_2944,N_311);
nand U4716 (N_4716,N_1713,N_2910);
nand U4717 (N_4717,N_202,N_2523);
xor U4718 (N_4718,N_787,N_2586);
nand U4719 (N_4719,N_1241,N_2887);
nand U4720 (N_4720,N_2895,N_2595);
nor U4721 (N_4721,N_2871,N_1540);
nand U4722 (N_4722,N_395,N_1025);
and U4723 (N_4723,N_2475,N_1809);
nand U4724 (N_4724,N_1764,N_481);
or U4725 (N_4725,N_2838,N_563);
or U4726 (N_4726,N_100,N_1820);
nor U4727 (N_4727,N_142,N_1604);
and U4728 (N_4728,N_1358,N_807);
nand U4729 (N_4729,N_1063,N_2692);
or U4730 (N_4730,N_2190,N_690);
nor U4731 (N_4731,N_659,N_1667);
nand U4732 (N_4732,N_1614,N_1372);
nand U4733 (N_4733,N_1730,N_2155);
nand U4734 (N_4734,N_1497,N_2980);
nand U4735 (N_4735,N_655,N_1322);
and U4736 (N_4736,N_1250,N_30);
and U4737 (N_4737,N_1770,N_2978);
or U4738 (N_4738,N_2317,N_1737);
nor U4739 (N_4739,N_1048,N_3050);
or U4740 (N_4740,N_1920,N_839);
and U4741 (N_4741,N_3105,N_352);
and U4742 (N_4742,N_234,N_458);
and U4743 (N_4743,N_2147,N_863);
nor U4744 (N_4744,N_2198,N_299);
or U4745 (N_4745,N_1044,N_2905);
xor U4746 (N_4746,N_137,N_2960);
xor U4747 (N_4747,N_2245,N_1299);
and U4748 (N_4748,N_52,N_2914);
nand U4749 (N_4749,N_1535,N_2812);
or U4750 (N_4750,N_1594,N_1152);
or U4751 (N_4751,N_3030,N_1216);
nor U4752 (N_4752,N_2005,N_320);
nor U4753 (N_4753,N_2120,N_1888);
nand U4754 (N_4754,N_2768,N_399);
nand U4755 (N_4755,N_360,N_766);
nor U4756 (N_4756,N_113,N_2023);
nor U4757 (N_4757,N_829,N_945);
nand U4758 (N_4758,N_2887,N_398);
nor U4759 (N_4759,N_2169,N_172);
nor U4760 (N_4760,N_1263,N_1753);
nor U4761 (N_4761,N_590,N_1475);
xnor U4762 (N_4762,N_2413,N_1847);
xor U4763 (N_4763,N_3032,N_222);
and U4764 (N_4764,N_428,N_499);
and U4765 (N_4765,N_22,N_2613);
or U4766 (N_4766,N_2696,N_2675);
nor U4767 (N_4767,N_1166,N_2842);
nand U4768 (N_4768,N_548,N_1763);
xor U4769 (N_4769,N_2147,N_215);
xnor U4770 (N_4770,N_2160,N_2669);
and U4771 (N_4771,N_1243,N_2799);
nand U4772 (N_4772,N_2416,N_1752);
xnor U4773 (N_4773,N_363,N_533);
and U4774 (N_4774,N_151,N_2699);
nor U4775 (N_4775,N_1392,N_1400);
nor U4776 (N_4776,N_967,N_1117);
and U4777 (N_4777,N_589,N_258);
nor U4778 (N_4778,N_2467,N_1398);
nand U4779 (N_4779,N_2030,N_1413);
nor U4780 (N_4780,N_1352,N_498);
xnor U4781 (N_4781,N_902,N_2864);
or U4782 (N_4782,N_2932,N_1043);
xnor U4783 (N_4783,N_3049,N_370);
nor U4784 (N_4784,N_2724,N_641);
or U4785 (N_4785,N_1739,N_288);
nand U4786 (N_4786,N_2420,N_2271);
or U4787 (N_4787,N_2879,N_2759);
nand U4788 (N_4788,N_707,N_99);
nand U4789 (N_4789,N_1487,N_2501);
and U4790 (N_4790,N_1746,N_2782);
or U4791 (N_4791,N_2180,N_534);
and U4792 (N_4792,N_2726,N_1418);
nor U4793 (N_4793,N_1284,N_549);
or U4794 (N_4794,N_1080,N_845);
xnor U4795 (N_4795,N_2554,N_410);
xor U4796 (N_4796,N_1282,N_679);
nand U4797 (N_4797,N_2524,N_417);
and U4798 (N_4798,N_1069,N_2894);
or U4799 (N_4799,N_2457,N_3050);
nand U4800 (N_4800,N_2522,N_1463);
nor U4801 (N_4801,N_468,N_2088);
nor U4802 (N_4802,N_2107,N_2291);
and U4803 (N_4803,N_2118,N_808);
and U4804 (N_4804,N_588,N_2509);
or U4805 (N_4805,N_1575,N_2147);
and U4806 (N_4806,N_2170,N_230);
xor U4807 (N_4807,N_199,N_2225);
nor U4808 (N_4808,N_858,N_293);
nand U4809 (N_4809,N_3037,N_890);
and U4810 (N_4810,N_440,N_125);
nand U4811 (N_4811,N_410,N_98);
nor U4812 (N_4812,N_2476,N_2433);
nor U4813 (N_4813,N_253,N_1983);
or U4814 (N_4814,N_2004,N_1377);
xnor U4815 (N_4815,N_3114,N_2141);
nor U4816 (N_4816,N_2276,N_1465);
nor U4817 (N_4817,N_1411,N_1622);
or U4818 (N_4818,N_717,N_1074);
or U4819 (N_4819,N_1395,N_344);
nand U4820 (N_4820,N_2003,N_2732);
and U4821 (N_4821,N_460,N_52);
and U4822 (N_4822,N_2696,N_2132);
nand U4823 (N_4823,N_3083,N_1198);
and U4824 (N_4824,N_2861,N_1514);
and U4825 (N_4825,N_35,N_846);
and U4826 (N_4826,N_1577,N_1627);
or U4827 (N_4827,N_2600,N_2438);
and U4828 (N_4828,N_1331,N_864);
or U4829 (N_4829,N_2857,N_1110);
or U4830 (N_4830,N_2707,N_3002);
xor U4831 (N_4831,N_2383,N_1949);
or U4832 (N_4832,N_1295,N_2442);
nor U4833 (N_4833,N_2736,N_1919);
nor U4834 (N_4834,N_2174,N_1635);
nor U4835 (N_4835,N_173,N_2008);
and U4836 (N_4836,N_1956,N_2285);
or U4837 (N_4837,N_2770,N_2076);
nand U4838 (N_4838,N_2568,N_1060);
xnor U4839 (N_4839,N_1629,N_2070);
or U4840 (N_4840,N_355,N_1689);
and U4841 (N_4841,N_2475,N_2392);
and U4842 (N_4842,N_2000,N_2293);
nand U4843 (N_4843,N_1681,N_1479);
or U4844 (N_4844,N_1951,N_410);
or U4845 (N_4845,N_913,N_901);
and U4846 (N_4846,N_2274,N_2823);
xor U4847 (N_4847,N_1509,N_823);
and U4848 (N_4848,N_1378,N_2341);
nor U4849 (N_4849,N_497,N_278);
or U4850 (N_4850,N_996,N_2204);
nor U4851 (N_4851,N_944,N_2623);
or U4852 (N_4852,N_1177,N_2252);
and U4853 (N_4853,N_2117,N_925);
and U4854 (N_4854,N_1320,N_337);
and U4855 (N_4855,N_1791,N_1032);
or U4856 (N_4856,N_772,N_2368);
nor U4857 (N_4857,N_3018,N_1876);
nand U4858 (N_4858,N_1159,N_2408);
or U4859 (N_4859,N_1240,N_1048);
and U4860 (N_4860,N_2861,N_961);
or U4861 (N_4861,N_2420,N_1452);
or U4862 (N_4862,N_732,N_1163);
nor U4863 (N_4863,N_2186,N_2428);
nor U4864 (N_4864,N_2220,N_3117);
nand U4865 (N_4865,N_2308,N_1143);
or U4866 (N_4866,N_139,N_377);
xnor U4867 (N_4867,N_1221,N_2659);
nand U4868 (N_4868,N_2943,N_1253);
and U4869 (N_4869,N_557,N_845);
or U4870 (N_4870,N_2712,N_1704);
and U4871 (N_4871,N_124,N_861);
xnor U4872 (N_4872,N_426,N_2066);
and U4873 (N_4873,N_2469,N_481);
nand U4874 (N_4874,N_1177,N_1882);
nand U4875 (N_4875,N_2912,N_979);
nor U4876 (N_4876,N_2759,N_1226);
or U4877 (N_4877,N_1689,N_2832);
nand U4878 (N_4878,N_2181,N_384);
nand U4879 (N_4879,N_1066,N_1167);
nand U4880 (N_4880,N_1673,N_668);
nand U4881 (N_4881,N_1758,N_1387);
and U4882 (N_4882,N_656,N_429);
nand U4883 (N_4883,N_2526,N_1210);
or U4884 (N_4884,N_627,N_221);
xnor U4885 (N_4885,N_706,N_743);
and U4886 (N_4886,N_655,N_2988);
nor U4887 (N_4887,N_569,N_2244);
or U4888 (N_4888,N_285,N_162);
and U4889 (N_4889,N_2564,N_1981);
xnor U4890 (N_4890,N_871,N_241);
xor U4891 (N_4891,N_1285,N_675);
xor U4892 (N_4892,N_1951,N_818);
or U4893 (N_4893,N_399,N_2407);
nand U4894 (N_4894,N_1404,N_124);
nand U4895 (N_4895,N_1525,N_872);
and U4896 (N_4896,N_725,N_530);
xnor U4897 (N_4897,N_2168,N_98);
or U4898 (N_4898,N_1492,N_1001);
nor U4899 (N_4899,N_1504,N_3008);
nand U4900 (N_4900,N_1309,N_1131);
and U4901 (N_4901,N_1806,N_1584);
nor U4902 (N_4902,N_1810,N_1327);
nand U4903 (N_4903,N_2289,N_524);
nand U4904 (N_4904,N_2658,N_389);
and U4905 (N_4905,N_1641,N_2382);
or U4906 (N_4906,N_2043,N_933);
nor U4907 (N_4907,N_1787,N_2814);
nor U4908 (N_4908,N_1953,N_2096);
nor U4909 (N_4909,N_2367,N_3031);
or U4910 (N_4910,N_925,N_425);
and U4911 (N_4911,N_294,N_894);
and U4912 (N_4912,N_1997,N_695);
or U4913 (N_4913,N_2452,N_1151);
nor U4914 (N_4914,N_2441,N_1479);
nand U4915 (N_4915,N_576,N_1717);
xnor U4916 (N_4916,N_1437,N_890);
or U4917 (N_4917,N_3065,N_3028);
nand U4918 (N_4918,N_1989,N_1920);
or U4919 (N_4919,N_1632,N_1038);
and U4920 (N_4920,N_882,N_2340);
xor U4921 (N_4921,N_2721,N_2139);
xnor U4922 (N_4922,N_116,N_226);
nand U4923 (N_4923,N_1830,N_914);
nor U4924 (N_4924,N_2988,N_2432);
nand U4925 (N_4925,N_2087,N_2042);
or U4926 (N_4926,N_2358,N_390);
or U4927 (N_4927,N_364,N_1715);
or U4928 (N_4928,N_2755,N_1012);
and U4929 (N_4929,N_2277,N_1227);
nor U4930 (N_4930,N_2,N_647);
nand U4931 (N_4931,N_2571,N_1633);
and U4932 (N_4932,N_169,N_2609);
nand U4933 (N_4933,N_7,N_2498);
nor U4934 (N_4934,N_914,N_2809);
nand U4935 (N_4935,N_991,N_2481);
and U4936 (N_4936,N_1742,N_118);
nor U4937 (N_4937,N_705,N_1874);
nor U4938 (N_4938,N_1080,N_2667);
xor U4939 (N_4939,N_1302,N_954);
nor U4940 (N_4940,N_2816,N_1701);
nor U4941 (N_4941,N_271,N_2031);
or U4942 (N_4942,N_1876,N_2802);
xor U4943 (N_4943,N_2110,N_332);
or U4944 (N_4944,N_2574,N_421);
nand U4945 (N_4945,N_2574,N_2830);
nor U4946 (N_4946,N_2970,N_2764);
nor U4947 (N_4947,N_2747,N_1206);
and U4948 (N_4948,N_239,N_188);
xor U4949 (N_4949,N_2973,N_227);
and U4950 (N_4950,N_2014,N_1066);
and U4951 (N_4951,N_2687,N_378);
xnor U4952 (N_4952,N_2595,N_1752);
or U4953 (N_4953,N_786,N_1620);
or U4954 (N_4954,N_330,N_2767);
and U4955 (N_4955,N_2882,N_1759);
or U4956 (N_4956,N_2172,N_1555);
nand U4957 (N_4957,N_834,N_503);
or U4958 (N_4958,N_2699,N_1207);
nand U4959 (N_4959,N_1369,N_1322);
and U4960 (N_4960,N_1055,N_23);
or U4961 (N_4961,N_1548,N_397);
and U4962 (N_4962,N_1415,N_678);
xnor U4963 (N_4963,N_2885,N_519);
nand U4964 (N_4964,N_2795,N_1933);
or U4965 (N_4965,N_1579,N_2718);
or U4966 (N_4966,N_1697,N_2701);
nor U4967 (N_4967,N_1221,N_1301);
nand U4968 (N_4968,N_568,N_3093);
nand U4969 (N_4969,N_1529,N_27);
nor U4970 (N_4970,N_1846,N_2703);
nor U4971 (N_4971,N_1874,N_2662);
or U4972 (N_4972,N_2362,N_1991);
or U4973 (N_4973,N_728,N_785);
nor U4974 (N_4974,N_200,N_2695);
or U4975 (N_4975,N_169,N_2433);
and U4976 (N_4976,N_2759,N_2772);
nand U4977 (N_4977,N_2374,N_1609);
nand U4978 (N_4978,N_2078,N_2311);
nor U4979 (N_4979,N_807,N_1476);
or U4980 (N_4980,N_1690,N_1883);
nor U4981 (N_4981,N_2909,N_2984);
xnor U4982 (N_4982,N_482,N_1294);
or U4983 (N_4983,N_2659,N_471);
nand U4984 (N_4984,N_2081,N_3004);
and U4985 (N_4985,N_1156,N_2228);
or U4986 (N_4986,N_2546,N_1914);
or U4987 (N_4987,N_613,N_1136);
nor U4988 (N_4988,N_2918,N_2947);
xnor U4989 (N_4989,N_476,N_2325);
xnor U4990 (N_4990,N_2182,N_2632);
nand U4991 (N_4991,N_1723,N_1027);
nor U4992 (N_4992,N_311,N_1809);
xor U4993 (N_4993,N_2215,N_1781);
nor U4994 (N_4994,N_1661,N_1458);
and U4995 (N_4995,N_240,N_1894);
nor U4996 (N_4996,N_2141,N_213);
or U4997 (N_4997,N_1012,N_3106);
xor U4998 (N_4998,N_2049,N_2717);
and U4999 (N_4999,N_98,N_2052);
nand U5000 (N_5000,N_480,N_2957);
nor U5001 (N_5001,N_2840,N_1642);
nor U5002 (N_5002,N_415,N_2077);
nand U5003 (N_5003,N_1222,N_2296);
xnor U5004 (N_5004,N_2750,N_1522);
nand U5005 (N_5005,N_2202,N_2499);
or U5006 (N_5006,N_1073,N_144);
xor U5007 (N_5007,N_2729,N_1676);
nand U5008 (N_5008,N_397,N_1146);
nor U5009 (N_5009,N_2954,N_1127);
and U5010 (N_5010,N_1151,N_877);
nand U5011 (N_5011,N_2708,N_1797);
or U5012 (N_5012,N_1096,N_558);
nor U5013 (N_5013,N_536,N_740);
or U5014 (N_5014,N_1363,N_2515);
nor U5015 (N_5015,N_2869,N_2209);
nand U5016 (N_5016,N_65,N_1493);
and U5017 (N_5017,N_2010,N_305);
nand U5018 (N_5018,N_1341,N_1930);
and U5019 (N_5019,N_359,N_1578);
or U5020 (N_5020,N_1924,N_671);
nand U5021 (N_5021,N_2277,N_793);
nand U5022 (N_5022,N_582,N_1821);
nand U5023 (N_5023,N_1785,N_1002);
xor U5024 (N_5024,N_240,N_2157);
nand U5025 (N_5025,N_1629,N_2701);
or U5026 (N_5026,N_1403,N_1925);
nand U5027 (N_5027,N_2328,N_2373);
nand U5028 (N_5028,N_534,N_2226);
and U5029 (N_5029,N_2676,N_1363);
nor U5030 (N_5030,N_1266,N_2977);
or U5031 (N_5031,N_2850,N_1899);
xnor U5032 (N_5032,N_2019,N_2981);
nand U5033 (N_5033,N_1793,N_2211);
or U5034 (N_5034,N_577,N_805);
nand U5035 (N_5035,N_939,N_2094);
nand U5036 (N_5036,N_1826,N_2671);
nor U5037 (N_5037,N_1888,N_292);
nand U5038 (N_5038,N_1089,N_2357);
or U5039 (N_5039,N_1963,N_815);
nand U5040 (N_5040,N_2308,N_1565);
and U5041 (N_5041,N_2697,N_2877);
or U5042 (N_5042,N_2136,N_500);
nand U5043 (N_5043,N_1159,N_658);
nor U5044 (N_5044,N_2514,N_2996);
and U5045 (N_5045,N_3120,N_922);
or U5046 (N_5046,N_2322,N_886);
nand U5047 (N_5047,N_1836,N_238);
and U5048 (N_5048,N_2956,N_1505);
nor U5049 (N_5049,N_2118,N_2683);
xnor U5050 (N_5050,N_549,N_2661);
nor U5051 (N_5051,N_395,N_1903);
and U5052 (N_5052,N_112,N_1141);
or U5053 (N_5053,N_2426,N_2725);
or U5054 (N_5054,N_1880,N_2237);
or U5055 (N_5055,N_2868,N_2328);
and U5056 (N_5056,N_457,N_788);
xor U5057 (N_5057,N_1246,N_1258);
nor U5058 (N_5058,N_781,N_1747);
or U5059 (N_5059,N_655,N_2982);
nor U5060 (N_5060,N_1118,N_1117);
nor U5061 (N_5061,N_1991,N_2809);
nand U5062 (N_5062,N_108,N_1056);
or U5063 (N_5063,N_3035,N_1247);
and U5064 (N_5064,N_2751,N_327);
nor U5065 (N_5065,N_2202,N_3049);
nand U5066 (N_5066,N_2034,N_2777);
nand U5067 (N_5067,N_2485,N_1171);
nor U5068 (N_5068,N_270,N_2503);
nor U5069 (N_5069,N_1665,N_555);
nor U5070 (N_5070,N_217,N_1093);
nand U5071 (N_5071,N_1844,N_182);
xor U5072 (N_5072,N_1176,N_1897);
or U5073 (N_5073,N_226,N_2984);
nand U5074 (N_5074,N_927,N_1831);
and U5075 (N_5075,N_551,N_2405);
and U5076 (N_5076,N_765,N_1224);
or U5077 (N_5077,N_120,N_573);
nand U5078 (N_5078,N_1485,N_1205);
xor U5079 (N_5079,N_2673,N_2310);
nor U5080 (N_5080,N_2852,N_2752);
nand U5081 (N_5081,N_1241,N_1660);
xnor U5082 (N_5082,N_1053,N_2834);
nor U5083 (N_5083,N_390,N_2073);
and U5084 (N_5084,N_2167,N_2492);
or U5085 (N_5085,N_2674,N_220);
xnor U5086 (N_5086,N_3063,N_3014);
and U5087 (N_5087,N_178,N_990);
xor U5088 (N_5088,N_2319,N_565);
nor U5089 (N_5089,N_2737,N_784);
or U5090 (N_5090,N_1497,N_2027);
nand U5091 (N_5091,N_2557,N_2903);
nand U5092 (N_5092,N_2554,N_2294);
nand U5093 (N_5093,N_2951,N_1269);
or U5094 (N_5094,N_295,N_3038);
xnor U5095 (N_5095,N_2931,N_1363);
and U5096 (N_5096,N_3077,N_2552);
nand U5097 (N_5097,N_2983,N_1538);
or U5098 (N_5098,N_101,N_575);
and U5099 (N_5099,N_2594,N_2702);
nand U5100 (N_5100,N_2151,N_2880);
and U5101 (N_5101,N_1596,N_711);
and U5102 (N_5102,N_2743,N_2151);
and U5103 (N_5103,N_2750,N_827);
or U5104 (N_5104,N_1102,N_781);
and U5105 (N_5105,N_2478,N_385);
nor U5106 (N_5106,N_530,N_2509);
nand U5107 (N_5107,N_2829,N_2045);
and U5108 (N_5108,N_2043,N_2629);
nand U5109 (N_5109,N_1747,N_1627);
and U5110 (N_5110,N_2171,N_1498);
nor U5111 (N_5111,N_1527,N_1751);
nand U5112 (N_5112,N_932,N_518);
nor U5113 (N_5113,N_279,N_120);
nand U5114 (N_5114,N_1687,N_931);
nand U5115 (N_5115,N_1303,N_2721);
or U5116 (N_5116,N_2796,N_587);
xnor U5117 (N_5117,N_3007,N_630);
or U5118 (N_5118,N_702,N_2209);
nand U5119 (N_5119,N_961,N_1406);
and U5120 (N_5120,N_3043,N_1083);
and U5121 (N_5121,N_1482,N_156);
nor U5122 (N_5122,N_2462,N_2386);
nand U5123 (N_5123,N_788,N_233);
nand U5124 (N_5124,N_1651,N_3094);
and U5125 (N_5125,N_1206,N_31);
and U5126 (N_5126,N_1186,N_275);
nand U5127 (N_5127,N_2463,N_2053);
or U5128 (N_5128,N_432,N_3057);
nand U5129 (N_5129,N_2642,N_2761);
nor U5130 (N_5130,N_2661,N_1247);
or U5131 (N_5131,N_2038,N_2028);
or U5132 (N_5132,N_2652,N_1824);
nor U5133 (N_5133,N_104,N_846);
nor U5134 (N_5134,N_625,N_2799);
nand U5135 (N_5135,N_312,N_654);
nand U5136 (N_5136,N_1934,N_2439);
xnor U5137 (N_5137,N_1197,N_30);
or U5138 (N_5138,N_135,N_1988);
or U5139 (N_5139,N_1557,N_2433);
nand U5140 (N_5140,N_2255,N_9);
nand U5141 (N_5141,N_1453,N_1170);
nand U5142 (N_5142,N_2564,N_1881);
and U5143 (N_5143,N_947,N_194);
nor U5144 (N_5144,N_2019,N_1395);
nor U5145 (N_5145,N_2857,N_588);
and U5146 (N_5146,N_2919,N_1004);
or U5147 (N_5147,N_1768,N_862);
nor U5148 (N_5148,N_2174,N_2812);
or U5149 (N_5149,N_2540,N_1131);
and U5150 (N_5150,N_2074,N_118);
xor U5151 (N_5151,N_2126,N_1251);
nor U5152 (N_5152,N_1329,N_36);
nand U5153 (N_5153,N_2751,N_1446);
and U5154 (N_5154,N_1674,N_1050);
nor U5155 (N_5155,N_2855,N_1179);
nand U5156 (N_5156,N_409,N_344);
nor U5157 (N_5157,N_1158,N_2463);
and U5158 (N_5158,N_443,N_2414);
or U5159 (N_5159,N_1911,N_630);
and U5160 (N_5160,N_2064,N_2465);
and U5161 (N_5161,N_2483,N_2769);
nand U5162 (N_5162,N_318,N_2622);
nand U5163 (N_5163,N_274,N_2962);
nand U5164 (N_5164,N_2995,N_2800);
and U5165 (N_5165,N_2827,N_703);
nor U5166 (N_5166,N_1704,N_490);
and U5167 (N_5167,N_2204,N_985);
or U5168 (N_5168,N_668,N_1224);
nor U5169 (N_5169,N_1646,N_1227);
and U5170 (N_5170,N_1887,N_482);
nand U5171 (N_5171,N_2591,N_611);
and U5172 (N_5172,N_632,N_245);
nand U5173 (N_5173,N_1754,N_2384);
nand U5174 (N_5174,N_2831,N_1496);
or U5175 (N_5175,N_149,N_1952);
and U5176 (N_5176,N_737,N_1676);
nand U5177 (N_5177,N_2385,N_116);
nand U5178 (N_5178,N_2121,N_1515);
nand U5179 (N_5179,N_983,N_812);
nand U5180 (N_5180,N_1571,N_2298);
nor U5181 (N_5181,N_1791,N_2587);
and U5182 (N_5182,N_841,N_675);
and U5183 (N_5183,N_2064,N_492);
or U5184 (N_5184,N_1663,N_1097);
nand U5185 (N_5185,N_747,N_1906);
or U5186 (N_5186,N_2680,N_2201);
nor U5187 (N_5187,N_1091,N_1042);
nor U5188 (N_5188,N_301,N_932);
and U5189 (N_5189,N_1228,N_637);
or U5190 (N_5190,N_1960,N_1425);
xnor U5191 (N_5191,N_2425,N_1546);
nand U5192 (N_5192,N_1646,N_2911);
nand U5193 (N_5193,N_597,N_653);
or U5194 (N_5194,N_555,N_411);
and U5195 (N_5195,N_2423,N_2969);
and U5196 (N_5196,N_2449,N_3102);
nor U5197 (N_5197,N_2684,N_1702);
and U5198 (N_5198,N_1231,N_2705);
and U5199 (N_5199,N_2233,N_2776);
nor U5200 (N_5200,N_1908,N_2444);
nand U5201 (N_5201,N_1366,N_665);
nor U5202 (N_5202,N_1282,N_1911);
nand U5203 (N_5203,N_1088,N_2298);
nand U5204 (N_5204,N_2093,N_1488);
nor U5205 (N_5205,N_1527,N_1806);
and U5206 (N_5206,N_2656,N_2376);
nand U5207 (N_5207,N_1123,N_1047);
nand U5208 (N_5208,N_203,N_678);
nand U5209 (N_5209,N_1926,N_2558);
or U5210 (N_5210,N_2348,N_1140);
nand U5211 (N_5211,N_2494,N_285);
xnor U5212 (N_5212,N_486,N_1354);
and U5213 (N_5213,N_2324,N_2782);
or U5214 (N_5214,N_619,N_2538);
or U5215 (N_5215,N_108,N_1657);
nor U5216 (N_5216,N_943,N_2576);
and U5217 (N_5217,N_449,N_314);
nand U5218 (N_5218,N_228,N_542);
and U5219 (N_5219,N_3,N_132);
and U5220 (N_5220,N_1086,N_1078);
or U5221 (N_5221,N_945,N_773);
nand U5222 (N_5222,N_251,N_2989);
nor U5223 (N_5223,N_1929,N_2738);
nand U5224 (N_5224,N_1759,N_2076);
or U5225 (N_5225,N_3023,N_2623);
xor U5226 (N_5226,N_2775,N_97);
nand U5227 (N_5227,N_2884,N_2942);
and U5228 (N_5228,N_1512,N_1560);
nand U5229 (N_5229,N_1332,N_1188);
nand U5230 (N_5230,N_1221,N_1262);
nor U5231 (N_5231,N_1180,N_2310);
nand U5232 (N_5232,N_1262,N_2101);
nand U5233 (N_5233,N_1806,N_1510);
and U5234 (N_5234,N_2285,N_2059);
nor U5235 (N_5235,N_49,N_1585);
and U5236 (N_5236,N_3062,N_874);
nand U5237 (N_5237,N_612,N_532);
or U5238 (N_5238,N_2329,N_982);
nand U5239 (N_5239,N_1225,N_808);
nor U5240 (N_5240,N_2364,N_2319);
or U5241 (N_5241,N_492,N_432);
and U5242 (N_5242,N_936,N_2295);
or U5243 (N_5243,N_2157,N_1904);
and U5244 (N_5244,N_1455,N_1012);
nand U5245 (N_5245,N_844,N_854);
or U5246 (N_5246,N_1198,N_2258);
nor U5247 (N_5247,N_499,N_1756);
and U5248 (N_5248,N_1098,N_2802);
nor U5249 (N_5249,N_86,N_2563);
or U5250 (N_5250,N_2842,N_2446);
and U5251 (N_5251,N_422,N_2970);
nor U5252 (N_5252,N_2034,N_2347);
xnor U5253 (N_5253,N_1566,N_107);
and U5254 (N_5254,N_725,N_3021);
xor U5255 (N_5255,N_1038,N_2422);
or U5256 (N_5256,N_1587,N_1512);
nand U5257 (N_5257,N_990,N_163);
or U5258 (N_5258,N_2366,N_735);
nand U5259 (N_5259,N_2770,N_347);
and U5260 (N_5260,N_95,N_1528);
xnor U5261 (N_5261,N_1617,N_2098);
or U5262 (N_5262,N_1295,N_510);
and U5263 (N_5263,N_1261,N_2349);
and U5264 (N_5264,N_111,N_745);
xor U5265 (N_5265,N_997,N_689);
nand U5266 (N_5266,N_209,N_1942);
nor U5267 (N_5267,N_1244,N_2302);
nor U5268 (N_5268,N_2635,N_262);
and U5269 (N_5269,N_224,N_705);
or U5270 (N_5270,N_1812,N_2212);
and U5271 (N_5271,N_108,N_779);
and U5272 (N_5272,N_458,N_2463);
and U5273 (N_5273,N_2817,N_2527);
or U5274 (N_5274,N_877,N_2205);
nand U5275 (N_5275,N_778,N_2759);
nor U5276 (N_5276,N_3061,N_1831);
nand U5277 (N_5277,N_3036,N_2406);
and U5278 (N_5278,N_1829,N_581);
or U5279 (N_5279,N_724,N_2547);
and U5280 (N_5280,N_441,N_2096);
nor U5281 (N_5281,N_2222,N_425);
and U5282 (N_5282,N_3109,N_607);
nor U5283 (N_5283,N_629,N_517);
or U5284 (N_5284,N_2673,N_1740);
nor U5285 (N_5285,N_1318,N_1030);
or U5286 (N_5286,N_230,N_613);
nor U5287 (N_5287,N_1189,N_928);
and U5288 (N_5288,N_434,N_1926);
and U5289 (N_5289,N_2362,N_1293);
nor U5290 (N_5290,N_3017,N_3091);
and U5291 (N_5291,N_2358,N_634);
nor U5292 (N_5292,N_969,N_324);
or U5293 (N_5293,N_2341,N_2079);
or U5294 (N_5294,N_2178,N_1292);
nand U5295 (N_5295,N_1549,N_2823);
xnor U5296 (N_5296,N_2853,N_1803);
nand U5297 (N_5297,N_486,N_1602);
and U5298 (N_5298,N_2330,N_3046);
nand U5299 (N_5299,N_1639,N_3022);
nor U5300 (N_5300,N_2576,N_1850);
nor U5301 (N_5301,N_2981,N_1681);
nor U5302 (N_5302,N_836,N_642);
and U5303 (N_5303,N_574,N_479);
nand U5304 (N_5304,N_838,N_2725);
nand U5305 (N_5305,N_1093,N_1768);
nand U5306 (N_5306,N_498,N_2833);
and U5307 (N_5307,N_2908,N_620);
or U5308 (N_5308,N_1223,N_2654);
and U5309 (N_5309,N_1777,N_225);
or U5310 (N_5310,N_2850,N_914);
xor U5311 (N_5311,N_824,N_646);
nand U5312 (N_5312,N_2883,N_2563);
nor U5313 (N_5313,N_1928,N_805);
nand U5314 (N_5314,N_1210,N_1086);
xor U5315 (N_5315,N_2155,N_2911);
nand U5316 (N_5316,N_845,N_2201);
and U5317 (N_5317,N_2221,N_3108);
and U5318 (N_5318,N_189,N_2694);
or U5319 (N_5319,N_2355,N_1086);
nor U5320 (N_5320,N_2649,N_2425);
or U5321 (N_5321,N_2451,N_1794);
or U5322 (N_5322,N_2980,N_735);
or U5323 (N_5323,N_178,N_922);
nand U5324 (N_5324,N_1746,N_843);
and U5325 (N_5325,N_1539,N_2962);
nand U5326 (N_5326,N_1022,N_1206);
and U5327 (N_5327,N_227,N_1393);
nand U5328 (N_5328,N_1796,N_58);
and U5329 (N_5329,N_2975,N_622);
nor U5330 (N_5330,N_330,N_2049);
nand U5331 (N_5331,N_2556,N_1625);
xnor U5332 (N_5332,N_1907,N_368);
and U5333 (N_5333,N_1691,N_1168);
nor U5334 (N_5334,N_2892,N_652);
nor U5335 (N_5335,N_2498,N_747);
nor U5336 (N_5336,N_2830,N_3014);
or U5337 (N_5337,N_1410,N_2753);
and U5338 (N_5338,N_367,N_738);
xor U5339 (N_5339,N_2238,N_1273);
xor U5340 (N_5340,N_1143,N_1950);
nor U5341 (N_5341,N_2063,N_1015);
nand U5342 (N_5342,N_1673,N_922);
nor U5343 (N_5343,N_820,N_888);
or U5344 (N_5344,N_2144,N_3056);
xor U5345 (N_5345,N_1287,N_1914);
nand U5346 (N_5346,N_594,N_1946);
nand U5347 (N_5347,N_278,N_1959);
nand U5348 (N_5348,N_532,N_2923);
nor U5349 (N_5349,N_514,N_2823);
nor U5350 (N_5350,N_2486,N_2909);
or U5351 (N_5351,N_1532,N_1735);
or U5352 (N_5352,N_965,N_1511);
and U5353 (N_5353,N_1861,N_1479);
nand U5354 (N_5354,N_1880,N_1218);
nand U5355 (N_5355,N_1224,N_190);
and U5356 (N_5356,N_1205,N_1071);
and U5357 (N_5357,N_139,N_503);
or U5358 (N_5358,N_1650,N_61);
and U5359 (N_5359,N_2745,N_62);
nor U5360 (N_5360,N_173,N_2795);
nor U5361 (N_5361,N_861,N_865);
nor U5362 (N_5362,N_1188,N_2029);
xnor U5363 (N_5363,N_1671,N_491);
or U5364 (N_5364,N_593,N_1813);
or U5365 (N_5365,N_299,N_2525);
and U5366 (N_5366,N_357,N_2563);
nor U5367 (N_5367,N_2896,N_2124);
nor U5368 (N_5368,N_17,N_2491);
nor U5369 (N_5369,N_279,N_181);
nand U5370 (N_5370,N_2573,N_1300);
or U5371 (N_5371,N_2206,N_64);
xnor U5372 (N_5372,N_1579,N_594);
xor U5373 (N_5373,N_3088,N_2866);
and U5374 (N_5374,N_2686,N_2770);
or U5375 (N_5375,N_1883,N_557);
nand U5376 (N_5376,N_2752,N_1945);
or U5377 (N_5377,N_1533,N_1515);
or U5378 (N_5378,N_2151,N_2309);
or U5379 (N_5379,N_1800,N_2883);
or U5380 (N_5380,N_771,N_660);
nor U5381 (N_5381,N_1487,N_1750);
xnor U5382 (N_5382,N_323,N_1953);
nor U5383 (N_5383,N_1712,N_1251);
and U5384 (N_5384,N_2731,N_1909);
or U5385 (N_5385,N_673,N_3024);
or U5386 (N_5386,N_720,N_436);
nand U5387 (N_5387,N_3031,N_1309);
or U5388 (N_5388,N_980,N_2574);
or U5389 (N_5389,N_529,N_2920);
nor U5390 (N_5390,N_2857,N_404);
nand U5391 (N_5391,N_643,N_1752);
and U5392 (N_5392,N_3094,N_2461);
and U5393 (N_5393,N_1431,N_1293);
and U5394 (N_5394,N_209,N_358);
and U5395 (N_5395,N_593,N_328);
nand U5396 (N_5396,N_1776,N_1691);
and U5397 (N_5397,N_1355,N_833);
nor U5398 (N_5398,N_754,N_109);
nand U5399 (N_5399,N_2410,N_1937);
nor U5400 (N_5400,N_1083,N_2393);
nand U5401 (N_5401,N_278,N_3031);
nand U5402 (N_5402,N_625,N_539);
xor U5403 (N_5403,N_2635,N_1656);
xnor U5404 (N_5404,N_2112,N_685);
nor U5405 (N_5405,N_1374,N_1801);
nor U5406 (N_5406,N_2591,N_1002);
nor U5407 (N_5407,N_1166,N_238);
nor U5408 (N_5408,N_2289,N_265);
nor U5409 (N_5409,N_985,N_2577);
nor U5410 (N_5410,N_1333,N_2281);
nand U5411 (N_5411,N_2838,N_2396);
and U5412 (N_5412,N_2085,N_1644);
nand U5413 (N_5413,N_595,N_2853);
nand U5414 (N_5414,N_2042,N_863);
nand U5415 (N_5415,N_629,N_2766);
and U5416 (N_5416,N_320,N_722);
xnor U5417 (N_5417,N_2889,N_1802);
nor U5418 (N_5418,N_1553,N_2525);
nor U5419 (N_5419,N_2227,N_2307);
and U5420 (N_5420,N_48,N_309);
and U5421 (N_5421,N_495,N_1100);
and U5422 (N_5422,N_2013,N_1096);
nor U5423 (N_5423,N_273,N_945);
nor U5424 (N_5424,N_2769,N_2244);
nand U5425 (N_5425,N_2855,N_2219);
or U5426 (N_5426,N_1287,N_319);
nand U5427 (N_5427,N_364,N_3104);
nor U5428 (N_5428,N_863,N_907);
xnor U5429 (N_5429,N_1680,N_224);
nor U5430 (N_5430,N_1951,N_789);
nand U5431 (N_5431,N_1751,N_2508);
nor U5432 (N_5432,N_2743,N_2635);
xnor U5433 (N_5433,N_52,N_316);
and U5434 (N_5434,N_182,N_2837);
nor U5435 (N_5435,N_2757,N_283);
nor U5436 (N_5436,N_1244,N_2128);
nor U5437 (N_5437,N_1092,N_1438);
xnor U5438 (N_5438,N_554,N_2378);
or U5439 (N_5439,N_1277,N_1619);
or U5440 (N_5440,N_2494,N_43);
or U5441 (N_5441,N_1762,N_1979);
or U5442 (N_5442,N_584,N_1615);
nor U5443 (N_5443,N_2351,N_637);
and U5444 (N_5444,N_2268,N_245);
or U5445 (N_5445,N_1084,N_3031);
or U5446 (N_5446,N_336,N_1438);
nor U5447 (N_5447,N_1756,N_2700);
nor U5448 (N_5448,N_1584,N_294);
and U5449 (N_5449,N_1297,N_2226);
nand U5450 (N_5450,N_2109,N_953);
nor U5451 (N_5451,N_2938,N_685);
or U5452 (N_5452,N_1629,N_1276);
or U5453 (N_5453,N_682,N_2532);
or U5454 (N_5454,N_974,N_1034);
xnor U5455 (N_5455,N_2324,N_1254);
or U5456 (N_5456,N_1751,N_1956);
nor U5457 (N_5457,N_2206,N_1920);
nor U5458 (N_5458,N_1769,N_2161);
xnor U5459 (N_5459,N_1260,N_679);
nor U5460 (N_5460,N_2319,N_77);
nor U5461 (N_5461,N_650,N_646);
nand U5462 (N_5462,N_221,N_2962);
and U5463 (N_5463,N_2903,N_684);
nor U5464 (N_5464,N_232,N_2263);
and U5465 (N_5465,N_2886,N_882);
or U5466 (N_5466,N_2806,N_2419);
nor U5467 (N_5467,N_1469,N_1348);
or U5468 (N_5468,N_1604,N_2306);
nand U5469 (N_5469,N_486,N_2717);
or U5470 (N_5470,N_403,N_2203);
nand U5471 (N_5471,N_818,N_2059);
nand U5472 (N_5472,N_195,N_981);
xnor U5473 (N_5473,N_126,N_901);
xnor U5474 (N_5474,N_1495,N_1104);
or U5475 (N_5475,N_2385,N_1267);
nor U5476 (N_5476,N_1229,N_2598);
nand U5477 (N_5477,N_1687,N_138);
or U5478 (N_5478,N_1096,N_992);
nor U5479 (N_5479,N_1420,N_2405);
and U5480 (N_5480,N_788,N_669);
or U5481 (N_5481,N_1579,N_295);
nand U5482 (N_5482,N_3016,N_1276);
and U5483 (N_5483,N_1173,N_703);
nor U5484 (N_5484,N_34,N_3103);
and U5485 (N_5485,N_1927,N_3055);
xnor U5486 (N_5486,N_2926,N_502);
and U5487 (N_5487,N_2560,N_647);
nor U5488 (N_5488,N_641,N_2334);
or U5489 (N_5489,N_1592,N_2226);
or U5490 (N_5490,N_591,N_1507);
xnor U5491 (N_5491,N_923,N_233);
nand U5492 (N_5492,N_2919,N_1930);
nor U5493 (N_5493,N_37,N_706);
or U5494 (N_5494,N_1789,N_409);
xor U5495 (N_5495,N_92,N_1147);
xnor U5496 (N_5496,N_2539,N_855);
nand U5497 (N_5497,N_2829,N_368);
and U5498 (N_5498,N_1257,N_2690);
xnor U5499 (N_5499,N_2038,N_334);
nor U5500 (N_5500,N_921,N_474);
and U5501 (N_5501,N_2388,N_2771);
xnor U5502 (N_5502,N_427,N_2875);
or U5503 (N_5503,N_993,N_8);
and U5504 (N_5504,N_2649,N_2467);
and U5505 (N_5505,N_146,N_1469);
xor U5506 (N_5506,N_1325,N_1964);
nor U5507 (N_5507,N_2805,N_746);
nand U5508 (N_5508,N_2726,N_856);
xnor U5509 (N_5509,N_2480,N_2244);
nand U5510 (N_5510,N_1646,N_629);
and U5511 (N_5511,N_2367,N_483);
and U5512 (N_5512,N_348,N_2915);
or U5513 (N_5513,N_2860,N_984);
and U5514 (N_5514,N_676,N_1468);
or U5515 (N_5515,N_123,N_572);
nor U5516 (N_5516,N_2950,N_9);
nor U5517 (N_5517,N_1117,N_528);
and U5518 (N_5518,N_2793,N_574);
xor U5519 (N_5519,N_496,N_1093);
nor U5520 (N_5520,N_287,N_385);
nand U5521 (N_5521,N_2126,N_862);
or U5522 (N_5522,N_1930,N_2634);
and U5523 (N_5523,N_386,N_1435);
nand U5524 (N_5524,N_1797,N_551);
or U5525 (N_5525,N_2994,N_1860);
nor U5526 (N_5526,N_1666,N_692);
nor U5527 (N_5527,N_241,N_1372);
xnor U5528 (N_5528,N_372,N_2349);
and U5529 (N_5529,N_866,N_3043);
or U5530 (N_5530,N_3091,N_2095);
nor U5531 (N_5531,N_3022,N_234);
and U5532 (N_5532,N_2915,N_511);
or U5533 (N_5533,N_450,N_3102);
xor U5534 (N_5534,N_1063,N_835);
and U5535 (N_5535,N_670,N_3059);
nand U5536 (N_5536,N_2646,N_1665);
nor U5537 (N_5537,N_1723,N_1775);
and U5538 (N_5538,N_1985,N_1168);
nor U5539 (N_5539,N_2492,N_575);
or U5540 (N_5540,N_2732,N_2476);
and U5541 (N_5541,N_1064,N_242);
or U5542 (N_5542,N_1032,N_2859);
nor U5543 (N_5543,N_2805,N_2282);
or U5544 (N_5544,N_2909,N_1681);
and U5545 (N_5545,N_469,N_2550);
nor U5546 (N_5546,N_2022,N_461);
xnor U5547 (N_5547,N_691,N_1577);
and U5548 (N_5548,N_442,N_306);
or U5549 (N_5549,N_1219,N_1837);
or U5550 (N_5550,N_2753,N_389);
and U5551 (N_5551,N_733,N_2380);
and U5552 (N_5552,N_286,N_541);
nor U5553 (N_5553,N_95,N_2183);
or U5554 (N_5554,N_2782,N_3046);
or U5555 (N_5555,N_202,N_2108);
or U5556 (N_5556,N_539,N_2547);
or U5557 (N_5557,N_1464,N_728);
nand U5558 (N_5558,N_2860,N_3053);
and U5559 (N_5559,N_3094,N_1571);
and U5560 (N_5560,N_1060,N_2564);
and U5561 (N_5561,N_309,N_1492);
nand U5562 (N_5562,N_2498,N_137);
nand U5563 (N_5563,N_440,N_473);
xnor U5564 (N_5564,N_635,N_1869);
and U5565 (N_5565,N_1391,N_1415);
and U5566 (N_5566,N_2735,N_830);
nor U5567 (N_5567,N_2219,N_3048);
nand U5568 (N_5568,N_2311,N_2003);
nor U5569 (N_5569,N_1541,N_2644);
xor U5570 (N_5570,N_322,N_2584);
and U5571 (N_5571,N_1101,N_3069);
or U5572 (N_5572,N_1989,N_2902);
or U5573 (N_5573,N_606,N_432);
nor U5574 (N_5574,N_1685,N_40);
and U5575 (N_5575,N_2724,N_1834);
and U5576 (N_5576,N_2204,N_1268);
and U5577 (N_5577,N_1636,N_2576);
nor U5578 (N_5578,N_459,N_460);
and U5579 (N_5579,N_1140,N_1312);
or U5580 (N_5580,N_2425,N_2752);
nor U5581 (N_5581,N_1101,N_713);
nand U5582 (N_5582,N_2012,N_366);
and U5583 (N_5583,N_1276,N_1183);
nand U5584 (N_5584,N_1984,N_2723);
or U5585 (N_5585,N_2599,N_1808);
xor U5586 (N_5586,N_68,N_623);
nand U5587 (N_5587,N_800,N_1635);
or U5588 (N_5588,N_766,N_2640);
and U5589 (N_5589,N_962,N_1059);
nand U5590 (N_5590,N_1150,N_350);
and U5591 (N_5591,N_2835,N_2745);
nand U5592 (N_5592,N_2204,N_1225);
or U5593 (N_5593,N_23,N_2195);
and U5594 (N_5594,N_2101,N_1903);
nor U5595 (N_5595,N_2625,N_2416);
nor U5596 (N_5596,N_306,N_1423);
nand U5597 (N_5597,N_977,N_774);
and U5598 (N_5598,N_1349,N_2955);
and U5599 (N_5599,N_448,N_237);
nor U5600 (N_5600,N_1668,N_2347);
nor U5601 (N_5601,N_966,N_1437);
xor U5602 (N_5602,N_2511,N_1209);
and U5603 (N_5603,N_1839,N_2584);
or U5604 (N_5604,N_556,N_328);
or U5605 (N_5605,N_845,N_2475);
and U5606 (N_5606,N_727,N_542);
or U5607 (N_5607,N_2310,N_2745);
nor U5608 (N_5608,N_1540,N_1449);
nand U5609 (N_5609,N_1586,N_1767);
nor U5610 (N_5610,N_51,N_1688);
or U5611 (N_5611,N_39,N_383);
or U5612 (N_5612,N_945,N_1022);
nor U5613 (N_5613,N_1392,N_1996);
nand U5614 (N_5614,N_1692,N_313);
nor U5615 (N_5615,N_2362,N_999);
and U5616 (N_5616,N_1973,N_1060);
and U5617 (N_5617,N_3099,N_1596);
or U5618 (N_5618,N_96,N_2245);
and U5619 (N_5619,N_1705,N_1457);
nand U5620 (N_5620,N_1813,N_2228);
and U5621 (N_5621,N_1043,N_1041);
and U5622 (N_5622,N_1637,N_24);
nand U5623 (N_5623,N_1275,N_270);
or U5624 (N_5624,N_3069,N_10);
xor U5625 (N_5625,N_2900,N_2189);
nand U5626 (N_5626,N_2597,N_2953);
and U5627 (N_5627,N_793,N_959);
and U5628 (N_5628,N_668,N_58);
and U5629 (N_5629,N_776,N_2766);
or U5630 (N_5630,N_2094,N_1106);
or U5631 (N_5631,N_686,N_1743);
nand U5632 (N_5632,N_1179,N_657);
or U5633 (N_5633,N_537,N_2853);
or U5634 (N_5634,N_1011,N_832);
nor U5635 (N_5635,N_2898,N_1628);
nor U5636 (N_5636,N_2444,N_2851);
nor U5637 (N_5637,N_1811,N_1813);
nor U5638 (N_5638,N_1436,N_1566);
nand U5639 (N_5639,N_1304,N_819);
nand U5640 (N_5640,N_1120,N_697);
nand U5641 (N_5641,N_448,N_1094);
and U5642 (N_5642,N_836,N_680);
or U5643 (N_5643,N_2893,N_2582);
and U5644 (N_5644,N_1589,N_1336);
and U5645 (N_5645,N_1018,N_3101);
nand U5646 (N_5646,N_2584,N_2471);
and U5647 (N_5647,N_2783,N_2691);
xnor U5648 (N_5648,N_2882,N_353);
or U5649 (N_5649,N_348,N_3017);
xor U5650 (N_5650,N_551,N_113);
nand U5651 (N_5651,N_2346,N_2299);
or U5652 (N_5652,N_2539,N_2188);
or U5653 (N_5653,N_1506,N_1840);
nor U5654 (N_5654,N_2692,N_1524);
or U5655 (N_5655,N_1596,N_721);
or U5656 (N_5656,N_226,N_2118);
or U5657 (N_5657,N_2368,N_1329);
or U5658 (N_5658,N_73,N_2613);
nand U5659 (N_5659,N_2848,N_1982);
nor U5660 (N_5660,N_405,N_2729);
or U5661 (N_5661,N_211,N_178);
nand U5662 (N_5662,N_3080,N_3053);
nand U5663 (N_5663,N_2689,N_398);
and U5664 (N_5664,N_2541,N_177);
nand U5665 (N_5665,N_864,N_1005);
and U5666 (N_5666,N_2813,N_2154);
nand U5667 (N_5667,N_2523,N_938);
and U5668 (N_5668,N_121,N_2592);
and U5669 (N_5669,N_1341,N_748);
and U5670 (N_5670,N_1663,N_1226);
nor U5671 (N_5671,N_28,N_541);
xor U5672 (N_5672,N_2090,N_488);
nor U5673 (N_5673,N_1164,N_1554);
nor U5674 (N_5674,N_1187,N_711);
or U5675 (N_5675,N_1083,N_598);
or U5676 (N_5676,N_335,N_281);
xor U5677 (N_5677,N_592,N_1655);
nand U5678 (N_5678,N_280,N_1072);
and U5679 (N_5679,N_1444,N_1465);
and U5680 (N_5680,N_1473,N_2355);
or U5681 (N_5681,N_2341,N_2131);
nand U5682 (N_5682,N_1028,N_1423);
nand U5683 (N_5683,N_2943,N_869);
nor U5684 (N_5684,N_2654,N_2513);
xor U5685 (N_5685,N_2076,N_607);
nand U5686 (N_5686,N_412,N_717);
nand U5687 (N_5687,N_2,N_3059);
nor U5688 (N_5688,N_1134,N_1262);
or U5689 (N_5689,N_2917,N_1255);
or U5690 (N_5690,N_142,N_373);
nor U5691 (N_5691,N_30,N_2667);
nand U5692 (N_5692,N_1093,N_874);
or U5693 (N_5693,N_1827,N_687);
nand U5694 (N_5694,N_1143,N_2907);
nor U5695 (N_5695,N_291,N_1019);
or U5696 (N_5696,N_83,N_1750);
nand U5697 (N_5697,N_3029,N_2086);
nor U5698 (N_5698,N_223,N_1330);
nand U5699 (N_5699,N_1563,N_2507);
and U5700 (N_5700,N_2881,N_997);
nor U5701 (N_5701,N_1410,N_962);
nand U5702 (N_5702,N_2956,N_1774);
or U5703 (N_5703,N_322,N_2258);
or U5704 (N_5704,N_1369,N_1017);
nand U5705 (N_5705,N_2099,N_2339);
or U5706 (N_5706,N_528,N_571);
and U5707 (N_5707,N_585,N_1933);
nor U5708 (N_5708,N_724,N_689);
nand U5709 (N_5709,N_1480,N_1895);
nor U5710 (N_5710,N_190,N_2325);
nor U5711 (N_5711,N_2361,N_1624);
and U5712 (N_5712,N_1514,N_963);
and U5713 (N_5713,N_1602,N_417);
or U5714 (N_5714,N_782,N_2258);
or U5715 (N_5715,N_2116,N_3022);
nor U5716 (N_5716,N_1080,N_890);
nor U5717 (N_5717,N_2611,N_1745);
xor U5718 (N_5718,N_2724,N_1760);
and U5719 (N_5719,N_2845,N_2317);
nor U5720 (N_5720,N_2087,N_1454);
and U5721 (N_5721,N_1609,N_363);
and U5722 (N_5722,N_467,N_1878);
nand U5723 (N_5723,N_507,N_1407);
nand U5724 (N_5724,N_481,N_684);
nor U5725 (N_5725,N_2386,N_2018);
nor U5726 (N_5726,N_1260,N_1127);
and U5727 (N_5727,N_2279,N_3017);
or U5728 (N_5728,N_2732,N_501);
and U5729 (N_5729,N_391,N_138);
nor U5730 (N_5730,N_2176,N_1734);
or U5731 (N_5731,N_1340,N_2667);
or U5732 (N_5732,N_1478,N_128);
nand U5733 (N_5733,N_1770,N_2964);
nor U5734 (N_5734,N_2452,N_1659);
or U5735 (N_5735,N_2261,N_2694);
nor U5736 (N_5736,N_898,N_885);
nor U5737 (N_5737,N_2652,N_826);
nand U5738 (N_5738,N_67,N_1545);
and U5739 (N_5739,N_1480,N_43);
nor U5740 (N_5740,N_2080,N_3061);
or U5741 (N_5741,N_1347,N_1025);
and U5742 (N_5742,N_2901,N_2768);
and U5743 (N_5743,N_1071,N_2885);
nand U5744 (N_5744,N_2578,N_1124);
nor U5745 (N_5745,N_2008,N_2436);
and U5746 (N_5746,N_375,N_688);
nor U5747 (N_5747,N_1683,N_810);
nor U5748 (N_5748,N_1206,N_2146);
or U5749 (N_5749,N_1489,N_1783);
nand U5750 (N_5750,N_779,N_2307);
xnor U5751 (N_5751,N_1362,N_296);
and U5752 (N_5752,N_2549,N_146);
and U5753 (N_5753,N_2563,N_1292);
and U5754 (N_5754,N_1828,N_2494);
and U5755 (N_5755,N_1798,N_180);
nor U5756 (N_5756,N_41,N_263);
nand U5757 (N_5757,N_1928,N_1880);
nand U5758 (N_5758,N_1659,N_2054);
nor U5759 (N_5759,N_3069,N_201);
nor U5760 (N_5760,N_1116,N_2378);
and U5761 (N_5761,N_2662,N_647);
or U5762 (N_5762,N_1744,N_2290);
and U5763 (N_5763,N_2812,N_626);
xor U5764 (N_5764,N_2152,N_2802);
or U5765 (N_5765,N_1082,N_2212);
and U5766 (N_5766,N_3080,N_1295);
and U5767 (N_5767,N_405,N_421);
xnor U5768 (N_5768,N_812,N_2660);
and U5769 (N_5769,N_1385,N_1866);
or U5770 (N_5770,N_1911,N_3040);
nor U5771 (N_5771,N_233,N_2644);
nand U5772 (N_5772,N_301,N_534);
nor U5773 (N_5773,N_2044,N_2423);
and U5774 (N_5774,N_2268,N_2746);
and U5775 (N_5775,N_3079,N_1963);
nor U5776 (N_5776,N_2975,N_1163);
xnor U5777 (N_5777,N_412,N_231);
nor U5778 (N_5778,N_2193,N_2885);
and U5779 (N_5779,N_607,N_2001);
or U5780 (N_5780,N_1121,N_763);
and U5781 (N_5781,N_2046,N_310);
nand U5782 (N_5782,N_428,N_855);
nand U5783 (N_5783,N_1973,N_1377);
nor U5784 (N_5784,N_1619,N_130);
or U5785 (N_5785,N_651,N_2269);
or U5786 (N_5786,N_1229,N_26);
or U5787 (N_5787,N_285,N_1094);
and U5788 (N_5788,N_2631,N_432);
xor U5789 (N_5789,N_1691,N_3042);
and U5790 (N_5790,N_1182,N_1897);
nand U5791 (N_5791,N_3018,N_2798);
or U5792 (N_5792,N_204,N_51);
and U5793 (N_5793,N_2740,N_1829);
nor U5794 (N_5794,N_770,N_1286);
nor U5795 (N_5795,N_1269,N_1042);
nand U5796 (N_5796,N_2285,N_1500);
or U5797 (N_5797,N_2621,N_2007);
or U5798 (N_5798,N_742,N_3101);
or U5799 (N_5799,N_1420,N_2089);
xor U5800 (N_5800,N_2197,N_1239);
xor U5801 (N_5801,N_1977,N_3058);
nor U5802 (N_5802,N_2952,N_603);
nor U5803 (N_5803,N_296,N_682);
and U5804 (N_5804,N_618,N_1186);
or U5805 (N_5805,N_464,N_1471);
xnor U5806 (N_5806,N_2276,N_1157);
or U5807 (N_5807,N_647,N_709);
or U5808 (N_5808,N_2799,N_656);
xnor U5809 (N_5809,N_699,N_2885);
or U5810 (N_5810,N_406,N_1834);
and U5811 (N_5811,N_2420,N_1832);
nor U5812 (N_5812,N_1980,N_1637);
or U5813 (N_5813,N_2038,N_164);
nand U5814 (N_5814,N_1985,N_268);
or U5815 (N_5815,N_2899,N_2342);
nand U5816 (N_5816,N_695,N_2456);
or U5817 (N_5817,N_2497,N_1);
and U5818 (N_5818,N_718,N_1880);
nand U5819 (N_5819,N_198,N_2409);
and U5820 (N_5820,N_657,N_2281);
and U5821 (N_5821,N_2321,N_475);
and U5822 (N_5822,N_1871,N_731);
and U5823 (N_5823,N_1150,N_394);
xor U5824 (N_5824,N_2222,N_2591);
nand U5825 (N_5825,N_727,N_2531);
or U5826 (N_5826,N_775,N_1727);
nand U5827 (N_5827,N_827,N_1180);
or U5828 (N_5828,N_2357,N_270);
nand U5829 (N_5829,N_1650,N_2150);
nand U5830 (N_5830,N_1349,N_1353);
nor U5831 (N_5831,N_1367,N_2825);
nand U5832 (N_5832,N_2973,N_1445);
xnor U5833 (N_5833,N_1033,N_1541);
nor U5834 (N_5834,N_2472,N_1739);
and U5835 (N_5835,N_736,N_653);
nor U5836 (N_5836,N_2926,N_1961);
xnor U5837 (N_5837,N_51,N_123);
or U5838 (N_5838,N_232,N_3104);
nor U5839 (N_5839,N_1345,N_49);
xor U5840 (N_5840,N_829,N_635);
or U5841 (N_5841,N_2399,N_974);
nor U5842 (N_5842,N_543,N_839);
and U5843 (N_5843,N_122,N_1172);
and U5844 (N_5844,N_1554,N_1291);
or U5845 (N_5845,N_1506,N_2112);
nand U5846 (N_5846,N_3086,N_3013);
or U5847 (N_5847,N_1235,N_2398);
and U5848 (N_5848,N_1616,N_991);
or U5849 (N_5849,N_57,N_1623);
or U5850 (N_5850,N_676,N_2262);
nand U5851 (N_5851,N_526,N_108);
nor U5852 (N_5852,N_1476,N_1093);
nand U5853 (N_5853,N_88,N_2727);
nand U5854 (N_5854,N_107,N_517);
or U5855 (N_5855,N_2530,N_2957);
and U5856 (N_5856,N_2439,N_336);
nand U5857 (N_5857,N_309,N_436);
or U5858 (N_5858,N_216,N_2641);
nor U5859 (N_5859,N_1471,N_2414);
and U5860 (N_5860,N_2296,N_2998);
or U5861 (N_5861,N_2926,N_2645);
nand U5862 (N_5862,N_799,N_1090);
or U5863 (N_5863,N_1997,N_828);
nor U5864 (N_5864,N_2604,N_1293);
nor U5865 (N_5865,N_2171,N_1056);
or U5866 (N_5866,N_1826,N_1758);
nand U5867 (N_5867,N_2058,N_3064);
or U5868 (N_5868,N_2658,N_1981);
xor U5869 (N_5869,N_316,N_1913);
xor U5870 (N_5870,N_596,N_1722);
nand U5871 (N_5871,N_2106,N_987);
nor U5872 (N_5872,N_2439,N_1693);
and U5873 (N_5873,N_1120,N_2339);
and U5874 (N_5874,N_1674,N_1141);
or U5875 (N_5875,N_666,N_1252);
nor U5876 (N_5876,N_2220,N_2505);
xnor U5877 (N_5877,N_1011,N_829);
nor U5878 (N_5878,N_2561,N_2856);
nor U5879 (N_5879,N_45,N_615);
and U5880 (N_5880,N_2556,N_892);
and U5881 (N_5881,N_631,N_913);
or U5882 (N_5882,N_709,N_2287);
or U5883 (N_5883,N_930,N_286);
nor U5884 (N_5884,N_1934,N_3006);
nand U5885 (N_5885,N_2601,N_1945);
xnor U5886 (N_5886,N_291,N_2903);
nand U5887 (N_5887,N_2410,N_2430);
nor U5888 (N_5888,N_1761,N_2543);
and U5889 (N_5889,N_1076,N_1147);
nor U5890 (N_5890,N_200,N_844);
nand U5891 (N_5891,N_2617,N_2178);
or U5892 (N_5892,N_1295,N_1895);
nand U5893 (N_5893,N_542,N_1436);
and U5894 (N_5894,N_3045,N_2237);
or U5895 (N_5895,N_18,N_758);
xnor U5896 (N_5896,N_1630,N_2793);
and U5897 (N_5897,N_2040,N_1576);
or U5898 (N_5898,N_1,N_1216);
and U5899 (N_5899,N_2219,N_390);
nand U5900 (N_5900,N_591,N_667);
and U5901 (N_5901,N_1713,N_652);
nor U5902 (N_5902,N_2823,N_2397);
nor U5903 (N_5903,N_3022,N_2474);
and U5904 (N_5904,N_1016,N_1432);
or U5905 (N_5905,N_2145,N_1209);
nor U5906 (N_5906,N_1710,N_2913);
nor U5907 (N_5907,N_2088,N_1509);
or U5908 (N_5908,N_86,N_352);
or U5909 (N_5909,N_2680,N_2090);
or U5910 (N_5910,N_2447,N_447);
and U5911 (N_5911,N_542,N_87);
nand U5912 (N_5912,N_1648,N_785);
nor U5913 (N_5913,N_2348,N_2120);
or U5914 (N_5914,N_871,N_2774);
and U5915 (N_5915,N_31,N_642);
or U5916 (N_5916,N_371,N_2922);
nor U5917 (N_5917,N_3079,N_2878);
xor U5918 (N_5918,N_260,N_1130);
or U5919 (N_5919,N_199,N_1954);
and U5920 (N_5920,N_2201,N_22);
nand U5921 (N_5921,N_1182,N_887);
and U5922 (N_5922,N_2947,N_1842);
or U5923 (N_5923,N_1542,N_933);
nor U5924 (N_5924,N_2042,N_138);
nor U5925 (N_5925,N_168,N_1092);
nor U5926 (N_5926,N_1366,N_2666);
nand U5927 (N_5927,N_1413,N_1326);
nor U5928 (N_5928,N_1546,N_2776);
or U5929 (N_5929,N_1133,N_1654);
xnor U5930 (N_5930,N_916,N_1090);
and U5931 (N_5931,N_2799,N_2208);
or U5932 (N_5932,N_1080,N_1829);
nor U5933 (N_5933,N_1634,N_127);
nand U5934 (N_5934,N_894,N_50);
or U5935 (N_5935,N_1769,N_843);
and U5936 (N_5936,N_257,N_1696);
and U5937 (N_5937,N_3121,N_152);
and U5938 (N_5938,N_860,N_239);
nand U5939 (N_5939,N_1285,N_279);
nand U5940 (N_5940,N_1919,N_2545);
nor U5941 (N_5941,N_2579,N_2732);
nor U5942 (N_5942,N_705,N_868);
nor U5943 (N_5943,N_2425,N_426);
and U5944 (N_5944,N_2605,N_1678);
or U5945 (N_5945,N_1052,N_2747);
or U5946 (N_5946,N_1304,N_2329);
nand U5947 (N_5947,N_365,N_1701);
and U5948 (N_5948,N_2174,N_2392);
or U5949 (N_5949,N_1971,N_1930);
and U5950 (N_5950,N_641,N_946);
and U5951 (N_5951,N_1431,N_2941);
or U5952 (N_5952,N_1204,N_1239);
nor U5953 (N_5953,N_2058,N_387);
nor U5954 (N_5954,N_1525,N_394);
and U5955 (N_5955,N_1875,N_1077);
or U5956 (N_5956,N_1186,N_2327);
or U5957 (N_5957,N_2367,N_2735);
nor U5958 (N_5958,N_747,N_959);
nand U5959 (N_5959,N_173,N_798);
xnor U5960 (N_5960,N_1260,N_844);
nand U5961 (N_5961,N_2225,N_1533);
nor U5962 (N_5962,N_1423,N_1368);
xnor U5963 (N_5963,N_2529,N_772);
nor U5964 (N_5964,N_3019,N_1470);
nand U5965 (N_5965,N_491,N_1313);
nor U5966 (N_5966,N_138,N_2986);
nand U5967 (N_5967,N_1276,N_566);
or U5968 (N_5968,N_275,N_3044);
and U5969 (N_5969,N_1958,N_980);
and U5970 (N_5970,N_702,N_575);
nor U5971 (N_5971,N_1031,N_2393);
and U5972 (N_5972,N_520,N_2593);
xnor U5973 (N_5973,N_2221,N_499);
and U5974 (N_5974,N_1223,N_3118);
xnor U5975 (N_5975,N_1404,N_1795);
or U5976 (N_5976,N_652,N_66);
xor U5977 (N_5977,N_277,N_2857);
nand U5978 (N_5978,N_1560,N_646);
and U5979 (N_5979,N_786,N_2035);
xnor U5980 (N_5980,N_380,N_1119);
or U5981 (N_5981,N_230,N_1343);
nand U5982 (N_5982,N_1820,N_1344);
xor U5983 (N_5983,N_317,N_1629);
nor U5984 (N_5984,N_1578,N_2308);
or U5985 (N_5985,N_2192,N_2493);
nor U5986 (N_5986,N_2163,N_1569);
and U5987 (N_5987,N_2700,N_63);
nor U5988 (N_5988,N_570,N_2282);
or U5989 (N_5989,N_741,N_1574);
xnor U5990 (N_5990,N_599,N_278);
and U5991 (N_5991,N_2100,N_1236);
xnor U5992 (N_5992,N_617,N_1294);
xor U5993 (N_5993,N_1598,N_1773);
or U5994 (N_5994,N_1195,N_1803);
nor U5995 (N_5995,N_1537,N_2635);
and U5996 (N_5996,N_1049,N_509);
or U5997 (N_5997,N_428,N_2635);
nand U5998 (N_5998,N_1219,N_958);
or U5999 (N_5999,N_264,N_1247);
nor U6000 (N_6000,N_2036,N_931);
xnor U6001 (N_6001,N_1780,N_1117);
nor U6002 (N_6002,N_2553,N_661);
nand U6003 (N_6003,N_2037,N_58);
nor U6004 (N_6004,N_2886,N_696);
nor U6005 (N_6005,N_3098,N_1545);
and U6006 (N_6006,N_669,N_2107);
nor U6007 (N_6007,N_553,N_2092);
or U6008 (N_6008,N_913,N_1123);
nor U6009 (N_6009,N_3094,N_1503);
nor U6010 (N_6010,N_1896,N_194);
nand U6011 (N_6011,N_3033,N_1313);
nand U6012 (N_6012,N_812,N_1295);
nor U6013 (N_6013,N_2603,N_2224);
or U6014 (N_6014,N_1687,N_2377);
nand U6015 (N_6015,N_3087,N_978);
or U6016 (N_6016,N_1100,N_392);
nand U6017 (N_6017,N_545,N_1877);
nor U6018 (N_6018,N_2229,N_2745);
nand U6019 (N_6019,N_2345,N_417);
or U6020 (N_6020,N_879,N_176);
xor U6021 (N_6021,N_1184,N_763);
xnor U6022 (N_6022,N_22,N_1151);
nand U6023 (N_6023,N_2839,N_663);
nor U6024 (N_6024,N_1934,N_2931);
nor U6025 (N_6025,N_688,N_2855);
nand U6026 (N_6026,N_2078,N_1344);
nand U6027 (N_6027,N_429,N_812);
nor U6028 (N_6028,N_865,N_1369);
nand U6029 (N_6029,N_1379,N_3004);
nor U6030 (N_6030,N_2858,N_619);
nor U6031 (N_6031,N_2069,N_863);
or U6032 (N_6032,N_2628,N_2277);
or U6033 (N_6033,N_629,N_775);
nand U6034 (N_6034,N_2936,N_2242);
xor U6035 (N_6035,N_1527,N_1931);
nand U6036 (N_6036,N_590,N_1053);
xor U6037 (N_6037,N_913,N_488);
or U6038 (N_6038,N_529,N_2913);
nand U6039 (N_6039,N_216,N_451);
and U6040 (N_6040,N_52,N_2383);
xor U6041 (N_6041,N_1234,N_1757);
and U6042 (N_6042,N_1209,N_1337);
and U6043 (N_6043,N_1244,N_1222);
xnor U6044 (N_6044,N_2621,N_2057);
or U6045 (N_6045,N_2186,N_2574);
nor U6046 (N_6046,N_1953,N_1720);
or U6047 (N_6047,N_2318,N_397);
nor U6048 (N_6048,N_973,N_743);
nor U6049 (N_6049,N_474,N_2405);
nand U6050 (N_6050,N_747,N_275);
nor U6051 (N_6051,N_2185,N_2588);
nand U6052 (N_6052,N_2944,N_1522);
nor U6053 (N_6053,N_2404,N_2481);
and U6054 (N_6054,N_548,N_282);
xnor U6055 (N_6055,N_1708,N_2366);
and U6056 (N_6056,N_70,N_45);
or U6057 (N_6057,N_694,N_1188);
or U6058 (N_6058,N_1778,N_2289);
and U6059 (N_6059,N_1621,N_3121);
and U6060 (N_6060,N_1101,N_1404);
and U6061 (N_6061,N_449,N_229);
nand U6062 (N_6062,N_0,N_2865);
nor U6063 (N_6063,N_2193,N_196);
xnor U6064 (N_6064,N_395,N_1300);
and U6065 (N_6065,N_1109,N_260);
xor U6066 (N_6066,N_1622,N_1399);
and U6067 (N_6067,N_1809,N_964);
or U6068 (N_6068,N_1278,N_3000);
xnor U6069 (N_6069,N_2570,N_515);
nand U6070 (N_6070,N_1231,N_1723);
or U6071 (N_6071,N_1858,N_2632);
nand U6072 (N_6072,N_1612,N_2390);
nor U6073 (N_6073,N_1427,N_1980);
or U6074 (N_6074,N_3088,N_1317);
nand U6075 (N_6075,N_2221,N_353);
and U6076 (N_6076,N_2706,N_319);
nor U6077 (N_6077,N_615,N_1895);
nand U6078 (N_6078,N_1829,N_2729);
or U6079 (N_6079,N_2665,N_2570);
and U6080 (N_6080,N_2082,N_1905);
nand U6081 (N_6081,N_2225,N_661);
nand U6082 (N_6082,N_640,N_1480);
nand U6083 (N_6083,N_2276,N_632);
and U6084 (N_6084,N_2441,N_1591);
and U6085 (N_6085,N_2019,N_2500);
and U6086 (N_6086,N_164,N_2016);
or U6087 (N_6087,N_1200,N_1211);
or U6088 (N_6088,N_1896,N_2678);
nand U6089 (N_6089,N_1357,N_534);
nand U6090 (N_6090,N_1376,N_1775);
and U6091 (N_6091,N_2943,N_56);
or U6092 (N_6092,N_308,N_1230);
or U6093 (N_6093,N_285,N_126);
and U6094 (N_6094,N_2078,N_646);
or U6095 (N_6095,N_2942,N_329);
and U6096 (N_6096,N_1623,N_14);
nand U6097 (N_6097,N_2199,N_3014);
nand U6098 (N_6098,N_2031,N_1763);
xnor U6099 (N_6099,N_1337,N_331);
nor U6100 (N_6100,N_763,N_208);
or U6101 (N_6101,N_791,N_1686);
or U6102 (N_6102,N_1198,N_234);
or U6103 (N_6103,N_1074,N_17);
nand U6104 (N_6104,N_1632,N_2762);
or U6105 (N_6105,N_1300,N_1266);
nor U6106 (N_6106,N_3029,N_2238);
nor U6107 (N_6107,N_1794,N_2986);
xnor U6108 (N_6108,N_976,N_2487);
or U6109 (N_6109,N_2599,N_2671);
nor U6110 (N_6110,N_1428,N_1949);
or U6111 (N_6111,N_2687,N_7);
and U6112 (N_6112,N_2079,N_992);
nor U6113 (N_6113,N_308,N_1549);
xnor U6114 (N_6114,N_380,N_3119);
nand U6115 (N_6115,N_19,N_172);
and U6116 (N_6116,N_2893,N_1883);
or U6117 (N_6117,N_694,N_11);
or U6118 (N_6118,N_2065,N_1030);
and U6119 (N_6119,N_2277,N_2040);
nand U6120 (N_6120,N_2397,N_3036);
and U6121 (N_6121,N_239,N_666);
and U6122 (N_6122,N_876,N_1151);
or U6123 (N_6123,N_803,N_1860);
nand U6124 (N_6124,N_24,N_1749);
or U6125 (N_6125,N_1688,N_2687);
and U6126 (N_6126,N_125,N_117);
nand U6127 (N_6127,N_1564,N_1030);
nand U6128 (N_6128,N_1326,N_2747);
and U6129 (N_6129,N_2304,N_2612);
nand U6130 (N_6130,N_2574,N_546);
or U6131 (N_6131,N_1596,N_2158);
nor U6132 (N_6132,N_1689,N_685);
nand U6133 (N_6133,N_245,N_2412);
and U6134 (N_6134,N_3077,N_1640);
nor U6135 (N_6135,N_1747,N_1218);
xnor U6136 (N_6136,N_2424,N_1846);
and U6137 (N_6137,N_2204,N_90);
nand U6138 (N_6138,N_326,N_2778);
or U6139 (N_6139,N_854,N_3080);
or U6140 (N_6140,N_1750,N_2618);
and U6141 (N_6141,N_452,N_417);
nand U6142 (N_6142,N_1386,N_794);
nor U6143 (N_6143,N_600,N_2675);
nor U6144 (N_6144,N_1467,N_705);
and U6145 (N_6145,N_1653,N_2541);
and U6146 (N_6146,N_1976,N_760);
xor U6147 (N_6147,N_1780,N_1081);
nor U6148 (N_6148,N_2586,N_373);
nor U6149 (N_6149,N_2630,N_2191);
nor U6150 (N_6150,N_335,N_1489);
or U6151 (N_6151,N_384,N_1858);
xor U6152 (N_6152,N_2279,N_2737);
nand U6153 (N_6153,N_111,N_2305);
nor U6154 (N_6154,N_618,N_2808);
nor U6155 (N_6155,N_53,N_1862);
xnor U6156 (N_6156,N_974,N_99);
and U6157 (N_6157,N_869,N_2595);
nand U6158 (N_6158,N_2626,N_906);
or U6159 (N_6159,N_1831,N_390);
nor U6160 (N_6160,N_1419,N_636);
or U6161 (N_6161,N_2758,N_1041);
and U6162 (N_6162,N_1760,N_174);
or U6163 (N_6163,N_190,N_80);
and U6164 (N_6164,N_1075,N_489);
nor U6165 (N_6165,N_1583,N_460);
nor U6166 (N_6166,N_2380,N_1359);
nand U6167 (N_6167,N_1943,N_1716);
nor U6168 (N_6168,N_731,N_2783);
and U6169 (N_6169,N_383,N_2965);
nand U6170 (N_6170,N_2307,N_1394);
xnor U6171 (N_6171,N_1198,N_2602);
and U6172 (N_6172,N_914,N_36);
nor U6173 (N_6173,N_1271,N_341);
nor U6174 (N_6174,N_2161,N_1690);
nor U6175 (N_6175,N_2124,N_1293);
nand U6176 (N_6176,N_1010,N_2302);
and U6177 (N_6177,N_1509,N_2580);
and U6178 (N_6178,N_401,N_424);
or U6179 (N_6179,N_1316,N_2946);
xor U6180 (N_6180,N_3032,N_2746);
or U6181 (N_6181,N_1807,N_2710);
xor U6182 (N_6182,N_1683,N_1936);
or U6183 (N_6183,N_2055,N_2469);
or U6184 (N_6184,N_1413,N_2481);
and U6185 (N_6185,N_2563,N_888);
xnor U6186 (N_6186,N_1045,N_276);
or U6187 (N_6187,N_3034,N_400);
and U6188 (N_6188,N_1394,N_2862);
or U6189 (N_6189,N_1643,N_923);
nor U6190 (N_6190,N_2757,N_957);
or U6191 (N_6191,N_1650,N_2048);
nand U6192 (N_6192,N_1078,N_2078);
nor U6193 (N_6193,N_1746,N_1355);
and U6194 (N_6194,N_2240,N_597);
and U6195 (N_6195,N_1687,N_834);
and U6196 (N_6196,N_36,N_1172);
or U6197 (N_6197,N_547,N_1200);
nor U6198 (N_6198,N_2726,N_739);
nand U6199 (N_6199,N_1779,N_457);
nor U6200 (N_6200,N_1077,N_2023);
or U6201 (N_6201,N_1317,N_1176);
nand U6202 (N_6202,N_731,N_789);
nor U6203 (N_6203,N_2669,N_764);
nand U6204 (N_6204,N_2959,N_379);
nand U6205 (N_6205,N_1769,N_2044);
nor U6206 (N_6206,N_759,N_932);
nand U6207 (N_6207,N_421,N_95);
or U6208 (N_6208,N_456,N_2007);
nor U6209 (N_6209,N_2341,N_1193);
or U6210 (N_6210,N_322,N_671);
and U6211 (N_6211,N_907,N_2633);
nor U6212 (N_6212,N_1381,N_2907);
and U6213 (N_6213,N_244,N_3043);
and U6214 (N_6214,N_372,N_2093);
nor U6215 (N_6215,N_1004,N_3116);
nor U6216 (N_6216,N_2382,N_978);
nor U6217 (N_6217,N_125,N_1015);
or U6218 (N_6218,N_2816,N_663);
xor U6219 (N_6219,N_2200,N_1634);
xnor U6220 (N_6220,N_1142,N_1262);
nand U6221 (N_6221,N_612,N_112);
or U6222 (N_6222,N_218,N_147);
nand U6223 (N_6223,N_2274,N_981);
and U6224 (N_6224,N_522,N_440);
and U6225 (N_6225,N_1908,N_2911);
nor U6226 (N_6226,N_1233,N_834);
and U6227 (N_6227,N_2178,N_97);
and U6228 (N_6228,N_2688,N_59);
or U6229 (N_6229,N_1255,N_3075);
xor U6230 (N_6230,N_1275,N_3045);
nand U6231 (N_6231,N_2159,N_2221);
and U6232 (N_6232,N_1066,N_76);
or U6233 (N_6233,N_1227,N_1624);
and U6234 (N_6234,N_2476,N_496);
and U6235 (N_6235,N_550,N_507);
and U6236 (N_6236,N_1261,N_397);
nor U6237 (N_6237,N_746,N_3021);
and U6238 (N_6238,N_2659,N_1177);
or U6239 (N_6239,N_1094,N_2323);
and U6240 (N_6240,N_686,N_1848);
nand U6241 (N_6241,N_2697,N_1526);
nor U6242 (N_6242,N_467,N_840);
or U6243 (N_6243,N_3087,N_2345);
or U6244 (N_6244,N_566,N_414);
and U6245 (N_6245,N_2458,N_2965);
and U6246 (N_6246,N_23,N_2170);
or U6247 (N_6247,N_998,N_3032);
or U6248 (N_6248,N_20,N_2463);
or U6249 (N_6249,N_1467,N_1122);
or U6250 (N_6250,N_3858,N_4017);
nand U6251 (N_6251,N_4787,N_6175);
and U6252 (N_6252,N_3566,N_3549);
nand U6253 (N_6253,N_4746,N_3291);
nor U6254 (N_6254,N_3957,N_6171);
or U6255 (N_6255,N_4918,N_6001);
nor U6256 (N_6256,N_5492,N_5097);
or U6257 (N_6257,N_3875,N_4485);
nor U6258 (N_6258,N_3892,N_3832);
nor U6259 (N_6259,N_5174,N_3516);
and U6260 (N_6260,N_3197,N_6204);
and U6261 (N_6261,N_4188,N_4340);
nand U6262 (N_6262,N_4734,N_3647);
xnor U6263 (N_6263,N_4264,N_3756);
xnor U6264 (N_6264,N_5814,N_3916);
nand U6265 (N_6265,N_4430,N_5919);
nor U6266 (N_6266,N_5441,N_4421);
and U6267 (N_6267,N_4969,N_3603);
nand U6268 (N_6268,N_3234,N_6231);
and U6269 (N_6269,N_3191,N_5094);
nand U6270 (N_6270,N_4982,N_4711);
xor U6271 (N_6271,N_6015,N_3551);
nand U6272 (N_6272,N_5754,N_3691);
nor U6273 (N_6273,N_5082,N_6058);
nand U6274 (N_6274,N_5678,N_3966);
nor U6275 (N_6275,N_4375,N_4577);
nor U6276 (N_6276,N_4939,N_3894);
xor U6277 (N_6277,N_5209,N_6153);
nor U6278 (N_6278,N_4554,N_5440);
nand U6279 (N_6279,N_4214,N_5085);
and U6280 (N_6280,N_4462,N_4432);
xnor U6281 (N_6281,N_5250,N_5914);
or U6282 (N_6282,N_4830,N_5732);
and U6283 (N_6283,N_3173,N_3141);
nor U6284 (N_6284,N_4946,N_3668);
and U6285 (N_6285,N_3153,N_3186);
nand U6286 (N_6286,N_4652,N_5080);
nand U6287 (N_6287,N_5634,N_4322);
or U6288 (N_6288,N_5220,N_4185);
and U6289 (N_6289,N_5452,N_3459);
nor U6290 (N_6290,N_5302,N_5834);
nor U6291 (N_6291,N_3819,N_6206);
nand U6292 (N_6292,N_5066,N_6156);
and U6293 (N_6293,N_3359,N_3783);
xnor U6294 (N_6294,N_4367,N_3730);
and U6295 (N_6295,N_5433,N_4046);
or U6296 (N_6296,N_5670,N_4549);
and U6297 (N_6297,N_3537,N_5093);
nand U6298 (N_6298,N_3754,N_5352);
nand U6299 (N_6299,N_4678,N_4945);
nand U6300 (N_6300,N_5524,N_4953);
and U6301 (N_6301,N_6236,N_5659);
nand U6302 (N_6302,N_3990,N_4476);
xor U6303 (N_6303,N_3198,N_6004);
nor U6304 (N_6304,N_4143,N_3740);
nand U6305 (N_6305,N_6076,N_4843);
nor U6306 (N_6306,N_3231,N_5824);
nand U6307 (N_6307,N_5833,N_5614);
nand U6308 (N_6308,N_5377,N_4628);
nand U6309 (N_6309,N_5325,N_5182);
xor U6310 (N_6310,N_3321,N_4045);
nor U6311 (N_6311,N_3736,N_4473);
nand U6312 (N_6312,N_3811,N_6192);
and U6313 (N_6313,N_5599,N_3673);
nor U6314 (N_6314,N_4030,N_3339);
or U6315 (N_6315,N_3642,N_6129);
or U6316 (N_6316,N_3637,N_4675);
nor U6317 (N_6317,N_3918,N_3974);
and U6318 (N_6318,N_4160,N_4908);
nor U6319 (N_6319,N_6123,N_4065);
nand U6320 (N_6320,N_4450,N_5455);
and U6321 (N_6321,N_3996,N_5024);
and U6322 (N_6322,N_4730,N_5436);
nand U6323 (N_6323,N_4791,N_5195);
or U6324 (N_6324,N_4378,N_3177);
and U6325 (N_6325,N_3865,N_4437);
or U6326 (N_6326,N_5029,N_3620);
or U6327 (N_6327,N_4433,N_4486);
or U6328 (N_6328,N_5846,N_5286);
and U6329 (N_6329,N_3480,N_5898);
xnor U6330 (N_6330,N_5362,N_5451);
or U6331 (N_6331,N_5616,N_4545);
xor U6332 (N_6332,N_5493,N_3347);
nor U6333 (N_6333,N_3542,N_6132);
nor U6334 (N_6334,N_5422,N_6089);
nor U6335 (N_6335,N_3268,N_5578);
nor U6336 (N_6336,N_3135,N_3728);
or U6337 (N_6337,N_4026,N_6131);
or U6338 (N_6338,N_3479,N_5995);
nor U6339 (N_6339,N_5326,N_4312);
nor U6340 (N_6340,N_6071,N_5811);
and U6341 (N_6341,N_5867,N_4125);
or U6342 (N_6342,N_4807,N_4496);
nor U6343 (N_6343,N_4077,N_6065);
and U6344 (N_6344,N_3567,N_5718);
or U6345 (N_6345,N_4698,N_3130);
nor U6346 (N_6346,N_4327,N_4548);
and U6347 (N_6347,N_3306,N_5546);
or U6348 (N_6348,N_4275,N_4977);
nand U6349 (N_6349,N_3494,N_4058);
or U6350 (N_6350,N_3632,N_4894);
nor U6351 (N_6351,N_3560,N_4820);
nor U6352 (N_6352,N_5936,N_5943);
or U6353 (N_6353,N_5582,N_3538);
and U6354 (N_6354,N_5866,N_3223);
nor U6355 (N_6355,N_4664,N_3677);
and U6356 (N_6356,N_3140,N_5620);
and U6357 (N_6357,N_5666,N_3945);
or U6358 (N_6358,N_4472,N_6144);
and U6359 (N_6359,N_4836,N_4303);
xnor U6360 (N_6360,N_4138,N_3482);
nor U6361 (N_6361,N_4226,N_5430);
or U6362 (N_6362,N_3839,N_4411);
nand U6363 (N_6363,N_4363,N_5380);
xnor U6364 (N_6364,N_3769,N_4742);
or U6365 (N_6365,N_4020,N_3350);
nor U6366 (N_6366,N_5393,N_5004);
nor U6367 (N_6367,N_6000,N_4636);
nand U6368 (N_6368,N_4137,N_4225);
or U6369 (N_6369,N_6224,N_3382);
nand U6370 (N_6370,N_5177,N_5548);
xnor U6371 (N_6371,N_5632,N_5555);
or U6372 (N_6372,N_5505,N_3574);
nor U6373 (N_6373,N_3834,N_3715);
nand U6374 (N_6374,N_3233,N_5015);
and U6375 (N_6375,N_3300,N_5984);
or U6376 (N_6376,N_5502,N_3443);
or U6377 (N_6377,N_5761,N_5396);
xnor U6378 (N_6378,N_3526,N_3963);
and U6379 (N_6379,N_5775,N_3596);
or U6380 (N_6380,N_5646,N_4521);
nand U6381 (N_6381,N_3388,N_3911);
nor U6382 (N_6382,N_3167,N_4876);
nor U6383 (N_6383,N_5682,N_3931);
or U6384 (N_6384,N_3638,N_4703);
nor U6385 (N_6385,N_3726,N_5645);
xnor U6386 (N_6386,N_5294,N_4447);
or U6387 (N_6387,N_3979,N_6111);
and U6388 (N_6388,N_5776,N_5355);
or U6389 (N_6389,N_4285,N_4621);
xnor U6390 (N_6390,N_6069,N_4000);
and U6391 (N_6391,N_5349,N_5590);
xor U6392 (N_6392,N_3266,N_4453);
and U6393 (N_6393,N_4705,N_3625);
xnor U6394 (N_6394,N_3744,N_3838);
and U6395 (N_6395,N_3840,N_5746);
or U6396 (N_6396,N_6041,N_5092);
and U6397 (N_6397,N_3271,N_5573);
nor U6398 (N_6398,N_5346,N_4480);
and U6399 (N_6399,N_5792,N_4282);
and U6400 (N_6400,N_3132,N_4248);
and U6401 (N_6401,N_4317,N_3855);
nor U6402 (N_6402,N_4262,N_3545);
nor U6403 (N_6403,N_4989,N_4382);
and U6404 (N_6404,N_5234,N_6057);
xnor U6405 (N_6405,N_4362,N_4934);
nand U6406 (N_6406,N_5348,N_3413);
nand U6407 (N_6407,N_4503,N_3485);
nand U6408 (N_6408,N_3866,N_5263);
or U6409 (N_6409,N_5685,N_5511);
and U6410 (N_6410,N_5575,N_5183);
and U6411 (N_6411,N_4872,N_4235);
nand U6412 (N_6412,N_3503,N_4003);
and U6413 (N_6413,N_5901,N_5588);
or U6414 (N_6414,N_4829,N_6221);
or U6415 (N_6415,N_3774,N_5817);
and U6416 (N_6416,N_4760,N_5394);
and U6417 (N_6417,N_6178,N_4154);
and U6418 (N_6418,N_5877,N_5860);
or U6419 (N_6419,N_5164,N_4469);
nand U6420 (N_6420,N_4096,N_3507);
nand U6421 (N_6421,N_5840,N_5930);
and U6422 (N_6422,N_4183,N_3397);
and U6423 (N_6423,N_3706,N_5300);
or U6424 (N_6424,N_5993,N_5468);
and U6425 (N_6425,N_5001,N_4803);
or U6426 (N_6426,N_5579,N_4558);
nand U6427 (N_6427,N_4716,N_3512);
or U6428 (N_6428,N_4580,N_4938);
nand U6429 (N_6429,N_5803,N_6093);
and U6430 (N_6430,N_3904,N_4333);
or U6431 (N_6431,N_3586,N_4550);
nand U6432 (N_6432,N_3786,N_4780);
nand U6433 (N_6433,N_5622,N_4646);
nor U6434 (N_6434,N_3711,N_5828);
xnor U6435 (N_6435,N_4048,N_3420);
nor U6436 (N_6436,N_4018,N_3409);
nand U6437 (N_6437,N_3983,N_5480);
or U6438 (N_6438,N_6003,N_3614);
nor U6439 (N_6439,N_3301,N_5257);
nand U6440 (N_6440,N_6052,N_3719);
or U6441 (N_6441,N_5844,N_3788);
nor U6442 (N_6442,N_4935,N_3320);
nor U6443 (N_6443,N_3442,N_5964);
or U6444 (N_6444,N_3188,N_3852);
nor U6445 (N_6445,N_4229,N_5063);
and U6446 (N_6446,N_5515,N_4933);
nand U6447 (N_6447,N_3572,N_4921);
or U6448 (N_6448,N_5946,N_3475);
nand U6449 (N_6449,N_3750,N_3532);
nor U6450 (N_6450,N_4533,N_4449);
and U6451 (N_6451,N_4852,N_3476);
nand U6452 (N_6452,N_4665,N_4148);
and U6453 (N_6453,N_3228,N_6228);
or U6454 (N_6454,N_6061,N_6039);
or U6455 (N_6455,N_3999,N_5594);
and U6456 (N_6456,N_5727,N_5766);
nand U6457 (N_6457,N_4344,N_6174);
nor U6458 (N_6458,N_6242,N_3854);
and U6459 (N_6459,N_4878,N_4044);
nand U6460 (N_6460,N_3242,N_3376);
nor U6461 (N_6461,N_4247,N_3600);
and U6462 (N_6462,N_3923,N_4713);
nor U6463 (N_6463,N_5163,N_3980);
nand U6464 (N_6464,N_3848,N_3798);
or U6465 (N_6465,N_4055,N_5042);
xor U6466 (N_6466,N_6104,N_4025);
or U6467 (N_6467,N_4896,N_4749);
or U6468 (N_6468,N_5795,N_4528);
and U6469 (N_6469,N_5071,N_3506);
and U6470 (N_6470,N_3988,N_3418);
or U6471 (N_6471,N_4607,N_5216);
or U6472 (N_6472,N_5981,N_5184);
and U6473 (N_6473,N_4592,N_3556);
nor U6474 (N_6474,N_4808,N_4861);
or U6475 (N_6475,N_3617,N_5412);
and U6476 (N_6476,N_4855,N_3787);
nand U6477 (N_6477,N_3995,N_5049);
xor U6478 (N_6478,N_4395,N_4885);
and U6479 (N_6479,N_4756,N_3899);
nand U6480 (N_6480,N_5020,N_6226);
nor U6481 (N_6481,N_4539,N_5595);
and U6482 (N_6482,N_4546,N_4740);
nor U6483 (N_6483,N_3484,N_3498);
nand U6484 (N_6484,N_5288,N_3954);
and U6485 (N_6485,N_5636,N_5457);
nor U6486 (N_6486,N_5601,N_4278);
nand U6487 (N_6487,N_5361,N_3913);
and U6488 (N_6488,N_4518,N_3951);
nor U6489 (N_6489,N_6074,N_4222);
or U6490 (N_6490,N_4391,N_4608);
nor U6491 (N_6491,N_5711,N_5320);
and U6492 (N_6492,N_6238,N_5008);
nand U6493 (N_6493,N_5251,N_3845);
or U6494 (N_6494,N_4374,N_5783);
and U6495 (N_6495,N_4640,N_6008);
or U6496 (N_6496,N_3535,N_4068);
or U6497 (N_6497,N_5664,N_4279);
nand U6498 (N_6498,N_3273,N_4602);
or U6499 (N_6499,N_5641,N_6233);
nand U6500 (N_6500,N_4793,N_4738);
nor U6501 (N_6501,N_6086,N_4634);
and U6502 (N_6502,N_4810,N_5338);
or U6503 (N_6503,N_4244,N_3561);
xor U6504 (N_6504,N_3212,N_4601);
nand U6505 (N_6505,N_4691,N_5970);
or U6506 (N_6506,N_3917,N_4258);
nor U6507 (N_6507,N_5961,N_4108);
nand U6508 (N_6508,N_4383,N_5559);
nand U6509 (N_6509,N_6198,N_3352);
or U6510 (N_6510,N_5083,N_3369);
nor U6511 (N_6511,N_4626,N_5985);
or U6512 (N_6512,N_3138,N_5035);
nor U6513 (N_6513,N_3410,N_4156);
nand U6514 (N_6514,N_6237,N_3696);
and U6515 (N_6515,N_5696,N_5966);
nand U6516 (N_6516,N_4530,N_4984);
nand U6517 (N_6517,N_4338,N_4342);
nor U6518 (N_6518,N_4165,N_5375);
and U6519 (N_6519,N_5003,N_5912);
xnor U6520 (N_6520,N_3569,N_5850);
and U6521 (N_6521,N_5988,N_6208);
nor U6522 (N_6522,N_4202,N_3763);
nand U6523 (N_6523,N_4463,N_4932);
or U6524 (N_6524,N_5038,N_4522);
nor U6525 (N_6525,N_4130,N_5612);
xnor U6526 (N_6526,N_3438,N_3310);
or U6527 (N_6527,N_5267,N_5528);
or U6528 (N_6528,N_4186,N_4647);
nand U6529 (N_6529,N_3679,N_3577);
nor U6530 (N_6530,N_4136,N_5295);
or U6531 (N_6531,N_4668,N_4440);
and U6532 (N_6532,N_3329,N_3692);
and U6533 (N_6533,N_3245,N_4859);
and U6534 (N_6534,N_3488,N_4565);
xor U6535 (N_6535,N_4571,N_3568);
nor U6536 (N_6536,N_5733,N_6092);
and U6537 (N_6537,N_5508,N_5378);
or U6538 (N_6538,N_5483,N_3161);
and U6539 (N_6539,N_3670,N_5141);
xnor U6540 (N_6540,N_3841,N_5117);
or U6541 (N_6541,N_5414,N_6148);
and U6542 (N_6542,N_3346,N_3623);
nor U6543 (N_6543,N_3348,N_5143);
or U6544 (N_6544,N_4388,N_4893);
or U6545 (N_6545,N_5437,N_5005);
nor U6546 (N_6546,N_6220,N_4866);
nor U6547 (N_6547,N_3776,N_5262);
nor U6548 (N_6548,N_3508,N_6072);
or U6549 (N_6549,N_5668,N_5976);
or U6550 (N_6550,N_3519,N_3587);
xnor U6551 (N_6551,N_4397,N_3361);
or U6552 (N_6552,N_3294,N_5968);
and U6553 (N_6553,N_4423,N_5058);
nand U6554 (N_6554,N_4336,N_3604);
nand U6555 (N_6555,N_5109,N_4770);
nor U6556 (N_6556,N_5818,N_5723);
nor U6557 (N_6557,N_5199,N_4039);
xnor U6558 (N_6558,N_5736,N_4999);
nand U6559 (N_6559,N_4805,N_5569);
nor U6560 (N_6560,N_4639,N_4105);
nand U6561 (N_6561,N_5387,N_3969);
and U6562 (N_6562,N_5046,N_5161);
nand U6563 (N_6563,N_4254,N_3912);
nand U6564 (N_6564,N_6169,N_5699);
and U6565 (N_6565,N_6037,N_4837);
and U6566 (N_6566,N_3779,N_6029);
and U6567 (N_6567,N_3707,N_6140);
and U6568 (N_6568,N_5535,N_5989);
or U6569 (N_6569,N_4699,N_4922);
nor U6570 (N_6570,N_3653,N_3939);
nor U6571 (N_6571,N_3505,N_5610);
nor U6572 (N_6572,N_3399,N_3164);
xnor U6573 (N_6573,N_4813,N_4723);
or U6574 (N_6574,N_3869,N_5841);
or U6575 (N_6575,N_4735,N_3635);
and U6576 (N_6576,N_5655,N_5978);
xnor U6577 (N_6577,N_4458,N_5434);
xnor U6578 (N_6578,N_4882,N_3741);
nor U6579 (N_6579,N_3725,N_5805);
and U6580 (N_6580,N_5246,N_4884);
and U6581 (N_6581,N_3861,N_3548);
and U6582 (N_6582,N_3651,N_3759);
nand U6583 (N_6583,N_3536,N_4833);
and U6584 (N_6584,N_5116,N_5929);
or U6585 (N_6585,N_5808,N_3664);
and U6586 (N_6586,N_4274,N_5934);
nor U6587 (N_6587,N_3955,N_5206);
and U6588 (N_6588,N_4063,N_3172);
nand U6589 (N_6589,N_3222,N_6120);
nor U6590 (N_6590,N_5619,N_3193);
nand U6591 (N_6591,N_5821,N_6067);
xor U6592 (N_6592,N_3477,N_3169);
xnor U6593 (N_6593,N_5025,N_4660);
and U6594 (N_6594,N_5462,N_5498);
nand U6595 (N_6595,N_6079,N_5779);
nand U6596 (N_6596,N_4455,N_5780);
and U6597 (N_6597,N_4109,N_4271);
or U6598 (N_6598,N_3766,N_3814);
or U6599 (N_6599,N_3981,N_5615);
nor U6600 (N_6600,N_5863,N_6043);
xor U6601 (N_6601,N_3760,N_3495);
nand U6602 (N_6602,N_4179,N_4663);
nor U6603 (N_6603,N_4253,N_6017);
nand U6604 (N_6604,N_5185,N_5425);
or U6605 (N_6605,N_5992,N_4215);
nor U6606 (N_6606,N_5996,N_5088);
nor U6607 (N_6607,N_5370,N_4578);
and U6608 (N_6608,N_4356,N_4069);
nand U6609 (N_6609,N_5747,N_4841);
and U6610 (N_6610,N_5854,N_4643);
nor U6611 (N_6611,N_4406,N_4627);
nand U6612 (N_6612,N_3335,N_3504);
nand U6613 (N_6613,N_4822,N_4702);
or U6614 (N_6614,N_5120,N_5525);
nand U6615 (N_6615,N_4587,N_4871);
or U6616 (N_6616,N_5734,N_4495);
or U6617 (N_6617,N_5899,N_5944);
nand U6618 (N_6618,N_5749,N_6038);
and U6619 (N_6619,N_5706,N_4107);
and U6620 (N_6620,N_4964,N_4428);
and U6621 (N_6621,N_4513,N_4874);
nand U6622 (N_6622,N_6101,N_5881);
xnor U6623 (N_6623,N_3770,N_5180);
and U6624 (N_6624,N_4732,N_5138);
or U6625 (N_6625,N_5456,N_4364);
or U6626 (N_6626,N_5170,N_5342);
nand U6627 (N_6627,N_4611,N_4697);
or U6628 (N_6628,N_5490,N_3390);
and U6629 (N_6629,N_3717,N_4210);
xor U6630 (N_6630,N_6217,N_3829);
nand U6631 (N_6631,N_4057,N_3773);
nand U6632 (N_6632,N_5214,N_5544);
or U6633 (N_6633,N_3380,N_5813);
and U6634 (N_6634,N_3395,N_4297);
nor U6635 (N_6635,N_6234,N_3288);
nand U6636 (N_6636,N_6152,N_4088);
nor U6637 (N_6637,N_3796,N_4266);
or U6638 (N_6638,N_3448,N_3263);
and U6639 (N_6639,N_4991,N_4347);
nor U6640 (N_6640,N_5918,N_4310);
or U6641 (N_6641,N_5526,N_3686);
nor U6642 (N_6642,N_6143,N_4191);
nor U6643 (N_6643,N_4047,N_3553);
nand U6644 (N_6644,N_6147,N_5197);
xor U6645 (N_6645,N_4722,N_5927);
or U6646 (N_6646,N_4692,N_3529);
nor U6647 (N_6647,N_5034,N_5924);
nand U6648 (N_6648,N_4824,N_5916);
xnor U6649 (N_6649,N_6044,N_3965);
nor U6650 (N_6650,N_3342,N_6030);
and U6651 (N_6651,N_3724,N_5397);
and U6652 (N_6652,N_5472,N_5376);
and U6653 (N_6653,N_5532,N_3304);
xor U6654 (N_6654,N_3684,N_5217);
nand U6655 (N_6655,N_3340,N_4071);
nand U6656 (N_6656,N_4209,N_3764);
or U6657 (N_6657,N_5991,N_3334);
nand U6658 (N_6658,N_5554,N_3927);
xnor U6659 (N_6659,N_3942,N_3846);
or U6660 (N_6660,N_4326,N_3330);
or U6661 (N_6661,N_3221,N_6040);
and U6662 (N_6662,N_4208,N_4757);
xor U6663 (N_6663,N_4540,N_4629);
nor U6664 (N_6664,N_4093,N_5392);
or U6665 (N_6665,N_4506,N_5110);
nand U6666 (N_6666,N_3515,N_6187);
or U6667 (N_6667,N_4267,N_5136);
nor U6668 (N_6668,N_5563,N_5602);
nand U6669 (N_6669,N_5293,N_4970);
nor U6670 (N_6670,N_5545,N_5640);
nor U6671 (N_6671,N_5181,N_5043);
and U6672 (N_6672,N_3772,N_4555);
and U6673 (N_6673,N_3297,N_3128);
nand U6674 (N_6674,N_5789,N_5304);
xor U6675 (N_6675,N_6240,N_5223);
or U6676 (N_6676,N_4307,N_4158);
and U6677 (N_6677,N_5429,N_4975);
nor U6678 (N_6678,N_6138,N_5690);
and U6679 (N_6679,N_5417,N_5710);
and U6680 (N_6680,N_5428,N_5576);
and U6681 (N_6681,N_4155,N_5331);
and U6682 (N_6682,N_4474,N_5705);
or U6683 (N_6683,N_3712,N_4369);
and U6684 (N_6684,N_4771,N_5770);
and U6685 (N_6685,N_4180,N_3472);
or U6686 (N_6686,N_4242,N_4637);
and U6687 (N_6687,N_5107,N_4309);
nand U6688 (N_6688,N_3752,N_4572);
nor U6689 (N_6689,N_5848,N_3650);
nor U6690 (N_6690,N_3274,N_5683);
nor U6691 (N_6691,N_4014,N_5772);
nor U6692 (N_6692,N_6199,N_5714);
nand U6693 (N_6693,N_4589,N_4149);
and U6694 (N_6694,N_4685,N_4979);
and U6695 (N_6695,N_5607,N_5345);
or U6696 (N_6696,N_4493,N_5297);
nand U6697 (N_6697,N_5371,N_5672);
or U6698 (N_6698,N_5306,N_5261);
nor U6699 (N_6699,N_5252,N_5227);
and U6700 (N_6700,N_5459,N_4051);
and U6701 (N_6701,N_5762,N_4371);
nor U6702 (N_6702,N_4029,N_3238);
and U6703 (N_6703,N_3601,N_5149);
or U6704 (N_6704,N_3908,N_5617);
nor U6705 (N_6705,N_5497,N_3224);
nor U6706 (N_6706,N_6135,N_4101);
nor U6707 (N_6707,N_3700,N_4456);
or U6708 (N_6708,N_5788,N_5904);
and U6709 (N_6709,N_4482,N_4033);
and U6710 (N_6710,N_4219,N_3777);
and U6711 (N_6711,N_4171,N_3435);
or U6712 (N_6712,N_4519,N_5385);
nor U6713 (N_6713,N_3950,N_3543);
or U6714 (N_6714,N_5507,N_4997);
or U6715 (N_6715,N_4390,N_3241);
nor U6716 (N_6716,N_6024,N_3155);
or U6717 (N_6717,N_3595,N_3791);
xnor U6718 (N_6718,N_4853,N_5745);
nor U6719 (N_6719,N_4858,N_3205);
and U6720 (N_6720,N_3964,N_3281);
or U6721 (N_6721,N_6195,N_4329);
or U6722 (N_6722,N_6212,N_5016);
xnor U6723 (N_6723,N_5002,N_4690);
nor U6724 (N_6724,N_4517,N_5022);
and U6725 (N_6725,N_6146,N_4763);
and U6726 (N_6726,N_5583,N_5374);
or U6727 (N_6727,N_5158,N_4584);
nor U6728 (N_6728,N_3471,N_4895);
and U6729 (N_6729,N_3194,N_6059);
xnor U6730 (N_6730,N_3363,N_3558);
xnor U6731 (N_6731,N_4263,N_3417);
nand U6732 (N_6732,N_4477,N_5339);
and U6733 (N_6733,N_3497,N_4251);
and U6734 (N_6734,N_4972,N_3160);
and U6735 (N_6735,N_5538,N_5892);
or U6736 (N_6736,N_5600,N_6075);
or U6737 (N_6737,N_3444,N_5675);
or U6738 (N_6738,N_3337,N_3972);
nor U6739 (N_6739,N_4373,N_3588);
nand U6740 (N_6740,N_4260,N_3824);
nor U6741 (N_6741,N_5909,N_3872);
or U6742 (N_6742,N_3441,N_3836);
or U6743 (N_6743,N_3247,N_5654);
and U6744 (N_6744,N_3422,N_5958);
nand U6745 (N_6745,N_4100,N_5077);
or U6746 (N_6746,N_3411,N_5757);
xor U6747 (N_6747,N_3844,N_4986);
or U6748 (N_6748,N_3733,N_5282);
and U6749 (N_6749,N_3565,N_4352);
and U6750 (N_6750,N_5006,N_3722);
or U6751 (N_6751,N_4325,N_6115);
nor U6752 (N_6752,N_4204,N_6121);
and U6753 (N_6753,N_5872,N_5774);
or U6754 (N_6754,N_4366,N_4553);
xor U6755 (N_6755,N_4281,N_4011);
and U6756 (N_6756,N_3389,N_6112);
nor U6757 (N_6757,N_5354,N_5994);
or U6758 (N_6758,N_5804,N_4087);
and U6759 (N_6759,N_4289,N_4931);
and U6760 (N_6760,N_4980,N_5771);
nand U6761 (N_6761,N_6096,N_5238);
nor U6762 (N_6762,N_4198,N_3227);
nor U6763 (N_6763,N_3421,N_5656);
or U6764 (N_6764,N_6002,N_6149);
and U6765 (N_6765,N_4710,N_5239);
nand U6766 (N_6766,N_3406,N_3778);
nand U6767 (N_6767,N_4689,N_3259);
nand U6768 (N_6768,N_4758,N_5543);
nor U6769 (N_6769,N_4142,N_4131);
nor U6770 (N_6770,N_4888,N_4750);
nand U6771 (N_6771,N_5598,N_5303);
nor U6772 (N_6772,N_4800,N_4674);
nand U6773 (N_6773,N_3737,N_5609);
or U6774 (N_6774,N_6036,N_3812);
and U6775 (N_6775,N_4902,N_5268);
nor U6776 (N_6776,N_3481,N_5778);
nor U6777 (N_6777,N_5915,N_4193);
nand U6778 (N_6778,N_6136,N_5680);
xor U6779 (N_6779,N_4720,N_4786);
nand U6780 (N_6780,N_4081,N_3137);
and U6781 (N_6781,N_5039,N_3439);
and U6782 (N_6782,N_3710,N_4062);
nand U6783 (N_6783,N_3293,N_4544);
and U6784 (N_6784,N_5530,N_3162);
and U6785 (N_6785,N_4870,N_4491);
nor U6786 (N_6786,N_5271,N_3518);
and U6787 (N_6787,N_4693,N_3436);
nand U6788 (N_6788,N_3163,N_4086);
or U6789 (N_6789,N_3509,N_5401);
nor U6790 (N_6790,N_3903,N_5301);
nand U6791 (N_6791,N_5611,N_5460);
nand U6792 (N_6792,N_3853,N_3258);
nand U6793 (N_6793,N_3997,N_4174);
or U6794 (N_6794,N_4079,N_3570);
nor U6795 (N_6795,N_5403,N_4681);
nand U6796 (N_6796,N_3804,N_5037);
or U6797 (N_6797,N_4315,N_4489);
nor U6798 (N_6798,N_5319,N_6026);
and U6799 (N_6799,N_4658,N_4562);
xnor U6800 (N_6800,N_4092,N_3468);
nand U6801 (N_6801,N_5529,N_5100);
nor U6802 (N_6802,N_6007,N_5756);
nand U6803 (N_6803,N_6248,N_5520);
xnor U6804 (N_6804,N_6047,N_4318);
and U6805 (N_6805,N_4925,N_3461);
or U6806 (N_6806,N_3134,N_4688);
and U6807 (N_6807,N_6010,N_5931);
nand U6808 (N_6808,N_5340,N_4976);
xnor U6809 (N_6809,N_5399,N_6014);
and U6810 (N_6810,N_4061,N_5305);
xnor U6811 (N_6811,N_3218,N_3914);
nor U6812 (N_6812,N_4413,N_5874);
nand U6813 (N_6813,N_5208,N_5477);
nor U6814 (N_6814,N_5312,N_4196);
nand U6815 (N_6815,N_4272,N_5050);
and U6816 (N_6816,N_3901,N_4427);
nand U6817 (N_6817,N_4140,N_6128);
or U6818 (N_6818,N_5160,N_5212);
and U6819 (N_6819,N_5017,N_3307);
nor U6820 (N_6820,N_3993,N_5837);
nor U6821 (N_6821,N_6155,N_5836);
and U6822 (N_6822,N_4487,N_5368);
xnor U6823 (N_6823,N_4122,N_3991);
nor U6824 (N_6824,N_3789,N_3364);
xor U6825 (N_6825,N_5215,N_5998);
nand U6826 (N_6826,N_4349,N_4049);
nor U6827 (N_6827,N_4488,N_5078);
and U6828 (N_6828,N_4028,N_6164);
and U6829 (N_6829,N_5900,N_4576);
nand U6830 (N_6830,N_5649,N_3547);
and U6831 (N_6831,N_4389,N_4543);
xnor U6832 (N_6832,N_3313,N_3278);
and U6833 (N_6833,N_4376,N_3308);
nor U6834 (N_6834,N_4298,N_5679);
nand U6835 (N_6835,N_5481,N_4733);
nor U6836 (N_6836,N_4346,N_5291);
nand U6837 (N_6837,N_5593,N_3762);
nand U6838 (N_6838,N_4203,N_4930);
nor U6839 (N_6839,N_5328,N_3678);
or U6840 (N_6840,N_3615,N_4891);
and U6841 (N_6841,N_4220,N_4955);
or U6842 (N_6842,N_4604,N_5264);
or U6843 (N_6843,N_5467,N_5819);
nand U6844 (N_6844,N_3491,N_4153);
nand U6845 (N_6845,N_4919,N_5550);
nand U6846 (N_6846,N_5255,N_5503);
nor U6847 (N_6847,N_5243,N_4694);
and U6848 (N_6848,N_5125,N_4270);
nor U6849 (N_6849,N_5299,N_4350);
and U6850 (N_6850,N_3400,N_3729);
xnor U6851 (N_6851,N_3185,N_5806);
and U6852 (N_6852,N_6207,N_3357);
and U6853 (N_6853,N_5628,N_3640);
xnor U6854 (N_6854,N_6006,N_5069);
nor U6855 (N_6855,N_6097,N_4737);
and U6856 (N_6856,N_5421,N_3249);
or U6857 (N_6857,N_4083,N_3156);
or U6858 (N_6858,N_4013,N_5704);
and U6859 (N_6859,N_5537,N_5887);
and U6860 (N_6860,N_4040,N_3947);
or U6861 (N_6861,N_4016,N_5830);
xnor U6862 (N_6862,N_4974,N_3755);
and U6863 (N_6863,N_4189,N_4761);
xnor U6864 (N_6864,N_5979,N_4785);
nor U6865 (N_6865,N_4036,N_5114);
xnor U6866 (N_6866,N_3575,N_5689);
and U6867 (N_6867,N_5883,N_5729);
and U6868 (N_6868,N_4911,N_5647);
and U6869 (N_6869,N_4332,N_5572);
or U6870 (N_6870,N_3718,N_4216);
or U6871 (N_6871,N_5353,N_6031);
xnor U6872 (N_6872,N_4920,N_4798);
nor U6873 (N_6873,N_5661,N_5489);
nand U6874 (N_6874,N_3502,N_4015);
nor U6875 (N_6875,N_3984,N_4089);
nor U6876 (N_6876,N_3285,N_5347);
nand U6877 (N_6877,N_3312,N_5987);
and U6878 (N_6878,N_5587,N_3431);
and U6879 (N_6879,N_5442,N_4541);
nor U6880 (N_6880,N_5265,N_4603);
or U6881 (N_6881,N_4330,N_5826);
nor U6882 (N_6882,N_3830,N_4616);
nand U6883 (N_6883,N_5698,N_3305);
nand U6884 (N_6884,N_5948,N_4112);
nand U6885 (N_6885,N_6054,N_5977);
and U6886 (N_6886,N_5191,N_6055);
xor U6887 (N_6887,N_4606,N_4118);
or U6888 (N_6888,N_5933,N_3631);
nand U6889 (N_6889,N_5012,N_3926);
nand U6890 (N_6890,N_3941,N_4814);
nor U6891 (N_6891,N_5218,N_4819);
and U6892 (N_6892,N_4060,N_5570);
nor U6893 (N_6893,N_4619,N_4434);
and U6894 (N_6894,N_5686,N_6196);
and U6895 (N_6895,N_4725,N_5852);
and U6896 (N_6896,N_3835,N_5959);
xnor U6897 (N_6897,N_5907,N_5233);
and U6898 (N_6898,N_5336,N_5581);
or U6899 (N_6899,N_3501,N_4128);
or U6900 (N_6900,N_6016,N_5127);
or U6901 (N_6901,N_3391,N_3768);
xnor U6902 (N_6902,N_4687,N_3597);
nor U6903 (N_6903,N_5449,N_5474);
nor U6904 (N_6904,N_5171,N_5928);
nor U6905 (N_6905,N_4890,N_6209);
or U6906 (N_6906,N_4605,N_4457);
nor U6907 (N_6907,N_5410,N_3856);
nor U6908 (N_6908,N_4886,N_5229);
or U6909 (N_6909,N_3131,N_4524);
xor U6910 (N_6910,N_3657,N_3489);
or U6911 (N_6911,N_3758,N_5652);
nor U6912 (N_6912,N_5603,N_5921);
and U6913 (N_6913,N_4638,N_5651);
and U6914 (N_6914,N_3534,N_4708);
nand U6915 (N_6915,N_4429,N_6189);
nand U6916 (N_6916,N_6241,N_3381);
nor U6917 (N_6917,N_3960,N_5957);
nand U6918 (N_6918,N_3254,N_5084);
nor U6919 (N_6919,N_4768,N_5728);
xnor U6920 (N_6920,N_3333,N_4968);
nand U6921 (N_6921,N_6124,N_3584);
nor U6922 (N_6922,N_4444,N_4952);
nand U6923 (N_6923,N_5903,N_5274);
and U6924 (N_6924,N_4067,N_4961);
nand U6925 (N_6925,N_4684,N_5982);
nand U6926 (N_6926,N_4066,N_5513);
nor U6927 (N_6927,N_5751,N_5021);
nor U6928 (N_6928,N_4410,N_5475);
nand U6929 (N_6929,N_3831,N_4990);
nand U6930 (N_6930,N_5875,N_5764);
nor U6931 (N_6931,N_4706,N_3362);
nand U6932 (N_6932,N_4257,N_5865);
nand U6933 (N_6933,N_4365,N_5962);
nand U6934 (N_6934,N_6099,N_4006);
or U6935 (N_6935,N_5222,N_5280);
nand U6936 (N_6936,N_5839,N_4967);
nor U6937 (N_6937,N_5781,N_5426);
or U6938 (N_6938,N_3462,N_4445);
and U6939 (N_6939,N_4073,N_4595);
and U6940 (N_6940,N_3810,N_5873);
nor U6941 (N_6941,N_3924,N_4995);
nor U6942 (N_6942,N_5986,N_3905);
and U6943 (N_6943,N_3978,N_5953);
nor U6944 (N_6944,N_4126,N_6184);
nor U6945 (N_6945,N_4948,N_4973);
or U6946 (N_6946,N_5439,N_5357);
and U6947 (N_6947,N_6145,N_3354);
nor U6948 (N_6948,N_3723,N_4557);
nor U6949 (N_6949,N_4027,N_4863);
nor U6950 (N_6950,N_5070,N_3994);
or U6951 (N_6951,N_3151,N_4645);
nor U6952 (N_6952,N_4414,N_4613);
and U6953 (N_6953,N_4653,N_6165);
or U6954 (N_6954,N_5724,N_3165);
nor U6955 (N_6955,N_4008,N_5404);
xor U6956 (N_6956,N_4245,N_3298);
or U6957 (N_6957,N_3289,N_4538);
and U6958 (N_6958,N_4212,N_3680);
xor U6959 (N_6959,N_5932,N_3262);
xnor U6960 (N_6960,N_3922,N_5169);
nor U6961 (N_6961,N_5266,N_5963);
nor U6962 (N_6962,N_3748,N_4502);
nor U6963 (N_6963,N_3257,N_3644);
nor U6964 (N_6964,N_5896,N_3344);
nand U6965 (N_6965,N_4662,N_5605);
nor U6966 (N_6966,N_5486,N_3219);
or U6967 (N_6967,N_4173,N_3415);
or U6968 (N_6968,N_4510,N_4825);
or U6969 (N_6969,N_5259,N_3745);
xnor U6970 (N_6970,N_4348,N_3784);
nand U6971 (N_6971,N_3687,N_4304);
nand U6972 (N_6972,N_6027,N_3434);
nor U6973 (N_6973,N_5226,N_5663);
xnor U6974 (N_6974,N_4211,N_4184);
or U6975 (N_6975,N_4915,N_3656);
nand U6976 (N_6976,N_5285,N_4358);
and U6977 (N_6977,N_5461,N_5975);
or U6978 (N_6978,N_3370,N_4368);
and U6979 (N_6979,N_5784,N_4642);
xnor U6980 (N_6980,N_3794,N_3619);
nor U6981 (N_6981,N_5323,N_3280);
and U6982 (N_6982,N_4941,N_4508);
or U6983 (N_6983,N_5007,N_3206);
nand U6984 (N_6984,N_6141,N_3987);
or U6985 (N_6985,N_6197,N_3714);
nor U6986 (N_6986,N_4119,N_3867);
nand U6987 (N_6987,N_3383,N_3237);
nand U6988 (N_6988,N_5485,N_3514);
or U6989 (N_6989,N_4151,N_4649);
nand U6990 (N_6990,N_5415,N_5488);
or U6991 (N_6991,N_6243,N_4754);
nor U6992 (N_6992,N_5389,N_5790);
nand U6993 (N_6993,N_6108,N_5853);
nand U6994 (N_6994,N_5205,N_3890);
nor U6995 (N_6995,N_3248,N_3385);
xnor U6996 (N_6996,N_6210,N_4514);
or U6997 (N_6997,N_3751,N_6194);
and U6998 (N_6998,N_4218,N_5878);
and U6999 (N_6999,N_5669,N_4454);
xnor U7000 (N_7000,N_5895,N_5232);
and U7001 (N_7001,N_5047,N_3429);
or U7002 (N_7002,N_5279,N_5221);
nand U7003 (N_7003,N_3676,N_3967);
or U7004 (N_7004,N_5955,N_5269);
nand U7005 (N_7005,N_4556,N_4178);
and U7006 (N_7006,N_4998,N_6222);
nand U7007 (N_7007,N_6018,N_3168);
or U7008 (N_7008,N_3244,N_4620);
nor U7009 (N_7009,N_3174,N_5692);
xor U7010 (N_7010,N_6019,N_4516);
and U7011 (N_7011,N_3426,N_4402);
nand U7012 (N_7012,N_4949,N_5091);
and U7013 (N_7013,N_3627,N_4936);
nand U7014 (N_7014,N_5684,N_5201);
and U7015 (N_7015,N_3782,N_4801);
xnor U7016 (N_7016,N_4899,N_5318);
nand U7017 (N_7017,N_4614,N_4021);
nand U7018 (N_7018,N_5738,N_5407);
nand U7019 (N_7019,N_5178,N_3761);
or U7020 (N_7020,N_5691,N_4759);
nor U7021 (N_7021,N_5687,N_4904);
and U7022 (N_7022,N_4426,N_4082);
and U7023 (N_7023,N_4717,N_5787);
nor U7024 (N_7024,N_6239,N_5241);
and U7025 (N_7025,N_5810,N_4847);
nor U7026 (N_7026,N_5351,N_4157);
xor U7027 (N_7027,N_4583,N_4959);
xor U7028 (N_7028,N_5750,N_4084);
nor U7029 (N_7029,N_3366,N_5635);
nand U7030 (N_7030,N_5148,N_5740);
nor U7031 (N_7031,N_5758,N_5767);
and U7032 (N_7032,N_4032,N_3743);
or U7033 (N_7033,N_6087,N_5843);
or U7034 (N_7034,N_4059,N_4361);
nand U7035 (N_7035,N_5518,N_4903);
nor U7036 (N_7036,N_5743,N_3734);
or U7037 (N_7037,N_3183,N_6142);
or U7038 (N_7038,N_3665,N_4162);
nor U7039 (N_7039,N_5522,N_4593);
nand U7040 (N_7040,N_4319,N_4838);
or U7041 (N_7041,N_4610,N_5019);
and U7042 (N_7042,N_6062,N_4788);
xor U7043 (N_7043,N_3573,N_4751);
nand U7044 (N_7044,N_5973,N_4360);
xnor U7045 (N_7045,N_6022,N_4091);
xor U7046 (N_7046,N_4052,N_5596);
or U7047 (N_7047,N_5741,N_4306);
or U7048 (N_7048,N_5695,N_5536);
and U7049 (N_7049,N_4372,N_6215);
and U7050 (N_7050,N_3253,N_3499);
or U7051 (N_7051,N_5408,N_4268);
nand U7052 (N_7052,N_5753,N_6203);
nor U7053 (N_7053,N_3368,N_4104);
or U7054 (N_7054,N_3583,N_3727);
and U7055 (N_7055,N_3136,N_3449);
nor U7056 (N_7056,N_3820,N_5861);
and U7057 (N_7057,N_4736,N_4849);
nor U7058 (N_7058,N_4288,N_3179);
nor U7059 (N_7059,N_4762,N_3379);
and U7060 (N_7060,N_4038,N_3367);
xor U7061 (N_7061,N_5584,N_4007);
and U7062 (N_7062,N_4147,N_3269);
nand U7063 (N_7063,N_4590,N_4192);
nand U7064 (N_7064,N_4906,N_3178);
and U7065 (N_7065,N_5202,N_4591);
or U7066 (N_7066,N_3267,N_4864);
nor U7067 (N_7067,N_5800,N_5341);
and U7068 (N_7068,N_5179,N_5832);
or U7069 (N_7069,N_4163,N_4789);
or U7070 (N_7070,N_4598,N_3467);
nor U7071 (N_7071,N_4826,N_4988);
nor U7072 (N_7072,N_4834,N_3946);
nor U7073 (N_7073,N_3324,N_5831);
nand U7074 (N_7074,N_4114,N_4335);
or U7075 (N_7075,N_5292,N_5384);
nand U7076 (N_7076,N_3492,N_5495);
nand U7077 (N_7077,N_3474,N_5032);
or U7078 (N_7078,N_5230,N_5947);
or U7079 (N_7079,N_4133,N_4860);
or U7080 (N_7080,N_3554,N_5521);
or U7081 (N_7081,N_4070,N_4507);
nand U7082 (N_7082,N_3881,N_5542);
nor U7083 (N_7083,N_4076,N_5662);
and U7084 (N_7084,N_5752,N_5917);
nand U7085 (N_7085,N_5424,N_5023);
and U7086 (N_7086,N_5911,N_3825);
nor U7087 (N_7087,N_4818,N_5284);
nand U7088 (N_7088,N_4320,N_5330);
nor U7089 (N_7089,N_5062,N_3458);
nand U7090 (N_7090,N_4393,N_4657);
xor U7091 (N_7091,N_4695,N_4534);
nand U7092 (N_7092,N_3493,N_4873);
nand U7093 (N_7093,N_5990,N_4600);
nand U7094 (N_7094,N_4781,N_5278);
or U7095 (N_7095,N_6200,N_3833);
nand U7096 (N_7096,N_6218,N_6213);
or U7097 (N_7097,N_5769,N_5708);
nand U7098 (N_7098,N_6012,N_5589);
nor U7099 (N_7099,N_5400,N_4909);
nand U7100 (N_7100,N_3859,N_4531);
and U7101 (N_7101,N_4287,N_3598);
and U7102 (N_7102,N_5258,N_6110);
and U7103 (N_7103,N_5871,N_3943);
xor U7104 (N_7104,N_3805,N_5406);
and U7105 (N_7105,N_5388,N_4236);
nor U7106 (N_7106,N_4095,N_4197);
nand U7107 (N_7107,N_5203,N_3432);
nor U7108 (N_7108,N_4942,N_3790);
xnor U7109 (N_7109,N_4672,N_3732);
or U7110 (N_7110,N_3469,N_4773);
nand U7111 (N_7111,N_5057,N_4981);
and U7112 (N_7112,N_5298,N_5009);
xor U7113 (N_7113,N_6180,N_5159);
nor U7114 (N_7114,N_4435,N_4525);
nand U7115 (N_7115,N_5207,N_3699);
xor U7116 (N_7116,N_5557,N_5054);
nand U7117 (N_7117,N_3888,N_3919);
nand U7118 (N_7118,N_3147,N_3276);
and U7119 (N_7119,N_4438,N_6105);
nor U7120 (N_7120,N_6046,N_3817);
or U7121 (N_7121,N_5275,N_5674);
or U7122 (N_7122,N_3871,N_5644);
or U7123 (N_7123,N_5010,N_3217);
or U7124 (N_7124,N_3171,N_3531);
nand U7125 (N_7125,N_5730,N_3286);
and U7126 (N_7126,N_6133,N_5822);
or U7127 (N_7127,N_4535,N_3886);
nor U7128 (N_7128,N_3878,N_6227);
or U7129 (N_7129,N_3821,N_5466);
or U7130 (N_7130,N_3314,N_6177);
and U7131 (N_7131,N_5245,N_5910);
and U7132 (N_7132,N_4129,N_5580);
nor U7133 (N_7133,N_4205,N_5254);
or U7134 (N_7134,N_3279,N_3332);
nor U7135 (N_7135,N_3694,N_4567);
or U7136 (N_7136,N_3564,N_3749);
xor U7137 (N_7137,N_6109,N_5124);
and U7138 (N_7138,N_5523,N_5864);
nand U7139 (N_7139,N_3201,N_3552);
and U7140 (N_7140,N_4797,N_3295);
nand U7141 (N_7141,N_3738,N_5128);
xor U7142 (N_7142,N_5721,N_4019);
or U7143 (N_7143,N_4385,N_3316);
nor U7144 (N_7144,N_4124,N_3689);
xor U7145 (N_7145,N_4408,N_5858);
nor U7146 (N_7146,N_4328,N_4526);
and U7147 (N_7147,N_5561,N_6211);
nor U7148 (N_7148,N_5132,N_4927);
nand U7149 (N_7149,N_4206,N_4043);
and U7150 (N_7150,N_5235,N_5102);
xnor U7151 (N_7151,N_4339,N_4676);
nor U7152 (N_7152,N_3454,N_6011);
nand U7153 (N_7153,N_4054,N_4625);
xnor U7154 (N_7154,N_4446,N_4542);
or U7155 (N_7155,N_3559,N_3192);
and U7156 (N_7156,N_5321,N_4570);
xnor U7157 (N_7157,N_4987,N_3393);
xnor U7158 (N_7158,N_3181,N_4779);
nor U7159 (N_7159,N_3803,N_6081);
or U7160 (N_7160,N_5494,N_3260);
or U7161 (N_7161,N_5920,N_3430);
xor U7162 (N_7162,N_5720,N_4492);
nor U7163 (N_7163,N_3986,N_3571);
and U7164 (N_7164,N_3920,N_4635);
xnor U7165 (N_7165,N_4701,N_4010);
or U7166 (N_7166,N_5956,N_4966);
or U7167 (N_7167,N_4451,N_5624);
and U7168 (N_7168,N_3655,N_3282);
nor U7169 (N_7169,N_4141,N_4499);
or U7170 (N_7170,N_5763,N_4794);
nor U7171 (N_7171,N_3407,N_4090);
nor U7172 (N_7172,N_6084,N_3159);
or U7173 (N_7173,N_3373,N_3404);
or U7174 (N_7174,N_4700,N_5033);
or U7175 (N_7175,N_4106,N_4386);
nor U7176 (N_7176,N_6245,N_4166);
xor U7177 (N_7177,N_3606,N_5086);
or U7178 (N_7178,N_4618,N_5395);
nand U7179 (N_7179,N_4085,N_5760);
nand U7180 (N_7180,N_4881,N_3496);
nor U7181 (N_7181,N_3879,N_5464);
or U7182 (N_7182,N_5068,N_6013);
nor U7183 (N_7183,N_3968,N_6070);
xnor U7184 (N_7184,N_4828,N_5786);
nor U7185 (N_7185,N_5123,N_4712);
and U7186 (N_7186,N_5923,N_4569);
or U7187 (N_7187,N_3528,N_3414);
xnor U7188 (N_7188,N_5618,N_5134);
nand U7189 (N_7189,N_4777,N_4962);
or U7190 (N_7190,N_5165,N_4442);
nor U7191 (N_7191,N_4900,N_4237);
and U7192 (N_7192,N_4256,N_5454);
nand U7193 (N_7193,N_4305,N_4954);
and U7194 (N_7194,N_5115,N_6172);
or U7195 (N_7195,N_6247,N_3125);
nand U7196 (N_7196,N_6068,N_5950);
nor U7197 (N_7197,N_3816,N_5157);
nand U7198 (N_7198,N_3142,N_4050);
nand U7199 (N_7199,N_5849,N_4897);
xor U7200 (N_7200,N_5052,N_3451);
nand U7201 (N_7201,N_4566,N_4850);
nand U7202 (N_7202,N_5627,N_3144);
xor U7203 (N_7203,N_3240,N_3938);
nand U7204 (N_7204,N_5386,N_4099);
or U7205 (N_7205,N_3936,N_5026);
nor U7206 (N_7206,N_5604,N_3675);
xor U7207 (N_7207,N_4947,N_3284);
nor U7208 (N_7208,N_4741,N_5725);
nand U7209 (N_7209,N_5512,N_4467);
or U7210 (N_7210,N_4034,N_5553);
and U7211 (N_7211,N_4585,N_5716);
and U7212 (N_7212,N_3539,N_4983);
or U7213 (N_7213,N_5673,N_4313);
xnor U7214 (N_7214,N_5623,N_5366);
nor U7215 (N_7215,N_5478,N_3251);
nand U7216 (N_7216,N_3277,N_3720);
and U7217 (N_7217,N_4023,N_4255);
and U7218 (N_7218,N_4337,N_5013);
nand U7219 (N_7219,N_4481,N_3645);
nor U7220 (N_7220,N_3563,N_5574);
and U7221 (N_7221,N_3970,N_3880);
or U7222 (N_7222,N_4116,N_5586);
nor U7223 (N_7223,N_4511,N_4851);
nand U7224 (N_7224,N_3862,N_6077);
or U7225 (N_7225,N_6158,N_5458);
nand U7226 (N_7226,N_5629,N_4351);
nand U7227 (N_7227,N_4441,N_3129);
and U7228 (N_7228,N_4283,N_5311);
nand U7229 (N_7229,N_5236,N_4123);
and U7230 (N_7230,N_4774,N_3721);
nand U7231 (N_7231,N_5869,N_4659);
nand U7232 (N_7232,N_4529,N_5500);
nor U7233 (N_7233,N_4669,N_6139);
and U7234 (N_7234,N_5137,N_5176);
and U7235 (N_7235,N_4929,N_5894);
nor U7236 (N_7236,N_4679,N_4334);
and U7237 (N_7237,N_5036,N_5785);
nor U7238 (N_7238,N_4755,N_3975);
or U7239 (N_7239,N_3662,N_3215);
nand U7240 (N_7240,N_3639,N_3154);
or U7241 (N_7241,N_3877,N_4294);
and U7242 (N_7242,N_3419,N_3296);
and U7243 (N_7243,N_4146,N_5713);
xnor U7244 (N_7244,N_4776,N_3387);
nor U7245 (N_7245,N_4221,N_5167);
and U7246 (N_7246,N_4802,N_5568);
nor U7247 (N_7247,N_6107,N_5835);
nor U7248 (N_7248,N_3483,N_5465);
nor U7249 (N_7249,N_5363,N_6083);
nand U7250 (N_7250,N_3906,N_3378);
nand U7251 (N_7251,N_4227,N_4588);
or U7252 (N_7252,N_3658,N_5560);
nand U7253 (N_7253,N_5855,N_5105);
and U7254 (N_7254,N_5231,N_3971);
nand U7255 (N_7255,N_4470,N_4880);
nand U7256 (N_7256,N_3701,N_5809);
and U7257 (N_7257,N_4164,N_5960);
xor U7258 (N_7258,N_5317,N_3170);
and U7259 (N_7259,N_5327,N_3377);
nor U7260 (N_7260,N_5815,N_3826);
nand U7261 (N_7261,N_3487,N_3149);
nand U7262 (N_7262,N_4686,N_3895);
nand U7263 (N_7263,N_3541,N_3150);
nand U7264 (N_7264,N_4609,N_5712);
or U7265 (N_7265,N_5228,N_5242);
nor U7266 (N_7266,N_5566,N_4958);
nand U7267 (N_7267,N_3742,N_3408);
xnor U7268 (N_7268,N_5650,N_5514);
and U7269 (N_7269,N_5122,N_5793);
nand U7270 (N_7270,N_5484,N_3319);
and U7271 (N_7271,N_5445,N_5420);
and U7272 (N_7272,N_5626,N_3230);
and U7273 (N_7273,N_5087,N_4889);
nand U7274 (N_7274,N_5281,N_5688);
and U7275 (N_7275,N_4599,N_6157);
nand U7276 (N_7276,N_5324,N_3909);
nor U7277 (N_7277,N_4387,N_5777);
nand U7278 (N_7278,N_5194,N_3962);
nor U7279 (N_7279,N_3126,N_3667);
and U7280 (N_7280,N_5360,N_4815);
xor U7281 (N_7281,N_3299,N_4134);
nand U7282 (N_7282,N_3594,N_4943);
nor U7283 (N_7283,N_5031,N_5028);
or U7284 (N_7284,N_5965,N_5027);
nand U7285 (N_7285,N_3562,N_3709);
nand U7286 (N_7286,N_5823,N_5450);
and U7287 (N_7287,N_3806,N_5625);
or U7288 (N_7288,N_5131,N_4494);
nor U7289 (N_7289,N_4002,N_4823);
and U7290 (N_7290,N_4419,N_4564);
nand U7291 (N_7291,N_5997,N_5531);
nand U7292 (N_7292,N_3864,N_4641);
nand U7293 (N_7293,N_5886,N_4024);
nand U7294 (N_7294,N_5565,N_5187);
and U7295 (N_7295,N_5048,N_5314);
nor U7296 (N_7296,N_5739,N_4213);
nor U7297 (N_7297,N_3456,N_4505);
xnor U7298 (N_7298,N_3345,N_3973);
xor U7299 (N_7299,N_6032,N_5558);
nand U7300 (N_7300,N_5735,N_3235);
nor U7301 (N_7301,N_4752,N_4848);
xor U7302 (N_7302,N_4957,N_5516);
and U7303 (N_7303,N_3851,N_3605);
or U7304 (N_7304,N_6225,N_3290);
xor U7305 (N_7305,N_3243,N_4115);
and U7306 (N_7306,N_5759,N_4394);
nor U7307 (N_7307,N_3460,N_4053);
or U7308 (N_7308,N_3898,N_4914);
and U7309 (N_7309,N_3611,N_4102);
and U7310 (N_7310,N_5130,N_4520);
nor U7311 (N_7311,N_6151,N_5089);
or U7312 (N_7312,N_3470,N_3809);
nand U7313 (N_7313,N_4671,N_6091);
nand U7314 (N_7314,N_5334,N_5889);
nand U7315 (N_7315,N_4078,N_4354);
and U7316 (N_7316,N_5694,N_6188);
nor U7317 (N_7317,N_4727,N_3523);
and U7318 (N_7318,N_3876,N_4816);
or U7319 (N_7319,N_4632,N_5967);
nor U7320 (N_7320,N_4579,N_5888);
xnor U7321 (N_7321,N_4113,N_6094);
nor U7322 (N_7322,N_5166,N_5954);
or U7323 (N_7323,N_4200,N_4181);
and U7324 (N_7324,N_5356,N_4291);
and U7325 (N_7325,N_5118,N_4560);
nor U7326 (N_7326,N_4624,N_5630);
nand U7327 (N_7327,N_3868,N_5715);
xnor U7328 (N_7328,N_4217,N_4452);
nand U7329 (N_7329,N_6106,N_5061);
or U7330 (N_7330,N_5527,N_5577);
nor U7331 (N_7331,N_3672,N_4407);
or U7332 (N_7332,N_3402,N_4575);
and U7333 (N_7333,N_5791,N_4224);
nor U7334 (N_7334,N_4001,N_3374);
nand U7335 (N_7335,N_5799,N_5247);
or U7336 (N_7336,N_5482,N_3145);
or U7337 (N_7337,N_5056,N_5359);
nand U7338 (N_7338,N_3341,N_4778);
nor U7339 (N_7339,N_3199,N_3592);
and U7340 (N_7340,N_6116,N_3196);
and U7341 (N_7341,N_4403,N_6159);
and U7342 (N_7342,N_3189,N_4246);
and U7343 (N_7343,N_3837,N_4552);
or U7344 (N_7344,N_5571,N_3896);
xnor U7345 (N_7345,N_5277,N_5073);
and U7346 (N_7346,N_4425,N_4644);
and U7347 (N_7347,N_3799,N_3593);
and U7348 (N_7348,N_5700,N_3464);
nor U7349 (N_7349,N_5657,N_4832);
and U7350 (N_7350,N_3513,N_5119);
xor U7351 (N_7351,N_4484,N_6161);
and U7352 (N_7352,N_5476,N_3590);
and U7353 (N_7353,N_4865,N_5156);
and U7354 (N_7354,N_5051,N_3843);
or U7355 (N_7355,N_3579,N_5862);
or U7356 (N_7356,N_4617,N_3127);
nor U7357 (N_7357,N_5562,N_3585);
and U7358 (N_7358,N_4321,N_3204);
nor U7359 (N_7359,N_6191,N_6082);
nor U7360 (N_7360,N_6201,N_4622);
nand U7361 (N_7361,N_4176,N_5365);
or U7362 (N_7362,N_4064,N_4110);
nor U7363 (N_7363,N_3925,N_4913);
nor U7364 (N_7364,N_5296,N_3445);
xnor U7365 (N_7365,N_4559,N_3934);
and U7366 (N_7366,N_5643,N_3708);
nor U7367 (N_7367,N_5642,N_4960);
nand U7368 (N_7368,N_3133,N_5310);
and U7369 (N_7369,N_4379,N_3275);
nand U7370 (N_7370,N_5801,N_3937);
nor U7371 (N_7371,N_5322,N_4724);
or U7372 (N_7372,N_3261,N_4478);
nor U7373 (N_7373,N_5446,N_4167);
nand U7374 (N_7374,N_6085,N_5608);
and U7375 (N_7375,N_5121,N_5190);
nor U7376 (N_7376,N_4806,N_4323);
nand U7377 (N_7377,N_4243,N_3416);
nor U7378 (N_7378,N_3807,N_3661);
xnor U7379 (N_7379,N_4439,N_5168);
xor U7380 (N_7380,N_3828,N_4682);
and U7381 (N_7381,N_3143,N_3336);
nand U7382 (N_7382,N_3187,N_4500);
nand U7383 (N_7383,N_4862,N_5974);
nand U7384 (N_7384,N_4299,N_4845);
and U7385 (N_7385,N_4654,N_4400);
and U7386 (N_7386,N_5945,N_5090);
or U7387 (N_7387,N_3386,N_3384);
or U7388 (N_7388,N_3283,N_4996);
and U7389 (N_7389,N_5902,N_5592);
nor U7390 (N_7390,N_5438,N_4661);
or U7391 (N_7391,N_4767,N_4459);
and U7392 (N_7392,N_4910,N_5983);
and U7393 (N_7393,N_4072,N_5369);
nand U7394 (N_7394,N_6117,N_3602);
nand U7395 (N_7395,N_5287,N_5192);
and U7396 (N_7396,N_3801,N_5856);
and U7397 (N_7397,N_3405,N_5315);
or U7398 (N_7398,N_5155,N_4269);
and U7399 (N_7399,N_4963,N_5079);
or U7400 (N_7400,N_6230,N_3478);
or U7401 (N_7401,N_4190,N_3303);
nor U7402 (N_7402,N_4840,N_4795);
or U7403 (N_7403,N_4461,N_4483);
or U7404 (N_7404,N_3349,N_3915);
and U7405 (N_7405,N_6066,N_4301);
nor U7406 (N_7406,N_4295,N_5798);
nor U7407 (N_7407,N_3634,N_3735);
nor U7408 (N_7408,N_5111,N_5551);
xnor U7409 (N_7409,N_4074,N_3857);
nor U7410 (N_7410,N_5726,N_3952);
and U7411 (N_7411,N_5104,N_3412);
or U7412 (N_7412,N_4586,N_5755);
and U7413 (N_7413,N_3815,N_4985);
or U7414 (N_7414,N_5189,N_5796);
and U7415 (N_7415,N_3450,N_5876);
nor U7416 (N_7416,N_4412,N_3190);
nor U7417 (N_7417,N_4944,N_3372);
and U7418 (N_7418,N_4292,N_4398);
nand U7419 (N_7419,N_3353,N_4744);
xnor U7420 (N_7420,N_3884,N_3265);
nor U7421 (N_7421,N_5044,N_4324);
or U7422 (N_7422,N_5040,N_5193);
xnor U7423 (N_7423,N_4504,N_3550);
nor U7424 (N_7424,N_5939,N_4265);
nand U7425 (N_7425,N_3207,N_4917);
nand U7426 (N_7426,N_5427,N_6216);
nand U7427 (N_7427,N_3530,N_6025);
xor U7428 (N_7428,N_3873,N_4696);
nand U7429 (N_7429,N_5667,N_5391);
nand U7430 (N_7430,N_5108,N_5140);
nor U7431 (N_7431,N_6179,N_5244);
or U7432 (N_7432,N_5075,N_5906);
xor U7433 (N_7433,N_4370,N_3325);
and U7434 (N_7434,N_4238,N_5885);
and U7435 (N_7435,N_4187,N_3682);
and U7436 (N_7436,N_6035,N_4170);
or U7437 (N_7437,N_4574,N_4842);
nand U7438 (N_7438,N_4547,N_3447);
or U7439 (N_7439,N_4201,N_4311);
nand U7440 (N_7440,N_3582,N_3326);
and U7441 (N_7441,N_6078,N_4844);
nor U7442 (N_7442,N_4443,N_5838);
and U7443 (N_7443,N_4905,N_3351);
nor U7444 (N_7444,N_4965,N_6021);
nor U7445 (N_7445,N_3961,N_4004);
nand U7446 (N_7446,N_3800,N_3220);
and U7447 (N_7447,N_4284,N_5289);
or U7448 (N_7448,N_3581,N_4630);
or U7449 (N_7449,N_5135,N_3309);
xnor U7450 (N_7450,N_4276,N_5470);
and U7451 (N_7451,N_3533,N_5030);
nor U7452 (N_7452,N_4879,N_4207);
and U7453 (N_7453,N_3935,N_5249);
and U7454 (N_7454,N_4790,N_3195);
or U7455 (N_7455,N_6048,N_4075);
nor U7456 (N_7456,N_3322,N_5637);
nor U7457 (N_7457,N_6193,N_6205);
nor U7458 (N_7458,N_4233,N_5213);
or U7459 (N_7459,N_4726,N_4673);
nor U7460 (N_7460,N_3427,N_3610);
or U7461 (N_7461,N_3666,N_5742);
nand U7462 (N_7462,N_3989,N_3630);
or U7463 (N_7463,N_4704,N_4721);
and U7464 (N_7464,N_4709,N_3910);
and U7465 (N_7465,N_3797,N_3775);
or U7466 (N_7466,N_4132,N_6080);
or U7467 (N_7467,N_3158,N_6056);
nand U7468 (N_7468,N_4308,N_5175);
or U7469 (N_7469,N_3690,N_3900);
xor U7470 (N_7470,N_5703,N_3287);
nand U7471 (N_7471,N_4887,N_4916);
nand U7472 (N_7472,N_5133,N_5106);
or U7473 (N_7473,N_4475,N_5765);
nor U7474 (N_7474,N_5335,N_3252);
and U7475 (N_7475,N_4515,N_4869);
nand U7476 (N_7476,N_4523,N_6166);
and U7477 (N_7477,N_6162,N_3203);
or U7478 (N_7478,N_3213,N_6126);
nor U7479 (N_7479,N_3659,N_3693);
nor U7480 (N_7480,N_5313,N_4417);
nor U7481 (N_7481,N_3521,N_5825);
xor U7482 (N_7482,N_4596,N_5547);
xor U7483 (N_7483,N_4230,N_3264);
nor U7484 (N_7484,N_4465,N_6098);
nor U7485 (N_7485,N_6127,N_5411);
or U7486 (N_7486,N_4764,N_4827);
or U7487 (N_7487,N_4651,N_5469);
nor U7488 (N_7488,N_5398,N_3705);
or U7489 (N_7489,N_6190,N_5702);
and U7490 (N_7490,N_4907,N_5188);
or U7491 (N_7491,N_4950,N_3490);
nand U7492 (N_7492,N_5126,N_3452);
nor U7493 (N_7493,N_5942,N_3209);
and U7494 (N_7494,N_5409,N_3208);
and U7495 (N_7495,N_5671,N_4745);
and U7496 (N_7496,N_3976,N_4293);
or U7497 (N_7497,N_3453,N_4835);
or U7498 (N_7498,N_5510,N_6103);
and U7499 (N_7499,N_4468,N_3182);
nor U7500 (N_7500,N_4937,N_3175);
and U7501 (N_7501,N_3863,N_5639);
nor U7502 (N_7502,N_4404,N_3510);
nor U7503 (N_7503,N_5519,N_5665);
and U7504 (N_7504,N_3681,N_3511);
nand U7505 (N_7505,N_4392,N_6073);
nand U7506 (N_7506,N_3486,N_5200);
and U7507 (N_7507,N_4753,N_3822);
nand U7508 (N_7508,N_6045,N_4821);
xor U7509 (N_7509,N_4839,N_5064);
and U7510 (N_7510,N_3500,N_3698);
nand U7511 (N_7511,N_5276,N_5390);
and U7512 (N_7512,N_5693,N_5224);
nand U7513 (N_7513,N_3466,N_3818);
nor U7514 (N_7514,N_3578,N_5879);
nor U7515 (N_7515,N_4409,N_3747);
or U7516 (N_7516,N_6020,N_5432);
xor U7517 (N_7517,N_4111,N_4241);
nand U7518 (N_7518,N_4537,N_3589);
nor U7519 (N_7519,N_3887,N_4792);
or U7520 (N_7520,N_6118,N_3902);
nand U7521 (N_7521,N_6185,N_5905);
nand U7522 (N_7522,N_4357,N_3932);
nand U7523 (N_7523,N_6049,N_4005);
nand U7524 (N_7524,N_6168,N_4714);
nor U7525 (N_7525,N_5709,N_5372);
or U7526 (N_7526,N_4035,N_4259);
nand U7527 (N_7527,N_5882,N_5941);
xnor U7528 (N_7528,N_4139,N_5333);
xor U7529 (N_7529,N_3428,N_5103);
nand U7530 (N_7530,N_5731,N_5564);
or U7531 (N_7531,N_6249,N_3757);
and U7532 (N_7532,N_3953,N_4536);
nor U7533 (N_7533,N_3546,N_3184);
and U7534 (N_7534,N_5969,N_3688);
nand U7535 (N_7535,N_4479,N_5951);
nand U7536 (N_7536,N_5631,N_5567);
and U7537 (N_7537,N_4951,N_4623);
and U7538 (N_7538,N_4249,N_3944);
nand U7539 (N_7539,N_4177,N_4117);
nand U7540 (N_7540,N_4121,N_5952);
and U7541 (N_7541,N_5621,N_4448);
nand U7542 (N_7542,N_5018,N_3827);
and U7543 (N_7543,N_3933,N_4331);
or U7544 (N_7544,N_5139,N_5147);
nand U7545 (N_7545,N_3343,N_3930);
nand U7546 (N_7546,N_3152,N_4353);
xor U7547 (N_7547,N_6053,N_5225);
or U7548 (N_7548,N_5290,N_6154);
nor U7549 (N_7549,N_5253,N_4127);
nor U7550 (N_7550,N_5940,N_4926);
nor U7551 (N_7551,N_5343,N_6005);
or U7552 (N_7552,N_4022,N_3540);
xor U7553 (N_7553,N_5447,N_5112);
or U7554 (N_7554,N_6114,N_3544);
or U7555 (N_7555,N_4341,N_3394);
or U7556 (N_7556,N_6042,N_3765);
nand U7557 (N_7557,N_5633,N_6183);
and U7558 (N_7558,N_4747,N_5196);
nand U7559 (N_7559,N_3660,N_5381);
nand U7560 (N_7560,N_6229,N_4471);
nor U7561 (N_7561,N_3870,N_5676);
and U7562 (N_7562,N_3157,N_5113);
nor U7563 (N_7563,N_5591,N_4994);
or U7564 (N_7564,N_4042,N_4405);
nand U7565 (N_7565,N_4563,N_4992);
xor U7566 (N_7566,N_3998,N_6050);
xor U7567 (N_7567,N_4420,N_3621);
nand U7568 (N_7568,N_6181,N_4831);
nor U7569 (N_7569,N_4715,N_4418);
or U7570 (N_7570,N_4175,N_5096);
xor U7571 (N_7571,N_4739,N_3977);
xor U7572 (N_7572,N_5539,N_4512);
xor U7573 (N_7573,N_4612,N_3889);
nor U7574 (N_7574,N_4314,N_3229);
nor U7575 (N_7575,N_3893,N_4796);
nand U7576 (N_7576,N_6244,N_3669);
nand U7577 (N_7577,N_5210,N_4568);
and U7578 (N_7578,N_3746,N_4993);
xnor U7579 (N_7579,N_4152,N_5448);
nor U7580 (N_7580,N_3695,N_6100);
and U7581 (N_7581,N_5405,N_6176);
nor U7582 (N_7582,N_5443,N_5556);
and U7583 (N_7583,N_4683,N_6064);
nor U7584 (N_7584,N_3629,N_4509);
or U7585 (N_7585,N_5925,N_3949);
and U7586 (N_7586,N_3850,N_3236);
or U7587 (N_7587,N_3180,N_5606);
or U7588 (N_7588,N_5913,N_4875);
nand U7589 (N_7589,N_3618,N_5501);
nand U7590 (N_7590,N_5868,N_3525);
nor U7591 (N_7591,N_3739,N_4956);
nand U7592 (N_7592,N_5499,N_3557);
and U7593 (N_7593,N_5794,N_4194);
and U7594 (N_7594,N_3371,N_3781);
nor U7595 (N_7595,N_3360,N_5095);
nor U7596 (N_7596,N_4150,N_6167);
nor U7597 (N_7597,N_5926,N_6130);
nand U7598 (N_7598,N_5812,N_4345);
and U7599 (N_7599,N_3702,N_5248);
nor U7600 (N_7600,N_4316,N_4277);
nor U7601 (N_7601,N_5658,N_4817);
or U7602 (N_7602,N_4135,N_6125);
nor U7603 (N_7603,N_3622,N_4145);
nor U7604 (N_7604,N_6034,N_4286);
and U7605 (N_7605,N_3216,N_5014);
nor U7606 (N_7606,N_4666,N_3270);
and U7607 (N_7607,N_6063,N_3424);
or U7608 (N_7608,N_5402,N_3891);
nor U7609 (N_7609,N_6009,N_4772);
xor U7610 (N_7610,N_3616,N_3771);
nor U7611 (N_7611,N_4551,N_4431);
xnor U7612 (N_7612,N_4094,N_3176);
xnor U7613 (N_7613,N_3148,N_5937);
nand U7614 (N_7614,N_5737,N_4182);
and U7615 (N_7615,N_3671,N_4809);
nor U7616 (N_7616,N_5435,N_5479);
nor U7617 (N_7617,N_3609,N_3874);
nor U7618 (N_7618,N_5367,N_3202);
nor U7619 (N_7619,N_3985,N_6214);
and U7620 (N_7620,N_5859,N_3929);
and U7621 (N_7621,N_4677,N_5890);
nor U7622 (N_7622,N_5379,N_4769);
nand U7623 (N_7623,N_5382,N_3704);
or U7624 (N_7624,N_3703,N_4498);
or U7625 (N_7625,N_5150,N_6150);
nand U7626 (N_7626,N_3473,N_4729);
and U7627 (N_7627,N_4868,N_4228);
or U7628 (N_7628,N_4928,N_6223);
nand U7629 (N_7629,N_5418,N_4680);
nor U7630 (N_7630,N_3959,N_4497);
nand U7631 (N_7631,N_5552,N_5768);
nor U7632 (N_7632,N_3328,N_3255);
nor U7633 (N_7633,N_5162,N_3624);
nor U7634 (N_7634,N_5172,N_3842);
nand U7635 (N_7635,N_5487,N_3823);
or U7636 (N_7636,N_3323,N_4401);
xnor U7637 (N_7637,N_4594,N_3338);
nand U7638 (N_7638,N_4597,N_5431);
xor U7639 (N_7639,N_3246,N_4811);
xor U7640 (N_7640,N_4144,N_3607);
nor U7641 (N_7641,N_4978,N_3628);
and U7642 (N_7642,N_6090,N_3375);
nand U7643 (N_7643,N_5332,N_3956);
nand U7644 (N_7644,N_5423,N_3555);
and U7645 (N_7645,N_4041,N_4355);
or U7646 (N_7646,N_4670,N_4250);
xor U7647 (N_7647,N_4097,N_3885);
nand U7648 (N_7648,N_3648,N_5797);
and U7649 (N_7649,N_4892,N_5055);
and U7650 (N_7650,N_4648,N_5719);
and U7651 (N_7651,N_3211,N_5081);
or U7652 (N_7652,N_6182,N_3649);
or U7653 (N_7653,N_5845,N_3398);
nand U7654 (N_7654,N_5880,N_4009);
and U7655 (N_7655,N_3302,N_4857);
and U7656 (N_7656,N_5744,N_5237);
nor U7657 (N_7657,N_3652,N_6095);
xnor U7658 (N_7658,N_5444,N_5153);
nor U7659 (N_7659,N_5000,N_4234);
nand U7660 (N_7660,N_5897,N_3897);
xnor U7661 (N_7661,N_5748,N_3907);
xor U7662 (N_7662,N_5540,N_5638);
xnor U7663 (N_7663,N_3795,N_5847);
nor U7664 (N_7664,N_5972,N_4436);
or U7665 (N_7665,N_4359,N_4466);
or U7666 (N_7666,N_5059,N_3465);
and U7667 (N_7667,N_5980,N_6232);
nor U7668 (N_7668,N_5517,N_3200);
nand U7669 (N_7669,N_4031,N_3446);
or U7670 (N_7670,N_6028,N_3808);
and U7671 (N_7671,N_6051,N_4923);
nor U7672 (N_7672,N_3958,N_3396);
nor U7673 (N_7673,N_4343,N_4120);
nor U7674 (N_7674,N_3437,N_4300);
xor U7675 (N_7675,N_4728,N_3256);
and U7676 (N_7676,N_3813,N_3663);
or U7677 (N_7677,N_6163,N_5722);
nand U7678 (N_7678,N_5677,N_5099);
or U7679 (N_7679,N_5463,N_4231);
and U7680 (N_7680,N_4296,N_3327);
nor U7681 (N_7681,N_3753,N_6134);
and U7682 (N_7682,N_4399,N_5496);
nand U7683 (N_7683,N_3731,N_5491);
nor U7684 (N_7684,N_4098,N_5219);
and U7685 (N_7685,N_6186,N_5707);
nand U7686 (N_7686,N_3166,N_5509);
or U7687 (N_7687,N_5533,N_6122);
nor U7688 (N_7688,N_5949,N_5851);
or U7689 (N_7689,N_5142,N_4460);
nor U7690 (N_7690,N_4239,N_5453);
nor U7691 (N_7691,N_5308,N_4415);
and U7692 (N_7692,N_3685,N_4223);
and U7693 (N_7693,N_5270,N_4527);
nand U7694 (N_7694,N_5549,N_4812);
or U7695 (N_7695,N_5473,N_5681);
nor U7696 (N_7696,N_3612,N_5782);
nor U7697 (N_7697,N_5329,N_4012);
nor U7698 (N_7698,N_5870,N_5471);
or U7699 (N_7699,N_3882,N_3643);
nand U7700 (N_7700,N_3674,N_5908);
or U7701 (N_7701,N_4867,N_5011);
xnor U7702 (N_7702,N_3940,N_4490);
and U7703 (N_7703,N_5857,N_3847);
or U7704 (N_7704,N_5935,N_3928);
and U7705 (N_7705,N_5613,N_3599);
nor U7706 (N_7706,N_3654,N_3315);
or U7707 (N_7707,N_3520,N_3992);
nor U7708 (N_7708,N_5041,N_4783);
and U7709 (N_7709,N_6160,N_4080);
or U7710 (N_7710,N_3457,N_5660);
or U7711 (N_7711,N_4159,N_3433);
nand U7712 (N_7712,N_4633,N_4784);
nand U7713 (N_7713,N_4766,N_4232);
nand U7714 (N_7714,N_4380,N_5773);
and U7715 (N_7715,N_5256,N_6113);
and U7716 (N_7716,N_3522,N_4883);
nand U7717 (N_7717,N_5971,N_5534);
and U7718 (N_7718,N_4273,N_5842);
nor U7719 (N_7719,N_4581,N_3626);
xor U7720 (N_7720,N_4655,N_5816);
or U7721 (N_7721,N_5045,N_4416);
nor U7722 (N_7722,N_5648,N_5211);
and U7723 (N_7723,N_3356,N_5307);
or U7724 (N_7724,N_5350,N_6033);
nand U7725 (N_7725,N_5072,N_4854);
or U7726 (N_7726,N_5146,N_5383);
or U7727 (N_7727,N_5076,N_5344);
xor U7728 (N_7728,N_5820,N_5802);
nor U7729 (N_7729,N_6246,N_4748);
and U7730 (N_7730,N_3713,N_4199);
and U7731 (N_7731,N_4804,N_6235);
nand U7732 (N_7732,N_5101,N_4924);
and U7733 (N_7733,N_5273,N_3524);
and U7734 (N_7734,N_4422,N_5316);
nor U7735 (N_7735,N_4901,N_5701);
or U7736 (N_7736,N_5697,N_3331);
xor U7737 (N_7737,N_3849,N_4743);
xnor U7738 (N_7738,N_4765,N_3463);
nand U7739 (N_7739,N_3982,N_3250);
or U7740 (N_7740,N_3403,N_3455);
and U7741 (N_7741,N_6137,N_3272);
or U7742 (N_7742,N_5922,N_3793);
nand U7743 (N_7743,N_3608,N_4195);
and U7744 (N_7744,N_3292,N_3365);
nand U7745 (N_7745,N_6173,N_4532);
nand U7746 (N_7746,N_3318,N_3239);
and U7747 (N_7747,N_3785,N_3576);
nand U7748 (N_7748,N_5717,N_4898);
xnor U7749 (N_7749,N_3355,N_3423);
and U7750 (N_7750,N_5204,N_4631);
or U7751 (N_7751,N_5597,N_4252);
or U7752 (N_7752,N_3311,N_3683);
and U7753 (N_7753,N_4056,N_3802);
nand U7754 (N_7754,N_3633,N_3527);
nand U7755 (N_7755,N_4377,N_4667);
nand U7756 (N_7756,N_5260,N_5129);
nor U7757 (N_7757,N_5283,N_4650);
nor U7758 (N_7758,N_5999,N_5186);
nand U7759 (N_7759,N_4561,N_4799);
nor U7760 (N_7760,N_6102,N_5198);
nor U7761 (N_7761,N_5065,N_5240);
nor U7762 (N_7762,N_3210,N_3401);
nor U7763 (N_7763,N_6088,N_3646);
nand U7764 (N_7764,N_5829,N_6023);
nand U7765 (N_7765,N_3214,N_4172);
nand U7766 (N_7766,N_3440,N_5151);
nor U7767 (N_7767,N_4707,N_4615);
nor U7768 (N_7768,N_3792,N_3232);
or U7769 (N_7769,N_5337,N_6219);
xor U7770 (N_7770,N_5272,N_5144);
xnor U7771 (N_7771,N_3146,N_3392);
and U7772 (N_7772,N_3716,N_4877);
nand U7773 (N_7773,N_5309,N_6060);
nand U7774 (N_7774,N_4240,N_4464);
or U7775 (N_7775,N_4161,N_5541);
nand U7776 (N_7776,N_4971,N_4396);
nor U7777 (N_7777,N_3225,N_6119);
and U7778 (N_7778,N_4582,N_4280);
and U7779 (N_7779,N_5413,N_3641);
nor U7780 (N_7780,N_5416,N_4384);
xor U7781 (N_7781,N_4846,N_4656);
or U7782 (N_7782,N_5504,N_3358);
and U7783 (N_7783,N_3517,N_4731);
nor U7784 (N_7784,N_5891,N_3226);
nor U7785 (N_7785,N_4103,N_5373);
or U7786 (N_7786,N_4168,N_4775);
xor U7787 (N_7787,N_5419,N_5067);
nand U7788 (N_7788,N_4381,N_4782);
nand U7789 (N_7789,N_5060,N_4501);
nor U7790 (N_7790,N_3425,N_3860);
or U7791 (N_7791,N_4424,N_4169);
or U7792 (N_7792,N_4718,N_3139);
nand U7793 (N_7793,N_5884,N_4940);
nand U7794 (N_7794,N_3948,N_5893);
nor U7795 (N_7795,N_3697,N_3317);
or U7796 (N_7796,N_4856,N_4037);
xnor U7797 (N_7797,N_5074,N_5358);
nor U7798 (N_7798,N_3613,N_4573);
nand U7799 (N_7799,N_6170,N_3883);
nand U7800 (N_7800,N_6202,N_5364);
and U7801 (N_7801,N_5807,N_5506);
nand U7802 (N_7802,N_5098,N_5152);
or U7803 (N_7803,N_3580,N_3636);
and U7804 (N_7804,N_5154,N_5653);
nor U7805 (N_7805,N_4912,N_3767);
and U7806 (N_7806,N_5938,N_5585);
xor U7807 (N_7807,N_5827,N_3780);
nand U7808 (N_7808,N_5053,N_5145);
or U7809 (N_7809,N_3921,N_4719);
nand U7810 (N_7810,N_4290,N_4302);
nor U7811 (N_7811,N_4261,N_3591);
or U7812 (N_7812,N_5173,N_5404);
or U7813 (N_7813,N_4998,N_5225);
or U7814 (N_7814,N_6011,N_6234);
nor U7815 (N_7815,N_5465,N_3323);
or U7816 (N_7816,N_5054,N_4667);
nand U7817 (N_7817,N_4649,N_5116);
nor U7818 (N_7818,N_5417,N_5813);
nand U7819 (N_7819,N_5927,N_5856);
and U7820 (N_7820,N_3732,N_3826);
nor U7821 (N_7821,N_5878,N_5131);
nand U7822 (N_7822,N_3727,N_4697);
and U7823 (N_7823,N_4967,N_5905);
nor U7824 (N_7824,N_3996,N_4592);
nor U7825 (N_7825,N_4492,N_4464);
or U7826 (N_7826,N_3476,N_3175);
or U7827 (N_7827,N_3723,N_3976);
and U7828 (N_7828,N_5722,N_3260);
xnor U7829 (N_7829,N_6214,N_3539);
xnor U7830 (N_7830,N_4599,N_5323);
and U7831 (N_7831,N_4422,N_4048);
and U7832 (N_7832,N_3177,N_5661);
or U7833 (N_7833,N_3963,N_5949);
or U7834 (N_7834,N_5879,N_3389);
xor U7835 (N_7835,N_4816,N_6229);
nand U7836 (N_7836,N_3256,N_3844);
nor U7837 (N_7837,N_3982,N_5899);
and U7838 (N_7838,N_4866,N_4019);
nand U7839 (N_7839,N_5678,N_4089);
and U7840 (N_7840,N_4011,N_5995);
or U7841 (N_7841,N_5140,N_4399);
or U7842 (N_7842,N_4967,N_3622);
and U7843 (N_7843,N_4563,N_5885);
or U7844 (N_7844,N_3821,N_5049);
or U7845 (N_7845,N_4060,N_5956);
or U7846 (N_7846,N_5294,N_4746);
and U7847 (N_7847,N_5567,N_4515);
and U7848 (N_7848,N_4329,N_4351);
or U7849 (N_7849,N_5079,N_4930);
nor U7850 (N_7850,N_5077,N_5643);
nand U7851 (N_7851,N_3883,N_4705);
nand U7852 (N_7852,N_5366,N_4564);
xor U7853 (N_7853,N_6157,N_5154);
or U7854 (N_7854,N_5627,N_5701);
nor U7855 (N_7855,N_3976,N_4900);
nor U7856 (N_7856,N_5353,N_3139);
or U7857 (N_7857,N_6235,N_5130);
and U7858 (N_7858,N_3800,N_5800);
nand U7859 (N_7859,N_6193,N_3305);
nand U7860 (N_7860,N_5269,N_6112);
nand U7861 (N_7861,N_5252,N_4351);
nor U7862 (N_7862,N_4308,N_3453);
nand U7863 (N_7863,N_3944,N_5959);
and U7864 (N_7864,N_5673,N_6173);
nand U7865 (N_7865,N_6057,N_4070);
or U7866 (N_7866,N_5072,N_5407);
and U7867 (N_7867,N_3838,N_5697);
and U7868 (N_7868,N_5896,N_5333);
nor U7869 (N_7869,N_3507,N_3863);
nor U7870 (N_7870,N_5184,N_5249);
and U7871 (N_7871,N_4764,N_5208);
and U7872 (N_7872,N_3967,N_5061);
and U7873 (N_7873,N_5006,N_6050);
or U7874 (N_7874,N_5191,N_4636);
nor U7875 (N_7875,N_4604,N_5322);
and U7876 (N_7876,N_4077,N_4529);
nor U7877 (N_7877,N_4410,N_3546);
or U7878 (N_7878,N_3274,N_3348);
nor U7879 (N_7879,N_4429,N_3490);
nand U7880 (N_7880,N_4544,N_5320);
or U7881 (N_7881,N_4687,N_4543);
nand U7882 (N_7882,N_4357,N_5968);
nand U7883 (N_7883,N_5401,N_3361);
nor U7884 (N_7884,N_3176,N_3125);
xor U7885 (N_7885,N_3371,N_3421);
nand U7886 (N_7886,N_4113,N_6139);
nand U7887 (N_7887,N_5778,N_4158);
and U7888 (N_7888,N_5304,N_4593);
nor U7889 (N_7889,N_4774,N_3291);
nor U7890 (N_7890,N_4948,N_5909);
nor U7891 (N_7891,N_6154,N_5459);
nor U7892 (N_7892,N_4674,N_4609);
or U7893 (N_7893,N_3885,N_5308);
and U7894 (N_7894,N_4537,N_4337);
or U7895 (N_7895,N_3268,N_5765);
and U7896 (N_7896,N_6161,N_4250);
nor U7897 (N_7897,N_5287,N_3181);
and U7898 (N_7898,N_4492,N_5560);
nand U7899 (N_7899,N_5437,N_5708);
and U7900 (N_7900,N_4215,N_3647);
nor U7901 (N_7901,N_4704,N_5083);
nor U7902 (N_7902,N_3592,N_4488);
nor U7903 (N_7903,N_4867,N_4880);
nor U7904 (N_7904,N_5337,N_5017);
or U7905 (N_7905,N_6199,N_3754);
or U7906 (N_7906,N_5864,N_3760);
or U7907 (N_7907,N_4860,N_4837);
or U7908 (N_7908,N_4449,N_4331);
nand U7909 (N_7909,N_5290,N_5215);
or U7910 (N_7910,N_4405,N_4472);
or U7911 (N_7911,N_5974,N_6131);
nor U7912 (N_7912,N_5997,N_5456);
nand U7913 (N_7913,N_4291,N_5191);
nand U7914 (N_7914,N_3965,N_4588);
and U7915 (N_7915,N_3310,N_3856);
nor U7916 (N_7916,N_3386,N_5422);
nand U7917 (N_7917,N_5408,N_5126);
or U7918 (N_7918,N_4557,N_6039);
nand U7919 (N_7919,N_3444,N_5839);
or U7920 (N_7920,N_4338,N_5081);
or U7921 (N_7921,N_5857,N_4954);
nand U7922 (N_7922,N_5136,N_3950);
nand U7923 (N_7923,N_4315,N_4878);
and U7924 (N_7924,N_5905,N_5290);
nor U7925 (N_7925,N_5395,N_5344);
or U7926 (N_7926,N_5781,N_3553);
nor U7927 (N_7927,N_4053,N_5562);
nor U7928 (N_7928,N_5158,N_4945);
or U7929 (N_7929,N_4564,N_4629);
nor U7930 (N_7930,N_4696,N_5679);
nand U7931 (N_7931,N_4908,N_3909);
nand U7932 (N_7932,N_3738,N_3185);
or U7933 (N_7933,N_3754,N_6040);
and U7934 (N_7934,N_3727,N_4943);
and U7935 (N_7935,N_5191,N_4281);
nor U7936 (N_7936,N_4710,N_6188);
and U7937 (N_7937,N_4066,N_3725);
xnor U7938 (N_7938,N_4481,N_3489);
or U7939 (N_7939,N_6106,N_4436);
xor U7940 (N_7940,N_3966,N_5933);
and U7941 (N_7941,N_4701,N_6242);
and U7942 (N_7942,N_5541,N_5197);
or U7943 (N_7943,N_4486,N_3687);
nand U7944 (N_7944,N_5513,N_3445);
nand U7945 (N_7945,N_4979,N_4932);
nand U7946 (N_7946,N_4224,N_4239);
or U7947 (N_7947,N_5904,N_3903);
xor U7948 (N_7948,N_5618,N_4058);
xor U7949 (N_7949,N_5873,N_5348);
or U7950 (N_7950,N_6000,N_5298);
and U7951 (N_7951,N_4134,N_5945);
nor U7952 (N_7952,N_3213,N_5770);
and U7953 (N_7953,N_6091,N_4622);
or U7954 (N_7954,N_6195,N_5322);
or U7955 (N_7955,N_3289,N_4736);
and U7956 (N_7956,N_4893,N_4982);
nand U7957 (N_7957,N_5164,N_3301);
nand U7958 (N_7958,N_3543,N_4823);
or U7959 (N_7959,N_6215,N_5697);
or U7960 (N_7960,N_4894,N_5605);
xor U7961 (N_7961,N_3318,N_4639);
nor U7962 (N_7962,N_4146,N_4577);
xor U7963 (N_7963,N_5830,N_3851);
and U7964 (N_7964,N_3973,N_4529);
or U7965 (N_7965,N_4419,N_4894);
and U7966 (N_7966,N_4824,N_4342);
nand U7967 (N_7967,N_4045,N_4788);
xnor U7968 (N_7968,N_3809,N_3153);
or U7969 (N_7969,N_4139,N_5877);
or U7970 (N_7970,N_4520,N_3155);
nand U7971 (N_7971,N_3315,N_4618);
and U7972 (N_7972,N_3490,N_5388);
and U7973 (N_7973,N_4533,N_4065);
nor U7974 (N_7974,N_5362,N_5917);
nor U7975 (N_7975,N_4311,N_6120);
nor U7976 (N_7976,N_5732,N_3561);
and U7977 (N_7977,N_5306,N_3599);
nand U7978 (N_7978,N_4657,N_4467);
and U7979 (N_7979,N_5306,N_5447);
nor U7980 (N_7980,N_3819,N_4459);
and U7981 (N_7981,N_4363,N_4246);
or U7982 (N_7982,N_4679,N_4572);
and U7983 (N_7983,N_4434,N_4056);
nand U7984 (N_7984,N_4940,N_5033);
nand U7985 (N_7985,N_4682,N_6067);
nor U7986 (N_7986,N_5622,N_3864);
nand U7987 (N_7987,N_5831,N_4313);
and U7988 (N_7988,N_5237,N_3941);
or U7989 (N_7989,N_5044,N_3840);
or U7990 (N_7990,N_6222,N_5917);
and U7991 (N_7991,N_5667,N_4737);
and U7992 (N_7992,N_3646,N_5784);
and U7993 (N_7993,N_4800,N_5639);
or U7994 (N_7994,N_4407,N_4770);
nor U7995 (N_7995,N_5000,N_5751);
nor U7996 (N_7996,N_5153,N_6141);
nand U7997 (N_7997,N_6102,N_5571);
nand U7998 (N_7998,N_4907,N_5199);
xor U7999 (N_7999,N_6120,N_3133);
or U8000 (N_8000,N_3193,N_5939);
or U8001 (N_8001,N_5525,N_5510);
or U8002 (N_8002,N_5836,N_3151);
or U8003 (N_8003,N_3770,N_5410);
and U8004 (N_8004,N_4481,N_4990);
nand U8005 (N_8005,N_4476,N_5432);
xnor U8006 (N_8006,N_5747,N_3993);
or U8007 (N_8007,N_3695,N_5517);
nand U8008 (N_8008,N_3144,N_3524);
and U8009 (N_8009,N_5560,N_5745);
or U8010 (N_8010,N_4061,N_3357);
nand U8011 (N_8011,N_3672,N_3919);
or U8012 (N_8012,N_4243,N_4620);
and U8013 (N_8013,N_4630,N_5003);
nor U8014 (N_8014,N_6003,N_4558);
xnor U8015 (N_8015,N_4745,N_3238);
xor U8016 (N_8016,N_5830,N_4223);
or U8017 (N_8017,N_5441,N_3790);
nand U8018 (N_8018,N_3426,N_6089);
nand U8019 (N_8019,N_4573,N_5113);
or U8020 (N_8020,N_5381,N_3620);
or U8021 (N_8021,N_4662,N_5163);
nor U8022 (N_8022,N_4335,N_4719);
nor U8023 (N_8023,N_3895,N_5905);
nor U8024 (N_8024,N_4843,N_5922);
nor U8025 (N_8025,N_3885,N_5262);
and U8026 (N_8026,N_3519,N_3723);
nand U8027 (N_8027,N_3491,N_3940);
or U8028 (N_8028,N_5367,N_5809);
and U8029 (N_8029,N_5919,N_6247);
and U8030 (N_8030,N_5511,N_5538);
or U8031 (N_8031,N_3269,N_4801);
nor U8032 (N_8032,N_5911,N_3213);
or U8033 (N_8033,N_4387,N_3196);
or U8034 (N_8034,N_4796,N_4357);
nand U8035 (N_8035,N_4202,N_5938);
xor U8036 (N_8036,N_5141,N_4273);
xnor U8037 (N_8037,N_5681,N_5464);
and U8038 (N_8038,N_3355,N_4237);
xor U8039 (N_8039,N_5645,N_4493);
nor U8040 (N_8040,N_3499,N_3515);
nand U8041 (N_8041,N_5928,N_6245);
nor U8042 (N_8042,N_3312,N_5526);
xor U8043 (N_8043,N_5766,N_4217);
and U8044 (N_8044,N_4888,N_3274);
and U8045 (N_8045,N_6185,N_4832);
nand U8046 (N_8046,N_5703,N_5046);
nor U8047 (N_8047,N_4269,N_3755);
or U8048 (N_8048,N_4453,N_5998);
xnor U8049 (N_8049,N_5999,N_4054);
and U8050 (N_8050,N_3812,N_5914);
xnor U8051 (N_8051,N_4347,N_5426);
and U8052 (N_8052,N_4132,N_4709);
or U8053 (N_8053,N_5795,N_5168);
nand U8054 (N_8054,N_4287,N_3717);
or U8055 (N_8055,N_4522,N_6200);
or U8056 (N_8056,N_5049,N_4264);
nor U8057 (N_8057,N_5798,N_5573);
and U8058 (N_8058,N_4373,N_3338);
and U8059 (N_8059,N_4522,N_4933);
nor U8060 (N_8060,N_5210,N_4113);
and U8061 (N_8061,N_4007,N_5549);
xnor U8062 (N_8062,N_5418,N_3672);
or U8063 (N_8063,N_5909,N_4044);
or U8064 (N_8064,N_3876,N_5605);
and U8065 (N_8065,N_3176,N_5893);
or U8066 (N_8066,N_5284,N_4713);
nand U8067 (N_8067,N_3495,N_4604);
nor U8068 (N_8068,N_4895,N_3998);
nand U8069 (N_8069,N_5190,N_5078);
or U8070 (N_8070,N_3728,N_4040);
or U8071 (N_8071,N_3393,N_5464);
nor U8072 (N_8072,N_4748,N_5321);
and U8073 (N_8073,N_3593,N_3442);
or U8074 (N_8074,N_3429,N_3932);
nand U8075 (N_8075,N_5510,N_5402);
and U8076 (N_8076,N_4367,N_5530);
nand U8077 (N_8077,N_4399,N_5954);
xor U8078 (N_8078,N_5957,N_3849);
nor U8079 (N_8079,N_4780,N_6235);
and U8080 (N_8080,N_5575,N_4538);
or U8081 (N_8081,N_3947,N_4455);
nand U8082 (N_8082,N_5939,N_4286);
and U8083 (N_8083,N_3268,N_5228);
nand U8084 (N_8084,N_4835,N_3771);
nand U8085 (N_8085,N_3267,N_5830);
and U8086 (N_8086,N_4698,N_4451);
and U8087 (N_8087,N_3530,N_5397);
or U8088 (N_8088,N_4397,N_3543);
nor U8089 (N_8089,N_5985,N_5211);
and U8090 (N_8090,N_3685,N_3287);
and U8091 (N_8091,N_3951,N_4985);
or U8092 (N_8092,N_4836,N_4801);
or U8093 (N_8093,N_5576,N_4709);
nor U8094 (N_8094,N_5013,N_5959);
nor U8095 (N_8095,N_4778,N_4234);
nor U8096 (N_8096,N_4760,N_3575);
nor U8097 (N_8097,N_3259,N_3423);
or U8098 (N_8098,N_5550,N_4500);
xnor U8099 (N_8099,N_5134,N_4077);
or U8100 (N_8100,N_4116,N_3751);
or U8101 (N_8101,N_4847,N_4549);
and U8102 (N_8102,N_3235,N_4071);
nand U8103 (N_8103,N_4524,N_4027);
or U8104 (N_8104,N_5921,N_4841);
xor U8105 (N_8105,N_4183,N_3216);
nand U8106 (N_8106,N_3655,N_5507);
nand U8107 (N_8107,N_4751,N_3363);
and U8108 (N_8108,N_4069,N_5548);
and U8109 (N_8109,N_3505,N_5222);
or U8110 (N_8110,N_3756,N_6038);
nor U8111 (N_8111,N_3697,N_6121);
nand U8112 (N_8112,N_4660,N_4279);
and U8113 (N_8113,N_3481,N_3494);
xor U8114 (N_8114,N_3747,N_6165);
nor U8115 (N_8115,N_5011,N_5987);
or U8116 (N_8116,N_4733,N_4367);
xnor U8117 (N_8117,N_4326,N_5266);
and U8118 (N_8118,N_3847,N_6068);
and U8119 (N_8119,N_4830,N_3949);
and U8120 (N_8120,N_3920,N_3198);
or U8121 (N_8121,N_4562,N_4391);
nand U8122 (N_8122,N_5060,N_5507);
and U8123 (N_8123,N_4366,N_4268);
nand U8124 (N_8124,N_3621,N_5914);
xor U8125 (N_8125,N_6175,N_6037);
and U8126 (N_8126,N_3986,N_6240);
nand U8127 (N_8127,N_5164,N_4899);
or U8128 (N_8128,N_4106,N_4762);
and U8129 (N_8129,N_4197,N_5890);
and U8130 (N_8130,N_5917,N_5593);
nand U8131 (N_8131,N_6144,N_6135);
xnor U8132 (N_8132,N_6072,N_4867);
or U8133 (N_8133,N_4585,N_5877);
or U8134 (N_8134,N_5173,N_4423);
nand U8135 (N_8135,N_5973,N_5162);
nand U8136 (N_8136,N_4792,N_5994);
or U8137 (N_8137,N_5791,N_4184);
and U8138 (N_8138,N_3692,N_4142);
and U8139 (N_8139,N_4722,N_3540);
and U8140 (N_8140,N_3705,N_3201);
or U8141 (N_8141,N_4149,N_4977);
and U8142 (N_8142,N_3831,N_4936);
nand U8143 (N_8143,N_5433,N_4860);
and U8144 (N_8144,N_5324,N_4309);
nor U8145 (N_8145,N_5464,N_5016);
nor U8146 (N_8146,N_5550,N_3961);
nand U8147 (N_8147,N_3973,N_5145);
or U8148 (N_8148,N_4331,N_3579);
and U8149 (N_8149,N_5525,N_4691);
and U8150 (N_8150,N_5789,N_3336);
nand U8151 (N_8151,N_3367,N_6159);
and U8152 (N_8152,N_3738,N_3542);
and U8153 (N_8153,N_3562,N_3754);
and U8154 (N_8154,N_5683,N_4546);
nand U8155 (N_8155,N_4926,N_3980);
and U8156 (N_8156,N_3880,N_5588);
or U8157 (N_8157,N_5555,N_4655);
or U8158 (N_8158,N_5772,N_5404);
nor U8159 (N_8159,N_5006,N_4331);
nor U8160 (N_8160,N_5527,N_4855);
and U8161 (N_8161,N_4738,N_5857);
nand U8162 (N_8162,N_5384,N_3598);
nand U8163 (N_8163,N_5938,N_5741);
nand U8164 (N_8164,N_4466,N_5176);
nor U8165 (N_8165,N_5814,N_5477);
nand U8166 (N_8166,N_5633,N_4220);
or U8167 (N_8167,N_3412,N_3676);
and U8168 (N_8168,N_3943,N_5942);
or U8169 (N_8169,N_4410,N_3932);
nand U8170 (N_8170,N_5235,N_4352);
xnor U8171 (N_8171,N_3977,N_4463);
nor U8172 (N_8172,N_4899,N_5272);
xor U8173 (N_8173,N_4988,N_6238);
nor U8174 (N_8174,N_5013,N_5000);
and U8175 (N_8175,N_5794,N_3217);
nand U8176 (N_8176,N_4248,N_5487);
nand U8177 (N_8177,N_3691,N_4546);
and U8178 (N_8178,N_4067,N_4986);
or U8179 (N_8179,N_3244,N_5552);
or U8180 (N_8180,N_5588,N_4345);
nand U8181 (N_8181,N_3200,N_4236);
nor U8182 (N_8182,N_4284,N_4035);
nand U8183 (N_8183,N_3430,N_3992);
or U8184 (N_8184,N_3295,N_5825);
nor U8185 (N_8185,N_4962,N_6115);
and U8186 (N_8186,N_3778,N_3944);
and U8187 (N_8187,N_5291,N_3304);
nor U8188 (N_8188,N_4632,N_4062);
or U8189 (N_8189,N_3557,N_3502);
nand U8190 (N_8190,N_4203,N_4279);
nand U8191 (N_8191,N_3779,N_3569);
and U8192 (N_8192,N_3176,N_4929);
and U8193 (N_8193,N_5231,N_5122);
nor U8194 (N_8194,N_4952,N_4490);
or U8195 (N_8195,N_4455,N_4544);
nand U8196 (N_8196,N_4642,N_3252);
or U8197 (N_8197,N_4755,N_3632);
or U8198 (N_8198,N_6009,N_3872);
xnor U8199 (N_8199,N_3797,N_5234);
and U8200 (N_8200,N_4850,N_5774);
and U8201 (N_8201,N_4741,N_5783);
and U8202 (N_8202,N_4166,N_5752);
nor U8203 (N_8203,N_3538,N_4149);
xnor U8204 (N_8204,N_3133,N_5728);
or U8205 (N_8205,N_5966,N_5653);
nand U8206 (N_8206,N_3600,N_5986);
xor U8207 (N_8207,N_4433,N_4006);
xnor U8208 (N_8208,N_3222,N_5422);
nand U8209 (N_8209,N_3392,N_5795);
or U8210 (N_8210,N_4791,N_4253);
and U8211 (N_8211,N_4189,N_4596);
or U8212 (N_8212,N_5431,N_3556);
and U8213 (N_8213,N_5642,N_3215);
nor U8214 (N_8214,N_5991,N_5864);
nor U8215 (N_8215,N_5145,N_4122);
nor U8216 (N_8216,N_5655,N_4500);
or U8217 (N_8217,N_4689,N_4139);
nand U8218 (N_8218,N_3443,N_5323);
and U8219 (N_8219,N_3130,N_4033);
nand U8220 (N_8220,N_3874,N_5442);
xnor U8221 (N_8221,N_5146,N_4041);
and U8222 (N_8222,N_5553,N_5976);
and U8223 (N_8223,N_3506,N_5714);
nor U8224 (N_8224,N_4718,N_3660);
nand U8225 (N_8225,N_4493,N_4610);
nand U8226 (N_8226,N_5540,N_3958);
nand U8227 (N_8227,N_3763,N_3951);
nor U8228 (N_8228,N_4294,N_5164);
nand U8229 (N_8229,N_3575,N_4182);
nor U8230 (N_8230,N_6239,N_5217);
or U8231 (N_8231,N_5793,N_4181);
nand U8232 (N_8232,N_6163,N_5892);
nor U8233 (N_8233,N_4313,N_3865);
and U8234 (N_8234,N_6209,N_3682);
xor U8235 (N_8235,N_6095,N_5653);
nor U8236 (N_8236,N_3286,N_3546);
nor U8237 (N_8237,N_6144,N_4606);
and U8238 (N_8238,N_4681,N_5676);
nor U8239 (N_8239,N_3437,N_5369);
nand U8240 (N_8240,N_3658,N_3996);
and U8241 (N_8241,N_5516,N_5378);
nor U8242 (N_8242,N_4343,N_5523);
and U8243 (N_8243,N_4445,N_5860);
nand U8244 (N_8244,N_4050,N_4898);
nor U8245 (N_8245,N_4179,N_5537);
nand U8246 (N_8246,N_5194,N_3717);
xnor U8247 (N_8247,N_4812,N_5195);
and U8248 (N_8248,N_4089,N_6143);
nand U8249 (N_8249,N_3155,N_3982);
nor U8250 (N_8250,N_3683,N_5692);
and U8251 (N_8251,N_3944,N_4853);
nor U8252 (N_8252,N_4909,N_3528);
nand U8253 (N_8253,N_5720,N_5261);
or U8254 (N_8254,N_4692,N_3246);
or U8255 (N_8255,N_3427,N_5762);
nand U8256 (N_8256,N_4028,N_3882);
or U8257 (N_8257,N_4331,N_5527);
nand U8258 (N_8258,N_4585,N_3363);
and U8259 (N_8259,N_6078,N_3650);
and U8260 (N_8260,N_3904,N_4191);
and U8261 (N_8261,N_4851,N_3260);
xor U8262 (N_8262,N_3687,N_4187);
nor U8263 (N_8263,N_3288,N_5511);
or U8264 (N_8264,N_5163,N_5335);
or U8265 (N_8265,N_4028,N_5474);
or U8266 (N_8266,N_5597,N_5120);
nor U8267 (N_8267,N_6140,N_5199);
nor U8268 (N_8268,N_4237,N_3221);
or U8269 (N_8269,N_3973,N_5828);
nor U8270 (N_8270,N_5395,N_6249);
nand U8271 (N_8271,N_5273,N_3755);
or U8272 (N_8272,N_5778,N_3817);
nand U8273 (N_8273,N_4635,N_3420);
and U8274 (N_8274,N_5717,N_4238);
nand U8275 (N_8275,N_4951,N_3958);
and U8276 (N_8276,N_4869,N_6078);
xor U8277 (N_8277,N_4385,N_4736);
nand U8278 (N_8278,N_4226,N_3425);
nand U8279 (N_8279,N_6188,N_5586);
or U8280 (N_8280,N_4760,N_4576);
nand U8281 (N_8281,N_4454,N_5657);
and U8282 (N_8282,N_4635,N_5403);
nand U8283 (N_8283,N_5933,N_5112);
nand U8284 (N_8284,N_6136,N_3431);
nor U8285 (N_8285,N_3203,N_4104);
nand U8286 (N_8286,N_3628,N_5702);
xnor U8287 (N_8287,N_5221,N_3484);
nand U8288 (N_8288,N_4763,N_3934);
nand U8289 (N_8289,N_5412,N_4819);
nor U8290 (N_8290,N_3431,N_5389);
or U8291 (N_8291,N_4304,N_3481);
xor U8292 (N_8292,N_3831,N_4714);
nor U8293 (N_8293,N_5053,N_5897);
and U8294 (N_8294,N_4407,N_3215);
or U8295 (N_8295,N_5023,N_3817);
nor U8296 (N_8296,N_5010,N_3245);
nand U8297 (N_8297,N_3805,N_5544);
nor U8298 (N_8298,N_5248,N_4559);
and U8299 (N_8299,N_5122,N_3479);
nor U8300 (N_8300,N_5669,N_3546);
nand U8301 (N_8301,N_5228,N_5805);
nand U8302 (N_8302,N_6101,N_4272);
nand U8303 (N_8303,N_4310,N_3659);
nand U8304 (N_8304,N_5247,N_5354);
nand U8305 (N_8305,N_6089,N_4112);
or U8306 (N_8306,N_3366,N_3747);
xor U8307 (N_8307,N_3210,N_5650);
or U8308 (N_8308,N_5468,N_4207);
or U8309 (N_8309,N_4199,N_4135);
nand U8310 (N_8310,N_4540,N_5629);
nor U8311 (N_8311,N_5889,N_5671);
and U8312 (N_8312,N_5765,N_5979);
and U8313 (N_8313,N_4495,N_5655);
nor U8314 (N_8314,N_3443,N_5228);
or U8315 (N_8315,N_4380,N_4889);
or U8316 (N_8316,N_5984,N_4937);
or U8317 (N_8317,N_3386,N_5932);
and U8318 (N_8318,N_4915,N_6236);
xnor U8319 (N_8319,N_3735,N_5672);
and U8320 (N_8320,N_5000,N_5466);
and U8321 (N_8321,N_4118,N_4164);
nor U8322 (N_8322,N_3173,N_4957);
xnor U8323 (N_8323,N_3382,N_5669);
and U8324 (N_8324,N_4869,N_5908);
or U8325 (N_8325,N_3157,N_5726);
nand U8326 (N_8326,N_3971,N_4079);
and U8327 (N_8327,N_3679,N_6137);
and U8328 (N_8328,N_4557,N_6038);
nor U8329 (N_8329,N_5839,N_5146);
nor U8330 (N_8330,N_3874,N_4172);
nand U8331 (N_8331,N_3269,N_5061);
and U8332 (N_8332,N_5956,N_5937);
nor U8333 (N_8333,N_3461,N_4508);
nand U8334 (N_8334,N_3528,N_5547);
xnor U8335 (N_8335,N_4153,N_4621);
nor U8336 (N_8336,N_5281,N_4652);
nand U8337 (N_8337,N_3793,N_5072);
xor U8338 (N_8338,N_5615,N_4521);
nor U8339 (N_8339,N_5772,N_6096);
nor U8340 (N_8340,N_4242,N_4891);
nand U8341 (N_8341,N_3408,N_3151);
nor U8342 (N_8342,N_4868,N_3672);
nand U8343 (N_8343,N_3232,N_4424);
and U8344 (N_8344,N_5451,N_3397);
or U8345 (N_8345,N_5445,N_5098);
or U8346 (N_8346,N_5390,N_3995);
or U8347 (N_8347,N_4860,N_4387);
or U8348 (N_8348,N_3522,N_5614);
xor U8349 (N_8349,N_5505,N_3913);
or U8350 (N_8350,N_3181,N_5449);
nor U8351 (N_8351,N_5950,N_5408);
or U8352 (N_8352,N_3126,N_6239);
and U8353 (N_8353,N_5978,N_3761);
and U8354 (N_8354,N_3537,N_4536);
nand U8355 (N_8355,N_4935,N_5080);
and U8356 (N_8356,N_3988,N_4504);
xor U8357 (N_8357,N_4822,N_4055);
nand U8358 (N_8358,N_5100,N_3545);
or U8359 (N_8359,N_5957,N_4110);
nand U8360 (N_8360,N_5384,N_5470);
nor U8361 (N_8361,N_5266,N_6093);
and U8362 (N_8362,N_5895,N_4970);
or U8363 (N_8363,N_5457,N_6119);
or U8364 (N_8364,N_5360,N_5551);
xnor U8365 (N_8365,N_3605,N_3689);
nand U8366 (N_8366,N_5557,N_4741);
nor U8367 (N_8367,N_5345,N_4892);
and U8368 (N_8368,N_4499,N_5072);
or U8369 (N_8369,N_5605,N_5707);
or U8370 (N_8370,N_5549,N_4756);
nand U8371 (N_8371,N_3722,N_4103);
or U8372 (N_8372,N_3591,N_4857);
xnor U8373 (N_8373,N_5207,N_5669);
and U8374 (N_8374,N_4492,N_3900);
and U8375 (N_8375,N_5873,N_4169);
or U8376 (N_8376,N_3976,N_5441);
or U8377 (N_8377,N_5596,N_5103);
or U8378 (N_8378,N_4310,N_3386);
or U8379 (N_8379,N_3214,N_3196);
nand U8380 (N_8380,N_4550,N_4818);
nand U8381 (N_8381,N_3220,N_5848);
and U8382 (N_8382,N_4263,N_5813);
and U8383 (N_8383,N_5157,N_5769);
or U8384 (N_8384,N_3924,N_4927);
nor U8385 (N_8385,N_6059,N_3256);
nand U8386 (N_8386,N_4590,N_5200);
and U8387 (N_8387,N_5598,N_3404);
or U8388 (N_8388,N_4874,N_4348);
nor U8389 (N_8389,N_5831,N_5118);
and U8390 (N_8390,N_6103,N_3347);
nand U8391 (N_8391,N_5864,N_3528);
xor U8392 (N_8392,N_6177,N_5004);
nand U8393 (N_8393,N_4558,N_3745);
and U8394 (N_8394,N_5188,N_5931);
or U8395 (N_8395,N_4396,N_3305);
or U8396 (N_8396,N_4640,N_3558);
nand U8397 (N_8397,N_3662,N_4592);
nor U8398 (N_8398,N_4186,N_4467);
nor U8399 (N_8399,N_5929,N_4505);
nor U8400 (N_8400,N_4578,N_5482);
xnor U8401 (N_8401,N_6091,N_4173);
nor U8402 (N_8402,N_3193,N_5691);
nor U8403 (N_8403,N_4843,N_4091);
and U8404 (N_8404,N_5252,N_4084);
nand U8405 (N_8405,N_3174,N_5009);
nand U8406 (N_8406,N_4197,N_5082);
nor U8407 (N_8407,N_3169,N_5055);
nand U8408 (N_8408,N_3258,N_5565);
or U8409 (N_8409,N_5004,N_3744);
and U8410 (N_8410,N_6045,N_3886);
or U8411 (N_8411,N_4788,N_5386);
or U8412 (N_8412,N_6245,N_6120);
nand U8413 (N_8413,N_3884,N_4918);
and U8414 (N_8414,N_4568,N_3264);
or U8415 (N_8415,N_6048,N_4456);
or U8416 (N_8416,N_4185,N_3562);
nor U8417 (N_8417,N_3394,N_3443);
and U8418 (N_8418,N_4349,N_5256);
nand U8419 (N_8419,N_4920,N_3660);
or U8420 (N_8420,N_3621,N_4323);
or U8421 (N_8421,N_4507,N_4657);
or U8422 (N_8422,N_5175,N_3856);
nor U8423 (N_8423,N_3834,N_3978);
nor U8424 (N_8424,N_5443,N_4889);
or U8425 (N_8425,N_6100,N_5003);
nor U8426 (N_8426,N_4938,N_5488);
nand U8427 (N_8427,N_3881,N_3837);
or U8428 (N_8428,N_3561,N_3770);
nor U8429 (N_8429,N_4800,N_3982);
nor U8430 (N_8430,N_3423,N_4893);
nor U8431 (N_8431,N_6232,N_5057);
nand U8432 (N_8432,N_3252,N_5986);
and U8433 (N_8433,N_4707,N_3737);
nand U8434 (N_8434,N_5052,N_6020);
nor U8435 (N_8435,N_4705,N_4034);
or U8436 (N_8436,N_3631,N_3461);
or U8437 (N_8437,N_3461,N_4167);
nor U8438 (N_8438,N_4639,N_4848);
or U8439 (N_8439,N_4117,N_3269);
nor U8440 (N_8440,N_4031,N_3302);
nor U8441 (N_8441,N_5957,N_4368);
xor U8442 (N_8442,N_4794,N_3540);
or U8443 (N_8443,N_4127,N_5168);
or U8444 (N_8444,N_3440,N_3279);
xnor U8445 (N_8445,N_4089,N_4037);
or U8446 (N_8446,N_4304,N_3147);
xnor U8447 (N_8447,N_4430,N_5602);
or U8448 (N_8448,N_5733,N_6227);
nor U8449 (N_8449,N_3672,N_5815);
and U8450 (N_8450,N_4138,N_4535);
nor U8451 (N_8451,N_4442,N_5833);
or U8452 (N_8452,N_4378,N_5106);
and U8453 (N_8453,N_5383,N_3465);
xnor U8454 (N_8454,N_4116,N_5489);
nor U8455 (N_8455,N_4174,N_4680);
and U8456 (N_8456,N_4092,N_5994);
or U8457 (N_8457,N_4492,N_3645);
and U8458 (N_8458,N_3635,N_5441);
nand U8459 (N_8459,N_3385,N_5242);
nor U8460 (N_8460,N_4962,N_3224);
nand U8461 (N_8461,N_3427,N_5533);
and U8462 (N_8462,N_5245,N_5515);
nor U8463 (N_8463,N_3416,N_5563);
or U8464 (N_8464,N_3682,N_4693);
and U8465 (N_8465,N_3225,N_5012);
xor U8466 (N_8466,N_5642,N_6209);
nor U8467 (N_8467,N_3185,N_3376);
xor U8468 (N_8468,N_4813,N_5412);
or U8469 (N_8469,N_5257,N_5420);
or U8470 (N_8470,N_3186,N_4082);
nor U8471 (N_8471,N_5090,N_6072);
nor U8472 (N_8472,N_3856,N_3398);
or U8473 (N_8473,N_4789,N_5528);
and U8474 (N_8474,N_3915,N_4064);
or U8475 (N_8475,N_3523,N_5162);
or U8476 (N_8476,N_5007,N_5741);
or U8477 (N_8477,N_3771,N_4568);
and U8478 (N_8478,N_5234,N_3882);
nand U8479 (N_8479,N_4840,N_3130);
nand U8480 (N_8480,N_3314,N_3871);
or U8481 (N_8481,N_4051,N_6058);
xnor U8482 (N_8482,N_3826,N_4715);
or U8483 (N_8483,N_5948,N_3632);
nand U8484 (N_8484,N_3420,N_3727);
or U8485 (N_8485,N_6014,N_4830);
xor U8486 (N_8486,N_3483,N_3893);
or U8487 (N_8487,N_4609,N_4928);
and U8488 (N_8488,N_4446,N_3266);
and U8489 (N_8489,N_4792,N_6209);
nor U8490 (N_8490,N_3201,N_3766);
or U8491 (N_8491,N_4158,N_4067);
nor U8492 (N_8492,N_6047,N_4416);
and U8493 (N_8493,N_5124,N_3950);
or U8494 (N_8494,N_5708,N_4562);
and U8495 (N_8495,N_5858,N_6058);
or U8496 (N_8496,N_3929,N_5635);
nand U8497 (N_8497,N_3555,N_3304);
nor U8498 (N_8498,N_4025,N_6214);
nor U8499 (N_8499,N_3459,N_3363);
nor U8500 (N_8500,N_5141,N_5589);
nor U8501 (N_8501,N_4304,N_3393);
and U8502 (N_8502,N_4798,N_4582);
and U8503 (N_8503,N_4955,N_4871);
or U8504 (N_8504,N_5383,N_5790);
and U8505 (N_8505,N_4901,N_4868);
nor U8506 (N_8506,N_3737,N_5722);
and U8507 (N_8507,N_5018,N_4820);
and U8508 (N_8508,N_6197,N_4134);
nand U8509 (N_8509,N_3231,N_3825);
nor U8510 (N_8510,N_4056,N_3882);
and U8511 (N_8511,N_3692,N_4596);
xnor U8512 (N_8512,N_6142,N_3559);
and U8513 (N_8513,N_3490,N_5595);
or U8514 (N_8514,N_4077,N_6110);
or U8515 (N_8515,N_3881,N_3227);
nor U8516 (N_8516,N_4902,N_3472);
and U8517 (N_8517,N_6175,N_3863);
and U8518 (N_8518,N_4926,N_3160);
nand U8519 (N_8519,N_5620,N_5999);
and U8520 (N_8520,N_3873,N_5651);
or U8521 (N_8521,N_4060,N_4599);
xnor U8522 (N_8522,N_3364,N_5894);
nor U8523 (N_8523,N_3712,N_4715);
nor U8524 (N_8524,N_3539,N_5350);
nand U8525 (N_8525,N_4343,N_5178);
nor U8526 (N_8526,N_4529,N_4609);
or U8527 (N_8527,N_3416,N_4681);
or U8528 (N_8528,N_5235,N_6037);
nand U8529 (N_8529,N_5939,N_3450);
nor U8530 (N_8530,N_4292,N_3236);
or U8531 (N_8531,N_3419,N_3567);
or U8532 (N_8532,N_4569,N_4753);
and U8533 (N_8533,N_6001,N_4746);
nand U8534 (N_8534,N_4519,N_5081);
or U8535 (N_8535,N_4390,N_4659);
or U8536 (N_8536,N_5858,N_3402);
nor U8537 (N_8537,N_3310,N_4765);
nor U8538 (N_8538,N_5483,N_6061);
nor U8539 (N_8539,N_5482,N_4079);
nor U8540 (N_8540,N_4845,N_4585);
nor U8541 (N_8541,N_5328,N_4051);
and U8542 (N_8542,N_6034,N_4342);
and U8543 (N_8543,N_5248,N_5114);
nand U8544 (N_8544,N_3480,N_3243);
nand U8545 (N_8545,N_5853,N_4311);
or U8546 (N_8546,N_5854,N_4133);
or U8547 (N_8547,N_3600,N_3253);
nand U8548 (N_8548,N_3552,N_3151);
and U8549 (N_8549,N_3540,N_3437);
nand U8550 (N_8550,N_5389,N_5157);
nand U8551 (N_8551,N_4617,N_4649);
or U8552 (N_8552,N_5542,N_3213);
or U8553 (N_8553,N_4553,N_5186);
or U8554 (N_8554,N_5555,N_5328);
and U8555 (N_8555,N_3472,N_5433);
nor U8556 (N_8556,N_3974,N_5115);
xnor U8557 (N_8557,N_5616,N_4343);
nor U8558 (N_8558,N_6246,N_4439);
nor U8559 (N_8559,N_5781,N_5927);
nand U8560 (N_8560,N_6237,N_5035);
nor U8561 (N_8561,N_5339,N_5720);
nand U8562 (N_8562,N_5504,N_5373);
nor U8563 (N_8563,N_3609,N_4750);
and U8564 (N_8564,N_5187,N_4334);
and U8565 (N_8565,N_5400,N_5318);
and U8566 (N_8566,N_6061,N_5981);
nor U8567 (N_8567,N_6115,N_4531);
nor U8568 (N_8568,N_4655,N_6135);
and U8569 (N_8569,N_6247,N_5950);
nand U8570 (N_8570,N_5711,N_5899);
or U8571 (N_8571,N_4343,N_4455);
nor U8572 (N_8572,N_5827,N_4738);
and U8573 (N_8573,N_3624,N_6180);
and U8574 (N_8574,N_3799,N_4977);
nand U8575 (N_8575,N_3515,N_4588);
nand U8576 (N_8576,N_3562,N_5479);
nor U8577 (N_8577,N_4187,N_5266);
nor U8578 (N_8578,N_3893,N_3583);
nand U8579 (N_8579,N_3900,N_5256);
nand U8580 (N_8580,N_5368,N_4300);
or U8581 (N_8581,N_4530,N_4601);
and U8582 (N_8582,N_5799,N_4578);
nand U8583 (N_8583,N_4739,N_3885);
or U8584 (N_8584,N_5452,N_5486);
or U8585 (N_8585,N_3973,N_3133);
nor U8586 (N_8586,N_5773,N_5745);
and U8587 (N_8587,N_5656,N_5434);
or U8588 (N_8588,N_5669,N_4436);
or U8589 (N_8589,N_5415,N_4509);
or U8590 (N_8590,N_5696,N_5184);
and U8591 (N_8591,N_3611,N_4352);
nor U8592 (N_8592,N_4924,N_6059);
nor U8593 (N_8593,N_4452,N_5244);
nor U8594 (N_8594,N_3284,N_5580);
nand U8595 (N_8595,N_5954,N_3669);
and U8596 (N_8596,N_5309,N_3159);
nor U8597 (N_8597,N_3312,N_4077);
nor U8598 (N_8598,N_3440,N_6137);
and U8599 (N_8599,N_4528,N_4947);
and U8600 (N_8600,N_5843,N_5893);
and U8601 (N_8601,N_4934,N_4415);
nand U8602 (N_8602,N_4063,N_5471);
nand U8603 (N_8603,N_3880,N_6138);
nand U8604 (N_8604,N_3274,N_5418);
or U8605 (N_8605,N_4126,N_4320);
or U8606 (N_8606,N_5585,N_5587);
nand U8607 (N_8607,N_6102,N_3463);
xor U8608 (N_8608,N_4721,N_4380);
xnor U8609 (N_8609,N_5249,N_4759);
nand U8610 (N_8610,N_3619,N_4872);
or U8611 (N_8611,N_4919,N_6171);
and U8612 (N_8612,N_4104,N_4641);
nor U8613 (N_8613,N_5304,N_4719);
and U8614 (N_8614,N_4209,N_5075);
nand U8615 (N_8615,N_4615,N_5166);
and U8616 (N_8616,N_4975,N_5120);
and U8617 (N_8617,N_3355,N_5735);
nand U8618 (N_8618,N_5701,N_4683);
xnor U8619 (N_8619,N_3638,N_5813);
nand U8620 (N_8620,N_5834,N_5446);
xnor U8621 (N_8621,N_6127,N_5468);
nor U8622 (N_8622,N_3383,N_6012);
and U8623 (N_8623,N_3172,N_6018);
and U8624 (N_8624,N_4223,N_3327);
nand U8625 (N_8625,N_4086,N_4475);
nand U8626 (N_8626,N_4917,N_3695);
or U8627 (N_8627,N_5773,N_5643);
and U8628 (N_8628,N_5087,N_3847);
xor U8629 (N_8629,N_6228,N_3605);
nand U8630 (N_8630,N_3652,N_4302);
or U8631 (N_8631,N_5076,N_5257);
xnor U8632 (N_8632,N_6178,N_3331);
nand U8633 (N_8633,N_6044,N_3802);
nand U8634 (N_8634,N_4966,N_5649);
or U8635 (N_8635,N_4319,N_4042);
and U8636 (N_8636,N_5361,N_4203);
and U8637 (N_8637,N_5468,N_5758);
nand U8638 (N_8638,N_3828,N_3272);
or U8639 (N_8639,N_3780,N_5789);
nor U8640 (N_8640,N_5329,N_5687);
xnor U8641 (N_8641,N_3287,N_5567);
and U8642 (N_8642,N_3434,N_4019);
and U8643 (N_8643,N_3184,N_5829);
xor U8644 (N_8644,N_5999,N_5366);
or U8645 (N_8645,N_5914,N_5304);
nand U8646 (N_8646,N_3823,N_3725);
nor U8647 (N_8647,N_5115,N_4390);
and U8648 (N_8648,N_6179,N_5572);
xnor U8649 (N_8649,N_5495,N_3573);
and U8650 (N_8650,N_5761,N_3823);
or U8651 (N_8651,N_5464,N_3403);
nor U8652 (N_8652,N_4542,N_4825);
xor U8653 (N_8653,N_3325,N_6155);
and U8654 (N_8654,N_5951,N_4433);
or U8655 (N_8655,N_3879,N_5044);
nand U8656 (N_8656,N_4931,N_3338);
or U8657 (N_8657,N_5608,N_4776);
xnor U8658 (N_8658,N_3586,N_4498);
and U8659 (N_8659,N_5878,N_3752);
nor U8660 (N_8660,N_5703,N_4004);
xor U8661 (N_8661,N_3645,N_5201);
and U8662 (N_8662,N_4960,N_4854);
nor U8663 (N_8663,N_4030,N_5954);
or U8664 (N_8664,N_3195,N_5701);
or U8665 (N_8665,N_3168,N_5290);
nor U8666 (N_8666,N_4694,N_4989);
or U8667 (N_8667,N_3699,N_4547);
or U8668 (N_8668,N_5879,N_5302);
nand U8669 (N_8669,N_4304,N_5434);
and U8670 (N_8670,N_5244,N_4930);
nor U8671 (N_8671,N_4305,N_4381);
nand U8672 (N_8672,N_3755,N_5512);
and U8673 (N_8673,N_3207,N_3357);
xnor U8674 (N_8674,N_5843,N_4722);
or U8675 (N_8675,N_6029,N_5342);
nor U8676 (N_8676,N_5502,N_3389);
or U8677 (N_8677,N_5792,N_5214);
nor U8678 (N_8678,N_4120,N_5124);
and U8679 (N_8679,N_5742,N_5725);
nor U8680 (N_8680,N_3665,N_5540);
xnor U8681 (N_8681,N_6145,N_5638);
nand U8682 (N_8682,N_5234,N_4918);
nand U8683 (N_8683,N_5074,N_3732);
or U8684 (N_8684,N_3636,N_3310);
or U8685 (N_8685,N_3506,N_5013);
or U8686 (N_8686,N_4177,N_4128);
nor U8687 (N_8687,N_4640,N_5531);
nor U8688 (N_8688,N_4255,N_5677);
or U8689 (N_8689,N_3797,N_4418);
nand U8690 (N_8690,N_3648,N_5862);
xnor U8691 (N_8691,N_4638,N_5984);
nor U8692 (N_8692,N_4066,N_3148);
and U8693 (N_8693,N_3294,N_5248);
nor U8694 (N_8694,N_4485,N_5068);
nor U8695 (N_8695,N_4258,N_3532);
nor U8696 (N_8696,N_5765,N_3512);
xnor U8697 (N_8697,N_5475,N_5327);
or U8698 (N_8698,N_4665,N_6175);
nor U8699 (N_8699,N_5688,N_5478);
or U8700 (N_8700,N_3502,N_5087);
and U8701 (N_8701,N_5639,N_3832);
and U8702 (N_8702,N_5524,N_5313);
xnor U8703 (N_8703,N_5537,N_6181);
or U8704 (N_8704,N_5211,N_5545);
or U8705 (N_8705,N_4436,N_4563);
and U8706 (N_8706,N_4237,N_5682);
or U8707 (N_8707,N_4919,N_4603);
or U8708 (N_8708,N_3339,N_3652);
or U8709 (N_8709,N_5915,N_5067);
xor U8710 (N_8710,N_3731,N_3634);
or U8711 (N_8711,N_5820,N_5503);
and U8712 (N_8712,N_5505,N_4903);
nand U8713 (N_8713,N_5333,N_3332);
and U8714 (N_8714,N_3331,N_4597);
and U8715 (N_8715,N_3961,N_5863);
or U8716 (N_8716,N_5913,N_5699);
nor U8717 (N_8717,N_4089,N_4768);
nand U8718 (N_8718,N_3740,N_5863);
nand U8719 (N_8719,N_5653,N_4369);
or U8720 (N_8720,N_5482,N_5036);
nor U8721 (N_8721,N_6111,N_3789);
nor U8722 (N_8722,N_5974,N_6031);
and U8723 (N_8723,N_4117,N_6130);
nand U8724 (N_8724,N_4666,N_6077);
or U8725 (N_8725,N_3375,N_4660);
or U8726 (N_8726,N_5485,N_3474);
and U8727 (N_8727,N_3897,N_3853);
nand U8728 (N_8728,N_3960,N_3715);
and U8729 (N_8729,N_4060,N_4609);
xor U8730 (N_8730,N_4785,N_6183);
or U8731 (N_8731,N_4051,N_5378);
nor U8732 (N_8732,N_5904,N_4327);
nand U8733 (N_8733,N_3784,N_5949);
and U8734 (N_8734,N_5477,N_4093);
and U8735 (N_8735,N_3434,N_6185);
nand U8736 (N_8736,N_5702,N_5512);
xnor U8737 (N_8737,N_5401,N_5018);
or U8738 (N_8738,N_3536,N_4730);
or U8739 (N_8739,N_5866,N_4407);
nand U8740 (N_8740,N_5761,N_3787);
and U8741 (N_8741,N_4482,N_3743);
nor U8742 (N_8742,N_3274,N_3856);
nand U8743 (N_8743,N_3839,N_3294);
nor U8744 (N_8744,N_3920,N_5387);
and U8745 (N_8745,N_5513,N_3176);
or U8746 (N_8746,N_5550,N_5530);
or U8747 (N_8747,N_4971,N_3905);
and U8748 (N_8748,N_4116,N_5674);
and U8749 (N_8749,N_4837,N_5916);
and U8750 (N_8750,N_3787,N_6078);
nand U8751 (N_8751,N_4447,N_5015);
nand U8752 (N_8752,N_3664,N_3723);
or U8753 (N_8753,N_4840,N_5135);
xnor U8754 (N_8754,N_3161,N_6050);
or U8755 (N_8755,N_5378,N_3443);
nor U8756 (N_8756,N_5481,N_5118);
or U8757 (N_8757,N_3838,N_4985);
nor U8758 (N_8758,N_3616,N_5594);
xnor U8759 (N_8759,N_3853,N_4556);
and U8760 (N_8760,N_4792,N_4036);
and U8761 (N_8761,N_4450,N_3819);
nand U8762 (N_8762,N_3776,N_6119);
nor U8763 (N_8763,N_3558,N_5861);
nor U8764 (N_8764,N_4051,N_3695);
nand U8765 (N_8765,N_3610,N_5804);
nand U8766 (N_8766,N_6065,N_3626);
xor U8767 (N_8767,N_3460,N_5877);
or U8768 (N_8768,N_3835,N_3611);
xor U8769 (N_8769,N_3545,N_3316);
and U8770 (N_8770,N_5144,N_5501);
or U8771 (N_8771,N_3824,N_5755);
nand U8772 (N_8772,N_3280,N_3320);
xor U8773 (N_8773,N_4671,N_4267);
and U8774 (N_8774,N_6107,N_3811);
and U8775 (N_8775,N_5106,N_5768);
nor U8776 (N_8776,N_4192,N_4757);
nand U8777 (N_8777,N_3401,N_4498);
nand U8778 (N_8778,N_6008,N_4114);
nor U8779 (N_8779,N_5859,N_4091);
xnor U8780 (N_8780,N_6104,N_4259);
xnor U8781 (N_8781,N_5429,N_3261);
and U8782 (N_8782,N_4879,N_3561);
or U8783 (N_8783,N_4451,N_3366);
nor U8784 (N_8784,N_3251,N_4216);
nor U8785 (N_8785,N_5338,N_4649);
nor U8786 (N_8786,N_4407,N_3892);
and U8787 (N_8787,N_4248,N_5060);
nand U8788 (N_8788,N_4334,N_4155);
nor U8789 (N_8789,N_3280,N_3880);
or U8790 (N_8790,N_3647,N_3465);
nor U8791 (N_8791,N_4882,N_4941);
and U8792 (N_8792,N_6106,N_3255);
nor U8793 (N_8793,N_5548,N_5728);
nor U8794 (N_8794,N_3218,N_6210);
nor U8795 (N_8795,N_6157,N_6039);
or U8796 (N_8796,N_5666,N_5524);
or U8797 (N_8797,N_5230,N_3850);
nor U8798 (N_8798,N_6198,N_3831);
nand U8799 (N_8799,N_3238,N_3531);
or U8800 (N_8800,N_3275,N_5110);
nor U8801 (N_8801,N_3506,N_5643);
xor U8802 (N_8802,N_5445,N_5213);
xnor U8803 (N_8803,N_3467,N_3812);
xnor U8804 (N_8804,N_6100,N_5809);
nand U8805 (N_8805,N_4537,N_5229);
or U8806 (N_8806,N_5392,N_5631);
xnor U8807 (N_8807,N_6066,N_4229);
and U8808 (N_8808,N_4819,N_3957);
nand U8809 (N_8809,N_6077,N_3621);
nor U8810 (N_8810,N_6071,N_3875);
or U8811 (N_8811,N_3678,N_4941);
and U8812 (N_8812,N_3203,N_3775);
nand U8813 (N_8813,N_4230,N_4349);
nor U8814 (N_8814,N_4494,N_3157);
and U8815 (N_8815,N_3922,N_5183);
nor U8816 (N_8816,N_4536,N_5026);
and U8817 (N_8817,N_3155,N_3744);
nor U8818 (N_8818,N_4680,N_4383);
or U8819 (N_8819,N_5614,N_5575);
nor U8820 (N_8820,N_5879,N_5996);
nor U8821 (N_8821,N_4754,N_5251);
nand U8822 (N_8822,N_4579,N_6116);
nand U8823 (N_8823,N_6124,N_5038);
or U8824 (N_8824,N_4038,N_5417);
or U8825 (N_8825,N_3839,N_3643);
nor U8826 (N_8826,N_4892,N_3315);
xor U8827 (N_8827,N_3752,N_5767);
xor U8828 (N_8828,N_4915,N_5988);
nor U8829 (N_8829,N_5160,N_3244);
xnor U8830 (N_8830,N_5774,N_4760);
or U8831 (N_8831,N_3332,N_3351);
nor U8832 (N_8832,N_4603,N_5739);
and U8833 (N_8833,N_5114,N_5700);
or U8834 (N_8834,N_4362,N_5384);
nand U8835 (N_8835,N_5353,N_5366);
and U8836 (N_8836,N_3300,N_4322);
or U8837 (N_8837,N_4953,N_4804);
or U8838 (N_8838,N_5567,N_4650);
xor U8839 (N_8839,N_4492,N_5530);
nor U8840 (N_8840,N_3260,N_4453);
or U8841 (N_8841,N_5804,N_4132);
xor U8842 (N_8842,N_5950,N_4720);
xnor U8843 (N_8843,N_5422,N_4581);
nor U8844 (N_8844,N_3285,N_3556);
nor U8845 (N_8845,N_5749,N_5391);
xor U8846 (N_8846,N_5992,N_5290);
xor U8847 (N_8847,N_4262,N_3745);
and U8848 (N_8848,N_4256,N_5091);
nor U8849 (N_8849,N_4166,N_4147);
nand U8850 (N_8850,N_5151,N_5830);
or U8851 (N_8851,N_5856,N_6236);
nand U8852 (N_8852,N_4157,N_3263);
or U8853 (N_8853,N_3193,N_5599);
nand U8854 (N_8854,N_4680,N_4375);
xor U8855 (N_8855,N_4363,N_3840);
nand U8856 (N_8856,N_6096,N_3881);
and U8857 (N_8857,N_6142,N_4523);
and U8858 (N_8858,N_3646,N_4368);
nand U8859 (N_8859,N_4749,N_5987);
xor U8860 (N_8860,N_3724,N_5410);
and U8861 (N_8861,N_4043,N_3899);
nor U8862 (N_8862,N_5719,N_5490);
xor U8863 (N_8863,N_5505,N_3365);
nor U8864 (N_8864,N_3151,N_5205);
or U8865 (N_8865,N_5340,N_5667);
or U8866 (N_8866,N_3653,N_4373);
or U8867 (N_8867,N_4547,N_4689);
or U8868 (N_8868,N_3483,N_5051);
nor U8869 (N_8869,N_4786,N_5884);
and U8870 (N_8870,N_5608,N_3263);
and U8871 (N_8871,N_5592,N_4393);
and U8872 (N_8872,N_4747,N_3315);
or U8873 (N_8873,N_5433,N_5778);
nand U8874 (N_8874,N_3980,N_4702);
nor U8875 (N_8875,N_5358,N_6248);
or U8876 (N_8876,N_4209,N_4789);
or U8877 (N_8877,N_4640,N_5231);
xor U8878 (N_8878,N_6155,N_4345);
nand U8879 (N_8879,N_5675,N_4411);
or U8880 (N_8880,N_4012,N_4771);
or U8881 (N_8881,N_4537,N_3770);
nor U8882 (N_8882,N_5832,N_4511);
nand U8883 (N_8883,N_4919,N_4028);
and U8884 (N_8884,N_5834,N_5641);
nor U8885 (N_8885,N_3868,N_4786);
nor U8886 (N_8886,N_4716,N_4708);
or U8887 (N_8887,N_4409,N_4579);
nor U8888 (N_8888,N_5990,N_5513);
nor U8889 (N_8889,N_5141,N_4619);
and U8890 (N_8890,N_4425,N_5388);
xnor U8891 (N_8891,N_3438,N_4410);
nand U8892 (N_8892,N_3392,N_4798);
nand U8893 (N_8893,N_5538,N_3136);
nand U8894 (N_8894,N_4344,N_4147);
nor U8895 (N_8895,N_4406,N_3372);
nand U8896 (N_8896,N_5952,N_3214);
nor U8897 (N_8897,N_5223,N_4627);
nor U8898 (N_8898,N_5504,N_6135);
and U8899 (N_8899,N_3388,N_5623);
xor U8900 (N_8900,N_3890,N_5359);
nand U8901 (N_8901,N_6114,N_3828);
nor U8902 (N_8902,N_3326,N_4694);
nand U8903 (N_8903,N_5050,N_4230);
or U8904 (N_8904,N_6146,N_4869);
nand U8905 (N_8905,N_3639,N_3963);
nor U8906 (N_8906,N_5343,N_5650);
nor U8907 (N_8907,N_3497,N_3381);
and U8908 (N_8908,N_5623,N_4280);
nand U8909 (N_8909,N_4238,N_5020);
nand U8910 (N_8910,N_4403,N_5003);
or U8911 (N_8911,N_3410,N_3910);
nor U8912 (N_8912,N_5557,N_3348);
and U8913 (N_8913,N_3615,N_4555);
and U8914 (N_8914,N_4762,N_5066);
nor U8915 (N_8915,N_4691,N_3383);
nor U8916 (N_8916,N_3579,N_3390);
and U8917 (N_8917,N_3566,N_5165);
or U8918 (N_8918,N_4575,N_3134);
and U8919 (N_8919,N_4716,N_4536);
and U8920 (N_8920,N_4593,N_5637);
or U8921 (N_8921,N_6155,N_4945);
nand U8922 (N_8922,N_4943,N_6208);
or U8923 (N_8923,N_3690,N_4416);
or U8924 (N_8924,N_3760,N_5104);
nand U8925 (N_8925,N_4537,N_3702);
xnor U8926 (N_8926,N_4683,N_5364);
nand U8927 (N_8927,N_4898,N_3910);
nand U8928 (N_8928,N_5765,N_6007);
nor U8929 (N_8929,N_3745,N_3149);
and U8930 (N_8930,N_4012,N_5829);
nor U8931 (N_8931,N_5917,N_5083);
and U8932 (N_8932,N_3484,N_4125);
or U8933 (N_8933,N_5748,N_5595);
or U8934 (N_8934,N_6158,N_6144);
nor U8935 (N_8935,N_3795,N_5345);
or U8936 (N_8936,N_3184,N_5487);
nand U8937 (N_8937,N_5958,N_4733);
nand U8938 (N_8938,N_4192,N_3662);
xor U8939 (N_8939,N_5133,N_3923);
and U8940 (N_8940,N_5141,N_3405);
or U8941 (N_8941,N_4990,N_4930);
nand U8942 (N_8942,N_4873,N_4605);
nand U8943 (N_8943,N_4865,N_3677);
and U8944 (N_8944,N_4648,N_5060);
nor U8945 (N_8945,N_3379,N_4649);
xnor U8946 (N_8946,N_4683,N_5780);
nor U8947 (N_8947,N_3311,N_6043);
or U8948 (N_8948,N_3172,N_5027);
nor U8949 (N_8949,N_5127,N_4915);
and U8950 (N_8950,N_3974,N_5326);
nor U8951 (N_8951,N_5914,N_5634);
nand U8952 (N_8952,N_5184,N_3473);
xnor U8953 (N_8953,N_4460,N_4774);
xor U8954 (N_8954,N_4164,N_3830);
nor U8955 (N_8955,N_6059,N_5200);
or U8956 (N_8956,N_5907,N_3942);
or U8957 (N_8957,N_3709,N_4754);
and U8958 (N_8958,N_3514,N_3412);
xnor U8959 (N_8959,N_4272,N_5150);
or U8960 (N_8960,N_3726,N_4975);
and U8961 (N_8961,N_6071,N_5767);
nand U8962 (N_8962,N_6087,N_4225);
nand U8963 (N_8963,N_4213,N_5052);
nor U8964 (N_8964,N_5641,N_6061);
nand U8965 (N_8965,N_3453,N_4550);
or U8966 (N_8966,N_5741,N_5221);
xor U8967 (N_8967,N_4730,N_6183);
nand U8968 (N_8968,N_5895,N_4838);
nor U8969 (N_8969,N_4961,N_5964);
and U8970 (N_8970,N_5412,N_5329);
xor U8971 (N_8971,N_5108,N_3653);
and U8972 (N_8972,N_3405,N_5372);
and U8973 (N_8973,N_5827,N_5191);
xor U8974 (N_8974,N_5842,N_5239);
nand U8975 (N_8975,N_4572,N_6208);
or U8976 (N_8976,N_3192,N_5300);
or U8977 (N_8977,N_3953,N_5291);
nor U8978 (N_8978,N_6205,N_3149);
nor U8979 (N_8979,N_6004,N_4693);
nand U8980 (N_8980,N_5745,N_4678);
and U8981 (N_8981,N_5838,N_4891);
and U8982 (N_8982,N_5881,N_4835);
or U8983 (N_8983,N_4164,N_3947);
nor U8984 (N_8984,N_3531,N_3988);
or U8985 (N_8985,N_3577,N_4683);
and U8986 (N_8986,N_5520,N_5309);
nor U8987 (N_8987,N_3227,N_3503);
nand U8988 (N_8988,N_3353,N_3771);
nand U8989 (N_8989,N_4313,N_3850);
nor U8990 (N_8990,N_4509,N_5088);
or U8991 (N_8991,N_4941,N_4445);
nor U8992 (N_8992,N_4097,N_5856);
nor U8993 (N_8993,N_6027,N_4709);
nor U8994 (N_8994,N_4357,N_4958);
and U8995 (N_8995,N_5178,N_4752);
or U8996 (N_8996,N_4226,N_3358);
and U8997 (N_8997,N_3163,N_3449);
nor U8998 (N_8998,N_5156,N_3532);
xnor U8999 (N_8999,N_4601,N_6231);
nand U9000 (N_9000,N_3480,N_3695);
or U9001 (N_9001,N_3934,N_6013);
xor U9002 (N_9002,N_5736,N_5472);
or U9003 (N_9003,N_5874,N_5570);
or U9004 (N_9004,N_3593,N_5115);
and U9005 (N_9005,N_4032,N_5800);
xor U9006 (N_9006,N_5205,N_3446);
nand U9007 (N_9007,N_4469,N_5229);
and U9008 (N_9008,N_3599,N_6034);
and U9009 (N_9009,N_4906,N_3252);
and U9010 (N_9010,N_3406,N_5747);
or U9011 (N_9011,N_4317,N_5268);
or U9012 (N_9012,N_4421,N_3222);
nor U9013 (N_9013,N_5934,N_5065);
or U9014 (N_9014,N_4139,N_3210);
nand U9015 (N_9015,N_4570,N_3484);
and U9016 (N_9016,N_4763,N_3672);
and U9017 (N_9017,N_5028,N_4377);
or U9018 (N_9018,N_5847,N_5965);
xor U9019 (N_9019,N_5596,N_6068);
nor U9020 (N_9020,N_5174,N_5621);
nor U9021 (N_9021,N_5518,N_3624);
and U9022 (N_9022,N_5999,N_4266);
or U9023 (N_9023,N_5009,N_5597);
or U9024 (N_9024,N_3355,N_5594);
or U9025 (N_9025,N_6035,N_3286);
nand U9026 (N_9026,N_6206,N_5203);
and U9027 (N_9027,N_4830,N_6038);
nor U9028 (N_9028,N_3644,N_5065);
nor U9029 (N_9029,N_4578,N_4713);
xor U9030 (N_9030,N_5217,N_4318);
xnor U9031 (N_9031,N_5416,N_5750);
and U9032 (N_9032,N_5273,N_5584);
and U9033 (N_9033,N_3199,N_5366);
nand U9034 (N_9034,N_5553,N_4303);
or U9035 (N_9035,N_3998,N_3446);
or U9036 (N_9036,N_3685,N_5171);
nor U9037 (N_9037,N_4991,N_3292);
nor U9038 (N_9038,N_4355,N_4847);
nand U9039 (N_9039,N_4949,N_4617);
and U9040 (N_9040,N_5316,N_5843);
xnor U9041 (N_9041,N_3160,N_3906);
or U9042 (N_9042,N_5450,N_4106);
xnor U9043 (N_9043,N_3494,N_3409);
and U9044 (N_9044,N_4166,N_5331);
and U9045 (N_9045,N_4150,N_6222);
nor U9046 (N_9046,N_5927,N_3658);
nor U9047 (N_9047,N_5627,N_3971);
and U9048 (N_9048,N_4469,N_4488);
nor U9049 (N_9049,N_3136,N_3636);
or U9050 (N_9050,N_3723,N_5665);
nor U9051 (N_9051,N_4791,N_3583);
and U9052 (N_9052,N_3546,N_3550);
or U9053 (N_9053,N_4626,N_3159);
nand U9054 (N_9054,N_3744,N_4899);
or U9055 (N_9055,N_5148,N_4424);
xnor U9056 (N_9056,N_5770,N_4782);
and U9057 (N_9057,N_4775,N_5923);
and U9058 (N_9058,N_4525,N_3145);
nand U9059 (N_9059,N_4513,N_5234);
nor U9060 (N_9060,N_5957,N_4531);
or U9061 (N_9061,N_5085,N_4863);
nand U9062 (N_9062,N_5833,N_3982);
nor U9063 (N_9063,N_3720,N_5065);
xnor U9064 (N_9064,N_3889,N_5354);
or U9065 (N_9065,N_5348,N_6140);
or U9066 (N_9066,N_5786,N_3531);
nand U9067 (N_9067,N_5462,N_5484);
or U9068 (N_9068,N_4109,N_4353);
nand U9069 (N_9069,N_5513,N_6116);
or U9070 (N_9070,N_3375,N_4264);
nor U9071 (N_9071,N_3151,N_4795);
nand U9072 (N_9072,N_3792,N_5906);
or U9073 (N_9073,N_3799,N_3990);
nand U9074 (N_9074,N_4780,N_4900);
nor U9075 (N_9075,N_4891,N_4121);
nand U9076 (N_9076,N_5956,N_3401);
nand U9077 (N_9077,N_4683,N_4303);
nor U9078 (N_9078,N_3200,N_4346);
nand U9079 (N_9079,N_6024,N_5934);
nor U9080 (N_9080,N_4787,N_4357);
and U9081 (N_9081,N_5958,N_5974);
nor U9082 (N_9082,N_3606,N_4480);
or U9083 (N_9083,N_5647,N_5554);
xnor U9084 (N_9084,N_3696,N_4656);
and U9085 (N_9085,N_4642,N_4531);
nand U9086 (N_9086,N_6210,N_6226);
nor U9087 (N_9087,N_5632,N_3319);
and U9088 (N_9088,N_6148,N_4297);
or U9089 (N_9089,N_4239,N_6115);
nand U9090 (N_9090,N_4527,N_4572);
or U9091 (N_9091,N_3334,N_4783);
and U9092 (N_9092,N_4323,N_3723);
or U9093 (N_9093,N_5275,N_3733);
nand U9094 (N_9094,N_4058,N_4373);
and U9095 (N_9095,N_3512,N_5474);
nand U9096 (N_9096,N_5939,N_4256);
xnor U9097 (N_9097,N_4733,N_4951);
and U9098 (N_9098,N_3817,N_5843);
nor U9099 (N_9099,N_5369,N_5119);
nand U9100 (N_9100,N_5801,N_5087);
nand U9101 (N_9101,N_3879,N_3999);
nor U9102 (N_9102,N_6109,N_5402);
nor U9103 (N_9103,N_4312,N_4255);
nand U9104 (N_9104,N_3684,N_3265);
and U9105 (N_9105,N_4158,N_4233);
and U9106 (N_9106,N_6178,N_5252);
nand U9107 (N_9107,N_6183,N_4680);
and U9108 (N_9108,N_3410,N_4335);
nand U9109 (N_9109,N_3789,N_3141);
and U9110 (N_9110,N_5126,N_4919);
nand U9111 (N_9111,N_4354,N_5015);
or U9112 (N_9112,N_3690,N_3921);
and U9113 (N_9113,N_4840,N_4669);
or U9114 (N_9114,N_5197,N_3895);
nor U9115 (N_9115,N_6040,N_5502);
nor U9116 (N_9116,N_3289,N_4059);
xnor U9117 (N_9117,N_3342,N_4626);
and U9118 (N_9118,N_4176,N_5631);
nand U9119 (N_9119,N_4897,N_4591);
nand U9120 (N_9120,N_3214,N_3351);
nor U9121 (N_9121,N_5997,N_6049);
nor U9122 (N_9122,N_5660,N_4022);
nor U9123 (N_9123,N_5163,N_5882);
or U9124 (N_9124,N_5022,N_5342);
and U9125 (N_9125,N_5402,N_3323);
nand U9126 (N_9126,N_3641,N_4256);
or U9127 (N_9127,N_4057,N_5672);
nor U9128 (N_9128,N_4437,N_3917);
nor U9129 (N_9129,N_6180,N_5996);
and U9130 (N_9130,N_3199,N_3789);
and U9131 (N_9131,N_4190,N_3375);
nor U9132 (N_9132,N_4194,N_5838);
and U9133 (N_9133,N_4227,N_5437);
and U9134 (N_9134,N_4977,N_6199);
or U9135 (N_9135,N_5200,N_4638);
or U9136 (N_9136,N_5388,N_3360);
or U9137 (N_9137,N_5385,N_5498);
xnor U9138 (N_9138,N_3920,N_4184);
nand U9139 (N_9139,N_5611,N_4568);
and U9140 (N_9140,N_5252,N_5671);
and U9141 (N_9141,N_3668,N_4715);
xor U9142 (N_9142,N_6121,N_4360);
nor U9143 (N_9143,N_6171,N_5451);
and U9144 (N_9144,N_4082,N_4131);
and U9145 (N_9145,N_4775,N_5910);
or U9146 (N_9146,N_5773,N_3447);
nand U9147 (N_9147,N_4007,N_3783);
nor U9148 (N_9148,N_5147,N_4091);
and U9149 (N_9149,N_5687,N_4022);
or U9150 (N_9150,N_3919,N_5328);
xnor U9151 (N_9151,N_4775,N_6181);
and U9152 (N_9152,N_5345,N_4305);
or U9153 (N_9153,N_3139,N_5364);
nand U9154 (N_9154,N_4542,N_3782);
nand U9155 (N_9155,N_3381,N_4343);
nand U9156 (N_9156,N_5162,N_5529);
nor U9157 (N_9157,N_4244,N_3799);
nand U9158 (N_9158,N_6201,N_4751);
or U9159 (N_9159,N_3416,N_6154);
and U9160 (N_9160,N_3516,N_6095);
xor U9161 (N_9161,N_4494,N_5704);
nor U9162 (N_9162,N_3383,N_3391);
nand U9163 (N_9163,N_5078,N_6181);
nand U9164 (N_9164,N_3705,N_5815);
nand U9165 (N_9165,N_4028,N_4829);
and U9166 (N_9166,N_5854,N_5937);
or U9167 (N_9167,N_3575,N_5363);
nand U9168 (N_9168,N_3746,N_4584);
and U9169 (N_9169,N_5373,N_3585);
or U9170 (N_9170,N_5753,N_4042);
nand U9171 (N_9171,N_4123,N_5540);
or U9172 (N_9172,N_5549,N_4584);
nand U9173 (N_9173,N_4271,N_5173);
or U9174 (N_9174,N_4098,N_5477);
and U9175 (N_9175,N_3951,N_5503);
and U9176 (N_9176,N_5354,N_5876);
and U9177 (N_9177,N_4512,N_5330);
nand U9178 (N_9178,N_4040,N_3916);
and U9179 (N_9179,N_3510,N_3167);
nand U9180 (N_9180,N_3372,N_3846);
and U9181 (N_9181,N_4814,N_4485);
nor U9182 (N_9182,N_3722,N_5154);
xor U9183 (N_9183,N_5418,N_4367);
and U9184 (N_9184,N_4702,N_4507);
and U9185 (N_9185,N_4269,N_5116);
nor U9186 (N_9186,N_4313,N_4463);
nand U9187 (N_9187,N_5665,N_3937);
or U9188 (N_9188,N_5729,N_4640);
or U9189 (N_9189,N_4762,N_5616);
nand U9190 (N_9190,N_5735,N_4726);
and U9191 (N_9191,N_5175,N_5395);
nand U9192 (N_9192,N_5594,N_5861);
nor U9193 (N_9193,N_5320,N_4596);
and U9194 (N_9194,N_4760,N_4775);
or U9195 (N_9195,N_3447,N_5394);
and U9196 (N_9196,N_3942,N_5683);
and U9197 (N_9197,N_5136,N_4359);
xor U9198 (N_9198,N_5065,N_5130);
xor U9199 (N_9199,N_5352,N_4641);
or U9200 (N_9200,N_4665,N_3131);
nor U9201 (N_9201,N_4076,N_5603);
nand U9202 (N_9202,N_3690,N_5152);
nand U9203 (N_9203,N_5273,N_5558);
or U9204 (N_9204,N_5455,N_6017);
or U9205 (N_9205,N_5115,N_3647);
nor U9206 (N_9206,N_3631,N_6152);
or U9207 (N_9207,N_5374,N_3539);
or U9208 (N_9208,N_5969,N_4128);
nand U9209 (N_9209,N_5990,N_5614);
and U9210 (N_9210,N_6040,N_3175);
nand U9211 (N_9211,N_4474,N_4877);
or U9212 (N_9212,N_3634,N_4495);
or U9213 (N_9213,N_5268,N_3785);
nand U9214 (N_9214,N_5564,N_5683);
nand U9215 (N_9215,N_3420,N_3701);
and U9216 (N_9216,N_5936,N_4232);
or U9217 (N_9217,N_6155,N_3967);
nand U9218 (N_9218,N_3492,N_4293);
nand U9219 (N_9219,N_5215,N_6187);
nor U9220 (N_9220,N_5067,N_5095);
nor U9221 (N_9221,N_3976,N_4634);
nand U9222 (N_9222,N_4703,N_3300);
nand U9223 (N_9223,N_4318,N_3957);
nand U9224 (N_9224,N_4028,N_3517);
or U9225 (N_9225,N_6227,N_3382);
or U9226 (N_9226,N_4008,N_3905);
and U9227 (N_9227,N_5102,N_3581);
or U9228 (N_9228,N_3180,N_3491);
and U9229 (N_9229,N_4881,N_4707);
and U9230 (N_9230,N_5697,N_4529);
or U9231 (N_9231,N_5018,N_6216);
and U9232 (N_9232,N_4615,N_3800);
nand U9233 (N_9233,N_5601,N_3293);
or U9234 (N_9234,N_4312,N_4072);
nand U9235 (N_9235,N_3865,N_3648);
nand U9236 (N_9236,N_5140,N_4039);
nand U9237 (N_9237,N_4185,N_4684);
xnor U9238 (N_9238,N_5889,N_3912);
nor U9239 (N_9239,N_4857,N_4861);
nor U9240 (N_9240,N_4493,N_5839);
or U9241 (N_9241,N_4591,N_4694);
and U9242 (N_9242,N_6078,N_3330);
xnor U9243 (N_9243,N_5980,N_3658);
nor U9244 (N_9244,N_4196,N_3763);
xor U9245 (N_9245,N_5963,N_4047);
and U9246 (N_9246,N_4952,N_5347);
nor U9247 (N_9247,N_5089,N_3185);
or U9248 (N_9248,N_5682,N_3287);
nor U9249 (N_9249,N_3170,N_3714);
and U9250 (N_9250,N_5264,N_4266);
nand U9251 (N_9251,N_6214,N_5194);
or U9252 (N_9252,N_5632,N_4014);
and U9253 (N_9253,N_5144,N_3386);
and U9254 (N_9254,N_4484,N_6083);
nor U9255 (N_9255,N_5060,N_3778);
or U9256 (N_9256,N_4042,N_3984);
and U9257 (N_9257,N_6213,N_4168);
xor U9258 (N_9258,N_4230,N_4288);
nand U9259 (N_9259,N_3451,N_4732);
and U9260 (N_9260,N_3628,N_4413);
or U9261 (N_9261,N_5633,N_3258);
nand U9262 (N_9262,N_3923,N_4678);
nor U9263 (N_9263,N_3983,N_3848);
and U9264 (N_9264,N_5221,N_3525);
and U9265 (N_9265,N_4962,N_4885);
nor U9266 (N_9266,N_3585,N_4811);
and U9267 (N_9267,N_3978,N_3414);
xnor U9268 (N_9268,N_5214,N_4334);
and U9269 (N_9269,N_6053,N_6228);
nand U9270 (N_9270,N_4239,N_5191);
or U9271 (N_9271,N_4242,N_5687);
and U9272 (N_9272,N_4474,N_5139);
and U9273 (N_9273,N_4051,N_4875);
nand U9274 (N_9274,N_6041,N_3469);
or U9275 (N_9275,N_4185,N_5230);
nor U9276 (N_9276,N_4702,N_5942);
nor U9277 (N_9277,N_5851,N_5739);
nor U9278 (N_9278,N_5223,N_4203);
nand U9279 (N_9279,N_3666,N_5565);
xnor U9280 (N_9280,N_3433,N_5040);
and U9281 (N_9281,N_3229,N_4510);
nand U9282 (N_9282,N_6139,N_5493);
nand U9283 (N_9283,N_5851,N_4012);
nor U9284 (N_9284,N_5113,N_6245);
nor U9285 (N_9285,N_5084,N_5122);
nor U9286 (N_9286,N_4485,N_6123);
or U9287 (N_9287,N_3755,N_6158);
or U9288 (N_9288,N_5351,N_4569);
and U9289 (N_9289,N_3534,N_4784);
nand U9290 (N_9290,N_3614,N_4637);
xnor U9291 (N_9291,N_3910,N_3394);
or U9292 (N_9292,N_4484,N_5359);
nor U9293 (N_9293,N_5701,N_5683);
or U9294 (N_9294,N_4604,N_3630);
nand U9295 (N_9295,N_4562,N_3455);
nor U9296 (N_9296,N_5817,N_4336);
nand U9297 (N_9297,N_3795,N_4770);
nand U9298 (N_9298,N_4080,N_5381);
or U9299 (N_9299,N_4502,N_5897);
or U9300 (N_9300,N_4438,N_5469);
and U9301 (N_9301,N_3217,N_4873);
nor U9302 (N_9302,N_6044,N_4759);
nand U9303 (N_9303,N_4139,N_3354);
or U9304 (N_9304,N_5101,N_3492);
or U9305 (N_9305,N_4038,N_6131);
and U9306 (N_9306,N_3326,N_4086);
nor U9307 (N_9307,N_5724,N_3742);
nand U9308 (N_9308,N_5662,N_3175);
or U9309 (N_9309,N_5029,N_3401);
nand U9310 (N_9310,N_4209,N_4899);
and U9311 (N_9311,N_5439,N_5964);
and U9312 (N_9312,N_4470,N_3512);
and U9313 (N_9313,N_4610,N_3996);
or U9314 (N_9314,N_5342,N_5903);
nand U9315 (N_9315,N_5320,N_5660);
xor U9316 (N_9316,N_4859,N_5123);
or U9317 (N_9317,N_3997,N_5542);
or U9318 (N_9318,N_5790,N_6076);
or U9319 (N_9319,N_4306,N_5776);
nor U9320 (N_9320,N_4339,N_4645);
nor U9321 (N_9321,N_4570,N_4190);
nand U9322 (N_9322,N_4064,N_5186);
nand U9323 (N_9323,N_3897,N_3375);
xor U9324 (N_9324,N_5768,N_4317);
nand U9325 (N_9325,N_4587,N_4933);
or U9326 (N_9326,N_5365,N_5543);
nor U9327 (N_9327,N_4736,N_3785);
nor U9328 (N_9328,N_4341,N_4415);
nand U9329 (N_9329,N_4179,N_4072);
xnor U9330 (N_9330,N_5178,N_5918);
nor U9331 (N_9331,N_4255,N_4819);
or U9332 (N_9332,N_3357,N_6148);
nor U9333 (N_9333,N_3460,N_4569);
and U9334 (N_9334,N_3603,N_3153);
or U9335 (N_9335,N_5185,N_6174);
nand U9336 (N_9336,N_3480,N_5269);
nand U9337 (N_9337,N_3220,N_3894);
or U9338 (N_9338,N_6205,N_4156);
nor U9339 (N_9339,N_5356,N_6248);
nor U9340 (N_9340,N_4140,N_5410);
xor U9341 (N_9341,N_6083,N_4813);
nor U9342 (N_9342,N_4251,N_5748);
or U9343 (N_9343,N_3781,N_5821);
nor U9344 (N_9344,N_4934,N_4006);
and U9345 (N_9345,N_4780,N_3494);
or U9346 (N_9346,N_3576,N_5987);
xnor U9347 (N_9347,N_5227,N_4944);
or U9348 (N_9348,N_5106,N_4125);
nor U9349 (N_9349,N_3542,N_4129);
or U9350 (N_9350,N_5897,N_4446);
or U9351 (N_9351,N_5235,N_5651);
and U9352 (N_9352,N_4852,N_4945);
or U9353 (N_9353,N_4825,N_5323);
nand U9354 (N_9354,N_4588,N_3432);
and U9355 (N_9355,N_3282,N_3914);
nor U9356 (N_9356,N_5186,N_3819);
nor U9357 (N_9357,N_5550,N_4431);
nor U9358 (N_9358,N_3512,N_4898);
or U9359 (N_9359,N_6248,N_3466);
or U9360 (N_9360,N_3873,N_5825);
nand U9361 (N_9361,N_5857,N_5789);
and U9362 (N_9362,N_4169,N_3649);
nand U9363 (N_9363,N_5676,N_4988);
nor U9364 (N_9364,N_3964,N_5801);
nor U9365 (N_9365,N_4126,N_5240);
nor U9366 (N_9366,N_3295,N_4627);
xor U9367 (N_9367,N_3280,N_5616);
and U9368 (N_9368,N_5988,N_3164);
xnor U9369 (N_9369,N_5292,N_4541);
or U9370 (N_9370,N_5081,N_6000);
nand U9371 (N_9371,N_3142,N_5633);
and U9372 (N_9372,N_3301,N_3173);
nand U9373 (N_9373,N_4993,N_6192);
nor U9374 (N_9374,N_4558,N_4914);
and U9375 (N_9375,N_8288,N_6344);
and U9376 (N_9376,N_6475,N_7542);
or U9377 (N_9377,N_6489,N_8338);
nor U9378 (N_9378,N_6274,N_7759);
or U9379 (N_9379,N_7595,N_6968);
nand U9380 (N_9380,N_7727,N_7691);
and U9381 (N_9381,N_7577,N_6350);
nand U9382 (N_9382,N_7621,N_7768);
and U9383 (N_9383,N_7706,N_7236);
or U9384 (N_9384,N_8611,N_7323);
nand U9385 (N_9385,N_8517,N_8905);
and U9386 (N_9386,N_8219,N_6850);
or U9387 (N_9387,N_6290,N_7290);
or U9388 (N_9388,N_7619,N_7710);
or U9389 (N_9389,N_7450,N_8968);
xnor U9390 (N_9390,N_9205,N_8590);
and U9391 (N_9391,N_6605,N_6785);
nand U9392 (N_9392,N_8064,N_6975);
and U9393 (N_9393,N_8986,N_8130);
xnor U9394 (N_9394,N_9179,N_8558);
or U9395 (N_9395,N_7413,N_6842);
or U9396 (N_9396,N_6745,N_8319);
and U9397 (N_9397,N_7735,N_6533);
nand U9398 (N_9398,N_6513,N_7658);
or U9399 (N_9399,N_7504,N_8753);
nor U9400 (N_9400,N_6469,N_9023);
nand U9401 (N_9401,N_8736,N_8058);
nor U9402 (N_9402,N_7563,N_9144);
and U9403 (N_9403,N_7137,N_8538);
or U9404 (N_9404,N_9087,N_8857);
nand U9405 (N_9405,N_7470,N_7113);
or U9406 (N_9406,N_7250,N_7221);
or U9407 (N_9407,N_7875,N_6281);
or U9408 (N_9408,N_8536,N_6947);
nor U9409 (N_9409,N_9268,N_8379);
and U9410 (N_9410,N_7535,N_6788);
nor U9411 (N_9411,N_6813,N_6560);
nand U9412 (N_9412,N_8705,N_8795);
nand U9413 (N_9413,N_7705,N_8474);
and U9414 (N_9414,N_9039,N_9364);
nor U9415 (N_9415,N_8061,N_8177);
nand U9416 (N_9416,N_7567,N_6267);
nand U9417 (N_9417,N_8835,N_8846);
or U9418 (N_9418,N_8443,N_9278);
and U9419 (N_9419,N_7270,N_7523);
or U9420 (N_9420,N_7093,N_7066);
and U9421 (N_9421,N_7274,N_6820);
and U9422 (N_9422,N_8455,N_7989);
or U9423 (N_9423,N_9090,N_8457);
or U9424 (N_9424,N_8133,N_6321);
nor U9425 (N_9425,N_8568,N_7019);
nand U9426 (N_9426,N_7394,N_8527);
nand U9427 (N_9427,N_8027,N_8083);
and U9428 (N_9428,N_8959,N_8132);
nor U9429 (N_9429,N_7639,N_8112);
or U9430 (N_9430,N_6926,N_9310);
or U9431 (N_9431,N_7215,N_8515);
or U9432 (N_9432,N_7089,N_7515);
and U9433 (N_9433,N_7483,N_7374);
nand U9434 (N_9434,N_7443,N_8943);
or U9435 (N_9435,N_8151,N_8648);
and U9436 (N_9436,N_8440,N_8283);
nand U9437 (N_9437,N_8211,N_7207);
nor U9438 (N_9438,N_7335,N_6561);
nand U9439 (N_9439,N_6995,N_6340);
nand U9440 (N_9440,N_7874,N_7338);
nor U9441 (N_9441,N_7712,N_7722);
or U9442 (N_9442,N_9164,N_7302);
xnor U9443 (N_9443,N_6633,N_9207);
xnor U9444 (N_9444,N_6728,N_6763);
xor U9445 (N_9445,N_7431,N_8250);
nor U9446 (N_9446,N_7564,N_8470);
nor U9447 (N_9447,N_8452,N_7540);
and U9448 (N_9448,N_7169,N_8799);
nand U9449 (N_9449,N_6473,N_6521);
and U9450 (N_9450,N_7162,N_8638);
and U9451 (N_9451,N_9271,N_6681);
and U9452 (N_9452,N_6634,N_7034);
nor U9453 (N_9453,N_8604,N_9221);
nor U9454 (N_9454,N_9254,N_6414);
and U9455 (N_9455,N_6609,N_9143);
nand U9456 (N_9456,N_7301,N_8144);
and U9457 (N_9457,N_7726,N_8892);
and U9458 (N_9458,N_7248,N_8302);
nand U9459 (N_9459,N_8547,N_7175);
xor U9460 (N_9460,N_7823,N_8758);
nor U9461 (N_9461,N_8624,N_8264);
and U9462 (N_9462,N_6811,N_7970);
or U9463 (N_9463,N_8370,N_8691);
xnor U9464 (N_9464,N_9238,N_9145);
and U9465 (N_9465,N_7913,N_8046);
nor U9466 (N_9466,N_6896,N_6250);
and U9467 (N_9467,N_6251,N_7001);
or U9468 (N_9468,N_8725,N_9022);
or U9469 (N_9469,N_8693,N_6464);
or U9470 (N_9470,N_7776,N_8883);
nor U9471 (N_9471,N_6574,N_6749);
nor U9472 (N_9472,N_9195,N_6640);
or U9473 (N_9473,N_6562,N_7841);
xor U9474 (N_9474,N_7956,N_8819);
nand U9475 (N_9475,N_8908,N_9089);
nand U9476 (N_9476,N_9163,N_7958);
or U9477 (N_9477,N_6596,N_8382);
nor U9478 (N_9478,N_8377,N_6752);
nand U9479 (N_9479,N_9313,N_7618);
and U9480 (N_9480,N_7486,N_7472);
and U9481 (N_9481,N_8350,N_8301);
and U9482 (N_9482,N_8872,N_7707);
and U9483 (N_9483,N_8769,N_8684);
nor U9484 (N_9484,N_6935,N_7798);
and U9485 (N_9485,N_8281,N_9015);
nand U9486 (N_9486,N_8496,N_8124);
xor U9487 (N_9487,N_7031,N_8494);
nor U9488 (N_9488,N_7231,N_7350);
or U9489 (N_9489,N_6747,N_9316);
nand U9490 (N_9490,N_8328,N_6392);
nand U9491 (N_9491,N_8954,N_6305);
and U9492 (N_9492,N_8561,N_7623);
nand U9493 (N_9493,N_6662,N_7312);
and U9494 (N_9494,N_8360,N_9199);
nand U9495 (N_9495,N_8808,N_8492);
nor U9496 (N_9496,N_6467,N_7008);
or U9497 (N_9497,N_7347,N_8717);
xnor U9498 (N_9498,N_8848,N_7683);
xor U9499 (N_9499,N_7369,N_6872);
and U9500 (N_9500,N_8263,N_8341);
nand U9501 (N_9501,N_8788,N_8078);
or U9502 (N_9502,N_8922,N_7636);
or U9503 (N_9503,N_7928,N_7141);
nand U9504 (N_9504,N_7140,N_7825);
nor U9505 (N_9505,N_6904,N_7033);
nor U9506 (N_9506,N_9257,N_8429);
nand U9507 (N_9507,N_7708,N_8489);
xnor U9508 (N_9508,N_9370,N_7490);
or U9509 (N_9509,N_6734,N_6461);
or U9510 (N_9510,N_6567,N_6621);
and U9511 (N_9511,N_7397,N_8444);
xor U9512 (N_9512,N_7204,N_9304);
and U9513 (N_9513,N_8395,N_8916);
xnor U9514 (N_9514,N_8564,N_6396);
or U9515 (N_9515,N_8111,N_8563);
nand U9516 (N_9516,N_8890,N_7056);
nand U9517 (N_9517,N_8314,N_8118);
xor U9518 (N_9518,N_6806,N_8394);
xor U9519 (N_9519,N_7822,N_6529);
or U9520 (N_9520,N_8179,N_8389);
nand U9521 (N_9521,N_7428,N_8269);
xnor U9522 (N_9522,N_6708,N_8204);
nand U9523 (N_9523,N_7931,N_7929);
nor U9524 (N_9524,N_7345,N_6337);
or U9525 (N_9525,N_6590,N_9160);
or U9526 (N_9526,N_9248,N_7884);
nor U9527 (N_9527,N_8958,N_7362);
nor U9528 (N_9528,N_6836,N_6351);
and U9529 (N_9529,N_8372,N_9121);
xor U9530 (N_9530,N_7367,N_7408);
or U9531 (N_9531,N_7600,N_8790);
nand U9532 (N_9532,N_8422,N_8294);
nor U9533 (N_9533,N_8679,N_6696);
and U9534 (N_9534,N_8800,N_6397);
and U9535 (N_9535,N_7295,N_7393);
and U9536 (N_9536,N_8217,N_7286);
nand U9537 (N_9537,N_6494,N_9009);
and U9538 (N_9538,N_6685,N_9214);
nor U9539 (N_9539,N_8742,N_6606);
nand U9540 (N_9540,N_6581,N_8096);
and U9541 (N_9541,N_9249,N_6415);
nand U9542 (N_9542,N_7084,N_8632);
or U9543 (N_9543,N_9171,N_8114);
nand U9544 (N_9544,N_6299,N_8791);
nor U9545 (N_9545,N_8893,N_8451);
and U9546 (N_9546,N_6722,N_8581);
nor U9547 (N_9547,N_8593,N_9369);
or U9548 (N_9548,N_8412,N_7488);
and U9549 (N_9549,N_8070,N_8598);
and U9550 (N_9550,N_6761,N_8775);
nor U9551 (N_9551,N_7499,N_7531);
or U9552 (N_9552,N_9020,N_6673);
and U9553 (N_9553,N_8562,N_7136);
or U9554 (N_9554,N_9103,N_7533);
nor U9555 (N_9555,N_9129,N_9234);
nor U9556 (N_9556,N_8170,N_6758);
or U9557 (N_9557,N_7593,N_7354);
or U9558 (N_9558,N_8765,N_8843);
xnor U9559 (N_9559,N_7261,N_8792);
nor U9560 (N_9560,N_9110,N_7607);
nand U9561 (N_9561,N_6316,N_7779);
or U9562 (N_9562,N_7608,N_8870);
nand U9563 (N_9563,N_6831,N_7580);
and U9564 (N_9564,N_6530,N_9032);
or U9565 (N_9565,N_7037,N_6952);
or U9566 (N_9566,N_8777,N_8191);
and U9567 (N_9567,N_6355,N_9050);
nand U9568 (N_9568,N_8471,N_7186);
and U9569 (N_9569,N_6262,N_6500);
or U9570 (N_9570,N_6538,N_9134);
nor U9571 (N_9571,N_8486,N_9201);
and U9572 (N_9572,N_6990,N_6411);
and U9573 (N_9573,N_9099,N_8266);
and U9574 (N_9574,N_9055,N_8384);
nand U9575 (N_9575,N_8094,N_6649);
nor U9576 (N_9576,N_6376,N_7087);
nand U9577 (N_9577,N_6864,N_9013);
or U9578 (N_9578,N_8738,N_8887);
or U9579 (N_9579,N_7665,N_7674);
or U9580 (N_9580,N_6965,N_7805);
nor U9581 (N_9581,N_8837,N_8131);
xor U9582 (N_9582,N_7660,N_7662);
nor U9583 (N_9583,N_7437,N_9077);
nor U9584 (N_9584,N_7571,N_7276);
nor U9585 (N_9585,N_6804,N_6720);
nor U9586 (N_9586,N_8122,N_6393);
nand U9587 (N_9587,N_8024,N_6568);
or U9588 (N_9588,N_7255,N_9166);
nor U9589 (N_9589,N_7349,N_6384);
nand U9590 (N_9590,N_8193,N_8347);
and U9591 (N_9591,N_6797,N_6751);
and U9592 (N_9592,N_7663,N_7234);
nand U9593 (N_9593,N_7208,N_8825);
or U9594 (N_9594,N_6943,N_8862);
nand U9595 (N_9595,N_8999,N_7506);
and U9596 (N_9596,N_6347,N_8012);
or U9597 (N_9597,N_7425,N_8498);
nor U9598 (N_9598,N_8618,N_9290);
xnor U9599 (N_9599,N_8866,N_8368);
nor U9600 (N_9600,N_7797,N_7919);
xnor U9601 (N_9601,N_7902,N_7685);
or U9602 (N_9602,N_7195,N_6724);
nor U9603 (N_9603,N_6774,N_8241);
nor U9604 (N_9604,N_8052,N_6525);
and U9605 (N_9605,N_8183,N_6900);
nor U9606 (N_9606,N_8493,N_7119);
and U9607 (N_9607,N_6424,N_8961);
or U9608 (N_9608,N_7632,N_8930);
and U9609 (N_9609,N_7733,N_7183);
nand U9610 (N_9610,N_8782,N_6981);
nor U9611 (N_9611,N_6725,N_7028);
and U9612 (N_9612,N_6795,N_7545);
nand U9613 (N_9613,N_6667,N_6508);
nand U9614 (N_9614,N_7570,N_8861);
and U9615 (N_9615,N_6729,N_7173);
nor U9616 (N_9616,N_7973,N_8582);
xor U9617 (N_9617,N_8841,N_8583);
nor U9618 (N_9618,N_7783,N_6933);
or U9619 (N_9619,N_9330,N_8724);
xor U9620 (N_9620,N_6284,N_7383);
nor U9621 (N_9621,N_8594,N_9016);
nor U9622 (N_9622,N_8567,N_7258);
or U9623 (N_9623,N_7435,N_7224);
nand U9624 (N_9624,N_7211,N_7481);
nor U9625 (N_9625,N_6268,N_8585);
nor U9626 (N_9626,N_6358,N_7620);
and U9627 (N_9627,N_8212,N_6466);
and U9628 (N_9628,N_6871,N_9085);
nor U9629 (N_9629,N_7824,N_8935);
nand U9630 (N_9630,N_6925,N_7288);
nand U9631 (N_9631,N_7793,N_7628);
and U9632 (N_9632,N_8352,N_8414);
and U9633 (N_9633,N_9049,N_9127);
nand U9634 (N_9634,N_7852,N_6520);
nor U9635 (N_9635,N_8692,N_7280);
or U9636 (N_9636,N_8316,N_7306);
nand U9637 (N_9637,N_8553,N_7452);
and U9638 (N_9638,N_8048,N_6471);
and U9639 (N_9639,N_6861,N_7401);
or U9640 (N_9640,N_8428,N_8362);
or U9641 (N_9641,N_9216,N_9117);
nor U9642 (N_9642,N_7149,N_6825);
nand U9643 (N_9643,N_8802,N_7441);
nor U9644 (N_9644,N_7802,N_8163);
xor U9645 (N_9645,N_6846,N_7878);
nor U9646 (N_9646,N_6913,N_8619);
xnor U9647 (N_9647,N_7667,N_8977);
and U9648 (N_9648,N_7879,N_7273);
nor U9649 (N_9649,N_7127,N_7760);
xnor U9650 (N_9650,N_9107,N_8912);
nor U9651 (N_9651,N_7122,N_9247);
nand U9652 (N_9652,N_9305,N_7867);
nor U9653 (N_9653,N_9230,N_7314);
or U9654 (N_9654,N_9031,N_6647);
and U9655 (N_9655,N_7903,N_7526);
or U9656 (N_9656,N_6378,N_9215);
nor U9657 (N_9657,N_7611,N_7055);
xor U9658 (N_9658,N_8107,N_9111);
or U9659 (N_9659,N_8859,N_8888);
nand U9660 (N_9660,N_8546,N_7922);
and U9661 (N_9661,N_8949,N_7921);
or U9662 (N_9662,N_8097,N_8853);
nor U9663 (N_9663,N_9133,N_7741);
or U9664 (N_9664,N_6931,N_7859);
and U9665 (N_9665,N_7990,N_6757);
and U9666 (N_9666,N_6873,N_8534);
xor U9667 (N_9667,N_7178,N_6556);
nand U9668 (N_9668,N_7512,N_7372);
and U9669 (N_9669,N_7709,N_7426);
or U9670 (N_9670,N_7686,N_6716);
nand U9671 (N_9671,N_8484,N_8655);
nand U9672 (N_9672,N_9296,N_6789);
nor U9673 (N_9673,N_6823,N_7510);
and U9674 (N_9674,N_8102,N_7099);
nand U9675 (N_9675,N_6840,N_6723);
or U9676 (N_9676,N_7151,N_7495);
nand U9677 (N_9677,N_8423,N_9182);
or U9678 (N_9678,N_9312,N_7230);
and U9679 (N_9679,N_8205,N_7023);
and U9680 (N_9680,N_8729,N_6519);
or U9681 (N_9681,N_9005,N_8544);
and U9682 (N_9682,N_8182,N_8188);
nand U9683 (N_9683,N_8974,N_8806);
nand U9684 (N_9684,N_6727,N_8672);
or U9685 (N_9685,N_6453,N_9357);
and U9686 (N_9686,N_7774,N_9261);
and U9687 (N_9687,N_6265,N_9322);
or U9688 (N_9688,N_6741,N_6571);
xnor U9689 (N_9689,N_8225,N_8067);
nor U9690 (N_9690,N_8522,N_7789);
nor U9691 (N_9691,N_8464,N_8821);
and U9692 (N_9692,N_8123,N_7134);
and U9693 (N_9693,N_6627,N_9035);
and U9694 (N_9694,N_8573,N_9102);
and U9695 (N_9695,N_9096,N_8727);
xnor U9696 (N_9696,N_8271,N_8774);
and U9697 (N_9697,N_6859,N_7461);
nor U9698 (N_9698,N_7171,N_7536);
nor U9699 (N_9699,N_8572,N_7364);
or U9700 (N_9700,N_6541,N_7749);
nor U9701 (N_9701,N_8458,N_6821);
nand U9702 (N_9702,N_7688,N_7359);
or U9703 (N_9703,N_7120,N_8432);
and U9704 (N_9704,N_6370,N_7344);
or U9705 (N_9705,N_9046,N_7615);
nor U9706 (N_9706,N_9292,N_9297);
nor U9707 (N_9707,N_7525,N_7676);
or U9708 (N_9708,N_6549,N_8086);
or U9709 (N_9709,N_8885,N_9209);
and U9710 (N_9710,N_9033,N_6956);
xor U9711 (N_9711,N_7521,N_7402);
nand U9712 (N_9712,N_7713,N_7039);
nand U9713 (N_9713,N_8715,N_8145);
or U9714 (N_9714,N_7163,N_6955);
or U9715 (N_9715,N_7924,N_8840);
or U9716 (N_9716,N_6684,N_8155);
xor U9717 (N_9717,N_8540,N_9122);
nor U9718 (N_9718,N_8010,N_9281);
or U9719 (N_9719,N_8026,N_7740);
xnor U9720 (N_9720,N_9233,N_6543);
nor U9721 (N_9721,N_9365,N_9367);
or U9722 (N_9722,N_8948,N_6781);
nand U9723 (N_9723,N_6504,N_9363);
nor U9724 (N_9724,N_6320,N_8303);
nand U9725 (N_9725,N_6712,N_8380);
nor U9726 (N_9726,N_7070,N_6579);
and U9727 (N_9727,N_7747,N_7761);
xor U9728 (N_9728,N_7769,N_9246);
nor U9729 (N_9729,N_6462,N_6887);
and U9730 (N_9730,N_8882,N_6570);
nor U9731 (N_9731,N_7478,N_6578);
and U9732 (N_9732,N_7750,N_8323);
xnor U9733 (N_9733,N_8981,N_8324);
or U9734 (N_9734,N_8577,N_7871);
nand U9735 (N_9735,N_7308,N_8374);
nand U9736 (N_9736,N_7539,N_7380);
nand U9737 (N_9737,N_7090,N_7101);
nor U9738 (N_9738,N_7612,N_6969);
and U9739 (N_9739,N_6330,N_6285);
nand U9740 (N_9740,N_8663,N_8056);
or U9741 (N_9741,N_9081,N_8673);
nand U9742 (N_9742,N_7240,N_6610);
and U9743 (N_9743,N_6550,N_9272);
xnor U9744 (N_9744,N_7910,N_7946);
and U9745 (N_9745,N_6275,N_6488);
or U9746 (N_9746,N_9206,N_9285);
nor U9747 (N_9747,N_7010,N_6452);
or U9748 (N_9748,N_7434,N_7115);
nand U9749 (N_9749,N_8780,N_7336);
nand U9750 (N_9750,N_7766,N_8392);
and U9751 (N_9751,N_7130,N_6730);
and U9752 (N_9752,N_8513,N_8939);
and U9753 (N_9753,N_7073,N_7080);
and U9754 (N_9754,N_7351,N_6402);
nor U9755 (N_9755,N_8393,N_9213);
and U9756 (N_9756,N_6356,N_9126);
nor U9757 (N_9757,N_7135,N_7319);
xor U9758 (N_9758,N_8349,N_8595);
or U9759 (N_9759,N_7745,N_6468);
and U9760 (N_9760,N_9208,N_8649);
nand U9761 (N_9761,N_7281,N_6819);
xor U9762 (N_9762,N_7527,N_6750);
and U9763 (N_9763,N_9181,N_6431);
and U9764 (N_9764,N_8654,N_9265);
or U9765 (N_9765,N_8039,N_7944);
and U9766 (N_9766,N_6436,N_6841);
or U9767 (N_9767,N_7724,N_6920);
or U9768 (N_9768,N_8924,N_9211);
and U9769 (N_9769,N_7209,N_7838);
xor U9770 (N_9770,N_9273,N_8243);
or U9771 (N_9771,N_7549,N_6474);
or U9772 (N_9772,N_8499,N_6256);
nand U9773 (N_9773,N_6834,N_8682);
nor U9774 (N_9774,N_6294,N_9139);
nand U9775 (N_9775,N_8442,N_6557);
and U9776 (N_9776,N_6671,N_6666);
or U9777 (N_9777,N_7496,N_7583);
or U9778 (N_9778,N_8626,N_8689);
or U9779 (N_9779,N_8969,N_7554);
nor U9780 (N_9780,N_6295,N_6688);
and U9781 (N_9781,N_8110,N_6863);
xor U9782 (N_9782,N_8928,N_6799);
nand U9783 (N_9783,N_8136,N_9183);
and U9784 (N_9784,N_7828,N_8164);
and U9785 (N_9785,N_8685,N_6537);
and U9786 (N_9786,N_7296,N_9004);
nand U9787 (N_9787,N_7916,N_6515);
or U9788 (N_9788,N_7888,N_7247);
nand U9789 (N_9789,N_9218,N_6989);
and U9790 (N_9790,N_9360,N_9041);
nand U9791 (N_9791,N_6585,N_7968);
and U9792 (N_9792,N_8702,N_8884);
nand U9793 (N_9793,N_7819,N_9161);
nand U9794 (N_9794,N_7839,N_7669);
and U9795 (N_9795,N_9098,N_8688);
nand U9796 (N_9796,N_8917,N_9186);
or U9797 (N_9797,N_7940,N_9054);
nor U9798 (N_9798,N_8817,N_8209);
nor U9799 (N_9799,N_8090,N_8004);
or U9800 (N_9800,N_6676,N_6406);
or U9801 (N_9801,N_8621,N_7972);
nand U9802 (N_9802,N_9176,N_9344);
or U9803 (N_9803,N_8129,N_9174);
nand U9804 (N_9804,N_8456,N_7444);
nand U9805 (N_9805,N_6619,N_9324);
nor U9806 (N_9806,N_7466,N_8268);
xor U9807 (N_9807,N_8106,N_8105);
or U9808 (N_9808,N_6260,N_6507);
nor U9809 (N_9809,N_8551,N_7899);
nand U9810 (N_9810,N_8698,N_8635);
or U9811 (N_9811,N_8506,N_7974);
xnor U9812 (N_9812,N_8172,N_7187);
or U9813 (N_9813,N_6252,N_7025);
nand U9814 (N_9814,N_6991,N_8326);
nor U9815 (N_9815,N_7960,N_8091);
and U9816 (N_9816,N_7943,N_9362);
nor U9817 (N_9817,N_7238,N_6369);
nor U9818 (N_9818,N_7763,N_7865);
and U9819 (N_9819,N_7589,N_8831);
nor U9820 (N_9820,N_6371,N_8313);
and U9821 (N_9821,N_8252,N_8956);
xnor U9822 (N_9822,N_8063,N_9000);
and U9823 (N_9823,N_8275,N_7330);
xor U9824 (N_9824,N_7965,N_7252);
nor U9825 (N_9825,N_8836,N_8253);
or U9826 (N_9826,N_7606,N_7352);
or U9827 (N_9827,N_7601,N_7049);
or U9828 (N_9828,N_7569,N_7588);
or U9829 (N_9829,N_7845,N_7313);
xor U9830 (N_9830,N_6930,N_9299);
xnor U9831 (N_9831,N_8200,N_8824);
nor U9832 (N_9832,N_7648,N_6743);
nor U9833 (N_9833,N_7457,N_6487);
xor U9834 (N_9834,N_8845,N_8365);
nand U9835 (N_9835,N_8050,N_6838);
nand U9836 (N_9836,N_8057,N_9073);
xnor U9837 (N_9837,N_8696,N_8147);
nor U9838 (N_9838,N_8849,N_6417);
and U9839 (N_9839,N_7266,N_8454);
and U9840 (N_9840,N_6848,N_6258);
nor U9841 (N_9841,N_7453,N_7263);
or U9842 (N_9842,N_8607,N_7894);
nand U9843 (N_9843,N_7937,N_8739);
xor U9844 (N_9844,N_8711,N_6440);
nand U9845 (N_9845,N_8669,N_7925);
nand U9846 (N_9846,N_8850,N_9335);
or U9847 (N_9847,N_7862,N_7616);
nand U9848 (N_9848,N_9120,N_7153);
or U9849 (N_9849,N_7388,N_7582);
nand U9850 (N_9850,N_7604,N_8827);
nand U9851 (N_9851,N_6755,N_8627);
and U9852 (N_9852,N_7047,N_6617);
nor U9853 (N_9853,N_8038,N_7505);
xor U9854 (N_9854,N_8224,N_7881);
and U9855 (N_9855,N_6993,N_8505);
xor U9856 (N_9856,N_8589,N_7734);
nor U9857 (N_9857,N_8985,N_6655);
xnor U9858 (N_9858,N_8420,N_8364);
or U9859 (N_9859,N_8921,N_9318);
and U9860 (N_9860,N_9132,N_8465);
nand U9861 (N_9861,N_7096,N_7764);
nand U9862 (N_9862,N_6664,N_7917);
nand U9863 (N_9863,N_7040,N_8699);
and U9864 (N_9864,N_6587,N_7245);
nor U9865 (N_9865,N_7553,N_6898);
or U9866 (N_9866,N_8645,N_7625);
nor U9867 (N_9867,N_8507,N_6308);
and U9868 (N_9868,N_6372,N_7840);
xnor U9869 (N_9869,N_7159,N_9348);
nor U9870 (N_9870,N_6428,N_7220);
nor U9871 (N_9871,N_7528,N_8975);
xnor U9872 (N_9872,N_8159,N_7659);
or U9873 (N_9873,N_8880,N_6959);
nand U9874 (N_9874,N_8359,N_9283);
nand U9875 (N_9875,N_8988,N_9036);
or U9876 (N_9876,N_6839,N_8941);
and U9877 (N_9877,N_8404,N_7873);
nand U9878 (N_9878,N_7237,N_8059);
nand U9879 (N_9879,N_6422,N_7718);
nor U9880 (N_9880,N_9196,N_8708);
and U9881 (N_9881,N_6780,N_9125);
nand U9882 (N_9882,N_8407,N_9224);
nor U9883 (N_9883,N_6707,N_7106);
and U9884 (N_9884,N_8529,N_9078);
and U9885 (N_9885,N_7020,N_7923);
nand U9886 (N_9886,N_9295,N_6924);
or U9887 (N_9887,N_8088,N_9353);
or U9888 (N_9888,N_7414,N_9010);
xor U9889 (N_9889,N_6495,N_7007);
and U9890 (N_9890,N_8896,N_6362);
or U9891 (N_9891,N_8502,N_8222);
xor U9892 (N_9892,N_6623,N_6867);
nand U9893 (N_9893,N_6348,N_7146);
nor U9894 (N_9894,N_8934,N_6784);
nand U9895 (N_9895,N_7051,N_7129);
nor U9896 (N_9896,N_8932,N_8022);
or U9897 (N_9897,N_7642,N_7386);
or U9898 (N_9898,N_6359,N_6903);
or U9899 (N_9899,N_9227,N_9284);
and U9900 (N_9900,N_8192,N_8524);
and U9901 (N_9901,N_9359,N_8901);
xor U9902 (N_9902,N_7633,N_7979);
xor U9903 (N_9903,N_7297,N_8278);
nand U9904 (N_9904,N_7081,N_7501);
and U9905 (N_9905,N_9235,N_8720);
nand U9906 (N_9906,N_9045,N_9346);
nand U9907 (N_9907,N_8023,N_9066);
xor U9908 (N_9908,N_7078,N_7703);
and U9909 (N_9909,N_6766,N_7456);
and U9910 (N_9910,N_6830,N_8113);
or U9911 (N_9911,N_9187,N_6631);
and U9912 (N_9912,N_8162,N_8891);
and U9913 (N_9913,N_9071,N_6803);
or U9914 (N_9914,N_6328,N_6291);
nor U9915 (N_9915,N_7200,N_8718);
xor U9916 (N_9916,N_6435,N_8721);
and U9917 (N_9917,N_7715,N_7725);
xor U9918 (N_9918,N_7176,N_8479);
and U9919 (N_9919,N_8449,N_6326);
and U9920 (N_9920,N_9113,N_9368);
nor U9921 (N_9921,N_7598,N_9006);
or U9922 (N_9922,N_7379,N_9100);
nor U9923 (N_9923,N_8545,N_6868);
nor U9924 (N_9924,N_8531,N_6472);
nor U9925 (N_9925,N_8274,N_7915);
and U9926 (N_9926,N_7933,N_6719);
or U9927 (N_9927,N_6894,N_7502);
and U9928 (N_9928,N_7216,N_7640);
nand U9929 (N_9929,N_7830,N_6865);
nor U9930 (N_9930,N_9298,N_8299);
and U9931 (N_9931,N_6922,N_8490);
nor U9932 (N_9932,N_7986,N_7389);
nor U9933 (N_9933,N_8847,N_9118);
or U9934 (N_9934,N_8757,N_9327);
nor U9935 (N_9935,N_8044,N_6272);
nand U9936 (N_9936,N_8475,N_7412);
nor U9937 (N_9937,N_7689,N_6885);
nand U9938 (N_9938,N_7948,N_7406);
and U9939 (N_9939,N_9263,N_6559);
and U9940 (N_9940,N_9255,N_7198);
xor U9941 (N_9941,N_6293,N_8869);
nand U9942 (N_9942,N_8321,N_6501);
or U9943 (N_9943,N_9021,N_7100);
or U9944 (N_9944,N_6646,N_6451);
nor U9945 (N_9945,N_6818,N_6446);
and U9946 (N_9946,N_7530,N_6432);
nor U9947 (N_9947,N_6297,N_7124);
nand U9948 (N_9948,N_8146,N_8704);
nand U9949 (N_9949,N_8526,N_8335);
nor U9950 (N_9950,N_7205,N_8525);
nand U9951 (N_9951,N_8355,N_8639);
nand U9952 (N_9952,N_7024,N_7143);
or U9953 (N_9953,N_8512,N_8631);
and U9954 (N_9954,N_8174,N_7860);
and U9955 (N_9955,N_9030,N_8330);
xor U9956 (N_9956,N_7189,N_7900);
nand U9957 (N_9957,N_6857,N_9343);
and U9958 (N_9958,N_8495,N_8279);
and U9959 (N_9959,N_8140,N_7684);
nand U9960 (N_9960,N_9243,N_6921);
nor U9961 (N_9961,N_6394,N_7719);
nand U9962 (N_9962,N_9326,N_7433);
and U9963 (N_9963,N_8103,N_9178);
or U9964 (N_9964,N_7584,N_9116);
nand U9965 (N_9965,N_7112,N_7666);
or U9966 (N_9966,N_7714,N_8189);
nor U9967 (N_9967,N_8436,N_6772);
and U9968 (N_9968,N_6794,N_6496);
and U9969 (N_9969,N_6882,N_8946);
and U9970 (N_9970,N_9079,N_6517);
nor U9971 (N_9971,N_6498,N_9237);
nor U9972 (N_9972,N_7482,N_6400);
and U9973 (N_9973,N_8397,N_8157);
nor U9974 (N_9974,N_8256,N_8646);
nand U9975 (N_9975,N_8353,N_7287);
nor U9976 (N_9976,N_6485,N_7544);
or U9977 (N_9977,N_8244,N_7914);
nand U9978 (N_9978,N_9372,N_7696);
nor U9979 (N_9979,N_9029,N_6641);
nor U9980 (N_9980,N_6336,N_8104);
or U9981 (N_9981,N_8863,N_9354);
xor U9982 (N_9982,N_6828,N_9065);
nand U9983 (N_9983,N_8482,N_7464);
xor U9984 (N_9984,N_6970,N_6917);
or U9985 (N_9985,N_8327,N_7356);
xnor U9986 (N_9986,N_6477,N_9095);
nor U9987 (N_9987,N_7404,N_8491);
nor U9988 (N_9988,N_8373,N_7353);
or U9989 (N_9989,N_7304,N_6941);
nand U9990 (N_9990,N_7011,N_7005);
nor U9991 (N_9991,N_6618,N_7337);
or U9992 (N_9992,N_8651,N_6620);
and U9993 (N_9993,N_6792,N_8722);
nor U9994 (N_9994,N_6445,N_8653);
or U9995 (N_9995,N_7299,N_7021);
or U9996 (N_9996,N_8852,N_9323);
or U9997 (N_9997,N_7375,N_6866);
nand U9998 (N_9998,N_6319,N_9194);
xnor U9999 (N_9999,N_6576,N_8783);
nor U10000 (N_10000,N_8983,N_8322);
or U10001 (N_10001,N_7500,N_7520);
nand U10002 (N_10002,N_8229,N_7118);
xnor U10003 (N_10003,N_6779,N_9229);
nor U10004 (N_10004,N_7184,N_7995);
nor U10005 (N_10005,N_9341,N_8864);
nor U10006 (N_10006,N_6849,N_7074);
nand U10007 (N_10007,N_8811,N_7664);
nor U10008 (N_10008,N_8623,N_8415);
nor U10009 (N_10009,N_6847,N_7826);
and U10010 (N_10010,N_7855,N_6739);
and U10011 (N_10011,N_8984,N_6817);
or U10012 (N_10012,N_7794,N_7614);
and U10013 (N_10013,N_7000,N_8992);
nor U10014 (N_10014,N_6616,N_8759);
xor U10015 (N_10015,N_8666,N_6764);
and U10016 (N_10016,N_6665,N_6663);
nor U10017 (N_10017,N_7532,N_8406);
or U10018 (N_10018,N_8697,N_6599);
or U10019 (N_10019,N_8000,N_9251);
and U10020 (N_10020,N_7720,N_7079);
xor U10021 (N_10021,N_9307,N_7752);
nand U10022 (N_10022,N_6787,N_7730);
nor U10023 (N_10023,N_6516,N_6699);
nor U10024 (N_10024,N_7110,N_6499);
nor U10025 (N_10025,N_6980,N_6628);
nor U10026 (N_10026,N_8045,N_7912);
nor U10027 (N_10027,N_6493,N_6746);
and U10028 (N_10028,N_7889,N_7188);
and U10029 (N_10029,N_8421,N_7006);
nand U10030 (N_10030,N_8911,N_7268);
and U10031 (N_10031,N_8900,N_7597);
nor U10032 (N_10032,N_6405,N_8592);
or U10033 (N_10033,N_8153,N_8637);
nor U10034 (N_10034,N_7849,N_9317);
and U10035 (N_10035,N_8933,N_7836);
and U10036 (N_10036,N_8767,N_7786);
nor U10037 (N_10037,N_6298,N_7243);
xnor U10038 (N_10038,N_9069,N_6540);
nor U10039 (N_10039,N_7909,N_9287);
nor U10040 (N_10040,N_8998,N_7256);
and U10041 (N_10041,N_6717,N_6979);
nor U10042 (N_10042,N_9056,N_8541);
and U10043 (N_10043,N_7107,N_7622);
or U10044 (N_10044,N_6674,N_6883);
xnor U10045 (N_10045,N_8509,N_6492);
or U10046 (N_10046,N_6270,N_6786);
and U10047 (N_10047,N_8405,N_7842);
xor U10048 (N_10048,N_6484,N_9308);
nand U10049 (N_10049,N_9172,N_8591);
or U10050 (N_10050,N_6845,N_7508);
nor U10051 (N_10051,N_8865,N_8223);
nor U10052 (N_10052,N_8731,N_8218);
nand U10053 (N_10053,N_8318,N_9266);
nand U10054 (N_10054,N_6998,N_8497);
and U10055 (N_10055,N_6768,N_9026);
nor U10056 (N_10056,N_7339,N_7160);
and U10057 (N_10057,N_7947,N_7366);
or U10058 (N_10058,N_8168,N_9142);
nor U10059 (N_10059,N_8745,N_8367);
nor U10060 (N_10060,N_6680,N_8938);
or U10061 (N_10061,N_6482,N_6607);
nor U10062 (N_10062,N_8716,N_9231);
and U10063 (N_10063,N_7309,N_8550);
and U10064 (N_10064,N_8014,N_8030);
and U10065 (N_10065,N_8240,N_6805);
nor U10066 (N_10066,N_7387,N_6869);
nand U10067 (N_10067,N_8747,N_7904);
nand U10068 (N_10068,N_8076,N_8606);
nand U10069 (N_10069,N_8674,N_8366);
or U10070 (N_10070,N_6310,N_6669);
or U10071 (N_10071,N_8035,N_8542);
nor U10072 (N_10072,N_7771,N_6465);
nand U10073 (N_10073,N_9105,N_7638);
nand U10074 (N_10074,N_7454,N_8630);
and U10075 (N_10075,N_7782,N_7572);
and U10076 (N_10076,N_7891,N_7744);
nand U10077 (N_10077,N_7951,N_8025);
and U10078 (N_10078,N_8886,N_8403);
nor U10079 (N_10079,N_8641,N_8796);
nand U10080 (N_10080,N_7926,N_7978);
or U10081 (N_10081,N_8979,N_6942);
and U10082 (N_10082,N_7785,N_6678);
nand U10083 (N_10083,N_7936,N_7803);
nand U10084 (N_10084,N_7650,N_6937);
xor U10085 (N_10085,N_6736,N_7599);
nand U10086 (N_10086,N_8856,N_6441);
nand U10087 (N_10087,N_9003,N_7858);
xor U10088 (N_10088,N_7448,N_7704);
nor U10089 (N_10089,N_7834,N_9152);
or U10090 (N_10090,N_7644,N_8336);
or U10091 (N_10091,N_8333,N_7065);
or U10092 (N_10092,N_6522,N_7590);
and U10093 (N_10093,N_8082,N_6837);
nor U10094 (N_10094,N_7799,N_6367);
or U10095 (N_10095,N_8109,N_8680);
or U10096 (N_10096,N_6895,N_6982);
or U10097 (N_10097,N_7778,N_6401);
and U10098 (N_10098,N_6523,N_6833);
nor U10099 (N_10099,N_6423,N_8376);
or U10100 (N_10100,N_7997,N_7668);
xnor U10101 (N_10101,N_6390,N_7790);
and U10102 (N_10102,N_8574,N_9040);
or U10103 (N_10103,N_9270,N_7325);
xnor U10104 (N_10104,N_8937,N_7473);
or U10105 (N_10105,N_7579,N_8923);
and U10106 (N_10106,N_6595,N_6563);
and U10107 (N_10107,N_7095,N_7548);
or U10108 (N_10108,N_9165,N_7594);
or U10109 (N_10109,N_8508,N_7645);
and U10110 (N_10110,N_6950,N_8161);
nand U10111 (N_10111,N_6703,N_6858);
or U10112 (N_10112,N_7210,N_8453);
nor U10113 (N_10113,N_7930,N_7983);
and U10114 (N_10114,N_7634,N_8794);
and U10115 (N_10115,N_7346,N_8272);
or U10116 (N_10116,N_8199,N_8476);
nor U10117 (N_10117,N_8137,N_6654);
nand U10118 (N_10118,N_7935,N_8424);
and U10119 (N_10119,N_8643,N_7156);
and U10120 (N_10120,N_9202,N_6706);
xnor U10121 (N_10121,N_7104,N_7228);
or U10122 (N_10122,N_7804,N_6808);
xnor U10123 (N_10123,N_8712,N_6782);
and U10124 (N_10124,N_8251,N_6977);
nor U10125 (N_10125,N_8143,N_6769);
or U10126 (N_10126,N_8391,N_6364);
nand U10127 (N_10127,N_9070,N_9112);
and U10128 (N_10128,N_9192,N_6800);
nand U10129 (N_10129,N_6360,N_7869);
and U10130 (N_10130,N_8095,N_6612);
or U10131 (N_10131,N_9159,N_6594);
and U10132 (N_10132,N_8019,N_8258);
xor U10133 (N_10133,N_6697,N_8752);
and U10134 (N_10134,N_7165,N_7487);
xor U10135 (N_10135,N_9222,N_9240);
nand U10136 (N_10136,N_8518,N_8763);
nand U10137 (N_10137,N_7770,N_6689);
nor U10138 (N_10138,N_6366,N_8273);
and U10139 (N_10139,N_8608,N_7509);
and U10140 (N_10140,N_8838,N_7223);
nor U10141 (N_10141,N_8603,N_8402);
nor U10142 (N_10142,N_6416,N_6510);
nand U10143 (N_10143,N_8519,N_8461);
nor U10144 (N_10144,N_7646,N_6698);
or U10145 (N_10145,N_7419,N_7576);
nand U10146 (N_10146,N_8537,N_7964);
nor U10147 (N_10147,N_6856,N_7832);
or U10148 (N_10148,N_8510,N_7272);
nor U10149 (N_10149,N_6822,N_9239);
and U10150 (N_10150,N_8580,N_8906);
nor U10151 (N_10151,N_8628,N_6906);
nor U10152 (N_10152,N_8198,N_8051);
nor U10153 (N_10153,N_6600,N_7293);
and U10154 (N_10154,N_9223,N_6434);
nor U10155 (N_10155,N_7057,N_7014);
or U10156 (N_10156,N_6760,N_7447);
nand U10157 (N_10157,N_8970,N_9371);
xor U10158 (N_10158,N_6983,N_7885);
and U10159 (N_10159,N_8480,N_9226);
nor U10160 (N_10160,N_8260,N_9064);
and U10161 (N_10161,N_8750,N_8297);
nor U10162 (N_10162,N_8254,N_8960);
and U10163 (N_10163,N_9124,N_6317);
nand U10164 (N_10164,N_7196,N_7812);
nand U10165 (N_10165,N_7068,N_9158);
nand U10166 (N_10166,N_8776,N_7267);
or U10167 (N_10167,N_6583,N_8918);
or U10168 (N_10168,N_9011,N_7154);
and U10169 (N_10169,N_7893,N_9151);
or U10170 (N_10170,N_7185,N_8277);
and U10171 (N_10171,N_7197,N_8610);
nand U10172 (N_10172,N_8005,N_7027);
nor U10173 (N_10173,N_7955,N_7998);
xor U10174 (N_10174,N_6790,N_8815);
and U10175 (N_10175,N_9320,N_7886);
and U10176 (N_10176,N_6656,N_9051);
or U10177 (N_10177,N_7442,N_6458);
nor U10178 (N_10178,N_6971,N_8210);
nor U10179 (N_10179,N_6586,N_7671);
xnor U10180 (N_10180,N_6373,N_9062);
nor U10181 (N_10181,N_7085,N_6954);
or U10182 (N_10182,N_9007,N_6409);
nor U10183 (N_10183,N_6615,N_7746);
or U10184 (N_10184,N_7788,N_8973);
nand U10185 (N_10185,N_6506,N_6597);
nor U10186 (N_10186,N_7460,N_9342);
nor U10187 (N_10187,N_9082,N_7476);
nor U10188 (N_10188,N_7232,N_7732);
or U10189 (N_10189,N_6826,N_7952);
nor U10190 (N_10190,N_7458,N_6449);
and U10191 (N_10191,N_8290,N_6388);
nand U10192 (N_10192,N_8614,N_8371);
nand U10193 (N_10193,N_8741,N_8221);
nand U10194 (N_10194,N_7284,N_8855);
or U10195 (N_10195,N_7911,N_8820);
nor U10196 (N_10196,N_7631,N_8233);
xor U10197 (N_10197,N_7182,N_7368);
or U10198 (N_10198,N_7170,N_8636);
or U10199 (N_10199,N_7217,N_6387);
nand U10200 (N_10200,N_8665,N_6338);
nand U10201 (N_10201,N_8036,N_7298);
nand U10202 (N_10202,N_7046,N_8416);
xor U10203 (N_10203,N_8190,N_6553);
nand U10204 (N_10204,N_8511,N_7069);
nand U10205 (N_10205,N_8990,N_7251);
nor U10206 (N_10206,N_9276,N_7181);
or U10207 (N_10207,N_6783,N_6886);
nor U10208 (N_10208,N_9333,N_8894);
and U10209 (N_10209,N_8695,N_6709);
or U10210 (N_10210,N_7294,N_8194);
or U10211 (N_10211,N_9328,N_6463);
or U10212 (N_10212,N_7203,N_6810);
nand U10213 (N_10213,N_8919,N_9097);
xnor U10214 (N_10214,N_8239,N_9180);
nor U10215 (N_10215,N_7702,N_8899);
nor U10216 (N_10216,N_8015,N_6324);
xor U10217 (N_10217,N_9329,N_8358);
or U10218 (N_10218,N_8125,N_9128);
nand U10219 (N_10219,N_9091,N_6919);
and U10220 (N_10220,N_9219,N_7680);
or U10221 (N_10221,N_6801,N_6648);
or U10222 (N_10222,N_7168,N_8772);
and U10223 (N_10223,N_9303,N_8068);
or U10224 (N_10224,N_8248,N_8735);
nor U10225 (N_10225,N_7123,N_7102);
or U10226 (N_10226,N_9177,N_7643);
xor U10227 (N_10227,N_7341,N_7275);
nor U10228 (N_10228,N_7514,N_7067);
nand U10229 (N_10229,N_7094,N_7637);
and U10230 (N_10230,N_9146,N_6809);
nor U10231 (N_10231,N_8073,N_7361);
and U10232 (N_10232,N_8195,N_6877);
and U10233 (N_10233,N_7052,N_9072);
nand U10234 (N_10234,N_8851,N_7489);
xnor U10235 (N_10235,N_9043,N_8468);
or U10236 (N_10236,N_6976,N_9115);
xnor U10237 (N_10237,N_6738,N_7498);
nand U10238 (N_10238,N_7229,N_7613);
nor U10239 (N_10239,N_6420,N_8430);
or U10240 (N_10240,N_8363,N_9061);
nor U10241 (N_10241,N_7132,N_8018);
nand U10242 (N_10242,N_8040,N_8343);
xnor U10243 (N_10243,N_6690,N_9157);
and U10244 (N_10244,N_6399,N_9162);
and U10245 (N_10245,N_7455,N_8633);
nor U10246 (N_10246,N_7700,N_8337);
and U10247 (N_10247,N_7029,N_6311);
and U10248 (N_10248,N_6588,N_7259);
and U10249 (N_10249,N_6447,N_7407);
or U10250 (N_10250,N_6907,N_7901);
or U10251 (N_10251,N_6481,N_7013);
or U10252 (N_10252,N_6715,N_7784);
and U10253 (N_10253,N_7847,N_8569);
xor U10254 (N_10254,N_6572,N_6704);
and U10255 (N_10255,N_8766,N_7038);
nor U10256 (N_10256,N_8657,N_9253);
nor U10257 (N_10257,N_7324,N_6604);
nand U10258 (N_10258,N_9109,N_7993);
and U10259 (N_10259,N_8889,N_7494);
and U10260 (N_10260,N_6276,N_7446);
nor U10261 (N_10261,N_8028,N_8431);
nor U10262 (N_10262,N_6683,N_7097);
nand U10263 (N_10263,N_8989,N_6261);
xnor U10264 (N_10264,N_9356,N_9220);
nand U10265 (N_10265,N_8761,N_7813);
nand U10266 (N_10266,N_7317,N_7322);
nor U10267 (N_10267,N_8947,N_8676);
or U10268 (N_10268,N_9150,N_7701);
nand U10269 (N_10269,N_8931,N_9123);
or U10270 (N_10270,N_8285,N_9058);
and U10271 (N_10271,N_8417,N_6335);
or U10272 (N_10272,N_8488,N_8009);
nand U10273 (N_10273,N_6389,N_6626);
and U10274 (N_10274,N_8400,N_6901);
nor U10275 (N_10275,N_9256,N_7092);
nand U10276 (N_10276,N_7398,N_9203);
xnor U10277 (N_10277,N_7307,N_8909);
and U10278 (N_10278,N_8419,N_8514);
or U10279 (N_10279,N_6460,N_7971);
and U10280 (N_10280,N_7365,N_7109);
xor U10281 (N_10281,N_7003,N_6632);
nand U10282 (N_10282,N_8520,N_8528);
xnor U10283 (N_10283,N_9137,N_6486);
or U10284 (N_10284,N_9358,N_6573);
or U10285 (N_10285,N_8746,N_6490);
nand U10286 (N_10286,N_8156,N_8267);
nor U10287 (N_10287,N_7883,N_7201);
nor U10288 (N_10288,N_9302,N_7373);
and U10289 (N_10289,N_6306,N_7098);
nor U10290 (N_10290,N_6997,N_9321);
and U10291 (N_10291,N_7179,N_8385);
and U10292 (N_10292,N_7980,N_9338);
and U10293 (N_10293,N_8242,N_9184);
nor U10294 (N_10294,N_7529,N_6948);
nand U10295 (N_10295,N_7043,N_8756);
nand U10296 (N_10296,N_8629,N_6343);
nand U10297 (N_10297,N_7762,N_6714);
or U10298 (N_10298,N_7626,N_7882);
xor U10299 (N_10299,N_7166,N_7491);
nand U10300 (N_10300,N_7681,N_7988);
nand U10301 (N_10301,N_8549,N_6374);
nand U10302 (N_10302,N_9037,N_7410);
and U10303 (N_10303,N_8351,N_6288);
nor U10304 (N_10304,N_7585,N_9057);
nand U10305 (N_10305,N_6759,N_7333);
nor U10306 (N_10306,N_7417,N_8232);
nor U10307 (N_10307,N_6835,N_9093);
and U10308 (N_10308,N_6386,N_8346);
nor U10309 (N_10309,N_9094,N_6309);
nor U10310 (N_10310,N_7172,N_8620);
and U10311 (N_10311,N_8270,N_7690);
or U10312 (N_10312,N_8662,N_6891);
nor U10313 (N_10313,N_8807,N_6491);
nor U10314 (N_10314,N_6286,N_7355);
and U10315 (N_10315,N_6622,N_6875);
or U10316 (N_10316,N_8160,N_7462);
and U10317 (N_10317,N_6592,N_9154);
and U10318 (N_10318,N_8823,N_6526);
nand U10319 (N_10319,N_7063,N_6413);
nand U10320 (N_10320,N_8570,N_7199);
and U10321 (N_10321,N_7315,N_7765);
or U10322 (N_10322,N_7918,N_8126);
nor U10323 (N_10323,N_8071,N_7316);
and U10324 (N_10324,N_7994,N_8049);
or U10325 (N_10325,N_7890,N_8805);
nand U10326 (N_10326,N_7927,N_7518);
and U10327 (N_10327,N_6395,N_7077);
nor U10328 (N_10328,N_7876,N_6829);
nand U10329 (N_10329,N_7987,N_7818);
and U10330 (N_10330,N_7045,N_9373);
nor U10331 (N_10331,N_8466,N_6972);
and U10332 (N_10332,N_8521,N_6292);
xor U10333 (N_10333,N_8007,N_8910);
or U10334 (N_10334,N_8425,N_8165);
nand U10335 (N_10335,N_6345,N_6613);
and U10336 (N_10336,N_7321,N_6548);
nor U10337 (N_10337,N_8317,N_6964);
or U10338 (N_10338,N_7898,N_8644);
or U10339 (N_10339,N_7610,N_7285);
nor U10340 (N_10340,N_7405,N_8361);
nand U10341 (N_10341,N_6511,N_8926);
or U10342 (N_10342,N_9170,N_8409);
nor U10343 (N_10343,N_9244,N_8448);
and U10344 (N_10344,N_6302,N_8139);
nor U10345 (N_10345,N_9025,N_7479);
xnor U10346 (N_10346,N_8809,N_8483);
nand U10347 (N_10347,N_6398,N_7202);
nor U10348 (N_10348,N_8435,N_6547);
nor U10349 (N_10349,N_8150,N_8197);
nand U10350 (N_10350,N_8357,N_7206);
nor U10351 (N_10351,N_8309,N_6742);
or U10352 (N_10352,N_8445,N_7905);
and U10353 (N_10353,N_8804,N_8797);
or U10354 (N_10354,N_8749,N_7880);
nor U10355 (N_10355,N_6427,N_8660);
nor U10356 (N_10356,N_6603,N_7657);
nor U10357 (N_10357,N_7575,N_8176);
nand U10358 (N_10358,N_7415,N_8875);
and U10359 (N_10359,N_6973,N_6731);
nand U10360 (N_10360,N_8167,N_6692);
and U10361 (N_10361,N_6927,N_8681);
or U10362 (N_10362,N_7655,N_6314);
and U10363 (N_10363,N_8398,N_7857);
and U10364 (N_10364,N_7164,N_9042);
and U10365 (N_10365,N_7326,N_8447);
or U10366 (N_10366,N_8433,N_6967);
and U10367 (N_10367,N_7843,N_8181);
nor U10368 (N_10368,N_6580,N_9068);
nand U10369 (N_10369,N_8356,N_7218);
and U10370 (N_10370,N_9155,N_8148);
nand U10371 (N_10371,N_9083,N_8115);
or U10372 (N_10372,N_7440,N_8559);
and U10373 (N_10373,N_6407,N_7739);
nor U10374 (N_10374,N_7378,N_6682);
and U10375 (N_10375,N_8043,N_7042);
and U10376 (N_10376,N_6914,N_6313);
nand U10377 (N_10377,N_6438,N_6264);
nand U10378 (N_10378,N_8077,N_8501);
nand U10379 (N_10379,N_8868,N_6702);
nor U10380 (N_10380,N_7088,N_7279);
or U10381 (N_10381,N_6470,N_9060);
nand U10382 (N_10382,N_8616,N_6514);
or U10383 (N_10383,N_8427,N_9315);
nand U10384 (N_10384,N_8867,N_8730);
or U10385 (N_10385,N_7474,N_9048);
and U10386 (N_10386,N_9140,N_6733);
nand U10387 (N_10387,N_9374,N_7485);
nand U10388 (N_10388,N_8876,N_8798);
nand U10389 (N_10389,N_9185,N_7192);
nand U10390 (N_10390,N_8149,N_9044);
xor U10391 (N_10391,N_6986,N_6814);
and U10392 (N_10392,N_8329,N_6289);
nor U10393 (N_10393,N_8265,N_6899);
nand U10394 (N_10394,N_7177,N_7152);
and U10395 (N_10395,N_8173,N_7550);
or U10396 (N_10396,N_8557,N_6269);
and U10397 (N_10397,N_9232,N_7833);
and U10398 (N_10398,N_9086,N_8381);
or U10399 (N_10399,N_6591,N_8950);
and U10400 (N_10400,N_6694,N_8964);
and U10401 (N_10401,N_8231,N_7030);
and U10402 (N_10402,N_7661,N_9027);
and U10403 (N_10403,N_8287,N_7780);
nand U10404 (N_10404,N_9210,N_8732);
nor U10405 (N_10405,N_6939,N_7241);
or U10406 (N_10406,N_7556,N_8032);
and U10407 (N_10407,N_6564,N_8089);
and U10408 (N_10408,N_6304,N_6598);
nand U10409 (N_10409,N_8305,N_9190);
xor U10410 (N_10410,N_9008,N_8099);
and U10411 (N_10411,N_9332,N_7418);
nand U10412 (N_10412,N_8874,N_8810);
nor U10413 (N_10413,N_6881,N_8860);
nand U10414 (N_10414,N_9135,N_8828);
or U10415 (N_10415,N_6807,N_8920);
nand U10416 (N_10416,N_8744,N_7111);
nor U10417 (N_10417,N_6726,N_7331);
nor U10418 (N_10418,N_8587,N_6916);
or U10419 (N_10419,N_9138,N_7934);
nand U10420 (N_10420,N_9288,N_8842);
or U10421 (N_10421,N_8311,N_6381);
nor U10422 (N_10422,N_9352,N_6403);
xnor U10423 (N_10423,N_6346,N_8208);
nor U10424 (N_10424,N_6860,N_9337);
or U10425 (N_10425,N_7015,N_6303);
nand U10426 (N_10426,N_8006,N_8781);
nor U10427 (N_10427,N_6996,N_7591);
nor U10428 (N_10428,N_6963,N_8535);
nand U10429 (N_10429,N_8962,N_7310);
nor U10430 (N_10430,N_8295,N_9228);
and U10431 (N_10431,N_8706,N_8108);
nand U10432 (N_10432,N_7800,N_8995);
nor U10433 (N_10433,N_7777,N_9200);
or U10434 (N_10434,N_8011,N_7041);
or U10435 (N_10435,N_7507,N_9156);
and U10436 (N_10436,N_8185,N_6672);
or U10437 (N_10437,N_7409,N_8257);
nand U10438 (N_10438,N_7654,N_6483);
or U10439 (N_10439,N_7370,N_7376);
or U10440 (N_10440,N_7117,N_8834);
nor U10441 (N_10441,N_6778,N_6691);
xor U10442 (N_10442,N_8261,N_7856);
and U10443 (N_10443,N_8652,N_7180);
or U10444 (N_10444,N_6601,N_9366);
nor U10445 (N_10445,N_9319,N_8467);
and U10446 (N_10446,N_8092,N_7503);
nor U10447 (N_10447,N_6645,N_7265);
nor U10448 (N_10448,N_7303,N_7076);
nor U10449 (N_10449,N_7305,N_7036);
nor U10450 (N_10450,N_7796,N_7729);
or U10451 (N_10451,N_7693,N_6307);
xnor U10452 (N_10452,N_8659,N_7128);
nor U10453 (N_10453,N_6798,N_6602);
nor U10454 (N_10454,N_6545,N_8134);
nand U10455 (N_10455,N_9014,N_7438);
or U10456 (N_10456,N_7053,N_6287);
nor U10457 (N_10457,N_8813,N_8987);
nand U10458 (N_10458,N_8760,N_8284);
or U10459 (N_10459,N_6892,N_6566);
nor U10460 (N_10460,N_6934,N_7754);
nand U10461 (N_10461,N_7291,N_7357);
and U10462 (N_10462,N_8310,N_8967);
nor U10463 (N_10463,N_8383,N_9012);
and U10464 (N_10464,N_7125,N_6480);
and U10465 (N_10465,N_8613,N_8881);
nor U10466 (N_10466,N_7811,N_6253);
and U10467 (N_10467,N_7985,N_8413);
nand U10468 (N_10468,N_6908,N_8694);
and U10469 (N_10469,N_8180,N_9147);
or U10470 (N_10470,N_8307,N_6582);
or U10471 (N_10471,N_8814,N_7519);
nand U10472 (N_10472,N_7524,N_9259);
nor U10473 (N_10473,N_8952,N_8778);
nor U10474 (N_10474,N_6705,N_8369);
xnor U10475 (N_10475,N_8762,N_8196);
nor U10476 (N_10476,N_9355,N_7465);
nand U10477 (N_10477,N_8152,N_8957);
nand U10478 (N_10478,N_9241,N_9197);
xor U10479 (N_10479,N_7682,N_6575);
nand U10480 (N_10480,N_6478,N_7949);
or U10481 (N_10481,N_8228,N_8135);
or U10482 (N_10482,N_7656,N_8054);
and U10483 (N_10483,N_6277,N_7787);
nor U10484 (N_10484,N_6851,N_8069);
xnor U10485 (N_10485,N_7233,N_7673);
and U10486 (N_10486,N_9347,N_7054);
xor U10487 (N_10487,N_8348,N_7371);
or U10488 (N_10488,N_6637,N_6765);
xor U10489 (N_10489,N_7781,N_8554);
or U10490 (N_10490,N_6554,N_6796);
or U10491 (N_10491,N_7062,N_6827);
and U10492 (N_10492,N_8074,N_9002);
and U10493 (N_10493,N_8138,N_7225);
or U10494 (N_10494,N_7938,N_8588);
nand U10495 (N_10495,N_7969,N_6419);
and U10496 (N_10496,N_7158,N_8280);
xnor U10497 (N_10497,N_9074,N_7967);
and U10498 (N_10498,N_6539,N_7213);
or U10499 (N_10499,N_6325,N_8354);
xor U10500 (N_10500,N_9250,N_7493);
nand U10501 (N_10501,N_7670,N_7574);
nand U10502 (N_10502,N_8292,N_7698);
and U10503 (N_10503,N_9106,N_6418);
and U10504 (N_10504,N_8477,N_8615);
or U10505 (N_10505,N_8543,N_7348);
or U10506 (N_10506,N_6949,N_8120);
or U10507 (N_10507,N_6668,N_9293);
nor U10508 (N_10508,N_6853,N_6383);
nand U10509 (N_10509,N_8955,N_7555);
xnor U10510 (N_10510,N_6855,N_7174);
or U10511 (N_10511,N_8186,N_9092);
or U10512 (N_10512,N_6735,N_8617);
nor U10513 (N_10513,N_8169,N_9314);
and U10514 (N_10514,N_8055,N_8214);
or U10515 (N_10515,N_8121,N_8236);
and U10516 (N_10516,N_7048,N_7558);
and U10517 (N_10517,N_7411,N_6368);
nor U10518 (N_10518,N_6430,N_6410);
nand U10519 (N_10519,N_7009,N_9339);
nand U10520 (N_10520,N_8533,N_8255);
or U10521 (N_10521,N_8779,N_7758);
and U10522 (N_10522,N_6754,N_6377);
and U10523 (N_10523,N_6693,N_8516);
or U10524 (N_10524,N_7573,N_6677);
nor U10525 (N_10525,N_7311,N_7103);
xor U10526 (N_10526,N_8332,N_7814);
nor U10527 (N_10527,N_6880,N_7578);
or U10528 (N_10528,N_8602,N_6748);
nand U10529 (N_10529,N_8980,N_8331);
or U10530 (N_10530,N_6923,N_8017);
or U10531 (N_10531,N_7868,N_8282);
nand U10532 (N_10532,N_7736,N_9024);
nor U10533 (N_10533,N_9047,N_6744);
nand U10534 (N_10534,N_8661,N_9300);
nand U10535 (N_10535,N_6994,N_6946);
or U10536 (N_10536,N_8556,N_8552);
or U10537 (N_10537,N_7560,N_8072);
nand U10538 (N_10538,N_6450,N_6936);
and U10539 (N_10539,N_8296,N_6957);
and U10540 (N_10540,N_6375,N_7629);
or U10541 (N_10541,N_7018,N_7292);
nor U10542 (N_10542,N_7451,N_6382);
nor U10543 (N_10543,N_8728,N_8060);
nand U10544 (N_10544,N_6259,N_8940);
nor U10545 (N_10545,N_8230,N_6629);
nand U10546 (N_10546,N_8784,N_6721);
or U10547 (N_10547,N_8816,N_6280);
xor U10548 (N_10548,N_8438,N_6263);
nor U10549 (N_10549,N_7975,N_6978);
nand U10550 (N_10550,N_8771,N_6852);
nand U10551 (N_10551,N_7139,N_7981);
or U10552 (N_10552,N_8723,N_7059);
or U10553 (N_10553,N_6802,N_7939);
nor U10554 (N_10554,N_8713,N_6497);
and U10555 (N_10555,N_9242,N_8504);
or U10556 (N_10556,N_6938,N_8184);
nor U10557 (N_10557,N_9258,N_8601);
nor U10558 (N_10558,N_7861,N_9289);
xor U10559 (N_10559,N_7126,N_8897);
or U10560 (N_10560,N_9245,N_9148);
or U10561 (N_10561,N_6426,N_6862);
and U10562 (N_10562,N_8858,N_9175);
nor U10563 (N_10563,N_6334,N_6650);
and U10564 (N_10564,N_8003,N_8675);
xnor U10565 (N_10565,N_7239,N_8387);
nand U10566 (N_10566,N_8822,N_8801);
or U10567 (N_10567,N_7945,N_8830);
nor U10568 (N_10568,N_6323,N_6380);
and U10569 (N_10569,N_7422,N_6657);
and U10570 (N_10570,N_8081,N_7678);
nand U10571 (N_10571,N_6611,N_8142);
nor U10572 (N_10572,N_8764,N_9334);
xor U10573 (N_10573,N_7942,N_7953);
or U10574 (N_10574,N_7907,N_7327);
nand U10575 (N_10575,N_7820,N_6278);
nand U10576 (N_10576,N_7775,N_8002);
nor U10577 (N_10577,N_7941,N_7144);
or U10578 (N_10578,N_7991,N_9168);
or U10579 (N_10579,N_6536,N_7977);
xnor U10580 (N_10580,N_6874,N_7635);
nor U10581 (N_10581,N_7756,N_8437);
or U10582 (N_10582,N_8158,N_6577);
nor U10583 (N_10583,N_6985,N_8463);
and U10584 (N_10584,N_9349,N_7244);
and U10585 (N_10585,N_7513,N_7131);
xor U10586 (N_10586,N_7219,N_8966);
xnor U10587 (N_10587,N_9279,N_9262);
and U10588 (N_10588,N_7511,N_9153);
or U10589 (N_10589,N_9193,N_8854);
nor U10590 (N_10590,N_7432,N_8344);
nand U10591 (N_10591,N_6832,N_8128);
or U10592 (N_10592,N_7872,N_8902);
or U10593 (N_10593,N_7329,N_6652);
xor U10594 (N_10594,N_6644,N_6753);
and U10595 (N_10595,N_7962,N_7844);
nor U10596 (N_10596,N_7358,N_8320);
or U10597 (N_10597,N_6546,N_7755);
xnor U10598 (N_10598,N_6966,N_8584);
or U10599 (N_10599,N_6661,N_7630);
nor U10600 (N_10600,N_8029,N_8596);
nor U10601 (N_10601,N_8640,N_7391);
or U10602 (N_10602,N_8234,N_7603);
and U10603 (N_10603,N_6888,N_8300);
nand U10604 (N_10604,N_6928,N_7133);
nor U10605 (N_10605,N_7517,N_7257);
and U10606 (N_10606,N_7161,N_7484);
or U10607 (N_10607,N_6518,N_6333);
and U10608 (N_10608,N_7672,N_7557);
and U10609 (N_10609,N_6296,N_6951);
nor U10610 (N_10610,N_6342,N_8579);
nor U10611 (N_10611,N_6897,N_7835);
or U10612 (N_10612,N_7091,N_7892);
nor U10613 (N_10613,N_7459,N_8116);
and U10614 (N_10614,N_6718,N_8021);
and U10615 (N_10615,N_7581,N_8084);
and U10616 (N_10616,N_7641,N_8216);
nor U10617 (N_10617,N_6974,N_8141);
nor U10618 (N_10618,N_7984,N_8879);
nand U10619 (N_10619,N_8500,N_9204);
and U10620 (N_10620,N_6815,N_8773);
xnor U10621 (N_10621,N_7602,N_8117);
and U10622 (N_10622,N_8936,N_8306);
and U10623 (N_10623,N_7748,N_6635);
or U10624 (N_10624,N_6670,N_7541);
nor U10625 (N_10625,N_8119,N_8399);
and U10626 (N_10626,N_6318,N_6824);
nor U10627 (N_10627,N_6589,N_6961);
or U10628 (N_10628,N_9275,N_7061);
or U10629 (N_10629,N_7190,N_7815);
xnor U10630 (N_10630,N_6412,N_8929);
nor U10631 (N_10631,N_8678,N_6544);
and U10632 (N_10632,N_8315,N_7381);
nand U10633 (N_10633,N_6732,N_8895);
and U10634 (N_10634,N_8291,N_8622);
and U10635 (N_10635,N_6361,N_7214);
nor U10636 (N_10636,N_7396,N_7277);
nor U10637 (N_10637,N_8065,N_8600);
nor U10638 (N_10638,N_7022,N_8903);
and U10639 (N_10639,N_7191,N_8473);
and U10640 (N_10640,N_6391,N_7283);
nand U10641 (N_10641,N_8386,N_7692);
or U10642 (N_10642,N_6902,N_6425);
nand U10643 (N_10643,N_7908,N_8246);
or U10644 (N_10644,N_7809,N_7534);
and U10645 (N_10645,N_7147,N_8215);
and U10646 (N_10646,N_6257,N_6944);
xnor U10647 (N_10647,N_6791,N_7609);
nor U10648 (N_10648,N_7429,N_6909);
or U10649 (N_10649,N_7961,N_6630);
xnor U10650 (N_10650,N_7721,N_7064);
or U10651 (N_10651,N_7050,N_8670);
and U10652 (N_10652,N_6984,N_7592);
nand U10653 (N_10653,N_8101,N_8293);
and U10654 (N_10654,N_7002,N_8737);
nor U10655 (N_10655,N_8818,N_8008);
or U10656 (N_10656,N_7226,N_8098);
nand U10657 (N_10657,N_8408,N_6762);
or U10658 (N_10658,N_8334,N_8080);
nand U10659 (N_10659,N_8560,N_9019);
nor U10660 (N_10660,N_8487,N_8575);
nand U10661 (N_10661,N_6322,N_6365);
and U10662 (N_10662,N_7060,N_7966);
and U10663 (N_10663,N_7155,N_8701);
nand U10664 (N_10664,N_8844,N_8671);
or U10665 (N_10665,N_8803,N_8375);
nand U10666 (N_10666,N_6551,N_9306);
xor U10667 (N_10667,N_7083,N_8997);
nor U10668 (N_10668,N_7463,N_8832);
nor U10669 (N_10669,N_6254,N_8053);
nor U10670 (N_10670,N_8667,N_7792);
nor U10671 (N_10671,N_6528,N_8175);
xor U10672 (N_10672,N_8664,N_6773);
or U10673 (N_10673,N_7568,N_7385);
nor U10674 (N_10674,N_7416,N_8220);
or U10675 (N_10675,N_6271,N_8472);
nor U10676 (N_10676,N_7791,N_7850);
nand U10677 (N_10677,N_7829,N_7649);
and U10678 (N_10678,N_7340,N_6558);
xnor U10679 (N_10679,N_9114,N_8904);
or U10680 (N_10680,N_8441,N_8325);
nand U10681 (N_10681,N_6992,N_7260);
or U10682 (N_10682,N_8993,N_8390);
or U10683 (N_10683,N_8249,N_7697);
nor U10684 (N_10684,N_7439,N_7827);
or U10685 (N_10685,N_8871,N_8787);
and U10686 (N_10686,N_9001,N_8450);
nor U10687 (N_10687,N_8033,N_8677);
or U10688 (N_10688,N_7653,N_8994);
or U10689 (N_10689,N_9173,N_6542);
nand U10690 (N_10690,N_8734,N_7016);
and U10691 (N_10691,N_7647,N_6352);
or U10692 (N_10692,N_6512,N_6624);
nor U10693 (N_10693,N_7497,N_9028);
or U10694 (N_10694,N_7343,N_6524);
nand U10695 (N_10695,N_6301,N_8710);
and U10696 (N_10696,N_8953,N_7012);
or U10697 (N_10697,N_7566,N_8079);
and U10698 (N_10698,N_7561,N_9191);
nor U10699 (N_10699,N_7932,N_7651);
nor U10700 (N_10700,N_7617,N_8927);
nand U10701 (N_10701,N_8839,N_7167);
nor U10702 (N_10702,N_6476,N_6363);
and U10703 (N_10703,N_8034,N_8555);
nand U10704 (N_10704,N_7846,N_7384);
nor U10705 (N_10705,N_8709,N_8754);
or U10706 (N_10706,N_7475,N_6816);
nand U10707 (N_10707,N_7377,N_7035);
or U10708 (N_10708,N_6889,N_6911);
or U10709 (N_10709,N_7896,N_6701);
nand U10710 (N_10710,N_7767,N_6660);
and U10711 (N_10711,N_7468,N_7837);
and U10712 (N_10712,N_7887,N_9108);
nand U10713 (N_10713,N_6341,N_7652);
nor U10714 (N_10714,N_6283,N_6878);
or U10715 (N_10715,N_6437,N_8247);
or U10716 (N_10716,N_7235,N_7723);
nor U10717 (N_10717,N_8751,N_6713);
nor U10718 (N_10718,N_8700,N_8719);
and U10719 (N_10719,N_8972,N_8187);
nor U10720 (N_10720,N_9018,N_7249);
or U10721 (N_10721,N_6266,N_7679);
nand U10722 (N_10722,N_8235,N_7058);
nand U10723 (N_10723,N_6593,N_7212);
or U10724 (N_10724,N_6444,N_7810);
and U10725 (N_10725,N_8945,N_8308);
nand U10726 (N_10726,N_7382,N_6929);
xnor U10727 (N_10727,N_9280,N_9063);
or U10728 (N_10728,N_7392,N_9130);
or U10729 (N_10729,N_6653,N_7424);
nand U10730 (N_10730,N_6915,N_8609);
and U10731 (N_10731,N_8748,N_8586);
nor U10732 (N_10732,N_8733,N_9188);
nor U10733 (N_10733,N_8485,N_7072);
or U10734 (N_10734,N_8001,N_8434);
or U10735 (N_10735,N_8976,N_7403);
nor U10736 (N_10736,N_6408,N_7004);
and U10737 (N_10737,N_7254,N_8411);
and U10738 (N_10738,N_9076,N_6312);
and U10739 (N_10739,N_8418,N_6890);
nand U10740 (N_10740,N_8262,N_9225);
nor U10741 (N_10741,N_7032,N_9119);
nor U10742 (N_10742,N_6455,N_8597);
or U10743 (N_10743,N_7395,N_6552);
nand U10744 (N_10744,N_6638,N_8100);
nor U10745 (N_10745,N_7264,N_7467);
nand U10746 (N_10746,N_8565,N_8996);
nor U10747 (N_10747,N_6658,N_6884);
nor U10748 (N_10748,N_9260,N_7552);
nor U10749 (N_10749,N_8786,N_8743);
and U10750 (N_10750,N_8245,N_7044);
and U10751 (N_10751,N_6442,N_7950);
nand U10752 (N_10752,N_7895,N_9067);
or U10753 (N_10753,N_6711,N_7421);
nor U10754 (N_10754,N_6457,N_7430);
or U10755 (N_10755,N_8942,N_8075);
or U10756 (N_10756,N_7363,N_7976);
nand U10757 (N_10757,N_7242,N_8785);
or U10758 (N_10758,N_7694,N_8768);
nand U10759 (N_10759,N_8037,N_8656);
nor U10760 (N_10760,N_8093,N_9034);
nor U10761 (N_10761,N_9167,N_8304);
nor U10762 (N_10762,N_8714,N_6953);
or U10763 (N_10763,N_7848,N_6625);
and U10764 (N_10764,N_9294,N_9038);
or U10765 (N_10765,N_7738,N_6532);
nand U10766 (N_10766,N_8833,N_6456);
and U10767 (N_10767,N_7522,N_8276);
and U10768 (N_10768,N_8378,N_7477);
nor U10769 (N_10769,N_7757,N_7017);
nor U10770 (N_10770,N_8826,N_6569);
or U10771 (N_10771,N_7071,N_8576);
xnor U10772 (N_10772,N_7449,N_8687);
xor U10773 (N_10773,N_7551,N_6255);
nor U10774 (N_10774,N_7423,N_6918);
and U10775 (N_10775,N_9075,N_7772);
nand U10776 (N_10776,N_7677,N_7121);
xnor U10777 (N_10777,N_8503,N_8481);
or U10778 (N_10778,N_8740,N_7546);
nand U10779 (N_10779,N_6534,N_8203);
nor U10780 (N_10780,N_8944,N_7105);
nor U10781 (N_10781,N_8658,N_8625);
nor U10782 (N_10782,N_8237,N_9101);
nand U10783 (N_10783,N_8201,N_6940);
or U10784 (N_10784,N_9264,N_7360);
or U10785 (N_10785,N_7471,N_7807);
nand U10786 (N_10786,N_6905,N_9274);
nand U10787 (N_10787,N_8532,N_7269);
and U10788 (N_10788,N_9336,N_6962);
and U10789 (N_10789,N_7586,N_6502);
nand U10790 (N_10790,N_8612,N_7806);
or U10791 (N_10791,N_9080,N_8925);
nand U10792 (N_10792,N_6433,N_6710);
nor U10793 (N_10793,N_7959,N_9149);
or U10794 (N_10794,N_8683,N_6443);
nand U10795 (N_10795,N_6756,N_9252);
nor U10796 (N_10796,N_7399,N_8401);
nor U10797 (N_10797,N_7328,N_9345);
and U10798 (N_10798,N_7728,N_7193);
and U10799 (N_10799,N_6332,N_8571);
or U10800 (N_10800,N_6503,N_9198);
nand U10801 (N_10801,N_7801,N_7821);
or U10802 (N_10802,N_9169,N_7262);
nor U10803 (N_10803,N_7142,N_6932);
and U10804 (N_10804,N_9104,N_9291);
nor U10805 (N_10805,N_9267,N_7864);
and U10806 (N_10806,N_8963,N_7870);
or U10807 (N_10807,N_6912,N_8207);
nand U10808 (N_10808,N_7282,N_9301);
or U10809 (N_10809,N_7537,N_9325);
xnor U10810 (N_10810,N_7920,N_6767);
nand U10811 (N_10811,N_8042,N_7086);
xnor U10812 (N_10812,N_8650,N_8478);
or U10813 (N_10813,N_8339,N_8047);
nand U10814 (N_10814,N_6812,N_7853);
or U10815 (N_10815,N_8016,N_7114);
xnor U10816 (N_10816,N_7562,N_8020);
or U10817 (N_10817,N_8460,N_8227);
xor U10818 (N_10818,N_6555,N_6945);
xor U10819 (N_10819,N_8578,N_7445);
nor U10820 (N_10820,N_6686,N_8289);
nor U10821 (N_10821,N_7675,N_8770);
or U10822 (N_10822,N_8238,N_7420);
xor U10823 (N_10823,N_8154,N_6379);
nor U10824 (N_10824,N_7717,N_7138);
nor U10825 (N_10825,N_7854,N_8789);
and U10826 (N_10826,N_7246,N_6776);
nor U10827 (N_10827,N_6354,N_8599);
and U10828 (N_10828,N_7150,N_8410);
or U10829 (N_10829,N_8878,N_9286);
or U10830 (N_10830,N_8340,N_7516);
nor U10831 (N_10831,N_7543,N_8755);
nand U10832 (N_10832,N_8041,N_7627);
and U10833 (N_10833,N_7605,N_7687);
and U10834 (N_10834,N_9361,N_7731);
nor U10835 (N_10835,N_6771,N_8213);
nand U10836 (N_10836,N_6509,N_8915);
nor U10837 (N_10837,N_8829,N_6282);
or U10838 (N_10838,N_7342,N_8642);
and U10839 (N_10839,N_6910,N_6659);
nor U10840 (N_10840,N_8686,N_8259);
nor U10841 (N_10841,N_9309,N_7116);
and U10842 (N_10842,N_8226,N_6843);
and U10843 (N_10843,N_6844,N_8342);
or U10844 (N_10844,N_8898,N_6651);
and U10845 (N_10845,N_9331,N_6958);
and U10846 (N_10846,N_6793,N_7737);
xnor U10847 (N_10847,N_7026,N_6893);
and U10848 (N_10848,N_8298,N_6999);
and U10849 (N_10849,N_8548,N_6339);
nor U10850 (N_10850,N_8793,N_8951);
and U10851 (N_10851,N_7587,N_8991);
and U10852 (N_10852,N_6329,N_7492);
or U10853 (N_10853,N_8539,N_7695);
or U10854 (N_10854,N_9059,N_6584);
nor U10855 (N_10855,N_7982,N_8202);
nor U10856 (N_10856,N_8530,N_7699);
or U10857 (N_10857,N_6687,N_8127);
and U10858 (N_10858,N_7596,N_6636);
and U10859 (N_10859,N_6960,N_6614);
nor U10860 (N_10860,N_7877,N_8345);
or U10861 (N_10861,N_8062,N_8388);
or U10862 (N_10862,N_6870,N_7547);
nand U10863 (N_10863,N_6357,N_6854);
or U10864 (N_10864,N_6527,N_7866);
nor U10865 (N_10865,N_8171,N_9052);
or U10866 (N_10866,N_9282,N_7194);
nand U10867 (N_10867,N_8469,N_7711);
nor U10868 (N_10868,N_6505,N_8066);
or U10869 (N_10869,N_7469,N_8647);
and U10870 (N_10870,N_9053,N_7753);
nand U10871 (N_10871,N_8703,N_7227);
nand U10872 (N_10872,N_8206,N_6775);
and U10873 (N_10873,N_7222,N_8726);
or U10874 (N_10874,N_7334,N_9212);
or U10875 (N_10875,N_8812,N_8396);
xor U10876 (N_10876,N_7320,N_9141);
xor U10877 (N_10877,N_8178,N_8982);
nor U10878 (N_10878,N_6675,N_7427);
nand U10879 (N_10879,N_6454,N_7271);
nor U10880 (N_10880,N_6879,N_7108);
or U10881 (N_10881,N_6353,N_8690);
or U10882 (N_10882,N_8914,N_7773);
nor U10883 (N_10883,N_6679,N_8286);
nand U10884 (N_10884,N_7716,N_6279);
nand U10885 (N_10885,N_9131,N_8668);
and U10886 (N_10886,N_6876,N_7992);
and U10887 (N_10887,N_7999,N_8707);
or U10888 (N_10888,N_8462,N_6421);
nand U10889 (N_10889,N_6385,N_6429);
or U10890 (N_10890,N_8913,N_7831);
and U10891 (N_10891,N_8439,N_7480);
or U10892 (N_10892,N_7816,N_8605);
or U10893 (N_10893,N_6448,N_7897);
nand U10894 (N_10894,N_6608,N_7300);
nor U10895 (N_10895,N_8166,N_8873);
nor U10896 (N_10896,N_7082,N_7075);
nand U10897 (N_10897,N_7148,N_8971);
nand U10898 (N_10898,N_7538,N_9217);
xor U10899 (N_10899,N_6535,N_6300);
and U10900 (N_10900,N_9236,N_9136);
or U10901 (N_10901,N_7624,N_8566);
or U10902 (N_10902,N_8031,N_7278);
and U10903 (N_10903,N_8085,N_6479);
and U10904 (N_10904,N_9269,N_9351);
or U10905 (N_10905,N_7817,N_7996);
or U10906 (N_10906,N_7332,N_7957);
nand U10907 (N_10907,N_8446,N_8013);
xor U10908 (N_10908,N_7742,N_9084);
and U10909 (N_10909,N_8634,N_6327);
or U10910 (N_10910,N_8312,N_6737);
and U10911 (N_10911,N_7253,N_6643);
or U10912 (N_10912,N_9340,N_9017);
xor U10913 (N_10913,N_6642,N_7318);
or U10914 (N_10914,N_6777,N_6439);
and U10915 (N_10915,N_7157,N_7400);
nand U10916 (N_10916,N_8965,N_6349);
nand U10917 (N_10917,N_8978,N_6565);
xor U10918 (N_10918,N_6700,N_8907);
and U10919 (N_10919,N_7559,N_6531);
and U10920 (N_10920,N_7751,N_7863);
nand U10921 (N_10921,N_6988,N_6740);
and U10922 (N_10922,N_7145,N_7289);
or U10923 (N_10923,N_7963,N_6770);
nor U10924 (N_10924,N_6404,N_6987);
and U10925 (N_10925,N_6315,N_6695);
nand U10926 (N_10926,N_8523,N_9277);
or U10927 (N_10927,N_7954,N_7565);
nor U10928 (N_10928,N_7808,N_8087);
and U10929 (N_10929,N_6459,N_9311);
and U10930 (N_10930,N_6639,N_9088);
and U10931 (N_10931,N_7436,N_7795);
and U10932 (N_10932,N_8426,N_7390);
nor U10933 (N_10933,N_9189,N_8459);
and U10934 (N_10934,N_7906,N_6273);
or U10935 (N_10935,N_6331,N_7743);
xor U10936 (N_10936,N_9350,N_7851);
nand U10937 (N_10937,N_8877,N_9195);
nand U10938 (N_10938,N_7009,N_7445);
xnor U10939 (N_10939,N_8101,N_8344);
xor U10940 (N_10940,N_7783,N_8475);
nor U10941 (N_10941,N_6929,N_8634);
and U10942 (N_10942,N_6922,N_7011);
and U10943 (N_10943,N_8051,N_7382);
or U10944 (N_10944,N_9061,N_9318);
nand U10945 (N_10945,N_7863,N_6592);
nor U10946 (N_10946,N_7136,N_9200);
and U10947 (N_10947,N_8857,N_7548);
or U10948 (N_10948,N_7592,N_6604);
or U10949 (N_10949,N_8107,N_6722);
and U10950 (N_10950,N_8090,N_8710);
nand U10951 (N_10951,N_7879,N_8339);
and U10952 (N_10952,N_6317,N_8019);
nor U10953 (N_10953,N_6670,N_7910);
nand U10954 (N_10954,N_7056,N_7500);
or U10955 (N_10955,N_7506,N_6828);
or U10956 (N_10956,N_8826,N_6585);
nand U10957 (N_10957,N_9083,N_8767);
nand U10958 (N_10958,N_7928,N_6546);
nor U10959 (N_10959,N_7563,N_6762);
or U10960 (N_10960,N_6454,N_7752);
nand U10961 (N_10961,N_9142,N_7759);
and U10962 (N_10962,N_7541,N_6307);
or U10963 (N_10963,N_7162,N_8508);
and U10964 (N_10964,N_7697,N_7317);
nand U10965 (N_10965,N_6923,N_6728);
nand U10966 (N_10966,N_6818,N_6930);
and U10967 (N_10967,N_7053,N_6560);
nor U10968 (N_10968,N_6279,N_7661);
or U10969 (N_10969,N_6992,N_6978);
and U10970 (N_10970,N_8096,N_6353);
nor U10971 (N_10971,N_8301,N_9078);
and U10972 (N_10972,N_6523,N_6560);
nor U10973 (N_10973,N_8398,N_8766);
or U10974 (N_10974,N_8740,N_8031);
nor U10975 (N_10975,N_6843,N_7453);
or U10976 (N_10976,N_8956,N_7739);
nand U10977 (N_10977,N_6626,N_8949);
or U10978 (N_10978,N_8825,N_7189);
or U10979 (N_10979,N_7800,N_7775);
and U10980 (N_10980,N_8981,N_7194);
xnor U10981 (N_10981,N_7268,N_7367);
nor U10982 (N_10982,N_8604,N_8700);
or U10983 (N_10983,N_9230,N_9157);
xor U10984 (N_10984,N_9343,N_8130);
nand U10985 (N_10985,N_7116,N_6442);
and U10986 (N_10986,N_7055,N_9017);
xor U10987 (N_10987,N_7451,N_6904);
and U10988 (N_10988,N_6902,N_9066);
nand U10989 (N_10989,N_6603,N_7142);
nor U10990 (N_10990,N_6431,N_9007);
nand U10991 (N_10991,N_7281,N_8210);
or U10992 (N_10992,N_6252,N_8063);
and U10993 (N_10993,N_7416,N_9085);
xor U10994 (N_10994,N_8149,N_7260);
nand U10995 (N_10995,N_7902,N_8497);
nand U10996 (N_10996,N_8469,N_7545);
nor U10997 (N_10997,N_6522,N_8904);
nor U10998 (N_10998,N_9272,N_8517);
nor U10999 (N_10999,N_9110,N_7731);
or U11000 (N_11000,N_8102,N_7343);
xnor U11001 (N_11001,N_6282,N_9012);
and U11002 (N_11002,N_9339,N_9071);
nand U11003 (N_11003,N_8040,N_8957);
nor U11004 (N_11004,N_7472,N_6981);
nor U11005 (N_11005,N_9035,N_6257);
nand U11006 (N_11006,N_8640,N_7104);
and U11007 (N_11007,N_8428,N_8183);
nor U11008 (N_11008,N_9281,N_8512);
or U11009 (N_11009,N_7604,N_7181);
and U11010 (N_11010,N_8826,N_6638);
nor U11011 (N_11011,N_8261,N_6287);
xor U11012 (N_11012,N_7005,N_7321);
nor U11013 (N_11013,N_9307,N_6544);
xor U11014 (N_11014,N_6430,N_9237);
and U11015 (N_11015,N_8024,N_7298);
xnor U11016 (N_11016,N_7891,N_6255);
and U11017 (N_11017,N_7089,N_7422);
and U11018 (N_11018,N_7449,N_6422);
nand U11019 (N_11019,N_8846,N_7713);
and U11020 (N_11020,N_7213,N_8678);
or U11021 (N_11021,N_7983,N_9348);
nand U11022 (N_11022,N_8227,N_6922);
nor U11023 (N_11023,N_6411,N_8717);
or U11024 (N_11024,N_8488,N_6999);
nor U11025 (N_11025,N_9216,N_7195);
or U11026 (N_11026,N_7216,N_8969);
nand U11027 (N_11027,N_6691,N_7830);
xnor U11028 (N_11028,N_7655,N_7886);
nor U11029 (N_11029,N_6509,N_7831);
nor U11030 (N_11030,N_7234,N_8170);
nor U11031 (N_11031,N_9262,N_7883);
or U11032 (N_11032,N_8523,N_6383);
or U11033 (N_11033,N_6630,N_7728);
and U11034 (N_11034,N_8439,N_8977);
nand U11035 (N_11035,N_6995,N_9306);
nand U11036 (N_11036,N_8881,N_7620);
nor U11037 (N_11037,N_8102,N_7137);
or U11038 (N_11038,N_8121,N_6410);
nand U11039 (N_11039,N_8305,N_8004);
and U11040 (N_11040,N_8433,N_8089);
or U11041 (N_11041,N_6632,N_8162);
or U11042 (N_11042,N_9199,N_7387);
and U11043 (N_11043,N_7081,N_7741);
and U11044 (N_11044,N_7799,N_8361);
or U11045 (N_11045,N_8138,N_8974);
nand U11046 (N_11046,N_6595,N_6565);
or U11047 (N_11047,N_8610,N_8262);
or U11048 (N_11048,N_8073,N_6731);
nand U11049 (N_11049,N_8299,N_7618);
nor U11050 (N_11050,N_8541,N_9215);
nor U11051 (N_11051,N_8180,N_8755);
nor U11052 (N_11052,N_9234,N_8272);
and U11053 (N_11053,N_9147,N_8858);
and U11054 (N_11054,N_8586,N_8198);
and U11055 (N_11055,N_9232,N_6994);
xnor U11056 (N_11056,N_6780,N_8720);
xnor U11057 (N_11057,N_7503,N_8831);
nor U11058 (N_11058,N_7893,N_8749);
and U11059 (N_11059,N_6463,N_7553);
xnor U11060 (N_11060,N_7847,N_8472);
nor U11061 (N_11061,N_6568,N_6749);
nor U11062 (N_11062,N_8416,N_8822);
xnor U11063 (N_11063,N_8118,N_7775);
and U11064 (N_11064,N_8218,N_9021);
and U11065 (N_11065,N_7176,N_7503);
or U11066 (N_11066,N_6554,N_8650);
or U11067 (N_11067,N_9330,N_7301);
nor U11068 (N_11068,N_7823,N_6612);
nor U11069 (N_11069,N_6762,N_6333);
nor U11070 (N_11070,N_6692,N_7941);
nor U11071 (N_11071,N_7580,N_7463);
nor U11072 (N_11072,N_6980,N_6366);
and U11073 (N_11073,N_6471,N_6704);
xor U11074 (N_11074,N_9247,N_8401);
nand U11075 (N_11075,N_8620,N_7499);
and U11076 (N_11076,N_7987,N_8344);
and U11077 (N_11077,N_7645,N_7526);
nor U11078 (N_11078,N_7713,N_6511);
nand U11079 (N_11079,N_7549,N_6441);
and U11080 (N_11080,N_8134,N_7273);
nand U11081 (N_11081,N_8396,N_8141);
and U11082 (N_11082,N_6337,N_6597);
nand U11083 (N_11083,N_7436,N_6764);
nor U11084 (N_11084,N_8517,N_9151);
and U11085 (N_11085,N_8513,N_8993);
nand U11086 (N_11086,N_6653,N_7369);
and U11087 (N_11087,N_8155,N_9174);
nand U11088 (N_11088,N_6425,N_8854);
and U11089 (N_11089,N_8473,N_7955);
and U11090 (N_11090,N_7509,N_9367);
and U11091 (N_11091,N_7739,N_8411);
or U11092 (N_11092,N_8800,N_9227);
or U11093 (N_11093,N_6926,N_7037);
nand U11094 (N_11094,N_8604,N_7837);
or U11095 (N_11095,N_8315,N_6777);
or U11096 (N_11096,N_6372,N_7463);
or U11097 (N_11097,N_7561,N_7322);
or U11098 (N_11098,N_6970,N_6563);
or U11099 (N_11099,N_8871,N_7284);
nor U11100 (N_11100,N_8729,N_7814);
nor U11101 (N_11101,N_9077,N_6450);
and U11102 (N_11102,N_7148,N_6355);
or U11103 (N_11103,N_9297,N_8405);
and U11104 (N_11104,N_6832,N_8104);
nor U11105 (N_11105,N_8435,N_8795);
nand U11106 (N_11106,N_7696,N_8983);
or U11107 (N_11107,N_8382,N_7514);
or U11108 (N_11108,N_8402,N_7466);
and U11109 (N_11109,N_7763,N_6416);
nand U11110 (N_11110,N_7962,N_8385);
or U11111 (N_11111,N_9357,N_7789);
and U11112 (N_11112,N_8241,N_9127);
and U11113 (N_11113,N_6936,N_7528);
and U11114 (N_11114,N_8503,N_7592);
nand U11115 (N_11115,N_8442,N_7210);
nor U11116 (N_11116,N_8778,N_9207);
nand U11117 (N_11117,N_8741,N_7858);
nor U11118 (N_11118,N_6300,N_7275);
or U11119 (N_11119,N_7748,N_9164);
or U11120 (N_11120,N_9021,N_6613);
or U11121 (N_11121,N_8390,N_9160);
nand U11122 (N_11122,N_7099,N_9221);
and U11123 (N_11123,N_9091,N_7646);
or U11124 (N_11124,N_8977,N_8635);
and U11125 (N_11125,N_6690,N_8020);
nor U11126 (N_11126,N_6832,N_7599);
and U11127 (N_11127,N_7696,N_6775);
nand U11128 (N_11128,N_8612,N_9211);
or U11129 (N_11129,N_8932,N_8346);
and U11130 (N_11130,N_8381,N_8156);
and U11131 (N_11131,N_8611,N_7080);
nor U11132 (N_11132,N_8483,N_6402);
or U11133 (N_11133,N_8028,N_6543);
nand U11134 (N_11134,N_7987,N_7674);
or U11135 (N_11135,N_8825,N_7700);
nand U11136 (N_11136,N_7910,N_7545);
nor U11137 (N_11137,N_8253,N_8509);
nor U11138 (N_11138,N_8339,N_6755);
nand U11139 (N_11139,N_6773,N_7696);
xnor U11140 (N_11140,N_7442,N_7125);
and U11141 (N_11141,N_7512,N_7373);
xnor U11142 (N_11142,N_9341,N_7615);
nand U11143 (N_11143,N_7246,N_7480);
nor U11144 (N_11144,N_8409,N_7347);
nor U11145 (N_11145,N_8726,N_7084);
nand U11146 (N_11146,N_8486,N_9335);
nor U11147 (N_11147,N_7853,N_8380);
or U11148 (N_11148,N_7903,N_7898);
nand U11149 (N_11149,N_8269,N_8389);
nor U11150 (N_11150,N_6427,N_6885);
nand U11151 (N_11151,N_8544,N_6705);
xor U11152 (N_11152,N_7143,N_9174);
or U11153 (N_11153,N_7254,N_7963);
nor U11154 (N_11154,N_9260,N_7077);
nand U11155 (N_11155,N_7397,N_9233);
or U11156 (N_11156,N_8470,N_9116);
or U11157 (N_11157,N_6531,N_6408);
or U11158 (N_11158,N_8870,N_8903);
nor U11159 (N_11159,N_8708,N_6530);
xnor U11160 (N_11160,N_7265,N_8165);
nor U11161 (N_11161,N_6498,N_7137);
nand U11162 (N_11162,N_9165,N_7283);
or U11163 (N_11163,N_6338,N_6414);
or U11164 (N_11164,N_7616,N_8238);
nor U11165 (N_11165,N_7173,N_7197);
or U11166 (N_11166,N_9221,N_8184);
nand U11167 (N_11167,N_9323,N_8958);
nand U11168 (N_11168,N_8517,N_9087);
nor U11169 (N_11169,N_8883,N_6853);
nand U11170 (N_11170,N_8796,N_7685);
or U11171 (N_11171,N_6906,N_8902);
xor U11172 (N_11172,N_9183,N_7717);
nor U11173 (N_11173,N_7009,N_6394);
nor U11174 (N_11174,N_6888,N_7966);
and U11175 (N_11175,N_9095,N_7291);
nand U11176 (N_11176,N_7263,N_6959);
nand U11177 (N_11177,N_6537,N_9305);
nor U11178 (N_11178,N_8091,N_8071);
nand U11179 (N_11179,N_6412,N_6373);
nand U11180 (N_11180,N_8268,N_6335);
or U11181 (N_11181,N_8470,N_9110);
and U11182 (N_11182,N_8014,N_7684);
xor U11183 (N_11183,N_7333,N_7289);
or U11184 (N_11184,N_6938,N_7400);
and U11185 (N_11185,N_8855,N_6553);
or U11186 (N_11186,N_7187,N_6825);
nand U11187 (N_11187,N_6780,N_7726);
nand U11188 (N_11188,N_8833,N_8578);
and U11189 (N_11189,N_6581,N_8364);
nor U11190 (N_11190,N_7094,N_8131);
and U11191 (N_11191,N_7110,N_8949);
and U11192 (N_11192,N_8916,N_7397);
nor U11193 (N_11193,N_7475,N_8904);
nand U11194 (N_11194,N_8751,N_8582);
and U11195 (N_11195,N_8127,N_7587);
or U11196 (N_11196,N_7587,N_6824);
nor U11197 (N_11197,N_6335,N_7593);
nor U11198 (N_11198,N_6979,N_7380);
or U11199 (N_11199,N_8265,N_7712);
xor U11200 (N_11200,N_8508,N_8772);
nand U11201 (N_11201,N_7346,N_7750);
or U11202 (N_11202,N_8313,N_6297);
nor U11203 (N_11203,N_6609,N_6666);
and U11204 (N_11204,N_8123,N_7052);
and U11205 (N_11205,N_7191,N_8146);
nand U11206 (N_11206,N_6291,N_6804);
xor U11207 (N_11207,N_7188,N_6447);
and U11208 (N_11208,N_7563,N_8784);
and U11209 (N_11209,N_7024,N_7978);
and U11210 (N_11210,N_7390,N_9114);
xnor U11211 (N_11211,N_8738,N_7355);
nor U11212 (N_11212,N_7212,N_7730);
nor U11213 (N_11213,N_6678,N_8447);
or U11214 (N_11214,N_9199,N_6969);
and U11215 (N_11215,N_8251,N_7325);
nor U11216 (N_11216,N_8232,N_9015);
nand U11217 (N_11217,N_6402,N_8142);
nor U11218 (N_11218,N_8034,N_7438);
nand U11219 (N_11219,N_7081,N_7699);
and U11220 (N_11220,N_8295,N_8088);
and U11221 (N_11221,N_6829,N_6390);
nor U11222 (N_11222,N_6707,N_8199);
and U11223 (N_11223,N_7859,N_8040);
nand U11224 (N_11224,N_8895,N_8649);
or U11225 (N_11225,N_7723,N_7847);
and U11226 (N_11226,N_8340,N_6426);
or U11227 (N_11227,N_6681,N_7791);
nor U11228 (N_11228,N_9122,N_7973);
or U11229 (N_11229,N_8899,N_9237);
nor U11230 (N_11230,N_7928,N_7393);
and U11231 (N_11231,N_9344,N_7254);
nand U11232 (N_11232,N_8282,N_8858);
and U11233 (N_11233,N_8338,N_7680);
nand U11234 (N_11234,N_9266,N_8117);
nand U11235 (N_11235,N_8469,N_7104);
nor U11236 (N_11236,N_6834,N_6829);
and U11237 (N_11237,N_7376,N_9043);
nand U11238 (N_11238,N_8812,N_8776);
nand U11239 (N_11239,N_8897,N_7534);
nor U11240 (N_11240,N_7913,N_8510);
and U11241 (N_11241,N_8605,N_6500);
and U11242 (N_11242,N_7199,N_7465);
xor U11243 (N_11243,N_8400,N_8548);
and U11244 (N_11244,N_9350,N_6833);
and U11245 (N_11245,N_8621,N_7481);
nor U11246 (N_11246,N_7064,N_8838);
nand U11247 (N_11247,N_8385,N_8052);
nand U11248 (N_11248,N_7267,N_8399);
or U11249 (N_11249,N_8281,N_7950);
nand U11250 (N_11250,N_9084,N_8523);
or U11251 (N_11251,N_8495,N_7553);
nand U11252 (N_11252,N_6892,N_6326);
and U11253 (N_11253,N_8374,N_7641);
and U11254 (N_11254,N_6697,N_6296);
nor U11255 (N_11255,N_7371,N_8403);
and U11256 (N_11256,N_8301,N_8871);
xor U11257 (N_11257,N_6740,N_8376);
or U11258 (N_11258,N_8713,N_7936);
xor U11259 (N_11259,N_7895,N_6742);
xor U11260 (N_11260,N_9254,N_8598);
nand U11261 (N_11261,N_7024,N_6378);
and U11262 (N_11262,N_7333,N_6264);
nand U11263 (N_11263,N_6261,N_8103);
nand U11264 (N_11264,N_7418,N_8196);
nand U11265 (N_11265,N_7846,N_7400);
and U11266 (N_11266,N_8713,N_8650);
or U11267 (N_11267,N_7574,N_8538);
xnor U11268 (N_11268,N_7098,N_8566);
nor U11269 (N_11269,N_6937,N_7904);
or U11270 (N_11270,N_8637,N_8244);
nand U11271 (N_11271,N_8688,N_8234);
nor U11272 (N_11272,N_6626,N_6965);
nand U11273 (N_11273,N_8063,N_7363);
nor U11274 (N_11274,N_9028,N_7544);
and U11275 (N_11275,N_7559,N_7616);
and U11276 (N_11276,N_6421,N_7784);
nor U11277 (N_11277,N_8955,N_7295);
nand U11278 (N_11278,N_8473,N_8387);
nor U11279 (N_11279,N_7101,N_8202);
nor U11280 (N_11280,N_9244,N_9196);
nor U11281 (N_11281,N_9334,N_9188);
nor U11282 (N_11282,N_8746,N_8219);
and U11283 (N_11283,N_9072,N_8820);
and U11284 (N_11284,N_7009,N_8291);
and U11285 (N_11285,N_7504,N_7725);
and U11286 (N_11286,N_8438,N_7259);
or U11287 (N_11287,N_8222,N_8118);
nand U11288 (N_11288,N_7587,N_7454);
xor U11289 (N_11289,N_6730,N_9050);
nor U11290 (N_11290,N_9030,N_9312);
or U11291 (N_11291,N_9139,N_8475);
nor U11292 (N_11292,N_7147,N_6818);
and U11293 (N_11293,N_7235,N_6435);
or U11294 (N_11294,N_8989,N_6553);
and U11295 (N_11295,N_9169,N_9285);
xnor U11296 (N_11296,N_9199,N_7455);
and U11297 (N_11297,N_7926,N_7747);
and U11298 (N_11298,N_7109,N_7099);
nand U11299 (N_11299,N_7482,N_9046);
nand U11300 (N_11300,N_8455,N_8060);
or U11301 (N_11301,N_8838,N_7765);
nor U11302 (N_11302,N_8880,N_9288);
nand U11303 (N_11303,N_7682,N_9272);
nor U11304 (N_11304,N_6849,N_7111);
nor U11305 (N_11305,N_6370,N_7354);
and U11306 (N_11306,N_7054,N_7110);
nor U11307 (N_11307,N_8980,N_8982);
or U11308 (N_11308,N_9148,N_7032);
nand U11309 (N_11309,N_8638,N_9260);
and U11310 (N_11310,N_7008,N_8780);
xnor U11311 (N_11311,N_6449,N_8104);
nor U11312 (N_11312,N_7719,N_7107);
or U11313 (N_11313,N_6835,N_7288);
xnor U11314 (N_11314,N_7377,N_6290);
nor U11315 (N_11315,N_8119,N_9202);
nand U11316 (N_11316,N_8054,N_7372);
nor U11317 (N_11317,N_8013,N_8283);
nor U11318 (N_11318,N_6349,N_7024);
nor U11319 (N_11319,N_8284,N_6287);
nor U11320 (N_11320,N_7929,N_7147);
or U11321 (N_11321,N_7545,N_8064);
nand U11322 (N_11322,N_6973,N_9300);
and U11323 (N_11323,N_8331,N_8563);
and U11324 (N_11324,N_8222,N_6673);
and U11325 (N_11325,N_7723,N_8963);
nor U11326 (N_11326,N_8353,N_8719);
nand U11327 (N_11327,N_7081,N_8635);
nor U11328 (N_11328,N_9353,N_8481);
and U11329 (N_11329,N_8357,N_8696);
nor U11330 (N_11330,N_8640,N_7722);
nand U11331 (N_11331,N_7476,N_8411);
and U11332 (N_11332,N_8590,N_8093);
xor U11333 (N_11333,N_9004,N_6429);
nor U11334 (N_11334,N_7297,N_6915);
and U11335 (N_11335,N_6448,N_9293);
and U11336 (N_11336,N_6279,N_7023);
or U11337 (N_11337,N_7366,N_7415);
nor U11338 (N_11338,N_6314,N_7017);
nand U11339 (N_11339,N_8451,N_6365);
nand U11340 (N_11340,N_9023,N_9308);
and U11341 (N_11341,N_8310,N_6668);
xnor U11342 (N_11342,N_6759,N_8795);
or U11343 (N_11343,N_6509,N_8728);
nand U11344 (N_11344,N_8261,N_8559);
or U11345 (N_11345,N_9161,N_8758);
nor U11346 (N_11346,N_8326,N_6587);
nor U11347 (N_11347,N_7849,N_6518);
nor U11348 (N_11348,N_7725,N_8107);
and U11349 (N_11349,N_6646,N_7126);
nor U11350 (N_11350,N_7464,N_8953);
nor U11351 (N_11351,N_7746,N_8881);
nand U11352 (N_11352,N_7271,N_6841);
or U11353 (N_11353,N_9091,N_9316);
or U11354 (N_11354,N_7344,N_8930);
and U11355 (N_11355,N_6857,N_6897);
or U11356 (N_11356,N_8378,N_8081);
and U11357 (N_11357,N_7739,N_6609);
or U11358 (N_11358,N_8336,N_8717);
and U11359 (N_11359,N_9237,N_7909);
and U11360 (N_11360,N_9343,N_7793);
and U11361 (N_11361,N_8991,N_6898);
nor U11362 (N_11362,N_7945,N_6332);
and U11363 (N_11363,N_8913,N_7048);
nand U11364 (N_11364,N_7970,N_7384);
nand U11365 (N_11365,N_8185,N_9367);
xor U11366 (N_11366,N_6485,N_8347);
nor U11367 (N_11367,N_7718,N_6309);
xor U11368 (N_11368,N_6959,N_8941);
or U11369 (N_11369,N_9112,N_9273);
nand U11370 (N_11370,N_8203,N_6657);
nor U11371 (N_11371,N_8211,N_7342);
or U11372 (N_11372,N_6699,N_8756);
and U11373 (N_11373,N_9352,N_7439);
nand U11374 (N_11374,N_6790,N_8897);
or U11375 (N_11375,N_7313,N_6494);
nand U11376 (N_11376,N_8650,N_8440);
nor U11377 (N_11377,N_7135,N_8506);
nand U11378 (N_11378,N_9364,N_7405);
nor U11379 (N_11379,N_7072,N_9009);
xnor U11380 (N_11380,N_7787,N_8915);
and U11381 (N_11381,N_9336,N_8144);
nand U11382 (N_11382,N_9350,N_7197);
and U11383 (N_11383,N_8523,N_8662);
nand U11384 (N_11384,N_7734,N_6663);
and U11385 (N_11385,N_8741,N_8658);
nand U11386 (N_11386,N_9304,N_8252);
nand U11387 (N_11387,N_6873,N_9028);
xor U11388 (N_11388,N_9213,N_8432);
or U11389 (N_11389,N_8222,N_9123);
xnor U11390 (N_11390,N_6251,N_9180);
and U11391 (N_11391,N_6514,N_6638);
and U11392 (N_11392,N_7613,N_7901);
or U11393 (N_11393,N_7837,N_6285);
or U11394 (N_11394,N_8310,N_8928);
nor U11395 (N_11395,N_7384,N_6262);
nor U11396 (N_11396,N_6980,N_7313);
nand U11397 (N_11397,N_7547,N_9150);
nand U11398 (N_11398,N_7910,N_8581);
nand U11399 (N_11399,N_9307,N_9221);
nor U11400 (N_11400,N_7473,N_6706);
nand U11401 (N_11401,N_7478,N_6655);
nor U11402 (N_11402,N_7636,N_8138);
nand U11403 (N_11403,N_7269,N_7132);
and U11404 (N_11404,N_6522,N_6351);
xor U11405 (N_11405,N_9325,N_8211);
and U11406 (N_11406,N_9271,N_7018);
nand U11407 (N_11407,N_6612,N_6929);
and U11408 (N_11408,N_8572,N_8796);
xor U11409 (N_11409,N_6873,N_7946);
and U11410 (N_11410,N_8882,N_8439);
nor U11411 (N_11411,N_6952,N_7662);
nand U11412 (N_11412,N_6614,N_9292);
nand U11413 (N_11413,N_8708,N_6569);
nand U11414 (N_11414,N_6817,N_7716);
nor U11415 (N_11415,N_6268,N_6526);
nand U11416 (N_11416,N_7032,N_7273);
xnor U11417 (N_11417,N_6621,N_7254);
and U11418 (N_11418,N_9146,N_9218);
nand U11419 (N_11419,N_8427,N_7494);
xor U11420 (N_11420,N_7639,N_6585);
nor U11421 (N_11421,N_8073,N_6751);
nand U11422 (N_11422,N_8220,N_8448);
or U11423 (N_11423,N_8264,N_6642);
nand U11424 (N_11424,N_8875,N_9032);
and U11425 (N_11425,N_6595,N_8883);
xnor U11426 (N_11426,N_7588,N_8257);
nand U11427 (N_11427,N_8818,N_6552);
and U11428 (N_11428,N_8063,N_7861);
or U11429 (N_11429,N_8172,N_7900);
nand U11430 (N_11430,N_6725,N_6908);
or U11431 (N_11431,N_9085,N_6766);
or U11432 (N_11432,N_6722,N_7652);
and U11433 (N_11433,N_7914,N_7828);
and U11434 (N_11434,N_6548,N_8665);
nor U11435 (N_11435,N_7508,N_9184);
or U11436 (N_11436,N_8014,N_8011);
nor U11437 (N_11437,N_9075,N_6597);
nor U11438 (N_11438,N_8444,N_6549);
or U11439 (N_11439,N_9179,N_8151);
or U11440 (N_11440,N_6385,N_7334);
nand U11441 (N_11441,N_7439,N_7601);
nor U11442 (N_11442,N_6468,N_8010);
and U11443 (N_11443,N_6837,N_6818);
nand U11444 (N_11444,N_8748,N_9347);
and U11445 (N_11445,N_8991,N_6771);
nor U11446 (N_11446,N_7330,N_7406);
nor U11447 (N_11447,N_9330,N_8622);
and U11448 (N_11448,N_7320,N_7483);
xor U11449 (N_11449,N_8777,N_8477);
or U11450 (N_11450,N_6998,N_8271);
nand U11451 (N_11451,N_8923,N_7399);
and U11452 (N_11452,N_9111,N_7555);
nor U11453 (N_11453,N_6250,N_8756);
and U11454 (N_11454,N_8355,N_6295);
and U11455 (N_11455,N_6426,N_7074);
nand U11456 (N_11456,N_7196,N_8847);
nor U11457 (N_11457,N_7957,N_8310);
nor U11458 (N_11458,N_7458,N_8540);
nand U11459 (N_11459,N_9040,N_6684);
and U11460 (N_11460,N_9163,N_6864);
nand U11461 (N_11461,N_6944,N_8112);
or U11462 (N_11462,N_6623,N_6465);
or U11463 (N_11463,N_6962,N_7587);
xor U11464 (N_11464,N_6653,N_7302);
or U11465 (N_11465,N_7972,N_6827);
or U11466 (N_11466,N_7589,N_7964);
and U11467 (N_11467,N_7549,N_7552);
and U11468 (N_11468,N_8390,N_7187);
or U11469 (N_11469,N_8064,N_8352);
nor U11470 (N_11470,N_7870,N_8087);
or U11471 (N_11471,N_7455,N_6254);
or U11472 (N_11472,N_8341,N_7296);
nor U11473 (N_11473,N_7331,N_7528);
or U11474 (N_11474,N_7919,N_7236);
and U11475 (N_11475,N_6347,N_8463);
and U11476 (N_11476,N_7132,N_7172);
nand U11477 (N_11477,N_6601,N_6728);
nand U11478 (N_11478,N_6563,N_7150);
xor U11479 (N_11479,N_6510,N_7717);
nor U11480 (N_11480,N_8075,N_8387);
or U11481 (N_11481,N_9218,N_8300);
nand U11482 (N_11482,N_8854,N_7720);
and U11483 (N_11483,N_8017,N_7607);
xnor U11484 (N_11484,N_9240,N_6736);
and U11485 (N_11485,N_7469,N_8318);
nand U11486 (N_11486,N_7331,N_7894);
nor U11487 (N_11487,N_6292,N_6940);
or U11488 (N_11488,N_9012,N_7852);
nand U11489 (N_11489,N_6922,N_7779);
xor U11490 (N_11490,N_6360,N_8869);
nor U11491 (N_11491,N_8669,N_7409);
nand U11492 (N_11492,N_8906,N_8080);
or U11493 (N_11493,N_6250,N_7151);
or U11494 (N_11494,N_7365,N_7183);
and U11495 (N_11495,N_7815,N_6819);
xnor U11496 (N_11496,N_8523,N_8200);
and U11497 (N_11497,N_9076,N_8615);
nor U11498 (N_11498,N_8981,N_6907);
xnor U11499 (N_11499,N_9119,N_6901);
and U11500 (N_11500,N_8808,N_7516);
and U11501 (N_11501,N_6385,N_8310);
nor U11502 (N_11502,N_7435,N_8340);
nand U11503 (N_11503,N_7098,N_6731);
nand U11504 (N_11504,N_7169,N_8947);
or U11505 (N_11505,N_8355,N_7137);
xnor U11506 (N_11506,N_7406,N_6876);
nand U11507 (N_11507,N_6941,N_9025);
or U11508 (N_11508,N_8944,N_7317);
and U11509 (N_11509,N_9349,N_7794);
nor U11510 (N_11510,N_6794,N_6850);
nor U11511 (N_11511,N_6834,N_9238);
nand U11512 (N_11512,N_8210,N_8031);
and U11513 (N_11513,N_6789,N_7110);
and U11514 (N_11514,N_7134,N_8143);
and U11515 (N_11515,N_6579,N_6332);
and U11516 (N_11516,N_8906,N_6363);
nand U11517 (N_11517,N_9355,N_8337);
nor U11518 (N_11518,N_8851,N_8088);
or U11519 (N_11519,N_6719,N_9065);
and U11520 (N_11520,N_7857,N_8803);
nand U11521 (N_11521,N_8339,N_8846);
nor U11522 (N_11522,N_8847,N_6255);
nand U11523 (N_11523,N_8970,N_7058);
nor U11524 (N_11524,N_6955,N_6344);
or U11525 (N_11525,N_9163,N_9068);
nand U11526 (N_11526,N_6651,N_7861);
nand U11527 (N_11527,N_8255,N_9329);
and U11528 (N_11528,N_6918,N_7542);
and U11529 (N_11529,N_7890,N_7181);
and U11530 (N_11530,N_6921,N_8916);
nand U11531 (N_11531,N_8439,N_6517);
nor U11532 (N_11532,N_9284,N_8944);
and U11533 (N_11533,N_7567,N_7100);
xor U11534 (N_11534,N_8641,N_9299);
nand U11535 (N_11535,N_8792,N_7192);
or U11536 (N_11536,N_8961,N_9127);
xnor U11537 (N_11537,N_7564,N_6385);
nor U11538 (N_11538,N_9127,N_9337);
xnor U11539 (N_11539,N_6463,N_8318);
xor U11540 (N_11540,N_7238,N_6585);
nor U11541 (N_11541,N_8188,N_7461);
nor U11542 (N_11542,N_9088,N_6747);
and U11543 (N_11543,N_8879,N_6994);
or U11544 (N_11544,N_7338,N_7193);
nand U11545 (N_11545,N_7364,N_6256);
nor U11546 (N_11546,N_8142,N_7886);
and U11547 (N_11547,N_8423,N_8756);
nor U11548 (N_11548,N_7330,N_7771);
or U11549 (N_11549,N_8978,N_8040);
and U11550 (N_11550,N_6774,N_7532);
xnor U11551 (N_11551,N_9008,N_6817);
or U11552 (N_11552,N_8001,N_8220);
nand U11553 (N_11553,N_8010,N_6798);
and U11554 (N_11554,N_7991,N_7286);
or U11555 (N_11555,N_9117,N_6813);
and U11556 (N_11556,N_7159,N_7590);
and U11557 (N_11557,N_9316,N_6714);
and U11558 (N_11558,N_7383,N_6805);
nand U11559 (N_11559,N_8259,N_8219);
nand U11560 (N_11560,N_8727,N_6893);
nor U11561 (N_11561,N_7466,N_7418);
or U11562 (N_11562,N_8334,N_6360);
and U11563 (N_11563,N_8695,N_9227);
nand U11564 (N_11564,N_9303,N_7889);
or U11565 (N_11565,N_7034,N_7621);
nor U11566 (N_11566,N_7035,N_8766);
or U11567 (N_11567,N_7302,N_8016);
and U11568 (N_11568,N_6759,N_7428);
nor U11569 (N_11569,N_7577,N_8650);
nand U11570 (N_11570,N_8377,N_8778);
nand U11571 (N_11571,N_8957,N_9305);
or U11572 (N_11572,N_8483,N_6715);
and U11573 (N_11573,N_6704,N_8114);
xnor U11574 (N_11574,N_7020,N_7675);
nor U11575 (N_11575,N_7853,N_7489);
nor U11576 (N_11576,N_9174,N_7045);
xnor U11577 (N_11577,N_8423,N_7074);
xnor U11578 (N_11578,N_6533,N_6897);
and U11579 (N_11579,N_8329,N_7047);
or U11580 (N_11580,N_6487,N_7061);
nor U11581 (N_11581,N_8269,N_7075);
or U11582 (N_11582,N_8035,N_7474);
nand U11583 (N_11583,N_9249,N_6679);
or U11584 (N_11584,N_7629,N_7397);
and U11585 (N_11585,N_7684,N_6622);
and U11586 (N_11586,N_7884,N_7756);
xor U11587 (N_11587,N_9078,N_9076);
nor U11588 (N_11588,N_8608,N_7052);
or U11589 (N_11589,N_8879,N_6820);
and U11590 (N_11590,N_8654,N_8354);
nand U11591 (N_11591,N_7096,N_8655);
nor U11592 (N_11592,N_7470,N_7829);
and U11593 (N_11593,N_6318,N_9142);
nand U11594 (N_11594,N_9348,N_8969);
nand U11595 (N_11595,N_6997,N_9293);
nand U11596 (N_11596,N_8353,N_7169);
or U11597 (N_11597,N_8996,N_8818);
or U11598 (N_11598,N_8156,N_6270);
xnor U11599 (N_11599,N_7317,N_7834);
and U11600 (N_11600,N_8801,N_9110);
and U11601 (N_11601,N_9109,N_8750);
nand U11602 (N_11602,N_8869,N_8581);
nand U11603 (N_11603,N_8888,N_7018);
xnor U11604 (N_11604,N_8297,N_9102);
or U11605 (N_11605,N_8455,N_7987);
or U11606 (N_11606,N_7123,N_6559);
or U11607 (N_11607,N_7756,N_8116);
nor U11608 (N_11608,N_7988,N_8579);
and U11609 (N_11609,N_8896,N_7831);
nor U11610 (N_11610,N_8491,N_6402);
and U11611 (N_11611,N_7292,N_8171);
nand U11612 (N_11612,N_8297,N_6784);
or U11613 (N_11613,N_7482,N_9204);
nor U11614 (N_11614,N_8354,N_7824);
nand U11615 (N_11615,N_7327,N_7922);
or U11616 (N_11616,N_6336,N_9075);
or U11617 (N_11617,N_7089,N_6795);
or U11618 (N_11618,N_8311,N_6493);
and U11619 (N_11619,N_8402,N_6800);
and U11620 (N_11620,N_6992,N_7749);
nand U11621 (N_11621,N_8231,N_7956);
nor U11622 (N_11622,N_7431,N_7388);
xor U11623 (N_11623,N_7888,N_9015);
and U11624 (N_11624,N_8254,N_8980);
and U11625 (N_11625,N_7766,N_9337);
nand U11626 (N_11626,N_6582,N_6837);
nand U11627 (N_11627,N_7628,N_8167);
or U11628 (N_11628,N_8788,N_7564);
nand U11629 (N_11629,N_6364,N_7145);
and U11630 (N_11630,N_7508,N_7681);
nand U11631 (N_11631,N_6980,N_7019);
or U11632 (N_11632,N_6431,N_8134);
nor U11633 (N_11633,N_6517,N_9230);
nand U11634 (N_11634,N_6979,N_6803);
nand U11635 (N_11635,N_6373,N_8110);
nand U11636 (N_11636,N_7346,N_6372);
nor U11637 (N_11637,N_8128,N_9062);
nand U11638 (N_11638,N_7872,N_8190);
nand U11639 (N_11639,N_6659,N_7595);
nand U11640 (N_11640,N_7101,N_6374);
nand U11641 (N_11641,N_8166,N_9097);
nand U11642 (N_11642,N_6893,N_8028);
nand U11643 (N_11643,N_7571,N_6435);
or U11644 (N_11644,N_6745,N_8533);
or U11645 (N_11645,N_7012,N_7890);
or U11646 (N_11646,N_7587,N_8569);
nor U11647 (N_11647,N_9220,N_7186);
and U11648 (N_11648,N_9055,N_8761);
and U11649 (N_11649,N_8225,N_7705);
or U11650 (N_11650,N_7086,N_6567);
or U11651 (N_11651,N_6786,N_7718);
nor U11652 (N_11652,N_6913,N_9194);
or U11653 (N_11653,N_7658,N_7966);
nand U11654 (N_11654,N_8879,N_9061);
nor U11655 (N_11655,N_8552,N_7504);
and U11656 (N_11656,N_7462,N_8069);
xnor U11657 (N_11657,N_6395,N_6716);
nor U11658 (N_11658,N_8481,N_8103);
or U11659 (N_11659,N_6405,N_8104);
and U11660 (N_11660,N_6991,N_7344);
and U11661 (N_11661,N_7304,N_8158);
or U11662 (N_11662,N_7306,N_9070);
nand U11663 (N_11663,N_7860,N_8628);
xor U11664 (N_11664,N_9109,N_7012);
nand U11665 (N_11665,N_8119,N_8059);
and U11666 (N_11666,N_7487,N_7507);
nor U11667 (N_11667,N_7887,N_7664);
or U11668 (N_11668,N_9215,N_8788);
nor U11669 (N_11669,N_8957,N_6692);
nand U11670 (N_11670,N_8439,N_6624);
and U11671 (N_11671,N_7966,N_7768);
and U11672 (N_11672,N_9225,N_7017);
and U11673 (N_11673,N_9368,N_6339);
nor U11674 (N_11674,N_8609,N_7960);
and U11675 (N_11675,N_9179,N_9256);
or U11676 (N_11676,N_6515,N_6604);
nor U11677 (N_11677,N_9081,N_8945);
nand U11678 (N_11678,N_6643,N_8829);
nor U11679 (N_11679,N_7880,N_7808);
nand U11680 (N_11680,N_7890,N_6481);
and U11681 (N_11681,N_8307,N_8202);
xor U11682 (N_11682,N_7935,N_6802);
or U11683 (N_11683,N_6432,N_7408);
nor U11684 (N_11684,N_6664,N_9041);
and U11685 (N_11685,N_8546,N_7654);
xnor U11686 (N_11686,N_7821,N_6280);
nor U11687 (N_11687,N_8589,N_7056);
nor U11688 (N_11688,N_7691,N_9067);
xor U11689 (N_11689,N_6529,N_6658);
or U11690 (N_11690,N_6275,N_8422);
nor U11691 (N_11691,N_7672,N_8893);
nor U11692 (N_11692,N_6268,N_8239);
nand U11693 (N_11693,N_8593,N_8801);
nor U11694 (N_11694,N_8704,N_9370);
or U11695 (N_11695,N_6989,N_8991);
or U11696 (N_11696,N_6450,N_7751);
xor U11697 (N_11697,N_9373,N_9005);
or U11698 (N_11698,N_6635,N_7098);
nand U11699 (N_11699,N_8521,N_6833);
and U11700 (N_11700,N_6587,N_7264);
or U11701 (N_11701,N_9047,N_7735);
or U11702 (N_11702,N_7294,N_7242);
nand U11703 (N_11703,N_8335,N_8301);
nand U11704 (N_11704,N_6897,N_8267);
nor U11705 (N_11705,N_6798,N_6459);
nor U11706 (N_11706,N_8555,N_7626);
or U11707 (N_11707,N_6580,N_7401);
nor U11708 (N_11708,N_8146,N_8193);
nand U11709 (N_11709,N_6690,N_6503);
nor U11710 (N_11710,N_9153,N_8268);
or U11711 (N_11711,N_7441,N_9304);
nor U11712 (N_11712,N_8641,N_6929);
or U11713 (N_11713,N_6373,N_6333);
and U11714 (N_11714,N_7094,N_6509);
and U11715 (N_11715,N_7280,N_6676);
or U11716 (N_11716,N_7835,N_7555);
nand U11717 (N_11717,N_7388,N_7505);
or U11718 (N_11718,N_7325,N_9170);
xnor U11719 (N_11719,N_6460,N_9166);
nor U11720 (N_11720,N_8925,N_7189);
or U11721 (N_11721,N_9052,N_8887);
and U11722 (N_11722,N_7936,N_6369);
nor U11723 (N_11723,N_7423,N_7185);
nand U11724 (N_11724,N_6582,N_7037);
and U11725 (N_11725,N_6831,N_7003);
nor U11726 (N_11726,N_8828,N_7319);
nand U11727 (N_11727,N_8446,N_6792);
xor U11728 (N_11728,N_8880,N_6344);
xnor U11729 (N_11729,N_6308,N_8831);
nand U11730 (N_11730,N_8607,N_8205);
nor U11731 (N_11731,N_8963,N_6990);
or U11732 (N_11732,N_7710,N_8612);
nand U11733 (N_11733,N_8754,N_7002);
and U11734 (N_11734,N_7875,N_8155);
xor U11735 (N_11735,N_6405,N_6912);
nand U11736 (N_11736,N_7984,N_6676);
or U11737 (N_11737,N_8875,N_8434);
nand U11738 (N_11738,N_9151,N_8322);
and U11739 (N_11739,N_8100,N_7490);
xor U11740 (N_11740,N_6550,N_7863);
or U11741 (N_11741,N_7101,N_7358);
xnor U11742 (N_11742,N_7350,N_8655);
and U11743 (N_11743,N_6741,N_8852);
nand U11744 (N_11744,N_6436,N_9142);
and U11745 (N_11745,N_9294,N_6695);
and U11746 (N_11746,N_8353,N_8990);
or U11747 (N_11747,N_8205,N_6851);
nand U11748 (N_11748,N_6905,N_8062);
xnor U11749 (N_11749,N_8381,N_9225);
or U11750 (N_11750,N_7356,N_7445);
xnor U11751 (N_11751,N_6273,N_7818);
nand U11752 (N_11752,N_7807,N_8117);
nand U11753 (N_11753,N_8582,N_9356);
and U11754 (N_11754,N_7292,N_7109);
and U11755 (N_11755,N_7628,N_9275);
nor U11756 (N_11756,N_7866,N_7401);
nand U11757 (N_11757,N_8481,N_7835);
and U11758 (N_11758,N_6835,N_6276);
or U11759 (N_11759,N_7620,N_7233);
and U11760 (N_11760,N_8642,N_7333);
xor U11761 (N_11761,N_8935,N_8872);
or U11762 (N_11762,N_6441,N_8377);
or U11763 (N_11763,N_8222,N_9045);
or U11764 (N_11764,N_8318,N_8503);
nand U11765 (N_11765,N_7715,N_6959);
or U11766 (N_11766,N_7805,N_8658);
nand U11767 (N_11767,N_7403,N_9039);
nand U11768 (N_11768,N_6475,N_7629);
nand U11769 (N_11769,N_8709,N_6461);
nor U11770 (N_11770,N_9367,N_8131);
nor U11771 (N_11771,N_7495,N_8245);
nand U11772 (N_11772,N_8401,N_7899);
nor U11773 (N_11773,N_7723,N_6933);
and U11774 (N_11774,N_7951,N_7633);
nor U11775 (N_11775,N_7287,N_7224);
nor U11776 (N_11776,N_9065,N_8020);
and U11777 (N_11777,N_7151,N_8297);
and U11778 (N_11778,N_8569,N_7951);
or U11779 (N_11779,N_7429,N_9352);
and U11780 (N_11780,N_7246,N_6407);
or U11781 (N_11781,N_8091,N_8963);
nand U11782 (N_11782,N_7972,N_7720);
and U11783 (N_11783,N_8616,N_8832);
nand U11784 (N_11784,N_8409,N_8270);
nor U11785 (N_11785,N_8325,N_8829);
nand U11786 (N_11786,N_6287,N_7312);
nand U11787 (N_11787,N_8293,N_6965);
xor U11788 (N_11788,N_7520,N_8140);
nor U11789 (N_11789,N_7774,N_6821);
nand U11790 (N_11790,N_9313,N_6493);
and U11791 (N_11791,N_9077,N_7897);
and U11792 (N_11792,N_8183,N_7599);
and U11793 (N_11793,N_6535,N_8290);
or U11794 (N_11794,N_8931,N_8945);
or U11795 (N_11795,N_7067,N_7607);
xor U11796 (N_11796,N_6354,N_8812);
nand U11797 (N_11797,N_6888,N_8187);
nand U11798 (N_11798,N_6329,N_7326);
nor U11799 (N_11799,N_6422,N_7959);
and U11800 (N_11800,N_7577,N_8384);
or U11801 (N_11801,N_7422,N_9081);
nor U11802 (N_11802,N_8310,N_8707);
nor U11803 (N_11803,N_8662,N_6361);
and U11804 (N_11804,N_8966,N_8436);
and U11805 (N_11805,N_6862,N_7676);
nand U11806 (N_11806,N_7754,N_7042);
and U11807 (N_11807,N_7347,N_8788);
and U11808 (N_11808,N_8394,N_8305);
nor U11809 (N_11809,N_7488,N_7384);
xor U11810 (N_11810,N_7766,N_8304);
nor U11811 (N_11811,N_7837,N_8929);
and U11812 (N_11812,N_6903,N_7765);
xor U11813 (N_11813,N_6426,N_6943);
or U11814 (N_11814,N_7973,N_9296);
and U11815 (N_11815,N_7767,N_8332);
nor U11816 (N_11816,N_7062,N_6729);
nor U11817 (N_11817,N_7375,N_8402);
or U11818 (N_11818,N_8605,N_8721);
nor U11819 (N_11819,N_7198,N_6462);
nor U11820 (N_11820,N_9316,N_7313);
xnor U11821 (N_11821,N_7175,N_8713);
or U11822 (N_11822,N_8601,N_9273);
or U11823 (N_11823,N_7074,N_7287);
nand U11824 (N_11824,N_6347,N_7013);
and U11825 (N_11825,N_8169,N_8249);
and U11826 (N_11826,N_8618,N_8893);
and U11827 (N_11827,N_7049,N_6721);
nand U11828 (N_11828,N_7845,N_8358);
nand U11829 (N_11829,N_7409,N_8364);
or U11830 (N_11830,N_6703,N_8585);
and U11831 (N_11831,N_6420,N_6324);
nand U11832 (N_11832,N_8147,N_8703);
nor U11833 (N_11833,N_6812,N_7111);
nand U11834 (N_11834,N_7522,N_7039);
nand U11835 (N_11835,N_7147,N_8749);
nand U11836 (N_11836,N_9082,N_6602);
or U11837 (N_11837,N_8897,N_7413);
or U11838 (N_11838,N_6275,N_7917);
nor U11839 (N_11839,N_6839,N_6470);
nand U11840 (N_11840,N_6791,N_7089);
nor U11841 (N_11841,N_7855,N_8832);
nor U11842 (N_11842,N_7346,N_9128);
nand U11843 (N_11843,N_7834,N_8015);
nor U11844 (N_11844,N_6401,N_7001);
or U11845 (N_11845,N_7505,N_8733);
nor U11846 (N_11846,N_7938,N_8024);
xor U11847 (N_11847,N_9257,N_6560);
xor U11848 (N_11848,N_7035,N_8778);
nand U11849 (N_11849,N_8930,N_9082);
and U11850 (N_11850,N_7115,N_8557);
or U11851 (N_11851,N_6284,N_6731);
nor U11852 (N_11852,N_7217,N_6503);
nand U11853 (N_11853,N_7991,N_8554);
or U11854 (N_11854,N_7848,N_7472);
nand U11855 (N_11855,N_7891,N_8245);
nor U11856 (N_11856,N_7424,N_6372);
or U11857 (N_11857,N_6699,N_7281);
or U11858 (N_11858,N_9339,N_7579);
or U11859 (N_11859,N_6664,N_8589);
or U11860 (N_11860,N_8640,N_8666);
and U11861 (N_11861,N_9172,N_8800);
xnor U11862 (N_11862,N_6638,N_7257);
or U11863 (N_11863,N_8658,N_7770);
or U11864 (N_11864,N_9161,N_7832);
nand U11865 (N_11865,N_8495,N_7340);
xor U11866 (N_11866,N_7527,N_8370);
nor U11867 (N_11867,N_6532,N_7487);
nand U11868 (N_11868,N_6384,N_7534);
nand U11869 (N_11869,N_8757,N_7157);
and U11870 (N_11870,N_8360,N_8405);
or U11871 (N_11871,N_8573,N_7161);
xnor U11872 (N_11872,N_6995,N_9351);
nor U11873 (N_11873,N_6621,N_7285);
nand U11874 (N_11874,N_7426,N_6689);
and U11875 (N_11875,N_6651,N_7130);
nor U11876 (N_11876,N_9335,N_8109);
or U11877 (N_11877,N_6545,N_9015);
nor U11878 (N_11878,N_9284,N_9286);
nand U11879 (N_11879,N_7984,N_6277);
xor U11880 (N_11880,N_6909,N_6344);
nor U11881 (N_11881,N_9168,N_7283);
nor U11882 (N_11882,N_6993,N_8974);
nor U11883 (N_11883,N_8798,N_6525);
nand U11884 (N_11884,N_8549,N_8490);
or U11885 (N_11885,N_8934,N_7073);
xor U11886 (N_11886,N_7481,N_6537);
nor U11887 (N_11887,N_6806,N_7123);
nand U11888 (N_11888,N_7100,N_8604);
nand U11889 (N_11889,N_9205,N_9297);
nor U11890 (N_11890,N_7311,N_7348);
nor U11891 (N_11891,N_8019,N_7821);
xnor U11892 (N_11892,N_9362,N_6511);
or U11893 (N_11893,N_6787,N_8476);
and U11894 (N_11894,N_8203,N_8375);
or U11895 (N_11895,N_8108,N_6891);
nor U11896 (N_11896,N_7100,N_9342);
and U11897 (N_11897,N_9161,N_8146);
xor U11898 (N_11898,N_8839,N_7614);
or U11899 (N_11899,N_7664,N_9242);
nor U11900 (N_11900,N_6895,N_8333);
and U11901 (N_11901,N_9035,N_6782);
and U11902 (N_11902,N_8505,N_7530);
nor U11903 (N_11903,N_6420,N_7040);
nor U11904 (N_11904,N_6668,N_6594);
and U11905 (N_11905,N_6889,N_7287);
nand U11906 (N_11906,N_7865,N_7178);
and U11907 (N_11907,N_9293,N_6906);
and U11908 (N_11908,N_7832,N_6592);
nor U11909 (N_11909,N_6719,N_8302);
or U11910 (N_11910,N_6346,N_6909);
xor U11911 (N_11911,N_6945,N_8120);
or U11912 (N_11912,N_8397,N_8448);
nand U11913 (N_11913,N_7390,N_6584);
nand U11914 (N_11914,N_8937,N_6645);
and U11915 (N_11915,N_9106,N_8306);
and U11916 (N_11916,N_7381,N_7644);
xnor U11917 (N_11917,N_6629,N_8776);
nor U11918 (N_11918,N_8076,N_8389);
nand U11919 (N_11919,N_8346,N_7928);
nand U11920 (N_11920,N_8549,N_7983);
nor U11921 (N_11921,N_8551,N_8258);
xnor U11922 (N_11922,N_7601,N_6431);
nand U11923 (N_11923,N_9048,N_9002);
nor U11924 (N_11924,N_7264,N_8049);
xnor U11925 (N_11925,N_7866,N_7749);
or U11926 (N_11926,N_6821,N_6328);
nand U11927 (N_11927,N_8663,N_7608);
and U11928 (N_11928,N_8153,N_9012);
nand U11929 (N_11929,N_6283,N_9015);
nor U11930 (N_11930,N_7894,N_8765);
nor U11931 (N_11931,N_7227,N_9079);
nor U11932 (N_11932,N_9159,N_7194);
xor U11933 (N_11933,N_6613,N_8197);
nor U11934 (N_11934,N_6329,N_9308);
nand U11935 (N_11935,N_8062,N_7999);
xnor U11936 (N_11936,N_7935,N_8509);
nor U11937 (N_11937,N_6577,N_7953);
nor U11938 (N_11938,N_8065,N_8525);
nand U11939 (N_11939,N_8612,N_7489);
nand U11940 (N_11940,N_7726,N_8814);
nor U11941 (N_11941,N_6714,N_8616);
nand U11942 (N_11942,N_7249,N_6252);
or U11943 (N_11943,N_7007,N_7778);
nor U11944 (N_11944,N_7965,N_8725);
and U11945 (N_11945,N_8668,N_8531);
or U11946 (N_11946,N_8014,N_7487);
nand U11947 (N_11947,N_7375,N_8782);
and U11948 (N_11948,N_6771,N_7351);
nor U11949 (N_11949,N_6449,N_6592);
xnor U11950 (N_11950,N_8602,N_6707);
nor U11951 (N_11951,N_8632,N_8782);
nand U11952 (N_11952,N_8585,N_7716);
nand U11953 (N_11953,N_8286,N_6995);
and U11954 (N_11954,N_7697,N_7714);
or U11955 (N_11955,N_6350,N_7087);
nor U11956 (N_11956,N_8410,N_8821);
xor U11957 (N_11957,N_8759,N_6897);
nor U11958 (N_11958,N_6759,N_7704);
nand U11959 (N_11959,N_8526,N_6396);
nor U11960 (N_11960,N_6544,N_6822);
nor U11961 (N_11961,N_7519,N_6363);
and U11962 (N_11962,N_8838,N_6681);
or U11963 (N_11963,N_8140,N_7123);
and U11964 (N_11964,N_7585,N_9111);
nand U11965 (N_11965,N_6703,N_6971);
or U11966 (N_11966,N_6703,N_7221);
and U11967 (N_11967,N_7374,N_9294);
nor U11968 (N_11968,N_8932,N_9366);
nor U11969 (N_11969,N_7448,N_8974);
and U11970 (N_11970,N_8425,N_8266);
xor U11971 (N_11971,N_6652,N_8976);
xor U11972 (N_11972,N_6916,N_7964);
or U11973 (N_11973,N_6882,N_8703);
or U11974 (N_11974,N_9035,N_7098);
or U11975 (N_11975,N_6431,N_9292);
nand U11976 (N_11976,N_7067,N_7100);
or U11977 (N_11977,N_8170,N_7936);
nand U11978 (N_11978,N_6844,N_7902);
xor U11979 (N_11979,N_8099,N_6314);
or U11980 (N_11980,N_8965,N_6455);
nand U11981 (N_11981,N_8921,N_6687);
or U11982 (N_11982,N_6387,N_8884);
nor U11983 (N_11983,N_7186,N_8488);
and U11984 (N_11984,N_8693,N_8449);
nand U11985 (N_11985,N_8898,N_8138);
nor U11986 (N_11986,N_7096,N_7514);
nand U11987 (N_11987,N_8635,N_8388);
nor U11988 (N_11988,N_7571,N_7864);
and U11989 (N_11989,N_7472,N_8819);
nor U11990 (N_11990,N_6452,N_8897);
xor U11991 (N_11991,N_7338,N_6815);
nand U11992 (N_11992,N_7208,N_7759);
nand U11993 (N_11993,N_9310,N_9317);
or U11994 (N_11994,N_7432,N_9198);
and U11995 (N_11995,N_7428,N_8147);
or U11996 (N_11996,N_6381,N_9275);
nor U11997 (N_11997,N_6870,N_6472);
and U11998 (N_11998,N_7803,N_7677);
and U11999 (N_11999,N_6911,N_7015);
nand U12000 (N_12000,N_8500,N_7283);
nand U12001 (N_12001,N_8242,N_6867);
nor U12002 (N_12002,N_6658,N_7113);
nand U12003 (N_12003,N_9284,N_6257);
nor U12004 (N_12004,N_9206,N_8133);
nand U12005 (N_12005,N_7902,N_9104);
and U12006 (N_12006,N_7076,N_9334);
nor U12007 (N_12007,N_8324,N_6788);
nand U12008 (N_12008,N_9083,N_6523);
nand U12009 (N_12009,N_7207,N_8824);
or U12010 (N_12010,N_6268,N_6433);
or U12011 (N_12011,N_7495,N_6669);
or U12012 (N_12012,N_6832,N_6836);
and U12013 (N_12013,N_7312,N_6445);
or U12014 (N_12014,N_8444,N_6452);
and U12015 (N_12015,N_8826,N_8984);
nor U12016 (N_12016,N_7219,N_7567);
or U12017 (N_12017,N_8259,N_8420);
and U12018 (N_12018,N_7665,N_7108);
or U12019 (N_12019,N_6855,N_7775);
xor U12020 (N_12020,N_7765,N_7562);
nor U12021 (N_12021,N_8836,N_8707);
nand U12022 (N_12022,N_8072,N_8766);
nor U12023 (N_12023,N_6449,N_6278);
or U12024 (N_12024,N_8595,N_7763);
nor U12025 (N_12025,N_9263,N_8177);
nand U12026 (N_12026,N_9208,N_8200);
or U12027 (N_12027,N_6697,N_8887);
and U12028 (N_12028,N_7650,N_7366);
nand U12029 (N_12029,N_6456,N_8203);
or U12030 (N_12030,N_7015,N_7010);
and U12031 (N_12031,N_6820,N_8912);
or U12032 (N_12032,N_6784,N_6814);
xor U12033 (N_12033,N_8917,N_8370);
or U12034 (N_12034,N_7511,N_7272);
nand U12035 (N_12035,N_8801,N_7167);
or U12036 (N_12036,N_8845,N_6680);
nand U12037 (N_12037,N_7610,N_7321);
nand U12038 (N_12038,N_6576,N_7501);
or U12039 (N_12039,N_9320,N_8638);
or U12040 (N_12040,N_6889,N_6336);
and U12041 (N_12041,N_8641,N_8839);
or U12042 (N_12042,N_7580,N_7650);
nand U12043 (N_12043,N_7652,N_8252);
or U12044 (N_12044,N_6402,N_7369);
or U12045 (N_12045,N_7942,N_6524);
nand U12046 (N_12046,N_7390,N_7631);
and U12047 (N_12047,N_7195,N_6691);
and U12048 (N_12048,N_7754,N_6995);
xnor U12049 (N_12049,N_6876,N_8558);
and U12050 (N_12050,N_7062,N_6840);
or U12051 (N_12051,N_7429,N_8010);
and U12052 (N_12052,N_6625,N_6828);
and U12053 (N_12053,N_8736,N_9294);
and U12054 (N_12054,N_8899,N_6325);
nand U12055 (N_12055,N_6750,N_7101);
nand U12056 (N_12056,N_6554,N_6275);
and U12057 (N_12057,N_6252,N_7141);
nor U12058 (N_12058,N_7702,N_7402);
nand U12059 (N_12059,N_7045,N_8203);
and U12060 (N_12060,N_6842,N_7524);
or U12061 (N_12061,N_7356,N_8674);
and U12062 (N_12062,N_8012,N_8339);
nor U12063 (N_12063,N_8588,N_9036);
nor U12064 (N_12064,N_8495,N_7520);
nor U12065 (N_12065,N_6379,N_6266);
nand U12066 (N_12066,N_8735,N_8186);
or U12067 (N_12067,N_6689,N_8315);
or U12068 (N_12068,N_8272,N_8354);
nor U12069 (N_12069,N_7003,N_9288);
or U12070 (N_12070,N_8429,N_7925);
nor U12071 (N_12071,N_7872,N_8695);
or U12072 (N_12072,N_6474,N_9178);
nor U12073 (N_12073,N_6812,N_8580);
and U12074 (N_12074,N_8310,N_7073);
nand U12075 (N_12075,N_6726,N_7375);
or U12076 (N_12076,N_7878,N_8760);
nand U12077 (N_12077,N_8667,N_7376);
nor U12078 (N_12078,N_8748,N_8546);
and U12079 (N_12079,N_7525,N_7270);
or U12080 (N_12080,N_7933,N_8169);
nor U12081 (N_12081,N_6962,N_8805);
or U12082 (N_12082,N_7991,N_9023);
nor U12083 (N_12083,N_8631,N_6448);
xor U12084 (N_12084,N_6529,N_9268);
nand U12085 (N_12085,N_6841,N_8992);
nor U12086 (N_12086,N_6841,N_6468);
and U12087 (N_12087,N_6400,N_7061);
and U12088 (N_12088,N_6944,N_6741);
or U12089 (N_12089,N_7131,N_6319);
nand U12090 (N_12090,N_8661,N_7612);
nand U12091 (N_12091,N_9180,N_8095);
and U12092 (N_12092,N_8705,N_7884);
nand U12093 (N_12093,N_7453,N_8892);
nand U12094 (N_12094,N_6802,N_8630);
and U12095 (N_12095,N_7179,N_9043);
nor U12096 (N_12096,N_8195,N_7277);
or U12097 (N_12097,N_9017,N_8376);
nor U12098 (N_12098,N_8315,N_7935);
nand U12099 (N_12099,N_8283,N_7662);
xnor U12100 (N_12100,N_6296,N_9233);
and U12101 (N_12101,N_8234,N_8255);
nand U12102 (N_12102,N_8282,N_9114);
nand U12103 (N_12103,N_8316,N_6507);
and U12104 (N_12104,N_6897,N_7264);
nand U12105 (N_12105,N_8617,N_7727);
nand U12106 (N_12106,N_7135,N_7718);
or U12107 (N_12107,N_7124,N_7692);
nand U12108 (N_12108,N_7775,N_6755);
nor U12109 (N_12109,N_7892,N_6997);
nor U12110 (N_12110,N_6492,N_7026);
or U12111 (N_12111,N_6891,N_8005);
nor U12112 (N_12112,N_9288,N_9158);
and U12113 (N_12113,N_6893,N_7193);
and U12114 (N_12114,N_9161,N_8345);
xor U12115 (N_12115,N_7374,N_6364);
or U12116 (N_12116,N_8853,N_6747);
nand U12117 (N_12117,N_8108,N_8307);
nand U12118 (N_12118,N_9262,N_8885);
or U12119 (N_12119,N_8123,N_9089);
xor U12120 (N_12120,N_8842,N_7482);
and U12121 (N_12121,N_7687,N_8470);
nand U12122 (N_12122,N_9217,N_8566);
and U12123 (N_12123,N_8358,N_6884);
nor U12124 (N_12124,N_9070,N_6892);
or U12125 (N_12125,N_7018,N_8904);
nand U12126 (N_12126,N_7375,N_7941);
or U12127 (N_12127,N_7471,N_8021);
nor U12128 (N_12128,N_6571,N_8416);
nor U12129 (N_12129,N_7182,N_6966);
or U12130 (N_12130,N_8777,N_7787);
nor U12131 (N_12131,N_8078,N_6815);
xnor U12132 (N_12132,N_7912,N_6607);
nand U12133 (N_12133,N_8540,N_9191);
nor U12134 (N_12134,N_7921,N_6589);
and U12135 (N_12135,N_6941,N_7085);
or U12136 (N_12136,N_8889,N_8952);
xnor U12137 (N_12137,N_9259,N_7222);
nor U12138 (N_12138,N_9123,N_9079);
nand U12139 (N_12139,N_8104,N_8482);
nor U12140 (N_12140,N_9184,N_8051);
or U12141 (N_12141,N_7582,N_6403);
nor U12142 (N_12142,N_7180,N_8421);
nand U12143 (N_12143,N_7775,N_7834);
nand U12144 (N_12144,N_8940,N_8348);
nor U12145 (N_12145,N_8367,N_6855);
and U12146 (N_12146,N_7553,N_6636);
nor U12147 (N_12147,N_9286,N_6924);
or U12148 (N_12148,N_8367,N_9364);
nor U12149 (N_12149,N_6459,N_8101);
nor U12150 (N_12150,N_9011,N_6372);
or U12151 (N_12151,N_6517,N_7643);
or U12152 (N_12152,N_8088,N_6546);
nor U12153 (N_12153,N_8093,N_7522);
xnor U12154 (N_12154,N_9075,N_6487);
or U12155 (N_12155,N_6757,N_8370);
or U12156 (N_12156,N_7554,N_8253);
or U12157 (N_12157,N_8681,N_6454);
and U12158 (N_12158,N_8636,N_6401);
nor U12159 (N_12159,N_8462,N_9189);
and U12160 (N_12160,N_8473,N_9322);
nand U12161 (N_12161,N_6568,N_7437);
and U12162 (N_12162,N_6779,N_6543);
and U12163 (N_12163,N_6754,N_6345);
or U12164 (N_12164,N_7558,N_8817);
nand U12165 (N_12165,N_7272,N_8659);
nor U12166 (N_12166,N_8715,N_6989);
and U12167 (N_12167,N_9065,N_7955);
and U12168 (N_12168,N_6659,N_6283);
nand U12169 (N_12169,N_6644,N_8275);
nor U12170 (N_12170,N_7100,N_9104);
nor U12171 (N_12171,N_6469,N_8282);
or U12172 (N_12172,N_8151,N_8640);
nand U12173 (N_12173,N_7950,N_8188);
xor U12174 (N_12174,N_8612,N_9043);
xor U12175 (N_12175,N_7292,N_6316);
and U12176 (N_12176,N_7878,N_7271);
nor U12177 (N_12177,N_7711,N_9366);
nor U12178 (N_12178,N_8758,N_8507);
or U12179 (N_12179,N_6269,N_8684);
nand U12180 (N_12180,N_8382,N_7834);
nor U12181 (N_12181,N_8991,N_6395);
nand U12182 (N_12182,N_7611,N_7674);
and U12183 (N_12183,N_6640,N_6971);
nand U12184 (N_12184,N_7796,N_7512);
nor U12185 (N_12185,N_7170,N_7631);
nand U12186 (N_12186,N_9048,N_6296);
nor U12187 (N_12187,N_7044,N_9163);
and U12188 (N_12188,N_6636,N_7175);
nor U12189 (N_12189,N_8674,N_8886);
nor U12190 (N_12190,N_8678,N_9304);
or U12191 (N_12191,N_8940,N_8054);
nand U12192 (N_12192,N_7453,N_7556);
nand U12193 (N_12193,N_7505,N_7115);
nor U12194 (N_12194,N_7996,N_9094);
nand U12195 (N_12195,N_6328,N_6482);
or U12196 (N_12196,N_8278,N_8320);
or U12197 (N_12197,N_7510,N_9120);
nand U12198 (N_12198,N_8847,N_6295);
nor U12199 (N_12199,N_8343,N_6362);
or U12200 (N_12200,N_7107,N_7390);
xor U12201 (N_12201,N_6815,N_7613);
or U12202 (N_12202,N_8105,N_7113);
xor U12203 (N_12203,N_7298,N_9003);
and U12204 (N_12204,N_6574,N_6942);
nor U12205 (N_12205,N_8219,N_7704);
or U12206 (N_12206,N_7142,N_8102);
or U12207 (N_12207,N_7863,N_6643);
nor U12208 (N_12208,N_6443,N_8310);
or U12209 (N_12209,N_9124,N_8601);
nand U12210 (N_12210,N_7303,N_8984);
or U12211 (N_12211,N_7408,N_7043);
nor U12212 (N_12212,N_7781,N_8853);
nand U12213 (N_12213,N_7667,N_9060);
nor U12214 (N_12214,N_9227,N_7363);
or U12215 (N_12215,N_7068,N_9289);
nor U12216 (N_12216,N_8540,N_6445);
nor U12217 (N_12217,N_8279,N_7708);
nor U12218 (N_12218,N_8277,N_7198);
and U12219 (N_12219,N_6674,N_8814);
nand U12220 (N_12220,N_9091,N_9008);
xor U12221 (N_12221,N_7959,N_8842);
or U12222 (N_12222,N_8209,N_8300);
nor U12223 (N_12223,N_9198,N_8667);
and U12224 (N_12224,N_7932,N_7544);
xnor U12225 (N_12225,N_8884,N_6959);
nor U12226 (N_12226,N_8499,N_7021);
and U12227 (N_12227,N_6607,N_7717);
nor U12228 (N_12228,N_6889,N_6811);
nand U12229 (N_12229,N_7892,N_9050);
xor U12230 (N_12230,N_8724,N_6828);
or U12231 (N_12231,N_7289,N_7679);
and U12232 (N_12232,N_8085,N_7052);
or U12233 (N_12233,N_8596,N_6641);
nor U12234 (N_12234,N_8144,N_7774);
nand U12235 (N_12235,N_8229,N_8749);
or U12236 (N_12236,N_6974,N_9033);
and U12237 (N_12237,N_7009,N_7366);
nand U12238 (N_12238,N_7743,N_7929);
xor U12239 (N_12239,N_8041,N_9055);
and U12240 (N_12240,N_9336,N_8375);
and U12241 (N_12241,N_6727,N_6735);
and U12242 (N_12242,N_9123,N_7185);
or U12243 (N_12243,N_8600,N_8694);
nand U12244 (N_12244,N_8775,N_7920);
nor U12245 (N_12245,N_8824,N_8541);
nand U12246 (N_12246,N_8189,N_6949);
or U12247 (N_12247,N_9189,N_7007);
and U12248 (N_12248,N_9078,N_8387);
nand U12249 (N_12249,N_9106,N_7103);
nor U12250 (N_12250,N_6869,N_8326);
nor U12251 (N_12251,N_9137,N_8019);
nand U12252 (N_12252,N_9348,N_9038);
nand U12253 (N_12253,N_8368,N_7669);
nand U12254 (N_12254,N_6419,N_9063);
or U12255 (N_12255,N_6422,N_8130);
nor U12256 (N_12256,N_7521,N_8424);
nor U12257 (N_12257,N_6299,N_7457);
nand U12258 (N_12258,N_8915,N_6853);
or U12259 (N_12259,N_8135,N_7267);
xnor U12260 (N_12260,N_9005,N_6314);
and U12261 (N_12261,N_6788,N_6580);
nand U12262 (N_12262,N_8909,N_8751);
nor U12263 (N_12263,N_8281,N_8769);
or U12264 (N_12264,N_8061,N_6504);
and U12265 (N_12265,N_8247,N_7741);
and U12266 (N_12266,N_7831,N_8789);
nor U12267 (N_12267,N_7834,N_7326);
nor U12268 (N_12268,N_7211,N_7197);
nand U12269 (N_12269,N_7238,N_7751);
or U12270 (N_12270,N_9151,N_6617);
or U12271 (N_12271,N_8326,N_7245);
nand U12272 (N_12272,N_9355,N_7284);
xnor U12273 (N_12273,N_7344,N_9348);
nor U12274 (N_12274,N_7362,N_7376);
xor U12275 (N_12275,N_8716,N_7163);
and U12276 (N_12276,N_8795,N_7061);
and U12277 (N_12277,N_7464,N_7888);
and U12278 (N_12278,N_9238,N_8987);
nand U12279 (N_12279,N_8459,N_9042);
nand U12280 (N_12280,N_7596,N_6931);
xnor U12281 (N_12281,N_8846,N_8287);
or U12282 (N_12282,N_7294,N_8174);
nor U12283 (N_12283,N_7105,N_7227);
nand U12284 (N_12284,N_7074,N_6415);
or U12285 (N_12285,N_8370,N_8155);
and U12286 (N_12286,N_9116,N_7272);
xor U12287 (N_12287,N_8243,N_7870);
nand U12288 (N_12288,N_7512,N_9191);
nand U12289 (N_12289,N_6269,N_8315);
and U12290 (N_12290,N_7823,N_8200);
nor U12291 (N_12291,N_7037,N_8533);
and U12292 (N_12292,N_8994,N_7436);
xnor U12293 (N_12293,N_7321,N_7257);
nor U12294 (N_12294,N_9237,N_8394);
nor U12295 (N_12295,N_7132,N_8627);
nor U12296 (N_12296,N_9299,N_7334);
xor U12297 (N_12297,N_7251,N_6400);
or U12298 (N_12298,N_8571,N_9038);
or U12299 (N_12299,N_6956,N_8406);
and U12300 (N_12300,N_7541,N_6481);
and U12301 (N_12301,N_6291,N_8055);
or U12302 (N_12302,N_6526,N_9311);
and U12303 (N_12303,N_8429,N_8548);
or U12304 (N_12304,N_6698,N_7655);
nand U12305 (N_12305,N_6349,N_7833);
nor U12306 (N_12306,N_6761,N_8810);
or U12307 (N_12307,N_7186,N_8691);
or U12308 (N_12308,N_7743,N_6912);
nor U12309 (N_12309,N_8708,N_8000);
or U12310 (N_12310,N_6703,N_8339);
nand U12311 (N_12311,N_6997,N_8335);
nor U12312 (N_12312,N_6572,N_9278);
xor U12313 (N_12313,N_8650,N_8967);
nor U12314 (N_12314,N_8248,N_8820);
and U12315 (N_12315,N_8915,N_8413);
nand U12316 (N_12316,N_8816,N_6294);
and U12317 (N_12317,N_9001,N_7692);
and U12318 (N_12318,N_6867,N_6505);
nor U12319 (N_12319,N_7122,N_8552);
nor U12320 (N_12320,N_7186,N_8660);
nor U12321 (N_12321,N_7770,N_7879);
and U12322 (N_12322,N_7780,N_6321);
nor U12323 (N_12323,N_8302,N_8506);
nor U12324 (N_12324,N_8607,N_6354);
and U12325 (N_12325,N_8274,N_6698);
and U12326 (N_12326,N_7567,N_7827);
and U12327 (N_12327,N_7131,N_7655);
and U12328 (N_12328,N_9138,N_7220);
and U12329 (N_12329,N_8679,N_8524);
nor U12330 (N_12330,N_7266,N_7020);
nand U12331 (N_12331,N_8742,N_9064);
or U12332 (N_12332,N_7705,N_8332);
xnor U12333 (N_12333,N_7627,N_8684);
and U12334 (N_12334,N_6400,N_8080);
or U12335 (N_12335,N_9106,N_7542);
nand U12336 (N_12336,N_8295,N_9020);
xor U12337 (N_12337,N_6271,N_8531);
xnor U12338 (N_12338,N_8935,N_9319);
xnor U12339 (N_12339,N_9126,N_8012);
and U12340 (N_12340,N_8046,N_8302);
nor U12341 (N_12341,N_7334,N_8436);
and U12342 (N_12342,N_8718,N_7955);
and U12343 (N_12343,N_6648,N_8489);
xor U12344 (N_12344,N_6332,N_7595);
or U12345 (N_12345,N_7226,N_7171);
or U12346 (N_12346,N_9314,N_7780);
xor U12347 (N_12347,N_7801,N_8824);
nor U12348 (N_12348,N_8603,N_8532);
nor U12349 (N_12349,N_7230,N_7421);
and U12350 (N_12350,N_7391,N_6616);
or U12351 (N_12351,N_9209,N_8078);
or U12352 (N_12352,N_9230,N_6628);
nand U12353 (N_12353,N_8213,N_7876);
or U12354 (N_12354,N_6940,N_6550);
nand U12355 (N_12355,N_6373,N_8552);
or U12356 (N_12356,N_7066,N_6558);
and U12357 (N_12357,N_9322,N_6898);
xor U12358 (N_12358,N_8959,N_6932);
nand U12359 (N_12359,N_9312,N_7253);
nand U12360 (N_12360,N_7615,N_6417);
and U12361 (N_12361,N_8217,N_6415);
nand U12362 (N_12362,N_7573,N_8446);
nand U12363 (N_12363,N_6723,N_7943);
nand U12364 (N_12364,N_6889,N_9262);
or U12365 (N_12365,N_7897,N_6540);
and U12366 (N_12366,N_8059,N_6761);
and U12367 (N_12367,N_6900,N_8333);
and U12368 (N_12368,N_6655,N_8425);
and U12369 (N_12369,N_7731,N_8423);
nand U12370 (N_12370,N_7989,N_7593);
nand U12371 (N_12371,N_7555,N_8619);
and U12372 (N_12372,N_7621,N_6765);
nand U12373 (N_12373,N_8672,N_7530);
and U12374 (N_12374,N_8055,N_8827);
or U12375 (N_12375,N_8865,N_6488);
nand U12376 (N_12376,N_7814,N_8121);
or U12377 (N_12377,N_6814,N_8682);
nand U12378 (N_12378,N_6631,N_8785);
and U12379 (N_12379,N_7652,N_8487);
nand U12380 (N_12380,N_6644,N_7152);
nand U12381 (N_12381,N_7483,N_7120);
and U12382 (N_12382,N_8797,N_6737);
or U12383 (N_12383,N_6367,N_7101);
and U12384 (N_12384,N_7693,N_6443);
or U12385 (N_12385,N_7500,N_7167);
nor U12386 (N_12386,N_8878,N_8163);
nor U12387 (N_12387,N_7852,N_6380);
and U12388 (N_12388,N_6807,N_9348);
nand U12389 (N_12389,N_8003,N_6477);
xnor U12390 (N_12390,N_8372,N_7662);
nor U12391 (N_12391,N_9064,N_8606);
xnor U12392 (N_12392,N_7039,N_8531);
or U12393 (N_12393,N_7793,N_6772);
xor U12394 (N_12394,N_9284,N_7669);
nand U12395 (N_12395,N_6739,N_8451);
nor U12396 (N_12396,N_7623,N_7409);
xor U12397 (N_12397,N_7292,N_7922);
nor U12398 (N_12398,N_6695,N_7949);
and U12399 (N_12399,N_8071,N_8238);
xor U12400 (N_12400,N_6267,N_6608);
and U12401 (N_12401,N_7197,N_8597);
and U12402 (N_12402,N_8091,N_9048);
or U12403 (N_12403,N_6644,N_8286);
xor U12404 (N_12404,N_6938,N_7647);
or U12405 (N_12405,N_6926,N_8439);
and U12406 (N_12406,N_8318,N_8249);
and U12407 (N_12407,N_8367,N_9164);
nor U12408 (N_12408,N_7659,N_6257);
nand U12409 (N_12409,N_8285,N_6436);
or U12410 (N_12410,N_7316,N_8857);
nor U12411 (N_12411,N_9290,N_7712);
nor U12412 (N_12412,N_9109,N_9171);
nand U12413 (N_12413,N_9338,N_7365);
nand U12414 (N_12414,N_6388,N_7691);
or U12415 (N_12415,N_6942,N_6702);
xor U12416 (N_12416,N_7905,N_7255);
or U12417 (N_12417,N_7035,N_8991);
nand U12418 (N_12418,N_6522,N_7160);
nor U12419 (N_12419,N_7009,N_8878);
or U12420 (N_12420,N_6325,N_8168);
and U12421 (N_12421,N_7680,N_7126);
nor U12422 (N_12422,N_7509,N_8461);
nor U12423 (N_12423,N_6824,N_6407);
and U12424 (N_12424,N_7107,N_6950);
nor U12425 (N_12425,N_9291,N_7312);
nand U12426 (N_12426,N_7750,N_8740);
nand U12427 (N_12427,N_8070,N_8571);
nand U12428 (N_12428,N_8653,N_8520);
or U12429 (N_12429,N_6750,N_8445);
nor U12430 (N_12430,N_8779,N_9310);
nor U12431 (N_12431,N_8896,N_7402);
nand U12432 (N_12432,N_7240,N_9126);
or U12433 (N_12433,N_7442,N_7970);
nor U12434 (N_12434,N_9090,N_9084);
nand U12435 (N_12435,N_6673,N_7577);
nor U12436 (N_12436,N_8847,N_6987);
nand U12437 (N_12437,N_8772,N_7654);
and U12438 (N_12438,N_7790,N_6335);
and U12439 (N_12439,N_7897,N_8406);
nand U12440 (N_12440,N_7072,N_9329);
or U12441 (N_12441,N_7622,N_9056);
and U12442 (N_12442,N_8979,N_6288);
and U12443 (N_12443,N_8246,N_9151);
and U12444 (N_12444,N_7539,N_9275);
nand U12445 (N_12445,N_6764,N_7950);
xor U12446 (N_12446,N_9107,N_9213);
or U12447 (N_12447,N_8484,N_8834);
nand U12448 (N_12448,N_7941,N_8766);
or U12449 (N_12449,N_6262,N_7662);
and U12450 (N_12450,N_7967,N_6985);
xor U12451 (N_12451,N_6906,N_9087);
nand U12452 (N_12452,N_6853,N_6258);
nor U12453 (N_12453,N_6554,N_6450);
nand U12454 (N_12454,N_8346,N_8762);
and U12455 (N_12455,N_6892,N_8495);
nor U12456 (N_12456,N_7307,N_6917);
or U12457 (N_12457,N_7961,N_6905);
nand U12458 (N_12458,N_8137,N_9269);
or U12459 (N_12459,N_7623,N_6292);
nand U12460 (N_12460,N_7851,N_8164);
nor U12461 (N_12461,N_7565,N_7562);
or U12462 (N_12462,N_7068,N_8759);
and U12463 (N_12463,N_7447,N_9240);
or U12464 (N_12464,N_6549,N_7038);
nand U12465 (N_12465,N_7076,N_7050);
xnor U12466 (N_12466,N_8065,N_7069);
xnor U12467 (N_12467,N_7734,N_7727);
xnor U12468 (N_12468,N_8610,N_6804);
and U12469 (N_12469,N_8033,N_7308);
and U12470 (N_12470,N_6756,N_6835);
nand U12471 (N_12471,N_7046,N_7336);
nor U12472 (N_12472,N_6340,N_8820);
nand U12473 (N_12473,N_6689,N_8194);
xor U12474 (N_12474,N_9036,N_8784);
and U12475 (N_12475,N_6914,N_8505);
nor U12476 (N_12476,N_7092,N_9073);
nand U12477 (N_12477,N_7182,N_6354);
nand U12478 (N_12478,N_8802,N_6572);
and U12479 (N_12479,N_6369,N_7464);
or U12480 (N_12480,N_6722,N_7059);
or U12481 (N_12481,N_6884,N_8160);
nand U12482 (N_12482,N_7405,N_9218);
nor U12483 (N_12483,N_8383,N_6958);
nor U12484 (N_12484,N_9263,N_8904);
or U12485 (N_12485,N_6825,N_6741);
and U12486 (N_12486,N_9052,N_6571);
or U12487 (N_12487,N_7595,N_8401);
or U12488 (N_12488,N_8339,N_9237);
nor U12489 (N_12489,N_8543,N_7528);
nor U12490 (N_12490,N_6870,N_8696);
and U12491 (N_12491,N_6514,N_8924);
nor U12492 (N_12492,N_6427,N_7809);
nand U12493 (N_12493,N_6996,N_7604);
xnor U12494 (N_12494,N_8061,N_6676);
nor U12495 (N_12495,N_7404,N_8579);
nor U12496 (N_12496,N_7269,N_8199);
and U12497 (N_12497,N_7961,N_8217);
or U12498 (N_12498,N_6765,N_8402);
nor U12499 (N_12499,N_6288,N_7207);
and U12500 (N_12500,N_12060,N_10417);
and U12501 (N_12501,N_11321,N_11175);
nor U12502 (N_12502,N_10444,N_10147);
and U12503 (N_12503,N_11888,N_11902);
and U12504 (N_12504,N_9865,N_12148);
and U12505 (N_12505,N_11935,N_11638);
nand U12506 (N_12506,N_10320,N_11217);
and U12507 (N_12507,N_12013,N_12031);
and U12508 (N_12508,N_9453,N_10152);
xnor U12509 (N_12509,N_11496,N_10921);
or U12510 (N_12510,N_11388,N_11130);
nor U12511 (N_12511,N_11096,N_12214);
xnor U12512 (N_12512,N_12302,N_11667);
nand U12513 (N_12513,N_10594,N_12047);
nand U12514 (N_12514,N_11529,N_11738);
and U12515 (N_12515,N_9950,N_12155);
nand U12516 (N_12516,N_11296,N_10616);
nand U12517 (N_12517,N_12299,N_10584);
nand U12518 (N_12518,N_10556,N_11358);
and U12519 (N_12519,N_10607,N_12254);
nand U12520 (N_12520,N_9910,N_10808);
or U12521 (N_12521,N_10934,N_11752);
or U12522 (N_12522,N_12297,N_11411);
nor U12523 (N_12523,N_11335,N_10819);
nor U12524 (N_12524,N_10781,N_12240);
and U12525 (N_12525,N_11796,N_11723);
and U12526 (N_12526,N_11917,N_9720);
and U12527 (N_12527,N_11025,N_9542);
nor U12528 (N_12528,N_10298,N_10522);
and U12529 (N_12529,N_12029,N_11813);
and U12530 (N_12530,N_11741,N_11979);
or U12531 (N_12531,N_9891,N_10567);
or U12532 (N_12532,N_10125,N_11019);
or U12533 (N_12533,N_10988,N_12475);
xor U12534 (N_12534,N_9468,N_9532);
xnor U12535 (N_12535,N_10318,N_10890);
and U12536 (N_12536,N_10553,N_9637);
or U12537 (N_12537,N_10762,N_11042);
and U12538 (N_12538,N_11870,N_10087);
nor U12539 (N_12539,N_12084,N_11823);
and U12540 (N_12540,N_10914,N_12159);
nor U12541 (N_12541,N_10712,N_10130);
or U12542 (N_12542,N_10515,N_10051);
or U12543 (N_12543,N_11736,N_11181);
xnor U12544 (N_12544,N_11029,N_9424);
nand U12545 (N_12545,N_10721,N_11415);
nand U12546 (N_12546,N_11374,N_11593);
and U12547 (N_12547,N_9899,N_11083);
nor U12548 (N_12548,N_9578,N_11879);
nor U12549 (N_12549,N_10433,N_11255);
nor U12550 (N_12550,N_10327,N_11760);
and U12551 (N_12551,N_9695,N_11474);
xnor U12552 (N_12552,N_10114,N_9837);
xor U12553 (N_12553,N_10123,N_12173);
nor U12554 (N_12554,N_10279,N_11419);
xnor U12555 (N_12555,N_10012,N_10590);
nand U12556 (N_12556,N_10221,N_10291);
nand U12557 (N_12557,N_10403,N_11595);
nor U12558 (N_12558,N_9987,N_11163);
and U12559 (N_12559,N_11174,N_10432);
nand U12560 (N_12560,N_9477,N_11924);
nor U12561 (N_12561,N_11500,N_10948);
or U12562 (N_12562,N_10927,N_10782);
nor U12563 (N_12563,N_9408,N_9996);
and U12564 (N_12564,N_9587,N_10027);
or U12565 (N_12565,N_9428,N_11471);
or U12566 (N_12566,N_11395,N_10053);
xnor U12567 (N_12567,N_11674,N_11624);
and U12568 (N_12568,N_10570,N_11768);
nor U12569 (N_12569,N_9631,N_10950);
xor U12570 (N_12570,N_9449,N_12014);
nor U12571 (N_12571,N_10095,N_12028);
or U12572 (N_12572,N_11905,N_9973);
xor U12573 (N_12573,N_11722,N_10600);
and U12574 (N_12574,N_9692,N_11584);
nand U12575 (N_12575,N_9828,N_10230);
nand U12576 (N_12576,N_9875,N_11837);
nand U12577 (N_12577,N_10835,N_9400);
xor U12578 (N_12578,N_11568,N_9502);
and U12579 (N_12579,N_10823,N_10943);
or U12580 (N_12580,N_9858,N_9434);
and U12581 (N_12581,N_10771,N_9783);
nand U12582 (N_12582,N_11880,N_10597);
or U12583 (N_12583,N_10818,N_9755);
nand U12584 (N_12584,N_11137,N_12382);
xnor U12585 (N_12585,N_9618,N_11835);
and U12586 (N_12586,N_10218,N_11060);
and U12587 (N_12587,N_12459,N_12243);
nand U12588 (N_12588,N_10375,N_10280);
or U12589 (N_12589,N_10655,N_9677);
and U12590 (N_12590,N_9616,N_11518);
nor U12591 (N_12591,N_10357,N_11819);
nand U12592 (N_12592,N_11754,N_11913);
nand U12593 (N_12593,N_11931,N_10962);
nor U12594 (N_12594,N_9398,N_11352);
nor U12595 (N_12595,N_11596,N_10270);
nand U12596 (N_12596,N_9665,N_9403);
and U12597 (N_12597,N_11273,N_11483);
or U12598 (N_12598,N_10732,N_10228);
nand U12599 (N_12599,N_9793,N_9597);
nand U12600 (N_12600,N_12094,N_10997);
and U12601 (N_12601,N_10376,N_11930);
nand U12602 (N_12602,N_12268,N_11489);
xor U12603 (N_12603,N_11330,N_11767);
and U12604 (N_12604,N_10811,N_9620);
or U12605 (N_12605,N_12193,N_10901);
or U12606 (N_12606,N_11550,N_9523);
nand U12607 (N_12607,N_9820,N_10408);
nand U12608 (N_12608,N_10677,N_10873);
nand U12609 (N_12609,N_10679,N_11460);
and U12610 (N_12610,N_9421,N_12386);
and U12611 (N_12611,N_10731,N_10705);
and U12612 (N_12612,N_9409,N_12183);
nand U12613 (N_12613,N_11574,N_9581);
and U12614 (N_12614,N_10586,N_12309);
nor U12615 (N_12615,N_11438,N_9739);
xnor U12616 (N_12616,N_9456,N_11322);
or U12617 (N_12617,N_11619,N_9507);
nand U12618 (N_12618,N_9498,N_12334);
nor U12619 (N_12619,N_11805,N_9876);
or U12620 (N_12620,N_11963,N_12341);
or U12621 (N_12621,N_11166,N_12153);
or U12622 (N_12622,N_11037,N_10973);
nand U12623 (N_12623,N_10702,N_11956);
nand U12624 (N_12624,N_11349,N_10879);
nand U12625 (N_12625,N_10502,N_9426);
nand U12626 (N_12626,N_10954,N_10529);
nor U12627 (N_12627,N_9638,N_11587);
nand U12628 (N_12628,N_10313,N_12172);
nand U12629 (N_12629,N_12336,N_10391);
and U12630 (N_12630,N_10370,N_12087);
or U12631 (N_12631,N_10420,N_10534);
and U12632 (N_12632,N_9853,N_11565);
or U12633 (N_12633,N_12121,N_10636);
nor U12634 (N_12634,N_12131,N_10812);
and U12635 (N_12635,N_11197,N_9981);
nand U12636 (N_12636,N_11633,N_11762);
or U12637 (N_12637,N_9656,N_10457);
or U12638 (N_12638,N_12467,N_11094);
nor U12639 (N_12639,N_10964,N_10955);
or U12640 (N_12640,N_11193,N_10458);
or U12641 (N_12641,N_12303,N_10929);
and U12642 (N_12642,N_11338,N_11729);
nand U12643 (N_12643,N_12204,N_11229);
or U12644 (N_12644,N_10387,N_11478);
nand U12645 (N_12645,N_10394,N_10525);
or U12646 (N_12646,N_11781,N_10648);
or U12647 (N_12647,N_12196,N_12317);
nor U12648 (N_12648,N_11831,N_9892);
nor U12649 (N_12649,N_10807,N_9433);
nor U12650 (N_12650,N_9903,N_10514);
or U12651 (N_12651,N_11287,N_11975);
nand U12652 (N_12652,N_11306,N_9405);
or U12653 (N_12653,N_11297,N_10512);
nand U12654 (N_12654,N_11728,N_11689);
and U12655 (N_12655,N_12406,N_12256);
and U12656 (N_12656,N_12053,N_10709);
or U12657 (N_12657,N_11146,N_11016);
xnor U12658 (N_12658,N_9738,N_11898);
nand U12659 (N_12659,N_10959,N_9741);
and U12660 (N_12660,N_12200,N_10090);
nand U12661 (N_12661,N_9752,N_9905);
nor U12662 (N_12662,N_12487,N_11551);
nor U12663 (N_12663,N_11090,N_10797);
or U12664 (N_12664,N_10212,N_9534);
or U12665 (N_12665,N_10855,N_12162);
and U12666 (N_12666,N_10490,N_9880);
nand U12667 (N_12667,N_11402,N_10776);
nand U12668 (N_12668,N_11095,N_11430);
nand U12669 (N_12669,N_9849,N_9926);
and U12670 (N_12670,N_12328,N_11301);
and U12671 (N_12671,N_9480,N_12215);
and U12672 (N_12672,N_10715,N_12481);
and U12673 (N_12673,N_12440,N_12206);
or U12674 (N_12674,N_9866,N_9606);
or U12675 (N_12675,N_12470,N_10034);
nand U12676 (N_12676,N_12128,N_9778);
and U12677 (N_12677,N_10231,N_11708);
and U12678 (N_12678,N_10595,N_9535);
nand U12679 (N_12679,N_10216,N_10907);
or U12680 (N_12680,N_9943,N_11262);
and U12681 (N_12681,N_12154,N_10926);
nor U12682 (N_12682,N_10219,N_12158);
xnor U12683 (N_12683,N_9816,N_10663);
nor U12684 (N_12684,N_11570,N_12147);
or U12685 (N_12685,N_12427,N_11490);
nor U12686 (N_12686,N_10018,N_11050);
nand U12687 (N_12687,N_12112,N_11607);
or U12688 (N_12688,N_12305,N_12451);
or U12689 (N_12689,N_12241,N_10085);
or U12690 (N_12690,N_11243,N_11364);
nor U12691 (N_12691,N_9844,N_10784);
or U12692 (N_12692,N_12192,N_12080);
nor U12693 (N_12693,N_10925,N_9696);
or U12694 (N_12694,N_9488,N_9661);
xnor U12695 (N_12695,N_10919,N_11101);
xnor U12696 (N_12696,N_10283,N_11598);
nor U12697 (N_12697,N_12006,N_11900);
nor U12698 (N_12698,N_11164,N_9727);
xnor U12699 (N_12699,N_11861,N_10754);
and U12700 (N_12700,N_10299,N_9956);
nor U12701 (N_12701,N_12021,N_12436);
nand U12702 (N_12702,N_12307,N_10739);
nand U12703 (N_12703,N_9617,N_9479);
xnor U12704 (N_12704,N_9676,N_11105);
nor U12705 (N_12705,N_12491,N_12486);
or U12706 (N_12706,N_11337,N_11613);
nor U12707 (N_12707,N_10100,N_11984);
and U12708 (N_12708,N_10166,N_11047);
nand U12709 (N_12709,N_9731,N_11452);
and U12710 (N_12710,N_11606,N_11921);
and U12711 (N_12711,N_9957,N_9985);
nand U12712 (N_12712,N_10742,N_11773);
or U12713 (N_12713,N_11332,N_9460);
and U12714 (N_12714,N_11148,N_12088);
nor U12715 (N_12715,N_10174,N_11571);
and U12716 (N_12716,N_10192,N_11662);
xnor U12717 (N_12717,N_11528,N_9413);
nor U12718 (N_12718,N_10535,N_10388);
and U12719 (N_12719,N_12034,N_9450);
nor U12720 (N_12720,N_9533,N_9571);
or U12721 (N_12721,N_11492,N_10442);
nor U12722 (N_12722,N_10608,N_9855);
nor U12723 (N_12723,N_11348,N_9660);
nand U12724 (N_12724,N_10990,N_9859);
nor U12725 (N_12725,N_10047,N_11999);
nand U12726 (N_12726,N_11808,N_11156);
nand U12727 (N_12727,N_11431,N_12439);
and U12728 (N_12728,N_11158,N_12433);
and U12729 (N_12729,N_9896,N_10466);
nor U12730 (N_12730,N_11311,N_9691);
or U12731 (N_12731,N_11525,N_10684);
nand U12732 (N_12732,N_10233,N_10530);
and U12733 (N_12733,N_10958,N_11734);
nor U12734 (N_12734,N_11782,N_11869);
nand U12735 (N_12735,N_12271,N_9548);
nand U12736 (N_12736,N_10076,N_11422);
xor U12737 (N_12737,N_10412,N_12346);
nor U12738 (N_12738,N_11686,N_11487);
xnor U12739 (N_12739,N_9930,N_12465);
nor U12740 (N_12740,N_11279,N_11413);
and U12741 (N_12741,N_12452,N_10257);
and U12742 (N_12742,N_11654,N_11997);
or U12743 (N_12743,N_10991,N_11780);
xnor U12744 (N_12744,N_9907,N_12207);
or U12745 (N_12745,N_9563,N_9651);
or U12746 (N_12746,N_11104,N_9962);
and U12747 (N_12747,N_9565,N_12211);
nor U12748 (N_12748,N_10194,N_10703);
and U12749 (N_12749,N_11108,N_10215);
nor U12750 (N_12750,N_11210,N_12431);
or U12751 (N_12751,N_9808,N_9906);
nand U12752 (N_12752,N_10789,N_10181);
nor U12753 (N_12753,N_10493,N_9522);
and U12754 (N_12754,N_10422,N_10575);
nor U12755 (N_12755,N_10416,N_12285);
nand U12756 (N_12756,N_11012,N_11820);
nand U12757 (N_12757,N_11610,N_9521);
or U12758 (N_12758,N_10867,N_12409);
nand U12759 (N_12759,N_9917,N_12203);
nor U12760 (N_12760,N_10509,N_9375);
nand U12761 (N_12761,N_11116,N_12058);
nand U12762 (N_12762,N_12267,N_11853);
or U12763 (N_12763,N_9472,N_9750);
or U12764 (N_12764,N_10912,N_9510);
nor U12765 (N_12765,N_10214,N_11240);
nand U12766 (N_12766,N_9715,N_10201);
nor U12767 (N_12767,N_11173,N_10956);
nand U12768 (N_12768,N_11787,N_11957);
nand U12769 (N_12769,N_11926,N_9941);
nand U12770 (N_12770,N_10725,N_11314);
or U12771 (N_12771,N_10942,N_11186);
nand U12772 (N_12772,N_9595,N_11258);
or U12773 (N_12773,N_11724,N_10714);
nor U12774 (N_12774,N_9402,N_11261);
or U12775 (N_12775,N_11825,N_10564);
nor U12776 (N_12776,N_12293,N_11549);
xor U12777 (N_12777,N_10286,N_9536);
xnor U12778 (N_12778,N_12490,N_12247);
or U12779 (N_12779,N_9455,N_12189);
or U12780 (N_12780,N_9952,N_9901);
nand U12781 (N_12781,N_11361,N_11511);
or U12782 (N_12782,N_9806,N_10109);
nand U12783 (N_12783,N_9714,N_11205);
and U12784 (N_12784,N_10385,N_9379);
and U12785 (N_12785,N_11766,N_11665);
or U12786 (N_12786,N_12485,N_10881);
nand U12787 (N_12787,N_12223,N_9701);
and U12788 (N_12788,N_10108,N_12375);
xor U12789 (N_12789,N_12322,N_11679);
or U12790 (N_12790,N_10870,N_10899);
and U12791 (N_12791,N_10918,N_11664);
nand U12792 (N_12792,N_10229,N_9596);
or U12793 (N_12793,N_12482,N_10278);
and U12794 (N_12794,N_9780,N_11838);
nor U12795 (N_12795,N_11849,N_10526);
nand U12796 (N_12796,N_10787,N_11038);
nand U12797 (N_12797,N_12417,N_11268);
nor U12798 (N_12798,N_10755,N_11069);
or U12799 (N_12799,N_11895,N_10399);
nand U12800 (N_12800,N_10665,N_10549);
and U12801 (N_12801,N_10048,N_12416);
and U12802 (N_12802,N_9777,N_11119);
and U12803 (N_12803,N_11989,N_11591);
and U12804 (N_12804,N_9585,N_10088);
or U12805 (N_12805,N_10809,N_12092);
or U12806 (N_12806,N_12413,N_11834);
and U12807 (N_12807,N_12478,N_11877);
and U12808 (N_12808,N_10694,N_12199);
nand U12809 (N_12809,N_9854,N_12428);
nor U12810 (N_12810,N_11818,N_11968);
nor U12811 (N_12811,N_9410,N_10871);
nor U12812 (N_12812,N_10492,N_11199);
or U12813 (N_12813,N_11098,N_10000);
nor U12814 (N_12814,N_10352,N_11809);
nor U12815 (N_12815,N_11073,N_11485);
or U12816 (N_12816,N_12370,N_9862);
xnor U12817 (N_12817,N_11188,N_12143);
xor U12818 (N_12818,N_12480,N_10126);
and U12819 (N_12819,N_9430,N_11676);
nor U12820 (N_12820,N_10837,N_10129);
and U12821 (N_12821,N_11439,N_10796);
or U12822 (N_12822,N_11244,N_11885);
or U12823 (N_12823,N_12472,N_11030);
nor U12824 (N_12824,N_10092,N_12349);
and U12825 (N_12825,N_12479,N_11715);
or U12826 (N_12826,N_12330,N_12408);
nor U12827 (N_12827,N_10972,N_10604);
nand U12828 (N_12828,N_11143,N_10136);
xnor U12829 (N_12829,N_10256,N_11546);
and U12830 (N_12830,N_12075,N_11278);
or U12831 (N_12831,N_9975,N_11732);
or U12832 (N_12832,N_10637,N_10200);
and U12833 (N_12833,N_10173,N_12244);
or U12834 (N_12834,N_12171,N_12221);
nand U12835 (N_12835,N_11757,N_11772);
nor U12836 (N_12836,N_10654,N_9628);
nand U12837 (N_12837,N_11407,N_11468);
and U12838 (N_12838,N_10987,N_11753);
nand U12839 (N_12839,N_11875,N_10380);
and U12840 (N_12840,N_11959,N_12137);
and U12841 (N_12841,N_11323,N_9749);
and U12842 (N_12842,N_11863,N_10435);
or U12843 (N_12843,N_10133,N_10961);
nor U12844 (N_12844,N_12105,N_11840);
or U12845 (N_12845,N_10993,N_10903);
nor U12846 (N_12846,N_11527,N_11378);
nor U12847 (N_12847,N_10379,N_11462);
or U12848 (N_12848,N_11467,N_10308);
and U12849 (N_12849,N_9490,N_12033);
or U12850 (N_12850,N_11085,N_11778);
and U12851 (N_12851,N_11687,N_11027);
xor U12852 (N_12852,N_11649,N_9894);
and U12853 (N_12853,N_12052,N_10355);
nand U12854 (N_12854,N_10261,N_10311);
and U12855 (N_12855,N_10029,N_10464);
and U12856 (N_12856,N_9448,N_12222);
nor U12857 (N_12857,N_10550,N_11319);
nand U12858 (N_12858,N_11333,N_11577);
xnor U12859 (N_12859,N_9439,N_9682);
or U12860 (N_12860,N_12186,N_9900);
nor U12861 (N_12861,N_10405,N_11932);
nor U12862 (N_12862,N_11138,N_9604);
and U12863 (N_12863,N_11429,N_11672);
nor U12864 (N_12864,N_11940,N_11582);
nand U12865 (N_12865,N_10552,N_12239);
nor U12866 (N_12866,N_12371,N_9625);
nor U12867 (N_12867,N_12444,N_11635);
or U12868 (N_12868,N_11035,N_10297);
or U12869 (N_12869,N_9721,N_10720);
and U12870 (N_12870,N_11510,N_12454);
nor U12871 (N_12871,N_11434,N_9852);
nor U12872 (N_12872,N_9505,N_11909);
and U12873 (N_12873,N_11678,N_12008);
nand U12874 (N_12874,N_11476,N_9785);
nor U12875 (N_12875,N_9553,N_11259);
or U12876 (N_12876,N_9757,N_12038);
nand U12877 (N_12877,N_9826,N_12339);
xnor U12878 (N_12878,N_10266,N_11717);
or U12879 (N_12879,N_12393,N_11925);
and U12880 (N_12880,N_10916,N_12048);
and U12881 (N_12881,N_11340,N_11960);
nand U12882 (N_12882,N_10227,N_9499);
and U12883 (N_12883,N_11969,N_11006);
and U12884 (N_12884,N_12387,N_11081);
or U12885 (N_12885,N_9923,N_11100);
xnor U12886 (N_12886,N_9441,N_10853);
or U12887 (N_12887,N_9577,N_9526);
or U12888 (N_12888,N_11346,N_11539);
nor U12889 (N_12889,N_11558,N_10559);
or U12890 (N_12890,N_10884,N_12359);
nand U12891 (N_12891,N_10625,N_11303);
xnor U12892 (N_12892,N_12493,N_10838);
or U12893 (N_12893,N_10440,N_11541);
and U12894 (N_12894,N_12333,N_10259);
nor U12895 (N_12895,N_9802,N_10748);
or U12896 (N_12896,N_10272,N_9846);
nor U12897 (N_12897,N_10676,N_9824);
nand U12898 (N_12898,N_10882,N_10699);
nand U12899 (N_12899,N_11974,N_11176);
or U12900 (N_12900,N_11789,N_10820);
or U12901 (N_12901,N_12265,N_10999);
nand U12902 (N_12902,N_9991,N_11418);
or U12903 (N_12903,N_10504,N_11142);
and U12904 (N_12904,N_9671,N_11614);
nand U12905 (N_12905,N_9603,N_10824);
nand U12906 (N_12906,N_11704,N_12499);
or U12907 (N_12907,N_11656,N_9995);
and U12908 (N_12908,N_10773,N_11800);
or U12909 (N_12909,N_12065,N_9636);
nor U12910 (N_12910,N_10054,N_9744);
xnor U12911 (N_12911,N_10825,N_12429);
nor U12912 (N_12912,N_10342,N_10941);
nand U12913 (N_12913,N_11859,N_10427);
and U12914 (N_12914,N_11162,N_9730);
or U12915 (N_12915,N_11727,N_11339);
and U12916 (N_12916,N_12025,N_11001);
or U12917 (N_12917,N_11713,N_10378);
nor U12918 (N_12918,N_11190,N_12165);
nand U12919 (N_12919,N_9685,N_10322);
or U12920 (N_12920,N_11118,N_10397);
or U12921 (N_12921,N_11891,N_9530);
or U12922 (N_12922,N_10462,N_12320);
xnor U12923 (N_12923,N_10546,N_11479);
and U12924 (N_12924,N_11764,N_11646);
nor U12925 (N_12925,N_12338,N_9774);
nor U12926 (N_12926,N_9728,N_11544);
nand U12927 (N_12927,N_11844,N_10198);
nor U12928 (N_12928,N_12016,N_10348);
and U12929 (N_12929,N_9458,N_11829);
and U12930 (N_12930,N_10040,N_11172);
nor U12931 (N_12931,N_11553,N_11293);
and U12932 (N_12932,N_9554,N_11718);
xor U12933 (N_12933,N_11347,N_9732);
and U12934 (N_12934,N_12396,N_10455);
nand U12935 (N_12935,N_12389,N_10722);
nand U12936 (N_12936,N_11308,N_10697);
nand U12937 (N_12937,N_11681,N_10507);
and U12938 (N_12938,N_11365,N_10591);
xor U12939 (N_12939,N_12078,N_11873);
or U12940 (N_12940,N_11583,N_9543);
or U12941 (N_12941,N_11636,N_11532);
nor U12942 (N_12942,N_10565,N_12455);
nor U12943 (N_12943,N_11230,N_9958);
nor U12944 (N_12944,N_11399,N_11153);
or U12945 (N_12945,N_11559,N_11473);
or U12946 (N_12946,N_11113,N_11436);
or U12947 (N_12947,N_10368,N_11435);
nand U12948 (N_12948,N_9809,N_10038);
nor U12949 (N_12949,N_10569,N_9961);
and U12950 (N_12950,N_9805,N_9787);
xor U12951 (N_12951,N_10976,N_10120);
nand U12952 (N_12952,N_9582,N_10863);
and U12953 (N_12953,N_10753,N_11107);
xor U12954 (N_12954,N_10202,N_12144);
and U12955 (N_12955,N_10056,N_9590);
and U12956 (N_12956,N_9540,N_10511);
or U12957 (N_12957,N_10801,N_9944);
or U12958 (N_12958,N_11482,N_11257);
and U12959 (N_12959,N_12212,N_12400);
and U12960 (N_12960,N_9949,N_11964);
nor U12961 (N_12961,N_12394,N_12353);
nor U12962 (N_12962,N_10293,N_9946);
nor U12963 (N_12963,N_11109,N_9570);
nor U12964 (N_12964,N_11222,N_10289);
nand U12965 (N_12965,N_10620,N_12024);
nand U12966 (N_12966,N_9766,N_12402);
nor U12967 (N_12967,N_11821,N_10169);
nand U12968 (N_12968,N_10083,N_11140);
or U12969 (N_12969,N_11842,N_10414);
nor U12970 (N_12970,N_9643,N_12040);
nor U12971 (N_12971,N_9994,N_11774);
xnor U12972 (N_12972,N_11032,N_11651);
nand U12973 (N_12973,N_10006,N_10850);
nand U12974 (N_12974,N_11031,N_10913);
nor U12975 (N_12975,N_12348,N_9951);
nor U12976 (N_12976,N_12146,N_10533);
nand U12977 (N_12977,N_11182,N_11421);
or U12978 (N_12978,N_11320,N_11045);
or U12979 (N_12979,N_9429,N_10418);
or U12980 (N_12980,N_10617,N_10062);
or U12981 (N_12981,N_10354,N_11264);
nand U12982 (N_12982,N_9870,N_11088);
and U12983 (N_12983,N_11131,N_9657);
nor U12984 (N_12984,N_10985,N_12198);
nand U12985 (N_12985,N_10685,N_12185);
nor U12986 (N_12986,N_10716,N_10346);
or U12987 (N_12987,N_11034,N_10264);
nor U12988 (N_12988,N_10178,N_12138);
and U12989 (N_12989,N_9927,N_11345);
or U12990 (N_12990,N_9629,N_11154);
nand U12991 (N_12991,N_11852,N_12259);
nor U12992 (N_12992,N_11215,N_11204);
nand U12993 (N_12993,N_10485,N_11171);
or U12994 (N_12994,N_9964,N_10184);
and U12995 (N_12995,N_11694,N_10247);
nand U12996 (N_12996,N_9861,N_12358);
nand U12997 (N_12997,N_9414,N_11097);
nand U12998 (N_12998,N_12066,N_9789);
or U12999 (N_12999,N_11342,N_9404);
or U13000 (N_13000,N_12201,N_10548);
xor U13001 (N_13001,N_12424,N_11248);
nand U13002 (N_13002,N_9392,N_10932);
and U13003 (N_13003,N_11192,N_11315);
and U13004 (N_13004,N_12498,N_10760);
and U13005 (N_13005,N_10708,N_9788);
nand U13006 (N_13006,N_9972,N_12030);
nand U13007 (N_13007,N_11071,N_10204);
nand U13008 (N_13008,N_12464,N_10618);
nor U13009 (N_13009,N_11384,N_10908);
nand U13010 (N_13010,N_11692,N_11742);
nand U13011 (N_13011,N_11621,N_11516);
and U13012 (N_13012,N_9653,N_11576);
or U13013 (N_13013,N_10471,N_11572);
or U13014 (N_13014,N_11669,N_11622);
or U13015 (N_13015,N_11836,N_10562);
nor U13016 (N_13016,N_9737,N_11198);
and U13017 (N_13017,N_9386,N_11826);
xnor U13018 (N_13018,N_10336,N_9982);
nor U13019 (N_13019,N_10592,N_9547);
nand U13020 (N_13020,N_11189,N_10052);
or U13021 (N_13021,N_11432,N_11507);
nor U13022 (N_13022,N_11867,N_11586);
nor U13023 (N_13023,N_10439,N_10067);
and U13024 (N_13024,N_10519,N_10605);
and U13025 (N_13025,N_9612,N_11615);
and U13026 (N_13026,N_12073,N_9960);
nand U13027 (N_13027,N_10419,N_10292);
or U13028 (N_13028,N_10079,N_10024);
or U13029 (N_13029,N_9501,N_10980);
xnor U13030 (N_13030,N_10145,N_10968);
xor U13031 (N_13031,N_10288,N_9719);
and U13032 (N_13032,N_10588,N_10058);
xnor U13033 (N_13033,N_10931,N_9976);
nor U13034 (N_13034,N_9594,N_11351);
or U13035 (N_13035,N_10122,N_10503);
or U13036 (N_13036,N_12176,N_10828);
nand U13037 (N_13037,N_11207,N_11941);
or U13038 (N_13038,N_11180,N_11286);
nand U13039 (N_13039,N_12213,N_9989);
or U13040 (N_13040,N_12169,N_11458);
nand U13041 (N_13041,N_11980,N_11139);
nor U13042 (N_13042,N_10640,N_11634);
and U13043 (N_13043,N_12083,N_10539);
or U13044 (N_13044,N_10603,N_11194);
xor U13045 (N_13045,N_12418,N_10643);
and U13046 (N_13046,N_11906,N_12456);
and U13047 (N_13047,N_12286,N_11526);
nor U13048 (N_13048,N_11747,N_10606);
or U13049 (N_13049,N_11866,N_12274);
nand U13050 (N_13050,N_9921,N_12106);
and U13051 (N_13051,N_11209,N_12395);
and U13052 (N_13052,N_10657,N_11359);
and U13053 (N_13053,N_10468,N_9819);
nand U13054 (N_13054,N_12249,N_11443);
nand U13055 (N_13055,N_10572,N_10082);
nor U13056 (N_13056,N_12093,N_10350);
xor U13057 (N_13057,N_12430,N_9613);
or U13058 (N_13058,N_11372,N_11958);
nor U13059 (N_13059,N_11160,N_9395);
or U13060 (N_13060,N_9856,N_11022);
or U13061 (N_13061,N_10306,N_11093);
nand U13062 (N_13062,N_12295,N_10876);
nand U13063 (N_13063,N_10790,N_9672);
and U13064 (N_13064,N_9799,N_10025);
and U13065 (N_13065,N_10104,N_11868);
nand U13066 (N_13066,N_11318,N_10315);
or U13067 (N_13067,N_11277,N_11699);
nand U13068 (N_13068,N_9918,N_9525);
nor U13069 (N_13069,N_11059,N_11401);
nor U13070 (N_13070,N_10452,N_10759);
nor U13071 (N_13071,N_11409,N_12129);
and U13072 (N_13072,N_12419,N_10923);
and U13073 (N_13073,N_9825,N_11122);
and U13074 (N_13074,N_10965,N_12027);
or U13075 (N_13075,N_11573,N_10365);
nor U13076 (N_13076,N_11981,N_10246);
nand U13077 (N_13077,N_9836,N_10946);
and U13078 (N_13078,N_10347,N_9493);
and U13079 (N_13079,N_9425,N_9632);
nor U13080 (N_13080,N_12076,N_9675);
nor U13081 (N_13081,N_11304,N_10335);
and U13082 (N_13082,N_10180,N_10847);
and U13083 (N_13083,N_11886,N_11099);
and U13084 (N_13084,N_12388,N_10695);
nand U13085 (N_13085,N_12410,N_12045);
or U13086 (N_13086,N_9610,N_11103);
nor U13087 (N_13087,N_11313,N_12364);
xor U13088 (N_13088,N_12231,N_11226);
nand U13089 (N_13089,N_11086,N_10602);
nor U13090 (N_13090,N_11334,N_10826);
and U13091 (N_13091,N_10282,N_10710);
and U13092 (N_13092,N_9935,N_12191);
or U13093 (N_13093,N_10651,N_12283);
or U13094 (N_13094,N_10393,N_11367);
and U13095 (N_13095,N_9467,N_12069);
xnor U13096 (N_13096,N_10171,N_10599);
nor U13097 (N_13097,N_11798,N_11201);
nand U13098 (N_13098,N_10382,N_11915);
nor U13099 (N_13099,N_11393,N_9909);
or U13100 (N_13100,N_10213,N_10571);
and U13101 (N_13101,N_11329,N_11196);
or U13102 (N_13102,N_9745,N_9939);
xor U13103 (N_13103,N_11440,N_11289);
and U13104 (N_13104,N_10619,N_10767);
nor U13105 (N_13105,N_11641,N_11275);
nand U13106 (N_13106,N_11994,N_10843);
nor U13107 (N_13107,N_10118,N_10099);
nor U13108 (N_13108,N_12111,N_11498);
or U13109 (N_13109,N_9833,N_12071);
or U13110 (N_13110,N_10713,N_11503);
or U13111 (N_13111,N_10893,N_11538);
xnor U13112 (N_13112,N_11331,N_10363);
nor U13113 (N_13113,N_10611,N_12296);
xnor U13114 (N_13114,N_12004,N_11177);
nand U13115 (N_13115,N_11720,N_10205);
xor U13116 (N_13116,N_10071,N_10170);
nand U13117 (N_13117,N_10478,N_12054);
xor U13118 (N_13118,N_11786,N_9725);
nor U13119 (N_13119,N_11874,N_11865);
nor U13120 (N_13120,N_11390,N_11260);
nor U13121 (N_13121,N_11657,N_11231);
nor U13122 (N_13122,N_9588,N_10159);
or U13123 (N_13123,N_10780,N_12278);
and U13124 (N_13124,N_9937,N_9517);
nor U13125 (N_13125,N_11883,N_10013);
and U13126 (N_13126,N_10224,N_9965);
nand U13127 (N_13127,N_9765,N_10413);
nor U13128 (N_13128,N_10473,N_12210);
nand U13129 (N_13129,N_10428,N_11495);
and U13130 (N_13130,N_12209,N_9415);
nor U13131 (N_13131,N_9557,N_11806);
nand U13132 (N_13132,N_10541,N_10007);
and U13133 (N_13133,N_11123,N_10917);
nand U13134 (N_13134,N_11761,N_12329);
and U13135 (N_13135,N_11112,N_11578);
or U13136 (N_13136,N_10329,N_11682);
nand U13137 (N_13137,N_12350,N_12179);
xnor U13138 (N_13138,N_11265,N_10974);
and U13139 (N_13139,N_10892,N_10560);
nor U13140 (N_13140,N_10817,N_11524);
nand U13141 (N_13141,N_11151,N_10177);
nor U13142 (N_13142,N_11791,N_11178);
and U13143 (N_13143,N_9697,N_9680);
nand U13144 (N_13144,N_12385,N_11850);
xor U13145 (N_13145,N_12074,N_10349);
nand U13146 (N_13146,N_10115,N_11563);
or U13147 (N_13147,N_10151,N_11280);
nand U13148 (N_13148,N_10041,N_11644);
xnor U13149 (N_13149,N_11461,N_9782);
or U13150 (N_13150,N_11851,N_10004);
nor U13151 (N_13151,N_10582,N_9998);
and U13152 (N_13152,N_12306,N_12365);
and U13153 (N_13153,N_10472,N_10070);
nand U13154 (N_13154,N_10840,N_12170);
nor U13155 (N_13155,N_9427,N_10642);
nor U13156 (N_13156,N_9516,N_11907);
nand U13157 (N_13157,N_10274,N_10690);
nand U13158 (N_13158,N_9442,N_11552);
or U13159 (N_13159,N_11366,N_10489);
xor U13160 (N_13160,N_9669,N_11627);
or U13161 (N_13161,N_10858,N_9838);
or U13162 (N_13162,N_11936,N_10121);
nor U13163 (N_13163,N_10127,N_11125);
nand U13164 (N_13164,N_11056,N_10532);
nand U13165 (N_13165,N_9767,N_11903);
and U13166 (N_13166,N_11161,N_12003);
nand U13167 (N_13167,N_11775,N_11428);
or U13168 (N_13168,N_9464,N_11946);
or U13169 (N_13169,N_11219,N_10447);
xor U13170 (N_13170,N_10316,N_10766);
and U13171 (N_13171,N_10717,N_10423);
and U13172 (N_13172,N_11934,N_11616);
nand U13173 (N_13173,N_11542,N_10922);
and U13174 (N_13174,N_12376,N_11792);
nor U13175 (N_13175,N_12378,N_11206);
nor U13176 (N_13176,N_11292,N_10207);
nor U13177 (N_13177,N_10183,N_10167);
nor U13178 (N_13178,N_10833,N_10505);
nand U13179 (N_13179,N_9485,N_11274);
nor U13180 (N_13180,N_12164,N_12383);
nand U13181 (N_13181,N_10459,N_12070);
xor U13182 (N_13182,N_10097,N_11952);
or U13183 (N_13183,N_9823,N_11893);
or U13184 (N_13184,N_10199,N_12236);
or U13185 (N_13185,N_9800,N_10528);
or U13186 (N_13186,N_10891,N_10255);
nor U13187 (N_13187,N_9851,N_10377);
or U13188 (N_13188,N_10704,N_12477);
nor U13189 (N_13189,N_9864,N_9779);
nor U13190 (N_13190,N_10268,N_12448);
xor U13191 (N_13191,N_9974,N_10888);
nor U13192 (N_13192,N_11677,N_11927);
nand U13193 (N_13193,N_9845,N_11242);
nand U13194 (N_13194,N_12290,N_11387);
nand U13195 (N_13195,N_9445,N_11793);
xnor U13196 (N_13196,N_11731,N_10911);
nor U13197 (N_13197,N_11414,N_10827);
xnor U13198 (N_13198,N_11993,N_11144);
or U13199 (N_13199,N_10894,N_12366);
nand U13200 (N_13200,N_10883,N_10624);
or U13201 (N_13201,N_10981,N_10573);
nor U13202 (N_13202,N_10621,N_9848);
or U13203 (N_13203,N_9630,N_11225);
xnor U13204 (N_13204,N_10906,N_11328);
nand U13205 (N_13205,N_9740,N_10967);
nand U13206 (N_13206,N_10186,N_10295);
and U13207 (N_13207,N_11464,N_9646);
and U13208 (N_13208,N_11380,N_11995);
xnor U13209 (N_13209,N_11523,N_10686);
and U13210 (N_13210,N_10737,N_10161);
nor U13211 (N_13211,N_10310,N_10467);
xor U13212 (N_13212,N_10463,N_9555);
or U13213 (N_13213,N_10073,N_10334);
xnor U13214 (N_13214,N_10469,N_12049);
nor U13215 (N_13215,N_11856,N_11475);
or U13216 (N_13216,N_10601,N_10324);
xor U13217 (N_13217,N_11847,N_9622);
nor U13218 (N_13218,N_10208,N_10683);
nand U13219 (N_13219,N_12059,N_11534);
and U13220 (N_13220,N_9662,N_10875);
nor U13221 (N_13221,N_11281,N_9496);
and U13222 (N_13222,N_10043,N_12238);
nor U13223 (N_13223,N_9418,N_10210);
nor U13224 (N_13224,N_11771,N_11354);
nor U13225 (N_13225,N_10203,N_11882);
nor U13226 (N_13226,N_11763,N_11276);
or U13227 (N_13227,N_10898,N_11737);
nor U13228 (N_13228,N_12135,N_9549);
and U13229 (N_13229,N_11996,N_11305);
nor U13230 (N_13230,N_11167,N_12381);
or U13231 (N_13231,N_12294,N_9623);
and U13232 (N_13232,N_12426,N_10889);
nor U13233 (N_13233,N_9877,N_11560);
or U13234 (N_13234,N_12404,N_10248);
or U13235 (N_13235,N_11536,N_10068);
nand U13236 (N_13236,N_10451,N_12347);
nand U13237 (N_13237,N_11637,N_10234);
and U13238 (N_13238,N_12085,N_10182);
xnor U13239 (N_13239,N_10805,N_11827);
or U13240 (N_13240,N_10689,N_10982);
nand U13241 (N_13241,N_10641,N_11755);
and U13242 (N_13242,N_10140,N_12446);
xnor U13243 (N_13243,N_10800,N_11777);
nor U13244 (N_13244,N_10566,N_10670);
and U13245 (N_13245,N_9560,N_10834);
nor U13246 (N_13246,N_9812,N_10077);
and U13247 (N_13247,N_9748,N_11247);
or U13248 (N_13248,N_11076,N_9659);
and U13249 (N_13249,N_9624,N_9478);
xnor U13250 (N_13250,N_9945,N_11547);
nand U13251 (N_13251,N_11072,N_10527);
nor U13252 (N_13252,N_10995,N_11725);
nand U13253 (N_13253,N_11919,N_9913);
xor U13254 (N_13254,N_10275,N_12352);
or U13255 (N_13255,N_12463,N_10226);
nand U13256 (N_13256,N_10583,N_10577);
nand U13257 (N_13257,N_11405,N_9544);
or U13258 (N_13258,N_10746,N_9599);
or U13259 (N_13259,N_9551,N_10992);
nand U13260 (N_13260,N_10520,N_12360);
nor U13261 (N_13261,N_12022,N_11494);
nand U13262 (N_13262,N_12081,N_9933);
xor U13263 (N_13263,N_11080,N_9494);
nand U13264 (N_13264,N_11499,N_12067);
nor U13265 (N_13265,N_12266,N_11594);
nor U13266 (N_13266,N_12460,N_10402);
nor U13267 (N_13267,N_11216,N_11671);
and U13268 (N_13268,N_12114,N_12403);
and U13269 (N_13269,N_12437,N_12327);
nor U13270 (N_13270,N_11472,N_9886);
nand U13271 (N_13271,N_10001,N_10975);
xnor U13272 (N_13272,N_11299,N_10540);
and U13273 (N_13273,N_11629,N_9598);
nand U13274 (N_13274,N_9763,N_11325);
nor U13275 (N_13275,N_10947,N_11392);
and U13276 (N_13276,N_10445,N_10842);
nor U13277 (N_13277,N_10373,N_11695);
nand U13278 (N_13278,N_11381,N_10680);
xor U13279 (N_13279,N_10287,N_10113);
and U13280 (N_13280,N_11183,N_9384);
and U13281 (N_13281,N_11191,N_9634);
nor U13282 (N_13282,N_11457,N_11223);
and U13283 (N_13283,N_9482,N_11540);
or U13284 (N_13284,N_10080,N_10341);
and U13285 (N_13285,N_10845,N_10794);
nand U13286 (N_13286,N_10696,N_11590);
or U13287 (N_13287,N_12438,N_10175);
or U13288 (N_13288,N_11067,N_10456);
nor U13289 (N_13289,N_9882,N_10337);
and U13290 (N_13290,N_9735,N_9486);
and U13291 (N_13291,N_11765,N_10132);
or U13292 (N_13292,N_10578,N_11739);
or U13293 (N_13293,N_9678,N_11872);
nand U13294 (N_13294,N_10969,N_11543);
xnor U13295 (N_13295,N_9614,N_9580);
nand U13296 (N_13296,N_12050,N_10146);
nor U13297 (N_13297,N_10242,N_10262);
and U13298 (N_13298,N_10749,N_10626);
and U13299 (N_13299,N_11795,N_12281);
or U13300 (N_13300,N_9411,N_9506);
nor U13301 (N_13301,N_10727,N_11253);
nor U13302 (N_13302,N_11815,N_12095);
nand U13303 (N_13303,N_9729,N_12284);
nor U13304 (N_13304,N_9666,N_10406);
nor U13305 (N_13305,N_11812,N_10750);
nand U13306 (N_13306,N_9983,N_9872);
nor U13307 (N_13307,N_12242,N_10267);
and U13308 (N_13308,N_11403,N_9959);
nand U13309 (N_13309,N_11520,N_9383);
nand U13310 (N_13310,N_11684,N_10250);
nor U13311 (N_13311,N_10940,N_12392);
xnor U13312 (N_13312,N_9431,N_10172);
or U13313 (N_13313,N_10538,N_10764);
and U13314 (N_13314,N_11744,N_10050);
nor U13315 (N_13315,N_11617,N_10644);
xor U13316 (N_13316,N_9524,N_10330);
or U13317 (N_13317,N_10486,N_12270);
nand U13318 (N_13318,N_9798,N_11051);
nand U13319 (N_13319,N_9843,N_12310);
nor U13320 (N_13320,N_9904,N_12257);
or U13321 (N_13321,N_11814,N_12041);
or U13322 (N_13322,N_10581,N_9489);
nor U13323 (N_13323,N_10747,N_11894);
and U13324 (N_13324,N_10830,N_12466);
and U13325 (N_13325,N_9664,N_11141);
nor U13326 (N_13326,N_10057,N_10944);
xor U13327 (N_13327,N_10074,N_9857);
and U13328 (N_13328,N_10551,N_11417);
or U13329 (N_13329,N_12272,N_12357);
nand U13330 (N_13330,N_9576,N_9761);
or U13331 (N_13331,N_11648,N_11531);
nand U13332 (N_13332,N_12434,N_12229);
nor U13333 (N_13333,N_11114,N_10886);
nor U13334 (N_13334,N_11135,N_9573);
and U13335 (N_13335,N_11521,N_12109);
or U13336 (N_13336,N_10150,N_11683);
nand U13337 (N_13337,N_9655,N_12497);
and U13338 (N_13338,N_10383,N_11864);
or U13339 (N_13339,N_11855,N_9929);
xor U13340 (N_13340,N_10815,N_10952);
and U13341 (N_13341,N_10615,N_11057);
nor U13342 (N_13342,N_12449,N_9471);
nor U13343 (N_13343,N_11881,N_12167);
or U13344 (N_13344,N_11858,N_10928);
or U13345 (N_13345,N_11716,N_10441);
or U13346 (N_13346,N_10909,N_9895);
nor U13347 (N_13347,N_11324,N_10488);
nor U13348 (N_13348,N_10933,N_11444);
nor U13349 (N_13349,N_10998,N_10966);
xor U13350 (N_13350,N_12156,N_11070);
and U13351 (N_13351,N_10996,N_11062);
and U13352 (N_13352,N_11290,N_9811);
nand U13353 (N_13353,N_10741,N_11609);
or U13354 (N_13354,N_11899,N_10769);
and U13355 (N_13355,N_9475,N_9564);
xnor U13356 (N_13356,N_10069,N_11688);
or U13357 (N_13357,N_10854,N_12130);
xnor U13358 (N_13358,N_11658,N_11632);
nand U13359 (N_13359,N_9734,N_9686);
and U13360 (N_13360,N_11832,N_9898);
nor U13361 (N_13361,N_10555,N_10970);
or U13362 (N_13362,N_10189,N_10682);
and U13363 (N_13363,N_11685,N_10792);
or U13364 (N_13364,N_11710,N_9733);
or U13365 (N_13365,N_9770,N_9642);
xor U13366 (N_13366,N_10016,N_9641);
xnor U13367 (N_13367,N_12288,N_11967);
nor U13368 (N_13368,N_10639,N_11224);
nor U13369 (N_13369,N_12090,N_11252);
and U13370 (N_13370,N_11133,N_11533);
xor U13371 (N_13371,N_11271,N_11579);
nor U13372 (N_13372,N_10103,N_10649);
nand U13373 (N_13373,N_11589,N_10343);
and U13374 (N_13374,N_11326,N_12002);
or U13375 (N_13375,N_9772,N_10531);
or U13376 (N_13376,N_11519,N_12251);
nor U13377 (N_13377,N_10238,N_10672);
nor U13378 (N_13378,N_11673,N_12492);
or U13379 (N_13379,N_11962,N_12217);
or U13380 (N_13380,N_10738,N_11555);
nand U13381 (N_13381,N_11561,N_12369);
or U13382 (N_13382,N_10091,N_10179);
nor U13383 (N_13383,N_9700,N_10351);
nand U13384 (N_13384,N_11451,N_11420);
nor U13385 (N_13385,N_10711,N_9829);
and U13386 (N_13386,N_11630,N_9797);
and U13387 (N_13387,N_9541,N_10778);
or U13388 (N_13388,N_9796,N_9842);
xor U13389 (N_13389,N_11650,N_10758);
nand U13390 (N_13390,N_11711,N_11501);
nand U13391 (N_13391,N_9670,N_10369);
or U13392 (N_13392,N_11269,N_12445);
nand U13393 (N_13393,N_12235,N_12220);
nand U13394 (N_13394,N_9572,N_10009);
xor U13395 (N_13395,N_9654,N_10028);
or U13396 (N_13396,N_9890,N_12098);
nor U13397 (N_13397,N_12115,N_10137);
nor U13398 (N_13398,N_12313,N_12230);
or U13399 (N_13399,N_9401,N_11522);
xor U13400 (N_13400,N_9419,N_10735);
or U13401 (N_13401,N_11213,N_12405);
or U13402 (N_13402,N_12421,N_10793);
xor U13403 (N_13403,N_10761,N_10561);
nand U13404 (N_13404,N_10740,N_9552);
and U13405 (N_13405,N_11841,N_11854);
nand U13406 (N_13406,N_11642,N_10772);
or U13407 (N_13407,N_9583,N_10666);
nor U13408 (N_13408,N_11748,N_9784);
xnor U13409 (N_13409,N_9868,N_11127);
and U13410 (N_13410,N_12342,N_11567);
nor U13411 (N_13411,N_10724,N_12314);
nand U13412 (N_13412,N_11652,N_11990);
and U13413 (N_13413,N_10576,N_10691);
or U13414 (N_13414,N_10003,N_10407);
and U13415 (N_13415,N_11600,N_11804);
or U13416 (N_13416,N_11232,N_10149);
or U13417 (N_13417,N_10107,N_10265);
and U13418 (N_13418,N_9713,N_10622);
and U13419 (N_13419,N_10613,N_9707);
nor U13420 (N_13420,N_10701,N_11049);
xnor U13421 (N_13421,N_9791,N_10206);
nor U13422 (N_13422,N_11839,N_10623);
nor U13423 (N_13423,N_12277,N_12091);
xnor U13424 (N_13424,N_11170,N_12262);
or U13425 (N_13425,N_11965,N_9942);
xnor U13426 (N_13426,N_11048,N_12234);
and U13427 (N_13427,N_11556,N_10362);
nand U13428 (N_13428,N_10390,N_9710);
nand U13429 (N_13429,N_12089,N_11040);
and U13430 (N_13430,N_11824,N_11947);
nor U13431 (N_13431,N_10187,N_11410);
and U13432 (N_13432,N_11237,N_11890);
nor U13433 (N_13433,N_10119,N_12100);
nand U13434 (N_13434,N_10638,N_11833);
or U13435 (N_13435,N_9454,N_11696);
nor U13436 (N_13436,N_9986,N_10160);
xnor U13437 (N_13437,N_9919,N_12441);
or U13438 (N_13438,N_11730,N_10328);
xnor U13439 (N_13439,N_11797,N_9703);
and U13440 (N_13440,N_9483,N_10046);
and U13441 (N_13441,N_11799,N_10188);
xnor U13442 (N_13442,N_10986,N_9940);
nand U13443 (N_13443,N_11134,N_10658);
and U13444 (N_13444,N_10579,N_10937);
and U13445 (N_13445,N_12246,N_9754);
or U13446 (N_13446,N_12337,N_10979);
and U13447 (N_13447,N_9936,N_9821);
nor U13448 (N_13448,N_9769,N_11666);
nor U13449 (N_13449,N_12255,N_9391);
nor U13450 (N_13450,N_11233,N_10296);
or U13451 (N_13451,N_11245,N_10936);
nor U13452 (N_13452,N_10791,N_11709);
nor U13453 (N_13453,N_11491,N_11480);
nor U13454 (N_13454,N_10983,N_9627);
and U13455 (N_13455,N_11425,N_12010);
nor U13456 (N_13456,N_11061,N_10358);
nor U13457 (N_13457,N_10277,N_11992);
and U13458 (N_13458,N_10915,N_12043);
xnor U13459 (N_13459,N_11668,N_11017);
or U13460 (N_13460,N_10831,N_9781);
or U13461 (N_13461,N_9484,N_12149);
or U13462 (N_13462,N_10963,N_11015);
nor U13463 (N_13463,N_11745,N_10660);
and U13464 (N_13464,N_11535,N_10195);
nand U13465 (N_13465,N_10669,N_9649);
and U13466 (N_13466,N_9650,N_10632);
and U13467 (N_13467,N_10303,N_12258);
nand U13468 (N_13468,N_9871,N_10094);
nand U13469 (N_13469,N_11988,N_12009);
nand U13470 (N_13470,N_11009,N_11843);
and U13471 (N_13471,N_10692,N_9652);
nor U13472 (N_13472,N_11147,N_9878);
and U13473 (N_13473,N_11618,N_11385);
nor U13474 (N_13474,N_12471,N_10404);
nand U13475 (N_13475,N_10730,N_11184);
and U13476 (N_13476,N_10217,N_9567);
nand U13477 (N_13477,N_12190,N_10930);
nand U13478 (N_13478,N_10263,N_11876);
xnor U13479 (N_13479,N_9481,N_10294);
nand U13480 (N_13480,N_12136,N_10896);
or U13481 (N_13481,N_11010,N_11871);
or U13482 (N_13482,N_9463,N_12178);
or U13483 (N_13483,N_11604,N_12453);
nand U13484 (N_13484,N_10344,N_11408);
nor U13485 (N_13485,N_10138,N_11272);
or U13486 (N_13486,N_12260,N_12397);
nor U13487 (N_13487,N_11128,N_11735);
nor U13488 (N_13488,N_10244,N_11447);
nand U13489 (N_13489,N_9736,N_9726);
nor U13490 (N_13490,N_10857,N_11822);
or U13491 (N_13491,N_9916,N_12373);
nor U13492 (N_13492,N_10802,N_10364);
or U13493 (N_13493,N_9461,N_12276);
nor U13494 (N_13494,N_12023,N_10832);
nor U13495 (N_13495,N_11626,N_12118);
and U13496 (N_13496,N_12468,N_10338);
nor U13497 (N_13497,N_10935,N_11285);
nand U13498 (N_13498,N_11066,N_10066);
xor U13499 (N_13499,N_10656,N_10372);
nor U13500 (N_13500,N_11557,N_11202);
xnor U13501 (N_13501,N_11484,N_10734);
nand U13502 (N_13502,N_12125,N_9706);
nor U13503 (N_13503,N_10736,N_12291);
or U13504 (N_13504,N_9815,N_12324);
or U13505 (N_13505,N_10756,N_11939);
nor U13506 (N_13506,N_11221,N_11726);
or U13507 (N_13507,N_9611,N_11985);
nor U13508 (N_13508,N_10587,N_10495);
or U13509 (N_13509,N_12300,N_9518);
or U13510 (N_13510,N_11961,N_12141);
or U13511 (N_13511,N_10185,N_10144);
nand U13512 (N_13512,N_11004,N_12133);
and U13513 (N_13513,N_10659,N_11659);
and U13514 (N_13514,N_10134,N_10949);
nor U13515 (N_13515,N_10673,N_10596);
and U13516 (N_13516,N_10360,N_10681);
and U13517 (N_13517,N_10667,N_10339);
and U13518 (N_13518,N_9922,N_9938);
nand U13519 (N_13519,N_11355,N_9495);
and U13520 (N_13520,N_10011,N_11055);
or U13521 (N_13521,N_11014,N_9751);
nor U13522 (N_13522,N_9762,N_11155);
or U13523 (N_13523,N_11588,N_11397);
or U13524 (N_13524,N_9984,N_10026);
nor U13525 (N_13525,N_12362,N_10249);
and U13526 (N_13526,N_11945,N_10904);
nand U13527 (N_13527,N_11039,N_12435);
nand U13528 (N_13528,N_9953,N_11991);
and U13529 (N_13529,N_12056,N_11246);
and U13530 (N_13530,N_11811,N_9683);
nand U13531 (N_13531,N_10153,N_9990);
nand U13532 (N_13532,N_12355,N_12318);
xor U13533 (N_13533,N_9435,N_12097);
nor U13534 (N_13534,N_11640,N_9810);
nand U13535 (N_13535,N_11497,N_10494);
and U13536 (N_13536,N_11052,N_9593);
nand U13537 (N_13537,N_11363,N_12390);
nand U13538 (N_13538,N_11203,N_9579);
xor U13539 (N_13539,N_11455,N_9545);
and U13540 (N_13540,N_9889,N_10498);
and U13541 (N_13541,N_10319,N_10497);
nand U13542 (N_13542,N_11929,N_12226);
nor U13543 (N_13543,N_11611,N_9500);
nand U13544 (N_13544,N_11136,N_12218);
nand U13545 (N_13545,N_11914,N_10044);
or U13546 (N_13546,N_10039,N_11758);
xor U13547 (N_13547,N_9978,N_10317);
and U13548 (N_13548,N_11195,N_10154);
or U13549 (N_13549,N_12216,N_10022);
or U13550 (N_13550,N_11675,N_10481);
nand U13551 (N_13551,N_10994,N_11955);
or U13552 (N_13552,N_12012,N_11058);
or U13553 (N_13553,N_10508,N_9743);
nand U13554 (N_13554,N_9827,N_11918);
nand U13555 (N_13555,N_9993,N_11845);
xor U13556 (N_13556,N_10897,N_10585);
nor U13557 (N_13557,N_12384,N_11703);
or U13558 (N_13558,N_10984,N_12325);
nand U13559 (N_13559,N_9795,N_11502);
and U13560 (N_13560,N_11470,N_11802);
or U13561 (N_13561,N_12264,N_11063);
nand U13562 (N_13562,N_10785,N_11944);
nor U13563 (N_13563,N_12253,N_10305);
or U13564 (N_13564,N_10240,N_11508);
nand U13565 (N_13565,N_10465,N_9704);
nand U13566 (N_13566,N_11691,N_12195);
and U13567 (N_13567,N_9528,N_10290);
and U13568 (N_13568,N_11920,N_10285);
nand U13569 (N_13569,N_9389,N_10111);
nand U13570 (N_13570,N_10544,N_10647);
xnor U13571 (N_13571,N_11298,N_10719);
or U13572 (N_13572,N_10728,N_11801);
and U13573 (N_13573,N_10084,N_11396);
and U13574 (N_13574,N_11515,N_10116);
or U13575 (N_13575,N_10191,N_10536);
xor U13576 (N_13576,N_9584,N_9378);
nand U13577 (N_13577,N_12101,N_9813);
or U13578 (N_13578,N_11904,N_9915);
xor U13579 (N_13579,N_11663,N_12495);
nor U13580 (N_13580,N_9873,N_11043);
nand U13581 (N_13581,N_11053,N_11803);
nor U13582 (N_13582,N_10222,N_9684);
and U13583 (N_13583,N_10117,N_12351);
and U13584 (N_13584,N_11370,N_11580);
and U13585 (N_13585,N_11670,N_11846);
or U13586 (N_13586,N_11449,N_12483);
xor U13587 (N_13587,N_11386,N_12096);
or U13588 (N_13588,N_9667,N_9546);
nand U13589 (N_13589,N_11283,N_12458);
nor U13590 (N_13590,N_10059,N_10939);
and U13591 (N_13591,N_10323,N_11698);
nor U13592 (N_13592,N_9626,N_11639);
or U13593 (N_13593,N_11608,N_11817);
nand U13594 (N_13594,N_9702,N_10698);
or U13595 (N_13595,N_9790,N_10436);
nand U13596 (N_13596,N_12232,N_11450);
or U13597 (N_13597,N_12103,N_9716);
and U13598 (N_13598,N_10848,N_10563);
xor U13599 (N_13599,N_11336,N_10627);
nand U13600 (N_13600,N_11023,N_11044);
nor U13601 (N_13601,N_11357,N_12237);
nor U13602 (N_13602,N_9561,N_10168);
nor U13603 (N_13603,N_10661,N_11998);
or U13604 (N_13604,N_10367,N_10938);
nor U13605 (N_13605,N_10143,N_10302);
and U13606 (N_13606,N_12140,N_10482);
or U13607 (N_13607,N_12086,N_12273);
or U13608 (N_13608,N_10821,N_10312);
nor U13609 (N_13609,N_12345,N_9814);
nand U13610 (N_13610,N_10037,N_9519);
and U13611 (N_13611,N_10693,N_12379);
nor U13612 (N_13612,N_10460,N_9925);
and U13613 (N_13613,N_12432,N_9459);
nor U13614 (N_13614,N_11719,N_10353);
nor U13615 (N_13615,N_10446,N_12319);
nand U13616 (N_13616,N_9508,N_12399);
xor U13617 (N_13617,N_10806,N_12184);
nand U13618 (N_13618,N_11647,N_11779);
nand U13619 (N_13619,N_10496,N_9681);
nand U13620 (N_13620,N_11830,N_10156);
nor U13621 (N_13621,N_12107,N_10448);
or U13622 (N_13622,N_10866,N_11316);
and U13623 (N_13623,N_10757,N_9970);
nor U13624 (N_13624,N_11966,N_10470);
and U13625 (N_13625,N_11317,N_12367);
or U13626 (N_13626,N_12415,N_12042);
nor U13627 (N_13627,N_11126,N_10055);
or U13628 (N_13628,N_9589,N_12037);
and U13629 (N_13629,N_10860,N_11916);
and U13630 (N_13630,N_9874,N_10580);
and U13631 (N_13631,N_10874,N_9747);
nand U13632 (N_13632,N_10978,N_12248);
or U13633 (N_13633,N_9924,N_11241);
or U13634 (N_13634,N_11465,N_9746);
xnor U13635 (N_13635,N_9615,N_9934);
xnor U13636 (N_13636,N_9971,N_10513);
nor U13637 (N_13637,N_11453,N_10321);
nor U13638 (N_13638,N_11469,N_12046);
nor U13639 (N_13639,N_10148,N_10953);
nor U13640 (N_13640,N_11889,N_10064);
or U13641 (N_13641,N_10031,N_10645);
nor U13642 (N_13642,N_9644,N_10971);
nor U13643 (N_13643,N_11706,N_10196);
nor U13644 (N_13644,N_11089,N_9963);
nand U13645 (N_13645,N_10864,N_10688);
and U13646 (N_13646,N_11208,N_9932);
or U13647 (N_13647,N_11770,N_10101);
nand U13648 (N_13648,N_10687,N_12150);
nand U13649 (N_13649,N_11701,N_11599);
nand U13650 (N_13650,N_12117,N_10777);
and U13651 (N_13651,N_9712,N_9839);
or U13652 (N_13652,N_9387,N_10718);
and U13653 (N_13653,N_10008,N_11788);
or U13654 (N_13654,N_9673,N_10841);
and U13655 (N_13655,N_12484,N_10431);
and U13656 (N_13656,N_9804,N_11441);
xnor U13657 (N_13657,N_10499,N_10743);
or U13658 (N_13658,N_10400,N_11693);
nand U13659 (N_13659,N_9465,N_11512);
nand U13660 (N_13660,N_9420,N_11977);
nand U13661 (N_13661,N_10241,N_11115);
or U13662 (N_13662,N_9503,N_10220);
and U13663 (N_13663,N_11908,N_9775);
or U13664 (N_13664,N_9711,N_9705);
or U13665 (N_13665,N_10036,N_10479);
nand U13666 (N_13666,N_9601,N_9968);
nor U13667 (N_13667,N_10671,N_10795);
nor U13668 (N_13668,N_11064,N_9658);
and U13669 (N_13669,N_11295,N_11810);
or U13670 (N_13670,N_10798,N_11235);
and U13671 (N_13671,N_11746,N_10045);
nand U13672 (N_13672,N_11493,N_11504);
nor U13673 (N_13673,N_11267,N_10652);
or U13674 (N_13674,N_11603,N_10829);
and U13675 (N_13675,N_12079,N_11733);
nand U13676 (N_13676,N_9834,N_12287);
or U13677 (N_13677,N_11371,N_9776);
and U13678 (N_13678,N_10706,N_11887);
xnor U13679 (N_13679,N_12461,N_10542);
nor U13680 (N_13680,N_9920,N_10872);
nor U13681 (N_13681,N_12000,N_9574);
or U13682 (N_13682,N_12019,N_11234);
nor U13683 (N_13683,N_12202,N_11445);
nand U13684 (N_13684,N_9841,N_9412);
xor U13685 (N_13685,N_9693,N_11712);
xnor U13686 (N_13686,N_11423,N_9753);
nand U13687 (N_13687,N_12275,N_9690);
nand U13688 (N_13688,N_12331,N_11660);
and U13689 (N_13689,N_10822,N_10332);
and U13690 (N_13690,N_12175,N_11106);
nor U13691 (N_13691,N_11394,N_12412);
xor U13692 (N_13692,N_11948,N_9648);
nand U13693 (N_13693,N_12015,N_10516);
nand U13694 (N_13694,N_11284,N_11404);
nand U13695 (N_13695,N_11084,N_11937);
nand U13696 (N_13696,N_11353,N_12177);
nand U13697 (N_13697,N_9674,N_10861);
nor U13698 (N_13698,N_11705,N_12228);
xor U13699 (N_13699,N_10042,N_10630);
or U13700 (N_13700,N_9432,N_9608);
nand U13701 (N_13701,N_10500,N_10844);
and U13702 (N_13702,N_10723,N_12356);
nand U13703 (N_13703,N_10063,N_10783);
nor U13704 (N_13704,N_9847,N_9881);
or U13705 (N_13705,N_9559,N_10284);
or U13706 (N_13706,N_10225,N_9717);
or U13707 (N_13707,N_11002,N_11075);
nor U13708 (N_13708,N_10633,N_12250);
nand U13709 (N_13709,N_11102,N_12473);
or U13710 (N_13710,N_12007,N_11424);
and U13711 (N_13711,N_9417,N_12315);
and U13712 (N_13712,N_9619,N_12489);
xnor U13713 (N_13713,N_11790,N_10510);
and U13714 (N_13714,N_10568,N_10135);
or U13715 (N_13715,N_11564,N_11350);
nand U13716 (N_13716,N_9640,N_10331);
and U13717 (N_13717,N_10251,N_11169);
xnor U13718 (N_13718,N_11003,N_9883);
or U13719 (N_13719,N_11214,N_10105);
or U13720 (N_13720,N_9807,N_10033);
or U13721 (N_13721,N_11159,N_10075);
xnor U13722 (N_13722,N_10162,N_9416);
or U13723 (N_13723,N_9452,N_12039);
or U13724 (N_13724,N_12181,N_11309);
and U13725 (N_13725,N_11702,N_12457);
and U13726 (N_13726,N_12062,N_10788);
nor U13727 (N_13727,N_11986,N_10015);
nand U13728 (N_13728,N_12001,N_9688);
nand U13729 (N_13729,N_12151,N_9832);
nor U13730 (N_13730,N_10614,N_12188);
nand U13731 (N_13731,N_10014,N_10035);
nor U13732 (N_13732,N_12126,N_11294);
and U13733 (N_13733,N_9887,N_9818);
or U13734 (N_13734,N_10910,N_9999);
and U13735 (N_13735,N_12252,N_10450);
nor U13736 (N_13736,N_12372,N_10002);
and U13737 (N_13737,N_12127,N_9562);
nor U13738 (N_13738,N_11942,N_9539);
or U13739 (N_13739,N_12032,N_11382);
or U13740 (N_13740,N_11597,N_11239);
or U13741 (N_13741,N_11690,N_11412);
nand U13742 (N_13742,N_11254,N_11157);
xor U13743 (N_13743,N_9511,N_10851);
or U13744 (N_13744,N_10093,N_11911);
and U13745 (N_13745,N_11655,N_9377);
nand U13746 (N_13746,N_11152,N_10017);
or U13747 (N_13747,N_10276,N_11680);
or U13748 (N_13748,N_10768,N_11700);
nand U13749 (N_13749,N_10634,N_12280);
or U13750 (N_13750,N_10361,N_10752);
xor U13751 (N_13751,N_12197,N_12312);
or U13752 (N_13752,N_9817,N_12168);
or U13753 (N_13753,N_10131,N_11756);
nand U13754 (N_13754,N_9436,N_12494);
and U13755 (N_13755,N_9422,N_10065);
xnor U13756 (N_13756,N_11220,N_10300);
and U13757 (N_13757,N_9792,N_11878);
and U13758 (N_13758,N_9967,N_12187);
nand U13759 (N_13759,N_11121,N_10650);
and U13760 (N_13760,N_12245,N_10434);
and U13761 (N_13761,N_10235,N_12261);
xnor U13762 (N_13762,N_12120,N_11149);
nor U13763 (N_13763,N_11033,N_9397);
nor U13764 (N_13764,N_11783,N_12269);
and U13765 (N_13765,N_10211,N_11008);
nand U13766 (N_13766,N_12289,N_11368);
nand U13767 (N_13767,N_10799,N_10193);
and U13768 (N_13768,N_11769,N_10518);
and U13769 (N_13769,N_11602,N_10176);
and U13770 (N_13770,N_11110,N_10421);
and U13771 (N_13771,N_10804,N_12205);
nor U13772 (N_13772,N_10258,N_9469);
nand U13773 (N_13773,N_12361,N_9724);
nor U13774 (N_13774,N_9497,N_10371);
nand U13775 (N_13775,N_11111,N_12282);
nor U13776 (N_13776,N_12108,N_12132);
or U13777 (N_13777,N_12036,N_11784);
nand U13778 (N_13778,N_11983,N_11200);
nor U13779 (N_13779,N_12142,N_11505);
nand U13780 (N_13780,N_10086,N_9801);
and U13781 (N_13781,N_11238,N_11426);
or U13782 (N_13782,N_10309,N_9708);
nand U13783 (N_13783,N_11400,N_12476);
xnor U13784 (N_13784,N_9768,N_11227);
nand U13785 (N_13785,N_11091,N_10021);
or U13786 (N_13786,N_11509,N_10900);
nand U13787 (N_13787,N_12363,N_11776);
xor U13788 (N_13788,N_10558,N_10245);
and U13789 (N_13789,N_12354,N_10765);
nor U13790 (N_13790,N_11389,N_11486);
nor U13791 (N_13791,N_12194,N_11750);
nand U13792 (N_13792,N_11343,N_10020);
nand U13793 (N_13793,N_10865,N_10098);
nor U13794 (N_13794,N_11653,N_11145);
nor U13795 (N_13795,N_10139,N_12316);
nor U13796 (N_13796,N_10269,N_11077);
xor U13797 (N_13797,N_11041,N_10461);
nor U13798 (N_13798,N_11369,N_11020);
and U13799 (N_13799,N_9709,N_10112);
nor U13800 (N_13800,N_10859,N_11605);
and U13801 (N_13801,N_11463,N_9850);
nand U13802 (N_13802,N_9566,N_11506);
or U13803 (N_13803,N_12407,N_11007);
or U13804 (N_13804,N_9912,N_12450);
nor U13805 (N_13805,N_12279,N_11481);
and U13806 (N_13806,N_9592,N_10155);
nand U13807 (N_13807,N_12321,N_10190);
and U13808 (N_13808,N_9948,N_10345);
or U13809 (N_13809,N_11282,N_11437);
nor U13810 (N_13810,N_11307,N_9621);
nor U13811 (N_13811,N_11087,N_9633);
nor U13812 (N_13812,N_11454,N_10598);
or U13813 (N_13813,N_12020,N_11212);
nor U13814 (N_13814,N_9437,N_10547);
nand U13815 (N_13815,N_10951,N_10304);
nor U13816 (N_13816,N_12026,N_10158);
nand U13817 (N_13817,N_9470,N_9759);
nand U13818 (N_13818,N_12163,N_9869);
and U13819 (N_13819,N_10707,N_10301);
nand U13820 (N_13820,N_9931,N_12055);
and U13821 (N_13821,N_11187,N_9609);
nand U13822 (N_13822,N_11554,N_10629);
and U13823 (N_13823,N_9831,N_12044);
and U13824 (N_13824,N_10868,N_9444);
and U13825 (N_13825,N_9635,N_10779);
xor U13826 (N_13826,N_9980,N_10675);
nor U13827 (N_13827,N_12263,N_11982);
nand U13828 (N_13828,N_11270,N_12005);
nor U13829 (N_13829,N_10089,N_11545);
nand U13830 (N_13830,N_10273,N_9699);
and U13831 (N_13831,N_10281,N_12332);
nor U13832 (N_13832,N_11749,N_9514);
and U13833 (N_13833,N_11344,N_10751);
nor U13834 (N_13834,N_11360,N_12311);
or U13835 (N_13835,N_11024,N_10197);
or U13836 (N_13836,N_10726,N_9760);
or U13837 (N_13837,N_12447,N_9897);
and U13838 (N_13838,N_9504,N_12323);
and U13839 (N_13839,N_9385,N_9474);
nor U13840 (N_13840,N_12123,N_12298);
xor U13841 (N_13841,N_10905,N_9914);
nand U13842 (N_13842,N_9381,N_9406);
nor U13843 (N_13843,N_11978,N_12166);
xor U13844 (N_13844,N_10443,N_11860);
or U13845 (N_13845,N_9491,N_10381);
or U13846 (N_13846,N_11129,N_10920);
nor U13847 (N_13847,N_12304,N_12425);
or U13848 (N_13848,N_10810,N_9531);
nand U13849 (N_13849,N_11928,N_11954);
and U13850 (N_13850,N_11000,N_9509);
and U13851 (N_13851,N_10814,N_11013);
nor U13852 (N_13852,N_9443,N_11011);
or U13853 (N_13853,N_11416,N_10729);
or U13854 (N_13854,N_10895,N_9399);
nand U13855 (N_13855,N_11569,N_11901);
or U13856 (N_13856,N_9908,N_12225);
nor U13857 (N_13857,N_11312,N_9988);
nor U13858 (N_13858,N_10612,N_9438);
nand U13859 (N_13859,N_9884,N_10260);
nor U13860 (N_13860,N_9679,N_11740);
xor U13861 (N_13861,N_10506,N_11291);
and U13862 (N_13862,N_12174,N_9764);
nor U13863 (N_13863,N_10243,N_9992);
nand U13864 (N_13864,N_10674,N_9382);
nor U13865 (N_13865,N_12145,N_9647);
nor U13866 (N_13866,N_11537,N_11356);
and U13867 (N_13867,N_12462,N_10501);
or U13868 (N_13868,N_12423,N_11079);
nor U13869 (N_13869,N_9568,N_12160);
xnor U13870 (N_13870,N_9440,N_12227);
and U13871 (N_13871,N_11816,N_11848);
and U13872 (N_13872,N_11251,N_10483);
nor U13873 (N_13873,N_10030,N_12116);
and U13874 (N_13874,N_10081,N_12340);
nor U13875 (N_13875,N_12398,N_12335);
nand U13876 (N_13876,N_10480,N_11018);
nor U13877 (N_13877,N_9396,N_12391);
and U13878 (N_13878,N_11150,N_10072);
xnor U13879 (N_13879,N_10437,N_11327);
nand U13880 (N_13880,N_10078,N_10340);
xnor U13881 (N_13881,N_10774,N_10678);
or U13882 (N_13882,N_9423,N_9668);
xor U13883 (N_13883,N_10325,N_11442);
nor U13884 (N_13884,N_11581,N_10454);
and U13885 (N_13885,N_10474,N_10862);
or U13886 (N_13886,N_11785,N_11065);
nand U13887 (N_13887,N_10646,N_10142);
nor U13888 (N_13888,N_12077,N_9457);
and U13889 (N_13889,N_10491,N_12488);
nor U13890 (N_13890,N_10653,N_10395);
or U13891 (N_13891,N_12035,N_10763);
and U13892 (N_13892,N_11021,N_9473);
nor U13893 (N_13893,N_12219,N_10989);
nand U13894 (N_13894,N_9388,N_12157);
nor U13895 (N_13895,N_10557,N_11046);
xor U13896 (N_13896,N_12082,N_9512);
nor U13897 (N_13897,N_11631,N_9879);
nand U13898 (N_13898,N_11953,N_11517);
and U13899 (N_13899,N_12420,N_9803);
or U13900 (N_13900,N_12122,N_10333);
or U13901 (N_13901,N_10836,N_10517);
xnor U13902 (N_13902,N_9773,N_9575);
xnor U13903 (N_13903,N_10366,N_9515);
xnor U13904 (N_13904,N_10252,N_9954);
nand U13905 (N_13905,N_11373,N_12018);
or U13906 (N_13906,N_9537,N_9390);
nand U13907 (N_13907,N_10453,N_11514);
nor U13908 (N_13908,N_10061,N_12233);
nand U13909 (N_13909,N_9466,N_11707);
nor U13910 (N_13910,N_10425,N_10049);
nor U13911 (N_13911,N_12061,N_9756);
nand U13912 (N_13912,N_12343,N_11310);
or U13913 (N_13913,N_10096,N_10476);
xor U13914 (N_13914,N_9694,N_11028);
nand U13915 (N_13915,N_9446,N_10449);
and U13916 (N_13916,N_10415,N_11938);
nand U13917 (N_13917,N_10786,N_10392);
and U13918 (N_13918,N_9947,N_9556);
nor U13919 (N_13919,N_11645,N_10253);
and U13920 (N_13920,N_12057,N_12182);
or U13921 (N_13921,N_9591,N_10424);
nand U13922 (N_13922,N_10609,N_11950);
and U13923 (N_13923,N_11976,N_11721);
and U13924 (N_13924,N_11643,N_10374);
and U13925 (N_13925,N_9722,N_11759);
or U13926 (N_13926,N_9527,N_10635);
nor U13927 (N_13927,N_11448,N_10384);
or U13928 (N_13928,N_12104,N_9966);
nor U13929 (N_13929,N_10396,N_9586);
and U13930 (N_13930,N_10398,N_10521);
or U13931 (N_13931,N_10163,N_11376);
nand U13932 (N_13932,N_10237,N_12344);
or U13933 (N_13933,N_9888,N_10005);
or U13934 (N_13934,N_11912,N_9538);
xnor U13935 (N_13935,N_9376,N_11971);
nand U13936 (N_13936,N_9698,N_9687);
nor U13937 (N_13937,N_12374,N_10856);
nor U13938 (N_13938,N_9663,N_9393);
or U13939 (N_13939,N_9718,N_9520);
or U13940 (N_13940,N_11391,N_10389);
or U13941 (N_13941,N_10411,N_9997);
and U13942 (N_13942,N_12099,N_11897);
or U13943 (N_13943,N_12308,N_11933);
nor U13944 (N_13944,N_10019,N_10128);
and U13945 (N_13945,N_9822,N_12301);
nand U13946 (N_13946,N_10977,N_10878);
nand U13947 (N_13947,N_11132,N_10744);
xor U13948 (N_13948,N_10164,N_11250);
or U13949 (N_13949,N_9689,N_10124);
and U13950 (N_13950,N_10554,N_9830);
nand U13951 (N_13951,N_10545,N_9840);
nor U13952 (N_13952,N_11398,N_12134);
and U13953 (N_13953,N_11661,N_9979);
nor U13954 (N_13954,N_10157,N_10102);
and U13955 (N_13955,N_11973,N_9771);
and U13956 (N_13956,N_12414,N_9569);
or U13957 (N_13957,N_11466,N_10877);
xnor U13958 (N_13958,N_9600,N_10429);
or U13959 (N_13959,N_9969,N_9786);
xnor U13960 (N_13960,N_11892,N_10610);
nand U13961 (N_13961,N_12292,N_10223);
nor U13962 (N_13962,N_11585,N_12411);
nand U13963 (N_13963,N_11459,N_10924);
nand U13964 (N_13964,N_10803,N_9513);
nand U13965 (N_13965,N_9893,N_9476);
nor U13966 (N_13966,N_9602,N_11078);
xor U13967 (N_13967,N_9723,N_10775);
nor U13968 (N_13968,N_10813,N_10668);
or U13969 (N_13969,N_10849,N_11117);
nor U13970 (N_13970,N_11179,N_11794);
nor U13971 (N_13971,N_11185,N_10106);
or U13972 (N_13972,N_11300,N_10664);
nand U13973 (N_13973,N_11383,N_11949);
or U13974 (N_13974,N_11406,N_10887);
or U13975 (N_13975,N_11477,N_10839);
and U13976 (N_13976,N_11456,N_11036);
or U13977 (N_13977,N_9758,N_10426);
and U13978 (N_13978,N_11625,N_9380);
and U13979 (N_13979,N_10271,N_12152);
nor U13980 (N_13980,N_11165,N_12443);
or U13981 (N_13981,N_10141,N_9558);
and U13982 (N_13982,N_10477,N_11026);
or U13983 (N_13983,N_9550,N_9911);
or U13984 (N_13984,N_11249,N_12442);
or U13985 (N_13985,N_10239,N_10524);
nor U13986 (N_13986,N_9860,N_10543);
nor U13987 (N_13987,N_11751,N_11256);
nand U13988 (N_13988,N_12496,N_10410);
nand U13989 (N_13989,N_11943,N_12011);
nand U13990 (N_13990,N_10487,N_11005);
nor U13991 (N_13991,N_11236,N_12474);
or U13992 (N_13992,N_9902,N_12326);
xor U13993 (N_13993,N_11218,N_11488);
and U13994 (N_13994,N_12368,N_11377);
and U13995 (N_13995,N_12051,N_11857);
nor U13996 (N_13996,N_10631,N_11743);
xor U13997 (N_13997,N_11092,N_11612);
nor U13998 (N_13998,N_11379,N_10254);
and U13999 (N_13999,N_9885,N_12113);
nor U14000 (N_14000,N_9492,N_12180);
nor U14001 (N_14001,N_10010,N_10484);
nand U14002 (N_14002,N_10662,N_11601);
or U14003 (N_14003,N_11896,N_10409);
nand U14004 (N_14004,N_11862,N_10957);
nor U14005 (N_14005,N_9605,N_11592);
or U14006 (N_14006,N_11082,N_9645);
nand U14007 (N_14007,N_10770,N_12063);
or U14008 (N_14008,N_11910,N_12422);
nor U14009 (N_14009,N_12068,N_11884);
or U14010 (N_14010,N_11362,N_12380);
or U14011 (N_14011,N_11427,N_11263);
or U14012 (N_14012,N_9487,N_11922);
nor U14013 (N_14013,N_11828,N_9451);
nand U14014 (N_14014,N_12124,N_10307);
nand U14015 (N_14015,N_9639,N_10110);
and U14016 (N_14016,N_10852,N_11124);
nand U14017 (N_14017,N_12224,N_11628);
or U14018 (N_14018,N_12119,N_11446);
nand U14019 (N_14019,N_11548,N_9928);
or U14020 (N_14020,N_10593,N_11288);
nor U14021 (N_14021,N_10438,N_10885);
and U14022 (N_14022,N_11068,N_12110);
nand U14023 (N_14023,N_9863,N_11266);
or U14024 (N_14024,N_11211,N_9607);
nand U14025 (N_14025,N_10733,N_10745);
or U14026 (N_14026,N_10880,N_10023);
or U14027 (N_14027,N_10628,N_11530);
or U14028 (N_14028,N_9529,N_12208);
nor U14029 (N_14029,N_10032,N_10475);
or U14030 (N_14030,N_10574,N_10960);
nand U14031 (N_14031,N_10430,N_10945);
or U14032 (N_14032,N_11972,N_9794);
or U14033 (N_14033,N_12161,N_10165);
and U14034 (N_14034,N_12064,N_11074);
nor U14035 (N_14035,N_10232,N_10236);
or U14036 (N_14036,N_10359,N_11951);
nand U14037 (N_14037,N_11302,N_9462);
xor U14038 (N_14038,N_10356,N_11697);
nand U14039 (N_14039,N_11620,N_9867);
nand U14040 (N_14040,N_11970,N_9407);
and U14041 (N_14041,N_11575,N_11566);
and U14042 (N_14042,N_10209,N_10326);
and U14043 (N_14043,N_12469,N_9977);
and U14044 (N_14044,N_10589,N_9447);
xnor U14045 (N_14045,N_9742,N_9955);
or U14046 (N_14046,N_10386,N_10401);
nor U14047 (N_14047,N_9394,N_10902);
xnor U14048 (N_14048,N_10537,N_12377);
or U14049 (N_14049,N_10700,N_11623);
or U14050 (N_14050,N_11341,N_11513);
nand U14051 (N_14051,N_11807,N_11375);
or U14052 (N_14052,N_11228,N_12017);
nand U14053 (N_14053,N_11168,N_10869);
nor U14054 (N_14054,N_10816,N_11562);
xor U14055 (N_14055,N_11714,N_11987);
or U14056 (N_14056,N_10846,N_9835);
xor U14057 (N_14057,N_12139,N_10314);
nor U14058 (N_14058,N_11923,N_11120);
nor U14059 (N_14059,N_12072,N_12102);
and U14060 (N_14060,N_10060,N_12401);
nor U14061 (N_14061,N_11054,N_11433);
and U14062 (N_14062,N_10523,N_11725);
nor U14063 (N_14063,N_10162,N_10844);
nand U14064 (N_14064,N_11263,N_10715);
or U14065 (N_14065,N_10829,N_12333);
and U14066 (N_14066,N_9866,N_10412);
or U14067 (N_14067,N_12275,N_10394);
nand U14068 (N_14068,N_12253,N_11429);
and U14069 (N_14069,N_10284,N_10736);
xor U14070 (N_14070,N_9694,N_10249);
or U14071 (N_14071,N_10197,N_10929);
and U14072 (N_14072,N_9432,N_11283);
nor U14073 (N_14073,N_11474,N_11422);
xor U14074 (N_14074,N_11553,N_12370);
and U14075 (N_14075,N_11698,N_9768);
or U14076 (N_14076,N_10019,N_11111);
and U14077 (N_14077,N_12453,N_9905);
nor U14078 (N_14078,N_11306,N_10260);
and U14079 (N_14079,N_10036,N_12438);
and U14080 (N_14080,N_11696,N_11525);
and U14081 (N_14081,N_10227,N_12480);
nor U14082 (N_14082,N_10148,N_10364);
nand U14083 (N_14083,N_11664,N_12449);
nand U14084 (N_14084,N_10891,N_11407);
xnor U14085 (N_14085,N_9660,N_11041);
nor U14086 (N_14086,N_9847,N_12061);
or U14087 (N_14087,N_11048,N_9873);
and U14088 (N_14088,N_11035,N_11962);
or U14089 (N_14089,N_9755,N_11087);
nand U14090 (N_14090,N_10295,N_11985);
and U14091 (N_14091,N_10542,N_12027);
nand U14092 (N_14092,N_10300,N_11877);
and U14093 (N_14093,N_11594,N_10361);
or U14094 (N_14094,N_9682,N_11532);
and U14095 (N_14095,N_12403,N_11892);
nor U14096 (N_14096,N_10022,N_12244);
xor U14097 (N_14097,N_10222,N_11092);
nor U14098 (N_14098,N_11197,N_11098);
nor U14099 (N_14099,N_12326,N_10934);
nor U14100 (N_14100,N_9896,N_12067);
or U14101 (N_14101,N_11438,N_11540);
nand U14102 (N_14102,N_9501,N_12246);
nor U14103 (N_14103,N_9402,N_11240);
xnor U14104 (N_14104,N_10359,N_10442);
and U14105 (N_14105,N_10513,N_10087);
or U14106 (N_14106,N_11257,N_10024);
nand U14107 (N_14107,N_12325,N_9602);
or U14108 (N_14108,N_11259,N_9445);
and U14109 (N_14109,N_10642,N_12209);
nor U14110 (N_14110,N_9477,N_11271);
and U14111 (N_14111,N_10165,N_12287);
and U14112 (N_14112,N_11759,N_10488);
and U14113 (N_14113,N_11669,N_12049);
and U14114 (N_14114,N_11156,N_11935);
or U14115 (N_14115,N_10261,N_11391);
and U14116 (N_14116,N_10778,N_10161);
nor U14117 (N_14117,N_10613,N_11766);
and U14118 (N_14118,N_11128,N_9495);
xnor U14119 (N_14119,N_9473,N_10253);
xnor U14120 (N_14120,N_10802,N_9826);
nand U14121 (N_14121,N_10266,N_9985);
nor U14122 (N_14122,N_9908,N_10592);
or U14123 (N_14123,N_9442,N_10020);
and U14124 (N_14124,N_10800,N_9550);
nand U14125 (N_14125,N_11667,N_10227);
nor U14126 (N_14126,N_10486,N_12009);
xnor U14127 (N_14127,N_12490,N_12427);
or U14128 (N_14128,N_12129,N_12435);
nor U14129 (N_14129,N_12482,N_9618);
and U14130 (N_14130,N_10475,N_11343);
and U14131 (N_14131,N_10587,N_9897);
nor U14132 (N_14132,N_12307,N_11532);
nand U14133 (N_14133,N_9984,N_11461);
or U14134 (N_14134,N_10857,N_11810);
and U14135 (N_14135,N_10732,N_10655);
and U14136 (N_14136,N_9525,N_11071);
or U14137 (N_14137,N_11154,N_10580);
and U14138 (N_14138,N_10943,N_12135);
and U14139 (N_14139,N_12190,N_12010);
nand U14140 (N_14140,N_11236,N_11962);
and U14141 (N_14141,N_9530,N_10734);
or U14142 (N_14142,N_11900,N_12207);
nand U14143 (N_14143,N_9509,N_11658);
or U14144 (N_14144,N_11295,N_12108);
nor U14145 (N_14145,N_12168,N_9457);
and U14146 (N_14146,N_11392,N_9897);
or U14147 (N_14147,N_11777,N_11199);
xor U14148 (N_14148,N_11966,N_10100);
nand U14149 (N_14149,N_11519,N_10485);
nor U14150 (N_14150,N_11693,N_11227);
nor U14151 (N_14151,N_10155,N_10385);
or U14152 (N_14152,N_12356,N_11142);
nor U14153 (N_14153,N_10749,N_9661);
xor U14154 (N_14154,N_11986,N_10140);
or U14155 (N_14155,N_9897,N_11262);
or U14156 (N_14156,N_10208,N_9417);
nor U14157 (N_14157,N_10055,N_10872);
xnor U14158 (N_14158,N_9751,N_10172);
nand U14159 (N_14159,N_11378,N_12360);
nand U14160 (N_14160,N_10032,N_10922);
nor U14161 (N_14161,N_10900,N_9411);
or U14162 (N_14162,N_10217,N_12341);
and U14163 (N_14163,N_9994,N_9885);
nor U14164 (N_14164,N_12175,N_11679);
or U14165 (N_14165,N_11387,N_9655);
and U14166 (N_14166,N_10267,N_11865);
nand U14167 (N_14167,N_10688,N_10573);
nand U14168 (N_14168,N_10028,N_10604);
and U14169 (N_14169,N_11363,N_9395);
nand U14170 (N_14170,N_10808,N_10023);
or U14171 (N_14171,N_12052,N_11443);
or U14172 (N_14172,N_12203,N_10889);
nor U14173 (N_14173,N_11840,N_10803);
or U14174 (N_14174,N_10572,N_10493);
nand U14175 (N_14175,N_11327,N_11739);
nor U14176 (N_14176,N_10245,N_9527);
nor U14177 (N_14177,N_11914,N_12160);
nand U14178 (N_14178,N_10164,N_10714);
nand U14179 (N_14179,N_10542,N_11180);
nor U14180 (N_14180,N_10365,N_12437);
or U14181 (N_14181,N_11711,N_10791);
nand U14182 (N_14182,N_9813,N_11035);
nand U14183 (N_14183,N_11162,N_11624);
xor U14184 (N_14184,N_12292,N_9658);
nor U14185 (N_14185,N_10311,N_11218);
and U14186 (N_14186,N_10303,N_11500);
and U14187 (N_14187,N_10204,N_10062);
nand U14188 (N_14188,N_11226,N_9447);
and U14189 (N_14189,N_11677,N_11223);
nand U14190 (N_14190,N_9700,N_9479);
and U14191 (N_14191,N_9852,N_10205);
or U14192 (N_14192,N_9561,N_10474);
nor U14193 (N_14193,N_9640,N_11486);
nor U14194 (N_14194,N_10879,N_9943);
nor U14195 (N_14195,N_10445,N_10957);
xor U14196 (N_14196,N_11994,N_9759);
and U14197 (N_14197,N_9589,N_11267);
and U14198 (N_14198,N_11087,N_10401);
and U14199 (N_14199,N_10703,N_10632);
nand U14200 (N_14200,N_10289,N_11579);
nor U14201 (N_14201,N_12189,N_10321);
nand U14202 (N_14202,N_10058,N_9568);
and U14203 (N_14203,N_12083,N_11281);
nand U14204 (N_14204,N_11371,N_10142);
nand U14205 (N_14205,N_10591,N_12402);
nor U14206 (N_14206,N_11768,N_9862);
or U14207 (N_14207,N_10754,N_11679);
nand U14208 (N_14208,N_12268,N_11076);
nand U14209 (N_14209,N_9910,N_9464);
or U14210 (N_14210,N_11985,N_9948);
and U14211 (N_14211,N_10140,N_12361);
nand U14212 (N_14212,N_12165,N_10039);
xnor U14213 (N_14213,N_12450,N_11134);
nor U14214 (N_14214,N_9707,N_11311);
and U14215 (N_14215,N_11959,N_10395);
or U14216 (N_14216,N_11869,N_10429);
or U14217 (N_14217,N_12140,N_9790);
or U14218 (N_14218,N_11561,N_10869);
and U14219 (N_14219,N_12357,N_9658);
and U14220 (N_14220,N_10740,N_12496);
and U14221 (N_14221,N_10786,N_11909);
xor U14222 (N_14222,N_10934,N_11139);
nand U14223 (N_14223,N_10117,N_9652);
nand U14224 (N_14224,N_10289,N_9824);
nand U14225 (N_14225,N_9509,N_10806);
xor U14226 (N_14226,N_9551,N_9897);
or U14227 (N_14227,N_10331,N_11437);
nor U14228 (N_14228,N_11714,N_9779);
nor U14229 (N_14229,N_10299,N_11704);
or U14230 (N_14230,N_9726,N_11368);
or U14231 (N_14231,N_11305,N_11986);
nand U14232 (N_14232,N_10355,N_11179);
or U14233 (N_14233,N_10862,N_11717);
or U14234 (N_14234,N_9502,N_9882);
nand U14235 (N_14235,N_9864,N_11676);
or U14236 (N_14236,N_11679,N_9592);
and U14237 (N_14237,N_10279,N_12249);
and U14238 (N_14238,N_11870,N_11748);
and U14239 (N_14239,N_12108,N_10537);
or U14240 (N_14240,N_10817,N_11003);
and U14241 (N_14241,N_11226,N_11275);
nand U14242 (N_14242,N_11708,N_9829);
xnor U14243 (N_14243,N_10266,N_11622);
or U14244 (N_14244,N_10489,N_10826);
or U14245 (N_14245,N_11970,N_10382);
nand U14246 (N_14246,N_9955,N_10955);
and U14247 (N_14247,N_11273,N_9582);
xor U14248 (N_14248,N_12061,N_11245);
or U14249 (N_14249,N_9718,N_12236);
nand U14250 (N_14250,N_9880,N_11804);
nor U14251 (N_14251,N_10776,N_11382);
nand U14252 (N_14252,N_11664,N_11560);
and U14253 (N_14253,N_9513,N_9691);
nor U14254 (N_14254,N_12136,N_10654);
or U14255 (N_14255,N_10807,N_10049);
and U14256 (N_14256,N_10933,N_10657);
or U14257 (N_14257,N_10852,N_11438);
and U14258 (N_14258,N_11793,N_9454);
or U14259 (N_14259,N_11623,N_9495);
xor U14260 (N_14260,N_10782,N_9758);
nor U14261 (N_14261,N_12048,N_11006);
nor U14262 (N_14262,N_11743,N_10856);
nor U14263 (N_14263,N_11524,N_11653);
and U14264 (N_14264,N_9542,N_10919);
xor U14265 (N_14265,N_9940,N_12095);
or U14266 (N_14266,N_12207,N_10564);
nor U14267 (N_14267,N_10120,N_10741);
nor U14268 (N_14268,N_11162,N_10786);
nor U14269 (N_14269,N_12342,N_11563);
and U14270 (N_14270,N_11421,N_10388);
nand U14271 (N_14271,N_11246,N_9791);
xnor U14272 (N_14272,N_12073,N_11152);
or U14273 (N_14273,N_10494,N_10072);
nor U14274 (N_14274,N_10550,N_11845);
and U14275 (N_14275,N_11547,N_10217);
and U14276 (N_14276,N_9453,N_9801);
nand U14277 (N_14277,N_10491,N_10054);
nor U14278 (N_14278,N_9698,N_12460);
and U14279 (N_14279,N_11194,N_10049);
nand U14280 (N_14280,N_10625,N_10915);
or U14281 (N_14281,N_11461,N_10726);
and U14282 (N_14282,N_11067,N_10613);
and U14283 (N_14283,N_10896,N_10995);
nand U14284 (N_14284,N_10700,N_9597);
and U14285 (N_14285,N_9723,N_10245);
nor U14286 (N_14286,N_10527,N_10337);
or U14287 (N_14287,N_10269,N_10934);
nor U14288 (N_14288,N_11675,N_12211);
nor U14289 (N_14289,N_11316,N_11307);
nor U14290 (N_14290,N_11062,N_11991);
xor U14291 (N_14291,N_12203,N_10478);
nand U14292 (N_14292,N_10662,N_9607);
nand U14293 (N_14293,N_10167,N_11417);
and U14294 (N_14294,N_10538,N_10825);
nor U14295 (N_14295,N_12096,N_9758);
and U14296 (N_14296,N_10956,N_11715);
nor U14297 (N_14297,N_9874,N_9589);
or U14298 (N_14298,N_12326,N_9408);
xor U14299 (N_14299,N_10908,N_10688);
and U14300 (N_14300,N_10507,N_10851);
xnor U14301 (N_14301,N_11657,N_10703);
or U14302 (N_14302,N_10524,N_11645);
nor U14303 (N_14303,N_10813,N_9805);
xor U14304 (N_14304,N_12044,N_11962);
or U14305 (N_14305,N_11933,N_9518);
nor U14306 (N_14306,N_11161,N_10525);
and U14307 (N_14307,N_11851,N_12136);
nor U14308 (N_14308,N_9761,N_10489);
nor U14309 (N_14309,N_11830,N_11106);
or U14310 (N_14310,N_11115,N_11377);
xnor U14311 (N_14311,N_12101,N_10173);
and U14312 (N_14312,N_10463,N_12151);
nand U14313 (N_14313,N_12097,N_12116);
nor U14314 (N_14314,N_9717,N_9627);
xnor U14315 (N_14315,N_9387,N_10203);
nand U14316 (N_14316,N_10352,N_12348);
or U14317 (N_14317,N_9445,N_11185);
xor U14318 (N_14318,N_11140,N_9950);
or U14319 (N_14319,N_9940,N_12156);
xor U14320 (N_14320,N_10113,N_11579);
nor U14321 (N_14321,N_9528,N_9905);
or U14322 (N_14322,N_12263,N_9814);
or U14323 (N_14323,N_11289,N_11537);
and U14324 (N_14324,N_9899,N_10127);
nor U14325 (N_14325,N_10141,N_11461);
or U14326 (N_14326,N_10687,N_12486);
and U14327 (N_14327,N_10293,N_11290);
nand U14328 (N_14328,N_10142,N_11991);
nor U14329 (N_14329,N_9454,N_11936);
and U14330 (N_14330,N_11983,N_11590);
nor U14331 (N_14331,N_12064,N_12309);
and U14332 (N_14332,N_9486,N_10310);
nor U14333 (N_14333,N_9985,N_10986);
nand U14334 (N_14334,N_10462,N_11062);
or U14335 (N_14335,N_12136,N_11349);
and U14336 (N_14336,N_10376,N_9793);
and U14337 (N_14337,N_11185,N_11384);
nor U14338 (N_14338,N_10229,N_12490);
nor U14339 (N_14339,N_12182,N_11938);
nand U14340 (N_14340,N_12088,N_12394);
nor U14341 (N_14341,N_11779,N_12103);
nand U14342 (N_14342,N_12419,N_12435);
xnor U14343 (N_14343,N_11810,N_11682);
nand U14344 (N_14344,N_9838,N_11261);
or U14345 (N_14345,N_9716,N_11010);
xnor U14346 (N_14346,N_9968,N_11367);
or U14347 (N_14347,N_11208,N_11752);
nor U14348 (N_14348,N_12261,N_9419);
and U14349 (N_14349,N_10894,N_10453);
and U14350 (N_14350,N_10290,N_11527);
and U14351 (N_14351,N_12009,N_11006);
xor U14352 (N_14352,N_11178,N_9769);
and U14353 (N_14353,N_9423,N_12031);
nor U14354 (N_14354,N_9440,N_11704);
or U14355 (N_14355,N_10416,N_11046);
and U14356 (N_14356,N_10769,N_11410);
nand U14357 (N_14357,N_10665,N_10159);
or U14358 (N_14358,N_10963,N_10009);
xor U14359 (N_14359,N_10658,N_11907);
nor U14360 (N_14360,N_9680,N_11041);
or U14361 (N_14361,N_10583,N_9956);
and U14362 (N_14362,N_11525,N_11164);
nand U14363 (N_14363,N_10082,N_11022);
nand U14364 (N_14364,N_12099,N_9852);
nor U14365 (N_14365,N_12027,N_11881);
or U14366 (N_14366,N_10658,N_10409);
and U14367 (N_14367,N_9529,N_10369);
or U14368 (N_14368,N_11271,N_12238);
nand U14369 (N_14369,N_11679,N_11397);
nand U14370 (N_14370,N_9744,N_11285);
nand U14371 (N_14371,N_12299,N_10166);
nor U14372 (N_14372,N_11901,N_10760);
or U14373 (N_14373,N_11442,N_10966);
or U14374 (N_14374,N_12287,N_11694);
nand U14375 (N_14375,N_11937,N_11026);
or U14376 (N_14376,N_11299,N_11871);
or U14377 (N_14377,N_10914,N_9666);
nor U14378 (N_14378,N_10161,N_10077);
and U14379 (N_14379,N_9989,N_10332);
xor U14380 (N_14380,N_11563,N_10201);
nand U14381 (N_14381,N_11399,N_12077);
or U14382 (N_14382,N_10749,N_12062);
and U14383 (N_14383,N_10543,N_11257);
and U14384 (N_14384,N_10114,N_11330);
nor U14385 (N_14385,N_9950,N_11150);
nand U14386 (N_14386,N_10949,N_10569);
nor U14387 (N_14387,N_11075,N_10912);
and U14388 (N_14388,N_12461,N_11468);
nor U14389 (N_14389,N_12383,N_10725);
or U14390 (N_14390,N_9837,N_10935);
nand U14391 (N_14391,N_10595,N_9595);
or U14392 (N_14392,N_10481,N_11927);
nor U14393 (N_14393,N_12159,N_9534);
and U14394 (N_14394,N_9684,N_12340);
xor U14395 (N_14395,N_11193,N_12113);
or U14396 (N_14396,N_11455,N_11904);
or U14397 (N_14397,N_10221,N_10961);
or U14398 (N_14398,N_11640,N_12434);
nand U14399 (N_14399,N_12220,N_10035);
and U14400 (N_14400,N_11761,N_11940);
and U14401 (N_14401,N_11176,N_11220);
nand U14402 (N_14402,N_9540,N_11404);
xnor U14403 (N_14403,N_11549,N_11759);
nand U14404 (N_14404,N_10218,N_9531);
and U14405 (N_14405,N_9816,N_9626);
nand U14406 (N_14406,N_11771,N_10663);
nor U14407 (N_14407,N_12423,N_11227);
nor U14408 (N_14408,N_12235,N_9525);
xnor U14409 (N_14409,N_12095,N_10623);
nor U14410 (N_14410,N_12085,N_11560);
or U14411 (N_14411,N_9649,N_11131);
or U14412 (N_14412,N_10904,N_11696);
xor U14413 (N_14413,N_10923,N_11390);
xnor U14414 (N_14414,N_11477,N_11339);
nand U14415 (N_14415,N_11225,N_10801);
nand U14416 (N_14416,N_9560,N_11349);
or U14417 (N_14417,N_9880,N_11922);
or U14418 (N_14418,N_10546,N_10796);
nor U14419 (N_14419,N_10741,N_10055);
nand U14420 (N_14420,N_10587,N_9995);
nand U14421 (N_14421,N_10697,N_10536);
nor U14422 (N_14422,N_11248,N_11425);
and U14423 (N_14423,N_11899,N_10365);
nor U14424 (N_14424,N_11060,N_12310);
and U14425 (N_14425,N_12405,N_9471);
nand U14426 (N_14426,N_10838,N_11250);
or U14427 (N_14427,N_11728,N_11371);
nand U14428 (N_14428,N_11104,N_11428);
nor U14429 (N_14429,N_11642,N_11846);
or U14430 (N_14430,N_10289,N_11685);
and U14431 (N_14431,N_12109,N_10668);
nor U14432 (N_14432,N_9632,N_12067);
nor U14433 (N_14433,N_12379,N_11896);
or U14434 (N_14434,N_11589,N_12382);
nand U14435 (N_14435,N_9773,N_11905);
or U14436 (N_14436,N_11826,N_11911);
xnor U14437 (N_14437,N_10381,N_9767);
and U14438 (N_14438,N_12153,N_9960);
or U14439 (N_14439,N_9510,N_9497);
and U14440 (N_14440,N_9411,N_11171);
xor U14441 (N_14441,N_9378,N_10157);
or U14442 (N_14442,N_10879,N_9845);
xnor U14443 (N_14443,N_11214,N_11396);
and U14444 (N_14444,N_10848,N_11521);
and U14445 (N_14445,N_11380,N_11278);
and U14446 (N_14446,N_9921,N_11587);
or U14447 (N_14447,N_11363,N_12340);
nand U14448 (N_14448,N_10533,N_11344);
and U14449 (N_14449,N_12105,N_9586);
nor U14450 (N_14450,N_11096,N_9768);
nor U14451 (N_14451,N_9589,N_12140);
nand U14452 (N_14452,N_11028,N_9693);
and U14453 (N_14453,N_11308,N_10727);
and U14454 (N_14454,N_12238,N_9773);
nand U14455 (N_14455,N_11041,N_10615);
nand U14456 (N_14456,N_9507,N_10944);
nand U14457 (N_14457,N_10405,N_10734);
or U14458 (N_14458,N_10498,N_10437);
and U14459 (N_14459,N_12469,N_12219);
xor U14460 (N_14460,N_10614,N_11248);
and U14461 (N_14461,N_11132,N_10221);
and U14462 (N_14462,N_9726,N_11780);
nor U14463 (N_14463,N_10524,N_11521);
and U14464 (N_14464,N_9672,N_10215);
and U14465 (N_14465,N_10874,N_10395);
nand U14466 (N_14466,N_9645,N_11622);
nand U14467 (N_14467,N_10641,N_9744);
and U14468 (N_14468,N_10077,N_11686);
or U14469 (N_14469,N_12496,N_10159);
or U14470 (N_14470,N_12236,N_12216);
nor U14471 (N_14471,N_11861,N_12457);
and U14472 (N_14472,N_12012,N_9990);
xor U14473 (N_14473,N_12211,N_10227);
nor U14474 (N_14474,N_9927,N_12307);
xor U14475 (N_14475,N_10524,N_11441);
nor U14476 (N_14476,N_11230,N_9470);
nor U14477 (N_14477,N_10004,N_11265);
nor U14478 (N_14478,N_11841,N_10716);
nor U14479 (N_14479,N_9823,N_10540);
and U14480 (N_14480,N_10252,N_11077);
nand U14481 (N_14481,N_12343,N_10687);
xnor U14482 (N_14482,N_10789,N_11934);
and U14483 (N_14483,N_9435,N_10029);
nor U14484 (N_14484,N_10348,N_12361);
nor U14485 (N_14485,N_9982,N_10128);
and U14486 (N_14486,N_11542,N_9457);
or U14487 (N_14487,N_10538,N_12142);
nor U14488 (N_14488,N_11964,N_11376);
nand U14489 (N_14489,N_11733,N_9866);
and U14490 (N_14490,N_10502,N_12375);
or U14491 (N_14491,N_11903,N_11688);
and U14492 (N_14492,N_10273,N_11178);
nor U14493 (N_14493,N_10498,N_9908);
and U14494 (N_14494,N_10843,N_10914);
nor U14495 (N_14495,N_9627,N_11206);
nor U14496 (N_14496,N_9794,N_10885);
xnor U14497 (N_14497,N_11490,N_12437);
nand U14498 (N_14498,N_10390,N_12309);
or U14499 (N_14499,N_10650,N_10056);
xnor U14500 (N_14500,N_9423,N_10046);
and U14501 (N_14501,N_10482,N_12085);
nor U14502 (N_14502,N_12365,N_10201);
or U14503 (N_14503,N_10725,N_12152);
xnor U14504 (N_14504,N_9439,N_11756);
or U14505 (N_14505,N_11813,N_9964);
nand U14506 (N_14506,N_10480,N_11193);
xor U14507 (N_14507,N_11805,N_12081);
nor U14508 (N_14508,N_10048,N_10749);
nand U14509 (N_14509,N_11903,N_10006);
nor U14510 (N_14510,N_10688,N_10467);
or U14511 (N_14511,N_11324,N_10450);
and U14512 (N_14512,N_11074,N_10595);
nand U14513 (N_14513,N_11771,N_11644);
nor U14514 (N_14514,N_9696,N_10879);
or U14515 (N_14515,N_10501,N_11966);
nand U14516 (N_14516,N_11740,N_11332);
nor U14517 (N_14517,N_11118,N_10291);
and U14518 (N_14518,N_12161,N_9942);
and U14519 (N_14519,N_9434,N_12464);
and U14520 (N_14520,N_10292,N_10144);
nand U14521 (N_14521,N_11865,N_12387);
nand U14522 (N_14522,N_10984,N_9560);
nor U14523 (N_14523,N_11854,N_12359);
nand U14524 (N_14524,N_11773,N_11432);
or U14525 (N_14525,N_11131,N_10085);
xor U14526 (N_14526,N_11876,N_12410);
nor U14527 (N_14527,N_11929,N_11448);
xor U14528 (N_14528,N_12425,N_11657);
nand U14529 (N_14529,N_10061,N_10430);
and U14530 (N_14530,N_10138,N_10729);
and U14531 (N_14531,N_9387,N_11777);
or U14532 (N_14532,N_11679,N_10255);
or U14533 (N_14533,N_11432,N_12322);
nor U14534 (N_14534,N_11495,N_10418);
nor U14535 (N_14535,N_11716,N_11456);
and U14536 (N_14536,N_10046,N_11321);
and U14537 (N_14537,N_9467,N_12028);
nand U14538 (N_14538,N_9489,N_9875);
and U14539 (N_14539,N_10397,N_11881);
xor U14540 (N_14540,N_10270,N_11831);
or U14541 (N_14541,N_10929,N_12327);
and U14542 (N_14542,N_10374,N_10096);
nand U14543 (N_14543,N_12385,N_12207);
xor U14544 (N_14544,N_11997,N_9435);
or U14545 (N_14545,N_11087,N_12112);
and U14546 (N_14546,N_11480,N_11190);
or U14547 (N_14547,N_11053,N_12313);
or U14548 (N_14548,N_11481,N_10031);
and U14549 (N_14549,N_10598,N_12190);
nand U14550 (N_14550,N_10758,N_11412);
nand U14551 (N_14551,N_9944,N_11320);
nor U14552 (N_14552,N_10609,N_10516);
and U14553 (N_14553,N_10606,N_10964);
nor U14554 (N_14554,N_9382,N_12117);
nor U14555 (N_14555,N_11294,N_10503);
or U14556 (N_14556,N_9474,N_10677);
or U14557 (N_14557,N_12410,N_9620);
or U14558 (N_14558,N_11506,N_10543);
or U14559 (N_14559,N_11936,N_9554);
xnor U14560 (N_14560,N_10053,N_11101);
nor U14561 (N_14561,N_10175,N_11633);
xnor U14562 (N_14562,N_11039,N_9395);
and U14563 (N_14563,N_11965,N_12042);
or U14564 (N_14564,N_10476,N_9406);
or U14565 (N_14565,N_10822,N_10042);
nand U14566 (N_14566,N_9923,N_12214);
nor U14567 (N_14567,N_11939,N_10528);
nand U14568 (N_14568,N_10323,N_11728);
or U14569 (N_14569,N_9746,N_12315);
nor U14570 (N_14570,N_9424,N_11446);
nor U14571 (N_14571,N_10029,N_10881);
and U14572 (N_14572,N_10293,N_9731);
nor U14573 (N_14573,N_10036,N_10853);
and U14574 (N_14574,N_11461,N_9968);
nor U14575 (N_14575,N_10806,N_10234);
or U14576 (N_14576,N_12151,N_10483);
nand U14577 (N_14577,N_12014,N_10606);
and U14578 (N_14578,N_9513,N_10135);
or U14579 (N_14579,N_12218,N_10265);
or U14580 (N_14580,N_9587,N_10176);
xnor U14581 (N_14581,N_11389,N_9713);
and U14582 (N_14582,N_11845,N_12152);
nand U14583 (N_14583,N_12341,N_12239);
nand U14584 (N_14584,N_10092,N_11075);
or U14585 (N_14585,N_10853,N_9524);
or U14586 (N_14586,N_10394,N_11533);
and U14587 (N_14587,N_9775,N_11313);
and U14588 (N_14588,N_11212,N_9655);
nor U14589 (N_14589,N_9830,N_9941);
and U14590 (N_14590,N_11457,N_10597);
nand U14591 (N_14591,N_10749,N_11687);
nand U14592 (N_14592,N_11140,N_10472);
nor U14593 (N_14593,N_10330,N_11119);
nand U14594 (N_14594,N_12400,N_10790);
and U14595 (N_14595,N_10931,N_12490);
and U14596 (N_14596,N_9970,N_10036);
or U14597 (N_14597,N_12093,N_10847);
and U14598 (N_14598,N_10898,N_10325);
and U14599 (N_14599,N_10549,N_10760);
and U14600 (N_14600,N_9473,N_9947);
nand U14601 (N_14601,N_11782,N_11069);
and U14602 (N_14602,N_10125,N_11482);
nand U14603 (N_14603,N_11475,N_12118);
nor U14604 (N_14604,N_11205,N_11319);
or U14605 (N_14605,N_11359,N_12116);
nand U14606 (N_14606,N_12041,N_12372);
nor U14607 (N_14607,N_11667,N_11080);
or U14608 (N_14608,N_10964,N_12487);
nand U14609 (N_14609,N_9995,N_11979);
nor U14610 (N_14610,N_9603,N_9446);
or U14611 (N_14611,N_11040,N_12010);
nand U14612 (N_14612,N_11823,N_12151);
and U14613 (N_14613,N_9567,N_9625);
or U14614 (N_14614,N_10664,N_10584);
nor U14615 (N_14615,N_11738,N_11631);
or U14616 (N_14616,N_10221,N_10558);
or U14617 (N_14617,N_12292,N_10879);
nand U14618 (N_14618,N_12420,N_10888);
xor U14619 (N_14619,N_9773,N_10497);
xor U14620 (N_14620,N_10469,N_10198);
or U14621 (N_14621,N_11672,N_12490);
or U14622 (N_14622,N_11851,N_9799);
nor U14623 (N_14623,N_9503,N_9468);
nand U14624 (N_14624,N_9595,N_11083);
and U14625 (N_14625,N_10855,N_10858);
or U14626 (N_14626,N_10200,N_11564);
xor U14627 (N_14627,N_11922,N_9873);
nand U14628 (N_14628,N_11148,N_12029);
or U14629 (N_14629,N_11556,N_11854);
nor U14630 (N_14630,N_10922,N_9721);
or U14631 (N_14631,N_10307,N_12459);
and U14632 (N_14632,N_9737,N_9575);
nand U14633 (N_14633,N_10403,N_10686);
nor U14634 (N_14634,N_10449,N_9971);
xor U14635 (N_14635,N_11008,N_10499);
nor U14636 (N_14636,N_9803,N_11704);
and U14637 (N_14637,N_9936,N_12302);
nand U14638 (N_14638,N_12161,N_9686);
and U14639 (N_14639,N_9708,N_10532);
and U14640 (N_14640,N_9690,N_12422);
or U14641 (N_14641,N_12245,N_9685);
and U14642 (N_14642,N_10524,N_12344);
and U14643 (N_14643,N_11902,N_10612);
or U14644 (N_14644,N_12460,N_12432);
nand U14645 (N_14645,N_11620,N_11309);
xor U14646 (N_14646,N_10461,N_9480);
and U14647 (N_14647,N_10619,N_11566);
or U14648 (N_14648,N_9857,N_12270);
or U14649 (N_14649,N_11493,N_10083);
and U14650 (N_14650,N_11378,N_10037);
or U14651 (N_14651,N_12041,N_9911);
or U14652 (N_14652,N_9828,N_12049);
nor U14653 (N_14653,N_10282,N_10769);
or U14654 (N_14654,N_11043,N_11757);
nor U14655 (N_14655,N_12190,N_10999);
nor U14656 (N_14656,N_9955,N_11948);
or U14657 (N_14657,N_11043,N_10559);
and U14658 (N_14658,N_10636,N_9667);
nor U14659 (N_14659,N_11629,N_11093);
nand U14660 (N_14660,N_11754,N_11786);
nor U14661 (N_14661,N_12176,N_10236);
nor U14662 (N_14662,N_12132,N_10416);
nor U14663 (N_14663,N_12436,N_11709);
xnor U14664 (N_14664,N_12263,N_9852);
or U14665 (N_14665,N_11790,N_9924);
nand U14666 (N_14666,N_10119,N_12437);
or U14667 (N_14667,N_9633,N_10477);
nor U14668 (N_14668,N_10514,N_9469);
or U14669 (N_14669,N_12054,N_10063);
and U14670 (N_14670,N_11844,N_12314);
nand U14671 (N_14671,N_12411,N_12116);
nand U14672 (N_14672,N_10823,N_10543);
nand U14673 (N_14673,N_10648,N_11807);
xor U14674 (N_14674,N_11937,N_9700);
and U14675 (N_14675,N_12459,N_9878);
or U14676 (N_14676,N_10088,N_11503);
nor U14677 (N_14677,N_10029,N_10302);
or U14678 (N_14678,N_12388,N_10712);
nand U14679 (N_14679,N_11115,N_11876);
and U14680 (N_14680,N_11999,N_9503);
nand U14681 (N_14681,N_12186,N_9821);
nand U14682 (N_14682,N_10985,N_9513);
nand U14683 (N_14683,N_9860,N_9830);
nand U14684 (N_14684,N_11566,N_10269);
and U14685 (N_14685,N_11288,N_11474);
xnor U14686 (N_14686,N_12347,N_12418);
and U14687 (N_14687,N_10803,N_10576);
or U14688 (N_14688,N_12324,N_10857);
or U14689 (N_14689,N_12207,N_10161);
and U14690 (N_14690,N_10277,N_10718);
and U14691 (N_14691,N_11275,N_11403);
or U14692 (N_14692,N_12282,N_9496);
or U14693 (N_14693,N_10226,N_12150);
or U14694 (N_14694,N_11392,N_11049);
or U14695 (N_14695,N_10472,N_10134);
nand U14696 (N_14696,N_11950,N_10055);
nor U14697 (N_14697,N_10596,N_11567);
nand U14698 (N_14698,N_12090,N_11381);
nand U14699 (N_14699,N_11312,N_10118);
or U14700 (N_14700,N_11134,N_12391);
nor U14701 (N_14701,N_11789,N_11882);
xor U14702 (N_14702,N_11064,N_10999);
xor U14703 (N_14703,N_11548,N_9891);
and U14704 (N_14704,N_10275,N_10429);
or U14705 (N_14705,N_12381,N_9600);
nand U14706 (N_14706,N_11769,N_11368);
or U14707 (N_14707,N_10512,N_9436);
or U14708 (N_14708,N_11152,N_10712);
nand U14709 (N_14709,N_11056,N_12012);
and U14710 (N_14710,N_10753,N_10870);
or U14711 (N_14711,N_11621,N_10081);
nor U14712 (N_14712,N_10667,N_11061);
nor U14713 (N_14713,N_9904,N_12434);
and U14714 (N_14714,N_11264,N_9805);
xnor U14715 (N_14715,N_10916,N_11158);
or U14716 (N_14716,N_12146,N_9465);
nand U14717 (N_14717,N_10272,N_9476);
or U14718 (N_14718,N_9547,N_10119);
nor U14719 (N_14719,N_10580,N_10955);
nand U14720 (N_14720,N_10604,N_9980);
or U14721 (N_14721,N_10373,N_9399);
xor U14722 (N_14722,N_12451,N_9600);
nand U14723 (N_14723,N_12357,N_11743);
and U14724 (N_14724,N_11671,N_11600);
xor U14725 (N_14725,N_9968,N_12310);
nor U14726 (N_14726,N_10765,N_9950);
nand U14727 (N_14727,N_12008,N_12217);
xnor U14728 (N_14728,N_12288,N_10812);
nand U14729 (N_14729,N_10811,N_12172);
nor U14730 (N_14730,N_10736,N_11687);
xor U14731 (N_14731,N_10761,N_12193);
xor U14732 (N_14732,N_9491,N_10595);
and U14733 (N_14733,N_9993,N_10272);
xnor U14734 (N_14734,N_11243,N_11644);
nand U14735 (N_14735,N_11674,N_11103);
nand U14736 (N_14736,N_11567,N_11924);
nor U14737 (N_14737,N_11043,N_10123);
or U14738 (N_14738,N_9730,N_10331);
or U14739 (N_14739,N_12101,N_11874);
nor U14740 (N_14740,N_11648,N_10276);
or U14741 (N_14741,N_10187,N_9648);
nor U14742 (N_14742,N_11983,N_11652);
nor U14743 (N_14743,N_11054,N_10125);
nand U14744 (N_14744,N_9434,N_10374);
nand U14745 (N_14745,N_11617,N_9958);
or U14746 (N_14746,N_11564,N_12361);
nand U14747 (N_14747,N_11418,N_12268);
or U14748 (N_14748,N_11205,N_11410);
or U14749 (N_14749,N_9547,N_9965);
and U14750 (N_14750,N_10449,N_11008);
and U14751 (N_14751,N_12060,N_11824);
nand U14752 (N_14752,N_9893,N_11838);
nand U14753 (N_14753,N_9495,N_12097);
nand U14754 (N_14754,N_9877,N_10382);
and U14755 (N_14755,N_11514,N_12376);
or U14756 (N_14756,N_10361,N_12479);
xor U14757 (N_14757,N_12037,N_10575);
nor U14758 (N_14758,N_12278,N_11287);
or U14759 (N_14759,N_9918,N_11532);
and U14760 (N_14760,N_12191,N_11675);
nand U14761 (N_14761,N_10376,N_9645);
or U14762 (N_14762,N_9674,N_11258);
nand U14763 (N_14763,N_11886,N_10743);
or U14764 (N_14764,N_12101,N_9596);
nor U14765 (N_14765,N_9745,N_11030);
xnor U14766 (N_14766,N_9674,N_10305);
or U14767 (N_14767,N_9590,N_12414);
or U14768 (N_14768,N_10742,N_9867);
nand U14769 (N_14769,N_11235,N_11511);
nand U14770 (N_14770,N_10118,N_9923);
nand U14771 (N_14771,N_11676,N_10242);
nor U14772 (N_14772,N_11800,N_9676);
nor U14773 (N_14773,N_12168,N_10191);
nand U14774 (N_14774,N_10050,N_10287);
and U14775 (N_14775,N_10570,N_12068);
nor U14776 (N_14776,N_10171,N_10307);
nor U14777 (N_14777,N_10395,N_11898);
and U14778 (N_14778,N_11360,N_11297);
xnor U14779 (N_14779,N_10376,N_11251);
xnor U14780 (N_14780,N_10492,N_11070);
and U14781 (N_14781,N_10268,N_12043);
and U14782 (N_14782,N_11495,N_9478);
nor U14783 (N_14783,N_9990,N_9402);
and U14784 (N_14784,N_10380,N_9673);
and U14785 (N_14785,N_11457,N_12285);
and U14786 (N_14786,N_11773,N_11658);
and U14787 (N_14787,N_9424,N_10409);
or U14788 (N_14788,N_11746,N_9517);
nand U14789 (N_14789,N_11173,N_10127);
or U14790 (N_14790,N_9742,N_9801);
nor U14791 (N_14791,N_12091,N_9766);
and U14792 (N_14792,N_10819,N_10281);
or U14793 (N_14793,N_11023,N_11898);
nor U14794 (N_14794,N_11563,N_12182);
nor U14795 (N_14795,N_12089,N_10481);
and U14796 (N_14796,N_9412,N_10817);
or U14797 (N_14797,N_12192,N_10585);
nor U14798 (N_14798,N_11252,N_11970);
or U14799 (N_14799,N_11852,N_11433);
or U14800 (N_14800,N_11284,N_10492);
or U14801 (N_14801,N_11355,N_11733);
nand U14802 (N_14802,N_11477,N_12144);
or U14803 (N_14803,N_11521,N_11459);
nor U14804 (N_14804,N_10511,N_11432);
nor U14805 (N_14805,N_11699,N_10052);
nand U14806 (N_14806,N_11055,N_11698);
nand U14807 (N_14807,N_10505,N_10646);
and U14808 (N_14808,N_9452,N_9705);
and U14809 (N_14809,N_9501,N_11537);
and U14810 (N_14810,N_10832,N_12095);
or U14811 (N_14811,N_10015,N_11916);
and U14812 (N_14812,N_11092,N_12230);
nor U14813 (N_14813,N_11555,N_11843);
nand U14814 (N_14814,N_9389,N_11094);
nor U14815 (N_14815,N_10568,N_10454);
and U14816 (N_14816,N_9540,N_10438);
and U14817 (N_14817,N_10106,N_10194);
nand U14818 (N_14818,N_12169,N_11386);
nand U14819 (N_14819,N_10743,N_10323);
nor U14820 (N_14820,N_10544,N_11338);
and U14821 (N_14821,N_12348,N_11153);
and U14822 (N_14822,N_10465,N_9951);
xor U14823 (N_14823,N_9609,N_11435);
nor U14824 (N_14824,N_10125,N_12233);
and U14825 (N_14825,N_10093,N_9866);
or U14826 (N_14826,N_11559,N_10494);
nand U14827 (N_14827,N_9835,N_11179);
and U14828 (N_14828,N_9963,N_11602);
nor U14829 (N_14829,N_12418,N_9810);
xor U14830 (N_14830,N_11291,N_10894);
nand U14831 (N_14831,N_11358,N_10309);
and U14832 (N_14832,N_11664,N_9400);
nand U14833 (N_14833,N_9726,N_9414);
or U14834 (N_14834,N_12436,N_10342);
nor U14835 (N_14835,N_9857,N_11553);
or U14836 (N_14836,N_10558,N_11971);
nand U14837 (N_14837,N_11278,N_11468);
nand U14838 (N_14838,N_12337,N_12154);
and U14839 (N_14839,N_11206,N_10297);
nand U14840 (N_14840,N_12429,N_11307);
and U14841 (N_14841,N_11774,N_11720);
nor U14842 (N_14842,N_10968,N_11062);
nor U14843 (N_14843,N_9647,N_11638);
and U14844 (N_14844,N_10570,N_9486);
or U14845 (N_14845,N_9683,N_12473);
and U14846 (N_14846,N_10618,N_11527);
or U14847 (N_14847,N_9681,N_10172);
nor U14848 (N_14848,N_10443,N_12009);
nor U14849 (N_14849,N_11507,N_11811);
or U14850 (N_14850,N_10583,N_9826);
nor U14851 (N_14851,N_12432,N_10731);
nor U14852 (N_14852,N_9839,N_11210);
nor U14853 (N_14853,N_9386,N_11633);
or U14854 (N_14854,N_10575,N_9777);
and U14855 (N_14855,N_10230,N_9875);
nand U14856 (N_14856,N_12177,N_10274);
nand U14857 (N_14857,N_9555,N_10227);
nand U14858 (N_14858,N_9885,N_11130);
nor U14859 (N_14859,N_12416,N_10548);
nand U14860 (N_14860,N_9786,N_9812);
nand U14861 (N_14861,N_10937,N_11287);
and U14862 (N_14862,N_9934,N_10119);
nand U14863 (N_14863,N_10042,N_12435);
and U14864 (N_14864,N_12410,N_9724);
nor U14865 (N_14865,N_10193,N_10209);
nor U14866 (N_14866,N_12314,N_12228);
or U14867 (N_14867,N_10953,N_11674);
nand U14868 (N_14868,N_12227,N_11387);
and U14869 (N_14869,N_12332,N_11376);
nand U14870 (N_14870,N_9838,N_11895);
nor U14871 (N_14871,N_9443,N_9577);
nand U14872 (N_14872,N_9926,N_10108);
nand U14873 (N_14873,N_10420,N_9601);
xor U14874 (N_14874,N_10843,N_12138);
or U14875 (N_14875,N_11264,N_12499);
and U14876 (N_14876,N_12085,N_11767);
nor U14877 (N_14877,N_11793,N_10548);
or U14878 (N_14878,N_10410,N_10210);
or U14879 (N_14879,N_10277,N_11414);
and U14880 (N_14880,N_12232,N_9550);
and U14881 (N_14881,N_12383,N_10140);
nand U14882 (N_14882,N_9432,N_12025);
nor U14883 (N_14883,N_10218,N_9664);
nor U14884 (N_14884,N_10113,N_11465);
xnor U14885 (N_14885,N_10265,N_9518);
nor U14886 (N_14886,N_10993,N_11342);
and U14887 (N_14887,N_12036,N_10583);
xnor U14888 (N_14888,N_11285,N_10436);
or U14889 (N_14889,N_11243,N_12270);
nor U14890 (N_14890,N_9933,N_9927);
nor U14891 (N_14891,N_10433,N_9713);
xnor U14892 (N_14892,N_12301,N_10971);
or U14893 (N_14893,N_11049,N_9590);
and U14894 (N_14894,N_10997,N_11889);
and U14895 (N_14895,N_10035,N_9541);
nor U14896 (N_14896,N_11440,N_12155);
nand U14897 (N_14897,N_10492,N_12460);
nor U14898 (N_14898,N_10633,N_11993);
and U14899 (N_14899,N_12301,N_9756);
nand U14900 (N_14900,N_9795,N_11076);
nand U14901 (N_14901,N_10280,N_11641);
or U14902 (N_14902,N_10181,N_11619);
nor U14903 (N_14903,N_9539,N_9471);
nor U14904 (N_14904,N_10096,N_9486);
or U14905 (N_14905,N_9452,N_9831);
or U14906 (N_14906,N_9729,N_9893);
or U14907 (N_14907,N_10012,N_11093);
and U14908 (N_14908,N_11800,N_11721);
nor U14909 (N_14909,N_9662,N_12142);
xor U14910 (N_14910,N_12404,N_9476);
xor U14911 (N_14911,N_9786,N_10163);
or U14912 (N_14912,N_12001,N_10051);
and U14913 (N_14913,N_11817,N_11129);
nor U14914 (N_14914,N_12277,N_9388);
xnor U14915 (N_14915,N_11483,N_11714);
nor U14916 (N_14916,N_10692,N_12447);
or U14917 (N_14917,N_10139,N_10272);
and U14918 (N_14918,N_9960,N_10111);
nor U14919 (N_14919,N_12373,N_11807);
nand U14920 (N_14920,N_12489,N_11338);
or U14921 (N_14921,N_9415,N_11459);
nor U14922 (N_14922,N_12100,N_11812);
and U14923 (N_14923,N_11138,N_10748);
and U14924 (N_14924,N_11973,N_12090);
and U14925 (N_14925,N_10774,N_11790);
nand U14926 (N_14926,N_11832,N_11117);
nand U14927 (N_14927,N_9879,N_10723);
and U14928 (N_14928,N_9778,N_9473);
or U14929 (N_14929,N_11139,N_10807);
and U14930 (N_14930,N_10151,N_11595);
nand U14931 (N_14931,N_11729,N_10109);
xor U14932 (N_14932,N_10638,N_11721);
or U14933 (N_14933,N_9557,N_11010);
nand U14934 (N_14934,N_10999,N_11621);
or U14935 (N_14935,N_10033,N_11410);
nor U14936 (N_14936,N_9505,N_11150);
or U14937 (N_14937,N_10706,N_9490);
nor U14938 (N_14938,N_10067,N_12444);
or U14939 (N_14939,N_11355,N_12031);
and U14940 (N_14940,N_9389,N_9990);
and U14941 (N_14941,N_9788,N_12458);
nor U14942 (N_14942,N_10478,N_9480);
nand U14943 (N_14943,N_12228,N_12191);
nand U14944 (N_14944,N_10132,N_12043);
nor U14945 (N_14945,N_10281,N_9997);
nand U14946 (N_14946,N_11928,N_10331);
xnor U14947 (N_14947,N_11834,N_12284);
or U14948 (N_14948,N_12206,N_9783);
nor U14949 (N_14949,N_10638,N_10310);
or U14950 (N_14950,N_10256,N_9528);
or U14951 (N_14951,N_10746,N_11356);
nand U14952 (N_14952,N_11191,N_10051);
or U14953 (N_14953,N_10781,N_10847);
nor U14954 (N_14954,N_12049,N_12452);
and U14955 (N_14955,N_11505,N_9837);
nand U14956 (N_14956,N_11007,N_10628);
and U14957 (N_14957,N_11886,N_10838);
and U14958 (N_14958,N_9738,N_12067);
xor U14959 (N_14959,N_11988,N_11100);
nor U14960 (N_14960,N_12111,N_12157);
or U14961 (N_14961,N_11220,N_9475);
and U14962 (N_14962,N_10577,N_9998);
nor U14963 (N_14963,N_9673,N_11501);
nor U14964 (N_14964,N_9667,N_12385);
or U14965 (N_14965,N_9480,N_11946);
nand U14966 (N_14966,N_11189,N_12205);
nor U14967 (N_14967,N_9767,N_10530);
nor U14968 (N_14968,N_10867,N_11372);
nor U14969 (N_14969,N_10227,N_10752);
nand U14970 (N_14970,N_12103,N_11765);
xnor U14971 (N_14971,N_10225,N_9939);
xor U14972 (N_14972,N_12243,N_10411);
nand U14973 (N_14973,N_11335,N_12464);
or U14974 (N_14974,N_11613,N_12360);
nor U14975 (N_14975,N_11429,N_10352);
nor U14976 (N_14976,N_11161,N_11622);
nor U14977 (N_14977,N_10245,N_10622);
nand U14978 (N_14978,N_9430,N_11377);
nor U14979 (N_14979,N_10841,N_11080);
nand U14980 (N_14980,N_10037,N_11879);
and U14981 (N_14981,N_10682,N_9795);
and U14982 (N_14982,N_9680,N_10593);
or U14983 (N_14983,N_11603,N_9674);
or U14984 (N_14984,N_11030,N_10003);
nor U14985 (N_14985,N_11717,N_12250);
nand U14986 (N_14986,N_11847,N_9525);
nand U14987 (N_14987,N_12189,N_12229);
or U14988 (N_14988,N_11625,N_12032);
xnor U14989 (N_14989,N_11462,N_10888);
and U14990 (N_14990,N_11518,N_9734);
or U14991 (N_14991,N_11396,N_10038);
nand U14992 (N_14992,N_11608,N_10296);
or U14993 (N_14993,N_12347,N_9741);
and U14994 (N_14994,N_11260,N_12330);
nor U14995 (N_14995,N_9618,N_11993);
nand U14996 (N_14996,N_11856,N_12460);
nor U14997 (N_14997,N_9905,N_10572);
nand U14998 (N_14998,N_9859,N_12268);
nand U14999 (N_14999,N_9875,N_11881);
nor U15000 (N_15000,N_10012,N_9598);
and U15001 (N_15001,N_9588,N_10574);
nand U15002 (N_15002,N_10876,N_9414);
or U15003 (N_15003,N_11573,N_12336);
and U15004 (N_15004,N_11545,N_12077);
and U15005 (N_15005,N_12206,N_9420);
or U15006 (N_15006,N_9875,N_10100);
or U15007 (N_15007,N_11369,N_10165);
and U15008 (N_15008,N_11961,N_9956);
and U15009 (N_15009,N_11906,N_12375);
xor U15010 (N_15010,N_11331,N_10544);
nor U15011 (N_15011,N_9731,N_11723);
xor U15012 (N_15012,N_9512,N_11986);
nor U15013 (N_15013,N_11384,N_9511);
and U15014 (N_15014,N_11952,N_11638);
or U15015 (N_15015,N_10531,N_12378);
nand U15016 (N_15016,N_9621,N_9650);
nor U15017 (N_15017,N_10234,N_10222);
nand U15018 (N_15018,N_10130,N_12228);
or U15019 (N_15019,N_11255,N_12263);
nand U15020 (N_15020,N_11157,N_12320);
and U15021 (N_15021,N_10604,N_12178);
or U15022 (N_15022,N_9543,N_11859);
xor U15023 (N_15023,N_12210,N_12356);
or U15024 (N_15024,N_10142,N_10305);
nand U15025 (N_15025,N_9497,N_10563);
xor U15026 (N_15026,N_11034,N_10656);
nor U15027 (N_15027,N_10532,N_11642);
or U15028 (N_15028,N_10088,N_11913);
and U15029 (N_15029,N_12153,N_10798);
xnor U15030 (N_15030,N_10145,N_10436);
and U15031 (N_15031,N_11382,N_10216);
or U15032 (N_15032,N_10394,N_11201);
or U15033 (N_15033,N_11495,N_11955);
and U15034 (N_15034,N_10316,N_11780);
nor U15035 (N_15035,N_10698,N_11799);
or U15036 (N_15036,N_10035,N_10448);
nor U15037 (N_15037,N_10474,N_10203);
nor U15038 (N_15038,N_9887,N_9389);
nand U15039 (N_15039,N_9791,N_12469);
nor U15040 (N_15040,N_11583,N_9968);
or U15041 (N_15041,N_9526,N_11585);
or U15042 (N_15042,N_11455,N_10686);
and U15043 (N_15043,N_10369,N_11554);
and U15044 (N_15044,N_10593,N_9903);
nor U15045 (N_15045,N_11534,N_9631);
or U15046 (N_15046,N_11227,N_11989);
and U15047 (N_15047,N_10329,N_9846);
nand U15048 (N_15048,N_12033,N_10439);
nor U15049 (N_15049,N_12136,N_12458);
and U15050 (N_15050,N_10689,N_11177);
nor U15051 (N_15051,N_9840,N_9747);
and U15052 (N_15052,N_11311,N_9584);
or U15053 (N_15053,N_11762,N_10993);
nand U15054 (N_15054,N_10951,N_12317);
nand U15055 (N_15055,N_12291,N_9403);
nor U15056 (N_15056,N_9569,N_11848);
nor U15057 (N_15057,N_10772,N_10097);
nand U15058 (N_15058,N_11695,N_10055);
nand U15059 (N_15059,N_12179,N_9675);
xnor U15060 (N_15060,N_10875,N_10439);
nor U15061 (N_15061,N_10074,N_11162);
nand U15062 (N_15062,N_11629,N_10866);
or U15063 (N_15063,N_9870,N_10216);
nor U15064 (N_15064,N_10543,N_11647);
or U15065 (N_15065,N_12478,N_12031);
nand U15066 (N_15066,N_10708,N_10817);
or U15067 (N_15067,N_11620,N_12097);
or U15068 (N_15068,N_10741,N_12450);
and U15069 (N_15069,N_11652,N_11474);
and U15070 (N_15070,N_10473,N_11183);
xor U15071 (N_15071,N_11588,N_12128);
nor U15072 (N_15072,N_11280,N_10722);
xnor U15073 (N_15073,N_11553,N_9868);
nor U15074 (N_15074,N_12068,N_9666);
or U15075 (N_15075,N_10077,N_11163);
and U15076 (N_15076,N_9705,N_11250);
nor U15077 (N_15077,N_10049,N_10129);
or U15078 (N_15078,N_11612,N_12457);
or U15079 (N_15079,N_12005,N_10899);
nor U15080 (N_15080,N_11184,N_9486);
or U15081 (N_15081,N_10716,N_11742);
nor U15082 (N_15082,N_10780,N_11968);
nor U15083 (N_15083,N_12444,N_9823);
and U15084 (N_15084,N_12215,N_9442);
and U15085 (N_15085,N_11562,N_11035);
nand U15086 (N_15086,N_12361,N_12256);
nand U15087 (N_15087,N_9839,N_11730);
nor U15088 (N_15088,N_10454,N_9875);
xnor U15089 (N_15089,N_10355,N_10886);
nor U15090 (N_15090,N_11249,N_10301);
nand U15091 (N_15091,N_9389,N_11516);
nor U15092 (N_15092,N_9773,N_9524);
and U15093 (N_15093,N_11036,N_11608);
xor U15094 (N_15094,N_12451,N_11220);
nand U15095 (N_15095,N_9440,N_11781);
xor U15096 (N_15096,N_10955,N_12426);
nor U15097 (N_15097,N_9937,N_11880);
nor U15098 (N_15098,N_11287,N_12305);
xnor U15099 (N_15099,N_11390,N_10078);
and U15100 (N_15100,N_10025,N_10856);
and U15101 (N_15101,N_9570,N_11039);
and U15102 (N_15102,N_11144,N_12138);
nor U15103 (N_15103,N_9874,N_10098);
or U15104 (N_15104,N_11813,N_10338);
xnor U15105 (N_15105,N_11699,N_10344);
nor U15106 (N_15106,N_10712,N_10078);
xor U15107 (N_15107,N_10859,N_9847);
and U15108 (N_15108,N_11274,N_11987);
nand U15109 (N_15109,N_11726,N_10178);
nor U15110 (N_15110,N_10695,N_9870);
nor U15111 (N_15111,N_11376,N_10621);
nand U15112 (N_15112,N_10570,N_10324);
nand U15113 (N_15113,N_10440,N_11693);
nand U15114 (N_15114,N_11249,N_10103);
nand U15115 (N_15115,N_11878,N_11787);
or U15116 (N_15116,N_11444,N_10130);
nor U15117 (N_15117,N_10688,N_10241);
or U15118 (N_15118,N_10018,N_12170);
and U15119 (N_15119,N_10561,N_11836);
nand U15120 (N_15120,N_9839,N_9590);
xor U15121 (N_15121,N_9538,N_10207);
and U15122 (N_15122,N_12281,N_11440);
nand U15123 (N_15123,N_10267,N_9752);
or U15124 (N_15124,N_11469,N_12173);
and U15125 (N_15125,N_12431,N_11134);
nor U15126 (N_15126,N_9780,N_12348);
nor U15127 (N_15127,N_11636,N_10581);
or U15128 (N_15128,N_11649,N_12398);
and U15129 (N_15129,N_10460,N_10426);
nand U15130 (N_15130,N_10061,N_9765);
nand U15131 (N_15131,N_9475,N_11803);
nor U15132 (N_15132,N_12274,N_11671);
nand U15133 (N_15133,N_11997,N_12331);
nand U15134 (N_15134,N_9789,N_11264);
or U15135 (N_15135,N_10666,N_11543);
or U15136 (N_15136,N_12397,N_9426);
nor U15137 (N_15137,N_11082,N_9669);
nor U15138 (N_15138,N_11821,N_10529);
or U15139 (N_15139,N_11772,N_9388);
and U15140 (N_15140,N_11217,N_11293);
or U15141 (N_15141,N_10982,N_9953);
and U15142 (N_15142,N_10668,N_11280);
or U15143 (N_15143,N_12281,N_12044);
nand U15144 (N_15144,N_10435,N_11391);
and U15145 (N_15145,N_11683,N_10930);
and U15146 (N_15146,N_10234,N_10634);
nand U15147 (N_15147,N_11710,N_10760);
nor U15148 (N_15148,N_10941,N_10742);
nand U15149 (N_15149,N_11635,N_11487);
or U15150 (N_15150,N_9991,N_9781);
or U15151 (N_15151,N_11667,N_12448);
or U15152 (N_15152,N_9465,N_11697);
and U15153 (N_15153,N_9589,N_10298);
nor U15154 (N_15154,N_9763,N_11475);
nor U15155 (N_15155,N_10307,N_9643);
or U15156 (N_15156,N_12033,N_9386);
xor U15157 (N_15157,N_11941,N_11560);
or U15158 (N_15158,N_10054,N_10883);
nand U15159 (N_15159,N_10901,N_10476);
nor U15160 (N_15160,N_10751,N_9705);
nand U15161 (N_15161,N_10367,N_9929);
nand U15162 (N_15162,N_11483,N_10104);
nand U15163 (N_15163,N_12239,N_10610);
nor U15164 (N_15164,N_11065,N_11461);
and U15165 (N_15165,N_12007,N_11248);
or U15166 (N_15166,N_10474,N_10165);
or U15167 (N_15167,N_11941,N_9567);
and U15168 (N_15168,N_11585,N_12210);
nand U15169 (N_15169,N_10223,N_9574);
and U15170 (N_15170,N_10418,N_11622);
and U15171 (N_15171,N_11977,N_12252);
nor U15172 (N_15172,N_9815,N_12214);
or U15173 (N_15173,N_9390,N_11848);
and U15174 (N_15174,N_9746,N_12448);
nor U15175 (N_15175,N_9401,N_10393);
nor U15176 (N_15176,N_10893,N_10289);
nor U15177 (N_15177,N_10496,N_9839);
or U15178 (N_15178,N_12322,N_9404);
or U15179 (N_15179,N_10701,N_10366);
nor U15180 (N_15180,N_10822,N_11465);
and U15181 (N_15181,N_11809,N_11787);
xor U15182 (N_15182,N_11326,N_11565);
and U15183 (N_15183,N_11070,N_10857);
or U15184 (N_15184,N_11067,N_9420);
nand U15185 (N_15185,N_12301,N_9953);
nor U15186 (N_15186,N_12378,N_12191);
nand U15187 (N_15187,N_11264,N_9409);
or U15188 (N_15188,N_12126,N_10280);
nor U15189 (N_15189,N_11352,N_12130);
nor U15190 (N_15190,N_10249,N_12300);
and U15191 (N_15191,N_11968,N_10197);
or U15192 (N_15192,N_11957,N_11557);
nor U15193 (N_15193,N_11950,N_12061);
or U15194 (N_15194,N_10882,N_11147);
nand U15195 (N_15195,N_10151,N_9897);
nand U15196 (N_15196,N_9737,N_12413);
or U15197 (N_15197,N_11620,N_11518);
and U15198 (N_15198,N_10875,N_9507);
nand U15199 (N_15199,N_11826,N_10488);
and U15200 (N_15200,N_12261,N_11263);
and U15201 (N_15201,N_11554,N_10540);
nand U15202 (N_15202,N_10440,N_10868);
nand U15203 (N_15203,N_9434,N_11868);
and U15204 (N_15204,N_12304,N_10532);
and U15205 (N_15205,N_12187,N_11202);
and U15206 (N_15206,N_10893,N_12160);
nor U15207 (N_15207,N_10829,N_12063);
nor U15208 (N_15208,N_10672,N_10181);
and U15209 (N_15209,N_11050,N_10226);
xnor U15210 (N_15210,N_9965,N_10951);
or U15211 (N_15211,N_10186,N_9484);
nand U15212 (N_15212,N_9653,N_11419);
and U15213 (N_15213,N_11908,N_10537);
and U15214 (N_15214,N_9959,N_9976);
or U15215 (N_15215,N_12189,N_11604);
and U15216 (N_15216,N_10507,N_11177);
nor U15217 (N_15217,N_9595,N_9884);
or U15218 (N_15218,N_9609,N_12119);
nor U15219 (N_15219,N_10619,N_10806);
or U15220 (N_15220,N_12242,N_9866);
nor U15221 (N_15221,N_10046,N_12210);
nor U15222 (N_15222,N_11936,N_11784);
and U15223 (N_15223,N_11859,N_12054);
xnor U15224 (N_15224,N_10460,N_11883);
and U15225 (N_15225,N_11359,N_9546);
and U15226 (N_15226,N_10557,N_11243);
nand U15227 (N_15227,N_11083,N_12075);
nor U15228 (N_15228,N_10178,N_11488);
nor U15229 (N_15229,N_11815,N_11405);
and U15230 (N_15230,N_11492,N_9780);
nand U15231 (N_15231,N_9908,N_12405);
nor U15232 (N_15232,N_10545,N_10823);
and U15233 (N_15233,N_9487,N_10916);
and U15234 (N_15234,N_10483,N_10731);
or U15235 (N_15235,N_9461,N_10876);
nand U15236 (N_15236,N_9381,N_10361);
or U15237 (N_15237,N_10469,N_12457);
nand U15238 (N_15238,N_10688,N_11194);
xor U15239 (N_15239,N_12197,N_12370);
and U15240 (N_15240,N_10815,N_11223);
and U15241 (N_15241,N_9613,N_10754);
nor U15242 (N_15242,N_12447,N_10602);
nor U15243 (N_15243,N_10018,N_9480);
and U15244 (N_15244,N_10742,N_12057);
xor U15245 (N_15245,N_10169,N_11194);
nand U15246 (N_15246,N_12443,N_11634);
xor U15247 (N_15247,N_12389,N_11395);
and U15248 (N_15248,N_10835,N_12408);
or U15249 (N_15249,N_12174,N_12404);
or U15250 (N_15250,N_10407,N_9417);
or U15251 (N_15251,N_11499,N_10404);
nand U15252 (N_15252,N_11485,N_11893);
or U15253 (N_15253,N_12377,N_10070);
nand U15254 (N_15254,N_11352,N_11999);
nand U15255 (N_15255,N_10758,N_11337);
nand U15256 (N_15256,N_10130,N_9462);
and U15257 (N_15257,N_11876,N_10024);
nand U15258 (N_15258,N_10999,N_9426);
xor U15259 (N_15259,N_11832,N_9725);
or U15260 (N_15260,N_11421,N_10971);
and U15261 (N_15261,N_11138,N_11786);
nor U15262 (N_15262,N_12130,N_9828);
nand U15263 (N_15263,N_11521,N_12247);
or U15264 (N_15264,N_10554,N_12119);
nand U15265 (N_15265,N_12385,N_11313);
or U15266 (N_15266,N_10435,N_10346);
nand U15267 (N_15267,N_11769,N_10885);
or U15268 (N_15268,N_10591,N_11544);
and U15269 (N_15269,N_10450,N_10076);
nand U15270 (N_15270,N_12299,N_9843);
nand U15271 (N_15271,N_10904,N_9876);
and U15272 (N_15272,N_11535,N_10525);
or U15273 (N_15273,N_12010,N_11654);
and U15274 (N_15274,N_11086,N_11612);
nor U15275 (N_15275,N_9549,N_10670);
and U15276 (N_15276,N_11877,N_10580);
xor U15277 (N_15277,N_9947,N_11594);
or U15278 (N_15278,N_9995,N_10995);
nor U15279 (N_15279,N_10988,N_10175);
and U15280 (N_15280,N_11782,N_10439);
or U15281 (N_15281,N_11947,N_11142);
or U15282 (N_15282,N_9688,N_11635);
nand U15283 (N_15283,N_11193,N_9391);
or U15284 (N_15284,N_9416,N_12359);
nor U15285 (N_15285,N_11682,N_9770);
nand U15286 (N_15286,N_10385,N_10080);
nor U15287 (N_15287,N_9962,N_10662);
nor U15288 (N_15288,N_10974,N_10851);
nand U15289 (N_15289,N_12251,N_9926);
nor U15290 (N_15290,N_11476,N_11880);
nand U15291 (N_15291,N_11247,N_10203);
and U15292 (N_15292,N_12315,N_12082);
xnor U15293 (N_15293,N_10721,N_12087);
and U15294 (N_15294,N_9931,N_12422);
nand U15295 (N_15295,N_12161,N_10471);
or U15296 (N_15296,N_9718,N_11465);
nand U15297 (N_15297,N_10699,N_9828);
nor U15298 (N_15298,N_10627,N_10928);
or U15299 (N_15299,N_9538,N_11156);
or U15300 (N_15300,N_11044,N_10927);
nor U15301 (N_15301,N_10351,N_10089);
or U15302 (N_15302,N_9534,N_12379);
nand U15303 (N_15303,N_12051,N_9525);
and U15304 (N_15304,N_12380,N_12383);
or U15305 (N_15305,N_11322,N_10622);
nor U15306 (N_15306,N_9687,N_11312);
and U15307 (N_15307,N_9993,N_10051);
or U15308 (N_15308,N_11093,N_11030);
nor U15309 (N_15309,N_9778,N_11843);
nand U15310 (N_15310,N_11740,N_10943);
nor U15311 (N_15311,N_10619,N_11200);
nor U15312 (N_15312,N_10787,N_10241);
and U15313 (N_15313,N_9545,N_9432);
or U15314 (N_15314,N_10369,N_11855);
nand U15315 (N_15315,N_11794,N_12012);
nor U15316 (N_15316,N_10846,N_12372);
nand U15317 (N_15317,N_10836,N_11933);
nand U15318 (N_15318,N_12049,N_12305);
nor U15319 (N_15319,N_12005,N_11493);
or U15320 (N_15320,N_9433,N_11074);
and U15321 (N_15321,N_11839,N_11192);
and U15322 (N_15322,N_10807,N_10432);
or U15323 (N_15323,N_10987,N_10514);
nand U15324 (N_15324,N_10543,N_10155);
nand U15325 (N_15325,N_11199,N_12007);
nand U15326 (N_15326,N_11792,N_11366);
or U15327 (N_15327,N_12124,N_12407);
and U15328 (N_15328,N_11360,N_11073);
or U15329 (N_15329,N_12441,N_11238);
nor U15330 (N_15330,N_12155,N_11531);
nand U15331 (N_15331,N_10208,N_11198);
and U15332 (N_15332,N_11312,N_10715);
nor U15333 (N_15333,N_10647,N_10607);
nand U15334 (N_15334,N_10183,N_10495);
and U15335 (N_15335,N_11184,N_11427);
or U15336 (N_15336,N_11078,N_11206);
or U15337 (N_15337,N_12113,N_9878);
or U15338 (N_15338,N_11268,N_9985);
xor U15339 (N_15339,N_12024,N_9380);
nand U15340 (N_15340,N_11225,N_11503);
or U15341 (N_15341,N_10292,N_10513);
or U15342 (N_15342,N_11104,N_11977);
and U15343 (N_15343,N_11863,N_11890);
or U15344 (N_15344,N_12423,N_11602);
or U15345 (N_15345,N_10287,N_10624);
nand U15346 (N_15346,N_9455,N_12447);
and U15347 (N_15347,N_10870,N_11996);
nand U15348 (N_15348,N_10045,N_11240);
nor U15349 (N_15349,N_10693,N_11753);
nor U15350 (N_15350,N_10389,N_9699);
nor U15351 (N_15351,N_11221,N_10808);
nand U15352 (N_15352,N_11911,N_12274);
or U15353 (N_15353,N_12104,N_9696);
and U15354 (N_15354,N_11618,N_10150);
or U15355 (N_15355,N_11125,N_11022);
or U15356 (N_15356,N_10984,N_11847);
xor U15357 (N_15357,N_9776,N_10559);
nand U15358 (N_15358,N_10012,N_12028);
nand U15359 (N_15359,N_12151,N_9488);
nand U15360 (N_15360,N_11175,N_9807);
nand U15361 (N_15361,N_10129,N_9461);
xor U15362 (N_15362,N_11289,N_11353);
nand U15363 (N_15363,N_12280,N_12241);
nand U15364 (N_15364,N_11444,N_11789);
or U15365 (N_15365,N_11825,N_9576);
nand U15366 (N_15366,N_9484,N_12388);
nand U15367 (N_15367,N_11822,N_11439);
xor U15368 (N_15368,N_10165,N_9839);
and U15369 (N_15369,N_11574,N_12115);
nor U15370 (N_15370,N_9912,N_11352);
or U15371 (N_15371,N_9752,N_10871);
or U15372 (N_15372,N_10692,N_11001);
nor U15373 (N_15373,N_10189,N_10463);
nor U15374 (N_15374,N_9684,N_10689);
nand U15375 (N_15375,N_10663,N_10276);
or U15376 (N_15376,N_9995,N_10218);
nor U15377 (N_15377,N_12469,N_11235);
and U15378 (N_15378,N_10176,N_11033);
nor U15379 (N_15379,N_11148,N_10190);
xnor U15380 (N_15380,N_11034,N_11688);
nor U15381 (N_15381,N_9586,N_11038);
nor U15382 (N_15382,N_12458,N_12449);
or U15383 (N_15383,N_12389,N_9937);
nor U15384 (N_15384,N_12370,N_10949);
nor U15385 (N_15385,N_11634,N_9602);
nand U15386 (N_15386,N_9684,N_9813);
or U15387 (N_15387,N_12242,N_10070);
nor U15388 (N_15388,N_11562,N_11801);
nor U15389 (N_15389,N_11053,N_9687);
or U15390 (N_15390,N_11076,N_12150);
or U15391 (N_15391,N_11319,N_10193);
nand U15392 (N_15392,N_9400,N_9427);
nor U15393 (N_15393,N_10905,N_10853);
nand U15394 (N_15394,N_10293,N_12101);
nand U15395 (N_15395,N_10030,N_10958);
and U15396 (N_15396,N_9913,N_9438);
xor U15397 (N_15397,N_9483,N_11976);
nand U15398 (N_15398,N_12293,N_11120);
nand U15399 (N_15399,N_10714,N_11507);
and U15400 (N_15400,N_11732,N_10967);
or U15401 (N_15401,N_10149,N_12073);
or U15402 (N_15402,N_10115,N_11566);
and U15403 (N_15403,N_10901,N_10003);
nor U15404 (N_15404,N_12027,N_10290);
nand U15405 (N_15405,N_11411,N_9801);
nor U15406 (N_15406,N_9520,N_10945);
or U15407 (N_15407,N_10100,N_9783);
and U15408 (N_15408,N_9986,N_10896);
nand U15409 (N_15409,N_10269,N_10315);
or U15410 (N_15410,N_12291,N_11732);
xor U15411 (N_15411,N_10990,N_11541);
nand U15412 (N_15412,N_11401,N_11422);
or U15413 (N_15413,N_9998,N_11287);
and U15414 (N_15414,N_10975,N_11663);
and U15415 (N_15415,N_11514,N_10064);
nand U15416 (N_15416,N_11938,N_9612);
and U15417 (N_15417,N_11710,N_11760);
xnor U15418 (N_15418,N_11282,N_12343);
and U15419 (N_15419,N_9526,N_9575);
nand U15420 (N_15420,N_10214,N_10454);
nand U15421 (N_15421,N_12415,N_12144);
xnor U15422 (N_15422,N_11759,N_11408);
xor U15423 (N_15423,N_10079,N_10094);
nand U15424 (N_15424,N_11087,N_11813);
nor U15425 (N_15425,N_9433,N_10058);
xnor U15426 (N_15426,N_11730,N_11585);
and U15427 (N_15427,N_11328,N_10352);
nor U15428 (N_15428,N_11893,N_11262);
nand U15429 (N_15429,N_10997,N_10164);
and U15430 (N_15430,N_11698,N_11548);
nand U15431 (N_15431,N_10911,N_11284);
and U15432 (N_15432,N_11929,N_12102);
and U15433 (N_15433,N_11069,N_11468);
nor U15434 (N_15434,N_12443,N_10121);
xor U15435 (N_15435,N_12435,N_11341);
nand U15436 (N_15436,N_11451,N_10950);
nand U15437 (N_15437,N_12190,N_10106);
and U15438 (N_15438,N_12254,N_11053);
nor U15439 (N_15439,N_11044,N_10010);
or U15440 (N_15440,N_12407,N_10234);
and U15441 (N_15441,N_11132,N_10369);
nand U15442 (N_15442,N_9945,N_10572);
and U15443 (N_15443,N_10880,N_12297);
xor U15444 (N_15444,N_11852,N_10212);
or U15445 (N_15445,N_10526,N_10444);
nand U15446 (N_15446,N_11037,N_9483);
and U15447 (N_15447,N_9418,N_10807);
or U15448 (N_15448,N_12077,N_10258);
nand U15449 (N_15449,N_11674,N_11844);
and U15450 (N_15450,N_10101,N_10444);
or U15451 (N_15451,N_10048,N_12272);
and U15452 (N_15452,N_10569,N_11337);
and U15453 (N_15453,N_9788,N_11414);
and U15454 (N_15454,N_10435,N_11818);
nor U15455 (N_15455,N_9959,N_11260);
and U15456 (N_15456,N_11480,N_10713);
xnor U15457 (N_15457,N_11801,N_10247);
nand U15458 (N_15458,N_10785,N_11480);
nand U15459 (N_15459,N_12390,N_10282);
and U15460 (N_15460,N_12084,N_11208);
and U15461 (N_15461,N_10384,N_11607);
and U15462 (N_15462,N_11159,N_10239);
nand U15463 (N_15463,N_11062,N_12371);
nor U15464 (N_15464,N_11560,N_10733);
or U15465 (N_15465,N_9844,N_11225);
and U15466 (N_15466,N_11845,N_10513);
nand U15467 (N_15467,N_11140,N_9764);
and U15468 (N_15468,N_12190,N_10691);
nand U15469 (N_15469,N_10955,N_9814);
and U15470 (N_15470,N_12429,N_10801);
nor U15471 (N_15471,N_11980,N_10064);
and U15472 (N_15472,N_10787,N_10271);
nand U15473 (N_15473,N_9859,N_10097);
and U15474 (N_15474,N_11066,N_12269);
and U15475 (N_15475,N_12166,N_10883);
or U15476 (N_15476,N_9433,N_11876);
nand U15477 (N_15477,N_9937,N_10349);
and U15478 (N_15478,N_10841,N_12080);
or U15479 (N_15479,N_11167,N_9984);
or U15480 (N_15480,N_10860,N_10748);
nand U15481 (N_15481,N_10035,N_9492);
and U15482 (N_15482,N_9578,N_9519);
nor U15483 (N_15483,N_10387,N_9873);
or U15484 (N_15484,N_10385,N_9727);
xnor U15485 (N_15485,N_10182,N_9997);
nand U15486 (N_15486,N_10797,N_11190);
or U15487 (N_15487,N_9963,N_12023);
or U15488 (N_15488,N_11140,N_11310);
xor U15489 (N_15489,N_9668,N_9672);
and U15490 (N_15490,N_10367,N_9972);
or U15491 (N_15491,N_12170,N_9587);
nand U15492 (N_15492,N_11557,N_10322);
or U15493 (N_15493,N_12419,N_10579);
and U15494 (N_15494,N_10814,N_10770);
or U15495 (N_15495,N_11359,N_10350);
nor U15496 (N_15496,N_9965,N_11932);
nor U15497 (N_15497,N_10682,N_10834);
or U15498 (N_15498,N_11675,N_9586);
and U15499 (N_15499,N_10857,N_10662);
nor U15500 (N_15500,N_11170,N_10698);
nor U15501 (N_15501,N_10764,N_9757);
and U15502 (N_15502,N_11727,N_12307);
and U15503 (N_15503,N_10480,N_12095);
or U15504 (N_15504,N_12240,N_10152);
nand U15505 (N_15505,N_11702,N_10873);
nor U15506 (N_15506,N_12094,N_11252);
or U15507 (N_15507,N_11316,N_11020);
and U15508 (N_15508,N_9816,N_12357);
xor U15509 (N_15509,N_10238,N_12471);
nor U15510 (N_15510,N_10623,N_11652);
nand U15511 (N_15511,N_10749,N_9626);
xor U15512 (N_15512,N_11792,N_9899);
nor U15513 (N_15513,N_10182,N_11143);
nor U15514 (N_15514,N_9678,N_10008);
nand U15515 (N_15515,N_10114,N_9866);
or U15516 (N_15516,N_11520,N_10743);
nand U15517 (N_15517,N_9567,N_12363);
or U15518 (N_15518,N_10647,N_11169);
nor U15519 (N_15519,N_11002,N_10828);
nor U15520 (N_15520,N_10796,N_11743);
nand U15521 (N_15521,N_10146,N_12426);
nor U15522 (N_15522,N_9435,N_10249);
nor U15523 (N_15523,N_12222,N_11822);
or U15524 (N_15524,N_10979,N_9845);
and U15525 (N_15525,N_9659,N_10219);
nor U15526 (N_15526,N_11701,N_9936);
or U15527 (N_15527,N_9703,N_9604);
nor U15528 (N_15528,N_10663,N_9875);
and U15529 (N_15529,N_11454,N_9714);
or U15530 (N_15530,N_9485,N_10930);
and U15531 (N_15531,N_10768,N_10961);
and U15532 (N_15532,N_11939,N_12249);
nor U15533 (N_15533,N_11830,N_10158);
and U15534 (N_15534,N_9844,N_11146);
and U15535 (N_15535,N_9778,N_10824);
or U15536 (N_15536,N_10350,N_11039);
and U15537 (N_15537,N_11917,N_9893);
and U15538 (N_15538,N_9432,N_10781);
nand U15539 (N_15539,N_11250,N_9575);
nor U15540 (N_15540,N_12303,N_10126);
nor U15541 (N_15541,N_11205,N_10681);
or U15542 (N_15542,N_10338,N_11881);
nor U15543 (N_15543,N_12241,N_11875);
nor U15544 (N_15544,N_12420,N_11411);
nor U15545 (N_15545,N_10121,N_9695);
or U15546 (N_15546,N_11183,N_10742);
nor U15547 (N_15547,N_10736,N_11324);
nand U15548 (N_15548,N_12281,N_10690);
nor U15549 (N_15549,N_9512,N_12015);
nand U15550 (N_15550,N_11691,N_11370);
or U15551 (N_15551,N_10566,N_11246);
nor U15552 (N_15552,N_10732,N_10901);
nand U15553 (N_15553,N_11236,N_10745);
and U15554 (N_15554,N_11391,N_10990);
and U15555 (N_15555,N_10463,N_10402);
nor U15556 (N_15556,N_9446,N_11552);
nand U15557 (N_15557,N_12302,N_12270);
nand U15558 (N_15558,N_12397,N_11793);
and U15559 (N_15559,N_12267,N_9876);
nor U15560 (N_15560,N_11944,N_10027);
nand U15561 (N_15561,N_12475,N_11313);
or U15562 (N_15562,N_12376,N_10998);
or U15563 (N_15563,N_12106,N_12058);
nor U15564 (N_15564,N_10192,N_10944);
nor U15565 (N_15565,N_10172,N_10231);
nor U15566 (N_15566,N_11329,N_9475);
xnor U15567 (N_15567,N_10885,N_12164);
nor U15568 (N_15568,N_10334,N_11165);
nand U15569 (N_15569,N_10580,N_12414);
xnor U15570 (N_15570,N_12388,N_10835);
and U15571 (N_15571,N_10328,N_12047);
or U15572 (N_15572,N_12272,N_11070);
xnor U15573 (N_15573,N_12119,N_10228);
xor U15574 (N_15574,N_11204,N_10402);
nor U15575 (N_15575,N_10204,N_10841);
nor U15576 (N_15576,N_10807,N_10563);
or U15577 (N_15577,N_10936,N_10469);
nor U15578 (N_15578,N_9851,N_12350);
or U15579 (N_15579,N_9530,N_10877);
and U15580 (N_15580,N_11703,N_11309);
or U15581 (N_15581,N_10897,N_12160);
nor U15582 (N_15582,N_11729,N_11182);
and U15583 (N_15583,N_12366,N_9845);
and U15584 (N_15584,N_11102,N_9725);
and U15585 (N_15585,N_11250,N_12012);
or U15586 (N_15586,N_10038,N_11944);
nor U15587 (N_15587,N_11492,N_9884);
xor U15588 (N_15588,N_12248,N_11955);
nor U15589 (N_15589,N_11572,N_12040);
nand U15590 (N_15590,N_10449,N_10450);
nand U15591 (N_15591,N_11660,N_11607);
nand U15592 (N_15592,N_10235,N_11024);
and U15593 (N_15593,N_11735,N_12450);
nand U15594 (N_15594,N_10230,N_12200);
or U15595 (N_15595,N_12208,N_10137);
and U15596 (N_15596,N_9564,N_11609);
xor U15597 (N_15597,N_12440,N_11894);
nand U15598 (N_15598,N_12390,N_9639);
nand U15599 (N_15599,N_9570,N_10746);
nor U15600 (N_15600,N_11531,N_11273);
and U15601 (N_15601,N_9401,N_10850);
nand U15602 (N_15602,N_10138,N_12265);
nand U15603 (N_15603,N_11651,N_10378);
nor U15604 (N_15604,N_11225,N_11265);
and U15605 (N_15605,N_9818,N_12417);
nand U15606 (N_15606,N_12112,N_10474);
xnor U15607 (N_15607,N_10583,N_10510);
xor U15608 (N_15608,N_9820,N_11005);
nor U15609 (N_15609,N_10535,N_10729);
or U15610 (N_15610,N_12468,N_10473);
nor U15611 (N_15611,N_9514,N_9996);
and U15612 (N_15612,N_9787,N_10269);
nor U15613 (N_15613,N_11743,N_11120);
nand U15614 (N_15614,N_12265,N_12187);
xor U15615 (N_15615,N_10429,N_10171);
nor U15616 (N_15616,N_11982,N_10117);
or U15617 (N_15617,N_11912,N_11277);
nand U15618 (N_15618,N_10866,N_10152);
or U15619 (N_15619,N_10154,N_9410);
nand U15620 (N_15620,N_9865,N_12233);
and U15621 (N_15621,N_10382,N_9576);
nor U15622 (N_15622,N_10009,N_9861);
and U15623 (N_15623,N_11126,N_10592);
nand U15624 (N_15624,N_10988,N_10046);
nand U15625 (N_15625,N_13303,N_14471);
xor U15626 (N_15626,N_13052,N_13718);
nand U15627 (N_15627,N_13637,N_13757);
and U15628 (N_15628,N_14981,N_14100);
nor U15629 (N_15629,N_13449,N_14166);
xor U15630 (N_15630,N_14107,N_15303);
or U15631 (N_15631,N_13998,N_15283);
and U15632 (N_15632,N_14150,N_15441);
and U15633 (N_15633,N_15431,N_14744);
and U15634 (N_15634,N_15197,N_12910);
xnor U15635 (N_15635,N_13825,N_15310);
nand U15636 (N_15636,N_13871,N_13463);
xnor U15637 (N_15637,N_13858,N_12514);
or U15638 (N_15638,N_14704,N_15457);
and U15639 (N_15639,N_12927,N_13209);
and U15640 (N_15640,N_15026,N_13831);
nor U15641 (N_15641,N_14985,N_13427);
nand U15642 (N_15642,N_14722,N_15616);
nor U15643 (N_15643,N_12717,N_13037);
and U15644 (N_15644,N_13280,N_13496);
and U15645 (N_15645,N_15612,N_14891);
nor U15646 (N_15646,N_12789,N_13768);
nor U15647 (N_15647,N_13863,N_14080);
nor U15648 (N_15648,N_12987,N_14119);
nor U15649 (N_15649,N_14134,N_14627);
nand U15650 (N_15650,N_14896,N_12507);
nor U15651 (N_15651,N_12813,N_12546);
nor U15652 (N_15652,N_15488,N_15450);
xnor U15653 (N_15653,N_12599,N_14784);
nand U15654 (N_15654,N_14738,N_14517);
and U15655 (N_15655,N_14193,N_15142);
and U15656 (N_15656,N_14795,N_12835);
or U15657 (N_15657,N_15069,N_14989);
and U15658 (N_15658,N_13343,N_14213);
nand U15659 (N_15659,N_14460,N_15330);
and U15660 (N_15660,N_13222,N_15273);
or U15661 (N_15661,N_14525,N_15136);
nor U15662 (N_15662,N_13801,N_13595);
nand U15663 (N_15663,N_14350,N_13015);
nor U15664 (N_15664,N_13295,N_14605);
nand U15665 (N_15665,N_12704,N_12685);
nor U15666 (N_15666,N_15478,N_14160);
nor U15667 (N_15667,N_13423,N_14701);
or U15668 (N_15668,N_15139,N_15272);
nand U15669 (N_15669,N_14562,N_13901);
and U15670 (N_15670,N_14415,N_14105);
nor U15671 (N_15671,N_13914,N_12660);
xnor U15672 (N_15672,N_14801,N_13018);
and U15673 (N_15673,N_14546,N_13542);
or U15674 (N_15674,N_14487,N_13421);
or U15675 (N_15675,N_15298,N_14163);
or U15676 (N_15676,N_12715,N_12994);
or U15677 (N_15677,N_14924,N_14096);
or U15678 (N_15678,N_13961,N_12637);
nand U15679 (N_15679,N_14061,N_14198);
or U15680 (N_15680,N_13741,N_15163);
nor U15681 (N_15681,N_13004,N_12547);
and U15682 (N_15682,N_13573,N_15129);
nor U15683 (N_15683,N_15104,N_13869);
nand U15684 (N_15684,N_13809,N_13736);
nand U15685 (N_15685,N_12710,N_14120);
nand U15686 (N_15686,N_13524,N_14805);
xnor U15687 (N_15687,N_13456,N_15153);
nor U15688 (N_15688,N_14216,N_14030);
nor U15689 (N_15689,N_13437,N_13007);
nand U15690 (N_15690,N_12879,N_13928);
nor U15691 (N_15691,N_15524,N_12743);
and U15692 (N_15692,N_14308,N_13604);
and U15693 (N_15693,N_15462,N_13548);
and U15694 (N_15694,N_14716,N_15332);
nor U15695 (N_15695,N_13168,N_12937);
nand U15696 (N_15696,N_15080,N_12884);
nand U15697 (N_15697,N_13239,N_14142);
nor U15698 (N_15698,N_15127,N_14933);
nor U15699 (N_15699,N_15401,N_14382);
nand U15700 (N_15700,N_12672,N_14063);
xnor U15701 (N_15701,N_14913,N_13078);
nand U15702 (N_15702,N_13515,N_15453);
or U15703 (N_15703,N_13795,N_13999);
or U15704 (N_15704,N_12712,N_13192);
xnor U15705 (N_15705,N_13849,N_13138);
xor U15706 (N_15706,N_14175,N_14938);
xnor U15707 (N_15707,N_12572,N_14332);
nand U15708 (N_15708,N_13762,N_15112);
nor U15709 (N_15709,N_14733,N_13461);
or U15710 (N_15710,N_13032,N_14688);
nor U15711 (N_15711,N_14697,N_13603);
nor U15712 (N_15712,N_13645,N_14653);
nor U15713 (N_15713,N_13953,N_13617);
xor U15714 (N_15714,N_15427,N_13157);
nand U15715 (N_15715,N_15046,N_14293);
and U15716 (N_15716,N_15528,N_13142);
and U15717 (N_15717,N_13465,N_12880);
nor U15718 (N_15718,N_12766,N_14541);
nor U15719 (N_15719,N_13674,N_13187);
nor U15720 (N_15720,N_14969,N_14448);
and U15721 (N_15721,N_12655,N_13300);
or U15722 (N_15722,N_12832,N_15154);
xnor U15723 (N_15723,N_15402,N_12550);
or U15724 (N_15724,N_14066,N_13845);
xnor U15725 (N_15725,N_13062,N_14141);
nor U15726 (N_15726,N_12512,N_15603);
and U15727 (N_15727,N_15291,N_14726);
xnor U15728 (N_15728,N_14990,N_12885);
and U15729 (N_15729,N_14632,N_12579);
nor U15730 (N_15730,N_15110,N_12955);
or U15731 (N_15731,N_12700,N_14024);
and U15732 (N_15732,N_13140,N_14077);
xnor U15733 (N_15733,N_13628,N_13931);
and U15734 (N_15734,N_13978,N_13357);
or U15735 (N_15735,N_14016,N_14189);
nor U15736 (N_15736,N_13445,N_15501);
nor U15737 (N_15737,N_14663,N_12658);
nor U15738 (N_15738,N_14219,N_14491);
nor U15739 (N_15739,N_13374,N_15351);
nand U15740 (N_15740,N_12619,N_14666);
or U15741 (N_15741,N_13213,N_13575);
or U15742 (N_15742,N_14789,N_13101);
nor U15743 (N_15743,N_14272,N_15206);
nor U15744 (N_15744,N_13048,N_14164);
and U15745 (N_15745,N_13436,N_12556);
or U15746 (N_15746,N_13266,N_14495);
nand U15747 (N_15747,N_14617,N_14366);
and U15748 (N_15748,N_14446,N_13511);
nand U15749 (N_15749,N_13410,N_15160);
xnor U15750 (N_15750,N_15525,N_13852);
nand U15751 (N_15751,N_13644,N_12582);
nand U15752 (N_15752,N_14537,N_12952);
and U15753 (N_15753,N_14770,N_15105);
or U15754 (N_15754,N_15436,N_15084);
nand U15755 (N_15755,N_13116,N_14354);
or U15756 (N_15756,N_13681,N_13093);
and U15757 (N_15757,N_13236,N_14387);
and U15758 (N_15758,N_14330,N_12600);
and U15759 (N_15759,N_14762,N_14231);
nor U15760 (N_15760,N_13586,N_13574);
nand U15761 (N_15761,N_14872,N_14835);
xor U15762 (N_15762,N_12644,N_14347);
and U15763 (N_15763,N_14118,N_15621);
and U15764 (N_15764,N_12935,N_13036);
and U15765 (N_15765,N_13879,N_14804);
or U15766 (N_15766,N_14612,N_13245);
and U15767 (N_15767,N_14528,N_15252);
xor U15768 (N_15768,N_13383,N_14549);
nand U15769 (N_15769,N_13118,N_15511);
nor U15770 (N_15770,N_14569,N_15366);
xnor U15771 (N_15771,N_12742,N_15352);
or U15772 (N_15772,N_14151,N_14881);
xnor U15773 (N_15773,N_12526,N_13751);
nand U15774 (N_15774,N_13419,N_14684);
or U15775 (N_15775,N_12777,N_13030);
nand U15776 (N_15776,N_15463,N_13925);
xor U15777 (N_15777,N_14021,N_15417);
and U15778 (N_15778,N_15338,N_13349);
nand U15779 (N_15779,N_15029,N_13550);
and U15780 (N_15780,N_12881,N_15128);
nor U15781 (N_15781,N_14638,N_15168);
nor U15782 (N_15782,N_13022,N_15063);
or U15783 (N_15783,N_13388,N_14966);
nor U15784 (N_15784,N_14402,N_14877);
or U15785 (N_15785,N_14004,N_14052);
and U15786 (N_15786,N_15367,N_14936);
and U15787 (N_15787,N_12652,N_14585);
nand U15788 (N_15788,N_12844,N_12862);
nand U15789 (N_15789,N_13003,N_12570);
and U15790 (N_15790,N_15238,N_13085);
or U15791 (N_15791,N_13360,N_13166);
and U15792 (N_15792,N_14391,N_14386);
nand U15793 (N_15793,N_15259,N_14509);
xor U15794 (N_15794,N_14081,N_12576);
nand U15795 (N_15795,N_12508,N_13875);
or U15796 (N_15796,N_14905,N_14453);
nand U15797 (N_15797,N_12867,N_13959);
nand U15798 (N_15798,N_15594,N_12820);
xnor U15799 (N_15799,N_13348,N_12569);
nand U15800 (N_15800,N_13703,N_14503);
nor U15801 (N_15801,N_14450,N_12774);
and U15802 (N_15802,N_12778,N_15073);
or U15803 (N_15803,N_14581,N_15204);
nand U15804 (N_15804,N_14311,N_14642);
and U15805 (N_15805,N_14480,N_12977);
and U15806 (N_15806,N_14616,N_12945);
and U15807 (N_15807,N_12634,N_14691);
and U15808 (N_15808,N_12960,N_15246);
or U15809 (N_15809,N_15543,N_13597);
or U15810 (N_15810,N_15487,N_13340);
nand U15811 (N_15811,N_14922,N_13540);
nand U15812 (N_15812,N_14147,N_15005);
or U15813 (N_15813,N_14333,N_15409);
nand U15814 (N_15814,N_15424,N_13218);
xnor U15815 (N_15815,N_13938,N_15389);
nor U15816 (N_15816,N_15025,N_13929);
nor U15817 (N_15817,N_15531,N_15514);
or U15818 (N_15818,N_14492,N_15593);
nor U15819 (N_15819,N_13927,N_12947);
xnor U15820 (N_15820,N_14619,N_14436);
and U15821 (N_15821,N_12703,N_14045);
or U15822 (N_15822,N_15510,N_13664);
nor U15823 (N_15823,N_13697,N_12830);
nand U15824 (N_15824,N_13194,N_14859);
nand U15825 (N_15825,N_14847,N_13792);
nor U15826 (N_15826,N_13273,N_15195);
or U15827 (N_15827,N_14582,N_14609);
and U15828 (N_15828,N_14793,N_15242);
nor U15829 (N_15829,N_15434,N_12590);
nand U15830 (N_15830,N_15185,N_14470);
or U15831 (N_15831,N_14740,N_15486);
nor U15832 (N_15832,N_12966,N_14615);
and U15833 (N_15833,N_13226,N_12536);
and U15834 (N_15834,N_15212,N_13397);
and U15835 (N_15835,N_14845,N_15465);
nor U15836 (N_15836,N_14679,N_14496);
and U15837 (N_15837,N_12868,N_15569);
or U15838 (N_15838,N_14978,N_13217);
or U15839 (N_15839,N_12971,N_12585);
nand U15840 (N_15840,N_13881,N_12523);
nor U15841 (N_15841,N_14370,N_12900);
nand U15842 (N_15842,N_13054,N_13943);
nand U15843 (N_15843,N_14056,N_13250);
or U15844 (N_15844,N_13319,N_13046);
and U15845 (N_15845,N_13313,N_13882);
nor U15846 (N_15846,N_12815,N_13560);
or U15847 (N_15847,N_14839,N_14786);
and U15848 (N_15848,N_14239,N_13123);
nor U15849 (N_15849,N_14048,N_14826);
or U15850 (N_15850,N_14959,N_14787);
xor U15851 (N_15851,N_13840,N_14817);
xnor U15852 (N_15852,N_13492,N_13316);
and U15853 (N_15853,N_12714,N_14128);
and U15854 (N_15854,N_12554,N_14458);
nand U15855 (N_15855,N_12964,N_14836);
and U15856 (N_15856,N_14785,N_14245);
nand U15857 (N_15857,N_14089,N_13296);
or U15858 (N_15858,N_14571,N_14490);
nand U15859 (N_15859,N_14428,N_12968);
nor U15860 (N_15860,N_15250,N_12709);
xor U15861 (N_15861,N_15047,N_12924);
or U15862 (N_15862,N_15287,N_12682);
and U15863 (N_15863,N_14346,N_13092);
nor U15864 (N_15864,N_14850,N_12728);
nor U15865 (N_15865,N_15152,N_13893);
and U15866 (N_15866,N_14713,N_14282);
nand U15867 (N_15867,N_14326,N_14328);
nand U15868 (N_15868,N_15432,N_12852);
and U15869 (N_15869,N_15349,N_13598);
xor U15870 (N_15870,N_15169,N_12756);
or U15871 (N_15871,N_13344,N_15233);
or U15872 (N_15872,N_13827,N_13873);
and U15873 (N_15873,N_13005,N_13872);
nor U15874 (N_15874,N_13447,N_12588);
nor U15875 (N_15875,N_13081,N_15591);
nor U15876 (N_15876,N_14814,N_14512);
or U15877 (N_15877,N_13988,N_12874);
nor U15878 (N_15878,N_15364,N_13384);
xnor U15879 (N_15879,N_14900,N_13038);
nand U15880 (N_15880,N_14778,N_12587);
or U15881 (N_15881,N_13124,N_13195);
and U15882 (N_15882,N_13017,N_13774);
nor U15883 (N_15883,N_15035,N_13089);
or U15884 (N_15884,N_13446,N_13727);
or U15885 (N_15885,N_14463,N_14079);
nand U15886 (N_15886,N_13474,N_12785);
or U15887 (N_15887,N_14379,N_15535);
nor U15888 (N_15888,N_15170,N_15395);
or U15889 (N_15889,N_12519,N_12779);
or U15890 (N_15890,N_15559,N_14940);
or U15891 (N_15891,N_13538,N_12916);
nor U15892 (N_15892,N_15052,N_12621);
nor U15893 (N_15893,N_14735,N_13663);
or U15894 (N_15894,N_14015,N_15408);
and U15895 (N_15895,N_14485,N_13534);
xor U15896 (N_15896,N_14920,N_12985);
nor U15897 (N_15897,N_12962,N_14305);
xnor U15898 (N_15898,N_14756,N_13094);
nand U15899 (N_15899,N_14515,N_15076);
xor U15900 (N_15900,N_12828,N_15467);
nor U15901 (N_15901,N_13691,N_13071);
nor U15902 (N_15902,N_15227,N_12936);
nor U15903 (N_15903,N_14739,N_12974);
nor U15904 (N_15904,N_13047,N_14218);
or U15905 (N_15905,N_14010,N_15201);
nand U15906 (N_15906,N_12842,N_13196);
and U15907 (N_15907,N_13522,N_13985);
nor U15908 (N_15908,N_13455,N_14685);
nand U15909 (N_15909,N_15159,N_15060);
nor U15910 (N_15910,N_13802,N_14340);
nor U15911 (N_15911,N_14675,N_15605);
nor U15912 (N_15912,N_15387,N_14906);
nand U15913 (N_15913,N_15053,N_13719);
and U15914 (N_15914,N_12817,N_14334);
and U15915 (N_15915,N_12539,N_14640);
and U15916 (N_15916,N_13365,N_14404);
nand U15917 (N_15917,N_14909,N_12689);
xor U15918 (N_15918,N_14136,N_14019);
nor U15919 (N_15919,N_12791,N_14047);
and U15920 (N_15920,N_14662,N_14182);
or U15921 (N_15921,N_14409,N_14676);
and U15922 (N_15922,N_13997,N_12782);
and U15923 (N_15923,N_13722,N_13278);
and U15924 (N_15924,N_14523,N_15499);
or U15925 (N_15925,N_14540,N_14466);
nand U15926 (N_15926,N_13987,N_14302);
or U15927 (N_15927,N_13509,N_13279);
and U15928 (N_15928,N_13439,N_13750);
nor U15929 (N_15929,N_14968,N_14344);
xor U15930 (N_15930,N_14860,N_15343);
or U15931 (N_15931,N_13761,N_15299);
and U15932 (N_15932,N_15507,N_15429);
nand U15933 (N_15933,N_12719,N_14337);
and U15934 (N_15934,N_14715,N_14618);
and U15935 (N_15935,N_14901,N_14037);
and U15936 (N_15936,N_14647,N_15393);
or U15937 (N_15937,N_12846,N_15164);
xnor U15938 (N_15938,N_12513,N_12559);
and U15939 (N_15939,N_14600,N_12839);
or U15940 (N_15940,N_15547,N_15082);
nor U15941 (N_15941,N_13412,N_15541);
nand U15942 (N_15942,N_14791,N_15439);
nand U15943 (N_15943,N_13561,N_12821);
nor U15944 (N_15944,N_14620,N_12608);
nand U15945 (N_15945,N_14846,N_13462);
nand U15946 (N_15946,N_13023,N_15526);
nor U15947 (N_15947,N_12873,N_15357);
and U15948 (N_15948,N_14204,N_13130);
nand U15949 (N_15949,N_12976,N_14290);
or U15950 (N_15950,N_14225,N_14320);
or U15951 (N_15951,N_13027,N_13654);
or U15952 (N_15952,N_15489,N_14518);
nor U15953 (N_15953,N_15613,N_14547);
nand U15954 (N_15954,N_14158,N_12921);
nor U15955 (N_15955,N_15515,N_12975);
and U15956 (N_15956,N_13921,N_13711);
or U15957 (N_15957,N_12598,N_13525);
and U15958 (N_15958,N_13473,N_13238);
or U15959 (N_15959,N_14601,N_15266);
nand U15960 (N_15960,N_13353,N_15406);
and U15961 (N_15961,N_14129,N_15070);
or U15962 (N_15962,N_14177,N_15589);
xor U15963 (N_15963,N_15325,N_15473);
nand U15964 (N_15964,N_13963,N_12631);
and U15965 (N_15965,N_14036,N_15058);
or U15966 (N_15966,N_12750,N_15057);
or U15967 (N_15967,N_13790,N_14194);
nand U15968 (N_15968,N_13165,N_13989);
and U15969 (N_15969,N_13315,N_15031);
and U15970 (N_15970,N_14455,N_14892);
nor U15971 (N_15971,N_14108,N_14763);
or U15972 (N_15972,N_14263,N_14751);
or U15973 (N_15973,N_13351,N_13002);
nor U15974 (N_15974,N_15567,N_14026);
and U15975 (N_15975,N_15010,N_14286);
and U15976 (N_15976,N_14809,N_12687);
nor U15977 (N_15977,N_14545,N_12995);
and U15978 (N_15978,N_12946,N_12515);
and U15979 (N_15979,N_14144,N_15100);
and U15980 (N_15980,N_14536,N_15041);
or U15981 (N_15981,N_13739,N_13390);
nor U15982 (N_15982,N_12573,N_12537);
and U15983 (N_15983,N_14017,N_14122);
nand U15984 (N_15984,N_13610,N_12959);
nand U15985 (N_15985,N_15032,N_13960);
nor U15986 (N_15986,N_13401,N_13075);
and U15987 (N_15987,N_14309,N_13744);
nand U15988 (N_15988,N_14777,N_15111);
and U15989 (N_15989,N_15231,N_14696);
nor U15990 (N_15990,N_15089,N_14964);
nand U15991 (N_15991,N_15248,N_14613);
and U15992 (N_15992,N_13571,N_13588);
nand U15993 (N_15993,N_14325,N_14092);
and U15994 (N_15994,N_12613,N_15302);
nand U15995 (N_15995,N_14230,N_12557);
nor U15996 (N_15996,N_13339,N_15203);
and U15997 (N_15997,N_14729,N_13899);
nand U15998 (N_15998,N_12929,N_14472);
nor U15999 (N_15999,N_12716,N_13188);
nor U16000 (N_16000,N_14068,N_13930);
and U16001 (N_16001,N_15324,N_15006);
nor U16002 (N_16002,N_15147,N_12713);
nor U16003 (N_16003,N_13778,N_13659);
nand U16004 (N_16004,N_13033,N_12811);
nor U16005 (N_16005,N_15433,N_14773);
nand U16006 (N_16006,N_15261,N_13621);
nor U16007 (N_16007,N_13889,N_14256);
and U16008 (N_16008,N_15297,N_13712);
and U16009 (N_16009,N_14228,N_15372);
nand U16010 (N_16010,N_14335,N_13570);
nand U16011 (N_16011,N_15295,N_15624);
and U16012 (N_16012,N_13748,N_15358);
nand U16013 (N_16013,N_13624,N_13887);
nor U16014 (N_16014,N_12906,N_14890);
nand U16015 (N_16015,N_14608,N_14291);
or U16016 (N_16016,N_13162,N_14479);
nand U16017 (N_16017,N_15506,N_13776);
or U16018 (N_16018,N_14067,N_12653);
xnor U16019 (N_16019,N_13133,N_13983);
nor U16020 (N_16020,N_12965,N_12659);
xor U16021 (N_16021,N_14400,N_14950);
or U16022 (N_16022,N_14539,N_13145);
nand U16023 (N_16023,N_13034,N_12577);
and U16024 (N_16024,N_12961,N_13008);
nor U16025 (N_16025,N_14693,N_14395);
or U16026 (N_16026,N_14887,N_13482);
or U16027 (N_16027,N_15336,N_12767);
xnor U16028 (N_16028,N_15173,N_12727);
nand U16029 (N_16029,N_15071,N_14780);
nand U16030 (N_16030,N_13454,N_14831);
nor U16031 (N_16031,N_13497,N_14630);
nor U16032 (N_16032,N_15456,N_14829);
nand U16033 (N_16033,N_13836,N_12905);
and U16034 (N_16034,N_13488,N_15377);
or U16035 (N_16035,N_14447,N_13345);
nand U16036 (N_16036,N_15239,N_13376);
or U16037 (N_16037,N_12847,N_14975);
or U16038 (N_16038,N_14110,N_13656);
or U16039 (N_16039,N_13520,N_14664);
nor U16040 (N_16040,N_12705,N_13111);
nor U16041 (N_16041,N_14898,N_13706);
and U16042 (N_16042,N_15210,N_15500);
nand U16043 (N_16043,N_13695,N_13521);
nand U16044 (N_16044,N_12702,N_15400);
xnor U16045 (N_16045,N_13063,N_13917);
xnor U16046 (N_16046,N_15421,N_14774);
nand U16047 (N_16047,N_14614,N_13884);
and U16048 (N_16048,N_15091,N_14610);
and U16049 (N_16049,N_13058,N_14866);
or U16050 (N_16050,N_15056,N_12612);
xor U16051 (N_16051,N_14465,N_13916);
or U16052 (N_16052,N_13077,N_14532);
nor U16053 (N_16053,N_13798,N_15037);
and U16054 (N_16054,N_14377,N_14645);
and U16055 (N_16055,N_12931,N_13688);
and U16056 (N_16056,N_13318,N_15097);
nand U16057 (N_16057,N_13948,N_13268);
nand U16058 (N_16058,N_12530,N_13641);
or U16059 (N_16059,N_13422,N_14488);
or U16060 (N_16060,N_13811,N_14375);
nand U16061 (N_16061,N_15245,N_13783);
or U16062 (N_16062,N_14734,N_14520);
or U16063 (N_16063,N_13532,N_13380);
and U16064 (N_16064,N_13584,N_14819);
nor U16065 (N_16065,N_15600,N_13231);
xnor U16066 (N_16066,N_14498,N_15015);
and U16067 (N_16067,N_14656,N_13600);
or U16068 (N_16068,N_12763,N_14552);
and U16069 (N_16069,N_13945,N_14345);
nand U16070 (N_16070,N_12963,N_13216);
or U16071 (N_16071,N_12648,N_14168);
nor U16072 (N_16072,N_14307,N_14051);
nand U16073 (N_16073,N_13627,N_15077);
or U16074 (N_16074,N_14790,N_12678);
nor U16075 (N_16075,N_14316,N_15183);
nand U16076 (N_16076,N_15419,N_15597);
nor U16077 (N_16077,N_14979,N_13487);
nand U16078 (N_16078,N_12892,N_13387);
nor U16079 (N_16079,N_14823,N_13633);
nand U16080 (N_16080,N_12509,N_12662);
and U16081 (N_16081,N_14992,N_12650);
and U16082 (N_16082,N_14069,N_13503);
or U16083 (N_16083,N_13336,N_12500);
or U16084 (N_16084,N_13844,N_15476);
nor U16085 (N_16085,N_13284,N_12748);
nand U16086 (N_16086,N_12969,N_12984);
nand U16087 (N_16087,N_15138,N_12849);
and U16088 (N_16088,N_15171,N_13108);
or U16089 (N_16089,N_12617,N_12810);
and U16090 (N_16090,N_14659,N_13174);
nand U16091 (N_16091,N_14965,N_15584);
or U16092 (N_16092,N_15444,N_15051);
or U16093 (N_16093,N_13459,N_14943);
nand U16094 (N_16094,N_13112,N_12816);
and U16095 (N_16095,N_12534,N_13724);
or U16096 (N_16096,N_12664,N_14806);
nor U16097 (N_16097,N_12795,N_13406);
nand U16098 (N_16098,N_14811,N_15296);
or U16099 (N_16099,N_15382,N_15546);
nand U16100 (N_16100,N_13740,N_12744);
and U16101 (N_16101,N_12551,N_13428);
or U16102 (N_16102,N_13682,N_13526);
nand U16103 (N_16103,N_13176,N_14639);
and U16104 (N_16104,N_14646,N_14669);
xnor U16105 (N_16105,N_13403,N_15240);
or U16106 (N_16106,N_14941,N_13854);
nor U16107 (N_16107,N_12610,N_13638);
nand U16108 (N_16108,N_14348,N_14449);
nand U16109 (N_16109,N_14511,N_15228);
nor U16110 (N_16110,N_14481,N_12555);
nand U16111 (N_16111,N_13211,N_14202);
nor U16112 (N_16112,N_14658,N_14956);
or U16113 (N_16113,N_14857,N_15008);
nand U16114 (N_16114,N_12567,N_12749);
and U16115 (N_16115,N_12772,N_13787);
nand U16116 (N_16116,N_13354,N_12630);
xnor U16117 (N_16117,N_14644,N_14904);
nand U16118 (N_16118,N_12657,N_12647);
nand U16119 (N_16119,N_14962,N_15443);
nor U16120 (N_16120,N_12616,N_14085);
nand U16121 (N_16121,N_13677,N_12601);
or U16122 (N_16122,N_14603,N_15512);
or U16123 (N_16123,N_14832,N_14882);
xor U16124 (N_16124,N_14258,N_12901);
nor U16125 (N_16125,N_12691,N_15549);
and U16126 (N_16126,N_15420,N_13764);
nand U16127 (N_16127,N_13936,N_15083);
or U16128 (N_16128,N_14815,N_13493);
and U16129 (N_16129,N_14923,N_13533);
or U16130 (N_16130,N_14533,N_13322);
nor U16131 (N_16131,N_13924,N_13755);
nor U16132 (N_16132,N_13072,N_12524);
nand U16133 (N_16133,N_13829,N_13060);
xnor U16134 (N_16134,N_14702,N_12690);
nor U16135 (N_16135,N_15038,N_12799);
nor U16136 (N_16136,N_14957,N_13941);
and U16137 (N_16137,N_14433,N_13708);
nor U16138 (N_16138,N_13992,N_13504);
xnor U16139 (N_16139,N_14671,N_15207);
or U16140 (N_16140,N_13651,N_14323);
and U16141 (N_16141,N_13678,N_14526);
or U16142 (N_16142,N_14628,N_13932);
and U16143 (N_16143,N_12997,N_14444);
nor U16144 (N_16144,N_13772,N_13786);
and U16145 (N_16145,N_14649,N_14214);
or U16146 (N_16146,N_13670,N_12646);
or U16147 (N_16147,N_14915,N_15007);
nand U16148 (N_16148,N_13311,N_13568);
nand U16149 (N_16149,N_15255,N_12988);
or U16150 (N_16150,N_13479,N_15306);
nor U16151 (N_16151,N_15184,N_13167);
or U16152 (N_16152,N_12798,N_12720);
or U16153 (N_16153,N_14893,N_13946);
nor U16154 (N_16154,N_14939,N_13649);
nand U16155 (N_16155,N_13257,N_15096);
and U16156 (N_16156,N_15576,N_14998);
nand U16157 (N_16157,N_13562,N_15378);
nand U16158 (N_16158,N_14102,N_13729);
and U16159 (N_16159,N_14871,N_15064);
nor U16160 (N_16160,N_12677,N_14279);
nor U16161 (N_16161,N_14970,N_14322);
nor U16162 (N_16162,N_13952,N_13274);
and U16163 (N_16163,N_15485,N_14631);
nor U16164 (N_16164,N_14139,N_13769);
and U16165 (N_16165,N_14131,N_12615);
nor U16166 (N_16166,N_13824,N_13347);
or U16167 (N_16167,N_15085,N_12746);
or U16168 (N_16168,N_14876,N_15368);
and U16169 (N_16169,N_14183,N_12845);
xnor U16170 (N_16170,N_14808,N_13745);
and U16171 (N_16171,N_13888,N_12869);
nand U16172 (N_16172,N_14953,N_14265);
nand U16173 (N_16173,N_13913,N_15373);
nand U16174 (N_16174,N_13480,N_15290);
and U16175 (N_16175,N_15042,N_14583);
nand U16176 (N_16176,N_13726,N_12629);
or U16177 (N_16177,N_13833,N_15107);
nand U16178 (N_16178,N_15274,N_12790);
nor U16179 (N_16179,N_14604,N_13232);
and U16180 (N_16180,N_13285,N_15571);
nor U16181 (N_16181,N_14554,N_15622);
nand U16182 (N_16182,N_13850,N_15209);
or U16183 (N_16183,N_14931,N_14457);
xnor U16184 (N_16184,N_13244,N_15361);
nor U16185 (N_16185,N_12754,N_14797);
or U16186 (N_16186,N_14314,N_14935);
nand U16187 (N_16187,N_13970,N_15012);
xnor U16188 (N_16188,N_13301,N_15321);
or U16189 (N_16189,N_13981,N_14897);
or U16190 (N_16190,N_14754,N_14262);
and U16191 (N_16191,N_13158,N_14753);
nor U16192 (N_16192,N_14925,N_12581);
or U16193 (N_16193,N_14556,N_13856);
nor U16194 (N_16194,N_13813,N_14889);
nor U16195 (N_16195,N_15529,N_14140);
or U16196 (N_16196,N_15619,N_15494);
and U16197 (N_16197,N_14201,N_14264);
or U16198 (N_16198,N_12893,N_13328);
nor U16199 (N_16199,N_15573,N_14281);
nand U16200 (N_16200,N_15004,N_13478);
nand U16201 (N_16201,N_14432,N_14721);
nor U16202 (N_16202,N_12943,N_14456);
nand U16203 (N_16203,N_14090,N_13483);
and U16204 (N_16204,N_12718,N_13966);
or U16205 (N_16205,N_13012,N_14779);
xor U16206 (N_16206,N_15043,N_13730);
and U16207 (N_16207,N_13519,N_14558);
or U16208 (N_16208,N_15354,N_12684);
nand U16209 (N_16209,N_13203,N_15162);
nor U16210 (N_16210,N_12980,N_13632);
or U16211 (N_16211,N_15502,N_14123);
and U16212 (N_16212,N_14430,N_14011);
xor U16213 (N_16213,N_14974,N_14971);
or U16214 (N_16214,N_14827,N_14462);
nand U16215 (N_16215,N_14440,N_14879);
or U16216 (N_16216,N_13214,N_12560);
and U16217 (N_16217,N_14083,N_13086);
xor U16218 (N_16218,N_13199,N_12865);
xnor U16219 (N_16219,N_15346,N_13470);
nor U16220 (N_16220,N_12566,N_12991);
or U16221 (N_16221,N_13883,N_14999);
nor U16222 (N_16222,N_13846,N_14411);
nand U16223 (N_16223,N_14544,N_12940);
nand U16224 (N_16224,N_13105,N_13206);
and U16225 (N_16225,N_13502,N_14486);
or U16226 (N_16226,N_12930,N_13594);
or U16227 (N_16227,N_15430,N_13450);
and U16228 (N_16228,N_14046,N_13716);
and U16229 (N_16229,N_14578,N_12641);
nand U16230 (N_16230,N_14499,N_13732);
and U16231 (N_16231,N_13171,N_13804);
nor U16232 (N_16232,N_14306,N_14180);
and U16233 (N_16233,N_14908,N_13352);
nand U16234 (N_16234,N_15277,N_13013);
nand U16235 (N_16235,N_15289,N_13263);
nand U16236 (N_16236,N_15123,N_13867);
and U16237 (N_16237,N_14972,N_12639);
or U16238 (N_16238,N_15208,N_15193);
nor U16239 (N_16239,N_12871,N_13705);
or U16240 (N_16240,N_14982,N_13227);
nor U16241 (N_16241,N_15570,N_13639);
or U16242 (N_16242,N_14802,N_14431);
or U16243 (N_16243,N_14874,N_14012);
xor U16244 (N_16244,N_15061,N_14994);
nor U16245 (N_16245,N_14519,N_13529);
and U16246 (N_16246,N_14339,N_15556);
or U16247 (N_16247,N_14072,N_13735);
xor U16248 (N_16248,N_13056,N_14186);
and U16249 (N_16249,N_15194,N_14765);
nor U16250 (N_16250,N_13942,N_14243);
xnor U16251 (N_16251,N_15544,N_14574);
or U16252 (N_16252,N_13779,N_14768);
nand U16253 (N_16253,N_13541,N_12792);
and U16254 (N_16254,N_15609,N_12732);
xnor U16255 (N_16255,N_14008,N_14426);
nand U16256 (N_16256,N_14208,N_15375);
nor U16257 (N_16257,N_15044,N_12752);
nor U16258 (N_16258,N_15258,N_14224);
or U16259 (N_16259,N_14174,N_14250);
xor U16260 (N_16260,N_12698,N_13020);
xor U16261 (N_16261,N_13902,N_13499);
and U16262 (N_16262,N_13233,N_13686);
xor U16263 (N_16263,N_12780,N_12620);
nor U16264 (N_16264,N_13964,N_15000);
and U16265 (N_16265,N_13259,N_14405);
xor U16266 (N_16266,N_13193,N_14318);
nor U16267 (N_16267,N_13874,N_14445);
or U16268 (N_16268,N_15217,N_15280);
or U16269 (N_16269,N_14295,N_13860);
or U16270 (N_16270,N_13127,N_13837);
and U16271 (N_16271,N_13143,N_15561);
nand U16272 (N_16272,N_13506,N_14624);
or U16273 (N_16273,N_15093,N_14407);
nor U16274 (N_16274,N_12797,N_13373);
nor U16275 (N_16275,N_15065,N_14476);
xnor U16276 (N_16276,N_13782,N_13746);
nand U16277 (N_16277,N_14563,N_13098);
nand U16278 (N_16278,N_13460,N_12898);
nand U16279 (N_16279,N_14543,N_13329);
nand U16280 (N_16280,N_15405,N_15001);
xor U16281 (N_16281,N_13894,N_14728);
nor U16282 (N_16282,N_12800,N_15319);
and U16283 (N_16283,N_13104,N_15394);
and U16284 (N_16284,N_13685,N_15229);
nand U16285 (N_16285,N_15519,N_13491);
nand U16286 (N_16286,N_14014,N_15523);
xnor U16287 (N_16287,N_13605,N_13781);
and U16288 (N_16288,N_13191,N_15021);
nor U16289 (N_16289,N_12680,N_13859);
and U16290 (N_16290,N_13000,N_15282);
and U16291 (N_16291,N_13453,N_14126);
and U16292 (N_16292,N_15144,N_14454);
nand U16293 (N_16293,N_13088,N_13702);
or U16294 (N_16294,N_13147,N_13163);
or U16295 (N_16295,N_13968,N_15224);
xor U16296 (N_16296,N_15318,N_13613);
and U16297 (N_16297,N_14727,N_13861);
xor U16298 (N_16298,N_14672,N_12541);
nand U16299 (N_16299,N_12517,N_14331);
xor U16300 (N_16300,N_14820,N_15265);
xor U16301 (N_16301,N_12505,N_14502);
and U16302 (N_16302,N_13069,N_12696);
nor U16303 (N_16303,N_13271,N_13413);
and U16304 (N_16304,N_15566,N_13601);
or U16305 (N_16305,N_15381,N_12808);
nor U16306 (N_16306,N_15604,N_14927);
or U16307 (N_16307,N_13558,N_14137);
xor U16308 (N_16308,N_12957,N_15410);
nand U16309 (N_16309,N_13405,N_13338);
or U16310 (N_16310,N_13255,N_15086);
nor U16311 (N_16311,N_13418,N_15254);
and U16312 (N_16312,N_12848,N_14260);
or U16313 (N_16313,N_14145,N_15610);
or U16314 (N_16314,N_12543,N_13200);
and U16315 (N_16315,N_12825,N_13399);
nand U16316 (N_16316,N_15016,N_13673);
and U16317 (N_16317,N_14719,N_13207);
and U16318 (N_16318,N_13544,N_14963);
nor U16319 (N_16319,N_12611,N_14022);
xnor U16320 (N_16320,N_15126,N_14570);
or U16321 (N_16321,N_15333,N_12903);
nor U16322 (N_16322,N_13415,N_13949);
nor U16323 (N_16323,N_15247,N_12838);
nand U16324 (N_16324,N_12506,N_14828);
and U16325 (N_16325,N_13070,N_14760);
and U16326 (N_16326,N_12920,N_14916);
or U16327 (N_16327,N_13177,N_15508);
or U16328 (N_16328,N_13619,N_14369);
nand U16329 (N_16329,N_13366,N_15607);
nand U16330 (N_16330,N_15284,N_14842);
and U16331 (N_16331,N_13229,N_12673);
or U16332 (N_16332,N_15268,N_13572);
or U16333 (N_16333,N_15308,N_14577);
nand U16334 (N_16334,N_15314,N_14967);
and U16335 (N_16335,N_13057,N_12733);
or U16336 (N_16336,N_12938,N_13103);
and U16337 (N_16337,N_13224,N_14268);
nor U16338 (N_16338,N_15281,N_13066);
or U16339 (N_16339,N_13016,N_12768);
nor U16340 (N_16340,N_15516,N_12899);
or U16341 (N_16341,N_13299,N_14775);
nand U16342 (N_16342,N_14741,N_14435);
nor U16343 (N_16343,N_14530,N_14643);
xnor U16344 (N_16344,N_14991,N_15099);
or U16345 (N_16345,N_13951,N_13918);
nand U16346 (N_16346,N_14712,N_14342);
nand U16347 (N_16347,N_14580,N_15305);
nand U16348 (N_16348,N_12914,N_12870);
nor U16349 (N_16349,N_12833,N_12973);
and U16350 (N_16350,N_13714,N_12604);
nand U16351 (N_16351,N_14686,N_12902);
or U16352 (N_16352,N_15596,N_15158);
nor U16353 (N_16353,N_13358,N_15518);
xnor U16354 (N_16354,N_12972,N_14223);
nor U16355 (N_16355,N_13976,N_13471);
or U16356 (N_16356,N_14976,N_13045);
nor U16357 (N_16357,N_15435,N_14508);
nor U16358 (N_16358,N_12671,N_15578);
or U16359 (N_16359,N_14414,N_15028);
or U16360 (N_16360,N_14199,N_13566);
nor U16361 (N_16361,N_14759,N_14594);
or U16362 (N_16362,N_13791,N_13053);
nand U16363 (N_16363,N_13747,N_15527);
and U16364 (N_16364,N_14363,N_12504);
nor U16365 (N_16365,N_15474,N_13234);
or U16366 (N_16366,N_14210,N_14222);
nor U16367 (N_16367,N_13289,N_15304);
or U16368 (N_16368,N_15461,N_12669);
nand U16369 (N_16369,N_12913,N_12887);
nand U16370 (N_16370,N_14961,N_15188);
or U16371 (N_16371,N_14681,N_14798);
or U16372 (N_16372,N_15562,N_13440);
xor U16373 (N_16373,N_14598,N_14113);
or U16374 (N_16374,N_14364,N_13490);
nand U16375 (N_16375,N_13583,N_15264);
nand U16376 (N_16376,N_13457,N_14737);
nand U16377 (N_16377,N_13495,N_13430);
or U16378 (N_16378,N_15390,N_12967);
and U16379 (N_16379,N_12759,N_14229);
or U16380 (N_16380,N_13201,N_14973);
or U16381 (N_16381,N_13475,N_14403);
nor U16382 (N_16382,N_15504,N_14687);
nand U16383 (N_16383,N_14474,N_13261);
nor U16384 (N_16384,N_13178,N_13508);
and U16385 (N_16385,N_14883,N_14338);
nand U16386 (N_16386,N_14853,N_13102);
nand U16387 (N_16387,N_13996,N_13725);
nand U16388 (N_16388,N_14075,N_14438);
and U16389 (N_16389,N_13580,N_13760);
nor U16390 (N_16390,N_14235,N_13675);
and U16391 (N_16391,N_15331,N_12805);
and U16392 (N_16392,N_14705,N_12622);
or U16393 (N_16393,N_15601,N_15532);
or U16394 (N_16394,N_15055,N_12950);
and U16395 (N_16395,N_12706,N_12624);
and U16396 (N_16396,N_15167,N_12731);
xor U16397 (N_16397,N_15220,N_15216);
nor U16398 (N_16398,N_15491,N_13923);
nand U16399 (N_16399,N_14718,N_13185);
or U16400 (N_16400,N_13276,N_15146);
or U16401 (N_16401,N_14093,N_14568);
or U16402 (N_16402,N_13051,N_14196);
or U16403 (N_16403,N_13982,N_14034);
xor U16404 (N_16404,N_14864,N_12683);
or U16405 (N_16405,N_14368,N_12738);
nand U16406 (N_16406,N_13839,N_12986);
nor U16407 (N_16407,N_13333,N_14091);
or U16408 (N_16408,N_13986,N_15425);
or U16409 (N_16409,N_14007,N_15572);
or U16410 (N_16410,N_14781,N_13129);
and U16411 (N_16411,N_13110,N_13050);
nor U16412 (N_16412,N_13665,N_13398);
nor U16413 (N_16413,N_12638,N_15180);
xor U16414 (N_16414,N_14947,N_13838);
nand U16415 (N_16415,N_13990,N_14694);
and U16416 (N_16416,N_14257,N_15013);
nor U16417 (N_16417,N_14641,N_13247);
and U16418 (N_16418,N_13106,N_12679);
nand U16419 (N_16419,N_15285,N_14944);
nand U16420 (N_16420,N_14534,N_13847);
or U16421 (N_16421,N_13417,N_13518);
and U16422 (N_16422,N_15440,N_13434);
nor U16423 (N_16423,N_13820,N_14167);
and U16424 (N_16424,N_13785,N_13608);
and U16425 (N_16425,N_15386,N_14220);
and U16426 (N_16426,N_12516,N_14413);
or U16427 (N_16427,N_15023,N_14009);
nor U16428 (N_16428,N_13467,N_13694);
and U16429 (N_16429,N_14668,N_14116);
and U16430 (N_16430,N_12596,N_14782);
or U16431 (N_16431,N_13306,N_12584);
and U16432 (N_16432,N_14948,N_15448);
and U16433 (N_16433,N_12753,N_13965);
or U16434 (N_16434,N_14750,N_13843);
nor U16435 (N_16435,N_14564,N_12531);
nor U16436 (N_16436,N_13485,N_14840);
or U16437 (N_16437,N_14524,N_15223);
xnor U16438 (N_16438,N_13636,N_13749);
and U16439 (N_16439,N_13246,N_15481);
and U16440 (N_16440,N_14551,N_13341);
xor U16441 (N_16441,N_14360,N_12535);
nand U16442 (N_16442,N_14548,N_13367);
nor U16443 (N_16443,N_13593,N_13717);
nand U16444 (N_16444,N_12699,N_12804);
and U16445 (N_16445,N_13876,N_14195);
and U16446 (N_16446,N_13737,N_12912);
nand U16447 (N_16447,N_13614,N_15106);
or U16448 (N_16448,N_14951,N_14254);
nand U16449 (N_16449,N_13155,N_15455);
or U16450 (N_16450,N_15263,N_13707);
or U16451 (N_16451,N_13184,N_12575);
or U16452 (N_16452,N_12803,N_12954);
nor U16453 (N_16453,N_14050,N_14792);
or U16454 (N_16454,N_14995,N_13933);
and U16455 (N_16455,N_12740,N_13817);
or U16456 (N_16456,N_15316,N_14133);
xor U16457 (N_16457,N_14482,N_13576);
xor U16458 (N_16458,N_14095,N_13363);
or U16459 (N_16459,N_13393,N_15340);
nand U16460 (N_16460,N_15027,N_15493);
or U16461 (N_16461,N_13464,N_13001);
and U16462 (N_16462,N_13683,N_13756);
or U16463 (N_16463,N_13539,N_14358);
nand U16464 (N_16464,N_13252,N_15020);
xor U16465 (N_16465,N_14478,N_13170);
nand U16466 (N_16466,N_15181,N_15222);
and U16467 (N_16467,N_13794,N_14535);
or U16468 (N_16468,N_15059,N_14902);
and U16469 (N_16469,N_14303,N_15363);
xnor U16470 (N_16470,N_15575,N_15145);
xor U16471 (N_16471,N_12812,N_13500);
or U16472 (N_16472,N_14112,N_14157);
nand U16473 (N_16473,N_13355,N_12922);
and U16474 (N_16474,N_14929,N_13283);
or U16475 (N_16475,N_15466,N_15369);
nor U16476 (N_16476,N_15034,N_13407);
nand U16477 (N_16477,N_14505,N_15548);
or U16478 (N_16478,N_13019,N_12525);
and U16479 (N_16479,N_14104,N_14682);
or U16480 (N_16480,N_15179,N_15286);
xnor U16481 (N_16481,N_12747,N_14852);
xnor U16482 (N_16482,N_14830,N_15550);
nand U16483 (N_16483,N_12918,N_15156);
nor U16484 (N_16484,N_15279,N_13832);
nor U16485 (N_16485,N_14217,N_13208);
nor U16486 (N_16486,N_15253,N_13202);
nor U16487 (N_16487,N_13035,N_12563);
and U16488 (N_16488,N_14497,N_13743);
xor U16489 (N_16489,N_15251,N_14825);
or U16490 (N_16490,N_14752,N_13323);
and U16491 (N_16491,N_15442,N_13179);
nand U16492 (N_16492,N_14918,N_14757);
nor U16493 (N_16493,N_13805,N_14031);
xnor U16494 (N_16494,N_12770,N_13149);
xnor U16495 (N_16495,N_14654,N_12688);
or U16496 (N_16496,N_13738,N_14720);
and U16497 (N_16497,N_15191,N_14410);
nor U16498 (N_16498,N_14917,N_13977);
nor U16499 (N_16499,N_14427,N_13629);
nor U16500 (N_16500,N_13909,N_14703);
nor U16501 (N_16501,N_15414,N_14667);
and U16502 (N_16502,N_14856,N_14115);
or U16503 (N_16503,N_14873,N_13626);
nor U16504 (N_16504,N_14602,N_15270);
nor U16505 (N_16505,N_12607,N_14156);
xor U16506 (N_16506,N_15392,N_15447);
nor U16507 (N_16507,N_13468,N_13489);
nand U16508 (N_16508,N_14117,N_12837);
xor U16509 (N_16509,N_14493,N_13535);
nand U16510 (N_16510,N_13159,N_13466);
or U16511 (N_16511,N_13152,N_15075);
and U16512 (N_16512,N_15141,N_13607);
nand U16513 (N_16513,N_13979,N_13173);
nand U16514 (N_16514,N_13369,N_13733);
xor U16515 (N_16515,N_13126,N_13087);
and U16516 (N_16516,N_13578,N_14420);
xnor U16517 (N_16517,N_14521,N_12583);
nand U16518 (N_16518,N_14599,N_13243);
nor U16519 (N_16519,N_15477,N_15334);
nor U16520 (N_16520,N_14181,N_13870);
nor U16521 (N_16521,N_12776,N_14287);
nor U16522 (N_16522,N_13569,N_13164);
nand U16523 (N_16523,N_14289,N_13680);
or U16524 (N_16524,N_14215,N_13679);
and U16525 (N_16525,N_12807,N_15530);
xor U16526 (N_16526,N_13661,N_12625);
or U16527 (N_16527,N_12735,N_13898);
and U16528 (N_16528,N_13657,N_13281);
nor U16529 (N_16529,N_12757,N_12998);
or U16530 (N_16530,N_13709,N_14648);
xor U16531 (N_16531,N_14849,N_15257);
and U16532 (N_16532,N_13853,N_13934);
or U16533 (N_16533,N_13073,N_14203);
nor U16534 (N_16534,N_13237,N_15189);
or U16535 (N_16535,N_14184,N_14838);
or U16536 (N_16536,N_14341,N_13400);
nand U16537 (N_16537,N_13230,N_13451);
or U16538 (N_16538,N_14278,N_15124);
nand U16539 (N_16539,N_14408,N_14023);
nand U16540 (N_16540,N_15177,N_13754);
or U16541 (N_16541,N_12697,N_14285);
nor U16542 (N_16542,N_13121,N_13715);
and U16543 (N_16543,N_14833,N_13821);
and U16544 (N_16544,N_15565,N_12875);
xor U16545 (N_16545,N_13312,N_15148);
nor U16546 (N_16546,N_14301,N_12956);
nand U16547 (N_16547,N_12635,N_14383);
nand U16548 (N_16548,N_13321,N_12796);
nand U16549 (N_16549,N_15090,N_12978);
and U16550 (N_16550,N_14858,N_13775);
nand U16551 (N_16551,N_12503,N_14452);
xnor U16552 (N_16552,N_14538,N_14381);
nand U16553 (N_16553,N_14699,N_12538);
and U16554 (N_16554,N_14221,N_13668);
nor U16555 (N_16555,N_14650,N_12522);
and U16556 (N_16556,N_13643,N_15307);
nor U16557 (N_16557,N_13922,N_13698);
xor U16558 (N_16558,N_15214,N_15019);
xnor U16559 (N_16559,N_15095,N_14053);
nand U16560 (N_16560,N_15359,N_14252);
and U16561 (N_16561,N_14003,N_13241);
nor U16562 (N_16562,N_13759,N_15134);
xor U16563 (N_16563,N_12618,N_14315);
or U16564 (N_16564,N_14895,N_14678);
nor U16565 (N_16565,N_13602,N_13010);
or U16566 (N_16566,N_13294,N_14042);
or U16567 (N_16567,N_15066,N_12723);
and U16568 (N_16568,N_14132,N_14353);
or U16569 (N_16569,N_13109,N_12532);
or U16570 (N_16570,N_13514,N_14070);
xor U16571 (N_16571,N_14557,N_12676);
and U16572 (N_16572,N_15294,N_12533);
and U16573 (N_16573,N_15079,N_14169);
nor U16574 (N_16574,N_13472,N_12890);
nand U16575 (N_16575,N_13557,N_13326);
nor U16576 (N_16576,N_14103,N_13623);
and U16577 (N_16577,N_14683,N_15564);
nand U16578 (N_16578,N_15538,N_15137);
or U16579 (N_16579,N_12872,N_15039);
nor U16580 (N_16580,N_13612,N_13609);
nor U16581 (N_16581,N_13270,N_14274);
and U16582 (N_16582,N_13452,N_13552);
or U16583 (N_16583,N_13061,N_13330);
xnor U16584 (N_16584,N_14038,N_14304);
and U16585 (N_16585,N_14575,N_15423);
nor U16586 (N_16586,N_14362,N_13758);
and U16587 (N_16587,N_15542,N_13646);
and U16588 (N_16588,N_13835,N_14783);
nand U16589 (N_16589,N_13517,N_13907);
nand U16590 (N_16590,N_13531,N_15024);
nor U16591 (N_16591,N_14561,N_14020);
nor U16592 (N_16592,N_13880,N_12806);
nor U16593 (N_16593,N_14028,N_14240);
or U16594 (N_16594,N_13120,N_14689);
nor U16595 (N_16595,N_12981,N_13994);
or U16596 (N_16596,N_13260,N_12856);
or U16597 (N_16597,N_15018,N_14266);
nand U16598 (N_16598,N_15350,N_13228);
xor U16599 (N_16599,N_15078,N_13549);
nor U16600 (N_16600,N_14355,N_13530);
nand U16601 (N_16601,N_12762,N_15337);
nor U16602 (N_16602,N_14439,N_12983);
xor U16603 (N_16603,N_12953,N_13432);
xor U16604 (N_16604,N_12932,N_13796);
nand U16605 (N_16605,N_15219,N_14596);
and U16606 (N_16606,N_14764,N_12970);
nand U16607 (N_16607,N_12558,N_15045);
nor U16608 (N_16608,N_15300,N_15030);
xor U16609 (N_16609,N_14510,N_13713);
or U16610 (N_16610,N_12784,N_15312);
or U16611 (N_16611,N_13269,N_14018);
nor U16612 (N_16612,N_13291,N_12606);
and U16613 (N_16613,N_14665,N_14854);
nand U16614 (N_16614,N_14468,N_12542);
nand U16615 (N_16615,N_14249,N_15114);
xnor U16616 (N_16616,N_15385,N_13848);
and U16617 (N_16617,N_13391,N_15490);
or U16618 (N_16618,N_13337,N_15237);
and U16619 (N_16619,N_13653,N_12578);
nand U16620 (N_16620,N_15278,N_13767);
nand U16621 (N_16621,N_13219,N_15033);
and U16622 (N_16622,N_14401,N_13672);
nand U16623 (N_16623,N_13096,N_12721);
nand U16624 (N_16624,N_14284,N_13864);
nor U16625 (N_16625,N_14711,N_14655);
or U16626 (N_16626,N_14692,N_14625);
xnor U16627 (N_16627,N_14932,N_15588);
or U16628 (N_16628,N_13251,N_14870);
nand U16629 (N_16629,N_14731,N_14980);
nor U16630 (N_16630,N_12878,N_13579);
or U16631 (N_16631,N_13404,N_14097);
nor U16632 (N_16632,N_14848,N_15348);
nand U16633 (N_16633,N_13763,N_15236);
nor U16634 (N_16634,N_13458,N_15438);
or U16635 (N_16635,N_14588,N_13438);
and U16636 (N_16636,N_13277,N_15470);
nand U16637 (N_16637,N_13780,N_15122);
and U16638 (N_16638,N_14300,N_14055);
nor U16639 (N_16639,N_13812,N_13980);
or U16640 (N_16640,N_15125,N_14984);
nor U16641 (N_16641,N_14399,N_15383);
nor U16642 (N_16642,N_14771,N_13648);
nand U16643 (N_16643,N_14500,N_12907);
xor U16644 (N_16644,N_13555,N_13091);
or U16645 (N_16645,N_14717,N_12917);
nor U16646 (N_16646,N_12602,N_13156);
or U16647 (N_16647,N_12540,N_15592);
or U16648 (N_16648,N_14589,N_13592);
nor U16649 (N_16649,N_15403,N_15449);
nor U16650 (N_16650,N_13204,N_12627);
or U16651 (N_16651,N_14170,N_13308);
nor U16652 (N_16652,N_12730,N_12632);
and U16653 (N_16653,N_14041,N_13414);
nand U16654 (N_16654,N_14758,N_14237);
or U16655 (N_16655,N_14794,N_14587);
and U16656 (N_16656,N_12864,N_13546);
nand U16657 (N_16657,N_14942,N_13039);
xor U16658 (N_16658,N_14277,N_13766);
or U16659 (N_16659,N_13240,N_14267);
or U16660 (N_16660,N_14810,N_13806);
nor U16661 (N_16661,N_13137,N_14297);
and U16662 (N_16662,N_13810,N_15459);
or U16663 (N_16663,N_14251,N_13896);
or U16664 (N_16664,N_14732,N_13908);
nand U16665 (N_16665,N_14422,N_12857);
nor U16666 (N_16666,N_14185,N_14986);
and U16667 (N_16667,N_12761,N_13119);
and U16668 (N_16668,N_12883,N_13287);
or U16669 (N_16669,N_12758,N_14001);
nand U16670 (N_16670,N_13693,N_13375);
nor U16671 (N_16671,N_13425,N_15241);
nand U16672 (N_16672,N_13469,N_14919);
nor U16673 (N_16673,N_15407,N_12894);
nor U16674 (N_16674,N_12520,N_12692);
nand U16675 (N_16675,N_14033,N_13731);
or U16676 (N_16676,N_15068,N_12889);
nor U16677 (N_16677,N_12854,N_14710);
and U16678 (N_16678,N_15101,N_14236);
and U16679 (N_16679,N_13314,N_14677);
and U16680 (N_16680,N_13215,N_14550);
and U16681 (N_16681,N_14190,N_13635);
and U16682 (N_16682,N_13721,N_13288);
or U16683 (N_16683,N_13797,N_12561);
nor U16684 (N_16684,N_12882,N_14273);
or U16685 (N_16685,N_14178,N_15537);
or U16686 (N_16686,N_15113,N_13915);
nor U16687 (N_16687,N_13834,N_12674);
or U16688 (N_16688,N_13082,N_13967);
and U16689 (N_16689,N_15445,N_15014);
nand U16690 (N_16690,N_15568,N_13379);
nor U16691 (N_16691,N_14238,N_12793);
nand U16692 (N_16692,N_14385,N_13947);
nand U16693 (N_16693,N_14724,N_15522);
xnor U16694 (N_16694,N_15115,N_13317);
and U16695 (N_16695,N_12861,N_15397);
nand U16696 (N_16696,N_14708,N_15011);
or U16697 (N_16697,N_13331,N_13773);
or U16698 (N_16698,N_14555,N_14321);
nor U16699 (N_16699,N_15539,N_14930);
nand U16700 (N_16700,N_13372,N_15341);
or U16701 (N_16701,N_12926,N_14622);
or U16702 (N_16702,N_13822,N_12663);
nor U16703 (N_16703,N_15460,N_13826);
and U16704 (N_16704,N_14209,N_12840);
nand U16705 (N_16705,N_14921,N_13342);
or U16706 (N_16706,N_14914,N_13364);
and U16707 (N_16707,N_15320,N_15560);
or U16708 (N_16708,N_12834,N_12786);
or U16709 (N_16709,N_14361,N_12518);
and U16710 (N_16710,N_13819,N_14078);
and U16711 (N_16711,N_13505,N_13180);
nand U16712 (N_16712,N_13841,N_15275);
or U16713 (N_16713,N_15399,N_13886);
nor U16714 (N_16714,N_14880,N_15505);
xor U16715 (N_16715,N_15315,N_12897);
and U16716 (N_16716,N_15586,N_15404);
nand U16717 (N_16717,N_14834,N_14029);
nand U16718 (N_16718,N_14125,N_13877);
or U16719 (N_16719,N_13476,N_12860);
nand U16720 (N_16720,N_15190,N_15067);
nand U16721 (N_16721,N_15416,N_15176);
nor U16722 (N_16722,N_13972,N_13868);
or U16723 (N_16723,N_15017,N_15269);
nor U16724 (N_16724,N_14035,N_12668);
and U16725 (N_16725,N_14434,N_15553);
nand U16726 (N_16726,N_15356,N_13723);
or U16727 (N_16727,N_14312,N_12666);
and U16728 (N_16728,N_12765,N_14246);
nor U16729 (N_16729,N_13161,N_13431);
nand U16730 (N_16730,N_13386,N_15211);
nor U16731 (N_16731,N_12549,N_14894);
nor U16732 (N_16732,N_13265,N_13146);
or U16733 (N_16733,N_12501,N_13028);
and U16734 (N_16734,N_13059,N_14987);
nor U16735 (N_16735,N_14390,N_14621);
or U16736 (N_16736,N_14483,N_12831);
or U16737 (N_16737,N_15574,N_14378);
or U16738 (N_16738,N_15412,N_14461);
and U16739 (N_16739,N_13113,N_12909);
nand U16740 (N_16740,N_15313,N_15327);
nor U16741 (N_16741,N_13132,N_12802);
nand U16742 (N_16742,N_14057,N_14197);
and U16743 (N_16743,N_12511,N_14173);
nor U16744 (N_16744,N_14813,N_15595);
xor U16745 (N_16745,N_13842,N_14869);
nand U16746 (N_16746,N_13248,N_14082);
nand U16747 (N_16747,N_13223,N_15602);
nor U16748 (N_16748,N_14928,N_15480);
nor U16749 (N_16749,N_14294,N_14586);
nor U16750 (N_16750,N_15215,N_14709);
xor U16751 (N_16751,N_14025,N_13937);
or U16752 (N_16752,N_12915,N_13547);
xor U16753 (N_16753,N_13523,N_13611);
xnor U16754 (N_16754,N_15098,N_14837);
nor U16755 (N_16755,N_13582,N_13382);
nand U16756 (N_16756,N_14242,N_15483);
or U16757 (N_16757,N_12643,N_13800);
nand U16758 (N_16758,N_14903,N_15555);
xor U16759 (N_16759,N_12925,N_13267);
nand U16760 (N_16760,N_13701,N_15022);
and U16761 (N_16761,N_14058,N_12855);
and U16762 (N_16762,N_13687,N_14165);
nor U16763 (N_16763,N_13442,N_15121);
nand U16764 (N_16764,N_12999,N_13684);
nand U16765 (N_16765,N_12670,N_14396);
or U16766 (N_16766,N_13097,N_14700);
nor U16767 (N_16767,N_13385,N_13904);
or U16768 (N_16768,N_14421,N_13634);
nor U16769 (N_16769,N_14475,N_14114);
nand U16770 (N_16770,N_13789,N_15175);
or U16771 (N_16771,N_13971,N_15611);
nor U16772 (N_16772,N_13197,N_13011);
and U16773 (N_16773,N_15552,N_12822);
nand U16774 (N_16774,N_13777,N_12958);
or U16775 (N_16775,N_13433,N_15365);
and U16776 (N_16776,N_13324,N_14637);
and U16777 (N_16777,N_14270,N_14442);
nand U16778 (N_16778,N_13816,N_14367);
and U16779 (N_16779,N_14205,N_15301);
and U16780 (N_16780,N_15225,N_13181);
xnor U16781 (N_16781,N_15422,N_12944);
nand U16782 (N_16782,N_13444,N_15581);
or U16783 (N_16783,N_14567,N_13136);
nor U16784 (N_16784,N_14027,N_14960);
nand U16785 (N_16785,N_13891,N_15103);
or U16786 (N_16786,N_15451,N_14380);
or U16787 (N_16787,N_13993,N_14247);
or U16788 (N_16788,N_14154,N_14124);
xor U16789 (N_16789,N_14372,N_13172);
nand U16790 (N_16790,N_15232,N_13567);
or U16791 (N_16791,N_14800,N_15094);
nand U16792 (N_16792,N_13378,N_14374);
nor U16793 (N_16793,N_12781,N_13615);
nand U16794 (N_16794,N_15545,N_15469);
and U16795 (N_16795,N_13182,N_13153);
nor U16796 (N_16796,N_12923,N_14566);
nor U16797 (N_16797,N_13512,N_15317);
or U16798 (N_16798,N_14155,N_14065);
nand U16799 (N_16799,N_13892,N_14723);
or U16800 (N_16800,N_14855,N_15396);
or U16801 (N_16801,N_12603,N_12708);
nor U16802 (N_16802,N_13494,N_15347);
xor U16803 (N_16803,N_15226,N_14952);
nand U16804 (N_16804,N_13630,N_13920);
and U16805 (N_16805,N_13090,N_14327);
nand U16806 (N_16806,N_15081,N_13564);
nand U16807 (N_16807,N_12841,N_12908);
and U16808 (N_16808,N_15454,N_12609);
xnor U16809 (N_16809,N_13067,N_15495);
nor U16810 (N_16810,N_14983,N_13307);
and U16811 (N_16811,N_13587,N_15437);
or U16812 (N_16812,N_14955,N_14271);
and U16813 (N_16813,N_14926,N_13900);
nand U16814 (N_16814,N_14232,N_14946);
nor U16815 (N_16815,N_15471,N_13099);
and U16816 (N_16816,N_13443,N_13320);
nand U16817 (N_16817,N_15249,N_14885);
xnor U16818 (N_16818,N_15335,N_15536);
and U16819 (N_16819,N_12527,N_13885);
xor U16820 (N_16820,N_14912,N_12982);
nand U16821 (N_16821,N_14861,N_14862);
nor U16822 (N_16822,N_15151,N_12773);
or U16823 (N_16823,N_13940,N_15617);
xnor U16824 (N_16824,N_14179,N_15411);
and U16825 (N_16825,N_14416,N_14868);
nor U16826 (N_16826,N_12729,N_14192);
and U16827 (N_16827,N_14076,N_12605);
nor U16828 (N_16828,N_14227,N_12564);
nand U16829 (N_16829,N_14606,N_14343);
and U16830 (N_16830,N_15276,N_13625);
nand U16831 (N_16831,N_12760,N_15418);
nand U16832 (N_16832,N_14516,N_14934);
nand U16833 (N_16833,N_12863,N_14807);
xnor U16834 (N_16834,N_15165,N_13728);
xnor U16835 (N_16835,N_13642,N_13362);
or U16836 (N_16836,N_15498,N_12593);
or U16837 (N_16837,N_15608,N_14062);
or U16838 (N_16838,N_15384,N_15267);
nand U16839 (N_16839,N_12649,N_12724);
nor U16840 (N_16840,N_13957,N_15503);
nor U16841 (N_16841,N_14988,N_13117);
xor U16842 (N_16842,N_14736,N_15150);
or U16843 (N_16843,N_15202,N_14553);
nor U16844 (N_16844,N_15618,N_14742);
and U16845 (N_16845,N_14626,N_15355);
or U16846 (N_16846,N_14743,N_14161);
nor U16847 (N_16847,N_12502,N_13394);
xnor U16848 (N_16848,N_15109,N_15497);
xor U16849 (N_16849,N_14389,N_15583);
nand U16850 (N_16850,N_13409,N_15345);
nand U16851 (N_16851,N_14371,N_12623);
or U16852 (N_16852,N_14088,N_15187);
nor U16853 (N_16853,N_14393,N_13984);
and U16854 (N_16854,N_12636,N_13662);
nor U16855 (N_16855,N_14584,N_15513);
xnor U16856 (N_16856,N_13006,N_13599);
nor U16857 (N_16857,N_14324,N_12667);
nor U16858 (N_16858,N_14406,N_13024);
xor U16859 (N_16859,N_13545,N_13290);
nor U16860 (N_16860,N_15200,N_15475);
nor U16861 (N_16861,N_14054,N_13402);
nand U16862 (N_16862,N_13585,N_13151);
or U16863 (N_16863,N_12553,N_12951);
nand U16864 (N_16864,N_13699,N_12993);
or U16865 (N_16865,N_12751,N_13258);
nor U16866 (N_16866,N_15623,N_13396);
and U16867 (N_16867,N_13356,N_13828);
nor U16868 (N_16868,N_14888,N_13865);
nor U16869 (N_16869,N_14611,N_15374);
nand U16870 (N_16870,N_13890,N_15428);
xnor U16871 (N_16871,N_15398,N_15178);
nor U16872 (N_16872,N_15244,N_14417);
nor U16873 (N_16873,N_15256,N_13944);
and U16874 (N_16874,N_12989,N_12764);
nand U16875 (N_16875,N_14844,N_13510);
and U16876 (N_16876,N_13420,N_14776);
nor U16877 (N_16877,N_13536,N_12694);
and U16878 (N_16878,N_13543,N_12829);
nand U16879 (N_16879,N_13793,N_12996);
and U16880 (N_16880,N_14772,N_12654);
nand U16881 (N_16881,N_12783,N_13652);
nand U16882 (N_16882,N_15563,N_15118);
nor U16883 (N_16883,N_13190,N_15130);
or U16884 (N_16884,N_12819,N_14993);
or U16885 (N_16885,N_14958,N_14725);
nand U16886 (N_16886,N_13590,N_13359);
or U16887 (N_16887,N_13189,N_14299);
and U16888 (N_16888,N_15140,N_15492);
nor U16889 (N_16889,N_13655,N_14746);
and U16890 (N_16890,N_15587,N_13807);
and U16891 (N_16891,N_15379,N_13830);
or U16892 (N_16892,N_15479,N_14748);
nor U16893 (N_16893,N_14049,N_13710);
or U16894 (N_16894,N_15271,N_14636);
nor U16895 (N_16895,N_13148,N_15050);
nor U16896 (N_16896,N_12939,N_14138);
nor U16897 (N_16897,N_12665,N_14886);
nand U16898 (N_16898,N_14531,N_12934);
and U16899 (N_16899,N_13309,N_14954);
or U16900 (N_16900,N_13565,N_14261);
or U16901 (N_16901,N_14680,N_14106);
nor U16902 (N_16902,N_15133,N_13064);
and U16903 (N_16903,N_15582,N_13435);
nor U16904 (N_16904,N_13974,N_13205);
and U16905 (N_16905,N_13411,N_14673);
nor U16906 (N_16906,N_14143,N_14506);
xor U16907 (N_16907,N_14146,N_13765);
nand U16908 (N_16908,N_13866,N_13903);
and U16909 (N_16909,N_14443,N_13381);
nand U16910 (N_16910,N_15323,N_14572);
nand U16911 (N_16911,N_13055,N_14130);
or U16912 (N_16912,N_13481,N_14560);
nor U16913 (N_16913,N_15606,N_13962);
xor U16914 (N_16914,N_13720,N_14084);
nand U16915 (N_16915,N_13014,N_13742);
and U16916 (N_16916,N_15322,N_12933);
and U16917 (N_16917,N_15149,N_13666);
nor U16918 (N_16918,N_15464,N_15157);
and U16919 (N_16919,N_12794,N_15509);
xor U16920 (N_16920,N_15072,N_13084);
nor U16921 (N_16921,N_13134,N_14359);
and U16922 (N_16922,N_14044,N_14148);
nand U16923 (N_16923,N_15580,N_15472);
and U16924 (N_16924,N_14269,N_15036);
xor U16925 (N_16925,N_13026,N_13253);
or U16926 (N_16926,N_13752,N_14288);
nand U16927 (N_16927,N_14899,N_12726);
nor U16928 (N_16928,N_13304,N_13416);
nand U16929 (N_16929,N_13676,N_15360);
nand U16930 (N_16930,N_13956,N_15533);
nor U16931 (N_16931,N_12628,N_13855);
or U16932 (N_16932,N_13818,N_15577);
nor U16933 (N_16933,N_13650,N_13076);
nor U16934 (N_16934,N_13771,N_15102);
or U16935 (N_16935,N_13950,N_12877);
and U16936 (N_16936,N_13074,N_14424);
nor U16937 (N_16937,N_14459,N_13851);
or U16938 (N_16938,N_14101,N_13955);
nor U16939 (N_16939,N_13429,N_13689);
nand U16940 (N_16940,N_13325,N_12741);
and U16941 (N_16941,N_13527,N_14188);
and U16942 (N_16942,N_13235,N_12739);
nand U16943 (N_16943,N_15342,N_14469);
xnor U16944 (N_16944,N_15376,N_13620);
nand U16945 (N_16945,N_15540,N_14714);
nand U16946 (N_16946,N_14336,N_12942);
xnor U16947 (N_16947,N_13788,N_13577);
or U16948 (N_16948,N_15615,N_13043);
nor U16949 (N_16949,N_13926,N_12574);
and U16950 (N_16950,N_12859,N_13100);
and U16951 (N_16951,N_13618,N_12769);
or U16952 (N_16952,N_15288,N_12529);
nor U16953 (N_16953,N_14074,N_13169);
nand U16954 (N_16954,N_15230,N_13528);
and U16955 (N_16955,N_13973,N_14949);
xnor U16956 (N_16956,N_15554,N_13210);
nand U16957 (N_16957,N_13912,N_13408);
xnor U16958 (N_16958,N_13031,N_14109);
nand U16959 (N_16959,N_13969,N_15579);
nor U16960 (N_16960,N_15002,N_14013);
nand U16961 (N_16961,N_12826,N_13025);
or U16962 (N_16962,N_14507,N_15218);
or U16963 (N_16963,N_12595,N_12775);
and U16964 (N_16964,N_13498,N_12645);
or U16965 (N_16965,N_15186,N_14135);
nand U16966 (N_16966,N_13150,N_14747);
nor U16967 (N_16967,N_15326,N_13911);
and U16968 (N_16968,N_14818,N_13220);
or U16969 (N_16969,N_13958,N_14248);
and U16970 (N_16970,N_13823,N_14425);
nor U16971 (N_16971,N_13305,N_13292);
nor U16972 (N_16972,N_15558,N_13905);
xnor U16973 (N_16973,N_14313,N_14200);
nor U16974 (N_16974,N_14937,N_14451);
nand U16975 (N_16975,N_14064,N_15292);
and U16976 (N_16976,N_14745,N_12876);
nor U16977 (N_16977,N_14749,N_13042);
nor U16978 (N_16978,N_14099,N_14816);
and U16979 (N_16979,N_15040,N_13441);
and U16980 (N_16980,N_15590,N_14397);
or U16981 (N_16981,N_14298,N_13264);
nor U16982 (N_16982,N_13667,N_14296);
and U16983 (N_16983,N_15182,N_13282);
or U16984 (N_16984,N_15620,N_14766);
or U16985 (N_16985,N_15062,N_12979);
and U16986 (N_16986,N_14878,N_14489);
nor U16987 (N_16987,N_13559,N_12651);
nand U16988 (N_16988,N_14317,N_12904);
and U16989 (N_16989,N_12544,N_13334);
nor U16990 (N_16990,N_12562,N_12571);
nor U16991 (N_16991,N_13371,N_12992);
or U16992 (N_16992,N_12858,N_15517);
nor U16993 (N_16993,N_14127,N_13424);
nor U16994 (N_16994,N_14875,N_14211);
and U16995 (N_16995,N_13878,N_13221);
nor U16996 (N_16996,N_14241,N_14945);
or U16997 (N_16997,N_13114,N_13302);
or U16998 (N_16998,N_13186,N_14086);
nand U16999 (N_16999,N_13808,N_13507);
and U17000 (N_17000,N_13368,N_13803);
xnor U17001 (N_17001,N_13065,N_12722);
nor U17002 (N_17002,N_15196,N_15262);
nor U17003 (N_17003,N_15446,N_12771);
nor U17004 (N_17004,N_12737,N_14429);
nor U17005 (N_17005,N_13897,N_13068);
nand U17006 (N_17006,N_15108,N_13392);
nand U17007 (N_17007,N_13183,N_15598);
or U17008 (N_17008,N_14292,N_12661);
nand U17009 (N_17009,N_12725,N_13815);
nand U17010 (N_17010,N_14040,N_15235);
nor U17011 (N_17011,N_12866,N_13589);
nand U17012 (N_17012,N_15119,N_14172);
and U17013 (N_17013,N_14437,N_13122);
nor U17014 (N_17014,N_14690,N_14527);
or U17015 (N_17015,N_15131,N_12787);
xnor U17016 (N_17016,N_13009,N_15198);
xor U17017 (N_17017,N_12736,N_13198);
or U17018 (N_17018,N_13954,N_13256);
and U17019 (N_17019,N_13049,N_12545);
and U17020 (N_17020,N_14821,N_14149);
or U17021 (N_17021,N_14607,N_13658);
or U17022 (N_17022,N_13591,N_12843);
or U17023 (N_17023,N_14002,N_14698);
nor U17024 (N_17024,N_14755,N_15484);
and U17025 (N_17025,N_15221,N_13671);
or U17026 (N_17026,N_13040,N_13700);
xor U17027 (N_17027,N_14843,N_12675);
nand U17028 (N_17028,N_14573,N_14060);
nand U17029 (N_17029,N_12656,N_12528);
and U17030 (N_17030,N_13606,N_14769);
nor U17031 (N_17031,N_14590,N_13477);
nand U17032 (N_17032,N_14841,N_13350);
nor U17033 (N_17033,N_12895,N_15370);
nand U17034 (N_17034,N_15088,N_14418);
or U17035 (N_17035,N_13021,N_12886);
nand U17036 (N_17036,N_12597,N_14005);
xnor U17037 (N_17037,N_14357,N_14073);
xnor U17038 (N_17038,N_15161,N_13095);
nand U17039 (N_17039,N_15309,N_14513);
or U17040 (N_17040,N_13041,N_13335);
nand U17041 (N_17041,N_14226,N_14504);
and U17042 (N_17042,N_13044,N_14280);
or U17043 (N_17043,N_15143,N_14803);
nor U17044 (N_17044,N_14629,N_14039);
or U17045 (N_17045,N_13272,N_15339);
nor U17046 (N_17046,N_15049,N_13225);
and U17047 (N_17047,N_14259,N_14514);
xnor U17048 (N_17048,N_13029,N_15371);
and U17049 (N_17049,N_15074,N_13995);
or U17050 (N_17050,N_14494,N_12614);
xnor U17051 (N_17051,N_13895,N_13537);
nor U17052 (N_17052,N_13556,N_12686);
or U17053 (N_17053,N_14660,N_13361);
or U17054 (N_17054,N_14191,N_15458);
or U17055 (N_17055,N_13581,N_13554);
or U17056 (N_17056,N_12521,N_15415);
nor U17057 (N_17057,N_12594,N_14253);
nor U17058 (N_17058,N_14398,N_14695);
and U17059 (N_17059,N_14674,N_14592);
nor U17060 (N_17060,N_13332,N_13935);
xor U17061 (N_17061,N_13563,N_14255);
nor U17062 (N_17062,N_13991,N_14623);
or U17063 (N_17063,N_12695,N_13128);
or U17064 (N_17064,N_14473,N_14761);
or U17065 (N_17065,N_13551,N_14000);
and U17066 (N_17066,N_13131,N_12928);
and U17067 (N_17067,N_15329,N_12949);
nor U17068 (N_17068,N_13080,N_14176);
nor U17069 (N_17069,N_13484,N_15380);
nand U17070 (N_17070,N_14319,N_13516);
nand U17071 (N_17071,N_13107,N_13249);
nor U17072 (N_17072,N_12809,N_14412);
or U17073 (N_17073,N_13501,N_12580);
nor U17074 (N_17074,N_13083,N_15585);
xnor U17075 (N_17075,N_15003,N_13596);
nand U17076 (N_17076,N_14997,N_14111);
nor U17077 (N_17077,N_15166,N_12818);
or U17078 (N_17078,N_15009,N_13275);
nand U17079 (N_17079,N_12941,N_14423);
nand U17080 (N_17080,N_13242,N_15426);
or U17081 (N_17081,N_14283,N_14388);
nor U17082 (N_17082,N_13346,N_14043);
nand U17083 (N_17083,N_14767,N_13631);
nand U17084 (N_17084,N_14121,N_14542);
nor U17085 (N_17085,N_13175,N_15205);
nand U17086 (N_17086,N_14032,N_12919);
nand U17087 (N_17087,N_12801,N_14863);
nand U17088 (N_17088,N_13079,N_15311);
nand U17089 (N_17089,N_13141,N_13692);
and U17090 (N_17090,N_12510,N_14593);
nor U17091 (N_17091,N_12853,N_12788);
and U17092 (N_17092,N_12734,N_14529);
and U17093 (N_17093,N_15132,N_15199);
and U17094 (N_17094,N_12591,N_14349);
nor U17095 (N_17095,N_13799,N_13377);
or U17096 (N_17096,N_15192,N_13297);
xnor U17097 (N_17097,N_12711,N_12592);
nand U17098 (N_17098,N_14275,N_12586);
nand U17099 (N_17099,N_14661,N_13975);
nand U17100 (N_17100,N_14206,N_14634);
or U17101 (N_17101,N_15468,N_13939);
nand U17102 (N_17102,N_12948,N_14799);
or U17103 (N_17103,N_15174,N_13327);
nand U17104 (N_17104,N_15234,N_14162);
and U17105 (N_17105,N_13640,N_13690);
nand U17106 (N_17106,N_14207,N_15599);
or U17107 (N_17107,N_13310,N_12990);
nand U17108 (N_17108,N_14635,N_14670);
or U17109 (N_17109,N_15213,N_15048);
or U17110 (N_17110,N_13254,N_13910);
nand U17111 (N_17111,N_13486,N_15243);
or U17112 (N_17112,N_15388,N_14977);
nor U17113 (N_17113,N_12827,N_14394);
nand U17114 (N_17114,N_14419,N_15362);
nand U17115 (N_17115,N_13704,N_14812);
and U17116 (N_17116,N_14851,N_13784);
nor U17117 (N_17117,N_15092,N_12896);
or U17118 (N_17118,N_15116,N_15120);
or U17119 (N_17119,N_14796,N_13513);
and U17120 (N_17120,N_12589,N_15614);
nor U17121 (N_17121,N_13906,N_12552);
nor U17122 (N_17122,N_14559,N_13370);
or U17123 (N_17123,N_12633,N_13389);
xnor U17124 (N_17124,N_14187,N_12707);
and U17125 (N_17125,N_14706,N_14365);
nor U17126 (N_17126,N_14171,N_15135);
xor U17127 (N_17127,N_14373,N_15520);
nand U17128 (N_17128,N_12642,N_14234);
or U17129 (N_17129,N_15087,N_14730);
and U17130 (N_17130,N_15260,N_13919);
nor U17131 (N_17131,N_12681,N_15054);
and U17132 (N_17132,N_13144,N_14392);
nor U17133 (N_17133,N_14087,N_12850);
or U17134 (N_17134,N_14633,N_13395);
nor U17135 (N_17135,N_12823,N_14651);
or U17136 (N_17136,N_13448,N_13262);
nand U17137 (N_17137,N_14094,N_14376);
or U17138 (N_17138,N_13298,N_14233);
nand U17139 (N_17139,N_13669,N_13125);
nand U17140 (N_17140,N_12814,N_14591);
nor U17141 (N_17141,N_13426,N_12891);
and U17142 (N_17142,N_14356,N_15413);
or U17143 (N_17143,N_13647,N_14565);
nand U17144 (N_17144,N_14501,N_15344);
or U17145 (N_17145,N_13857,N_14477);
xor U17146 (N_17146,N_13293,N_13660);
and U17147 (N_17147,N_13139,N_15155);
nand U17148 (N_17148,N_14824,N_12745);
nor U17149 (N_17149,N_14707,N_14276);
and U17150 (N_17150,N_14351,N_14071);
or U17151 (N_17151,N_15293,N_14059);
nand U17152 (N_17152,N_14788,N_14006);
nor U17153 (N_17153,N_15452,N_14352);
nand U17154 (N_17154,N_14152,N_14212);
nand U17155 (N_17155,N_14522,N_12824);
nand U17156 (N_17156,N_13135,N_12568);
and U17157 (N_17157,N_14153,N_12693);
and U17158 (N_17158,N_14244,N_15391);
nor U17159 (N_17159,N_13814,N_14464);
or U17160 (N_17160,N_13862,N_14597);
nor U17161 (N_17161,N_13622,N_15482);
and U17162 (N_17162,N_12755,N_14907);
or U17163 (N_17163,N_14159,N_13770);
nor U17164 (N_17164,N_13115,N_13553);
nand U17165 (N_17165,N_12836,N_13160);
and U17166 (N_17166,N_14384,N_14867);
or U17167 (N_17167,N_12888,N_12548);
nor U17168 (N_17168,N_15117,N_14822);
nand U17169 (N_17169,N_14579,N_15496);
nor U17170 (N_17170,N_15557,N_12626);
nor U17171 (N_17171,N_15353,N_14576);
or U17172 (N_17172,N_14441,N_15534);
nor U17173 (N_17173,N_14484,N_14652);
or U17174 (N_17174,N_14098,N_15551);
nand U17175 (N_17175,N_13154,N_12640);
nand U17176 (N_17176,N_12701,N_15521);
or U17177 (N_17177,N_13212,N_14467);
nand U17178 (N_17178,N_14884,N_13734);
and U17179 (N_17179,N_12851,N_14310);
and U17180 (N_17180,N_13286,N_13616);
nand U17181 (N_17181,N_14911,N_15172);
nand U17182 (N_17182,N_15328,N_14865);
xnor U17183 (N_17183,N_14910,N_14595);
nor U17184 (N_17184,N_12565,N_14996);
and U17185 (N_17185,N_13696,N_14329);
nor U17186 (N_17186,N_14657,N_12911);
or U17187 (N_17187,N_13753,N_12885);
and U17188 (N_17188,N_12593,N_14088);
nor U17189 (N_17189,N_13255,N_13797);
or U17190 (N_17190,N_13989,N_14142);
or U17191 (N_17191,N_12657,N_12915);
xnor U17192 (N_17192,N_14797,N_13717);
nand U17193 (N_17193,N_14157,N_13613);
nand U17194 (N_17194,N_14245,N_13628);
nor U17195 (N_17195,N_12594,N_13378);
and U17196 (N_17196,N_15031,N_14458);
xnor U17197 (N_17197,N_13805,N_14101);
nand U17198 (N_17198,N_13391,N_14790);
nor U17199 (N_17199,N_13377,N_12960);
or U17200 (N_17200,N_12551,N_14944);
nand U17201 (N_17201,N_12540,N_14909);
xnor U17202 (N_17202,N_14067,N_14063);
nor U17203 (N_17203,N_14517,N_15091);
nor U17204 (N_17204,N_13777,N_13489);
nand U17205 (N_17205,N_13321,N_15438);
and U17206 (N_17206,N_13287,N_13548);
nand U17207 (N_17207,N_13136,N_12739);
and U17208 (N_17208,N_13333,N_14646);
nand U17209 (N_17209,N_13531,N_13044);
nor U17210 (N_17210,N_13227,N_15197);
nor U17211 (N_17211,N_12739,N_15427);
and U17212 (N_17212,N_14800,N_14411);
nand U17213 (N_17213,N_13254,N_13651);
nor U17214 (N_17214,N_12538,N_14646);
nor U17215 (N_17215,N_12684,N_15310);
and U17216 (N_17216,N_13521,N_15394);
and U17217 (N_17217,N_13346,N_13951);
or U17218 (N_17218,N_13785,N_15303);
and U17219 (N_17219,N_15019,N_12795);
and U17220 (N_17220,N_14616,N_12707);
and U17221 (N_17221,N_14232,N_14879);
and U17222 (N_17222,N_15565,N_14707);
and U17223 (N_17223,N_14283,N_13882);
or U17224 (N_17224,N_13872,N_13778);
and U17225 (N_17225,N_12982,N_15552);
and U17226 (N_17226,N_12733,N_13506);
nor U17227 (N_17227,N_14708,N_15084);
and U17228 (N_17228,N_14587,N_15518);
xor U17229 (N_17229,N_13637,N_13242);
or U17230 (N_17230,N_14233,N_14156);
or U17231 (N_17231,N_15591,N_14125);
nand U17232 (N_17232,N_13089,N_15499);
or U17233 (N_17233,N_14401,N_14593);
nand U17234 (N_17234,N_14437,N_14287);
nand U17235 (N_17235,N_15493,N_15005);
nand U17236 (N_17236,N_14903,N_13827);
nand U17237 (N_17237,N_13064,N_13684);
nand U17238 (N_17238,N_13892,N_14664);
or U17239 (N_17239,N_13507,N_14705);
nor U17240 (N_17240,N_13082,N_13317);
nor U17241 (N_17241,N_13720,N_14410);
or U17242 (N_17242,N_14639,N_14655);
and U17243 (N_17243,N_15119,N_13946);
or U17244 (N_17244,N_14779,N_13738);
and U17245 (N_17245,N_15029,N_14967);
or U17246 (N_17246,N_15250,N_15366);
xor U17247 (N_17247,N_13616,N_14057);
nor U17248 (N_17248,N_15613,N_13398);
or U17249 (N_17249,N_14598,N_14120);
or U17250 (N_17250,N_14826,N_14034);
nor U17251 (N_17251,N_14381,N_14761);
or U17252 (N_17252,N_12881,N_12535);
and U17253 (N_17253,N_12883,N_14036);
nor U17254 (N_17254,N_13915,N_13114);
nor U17255 (N_17255,N_14225,N_14430);
xor U17256 (N_17256,N_13215,N_15440);
nand U17257 (N_17257,N_13592,N_14613);
nor U17258 (N_17258,N_14594,N_14395);
or U17259 (N_17259,N_12925,N_13598);
nor U17260 (N_17260,N_14284,N_13298);
or U17261 (N_17261,N_14883,N_13169);
and U17262 (N_17262,N_13375,N_14157);
and U17263 (N_17263,N_14181,N_15274);
nand U17264 (N_17264,N_14005,N_14218);
or U17265 (N_17265,N_13316,N_13391);
nor U17266 (N_17266,N_13196,N_14639);
or U17267 (N_17267,N_12607,N_14329);
nand U17268 (N_17268,N_14156,N_14637);
nor U17269 (N_17269,N_14614,N_14378);
and U17270 (N_17270,N_14100,N_14562);
xor U17271 (N_17271,N_14494,N_15530);
or U17272 (N_17272,N_15075,N_13262);
nand U17273 (N_17273,N_15236,N_14855);
and U17274 (N_17274,N_15550,N_15228);
xnor U17275 (N_17275,N_12913,N_14346);
nand U17276 (N_17276,N_14081,N_12815);
and U17277 (N_17277,N_13682,N_14139);
nand U17278 (N_17278,N_13696,N_13165);
nand U17279 (N_17279,N_13846,N_14700);
and U17280 (N_17280,N_13870,N_14250);
or U17281 (N_17281,N_14187,N_12639);
nand U17282 (N_17282,N_15166,N_13329);
and U17283 (N_17283,N_13781,N_12673);
xor U17284 (N_17284,N_14892,N_15166);
xnor U17285 (N_17285,N_13602,N_14440);
and U17286 (N_17286,N_14038,N_14632);
and U17287 (N_17287,N_15616,N_15509);
and U17288 (N_17288,N_14461,N_14069);
and U17289 (N_17289,N_12994,N_14068);
nand U17290 (N_17290,N_13875,N_13272);
or U17291 (N_17291,N_13350,N_14007);
and U17292 (N_17292,N_12685,N_13265);
and U17293 (N_17293,N_14776,N_13323);
and U17294 (N_17294,N_15459,N_13922);
xnor U17295 (N_17295,N_12799,N_13872);
and U17296 (N_17296,N_14497,N_12870);
nor U17297 (N_17297,N_14464,N_14866);
nor U17298 (N_17298,N_13886,N_13194);
nand U17299 (N_17299,N_13157,N_13824);
or U17300 (N_17300,N_14983,N_12954);
or U17301 (N_17301,N_13010,N_15281);
nor U17302 (N_17302,N_12773,N_15093);
or U17303 (N_17303,N_15064,N_14948);
xnor U17304 (N_17304,N_14491,N_15583);
or U17305 (N_17305,N_15393,N_13421);
and U17306 (N_17306,N_15587,N_14968);
nor U17307 (N_17307,N_15051,N_14049);
nor U17308 (N_17308,N_14971,N_13994);
or U17309 (N_17309,N_13444,N_13808);
nand U17310 (N_17310,N_15318,N_12816);
xnor U17311 (N_17311,N_14717,N_13349);
nand U17312 (N_17312,N_13345,N_14579);
and U17313 (N_17313,N_14655,N_15108);
nor U17314 (N_17314,N_14481,N_14570);
or U17315 (N_17315,N_13476,N_13368);
nand U17316 (N_17316,N_14554,N_15008);
and U17317 (N_17317,N_12856,N_13827);
or U17318 (N_17318,N_13587,N_14586);
nor U17319 (N_17319,N_14861,N_14061);
nor U17320 (N_17320,N_15335,N_14156);
nand U17321 (N_17321,N_13021,N_13712);
nor U17322 (N_17322,N_14920,N_15499);
and U17323 (N_17323,N_12801,N_12589);
nand U17324 (N_17324,N_14312,N_14170);
xnor U17325 (N_17325,N_14853,N_14608);
nand U17326 (N_17326,N_13608,N_15240);
or U17327 (N_17327,N_12757,N_15445);
nor U17328 (N_17328,N_13378,N_13367);
nand U17329 (N_17329,N_13766,N_14091);
or U17330 (N_17330,N_15150,N_13994);
and U17331 (N_17331,N_13711,N_14644);
nand U17332 (N_17332,N_12670,N_13588);
nand U17333 (N_17333,N_12905,N_14535);
nor U17334 (N_17334,N_13921,N_12791);
nand U17335 (N_17335,N_13562,N_14922);
and U17336 (N_17336,N_12785,N_15311);
or U17337 (N_17337,N_12847,N_14566);
or U17338 (N_17338,N_13391,N_12529);
nand U17339 (N_17339,N_13286,N_15034);
nand U17340 (N_17340,N_12740,N_13389);
nor U17341 (N_17341,N_13673,N_14401);
nand U17342 (N_17342,N_15610,N_14552);
or U17343 (N_17343,N_13505,N_14464);
xnor U17344 (N_17344,N_13312,N_15102);
xor U17345 (N_17345,N_15085,N_13402);
nand U17346 (N_17346,N_14190,N_12723);
and U17347 (N_17347,N_13756,N_13640);
nand U17348 (N_17348,N_13450,N_13170);
xnor U17349 (N_17349,N_14958,N_13202);
xnor U17350 (N_17350,N_12730,N_13668);
or U17351 (N_17351,N_14335,N_14567);
and U17352 (N_17352,N_12850,N_12597);
or U17353 (N_17353,N_13176,N_13562);
and U17354 (N_17354,N_14562,N_15057);
xnor U17355 (N_17355,N_14599,N_14250);
xnor U17356 (N_17356,N_14914,N_15177);
xor U17357 (N_17357,N_15561,N_13180);
and U17358 (N_17358,N_13821,N_13293);
or U17359 (N_17359,N_12746,N_12683);
nand U17360 (N_17360,N_14752,N_12853);
and U17361 (N_17361,N_12742,N_12527);
or U17362 (N_17362,N_12797,N_14667);
and U17363 (N_17363,N_13822,N_13770);
nand U17364 (N_17364,N_14743,N_13692);
and U17365 (N_17365,N_15283,N_13940);
xor U17366 (N_17366,N_14058,N_13752);
xor U17367 (N_17367,N_13541,N_15569);
or U17368 (N_17368,N_15591,N_12799);
nor U17369 (N_17369,N_13301,N_12979);
or U17370 (N_17370,N_15226,N_14192);
and U17371 (N_17371,N_13458,N_15433);
or U17372 (N_17372,N_14948,N_15278);
nor U17373 (N_17373,N_14699,N_15115);
xor U17374 (N_17374,N_12675,N_15359);
nand U17375 (N_17375,N_13462,N_15472);
and U17376 (N_17376,N_13232,N_15601);
and U17377 (N_17377,N_13508,N_13284);
xor U17378 (N_17378,N_13367,N_13856);
and U17379 (N_17379,N_13391,N_14221);
nor U17380 (N_17380,N_14496,N_15205);
nand U17381 (N_17381,N_15172,N_14735);
nor U17382 (N_17382,N_13469,N_14040);
nor U17383 (N_17383,N_13168,N_14125);
or U17384 (N_17384,N_13580,N_12502);
nand U17385 (N_17385,N_13419,N_14092);
xnor U17386 (N_17386,N_15050,N_14311);
nor U17387 (N_17387,N_13605,N_14043);
xor U17388 (N_17388,N_12810,N_14692);
and U17389 (N_17389,N_15109,N_12878);
nand U17390 (N_17390,N_13100,N_14847);
nand U17391 (N_17391,N_13246,N_13334);
nand U17392 (N_17392,N_13263,N_15499);
and U17393 (N_17393,N_12640,N_14005);
or U17394 (N_17394,N_13157,N_14629);
nand U17395 (N_17395,N_14335,N_15028);
and U17396 (N_17396,N_15480,N_14489);
xnor U17397 (N_17397,N_14757,N_13804);
and U17398 (N_17398,N_13783,N_15505);
or U17399 (N_17399,N_14732,N_13195);
or U17400 (N_17400,N_13377,N_14569);
xor U17401 (N_17401,N_12867,N_13129);
nand U17402 (N_17402,N_13690,N_14018);
or U17403 (N_17403,N_13685,N_14927);
or U17404 (N_17404,N_14046,N_13371);
xnor U17405 (N_17405,N_12523,N_15151);
nand U17406 (N_17406,N_15492,N_14627);
and U17407 (N_17407,N_13829,N_14584);
or U17408 (N_17408,N_14205,N_14325);
nand U17409 (N_17409,N_14893,N_15063);
or U17410 (N_17410,N_13218,N_14883);
nand U17411 (N_17411,N_14280,N_15048);
and U17412 (N_17412,N_15601,N_14300);
nor U17413 (N_17413,N_14292,N_13371);
nor U17414 (N_17414,N_15236,N_14619);
or U17415 (N_17415,N_15487,N_15599);
nand U17416 (N_17416,N_14678,N_12672);
nor U17417 (N_17417,N_13111,N_14075);
nor U17418 (N_17418,N_13277,N_14148);
nor U17419 (N_17419,N_13388,N_12761);
nand U17420 (N_17420,N_14984,N_15380);
and U17421 (N_17421,N_15580,N_14809);
nand U17422 (N_17422,N_13839,N_13773);
nor U17423 (N_17423,N_14258,N_15133);
or U17424 (N_17424,N_14566,N_14534);
and U17425 (N_17425,N_14122,N_13625);
xnor U17426 (N_17426,N_13513,N_12953);
nor U17427 (N_17427,N_15191,N_13639);
xnor U17428 (N_17428,N_14173,N_15115);
xnor U17429 (N_17429,N_13775,N_13530);
and U17430 (N_17430,N_13818,N_15507);
nor U17431 (N_17431,N_15201,N_13433);
nor U17432 (N_17432,N_13744,N_15569);
or U17433 (N_17433,N_14422,N_14133);
and U17434 (N_17434,N_14869,N_12726);
nor U17435 (N_17435,N_15494,N_15412);
nor U17436 (N_17436,N_14136,N_15569);
nand U17437 (N_17437,N_14521,N_13478);
and U17438 (N_17438,N_13081,N_14006);
nor U17439 (N_17439,N_13680,N_14037);
nand U17440 (N_17440,N_14950,N_15500);
nand U17441 (N_17441,N_12990,N_14157);
and U17442 (N_17442,N_13538,N_13331);
and U17443 (N_17443,N_13347,N_13311);
and U17444 (N_17444,N_15309,N_13582);
xnor U17445 (N_17445,N_14398,N_13884);
nor U17446 (N_17446,N_14273,N_14749);
or U17447 (N_17447,N_15321,N_13491);
xnor U17448 (N_17448,N_12998,N_13566);
and U17449 (N_17449,N_14657,N_13322);
nand U17450 (N_17450,N_14694,N_15326);
and U17451 (N_17451,N_14561,N_15347);
xor U17452 (N_17452,N_14576,N_12652);
nand U17453 (N_17453,N_14209,N_14300);
and U17454 (N_17454,N_12552,N_13964);
and U17455 (N_17455,N_14413,N_14758);
nand U17456 (N_17456,N_13241,N_14424);
nand U17457 (N_17457,N_15538,N_13889);
or U17458 (N_17458,N_13817,N_14583);
nor U17459 (N_17459,N_13006,N_14259);
or U17460 (N_17460,N_13979,N_13111);
nand U17461 (N_17461,N_12755,N_13885);
xor U17462 (N_17462,N_12898,N_14276);
or U17463 (N_17463,N_12701,N_15078);
or U17464 (N_17464,N_12614,N_15241);
nand U17465 (N_17465,N_15457,N_12695);
or U17466 (N_17466,N_15366,N_14187);
nor U17467 (N_17467,N_15252,N_15139);
or U17468 (N_17468,N_14352,N_14094);
nand U17469 (N_17469,N_15570,N_13676);
and U17470 (N_17470,N_13607,N_14328);
nor U17471 (N_17471,N_15247,N_13912);
or U17472 (N_17472,N_13748,N_14238);
or U17473 (N_17473,N_14196,N_15001);
and U17474 (N_17474,N_12794,N_14269);
or U17475 (N_17475,N_15030,N_13515);
or U17476 (N_17476,N_15436,N_13460);
nand U17477 (N_17477,N_13292,N_13693);
and U17478 (N_17478,N_13782,N_14763);
nor U17479 (N_17479,N_13718,N_15504);
and U17480 (N_17480,N_14470,N_14293);
and U17481 (N_17481,N_13211,N_15264);
xor U17482 (N_17482,N_14517,N_14896);
and U17483 (N_17483,N_12736,N_14211);
nand U17484 (N_17484,N_14242,N_12744);
nor U17485 (N_17485,N_12654,N_15295);
and U17486 (N_17486,N_12793,N_14669);
and U17487 (N_17487,N_15228,N_13906);
nor U17488 (N_17488,N_12661,N_14047);
or U17489 (N_17489,N_15159,N_14925);
and U17490 (N_17490,N_12902,N_13208);
or U17491 (N_17491,N_15276,N_12825);
and U17492 (N_17492,N_13357,N_13257);
nor U17493 (N_17493,N_15411,N_15247);
nor U17494 (N_17494,N_14028,N_15533);
or U17495 (N_17495,N_13927,N_14937);
or U17496 (N_17496,N_15221,N_13935);
or U17497 (N_17497,N_14729,N_15419);
or U17498 (N_17498,N_12785,N_12792);
and U17499 (N_17499,N_13209,N_14818);
and U17500 (N_17500,N_14256,N_12616);
nor U17501 (N_17501,N_14770,N_13637);
nand U17502 (N_17502,N_15428,N_15272);
or U17503 (N_17503,N_15091,N_13617);
or U17504 (N_17504,N_15157,N_14103);
xor U17505 (N_17505,N_12660,N_13922);
or U17506 (N_17506,N_13771,N_14994);
nor U17507 (N_17507,N_13693,N_13289);
or U17508 (N_17508,N_14496,N_13034);
nand U17509 (N_17509,N_14923,N_14279);
and U17510 (N_17510,N_15297,N_13164);
nand U17511 (N_17511,N_15270,N_13298);
nand U17512 (N_17512,N_12712,N_15184);
or U17513 (N_17513,N_14246,N_14586);
nand U17514 (N_17514,N_15334,N_12771);
xnor U17515 (N_17515,N_13376,N_12548);
nor U17516 (N_17516,N_15108,N_15458);
or U17517 (N_17517,N_12581,N_15181);
or U17518 (N_17518,N_12795,N_14231);
or U17519 (N_17519,N_15457,N_12711);
or U17520 (N_17520,N_13867,N_14278);
or U17521 (N_17521,N_12717,N_14163);
and U17522 (N_17522,N_13256,N_12805);
nor U17523 (N_17523,N_15586,N_13025);
nand U17524 (N_17524,N_12994,N_13362);
nor U17525 (N_17525,N_15149,N_14579);
and U17526 (N_17526,N_13868,N_15606);
or U17527 (N_17527,N_12949,N_14478);
nand U17528 (N_17528,N_12998,N_15572);
nand U17529 (N_17529,N_14220,N_15479);
or U17530 (N_17530,N_15263,N_13494);
or U17531 (N_17531,N_13329,N_12995);
or U17532 (N_17532,N_13420,N_14447);
nand U17533 (N_17533,N_14788,N_13853);
xor U17534 (N_17534,N_15223,N_13560);
or U17535 (N_17535,N_15551,N_13746);
nand U17536 (N_17536,N_12811,N_15492);
and U17537 (N_17537,N_12779,N_12546);
or U17538 (N_17538,N_14592,N_15215);
or U17539 (N_17539,N_14998,N_13735);
nor U17540 (N_17540,N_12721,N_13226);
xnor U17541 (N_17541,N_14211,N_15117);
xor U17542 (N_17542,N_14377,N_13196);
and U17543 (N_17543,N_14110,N_15474);
or U17544 (N_17544,N_12849,N_13966);
nand U17545 (N_17545,N_13688,N_14891);
and U17546 (N_17546,N_12602,N_13088);
or U17547 (N_17547,N_14311,N_14972);
nor U17548 (N_17548,N_13759,N_14097);
nor U17549 (N_17549,N_15413,N_15619);
nand U17550 (N_17550,N_13166,N_15550);
nor U17551 (N_17551,N_13032,N_13344);
nor U17552 (N_17552,N_15511,N_14536);
nor U17553 (N_17553,N_13951,N_12696);
and U17554 (N_17554,N_15460,N_14378);
or U17555 (N_17555,N_14304,N_14138);
nor U17556 (N_17556,N_14163,N_12933);
and U17557 (N_17557,N_14380,N_13995);
xnor U17558 (N_17558,N_14579,N_12970);
and U17559 (N_17559,N_13026,N_13894);
or U17560 (N_17560,N_12871,N_15000);
and U17561 (N_17561,N_13746,N_13006);
nand U17562 (N_17562,N_14352,N_14458);
xor U17563 (N_17563,N_15151,N_15621);
xor U17564 (N_17564,N_15226,N_14861);
nand U17565 (N_17565,N_13137,N_14642);
nand U17566 (N_17566,N_13014,N_12813);
nor U17567 (N_17567,N_14838,N_14883);
or U17568 (N_17568,N_14013,N_14562);
nand U17569 (N_17569,N_12654,N_14843);
and U17570 (N_17570,N_13396,N_13649);
nor U17571 (N_17571,N_12656,N_12683);
nand U17572 (N_17572,N_15028,N_14093);
nor U17573 (N_17573,N_13617,N_13015);
and U17574 (N_17574,N_12769,N_13209);
or U17575 (N_17575,N_15317,N_12769);
nor U17576 (N_17576,N_12626,N_13001);
and U17577 (N_17577,N_13466,N_14610);
nand U17578 (N_17578,N_13592,N_15025);
and U17579 (N_17579,N_15537,N_14722);
and U17580 (N_17580,N_13409,N_14800);
nand U17581 (N_17581,N_13450,N_13016);
or U17582 (N_17582,N_14479,N_15228);
and U17583 (N_17583,N_14167,N_14903);
or U17584 (N_17584,N_15145,N_15479);
and U17585 (N_17585,N_12949,N_15227);
or U17586 (N_17586,N_14535,N_14293);
or U17587 (N_17587,N_12955,N_15100);
nand U17588 (N_17588,N_15231,N_13292);
nor U17589 (N_17589,N_13388,N_14838);
nand U17590 (N_17590,N_12632,N_13811);
or U17591 (N_17591,N_14383,N_14103);
nand U17592 (N_17592,N_14677,N_15117);
nand U17593 (N_17593,N_12622,N_14464);
or U17594 (N_17594,N_15224,N_13771);
or U17595 (N_17595,N_15597,N_14006);
nand U17596 (N_17596,N_13049,N_14246);
or U17597 (N_17597,N_14066,N_14455);
nor U17598 (N_17598,N_15253,N_15033);
or U17599 (N_17599,N_14843,N_13796);
or U17600 (N_17600,N_12616,N_13973);
nand U17601 (N_17601,N_14440,N_14069);
nor U17602 (N_17602,N_12646,N_13047);
xor U17603 (N_17603,N_12787,N_12855);
or U17604 (N_17604,N_15144,N_14546);
or U17605 (N_17605,N_12626,N_14359);
nand U17606 (N_17606,N_14030,N_14011);
or U17607 (N_17607,N_13318,N_12666);
and U17608 (N_17608,N_13119,N_13316);
or U17609 (N_17609,N_14737,N_13148);
nor U17610 (N_17610,N_15157,N_13039);
xor U17611 (N_17611,N_14521,N_14830);
nand U17612 (N_17612,N_12570,N_12989);
nor U17613 (N_17613,N_15205,N_12805);
xnor U17614 (N_17614,N_15576,N_14491);
nand U17615 (N_17615,N_14184,N_13390);
nor U17616 (N_17616,N_13160,N_14774);
nand U17617 (N_17617,N_12532,N_14338);
or U17618 (N_17618,N_14659,N_12720);
and U17619 (N_17619,N_13019,N_15020);
and U17620 (N_17620,N_13208,N_15488);
nor U17621 (N_17621,N_15357,N_13659);
or U17622 (N_17622,N_14238,N_13772);
nor U17623 (N_17623,N_14256,N_13358);
nor U17624 (N_17624,N_15560,N_14376);
nand U17625 (N_17625,N_14519,N_13192);
nand U17626 (N_17626,N_14350,N_13507);
xnor U17627 (N_17627,N_14754,N_13012);
nand U17628 (N_17628,N_14591,N_12522);
and U17629 (N_17629,N_15354,N_13965);
and U17630 (N_17630,N_13705,N_14195);
nor U17631 (N_17631,N_12988,N_13719);
xor U17632 (N_17632,N_13441,N_13213);
or U17633 (N_17633,N_13404,N_15249);
nor U17634 (N_17634,N_13361,N_14032);
or U17635 (N_17635,N_12562,N_13879);
nor U17636 (N_17636,N_14171,N_13387);
xnor U17637 (N_17637,N_15210,N_15059);
nor U17638 (N_17638,N_13002,N_14723);
and U17639 (N_17639,N_14109,N_14982);
or U17640 (N_17640,N_15513,N_14515);
or U17641 (N_17641,N_15183,N_14209);
and U17642 (N_17642,N_13062,N_13730);
nand U17643 (N_17643,N_12530,N_15407);
and U17644 (N_17644,N_13113,N_14648);
and U17645 (N_17645,N_13344,N_13121);
nor U17646 (N_17646,N_15143,N_13976);
and U17647 (N_17647,N_13353,N_14509);
or U17648 (N_17648,N_14746,N_15242);
or U17649 (N_17649,N_13493,N_14805);
and U17650 (N_17650,N_13880,N_14264);
and U17651 (N_17651,N_13644,N_13996);
and U17652 (N_17652,N_13515,N_12769);
nor U17653 (N_17653,N_15219,N_13882);
or U17654 (N_17654,N_13672,N_15289);
nor U17655 (N_17655,N_13736,N_14977);
nor U17656 (N_17656,N_14733,N_13378);
nand U17657 (N_17657,N_15393,N_12982);
xnor U17658 (N_17658,N_14517,N_13320);
or U17659 (N_17659,N_14078,N_12938);
and U17660 (N_17660,N_13770,N_13785);
and U17661 (N_17661,N_13729,N_14666);
and U17662 (N_17662,N_15105,N_14455);
or U17663 (N_17663,N_13797,N_13337);
nand U17664 (N_17664,N_13197,N_14384);
xnor U17665 (N_17665,N_13895,N_12909);
xor U17666 (N_17666,N_13316,N_12599);
or U17667 (N_17667,N_13577,N_13573);
nor U17668 (N_17668,N_14475,N_12914);
nand U17669 (N_17669,N_14775,N_14308);
nor U17670 (N_17670,N_15322,N_13349);
xor U17671 (N_17671,N_12911,N_13301);
xnor U17672 (N_17672,N_12614,N_15413);
nor U17673 (N_17673,N_13840,N_14444);
xor U17674 (N_17674,N_15224,N_14653);
nand U17675 (N_17675,N_13423,N_15165);
nor U17676 (N_17676,N_15110,N_13284);
nand U17677 (N_17677,N_14558,N_12562);
nand U17678 (N_17678,N_14409,N_15035);
nor U17679 (N_17679,N_13822,N_15061);
and U17680 (N_17680,N_15063,N_13305);
nand U17681 (N_17681,N_14281,N_12884);
and U17682 (N_17682,N_15168,N_13098);
and U17683 (N_17683,N_13043,N_15494);
nand U17684 (N_17684,N_14134,N_13967);
nor U17685 (N_17685,N_14485,N_12885);
nor U17686 (N_17686,N_13816,N_15186);
xor U17687 (N_17687,N_13329,N_15085);
and U17688 (N_17688,N_12759,N_15145);
and U17689 (N_17689,N_14350,N_13865);
and U17690 (N_17690,N_12792,N_13980);
nor U17691 (N_17691,N_13903,N_13859);
nor U17692 (N_17692,N_13835,N_12969);
nand U17693 (N_17693,N_14145,N_14941);
xnor U17694 (N_17694,N_13000,N_13594);
nand U17695 (N_17695,N_12532,N_12638);
and U17696 (N_17696,N_15329,N_13747);
nand U17697 (N_17697,N_15143,N_13974);
nor U17698 (N_17698,N_15115,N_14024);
or U17699 (N_17699,N_13307,N_14625);
nand U17700 (N_17700,N_12942,N_13912);
nor U17701 (N_17701,N_12789,N_14320);
or U17702 (N_17702,N_13088,N_12969);
nor U17703 (N_17703,N_12912,N_14955);
nor U17704 (N_17704,N_15164,N_12501);
nand U17705 (N_17705,N_12856,N_14895);
xnor U17706 (N_17706,N_13917,N_14381);
nand U17707 (N_17707,N_14902,N_13981);
and U17708 (N_17708,N_13681,N_15230);
or U17709 (N_17709,N_12513,N_14398);
nor U17710 (N_17710,N_13457,N_15416);
nand U17711 (N_17711,N_14115,N_15529);
nand U17712 (N_17712,N_14739,N_14417);
nor U17713 (N_17713,N_14854,N_12503);
nor U17714 (N_17714,N_14685,N_13979);
or U17715 (N_17715,N_14472,N_13499);
nand U17716 (N_17716,N_15209,N_14177);
nand U17717 (N_17717,N_12639,N_15322);
xor U17718 (N_17718,N_13544,N_13868);
nand U17719 (N_17719,N_14047,N_12780);
or U17720 (N_17720,N_14148,N_15574);
or U17721 (N_17721,N_12911,N_14759);
and U17722 (N_17722,N_13193,N_15261);
and U17723 (N_17723,N_13172,N_13011);
xnor U17724 (N_17724,N_14570,N_14776);
nand U17725 (N_17725,N_15077,N_14636);
nand U17726 (N_17726,N_15224,N_13329);
or U17727 (N_17727,N_13782,N_14552);
nor U17728 (N_17728,N_13875,N_15009);
and U17729 (N_17729,N_12535,N_13525);
and U17730 (N_17730,N_14171,N_15543);
nor U17731 (N_17731,N_12959,N_13936);
or U17732 (N_17732,N_12731,N_15297);
nand U17733 (N_17733,N_13352,N_14034);
nor U17734 (N_17734,N_12622,N_14301);
nand U17735 (N_17735,N_13979,N_14605);
and U17736 (N_17736,N_13549,N_14079);
nor U17737 (N_17737,N_15520,N_13601);
or U17738 (N_17738,N_15528,N_14666);
or U17739 (N_17739,N_13580,N_13255);
and U17740 (N_17740,N_13529,N_14627);
nor U17741 (N_17741,N_14259,N_13350);
nor U17742 (N_17742,N_14994,N_15150);
or U17743 (N_17743,N_13931,N_15331);
or U17744 (N_17744,N_14004,N_13183);
or U17745 (N_17745,N_14527,N_14977);
nand U17746 (N_17746,N_14328,N_14324);
nand U17747 (N_17747,N_13294,N_14469);
and U17748 (N_17748,N_15270,N_15423);
nand U17749 (N_17749,N_15253,N_13048);
or U17750 (N_17750,N_14773,N_13042);
and U17751 (N_17751,N_13159,N_13150);
or U17752 (N_17752,N_13150,N_13701);
nor U17753 (N_17753,N_13233,N_13253);
and U17754 (N_17754,N_14908,N_13951);
nand U17755 (N_17755,N_14485,N_14935);
nand U17756 (N_17756,N_12571,N_13516);
nand U17757 (N_17757,N_12717,N_14362);
nand U17758 (N_17758,N_12855,N_13516);
xor U17759 (N_17759,N_14523,N_13747);
nand U17760 (N_17760,N_14671,N_15131);
nand U17761 (N_17761,N_15486,N_12546);
nand U17762 (N_17762,N_12657,N_13012);
or U17763 (N_17763,N_13127,N_14692);
or U17764 (N_17764,N_12538,N_12716);
nor U17765 (N_17765,N_15421,N_13041);
or U17766 (N_17766,N_14676,N_13677);
and U17767 (N_17767,N_15440,N_12894);
xnor U17768 (N_17768,N_13925,N_14478);
and U17769 (N_17769,N_14937,N_13055);
or U17770 (N_17770,N_15158,N_12997);
nor U17771 (N_17771,N_15437,N_13355);
or U17772 (N_17772,N_13151,N_14669);
nor U17773 (N_17773,N_14638,N_12633);
or U17774 (N_17774,N_15496,N_15094);
nand U17775 (N_17775,N_15081,N_12940);
nor U17776 (N_17776,N_12811,N_12947);
or U17777 (N_17777,N_14198,N_12910);
nor U17778 (N_17778,N_14984,N_14217);
nor U17779 (N_17779,N_13093,N_14740);
or U17780 (N_17780,N_13069,N_13065);
and U17781 (N_17781,N_13858,N_13649);
nand U17782 (N_17782,N_15146,N_13666);
and U17783 (N_17783,N_13589,N_13052);
and U17784 (N_17784,N_13058,N_13083);
and U17785 (N_17785,N_14596,N_14624);
xnor U17786 (N_17786,N_13273,N_14236);
nor U17787 (N_17787,N_12731,N_15470);
nand U17788 (N_17788,N_13165,N_14060);
or U17789 (N_17789,N_13437,N_13378);
nor U17790 (N_17790,N_12980,N_13874);
or U17791 (N_17791,N_14235,N_13031);
nand U17792 (N_17792,N_14134,N_13906);
nand U17793 (N_17793,N_15610,N_13132);
xnor U17794 (N_17794,N_13779,N_14250);
or U17795 (N_17795,N_13885,N_13218);
nand U17796 (N_17796,N_13919,N_13116);
nand U17797 (N_17797,N_15009,N_13594);
nor U17798 (N_17798,N_14011,N_14047);
nor U17799 (N_17799,N_15529,N_14400);
and U17800 (N_17800,N_14345,N_12816);
or U17801 (N_17801,N_14593,N_14180);
or U17802 (N_17802,N_14092,N_13483);
or U17803 (N_17803,N_12613,N_14524);
or U17804 (N_17804,N_13848,N_15372);
xnor U17805 (N_17805,N_14442,N_13880);
nand U17806 (N_17806,N_14130,N_15412);
nand U17807 (N_17807,N_12853,N_14782);
nand U17808 (N_17808,N_12586,N_13069);
nor U17809 (N_17809,N_12661,N_14561);
or U17810 (N_17810,N_14752,N_13579);
and U17811 (N_17811,N_13028,N_14387);
nand U17812 (N_17812,N_15072,N_13471);
xor U17813 (N_17813,N_15219,N_12516);
or U17814 (N_17814,N_15336,N_13154);
nand U17815 (N_17815,N_15309,N_14309);
or U17816 (N_17816,N_12910,N_14954);
nand U17817 (N_17817,N_13085,N_14638);
or U17818 (N_17818,N_15479,N_13405);
or U17819 (N_17819,N_12652,N_15581);
and U17820 (N_17820,N_14199,N_13082);
or U17821 (N_17821,N_13883,N_14252);
or U17822 (N_17822,N_13619,N_14966);
or U17823 (N_17823,N_15463,N_13040);
xor U17824 (N_17824,N_15141,N_13166);
or U17825 (N_17825,N_15365,N_15303);
nand U17826 (N_17826,N_14234,N_14866);
nor U17827 (N_17827,N_13699,N_13481);
and U17828 (N_17828,N_12810,N_14058);
xor U17829 (N_17829,N_12503,N_12548);
nand U17830 (N_17830,N_14301,N_13476);
or U17831 (N_17831,N_13652,N_12615);
nor U17832 (N_17832,N_14632,N_12732);
nor U17833 (N_17833,N_12531,N_14377);
xnor U17834 (N_17834,N_13881,N_12753);
nor U17835 (N_17835,N_15468,N_15564);
or U17836 (N_17836,N_14368,N_13467);
nand U17837 (N_17837,N_13909,N_14609);
or U17838 (N_17838,N_14184,N_13742);
and U17839 (N_17839,N_15204,N_14704);
nand U17840 (N_17840,N_13404,N_14877);
and U17841 (N_17841,N_15577,N_13424);
or U17842 (N_17842,N_12596,N_12812);
and U17843 (N_17843,N_13418,N_13944);
or U17844 (N_17844,N_14380,N_15183);
nor U17845 (N_17845,N_14250,N_13194);
or U17846 (N_17846,N_14334,N_15442);
xor U17847 (N_17847,N_14215,N_12585);
and U17848 (N_17848,N_14429,N_12638);
nor U17849 (N_17849,N_13059,N_12642);
xnor U17850 (N_17850,N_13051,N_13317);
nor U17851 (N_17851,N_14015,N_14660);
or U17852 (N_17852,N_14288,N_14715);
or U17853 (N_17853,N_15408,N_14046);
nor U17854 (N_17854,N_13780,N_14229);
xnor U17855 (N_17855,N_14700,N_13402);
nand U17856 (N_17856,N_14145,N_15089);
or U17857 (N_17857,N_14965,N_13822);
nor U17858 (N_17858,N_14965,N_15353);
or U17859 (N_17859,N_14071,N_15117);
or U17860 (N_17860,N_13592,N_14665);
or U17861 (N_17861,N_13973,N_14161);
or U17862 (N_17862,N_13258,N_14738);
or U17863 (N_17863,N_14452,N_15554);
nor U17864 (N_17864,N_14794,N_14977);
nor U17865 (N_17865,N_13817,N_13216);
and U17866 (N_17866,N_14654,N_14365);
and U17867 (N_17867,N_14002,N_14372);
xor U17868 (N_17868,N_13393,N_13637);
and U17869 (N_17869,N_14715,N_15266);
or U17870 (N_17870,N_14694,N_13176);
nor U17871 (N_17871,N_13173,N_13214);
xnor U17872 (N_17872,N_14470,N_12577);
nand U17873 (N_17873,N_14417,N_15265);
or U17874 (N_17874,N_13330,N_12735);
xnor U17875 (N_17875,N_12894,N_15582);
nor U17876 (N_17876,N_12742,N_14042);
nand U17877 (N_17877,N_12848,N_13620);
nand U17878 (N_17878,N_14738,N_14673);
nor U17879 (N_17879,N_15115,N_12864);
nor U17880 (N_17880,N_14529,N_12567);
nand U17881 (N_17881,N_15036,N_15088);
and U17882 (N_17882,N_14934,N_15096);
and U17883 (N_17883,N_14596,N_14891);
xnor U17884 (N_17884,N_12722,N_14400);
and U17885 (N_17885,N_14493,N_13094);
xnor U17886 (N_17886,N_13473,N_13813);
or U17887 (N_17887,N_13223,N_14421);
and U17888 (N_17888,N_14681,N_13340);
nor U17889 (N_17889,N_13427,N_14716);
or U17890 (N_17890,N_14427,N_12737);
nor U17891 (N_17891,N_14527,N_14933);
and U17892 (N_17892,N_14903,N_14914);
and U17893 (N_17893,N_14170,N_14240);
nand U17894 (N_17894,N_13790,N_14820);
nand U17895 (N_17895,N_12900,N_15566);
or U17896 (N_17896,N_13517,N_13787);
or U17897 (N_17897,N_13669,N_12590);
xnor U17898 (N_17898,N_14507,N_13083);
nor U17899 (N_17899,N_15311,N_13913);
nor U17900 (N_17900,N_13225,N_14323);
nor U17901 (N_17901,N_13134,N_13809);
nand U17902 (N_17902,N_14410,N_14989);
nor U17903 (N_17903,N_13071,N_13139);
nand U17904 (N_17904,N_12947,N_15528);
or U17905 (N_17905,N_14960,N_13390);
nand U17906 (N_17906,N_12941,N_15299);
or U17907 (N_17907,N_13537,N_13904);
nor U17908 (N_17908,N_12728,N_12787);
nand U17909 (N_17909,N_13627,N_13009);
or U17910 (N_17910,N_12760,N_13861);
nand U17911 (N_17911,N_13528,N_14222);
nand U17912 (N_17912,N_12987,N_15303);
nand U17913 (N_17913,N_14320,N_14899);
or U17914 (N_17914,N_12618,N_13796);
and U17915 (N_17915,N_14077,N_14975);
nand U17916 (N_17916,N_15395,N_12603);
nand U17917 (N_17917,N_14333,N_14276);
or U17918 (N_17918,N_13006,N_14551);
and U17919 (N_17919,N_12830,N_12550);
and U17920 (N_17920,N_13561,N_12688);
and U17921 (N_17921,N_12617,N_13380);
and U17922 (N_17922,N_15256,N_15365);
nand U17923 (N_17923,N_14284,N_12743);
or U17924 (N_17924,N_14223,N_13326);
and U17925 (N_17925,N_15462,N_12784);
or U17926 (N_17926,N_12898,N_13263);
nand U17927 (N_17927,N_12948,N_14377);
nor U17928 (N_17928,N_14216,N_12777);
nor U17929 (N_17929,N_13414,N_15047);
or U17930 (N_17930,N_12770,N_13699);
and U17931 (N_17931,N_13208,N_12869);
and U17932 (N_17932,N_13982,N_12869);
or U17933 (N_17933,N_13279,N_14375);
nor U17934 (N_17934,N_13686,N_13226);
and U17935 (N_17935,N_15595,N_15523);
nor U17936 (N_17936,N_13841,N_15220);
nor U17937 (N_17937,N_13516,N_14083);
or U17938 (N_17938,N_14305,N_15559);
nand U17939 (N_17939,N_13526,N_13546);
and U17940 (N_17940,N_15447,N_14593);
or U17941 (N_17941,N_14171,N_14008);
or U17942 (N_17942,N_13222,N_12896);
or U17943 (N_17943,N_12696,N_13093);
or U17944 (N_17944,N_13955,N_12960);
nand U17945 (N_17945,N_14971,N_15424);
nor U17946 (N_17946,N_14571,N_13828);
or U17947 (N_17947,N_15277,N_14121);
nor U17948 (N_17948,N_12813,N_14627);
or U17949 (N_17949,N_12986,N_13113);
nand U17950 (N_17950,N_15251,N_14017);
and U17951 (N_17951,N_15135,N_13549);
and U17952 (N_17952,N_12859,N_15576);
nand U17953 (N_17953,N_14552,N_15205);
and U17954 (N_17954,N_15525,N_14320);
nand U17955 (N_17955,N_14985,N_13293);
or U17956 (N_17956,N_13107,N_15143);
nand U17957 (N_17957,N_14456,N_14330);
and U17958 (N_17958,N_13170,N_13355);
nor U17959 (N_17959,N_14641,N_13085);
nor U17960 (N_17960,N_14342,N_15410);
nand U17961 (N_17961,N_14076,N_14865);
nand U17962 (N_17962,N_14138,N_14010);
or U17963 (N_17963,N_15108,N_12798);
xor U17964 (N_17964,N_15514,N_12795);
and U17965 (N_17965,N_13816,N_14163);
nor U17966 (N_17966,N_14904,N_15128);
or U17967 (N_17967,N_15100,N_15159);
and U17968 (N_17968,N_13496,N_12671);
nor U17969 (N_17969,N_12960,N_13858);
nand U17970 (N_17970,N_14755,N_14150);
or U17971 (N_17971,N_14833,N_12528);
and U17972 (N_17972,N_14111,N_15486);
or U17973 (N_17973,N_13920,N_13434);
and U17974 (N_17974,N_15435,N_15521);
nor U17975 (N_17975,N_14940,N_12765);
nor U17976 (N_17976,N_14038,N_12848);
or U17977 (N_17977,N_13907,N_14638);
nor U17978 (N_17978,N_13283,N_14669);
nor U17979 (N_17979,N_14212,N_14960);
and U17980 (N_17980,N_13646,N_15428);
or U17981 (N_17981,N_14645,N_14072);
xor U17982 (N_17982,N_13679,N_15188);
nor U17983 (N_17983,N_15442,N_12995);
nand U17984 (N_17984,N_14404,N_13320);
nor U17985 (N_17985,N_13309,N_14546);
and U17986 (N_17986,N_12679,N_12747);
nand U17987 (N_17987,N_14397,N_15318);
xnor U17988 (N_17988,N_14740,N_14857);
nand U17989 (N_17989,N_15422,N_13061);
and U17990 (N_17990,N_13573,N_15519);
nor U17991 (N_17991,N_15084,N_15381);
nand U17992 (N_17992,N_15474,N_13951);
and U17993 (N_17993,N_14878,N_13173);
nand U17994 (N_17994,N_13111,N_14204);
or U17995 (N_17995,N_15500,N_13519);
and U17996 (N_17996,N_14385,N_13649);
nor U17997 (N_17997,N_12833,N_12538);
nor U17998 (N_17998,N_12612,N_12684);
xor U17999 (N_17999,N_13168,N_12827);
nand U18000 (N_18000,N_13602,N_12883);
or U18001 (N_18001,N_12637,N_13463);
xor U18002 (N_18002,N_15222,N_15086);
nand U18003 (N_18003,N_13602,N_13035);
and U18004 (N_18004,N_15239,N_15380);
or U18005 (N_18005,N_13895,N_14191);
nand U18006 (N_18006,N_13190,N_12887);
or U18007 (N_18007,N_13085,N_14036);
nand U18008 (N_18008,N_14562,N_14489);
and U18009 (N_18009,N_13249,N_14272);
or U18010 (N_18010,N_13780,N_14500);
or U18011 (N_18011,N_14003,N_14788);
and U18012 (N_18012,N_13225,N_15444);
nand U18013 (N_18013,N_15209,N_14099);
or U18014 (N_18014,N_13630,N_13082);
and U18015 (N_18015,N_13557,N_15010);
nor U18016 (N_18016,N_12733,N_14229);
or U18017 (N_18017,N_14280,N_15061);
or U18018 (N_18018,N_14705,N_13317);
or U18019 (N_18019,N_12714,N_12722);
nor U18020 (N_18020,N_14746,N_14162);
and U18021 (N_18021,N_13122,N_15347);
and U18022 (N_18022,N_14153,N_15287);
nor U18023 (N_18023,N_14308,N_12513);
nor U18024 (N_18024,N_12892,N_15308);
and U18025 (N_18025,N_14201,N_15282);
xnor U18026 (N_18026,N_12689,N_13490);
nor U18027 (N_18027,N_15308,N_15186);
nor U18028 (N_18028,N_14906,N_13826);
or U18029 (N_18029,N_14690,N_13515);
nor U18030 (N_18030,N_15553,N_14325);
xor U18031 (N_18031,N_12595,N_14047);
nand U18032 (N_18032,N_12521,N_14855);
nand U18033 (N_18033,N_14559,N_15357);
xor U18034 (N_18034,N_15279,N_13586);
nand U18035 (N_18035,N_13215,N_13528);
and U18036 (N_18036,N_15067,N_14235);
nor U18037 (N_18037,N_13766,N_15234);
and U18038 (N_18038,N_14693,N_13183);
and U18039 (N_18039,N_13947,N_14129);
or U18040 (N_18040,N_14439,N_13634);
and U18041 (N_18041,N_12929,N_14267);
and U18042 (N_18042,N_12523,N_14248);
and U18043 (N_18043,N_14575,N_12999);
xor U18044 (N_18044,N_13840,N_13205);
xor U18045 (N_18045,N_14318,N_14357);
nor U18046 (N_18046,N_15142,N_14065);
nor U18047 (N_18047,N_12576,N_13850);
and U18048 (N_18048,N_14239,N_15605);
or U18049 (N_18049,N_13579,N_15603);
nand U18050 (N_18050,N_15137,N_12817);
nand U18051 (N_18051,N_12995,N_14461);
nand U18052 (N_18052,N_14009,N_14220);
or U18053 (N_18053,N_14489,N_13573);
nand U18054 (N_18054,N_13771,N_13395);
or U18055 (N_18055,N_15320,N_14533);
or U18056 (N_18056,N_13274,N_15469);
or U18057 (N_18057,N_12940,N_15188);
and U18058 (N_18058,N_13485,N_15138);
nor U18059 (N_18059,N_13298,N_14581);
xnor U18060 (N_18060,N_15534,N_13181);
nand U18061 (N_18061,N_15201,N_14244);
xor U18062 (N_18062,N_15343,N_13228);
nand U18063 (N_18063,N_13257,N_13964);
xor U18064 (N_18064,N_14951,N_13837);
nor U18065 (N_18065,N_15137,N_12667);
nor U18066 (N_18066,N_12523,N_15103);
nand U18067 (N_18067,N_14334,N_13989);
and U18068 (N_18068,N_12824,N_15483);
xor U18069 (N_18069,N_15323,N_14147);
nor U18070 (N_18070,N_13531,N_15177);
nor U18071 (N_18071,N_13178,N_14720);
nand U18072 (N_18072,N_13797,N_14762);
nor U18073 (N_18073,N_15177,N_12861);
and U18074 (N_18074,N_15191,N_14456);
and U18075 (N_18075,N_14030,N_13166);
or U18076 (N_18076,N_14191,N_13134);
and U18077 (N_18077,N_13906,N_14657);
or U18078 (N_18078,N_13651,N_13509);
xor U18079 (N_18079,N_14396,N_14458);
nand U18080 (N_18080,N_12656,N_13696);
or U18081 (N_18081,N_14547,N_14773);
nand U18082 (N_18082,N_13575,N_13562);
and U18083 (N_18083,N_14479,N_15536);
nand U18084 (N_18084,N_13481,N_13515);
xor U18085 (N_18085,N_13488,N_12564);
nor U18086 (N_18086,N_14628,N_14095);
and U18087 (N_18087,N_14552,N_14375);
or U18088 (N_18088,N_12710,N_14238);
or U18089 (N_18089,N_13213,N_12574);
nor U18090 (N_18090,N_12522,N_14432);
or U18091 (N_18091,N_13960,N_14792);
xor U18092 (N_18092,N_15131,N_13165);
xnor U18093 (N_18093,N_13269,N_14878);
nand U18094 (N_18094,N_14447,N_12718);
nand U18095 (N_18095,N_15557,N_13247);
nand U18096 (N_18096,N_12693,N_14983);
xor U18097 (N_18097,N_13742,N_13344);
and U18098 (N_18098,N_13277,N_15494);
xnor U18099 (N_18099,N_12954,N_14056);
xnor U18100 (N_18100,N_13410,N_12847);
nand U18101 (N_18101,N_13776,N_14700);
xor U18102 (N_18102,N_13189,N_12983);
or U18103 (N_18103,N_13084,N_12618);
or U18104 (N_18104,N_13448,N_13334);
and U18105 (N_18105,N_15235,N_12727);
nand U18106 (N_18106,N_14522,N_14108);
nand U18107 (N_18107,N_14669,N_13223);
and U18108 (N_18108,N_15289,N_13143);
nand U18109 (N_18109,N_14359,N_14826);
xor U18110 (N_18110,N_13533,N_13526);
and U18111 (N_18111,N_13049,N_14291);
nand U18112 (N_18112,N_12860,N_12592);
and U18113 (N_18113,N_15371,N_15370);
nor U18114 (N_18114,N_14180,N_15456);
xor U18115 (N_18115,N_15452,N_13677);
or U18116 (N_18116,N_14038,N_13003);
or U18117 (N_18117,N_14178,N_14482);
xor U18118 (N_18118,N_13157,N_12801);
or U18119 (N_18119,N_13065,N_13058);
nand U18120 (N_18120,N_14590,N_15555);
or U18121 (N_18121,N_13260,N_14349);
nand U18122 (N_18122,N_14695,N_15151);
or U18123 (N_18123,N_14301,N_12864);
and U18124 (N_18124,N_14928,N_14088);
and U18125 (N_18125,N_14317,N_13481);
nor U18126 (N_18126,N_12821,N_14152);
and U18127 (N_18127,N_14582,N_15358);
nor U18128 (N_18128,N_13503,N_13841);
and U18129 (N_18129,N_13648,N_12945);
nand U18130 (N_18130,N_15199,N_14712);
or U18131 (N_18131,N_14337,N_15103);
and U18132 (N_18132,N_13898,N_13754);
nand U18133 (N_18133,N_13316,N_14737);
nand U18134 (N_18134,N_13561,N_14183);
xnor U18135 (N_18135,N_13630,N_15618);
or U18136 (N_18136,N_13578,N_14996);
and U18137 (N_18137,N_14561,N_13557);
and U18138 (N_18138,N_13765,N_14700);
xnor U18139 (N_18139,N_14213,N_14892);
xor U18140 (N_18140,N_14719,N_14038);
nand U18141 (N_18141,N_15583,N_13596);
nand U18142 (N_18142,N_13911,N_13813);
xnor U18143 (N_18143,N_14007,N_14503);
or U18144 (N_18144,N_13146,N_14706);
or U18145 (N_18145,N_15348,N_14531);
nor U18146 (N_18146,N_13457,N_15135);
nor U18147 (N_18147,N_14190,N_14284);
nor U18148 (N_18148,N_12828,N_13924);
and U18149 (N_18149,N_13871,N_15260);
nand U18150 (N_18150,N_15460,N_14197);
nor U18151 (N_18151,N_13335,N_13255);
and U18152 (N_18152,N_15363,N_13087);
and U18153 (N_18153,N_12670,N_13034);
or U18154 (N_18154,N_13874,N_13859);
or U18155 (N_18155,N_13664,N_14622);
nor U18156 (N_18156,N_14530,N_15516);
nor U18157 (N_18157,N_13439,N_14740);
nand U18158 (N_18158,N_13033,N_14710);
nor U18159 (N_18159,N_13313,N_13250);
nor U18160 (N_18160,N_14785,N_13013);
or U18161 (N_18161,N_15185,N_14756);
xor U18162 (N_18162,N_13934,N_14139);
and U18163 (N_18163,N_13599,N_15593);
nand U18164 (N_18164,N_15465,N_13973);
nor U18165 (N_18165,N_12963,N_13381);
nor U18166 (N_18166,N_12572,N_13404);
nand U18167 (N_18167,N_14591,N_14975);
xnor U18168 (N_18168,N_12688,N_14556);
nor U18169 (N_18169,N_13786,N_15042);
nand U18170 (N_18170,N_13450,N_14418);
nor U18171 (N_18171,N_13732,N_14071);
nor U18172 (N_18172,N_13984,N_15470);
nor U18173 (N_18173,N_13056,N_13546);
nor U18174 (N_18174,N_12888,N_12956);
or U18175 (N_18175,N_13056,N_14128);
nand U18176 (N_18176,N_13238,N_15380);
nand U18177 (N_18177,N_13404,N_15256);
and U18178 (N_18178,N_12588,N_12947);
nor U18179 (N_18179,N_14164,N_15028);
nand U18180 (N_18180,N_13941,N_13820);
or U18181 (N_18181,N_13707,N_15270);
and U18182 (N_18182,N_14421,N_13421);
nand U18183 (N_18183,N_15380,N_15555);
nor U18184 (N_18184,N_14455,N_15350);
nor U18185 (N_18185,N_15186,N_13669);
xnor U18186 (N_18186,N_12555,N_13522);
nor U18187 (N_18187,N_13337,N_15357);
and U18188 (N_18188,N_14529,N_14844);
nand U18189 (N_18189,N_13767,N_13482);
nor U18190 (N_18190,N_12960,N_15597);
nor U18191 (N_18191,N_14299,N_14898);
and U18192 (N_18192,N_14665,N_14993);
nor U18193 (N_18193,N_15027,N_13913);
nor U18194 (N_18194,N_13167,N_14824);
and U18195 (N_18195,N_14671,N_15252);
nor U18196 (N_18196,N_14342,N_13384);
xor U18197 (N_18197,N_14018,N_14706);
or U18198 (N_18198,N_14389,N_13196);
nand U18199 (N_18199,N_15285,N_12922);
nand U18200 (N_18200,N_15199,N_13427);
nor U18201 (N_18201,N_14749,N_12974);
nand U18202 (N_18202,N_12682,N_14643);
and U18203 (N_18203,N_15401,N_12825);
or U18204 (N_18204,N_13071,N_14406);
or U18205 (N_18205,N_14341,N_15174);
nand U18206 (N_18206,N_12911,N_14335);
nor U18207 (N_18207,N_15283,N_15119);
nor U18208 (N_18208,N_13963,N_15372);
or U18209 (N_18209,N_15128,N_13425);
nor U18210 (N_18210,N_13029,N_15186);
or U18211 (N_18211,N_14338,N_12657);
nand U18212 (N_18212,N_12615,N_13903);
and U18213 (N_18213,N_14651,N_13560);
or U18214 (N_18214,N_13729,N_15332);
and U18215 (N_18215,N_14538,N_13060);
nand U18216 (N_18216,N_13975,N_14267);
nand U18217 (N_18217,N_15335,N_15281);
or U18218 (N_18218,N_13876,N_13981);
or U18219 (N_18219,N_12687,N_13301);
or U18220 (N_18220,N_14584,N_13150);
nor U18221 (N_18221,N_15379,N_14407);
nand U18222 (N_18222,N_13065,N_14893);
nand U18223 (N_18223,N_14304,N_15597);
nand U18224 (N_18224,N_13501,N_13221);
xnor U18225 (N_18225,N_14122,N_12689);
and U18226 (N_18226,N_13792,N_13630);
nor U18227 (N_18227,N_13948,N_14350);
and U18228 (N_18228,N_14394,N_14590);
nand U18229 (N_18229,N_12932,N_14032);
nand U18230 (N_18230,N_14526,N_15355);
and U18231 (N_18231,N_14555,N_15495);
xor U18232 (N_18232,N_14345,N_14360);
xnor U18233 (N_18233,N_14090,N_13587);
and U18234 (N_18234,N_14269,N_13967);
xor U18235 (N_18235,N_14339,N_15553);
or U18236 (N_18236,N_15041,N_14057);
nand U18237 (N_18237,N_14100,N_12995);
nand U18238 (N_18238,N_15271,N_13880);
nor U18239 (N_18239,N_12529,N_14896);
or U18240 (N_18240,N_14239,N_14988);
nand U18241 (N_18241,N_14338,N_12868);
nand U18242 (N_18242,N_14265,N_12827);
or U18243 (N_18243,N_14476,N_12646);
and U18244 (N_18244,N_15594,N_14312);
nand U18245 (N_18245,N_13791,N_12818);
and U18246 (N_18246,N_13397,N_13671);
xnor U18247 (N_18247,N_14536,N_14205);
xnor U18248 (N_18248,N_12740,N_14433);
nand U18249 (N_18249,N_14832,N_13139);
or U18250 (N_18250,N_13365,N_14184);
nand U18251 (N_18251,N_12522,N_15597);
nand U18252 (N_18252,N_14583,N_12835);
nand U18253 (N_18253,N_14989,N_13176);
nand U18254 (N_18254,N_13863,N_12561);
and U18255 (N_18255,N_15152,N_14444);
or U18256 (N_18256,N_15591,N_12646);
xnor U18257 (N_18257,N_14032,N_13405);
nor U18258 (N_18258,N_12735,N_15489);
or U18259 (N_18259,N_12776,N_12582);
and U18260 (N_18260,N_14386,N_13132);
nand U18261 (N_18261,N_12847,N_14859);
xor U18262 (N_18262,N_14924,N_15021);
or U18263 (N_18263,N_15456,N_14576);
or U18264 (N_18264,N_13553,N_12895);
and U18265 (N_18265,N_14350,N_14131);
nor U18266 (N_18266,N_13884,N_14586);
or U18267 (N_18267,N_14624,N_13455);
xnor U18268 (N_18268,N_15308,N_13993);
and U18269 (N_18269,N_13445,N_15414);
and U18270 (N_18270,N_15194,N_14370);
or U18271 (N_18271,N_13869,N_14934);
or U18272 (N_18272,N_13781,N_12918);
nor U18273 (N_18273,N_13764,N_13939);
or U18274 (N_18274,N_14911,N_12874);
nor U18275 (N_18275,N_15048,N_14133);
and U18276 (N_18276,N_14674,N_15031);
nor U18277 (N_18277,N_13189,N_12833);
nor U18278 (N_18278,N_14022,N_15288);
nand U18279 (N_18279,N_14684,N_13375);
or U18280 (N_18280,N_14546,N_15335);
nor U18281 (N_18281,N_14198,N_13198);
nor U18282 (N_18282,N_13810,N_14272);
or U18283 (N_18283,N_15054,N_14769);
nand U18284 (N_18284,N_15398,N_12900);
or U18285 (N_18285,N_13297,N_14845);
and U18286 (N_18286,N_15456,N_14409);
nor U18287 (N_18287,N_15305,N_15223);
and U18288 (N_18288,N_13716,N_12691);
and U18289 (N_18289,N_13225,N_14689);
and U18290 (N_18290,N_14435,N_13707);
or U18291 (N_18291,N_13751,N_13458);
nor U18292 (N_18292,N_14134,N_13781);
and U18293 (N_18293,N_13574,N_14623);
or U18294 (N_18294,N_15061,N_13907);
and U18295 (N_18295,N_13516,N_14215);
or U18296 (N_18296,N_15067,N_12838);
nand U18297 (N_18297,N_13031,N_14143);
xnor U18298 (N_18298,N_14610,N_14749);
and U18299 (N_18299,N_12884,N_14450);
nand U18300 (N_18300,N_12904,N_13322);
nor U18301 (N_18301,N_15160,N_13056);
nor U18302 (N_18302,N_15409,N_13770);
or U18303 (N_18303,N_12885,N_12908);
nor U18304 (N_18304,N_12611,N_14887);
and U18305 (N_18305,N_13365,N_14637);
nor U18306 (N_18306,N_14659,N_14789);
and U18307 (N_18307,N_12656,N_13760);
or U18308 (N_18308,N_15237,N_15372);
and U18309 (N_18309,N_12847,N_13158);
nand U18310 (N_18310,N_15387,N_14860);
or U18311 (N_18311,N_13273,N_14861);
and U18312 (N_18312,N_13063,N_15156);
nand U18313 (N_18313,N_13291,N_13175);
nor U18314 (N_18314,N_14712,N_14543);
nand U18315 (N_18315,N_14298,N_14804);
xnor U18316 (N_18316,N_12699,N_13462);
nor U18317 (N_18317,N_13781,N_12742);
or U18318 (N_18318,N_14907,N_14033);
nand U18319 (N_18319,N_12552,N_13944);
xnor U18320 (N_18320,N_14090,N_13124);
and U18321 (N_18321,N_13592,N_14144);
nor U18322 (N_18322,N_13694,N_12696);
nor U18323 (N_18323,N_15341,N_12553);
or U18324 (N_18324,N_15523,N_14272);
or U18325 (N_18325,N_13199,N_14808);
or U18326 (N_18326,N_13972,N_12841);
nand U18327 (N_18327,N_13802,N_14705);
nor U18328 (N_18328,N_13564,N_13344);
and U18329 (N_18329,N_12642,N_12914);
and U18330 (N_18330,N_15571,N_15026);
and U18331 (N_18331,N_15348,N_13036);
nand U18332 (N_18332,N_14007,N_15548);
or U18333 (N_18333,N_15287,N_12961);
and U18334 (N_18334,N_14966,N_12877);
nand U18335 (N_18335,N_15459,N_12708);
nor U18336 (N_18336,N_15210,N_14806);
nor U18337 (N_18337,N_13033,N_13111);
nand U18338 (N_18338,N_13578,N_12712);
or U18339 (N_18339,N_14207,N_13783);
xnor U18340 (N_18340,N_14557,N_12733);
nor U18341 (N_18341,N_14583,N_13980);
nand U18342 (N_18342,N_12633,N_13120);
or U18343 (N_18343,N_12520,N_13822);
nor U18344 (N_18344,N_12631,N_13568);
nand U18345 (N_18345,N_15214,N_12560);
or U18346 (N_18346,N_12610,N_12908);
and U18347 (N_18347,N_12702,N_12887);
and U18348 (N_18348,N_13848,N_13901);
or U18349 (N_18349,N_13898,N_12852);
nand U18350 (N_18350,N_14534,N_15565);
nor U18351 (N_18351,N_15498,N_14287);
nand U18352 (N_18352,N_12952,N_12800);
nand U18353 (N_18353,N_12712,N_13974);
nand U18354 (N_18354,N_12682,N_12888);
or U18355 (N_18355,N_14167,N_15465);
or U18356 (N_18356,N_15548,N_15320);
or U18357 (N_18357,N_14792,N_12592);
nand U18358 (N_18358,N_15485,N_13585);
or U18359 (N_18359,N_14120,N_13815);
nor U18360 (N_18360,N_15125,N_12656);
or U18361 (N_18361,N_14639,N_15213);
nor U18362 (N_18362,N_13860,N_14151);
nor U18363 (N_18363,N_12969,N_14588);
or U18364 (N_18364,N_12783,N_14070);
nor U18365 (N_18365,N_14456,N_13109);
or U18366 (N_18366,N_13355,N_12634);
nor U18367 (N_18367,N_13567,N_13217);
or U18368 (N_18368,N_13861,N_15415);
nor U18369 (N_18369,N_15401,N_13949);
nand U18370 (N_18370,N_14677,N_15047);
xor U18371 (N_18371,N_13869,N_12946);
nor U18372 (N_18372,N_14146,N_12697);
nand U18373 (N_18373,N_14519,N_13179);
xor U18374 (N_18374,N_14631,N_13835);
xor U18375 (N_18375,N_14389,N_12505);
nor U18376 (N_18376,N_12605,N_14872);
nand U18377 (N_18377,N_13477,N_13708);
or U18378 (N_18378,N_14052,N_13271);
nand U18379 (N_18379,N_13942,N_14280);
nand U18380 (N_18380,N_13743,N_15168);
and U18381 (N_18381,N_14049,N_13589);
nand U18382 (N_18382,N_13624,N_14485);
xor U18383 (N_18383,N_13549,N_14927);
and U18384 (N_18384,N_12885,N_14430);
nor U18385 (N_18385,N_14580,N_15145);
or U18386 (N_18386,N_14527,N_13786);
nand U18387 (N_18387,N_13221,N_15458);
or U18388 (N_18388,N_14773,N_15009);
nor U18389 (N_18389,N_14355,N_13663);
nor U18390 (N_18390,N_13200,N_14766);
and U18391 (N_18391,N_14598,N_13840);
or U18392 (N_18392,N_15079,N_14517);
nor U18393 (N_18393,N_13615,N_14229);
and U18394 (N_18394,N_15369,N_15385);
or U18395 (N_18395,N_14211,N_13511);
or U18396 (N_18396,N_14140,N_13608);
nor U18397 (N_18397,N_12660,N_12501);
nand U18398 (N_18398,N_14756,N_13065);
nand U18399 (N_18399,N_12780,N_14549);
or U18400 (N_18400,N_13849,N_14115);
and U18401 (N_18401,N_12569,N_13171);
nand U18402 (N_18402,N_13357,N_14599);
xnor U18403 (N_18403,N_15592,N_13523);
and U18404 (N_18404,N_13679,N_13269);
nand U18405 (N_18405,N_13083,N_14273);
and U18406 (N_18406,N_14485,N_12532);
and U18407 (N_18407,N_13514,N_15563);
nand U18408 (N_18408,N_12828,N_12859);
xnor U18409 (N_18409,N_12731,N_15346);
nand U18410 (N_18410,N_12710,N_14295);
or U18411 (N_18411,N_12846,N_15002);
or U18412 (N_18412,N_13328,N_14741);
or U18413 (N_18413,N_13081,N_13225);
nand U18414 (N_18414,N_14142,N_13420);
and U18415 (N_18415,N_14207,N_14984);
or U18416 (N_18416,N_14277,N_14243);
or U18417 (N_18417,N_12638,N_15425);
nor U18418 (N_18418,N_14578,N_13664);
nor U18419 (N_18419,N_15526,N_14438);
and U18420 (N_18420,N_14659,N_13021);
nor U18421 (N_18421,N_14884,N_15157);
nor U18422 (N_18422,N_14336,N_13790);
nor U18423 (N_18423,N_14296,N_12954);
and U18424 (N_18424,N_14426,N_14363);
nor U18425 (N_18425,N_12691,N_15020);
nor U18426 (N_18426,N_14725,N_14818);
and U18427 (N_18427,N_13967,N_13539);
or U18428 (N_18428,N_13503,N_14464);
and U18429 (N_18429,N_14391,N_14536);
nor U18430 (N_18430,N_13589,N_14345);
and U18431 (N_18431,N_13390,N_13021);
xnor U18432 (N_18432,N_12771,N_12744);
and U18433 (N_18433,N_14089,N_13130);
nor U18434 (N_18434,N_14326,N_15241);
and U18435 (N_18435,N_14749,N_12726);
nand U18436 (N_18436,N_13024,N_13654);
and U18437 (N_18437,N_14641,N_15164);
nand U18438 (N_18438,N_13544,N_13293);
or U18439 (N_18439,N_12550,N_15382);
nand U18440 (N_18440,N_14489,N_13516);
or U18441 (N_18441,N_13034,N_15114);
nor U18442 (N_18442,N_13095,N_14282);
xor U18443 (N_18443,N_13187,N_13062);
xnor U18444 (N_18444,N_13730,N_14985);
and U18445 (N_18445,N_13674,N_14347);
or U18446 (N_18446,N_14348,N_13517);
xnor U18447 (N_18447,N_15452,N_14151);
and U18448 (N_18448,N_15350,N_12754);
nor U18449 (N_18449,N_13355,N_15384);
nor U18450 (N_18450,N_15117,N_15598);
or U18451 (N_18451,N_14749,N_14220);
xnor U18452 (N_18452,N_12808,N_13430);
or U18453 (N_18453,N_14747,N_15056);
nand U18454 (N_18454,N_15399,N_15191);
nand U18455 (N_18455,N_13542,N_14191);
nand U18456 (N_18456,N_15220,N_14305);
nand U18457 (N_18457,N_13113,N_12533);
nand U18458 (N_18458,N_15391,N_12758);
nand U18459 (N_18459,N_12506,N_13618);
or U18460 (N_18460,N_14134,N_13860);
nand U18461 (N_18461,N_13963,N_13531);
nand U18462 (N_18462,N_12815,N_14041);
and U18463 (N_18463,N_13649,N_14819);
xor U18464 (N_18464,N_12806,N_12537);
nand U18465 (N_18465,N_14953,N_13392);
nor U18466 (N_18466,N_13551,N_12564);
or U18467 (N_18467,N_12965,N_15500);
and U18468 (N_18468,N_15330,N_14499);
and U18469 (N_18469,N_13445,N_13596);
nand U18470 (N_18470,N_15596,N_13115);
nand U18471 (N_18471,N_12699,N_14950);
and U18472 (N_18472,N_15351,N_13827);
nand U18473 (N_18473,N_15380,N_15598);
nor U18474 (N_18474,N_13120,N_14250);
nor U18475 (N_18475,N_14409,N_14364);
xnor U18476 (N_18476,N_13366,N_13602);
or U18477 (N_18477,N_14189,N_13876);
nor U18478 (N_18478,N_13547,N_14049);
or U18479 (N_18479,N_15284,N_13611);
nor U18480 (N_18480,N_13737,N_13430);
and U18481 (N_18481,N_14754,N_15209);
and U18482 (N_18482,N_15248,N_12640);
nand U18483 (N_18483,N_14163,N_15021);
nand U18484 (N_18484,N_14737,N_13245);
nand U18485 (N_18485,N_15199,N_13932);
or U18486 (N_18486,N_13229,N_14520);
nor U18487 (N_18487,N_14275,N_12813);
and U18488 (N_18488,N_14979,N_15460);
or U18489 (N_18489,N_15037,N_14778);
xnor U18490 (N_18490,N_15093,N_15287);
nor U18491 (N_18491,N_13942,N_13223);
nor U18492 (N_18492,N_14896,N_15543);
or U18493 (N_18493,N_12997,N_15427);
or U18494 (N_18494,N_13850,N_14288);
or U18495 (N_18495,N_12742,N_13178);
xor U18496 (N_18496,N_13725,N_14257);
nand U18497 (N_18497,N_12884,N_14158);
nor U18498 (N_18498,N_15516,N_12967);
xnor U18499 (N_18499,N_13709,N_13129);
and U18500 (N_18500,N_15021,N_13243);
nor U18501 (N_18501,N_13452,N_13137);
nand U18502 (N_18502,N_14062,N_12863);
and U18503 (N_18503,N_15277,N_14043);
and U18504 (N_18504,N_15022,N_12514);
and U18505 (N_18505,N_15395,N_15324);
xnor U18506 (N_18506,N_13433,N_13572);
and U18507 (N_18507,N_13349,N_13565);
nand U18508 (N_18508,N_14169,N_15474);
nand U18509 (N_18509,N_14653,N_15045);
nand U18510 (N_18510,N_14080,N_14148);
nor U18511 (N_18511,N_13166,N_14659);
nor U18512 (N_18512,N_15600,N_15375);
or U18513 (N_18513,N_13305,N_14973);
nand U18514 (N_18514,N_13314,N_14999);
nor U18515 (N_18515,N_13756,N_15395);
nor U18516 (N_18516,N_13772,N_12906);
or U18517 (N_18517,N_14398,N_14673);
nand U18518 (N_18518,N_12788,N_14671);
or U18519 (N_18519,N_12698,N_13526);
nand U18520 (N_18520,N_14567,N_12842);
nor U18521 (N_18521,N_13740,N_12858);
nor U18522 (N_18522,N_15107,N_13791);
or U18523 (N_18523,N_13709,N_12663);
or U18524 (N_18524,N_12931,N_14021);
xor U18525 (N_18525,N_13585,N_15294);
nand U18526 (N_18526,N_13705,N_13804);
xor U18527 (N_18527,N_12687,N_13618);
or U18528 (N_18528,N_12685,N_14344);
or U18529 (N_18529,N_15556,N_14221);
nand U18530 (N_18530,N_15620,N_14774);
or U18531 (N_18531,N_15214,N_13058);
nand U18532 (N_18532,N_14491,N_12885);
and U18533 (N_18533,N_13874,N_14206);
xnor U18534 (N_18534,N_14742,N_14630);
xor U18535 (N_18535,N_13029,N_14464);
and U18536 (N_18536,N_13133,N_14869);
nor U18537 (N_18537,N_12714,N_14865);
and U18538 (N_18538,N_13849,N_12863);
nand U18539 (N_18539,N_12567,N_13850);
xnor U18540 (N_18540,N_14701,N_12623);
nand U18541 (N_18541,N_14775,N_13687);
nand U18542 (N_18542,N_14526,N_12899);
nor U18543 (N_18543,N_13338,N_12761);
nor U18544 (N_18544,N_12500,N_15354);
or U18545 (N_18545,N_13999,N_14566);
xor U18546 (N_18546,N_15410,N_15282);
nor U18547 (N_18547,N_15046,N_12851);
and U18548 (N_18548,N_13851,N_14926);
nor U18549 (N_18549,N_15551,N_14566);
nand U18550 (N_18550,N_12596,N_12870);
or U18551 (N_18551,N_14714,N_14962);
xnor U18552 (N_18552,N_14882,N_13262);
or U18553 (N_18553,N_14519,N_15250);
or U18554 (N_18554,N_13562,N_13916);
and U18555 (N_18555,N_12843,N_15160);
and U18556 (N_18556,N_15543,N_14076);
and U18557 (N_18557,N_14852,N_14956);
or U18558 (N_18558,N_14948,N_13872);
and U18559 (N_18559,N_14304,N_15520);
xor U18560 (N_18560,N_14418,N_14107);
and U18561 (N_18561,N_14881,N_14223);
nand U18562 (N_18562,N_13079,N_14949);
and U18563 (N_18563,N_13644,N_13233);
nand U18564 (N_18564,N_14897,N_13538);
or U18565 (N_18565,N_13347,N_12695);
or U18566 (N_18566,N_13946,N_12840);
or U18567 (N_18567,N_12916,N_14922);
and U18568 (N_18568,N_13216,N_14888);
and U18569 (N_18569,N_13755,N_13015);
nand U18570 (N_18570,N_15271,N_14175);
and U18571 (N_18571,N_14874,N_14957);
nor U18572 (N_18572,N_12655,N_13967);
and U18573 (N_18573,N_14675,N_13641);
and U18574 (N_18574,N_15507,N_13434);
nand U18575 (N_18575,N_12858,N_12686);
xor U18576 (N_18576,N_14403,N_14817);
nand U18577 (N_18577,N_14612,N_12835);
and U18578 (N_18578,N_14153,N_13445);
or U18579 (N_18579,N_14431,N_13243);
and U18580 (N_18580,N_14760,N_14131);
nor U18581 (N_18581,N_14282,N_13211);
or U18582 (N_18582,N_14897,N_12721);
nor U18583 (N_18583,N_14922,N_12556);
or U18584 (N_18584,N_14941,N_12550);
and U18585 (N_18585,N_15449,N_13572);
and U18586 (N_18586,N_14806,N_13516);
or U18587 (N_18587,N_12850,N_15498);
nor U18588 (N_18588,N_12689,N_15567);
nor U18589 (N_18589,N_12867,N_12586);
nor U18590 (N_18590,N_15012,N_12570);
nor U18591 (N_18591,N_15407,N_13195);
nand U18592 (N_18592,N_15617,N_14135);
and U18593 (N_18593,N_14298,N_13703);
or U18594 (N_18594,N_13934,N_13047);
nand U18595 (N_18595,N_15412,N_12743);
and U18596 (N_18596,N_12857,N_13006);
nor U18597 (N_18597,N_14939,N_12689);
nand U18598 (N_18598,N_15416,N_14284);
and U18599 (N_18599,N_13556,N_14115);
nor U18600 (N_18600,N_13928,N_15445);
nor U18601 (N_18601,N_14948,N_13581);
and U18602 (N_18602,N_14338,N_14342);
nor U18603 (N_18603,N_12680,N_13020);
and U18604 (N_18604,N_15157,N_14529);
xor U18605 (N_18605,N_15513,N_13245);
or U18606 (N_18606,N_13822,N_14112);
and U18607 (N_18607,N_13512,N_14953);
nand U18608 (N_18608,N_14206,N_14892);
or U18609 (N_18609,N_14271,N_12581);
nand U18610 (N_18610,N_14799,N_13965);
nor U18611 (N_18611,N_14252,N_15071);
xnor U18612 (N_18612,N_15085,N_15424);
xnor U18613 (N_18613,N_13630,N_14243);
or U18614 (N_18614,N_14170,N_13856);
nand U18615 (N_18615,N_14093,N_15333);
nand U18616 (N_18616,N_13559,N_15283);
nor U18617 (N_18617,N_14802,N_15478);
nor U18618 (N_18618,N_14658,N_12741);
xor U18619 (N_18619,N_13980,N_14207);
nor U18620 (N_18620,N_13062,N_14719);
or U18621 (N_18621,N_13942,N_13945);
nor U18622 (N_18622,N_15275,N_15582);
and U18623 (N_18623,N_13381,N_14465);
nor U18624 (N_18624,N_14988,N_15288);
nor U18625 (N_18625,N_14243,N_15022);
nor U18626 (N_18626,N_14607,N_13132);
nor U18627 (N_18627,N_12540,N_14514);
nand U18628 (N_18628,N_14948,N_13997);
xnor U18629 (N_18629,N_15097,N_13103);
nor U18630 (N_18630,N_13355,N_14294);
or U18631 (N_18631,N_13089,N_14695);
and U18632 (N_18632,N_15408,N_14525);
and U18633 (N_18633,N_14945,N_13453);
nor U18634 (N_18634,N_13399,N_13610);
and U18635 (N_18635,N_14737,N_14863);
xnor U18636 (N_18636,N_14364,N_12553);
or U18637 (N_18637,N_12819,N_12733);
or U18638 (N_18638,N_14305,N_14004);
xnor U18639 (N_18639,N_15493,N_13757);
or U18640 (N_18640,N_13615,N_13134);
nand U18641 (N_18641,N_14850,N_13209);
nand U18642 (N_18642,N_13363,N_12803);
or U18643 (N_18643,N_13578,N_14471);
and U18644 (N_18644,N_15435,N_14108);
nor U18645 (N_18645,N_12601,N_13012);
nand U18646 (N_18646,N_13158,N_14058);
or U18647 (N_18647,N_15111,N_12588);
and U18648 (N_18648,N_15478,N_14153);
and U18649 (N_18649,N_15313,N_14463);
or U18650 (N_18650,N_15285,N_15260);
or U18651 (N_18651,N_12758,N_13010);
nor U18652 (N_18652,N_13597,N_12505);
nand U18653 (N_18653,N_15351,N_14410);
or U18654 (N_18654,N_14906,N_12661);
or U18655 (N_18655,N_13046,N_14057);
nand U18656 (N_18656,N_12572,N_13773);
nor U18657 (N_18657,N_13702,N_13979);
or U18658 (N_18658,N_13183,N_13628);
nand U18659 (N_18659,N_14563,N_14415);
and U18660 (N_18660,N_13716,N_12786);
nand U18661 (N_18661,N_14633,N_15424);
nand U18662 (N_18662,N_15503,N_13368);
nand U18663 (N_18663,N_13142,N_12630);
nand U18664 (N_18664,N_14836,N_13441);
or U18665 (N_18665,N_14388,N_13934);
or U18666 (N_18666,N_12771,N_14224);
or U18667 (N_18667,N_14627,N_12974);
and U18668 (N_18668,N_14032,N_13018);
and U18669 (N_18669,N_15502,N_14078);
nor U18670 (N_18670,N_13009,N_14422);
xnor U18671 (N_18671,N_14139,N_14449);
and U18672 (N_18672,N_12819,N_12745);
xor U18673 (N_18673,N_14121,N_15097);
nor U18674 (N_18674,N_14322,N_12700);
nand U18675 (N_18675,N_13619,N_12842);
nand U18676 (N_18676,N_15575,N_13757);
and U18677 (N_18677,N_13950,N_13502);
or U18678 (N_18678,N_14644,N_13781);
and U18679 (N_18679,N_13917,N_15081);
nand U18680 (N_18680,N_15203,N_12878);
and U18681 (N_18681,N_14362,N_14912);
and U18682 (N_18682,N_12797,N_13283);
nor U18683 (N_18683,N_14366,N_13441);
or U18684 (N_18684,N_14795,N_14645);
xnor U18685 (N_18685,N_15409,N_14941);
nand U18686 (N_18686,N_13228,N_14139);
xor U18687 (N_18687,N_14556,N_13443);
nor U18688 (N_18688,N_14763,N_14838);
and U18689 (N_18689,N_15235,N_13727);
or U18690 (N_18690,N_14305,N_14214);
or U18691 (N_18691,N_15419,N_14714);
or U18692 (N_18692,N_12664,N_12884);
and U18693 (N_18693,N_14155,N_14813);
or U18694 (N_18694,N_13638,N_14241);
and U18695 (N_18695,N_13423,N_13333);
or U18696 (N_18696,N_13588,N_14328);
and U18697 (N_18697,N_14220,N_13471);
nor U18698 (N_18698,N_13965,N_13894);
and U18699 (N_18699,N_13797,N_14657);
nor U18700 (N_18700,N_13442,N_13510);
nand U18701 (N_18701,N_13285,N_14499);
and U18702 (N_18702,N_13026,N_12970);
nor U18703 (N_18703,N_13493,N_14718);
nor U18704 (N_18704,N_14209,N_15125);
xor U18705 (N_18705,N_15441,N_12890);
and U18706 (N_18706,N_12689,N_14081);
nor U18707 (N_18707,N_12639,N_14057);
nor U18708 (N_18708,N_14769,N_13623);
and U18709 (N_18709,N_14404,N_14211);
and U18710 (N_18710,N_14848,N_13578);
or U18711 (N_18711,N_15502,N_13047);
or U18712 (N_18712,N_13224,N_13048);
or U18713 (N_18713,N_13927,N_13824);
nor U18714 (N_18714,N_12640,N_15044);
or U18715 (N_18715,N_13881,N_15228);
or U18716 (N_18716,N_15195,N_13034);
nand U18717 (N_18717,N_13626,N_12687);
or U18718 (N_18718,N_14352,N_13916);
nand U18719 (N_18719,N_14240,N_13993);
nand U18720 (N_18720,N_13867,N_13579);
nor U18721 (N_18721,N_13683,N_15536);
or U18722 (N_18722,N_15364,N_13718);
and U18723 (N_18723,N_15471,N_15508);
and U18724 (N_18724,N_15049,N_15505);
nand U18725 (N_18725,N_14538,N_14176);
or U18726 (N_18726,N_13242,N_13108);
and U18727 (N_18727,N_13892,N_13190);
xor U18728 (N_18728,N_14866,N_14789);
and U18729 (N_18729,N_13842,N_13366);
nor U18730 (N_18730,N_14814,N_13240);
or U18731 (N_18731,N_12904,N_14187);
xor U18732 (N_18732,N_14853,N_13508);
nor U18733 (N_18733,N_14328,N_15371);
or U18734 (N_18734,N_15588,N_14925);
nor U18735 (N_18735,N_13411,N_15120);
and U18736 (N_18736,N_12591,N_12753);
nor U18737 (N_18737,N_14305,N_14104);
xor U18738 (N_18738,N_15104,N_13733);
xor U18739 (N_18739,N_14881,N_12615);
or U18740 (N_18740,N_13293,N_13383);
or U18741 (N_18741,N_12684,N_15249);
or U18742 (N_18742,N_14959,N_14134);
xnor U18743 (N_18743,N_14597,N_15545);
or U18744 (N_18744,N_13270,N_13321);
nand U18745 (N_18745,N_14520,N_12816);
nor U18746 (N_18746,N_14687,N_13040);
nand U18747 (N_18747,N_13365,N_15576);
xnor U18748 (N_18748,N_13651,N_12604);
nor U18749 (N_18749,N_13966,N_15304);
nand U18750 (N_18750,N_17329,N_15868);
nor U18751 (N_18751,N_17622,N_18676);
nor U18752 (N_18752,N_17276,N_17331);
or U18753 (N_18753,N_16975,N_17980);
nand U18754 (N_18754,N_17448,N_18056);
and U18755 (N_18755,N_15823,N_17242);
nand U18756 (N_18756,N_17846,N_16244);
and U18757 (N_18757,N_15727,N_18232);
or U18758 (N_18758,N_16196,N_18384);
nand U18759 (N_18759,N_16703,N_18455);
or U18760 (N_18760,N_18543,N_16722);
nand U18761 (N_18761,N_18339,N_18406);
nand U18762 (N_18762,N_15809,N_17761);
and U18763 (N_18763,N_18637,N_16598);
or U18764 (N_18764,N_17476,N_16659);
or U18765 (N_18765,N_15648,N_16570);
nor U18766 (N_18766,N_16629,N_17571);
and U18767 (N_18767,N_16061,N_18510);
or U18768 (N_18768,N_16469,N_18053);
nor U18769 (N_18769,N_18545,N_18358);
xor U18770 (N_18770,N_16769,N_15659);
xor U18771 (N_18771,N_16476,N_15704);
or U18772 (N_18772,N_18297,N_16658);
nand U18773 (N_18773,N_17990,N_18018);
nor U18774 (N_18774,N_16094,N_15942);
or U18775 (N_18775,N_15834,N_16983);
or U18776 (N_18776,N_17012,N_16102);
nand U18777 (N_18777,N_16202,N_18307);
nand U18778 (N_18778,N_16153,N_16470);
nor U18779 (N_18779,N_15751,N_18569);
and U18780 (N_18780,N_18480,N_18489);
and U18781 (N_18781,N_17591,N_15780);
or U18782 (N_18782,N_17213,N_15803);
and U18783 (N_18783,N_17303,N_16155);
or U18784 (N_18784,N_18405,N_16784);
or U18785 (N_18785,N_16279,N_16446);
nand U18786 (N_18786,N_18310,N_16667);
nor U18787 (N_18787,N_16529,N_15762);
or U18788 (N_18788,N_17562,N_16489);
and U18789 (N_18789,N_16661,N_18004);
and U18790 (N_18790,N_17743,N_16370);
xor U18791 (N_18791,N_17139,N_15987);
or U18792 (N_18792,N_16323,N_17458);
nor U18793 (N_18793,N_15685,N_16430);
nor U18794 (N_18794,N_17533,N_16653);
or U18795 (N_18795,N_15796,N_18334);
nor U18796 (N_18796,N_17466,N_18642);
and U18797 (N_18797,N_16393,N_16145);
and U18798 (N_18798,N_16282,N_18498);
nor U18799 (N_18799,N_16542,N_18226);
nand U18800 (N_18800,N_17350,N_16727);
or U18801 (N_18801,N_15705,N_18397);
and U18802 (N_18802,N_17346,N_17515);
nand U18803 (N_18803,N_18620,N_16358);
nand U18804 (N_18804,N_16278,N_16862);
nor U18805 (N_18805,N_15862,N_18281);
xor U18806 (N_18806,N_15958,N_17143);
nand U18807 (N_18807,N_16204,N_17689);
nand U18808 (N_18808,N_15883,N_15943);
and U18809 (N_18809,N_16112,N_16432);
nand U18810 (N_18810,N_18689,N_17048);
and U18811 (N_18811,N_17240,N_16031);
nor U18812 (N_18812,N_16456,N_17472);
nor U18813 (N_18813,N_15725,N_15636);
nand U18814 (N_18814,N_17264,N_18114);
nor U18815 (N_18815,N_18693,N_18598);
or U18816 (N_18816,N_16406,N_16685);
nand U18817 (N_18817,N_17419,N_17899);
nand U18818 (N_18818,N_16097,N_15793);
nor U18819 (N_18819,N_15973,N_18286);
or U18820 (N_18820,N_17391,N_16780);
nand U18821 (N_18821,N_15989,N_16675);
nand U18822 (N_18822,N_16616,N_17860);
nor U18823 (N_18823,N_16807,N_17808);
or U18824 (N_18824,N_18321,N_17341);
or U18825 (N_18825,N_17183,N_15820);
nor U18826 (N_18826,N_15983,N_17018);
nor U18827 (N_18827,N_18547,N_16338);
and U18828 (N_18828,N_17325,N_16638);
nor U18829 (N_18829,N_17982,N_18097);
and U18830 (N_18830,N_18675,N_17769);
nor U18831 (N_18831,N_17559,N_15911);
and U18832 (N_18832,N_16054,N_18533);
or U18833 (N_18833,N_16263,N_16090);
xnor U18834 (N_18834,N_16166,N_17411);
or U18835 (N_18835,N_16836,N_16093);
nor U18836 (N_18836,N_17539,N_17468);
nor U18837 (N_18837,N_16396,N_18695);
nor U18838 (N_18838,N_15927,N_17068);
or U18839 (N_18839,N_15992,N_16036);
and U18840 (N_18840,N_18218,N_16644);
nor U18841 (N_18841,N_18118,N_18263);
nand U18842 (N_18842,N_17861,N_16778);
nand U18843 (N_18843,N_16173,N_16201);
nor U18844 (N_18844,N_17995,N_16003);
or U18845 (N_18845,N_18298,N_17198);
nor U18846 (N_18846,N_17713,N_17505);
nor U18847 (N_18847,N_18707,N_17101);
or U18848 (N_18848,N_15741,N_16705);
and U18849 (N_18849,N_17003,N_18440);
xor U18850 (N_18850,N_15890,N_17858);
nor U18851 (N_18851,N_18579,N_17741);
nor U18852 (N_18852,N_16070,N_17330);
and U18853 (N_18853,N_18368,N_15967);
or U18854 (N_18854,N_18199,N_18668);
nand U18855 (N_18855,N_15692,N_17053);
nor U18856 (N_18856,N_15896,N_16325);
and U18857 (N_18857,N_17035,N_17895);
nand U18858 (N_18858,N_17919,N_16940);
or U18859 (N_18859,N_17480,N_17932);
nor U18860 (N_18860,N_17520,N_17088);
or U18861 (N_18861,N_15631,N_18463);
or U18862 (N_18862,N_17024,N_15900);
nand U18863 (N_18863,N_16458,N_15966);
or U18864 (N_18864,N_16952,N_17940);
nor U18865 (N_18865,N_18402,N_17140);
nand U18866 (N_18866,N_17586,N_18472);
nand U18867 (N_18867,N_15728,N_17377);
and U18868 (N_18868,N_16122,N_16682);
xnor U18869 (N_18869,N_17913,N_16422);
nand U18870 (N_18870,N_17361,N_16042);
and U18871 (N_18871,N_17582,N_16146);
nor U18872 (N_18872,N_17510,N_16010);
xnor U18873 (N_18873,N_15691,N_18430);
xor U18874 (N_18874,N_16979,N_16158);
and U18875 (N_18875,N_17395,N_16231);
or U18876 (N_18876,N_16230,N_17939);
and U18877 (N_18877,N_18619,N_15652);
nand U18878 (N_18878,N_18178,N_17208);
or U18879 (N_18879,N_15975,N_16259);
and U18880 (N_18880,N_16310,N_17518);
or U18881 (N_18881,N_16363,N_17031);
or U18882 (N_18882,N_16591,N_16372);
nand U18883 (N_18883,N_17760,N_18703);
and U18884 (N_18884,N_16110,N_17798);
and U18885 (N_18885,N_16630,N_16072);
or U18886 (N_18886,N_18108,N_17216);
nand U18887 (N_18887,N_15821,N_18058);
or U18888 (N_18888,N_17725,N_16413);
nor U18889 (N_18889,N_16418,N_18006);
or U18890 (N_18890,N_16976,N_16283);
or U18891 (N_18891,N_16861,N_17668);
nand U18892 (N_18892,N_15937,N_18445);
and U18893 (N_18893,N_17594,N_15882);
nor U18894 (N_18894,N_17112,N_17127);
and U18895 (N_18895,N_17202,N_17948);
nand U18896 (N_18896,N_16852,N_16198);
nand U18897 (N_18897,N_17179,N_17815);
or U18898 (N_18898,N_17171,N_17495);
or U18899 (N_18899,N_18153,N_17827);
or U18900 (N_18900,N_17454,N_18170);
nand U18901 (N_18901,N_18205,N_16702);
or U18902 (N_18902,N_15847,N_18179);
and U18903 (N_18903,N_16760,N_18089);
nor U18904 (N_18904,N_15644,N_16157);
and U18905 (N_18905,N_17842,N_18048);
nor U18906 (N_18906,N_16210,N_18664);
nor U18907 (N_18907,N_16232,N_17872);
and U18908 (N_18908,N_18554,N_17188);
nand U18909 (N_18909,N_17768,N_15657);
or U18910 (N_18910,N_17925,N_16127);
xnor U18911 (N_18911,N_18016,N_15976);
and U18912 (N_18912,N_17473,N_15650);
nor U18913 (N_18913,N_18119,N_16447);
xor U18914 (N_18914,N_16104,N_16039);
nor U18915 (N_18915,N_18403,N_16512);
nand U18916 (N_18916,N_18528,N_16123);
nor U18917 (N_18917,N_18129,N_17151);
nor U18918 (N_18918,N_18191,N_15646);
xor U18919 (N_18919,N_17380,N_18509);
xor U18920 (N_18920,N_17663,N_18336);
and U18921 (N_18921,N_15717,N_16203);
or U18922 (N_18922,N_16929,N_16240);
or U18923 (N_18923,N_16657,N_17349);
and U18924 (N_18924,N_17791,N_17444);
or U18925 (N_18925,N_16497,N_16656);
and U18926 (N_18926,N_16872,N_18641);
and U18927 (N_18927,N_17737,N_17991);
and U18928 (N_18928,N_17609,N_17356);
xor U18929 (N_18929,N_18540,N_16592);
or U18930 (N_18930,N_16357,N_18366);
nor U18931 (N_18931,N_17837,N_16193);
and U18932 (N_18932,N_16991,N_18364);
nand U18933 (N_18933,N_18107,N_18067);
or U18934 (N_18934,N_16544,N_15649);
nor U18935 (N_18935,N_16774,N_17578);
or U18936 (N_18936,N_18433,N_18019);
nor U18937 (N_18937,N_17707,N_17916);
nand U18938 (N_18938,N_17993,N_17706);
xor U18939 (N_18939,N_17211,N_17886);
or U18940 (N_18940,N_18376,N_17593);
and U18941 (N_18941,N_17189,N_17884);
nor U18942 (N_18942,N_16618,N_16139);
xor U18943 (N_18943,N_18544,N_16669);
nor U18944 (N_18944,N_18370,N_17796);
and U18945 (N_18945,N_18135,N_18106);
and U18946 (N_18946,N_18456,N_16756);
and U18947 (N_18947,N_16663,N_18233);
nor U18948 (N_18948,N_17783,N_17855);
nand U18949 (N_18949,N_18269,N_16842);
and U18950 (N_18950,N_18140,N_16908);
or U18951 (N_18951,N_16297,N_17440);
nor U18952 (N_18952,N_17822,N_18197);
nand U18953 (N_18953,N_16923,N_16893);
or U18954 (N_18954,N_18407,N_17339);
and U18955 (N_18955,N_18473,N_16188);
and U18956 (N_18956,N_17381,N_18512);
nor U18957 (N_18957,N_18080,N_18266);
nand U18958 (N_18958,N_17271,N_17459);
nor U18959 (N_18959,N_17109,N_16850);
and U18960 (N_18960,N_18568,N_16351);
xor U18961 (N_18961,N_17045,N_15753);
and U18962 (N_18962,N_16251,N_17635);
nand U18963 (N_18963,N_15641,N_17650);
nand U18964 (N_18964,N_16462,N_18736);
nor U18965 (N_18965,N_17320,N_17897);
or U18966 (N_18966,N_18317,N_17723);
and U18967 (N_18967,N_18603,N_16346);
xnor U18968 (N_18968,N_16848,N_16977);
nor U18969 (N_18969,N_16967,N_16748);
nor U18970 (N_18970,N_18229,N_18157);
xnor U18971 (N_18971,N_17138,N_16239);
nand U18972 (N_18972,N_16568,N_16066);
nor U18973 (N_18973,N_17898,N_18494);
and U18974 (N_18974,N_15804,N_16319);
and U18975 (N_18975,N_18529,N_15901);
or U18976 (N_18976,N_17947,N_17166);
nor U18977 (N_18977,N_17445,N_17751);
or U18978 (N_18978,N_18502,N_16264);
or U18979 (N_18979,N_18166,N_18274);
and U18980 (N_18980,N_16563,N_16766);
nor U18981 (N_18981,N_15663,N_17008);
nand U18982 (N_18982,N_18657,N_15988);
and U18983 (N_18983,N_17731,N_16015);
and U18984 (N_18984,N_18162,N_18511);
and U18985 (N_18985,N_18388,N_15895);
and U18986 (N_18986,N_17661,N_15682);
nand U18987 (N_18987,N_16341,N_16701);
xor U18988 (N_18988,N_18694,N_17327);
nand U18989 (N_18989,N_17298,N_17836);
nor U18990 (N_18990,N_17283,N_18416);
and U18991 (N_18991,N_16582,N_18690);
or U18992 (N_18992,N_18238,N_17435);
and U18993 (N_18993,N_18168,N_16628);
nand U18994 (N_18994,N_15971,N_17522);
or U18995 (N_18995,N_15830,N_16691);
or U18996 (N_18996,N_16109,N_18589);
and U18997 (N_18997,N_18417,N_15813);
nor U18998 (N_18998,N_18553,N_15656);
and U18999 (N_18999,N_15739,N_18055);
and U19000 (N_19000,N_16806,N_18742);
or U19001 (N_19001,N_17104,N_17976);
nand U19002 (N_19002,N_17747,N_17811);
xnor U19003 (N_19003,N_16603,N_16599);
or U19004 (N_19004,N_16814,N_17431);
or U19005 (N_19005,N_16830,N_15977);
xor U19006 (N_19006,N_16348,N_16532);
nand U19007 (N_19007,N_18306,N_15959);
nand U19008 (N_19008,N_16419,N_18651);
nor U19009 (N_19009,N_16622,N_18715);
or U19010 (N_19010,N_17201,N_15950);
nand U19011 (N_19011,N_18063,N_16474);
nand U19012 (N_19012,N_15635,N_17504);
nor U19013 (N_19013,N_17296,N_17810);
nand U19014 (N_19014,N_17187,N_16607);
nand U19015 (N_19015,N_15894,N_17375);
or U19016 (N_19016,N_18409,N_16546);
or U19017 (N_19017,N_17513,N_18222);
and U19018 (N_19018,N_18017,N_18148);
and U19019 (N_19019,N_15969,N_16641);
nand U19020 (N_19020,N_15714,N_17499);
nor U19021 (N_19021,N_18046,N_16538);
and U19022 (N_19022,N_16725,N_17629);
and U19023 (N_19023,N_15906,N_17696);
or U19024 (N_19024,N_17519,N_16245);
or U19025 (N_19025,N_16808,N_16414);
nor U19026 (N_19026,N_17058,N_17086);
xor U19027 (N_19027,N_18284,N_17758);
nand U19028 (N_19028,N_17022,N_17358);
nand U19029 (N_19029,N_16524,N_15708);
nand U19030 (N_19030,N_18630,N_18361);
xnor U19031 (N_19031,N_18071,N_16790);
nor U19032 (N_19032,N_16941,N_16400);
nand U19033 (N_19033,N_17011,N_18289);
or U19034 (N_19034,N_17483,N_17098);
and U19035 (N_19035,N_16148,N_18186);
or U19036 (N_19036,N_16194,N_15805);
or U19037 (N_19037,N_16617,N_18239);
or U19038 (N_19038,N_16525,N_15738);
and U19039 (N_19039,N_17215,N_17918);
and U19040 (N_19040,N_17042,N_16343);
nor U19041 (N_19041,N_16534,N_17887);
or U19042 (N_19042,N_15846,N_17590);
nor U19043 (N_19043,N_15788,N_16475);
nor U19044 (N_19044,N_17945,N_16825);
and U19045 (N_19045,N_16886,N_17611);
and U19046 (N_19046,N_17038,N_17905);
nor U19047 (N_19047,N_17234,N_16087);
nand U19048 (N_19048,N_16133,N_17926);
nor U19049 (N_19049,N_18485,N_18078);
nor U19050 (N_19050,N_18315,N_18200);
nand U19051 (N_19051,N_17155,N_17805);
or U19052 (N_19052,N_17718,N_18708);
or U19053 (N_19053,N_17524,N_17389);
nand U19054 (N_19054,N_17543,N_16179);
nand U19055 (N_19055,N_18219,N_16938);
nand U19056 (N_19056,N_17604,N_17268);
nand U19057 (N_19057,N_17238,N_16096);
or U19058 (N_19058,N_15684,N_18597);
and U19059 (N_19059,N_17669,N_15961);
nand U19060 (N_19060,N_15784,N_16815);
nor U19061 (N_19061,N_18648,N_17508);
xor U19062 (N_19062,N_18527,N_16314);
nor U19063 (N_19063,N_15736,N_16337);
or U19064 (N_19064,N_18049,N_16295);
or U19065 (N_19065,N_15863,N_18185);
and U19066 (N_19066,N_16519,N_16738);
nand U19067 (N_19067,N_16350,N_18088);
or U19068 (N_19068,N_17549,N_17800);
xnor U19069 (N_19069,N_16687,N_17653);
or U19070 (N_19070,N_18696,N_16833);
or U19071 (N_19071,N_16009,N_16557);
xor U19072 (N_19072,N_16533,N_18497);
nor U19073 (N_19073,N_18549,N_17809);
and U19074 (N_19074,N_18125,N_18037);
nor U19075 (N_19075,N_16936,N_18189);
and U19076 (N_19076,N_18209,N_18206);
xnor U19077 (N_19077,N_18177,N_15836);
nand U19078 (N_19078,N_17693,N_18685);
nand U19079 (N_19079,N_15754,N_18287);
or U19080 (N_19080,N_15880,N_16987);
and U19081 (N_19081,N_16881,N_15791);
or U19082 (N_19082,N_17966,N_17540);
nor U19083 (N_19083,N_15729,N_18660);
nor U19084 (N_19084,N_15910,N_16785);
nor U19085 (N_19085,N_16027,N_15768);
or U19086 (N_19086,N_18246,N_17462);
or U19087 (N_19087,N_17688,N_17062);
and U19088 (N_19088,N_18060,N_17971);
nand U19089 (N_19089,N_17163,N_18007);
nor U19090 (N_19090,N_18571,N_16716);
nand U19091 (N_19091,N_16854,N_17700);
nor U19092 (N_19092,N_16365,N_16498);
nand U19093 (N_19093,N_17365,N_16421);
nor U19094 (N_19094,N_16601,N_17658);
nand U19095 (N_19095,N_16799,N_18094);
nand U19096 (N_19096,N_16420,N_17367);
nand U19097 (N_19097,N_15914,N_16455);
and U19098 (N_19098,N_18670,N_16266);
nand U19099 (N_19099,N_17778,N_16998);
and U19100 (N_19100,N_15926,N_16083);
nand U19101 (N_19101,N_17154,N_18175);
nor U19102 (N_19102,N_18507,N_16482);
nand U19103 (N_19103,N_16646,N_16920);
and U19104 (N_19104,N_18220,N_17705);
and U19105 (N_19105,N_17430,N_18328);
and U19106 (N_19106,N_16942,N_18699);
nor U19107 (N_19107,N_16209,N_17221);
nor U19108 (N_19108,N_16270,N_16294);
nor U19109 (N_19109,N_18204,N_18044);
and U19110 (N_19110,N_18247,N_17040);
nor U19111 (N_19111,N_16043,N_16997);
and U19112 (N_19112,N_16345,N_16496);
xor U19113 (N_19113,N_16905,N_17259);
or U19114 (N_19114,N_16781,N_18558);
nor U19115 (N_19115,N_17636,N_18225);
nor U19116 (N_19116,N_17099,N_18330);
nor U19117 (N_19117,N_17660,N_17083);
nand U19118 (N_19118,N_17854,N_16890);
nor U19119 (N_19119,N_16246,N_15946);
or U19120 (N_19120,N_16080,N_16129);
or U19121 (N_19121,N_18688,N_16499);
xor U19122 (N_19122,N_17450,N_18322);
nor U19123 (N_19123,N_17826,N_16017);
nand U19124 (N_19124,N_16856,N_17383);
or U19125 (N_19125,N_16473,N_18365);
and U19126 (N_19126,N_18158,N_16824);
or U19127 (N_19127,N_18038,N_18556);
nor U19128 (N_19128,N_17147,N_16897);
or U19129 (N_19129,N_16863,N_17665);
nand U19130 (N_19130,N_18398,N_16437);
nor U19131 (N_19131,N_16569,N_16980);
nand U19132 (N_19132,N_15661,N_16957);
nand U19133 (N_19133,N_17790,N_18681);
or U19134 (N_19134,N_16220,N_16523);
or U19135 (N_19135,N_16804,N_18749);
and U19136 (N_19136,N_17424,N_17674);
nor U19137 (N_19137,N_17799,N_15695);
or U19138 (N_19138,N_16913,N_18745);
and U19139 (N_19139,N_16032,N_15839);
nor U19140 (N_19140,N_18352,N_18419);
nor U19141 (N_19141,N_17030,N_15848);
or U19142 (N_19142,N_16739,N_18679);
and U19143 (N_19143,N_15929,N_16958);
and U19144 (N_19144,N_16047,N_16505);
xnor U19145 (N_19145,N_16626,N_17108);
and U19146 (N_19146,N_16966,N_18112);
nor U19147 (N_19147,N_17004,N_16688);
xnor U19148 (N_19148,N_16164,N_15897);
nor U19149 (N_19149,N_17906,N_15843);
nand U19150 (N_19150,N_18264,N_18737);
or U19151 (N_19151,N_17106,N_17773);
or U19152 (N_19152,N_18032,N_16186);
nor U19153 (N_19153,N_15790,N_17255);
nor U19154 (N_19154,N_18001,N_16312);
nand U19155 (N_19155,N_17293,N_17670);
or U19156 (N_19156,N_18500,N_15683);
or U19157 (N_19157,N_17054,N_16354);
or U19158 (N_19158,N_17061,N_16819);
nor U19159 (N_19159,N_17479,N_16069);
and U19160 (N_19160,N_16789,N_18329);
nor U19161 (N_19161,N_17409,N_18577);
nor U19162 (N_19162,N_16768,N_16999);
nand U19163 (N_19163,N_18565,N_18677);
or U19164 (N_19164,N_16857,N_17020);
or U19165 (N_19165,N_18267,N_18081);
nand U19166 (N_19166,N_16973,N_17623);
or U19167 (N_19167,N_17775,N_17025);
xor U19168 (N_19168,N_18534,N_16671);
nand U19169 (N_19169,N_16255,N_16613);
nand U19170 (N_19170,N_16490,N_16448);
or U19171 (N_19171,N_16029,N_16288);
nand U19172 (N_19172,N_16693,N_16214);
nor U19173 (N_19173,N_16621,N_16404);
or U19174 (N_19174,N_17942,N_15720);
and U19175 (N_19175,N_18325,N_15643);
and U19176 (N_19176,N_18012,N_18131);
or U19177 (N_19177,N_18729,N_17986);
xor U19178 (N_19178,N_16452,N_18709);
nand U19179 (N_19179,N_15642,N_16386);
nor U19180 (N_19180,N_16590,N_16285);
nor U19181 (N_19181,N_18400,N_16649);
nor U19182 (N_19182,N_17920,N_16556);
or U19183 (N_19183,N_16327,N_16060);
nor U19184 (N_19184,N_16144,N_17941);
xor U19185 (N_19185,N_15690,N_17802);
nor U19186 (N_19186,N_17825,N_16019);
xnor U19187 (N_19187,N_18174,N_17481);
and U19188 (N_19188,N_18662,N_17588);
and U19189 (N_19189,N_18518,N_16812);
or U19190 (N_19190,N_17376,N_16011);
or U19191 (N_19191,N_18033,N_16301);
and U19192 (N_19192,N_18541,N_18578);
xnor U19193 (N_19193,N_16329,N_18726);
nor U19194 (N_19194,N_16318,N_15798);
and U19195 (N_19195,N_17455,N_17818);
nand U19196 (N_19196,N_16442,N_17606);
or U19197 (N_19197,N_17252,N_18522);
nand U19198 (N_19198,N_18002,N_15854);
xnor U19199 (N_19199,N_16241,N_17418);
or U19200 (N_19200,N_18035,N_17368);
and U19201 (N_19201,N_18661,N_16652);
xnor U19202 (N_19202,N_17605,N_15746);
or U19203 (N_19203,N_15956,N_16369);
or U19204 (N_19204,N_17348,N_16755);
and U19205 (N_19205,N_17452,N_17962);
nor U19206 (N_19206,N_17353,N_16614);
and U19207 (N_19207,N_16879,N_16627);
xor U19208 (N_19208,N_17795,N_15865);
or U19209 (N_19209,N_17206,N_17512);
xor U19210 (N_19210,N_17486,N_15700);
nor U19211 (N_19211,N_18230,N_17771);
nor U19212 (N_19212,N_17579,N_16021);
or U19213 (N_19213,N_18308,N_17118);
and U19214 (N_19214,N_16639,N_16805);
xnor U19215 (N_19215,N_17672,N_15870);
nor U19216 (N_19216,N_17681,N_15778);
xnor U19217 (N_19217,N_18583,N_15688);
and U19218 (N_19218,N_18610,N_17241);
or U19219 (N_19219,N_18691,N_18652);
xor U19220 (N_19220,N_15954,N_16562);
and U19221 (N_19221,N_17789,N_17235);
or U19222 (N_19222,N_18160,N_18280);
and U19223 (N_19223,N_17845,N_15711);
nor U19224 (N_19224,N_18074,N_16501);
nor U19225 (N_19225,N_18214,N_15756);
xor U19226 (N_19226,N_17757,N_18327);
nor U19227 (N_19227,N_17194,N_16368);
nor U19228 (N_19228,N_18724,N_15669);
nand U19229 (N_19229,N_16878,N_18235);
and U19230 (N_19230,N_18536,N_16567);
or U19231 (N_19231,N_18656,N_17888);
and U19232 (N_19232,N_18077,N_15899);
nor U19233 (N_19233,N_16035,N_16916);
and U19234 (N_19234,N_18605,N_16892);
nor U19235 (N_19235,N_16082,N_18710);
xor U19236 (N_19236,N_15775,N_17484);
xnor U19237 (N_19237,N_17923,N_16091);
nor U19238 (N_19238,N_18045,N_18588);
nor U19239 (N_19239,N_17978,N_18011);
nor U19240 (N_19240,N_18025,N_18495);
and U19241 (N_19241,N_16005,N_18367);
nand U19242 (N_19242,N_18377,N_16394);
nand U19243 (N_19243,N_18095,N_17460);
nand U19244 (N_19244,N_16704,N_17721);
nor U19245 (N_19245,N_18748,N_18505);
nor U19246 (N_19246,N_17378,N_16559);
or U19247 (N_19247,N_17333,N_17056);
nand U19248 (N_19248,N_17560,N_16565);
nor U19249 (N_19249,N_16655,N_17269);
nand U19250 (N_19250,N_16377,N_18010);
nor U19251 (N_19251,N_15957,N_18477);
nor U19252 (N_19252,N_17028,N_18293);
and U19253 (N_19253,N_18649,N_18193);
or U19254 (N_19254,N_16896,N_15907);
nand U19255 (N_19255,N_18692,N_18423);
and U19256 (N_19256,N_17278,N_15889);
or U19257 (N_19257,N_17404,N_16371);
and U19258 (N_19258,N_18457,N_17408);
or U19259 (N_19259,N_17291,N_18275);
nand U19260 (N_19260,N_18351,N_16541);
or U19261 (N_19261,N_18090,N_18435);
or U19262 (N_19262,N_17477,N_16680);
nor U19263 (N_19263,N_18151,N_17322);
nand U19264 (N_19264,N_18169,N_16062);
nand U19265 (N_19265,N_16612,N_18481);
or U19266 (N_19266,N_17148,N_18282);
or U19267 (N_19267,N_16076,N_16584);
or U19268 (N_19268,N_16284,N_18326);
and U19269 (N_19269,N_17853,N_15666);
and U19270 (N_19270,N_18182,N_16189);
and U19271 (N_19271,N_16436,N_16885);
or U19272 (N_19272,N_18718,N_17134);
and U19273 (N_19273,N_17398,N_17117);
nor U19274 (N_19274,N_15871,N_17891);
and U19275 (N_19275,N_18324,N_18192);
xor U19276 (N_19276,N_18720,N_17229);
nor U19277 (N_19277,N_17082,N_16160);
xnor U19278 (N_19278,N_15716,N_16461);
nand U19279 (N_19279,N_17726,N_18173);
and U19280 (N_19280,N_18309,N_16964);
or U19281 (N_19281,N_16170,N_17651);
nor U19282 (N_19282,N_17714,N_18705);
xnor U19283 (N_19283,N_15913,N_15884);
or U19284 (N_19284,N_16492,N_15726);
or U19285 (N_19285,N_16514,N_18156);
or U19286 (N_19286,N_16798,N_17843);
and U19287 (N_19287,N_16092,N_17277);
nand U19288 (N_19288,N_17223,N_18154);
nand U19289 (N_19289,N_15861,N_16536);
and U19290 (N_19290,N_16443,N_18343);
and U19291 (N_19291,N_18475,N_18138);
and U19292 (N_19292,N_17181,N_18380);
nor U19293 (N_19293,N_18567,N_18381);
nor U19294 (N_19294,N_17911,N_16692);
and U19295 (N_19295,N_17357,N_17249);
nor U19296 (N_19296,N_16550,N_17506);
and U19297 (N_19297,N_17461,N_16412);
or U19298 (N_19298,N_15968,N_17695);
nand U19299 (N_19299,N_18628,N_16552);
or U19300 (N_19300,N_16375,N_17632);
or U19301 (N_19301,N_16012,N_16378);
and U19302 (N_19302,N_17116,N_18744);
nor U19303 (N_19303,N_17955,N_17261);
or U19304 (N_19304,N_15779,N_16126);
nor U19305 (N_19305,N_17039,N_16606);
nor U19306 (N_19306,N_17770,N_15679);
nor U19307 (N_19307,N_17882,N_16185);
nor U19308 (N_19308,N_16796,N_17414);
xor U19309 (N_19309,N_17755,N_17954);
xor U19310 (N_19310,N_16978,N_16366);
nand U19311 (N_19311,N_18504,N_16993);
or U19312 (N_19312,N_16373,N_18747);
or U19313 (N_19313,N_17265,N_16034);
and U19314 (N_19314,N_17994,N_17317);
nand U19315 (N_19315,N_16178,N_16635);
or U19316 (N_19316,N_17946,N_16677);
and U19317 (N_19317,N_18356,N_16788);
xor U19318 (N_19318,N_17753,N_17820);
nand U19319 (N_19319,N_18115,N_16374);
or U19320 (N_19320,N_18486,N_17232);
nand U19321 (N_19321,N_15757,N_17733);
nand U19322 (N_19322,N_17866,N_17111);
nand U19323 (N_19323,N_17927,N_18150);
xnor U19324 (N_19324,N_16746,N_17316);
nor U19325 (N_19325,N_16433,N_17070);
nor U19326 (N_19326,N_18085,N_16467);
nand U19327 (N_19327,N_15794,N_16030);
or U19328 (N_19328,N_18337,N_18484);
and U19329 (N_19329,N_16909,N_15940);
nor U19330 (N_19330,N_16269,N_17840);
xor U19331 (N_19331,N_16959,N_18513);
or U19332 (N_19332,N_17149,N_18161);
or U19333 (N_19333,N_18015,N_17687);
or U19334 (N_19334,N_15637,N_17956);
and U19335 (N_19335,N_17517,N_17873);
and U19336 (N_19336,N_16233,N_17304);
xor U19337 (N_19337,N_17617,N_16791);
or U19338 (N_19338,N_16485,N_15879);
or U19339 (N_19339,N_16743,N_17172);
and U19340 (N_19340,N_17231,N_18414);
xnor U19341 (N_19341,N_18350,N_17677);
nor U19342 (N_19342,N_16152,N_15891);
nand U19343 (N_19343,N_17710,N_16566);
nor U19344 (N_19344,N_18181,N_16801);
or U19345 (N_19345,N_16887,N_18422);
and U19346 (N_19346,N_18706,N_16829);
xor U19347 (N_19347,N_18608,N_16438);
or U19348 (N_19348,N_18277,N_17286);
and U19349 (N_19349,N_17233,N_18474);
nand U19350 (N_19350,N_17865,N_15785);
and U19351 (N_19351,N_17752,N_16740);
or U19352 (N_19352,N_18454,N_16509);
nand U19353 (N_19353,N_16934,N_18727);
nand U19354 (N_19354,N_17985,N_18450);
and U19355 (N_19355,N_17279,N_16234);
or U19356 (N_19356,N_17550,N_18469);
and U19357 (N_19357,N_15825,N_18143);
or U19358 (N_19358,N_16875,N_16281);
nand U19359 (N_19359,N_17314,N_17652);
nand U19360 (N_19360,N_18444,N_16121);
xnor U19361 (N_19361,N_16877,N_17821);
nand U19362 (N_19362,N_15748,N_18299);
and U19363 (N_19363,N_17615,N_17984);
nand U19364 (N_19364,N_17128,N_16678);
or U19365 (N_19365,N_16894,N_18447);
and U19366 (N_19366,N_18586,N_17441);
and U19367 (N_19367,N_16953,N_17585);
xnor U19368 (N_19368,N_15919,N_15928);
or U19369 (N_19369,N_17979,N_15777);
and U19370 (N_19370,N_18663,N_18383);
and U19371 (N_19371,N_16597,N_16340);
nor U19372 (N_19372,N_15921,N_17185);
nor U19373 (N_19373,N_18096,N_16376);
xor U19374 (N_19374,N_16634,N_15693);
xnor U19375 (N_19375,N_17885,N_15712);
nand U19376 (N_19376,N_17173,N_17299);
nor U19377 (N_19377,N_17161,N_16480);
or U19378 (N_19378,N_17126,N_15626);
or U19379 (N_19379,N_15689,N_16408);
nand U19380 (N_19380,N_17059,N_16308);
and U19381 (N_19381,N_17780,N_18658);
nand U19382 (N_19382,N_18113,N_17284);
nand U19383 (N_19383,N_15698,N_17195);
and U19384 (N_19384,N_15655,N_16954);
or U19385 (N_19385,N_17835,N_15782);
and U19386 (N_19386,N_18723,N_18047);
nand U19387 (N_19387,N_17010,N_16397);
nor U19388 (N_19388,N_15934,N_16792);
or U19389 (N_19389,N_18292,N_17542);
xnor U19390 (N_19390,N_18331,N_18566);
or U19391 (N_19391,N_17788,N_15945);
or U19392 (N_19392,N_17037,N_16718);
nor U19393 (N_19393,N_18573,N_16813);
nand U19394 (N_19394,N_17639,N_17857);
nand U19395 (N_19395,N_18194,N_16944);
nor U19396 (N_19396,N_16040,N_18283);
or U19397 (N_19397,N_16360,N_16389);
nand U19398 (N_19398,N_18146,N_17572);
and U19399 (N_19399,N_16648,N_16291);
nand U19400 (N_19400,N_16974,N_17692);
xnor U19401 (N_19401,N_16947,N_18300);
or U19402 (N_19402,N_18404,N_16073);
and U19403 (N_19403,N_18714,N_18024);
nor U19404 (N_19404,N_15702,N_17766);
nand U19405 (N_19405,N_18210,N_18735);
and U19406 (N_19406,N_16405,N_17961);
nand U19407 (N_19407,N_17953,N_16864);
nor U19408 (N_19408,N_16426,N_16272);
nand U19409 (N_19409,N_18531,N_16581);
and U19410 (N_19410,N_15707,N_18555);
nand U19411 (N_19411,N_15699,N_16786);
nand U19412 (N_19412,N_18183,N_18147);
nor U19413 (N_19413,N_17425,N_16504);
or U19414 (N_19414,N_18304,N_18491);
and U19415 (N_19415,N_18538,N_17007);
or U19416 (N_19416,N_17599,N_17167);
xor U19417 (N_19417,N_16924,N_17534);
or U19418 (N_19418,N_17570,N_18451);
nand U19419 (N_19419,N_17744,N_17933);
or U19420 (N_19420,N_16435,N_16816);
and U19421 (N_19421,N_17204,N_18520);
and U19422 (N_19422,N_17694,N_16883);
and U19423 (N_19423,N_15972,N_17625);
and U19424 (N_19424,N_17199,N_16391);
nor U19425 (N_19425,N_17080,N_17230);
or U19426 (N_19426,N_17014,N_17340);
nor U19427 (N_19427,N_16226,N_17072);
nor U19428 (N_19428,N_16633,N_18362);
or U19429 (N_19429,N_17345,N_18570);
or U19430 (N_19430,N_16445,N_17087);
or U19431 (N_19431,N_16051,N_17405);
or U19432 (N_19432,N_18612,N_16478);
xnor U19433 (N_19433,N_16921,N_16965);
or U19434 (N_19434,N_16845,N_16625);
nand U19435 (N_19435,N_18149,N_16679);
nor U19436 (N_19436,N_15877,N_16424);
nand U19437 (N_19437,N_17892,N_17523);
nor U19438 (N_19438,N_17988,N_16580);
nand U19439 (N_19439,N_15875,N_18190);
or U19440 (N_19440,N_18252,N_18087);
nor U19441 (N_19441,N_16911,N_16860);
xnor U19442 (N_19442,N_17342,N_16931);
nand U19443 (N_19443,N_17036,N_16225);
nor U19444 (N_19444,N_16577,N_17027);
and U19445 (N_19445,N_18524,N_17175);
or U19446 (N_19446,N_16049,N_16714);
and U19447 (N_19447,N_18249,N_18372);
nand U19448 (N_19448,N_16935,N_18611);
nor U19449 (N_19449,N_16187,N_18215);
and U19450 (N_19450,N_16243,N_16620);
or U19451 (N_19451,N_18600,N_16162);
nor U19452 (N_19452,N_16930,N_18448);
and U19453 (N_19453,N_18139,N_17727);
nand U19454 (N_19454,N_17060,N_17545);
xnor U19455 (N_19455,N_18121,N_17970);
nor U19456 (N_19456,N_15970,N_17659);
nand U19457 (N_19457,N_15835,N_18375);
or U19458 (N_19458,N_16971,N_15864);
nor U19459 (N_19459,N_16238,N_17415);
and U19460 (N_19460,N_17614,N_18101);
and U19461 (N_19461,N_18643,N_16028);
nand U19462 (N_19462,N_15941,N_17896);
and U19463 (N_19463,N_15677,N_17581);
or U19464 (N_19464,N_16046,N_15737);
or U19465 (N_19465,N_16828,N_17627);
or U19466 (N_19466,N_15651,N_15962);
or U19467 (N_19467,N_17558,N_18051);
and U19468 (N_19468,N_15776,N_16107);
nand U19469 (N_19469,N_16593,N_17745);
or U19470 (N_19470,N_17680,N_18253);
nor U19471 (N_19471,N_16664,N_18031);
nand U19472 (N_19472,N_17868,N_16268);
and U19473 (N_19473,N_18700,N_17748);
nor U19474 (N_19474,N_16901,N_16484);
nor U19475 (N_19475,N_18184,N_18650);
or U19476 (N_19476,N_16555,N_16392);
and U19477 (N_19477,N_16605,N_15765);
nor U19478 (N_19478,N_16585,N_16417);
or U19479 (N_19479,N_17493,N_18268);
and U19480 (N_19480,N_18390,N_18008);
and U19481 (N_19481,N_15986,N_18110);
xor U19482 (N_19482,N_18604,N_17881);
or U19483 (N_19483,N_16945,N_18666);
xnor U19484 (N_19484,N_15710,N_17121);
nor U19485 (N_19485,N_17921,N_15633);
and U19486 (N_19486,N_16217,N_18683);
or U19487 (N_19487,N_16206,N_16199);
and U19488 (N_19488,N_18136,N_18379);
or U19489 (N_19489,N_17359,N_17422);
and U19490 (N_19490,N_16292,N_16912);
and U19491 (N_19491,N_18669,N_17122);
xnor U19492 (N_19492,N_17619,N_15831);
nor U19493 (N_19493,N_16483,N_17655);
and U19494 (N_19494,N_17457,N_18124);
and U19495 (N_19495,N_17052,N_17525);
nor U19496 (N_19496,N_17453,N_16948);
or U19497 (N_19497,N_17478,N_15802);
or U19498 (N_19498,N_18686,N_16583);
and U19499 (N_19499,N_17097,N_15703);
xnor U19500 (N_19500,N_18242,N_16088);
or U19501 (N_19501,N_16398,N_16673);
nor U19502 (N_19502,N_15904,N_18243);
nor U19503 (N_19503,N_18439,N_16619);
nor U19504 (N_19504,N_15749,N_16222);
nor U19505 (N_19505,N_16608,N_16694);
or U19506 (N_19506,N_16624,N_18741);
or U19507 (N_19507,N_17589,N_16457);
or U19508 (N_19508,N_15743,N_18731);
and U19509 (N_19509,N_17566,N_18678);
and U19510 (N_19510,N_18203,N_15949);
and U19511 (N_19511,N_17548,N_17924);
or U19512 (N_19512,N_16554,N_16946);
nand U19513 (N_19513,N_16870,N_15938);
nand U19514 (N_19514,N_17399,N_17260);
nor U19515 (N_19515,N_17749,N_16683);
nor U19516 (N_19516,N_18462,N_16300);
or U19517 (N_19517,N_17526,N_18311);
nor U19518 (N_19518,N_17412,N_18100);
or U19519 (N_19519,N_15869,N_16379);
nand U19520 (N_19520,N_16925,N_17634);
or U19521 (N_19521,N_16174,N_15939);
nand U19522 (N_19522,N_17666,N_17645);
nor U19523 (N_19523,N_18262,N_18013);
or U19524 (N_19524,N_15806,N_17867);
xor U19525 (N_19525,N_17934,N_18270);
nand U19526 (N_19526,N_16333,N_17633);
and U19527 (N_19527,N_16903,N_18672);
nor U19528 (N_19528,N_17569,N_15801);
nand U19529 (N_19529,N_15898,N_17237);
and U19530 (N_19530,N_17094,N_18446);
xnor U19531 (N_19531,N_16399,N_17641);
or U19532 (N_19532,N_16402,N_16726);
nand U19533 (N_19533,N_17830,N_18340);
or U19534 (N_19534,N_17372,N_16898);
and U19535 (N_19535,N_17363,N_18479);
nor U19536 (N_19536,N_16481,N_16181);
nand U19537 (N_19537,N_15687,N_15925);
nor U19538 (N_19538,N_15771,N_15670);
nor U19539 (N_19539,N_17434,N_15965);
or U19540 (N_19540,N_16986,N_17794);
or U19541 (N_19541,N_16384,N_15860);
nand U19542 (N_19542,N_15745,N_17043);
or U19543 (N_19543,N_16817,N_17076);
nor U19544 (N_19544,N_18039,N_17463);
nor U19545 (N_19545,N_16643,N_17382);
nor U19546 (N_19546,N_18079,N_17160);
or U19547 (N_19547,N_17123,N_17567);
and U19548 (N_19548,N_18248,N_16055);
nand U19549 (N_19549,N_16561,N_18614);
nand U19550 (N_19550,N_15722,N_17613);
and U19551 (N_19551,N_18465,N_17912);
and U19552 (N_19552,N_17439,N_17464);
or U19553 (N_19553,N_16116,N_16549);
nor U19554 (N_19554,N_15660,N_15795);
and U19555 (N_19555,N_16316,N_15981);
or U19556 (N_19556,N_17803,N_16834);
or U19557 (N_19557,N_18739,N_15979);
and U19558 (N_19558,N_16985,N_17218);
nand U19559 (N_19559,N_17797,N_18449);
nand U19560 (N_19560,N_16821,N_17385);
nor U19561 (N_19561,N_18320,N_16721);
or U19562 (N_19562,N_17436,N_18104);
and U19563 (N_19563,N_15858,N_17644);
nand U19564 (N_19564,N_16674,N_16914);
and U19565 (N_19565,N_16818,N_17728);
nand U19566 (N_19566,N_16115,N_16395);
xor U19567 (N_19567,N_17388,N_17497);
nor U19568 (N_19568,N_16956,N_17470);
nor U19569 (N_19569,N_17987,N_17266);
or U19570 (N_19570,N_18561,N_18021);
nand U19571 (N_19571,N_17257,N_17120);
or U19572 (N_19572,N_16720,N_18086);
nor U19573 (N_19573,N_17214,N_18634);
or U19574 (N_19574,N_17203,N_16723);
nand U19575 (N_19575,N_18582,N_18062);
nor U19576 (N_19576,N_16797,N_17724);
or U19577 (N_19577,N_18290,N_17397);
or U19578 (N_19578,N_17219,N_17227);
xor U19579 (N_19579,N_15724,N_16771);
nand U19580 (N_19580,N_15953,N_17928);
or U19581 (N_19581,N_17256,N_16183);
nand U19582 (N_19582,N_17907,N_15671);
xnor U19583 (N_19583,N_18257,N_16516);
or U19584 (N_19584,N_17959,N_17423);
and U19585 (N_19585,N_17977,N_17552);
nand U19586 (N_19586,N_16101,N_17193);
nand U19587 (N_19587,N_17900,N_16918);
or U19588 (N_19588,N_17812,N_17490);
or U19589 (N_19589,N_17875,N_16902);
nor U19590 (N_19590,N_16041,N_18746);
and U19591 (N_19591,N_18227,N_18557);
or U19592 (N_19592,N_15881,N_16522);
nor U19593 (N_19593,N_16142,N_18434);
and U19594 (N_19594,N_16927,N_15634);
xnor U19595 (N_19595,N_18082,N_17467);
or U19596 (N_19596,N_15920,N_15999);
and U19597 (N_19597,N_16184,N_16749);
and U19598 (N_19598,N_15800,N_17894);
nand U19599 (N_19599,N_18483,N_16889);
or U19600 (N_19600,N_16631,N_16707);
nand U19601 (N_19601,N_15752,N_18261);
xor U19602 (N_19602,N_16513,N_16731);
nor U19603 (N_19603,N_17323,N_15824);
nor U19604 (N_19604,N_18631,N_18722);
and U19605 (N_19605,N_18426,N_18622);
nor U19606 (N_19606,N_17096,N_16014);
nor U19607 (N_19607,N_18421,N_16388);
and U19608 (N_19608,N_15909,N_17717);
nor U19609 (N_19609,N_16609,N_16904);
nor U19610 (N_19610,N_18341,N_16803);
nand U19611 (N_19611,N_16752,N_16763);
xor U19612 (N_19612,N_17152,N_18164);
nand U19613 (N_19613,N_17498,N_17711);
and U19614 (N_19614,N_15755,N_18523);
xnor U19615 (N_19615,N_15668,N_16949);
nor U19616 (N_19616,N_18228,N_17328);
xor U19617 (N_19617,N_17403,N_17078);
nor U19618 (N_19618,N_18437,N_18438);
nand U19619 (N_19619,N_16510,N_16859);
nor U19620 (N_19620,N_18323,N_17878);
nor U19621 (N_19621,N_18014,N_16880);
xor U19622 (N_19622,N_18581,N_18517);
and U19623 (N_19623,N_16793,N_17302);
and U19624 (N_19624,N_16267,N_17704);
nand U19625 (N_19625,N_16917,N_18550);
nor U19626 (N_19626,N_15893,N_15639);
and U19627 (N_19627,N_16961,N_18460);
and U19628 (N_19628,N_15947,N_17190);
nor U19629 (N_19629,N_17511,N_15718);
and U19630 (N_19630,N_15888,N_18453);
and U19631 (N_19631,N_17626,N_17485);
nand U19632 (N_19632,N_15658,N_18595);
or U19633 (N_19633,N_16735,N_15665);
or U19634 (N_19634,N_17640,N_18654);
xor U19635 (N_19635,N_18132,N_16105);
or U19636 (N_19636,N_16662,N_17420);
and U19637 (N_19637,N_18123,N_17965);
and U19638 (N_19638,N_18276,N_16744);
or U19639 (N_19639,N_17879,N_18305);
nor U19640 (N_19640,N_17556,N_17575);
xor U19641 (N_19641,N_16963,N_18740);
and U19642 (N_19642,N_17079,N_16191);
and U19643 (N_19643,N_16668,N_16713);
nand U19644 (N_19644,N_17541,N_18734);
xor U19645 (N_19645,N_18514,N_15817);
and U19646 (N_19646,N_15851,N_16108);
or U19647 (N_19647,N_17529,N_17675);
and U19648 (N_19648,N_16059,N_17958);
or U19649 (N_19649,N_18492,N_17496);
nand U19650 (N_19650,N_15759,N_18133);
nand U19651 (N_19651,N_17446,N_18519);
nor U19652 (N_19652,N_18237,N_15742);
nand U19653 (N_19653,N_17132,N_16895);
and U19654 (N_19654,N_15662,N_16106);
nand U19655 (N_19655,N_15930,N_17006);
or U19656 (N_19656,N_17180,N_17904);
nand U19657 (N_19657,N_17685,N_17877);
nand U19658 (N_19658,N_18059,N_16472);
nor U19659 (N_19659,N_16381,N_16506);
nor U19660 (N_19660,N_16955,N_16545);
and U19661 (N_19661,N_17200,N_17312);
and U19662 (N_19662,N_17779,N_17013);
or U19663 (N_19663,N_16001,N_17029);
nor U19664 (N_19664,N_18068,N_16745);
or U19665 (N_19665,N_15998,N_16962);
nor U19666 (N_19666,N_15980,N_17245);
and U19667 (N_19667,N_16530,N_17475);
nor U19668 (N_19668,N_18126,N_18711);
xor U19669 (N_19669,N_18441,N_15878);
and U19670 (N_19670,N_16307,N_16695);
nand U19671 (N_19671,N_18730,N_17057);
and U19672 (N_19672,N_17841,N_17026);
and U19673 (N_19673,N_18704,N_18548);
and U19674 (N_19674,N_18508,N_16876);
nand U19675 (N_19675,N_18050,N_16444);
or U19676 (N_19676,N_16180,N_16982);
nand U19677 (N_19677,N_17285,N_17426);
nor U19678 (N_19678,N_18036,N_17851);
and U19679 (N_19679,N_16751,N_16776);
nand U19680 (N_19680,N_15814,N_16286);
or U19681 (N_19681,N_16665,N_16576);
and U19682 (N_19682,N_16697,N_17630);
or U19683 (N_19683,N_17682,N_16454);
nor U19684 (N_19684,N_18335,N_16216);
and U19685 (N_19685,N_17442,N_15874);
and U19686 (N_19686,N_16163,N_15856);
nor U19687 (N_19687,N_17471,N_17021);
nor U19688 (N_19688,N_17786,N_18312);
nor U19689 (N_19689,N_17801,N_16298);
nand U19690 (N_19690,N_17902,N_16647);
nand U19691 (N_19691,N_16636,N_16223);
or U19692 (N_19692,N_18591,N_18273);
nor U19693 (N_19693,N_17968,N_17311);
and U19694 (N_19694,N_16610,N_15841);
and U19695 (N_19695,N_16321,N_17428);
and U19696 (N_19696,N_17616,N_17192);
or U19697 (N_19697,N_18429,N_15797);
or U19698 (N_19698,N_17191,N_17487);
or U19699 (N_19699,N_18606,N_16410);
and U19700 (N_19700,N_16873,N_16254);
or U19701 (N_19701,N_15761,N_15675);
and U19702 (N_19702,N_17889,N_17649);
nand U19703 (N_19703,N_18075,N_16459);
nand U19704 (N_19704,N_16274,N_18532);
nand U19705 (N_19705,N_16328,N_17135);
nand U19706 (N_19706,N_17553,N_17762);
nor U19707 (N_19707,N_17396,N_17859);
or U19708 (N_19708,N_17307,N_17804);
nor U19709 (N_19709,N_16712,N_18418);
nand U19710 (N_19710,N_18560,N_17406);
nor U19711 (N_19711,N_16615,N_16064);
or U19712 (N_19712,N_17564,N_17624);
xnor U19713 (N_19713,N_16218,N_18496);
or U19714 (N_19714,N_17110,N_16795);
xor U19715 (N_19715,N_16065,N_18128);
nor U19716 (N_19716,N_17170,N_17750);
nor U19717 (N_19717,N_17051,N_17501);
nor U19718 (N_19718,N_18250,N_18488);
nor U19719 (N_19719,N_18295,N_17292);
nor U19720 (N_19720,N_16411,N_18109);
nand U19721 (N_19721,N_17951,N_16640);
or U19722 (N_19722,N_16063,N_17538);
and U19723 (N_19723,N_16171,N_18172);
nor U19724 (N_19724,N_17354,N_17334);
xnor U19725 (N_19725,N_18392,N_17366);
or U19726 (N_19726,N_17729,N_15872);
and U19727 (N_19727,N_17220,N_16361);
and U19728 (N_19728,N_16081,N_17437);
and U19729 (N_19729,N_16724,N_17708);
xnor U19730 (N_19730,N_18443,N_15873);
or U19731 (N_19731,N_16290,N_18616);
and U19732 (N_19732,N_15951,N_15905);
or U19733 (N_19733,N_16111,N_16822);
or U19734 (N_19734,N_16058,N_16156);
and U19735 (N_19735,N_16528,N_16002);
or U19736 (N_19736,N_17301,N_16874);
nand U19737 (N_19737,N_16866,N_16271);
or U19738 (N_19738,N_17527,N_16151);
nor U19739 (N_19739,N_15844,N_17273);
nand U19740 (N_19740,N_17716,N_17482);
nand U19741 (N_19741,N_17699,N_18673);
nor U19742 (N_19742,N_16696,N_16741);
or U19743 (N_19743,N_16779,N_17168);
nor U19744 (N_19744,N_17090,N_16709);
nor U19745 (N_19745,N_17451,N_15932);
xor U19746 (N_19746,N_18005,N_16910);
nand U19747 (N_19747,N_17336,N_16820);
nand U19748 (N_19748,N_16098,N_16332);
nand U19749 (N_19749,N_16479,N_17819);
xnor U19750 (N_19750,N_16558,N_18386);
or U19751 (N_19751,N_17679,N_18733);
nor U19752 (N_19752,N_18105,N_15845);
nand U19753 (N_19753,N_18196,N_17319);
or U19754 (N_19754,N_16835,N_17491);
and U19755 (N_19755,N_16339,N_17862);
xnor U19756 (N_19756,N_17929,N_17244);
xor U19757 (N_19757,N_17306,N_17943);
or U19758 (N_19758,N_18625,N_16228);
or U19759 (N_19759,N_16700,N_17844);
nand U19760 (N_19760,N_17224,N_17598);
nand U19761 (N_19761,N_16871,N_15653);
nor U19762 (N_19762,N_18525,N_18165);
and U19763 (N_19763,N_18076,N_18303);
nor U19764 (N_19764,N_17174,N_17577);
nand U19765 (N_19765,N_15997,N_16276);
nor U19766 (N_19766,N_16632,N_16229);
xnor U19767 (N_19767,N_17847,N_18701);
or U19768 (N_19768,N_15819,N_18294);
or U19769 (N_19769,N_18073,N_18621);
or U19770 (N_19770,N_15876,N_18028);
nor U19771 (N_19771,N_15960,N_16293);
nor U19772 (N_19772,N_17217,N_16453);
nand U19773 (N_19773,N_15783,N_18102);
nor U19774 (N_19774,N_17537,N_15627);
or U19775 (N_19775,N_17602,N_18539);
nor U19776 (N_19776,N_17824,N_16326);
nor U19777 (N_19777,N_17379,N_17686);
nor U19778 (N_19778,N_18354,N_17410);
nand U19779 (N_19779,N_18093,N_15826);
or U19780 (N_19780,N_15680,N_17212);
nand U19781 (N_19781,N_17503,N_18130);
nor U19782 (N_19782,N_17263,N_17041);
and U19783 (N_19783,N_17274,N_16508);
nand U19784 (N_19784,N_16013,N_18626);
nor U19785 (N_19785,N_17730,N_18640);
or U19786 (N_19786,N_18424,N_18467);
nor U19787 (N_19787,N_17500,N_18627);
nor U19788 (N_19788,N_17005,N_18680);
and U19789 (N_19789,N_18659,N_17210);
and U19790 (N_19790,N_17664,N_16450);
nand U19791 (N_19791,N_18034,N_17023);
or U19792 (N_19792,N_17785,N_16197);
nor U19793 (N_19793,N_17321,N_18026);
or U19794 (N_19794,N_16754,N_15917);
nand U19795 (N_19795,N_18385,N_18646);
or U19796 (N_19796,N_16026,N_17715);
xnor U19797 (N_19797,N_16221,N_15833);
and U19798 (N_19798,N_16838,N_15923);
nor U19799 (N_19799,N_17952,N_17712);
nand U19800 (N_19800,N_15706,N_18395);
xnor U19801 (N_19801,N_17583,N_17081);
and U19802 (N_19802,N_17075,N_16737);
nor U19803 (N_19803,N_17158,N_17930);
nand U19804 (N_19804,N_16077,N_16247);
or U19805 (N_19805,N_16463,N_17067);
or U19806 (N_19806,N_16000,N_18363);
and U19807 (N_19807,N_16175,N_17502);
nor U19808 (N_19808,N_18052,N_18499);
nand U19809 (N_19809,N_16025,N_16248);
nand U19810 (N_19810,N_15859,N_16331);
nor U19811 (N_19811,N_18607,N_17972);
nand U19812 (N_19812,N_17607,N_17691);
nand U19813 (N_19813,N_17702,N_16732);
nand U19814 (N_19814,N_18401,N_16304);
xnor U19815 (N_19815,N_17196,N_17648);
nor U19816 (N_19816,N_16169,N_17957);
nor U19817 (N_19817,N_16660,N_18092);
nand U19818 (N_19818,N_18674,N_16344);
nor U19819 (N_19819,N_18180,N_17222);
or U19820 (N_19820,N_17671,N_16079);
and U19821 (N_19821,N_17162,N_15723);
nand U19822 (N_19822,N_16734,N_16666);
and U19823 (N_19823,N_18057,N_16434);
or U19824 (N_19824,N_18342,N_16460);
nand U19825 (N_19825,N_18023,N_15764);
nand U19826 (N_19826,N_18020,N_17735);
nor U19827 (N_19827,N_17295,N_17949);
nor U19828 (N_19828,N_15719,N_16736);
nor U19829 (N_19829,N_15730,N_15816);
nand U19830 (N_19830,N_17684,N_18302);
nor U19831 (N_19831,N_17103,N_15713);
or U19832 (N_19832,N_16023,N_16124);
nor U19833 (N_19833,N_16759,N_17084);
xor U19834 (N_19834,N_17016,N_17983);
nand U19835 (N_19835,N_17981,N_16355);
and U19836 (N_19836,N_16167,N_18040);
and U19837 (N_19837,N_17063,N_17999);
nand U19838 (N_19838,N_16257,N_17621);
nand U19839 (N_19839,N_17807,N_17828);
or U19840 (N_19840,N_17698,N_15781);
nor U19841 (N_19841,N_16711,N_15732);
nand U19842 (N_19842,N_18098,N_18159);
or U19843 (N_19843,N_17754,N_18624);
nand U19844 (N_19844,N_16095,N_16867);
nor U19845 (N_19845,N_15867,N_16252);
and U19846 (N_19846,N_16085,N_16984);
nand U19847 (N_19847,N_17413,N_16165);
nor U19848 (N_19848,N_16783,N_17863);
and U19849 (N_19849,N_16782,N_18665);
nand U19850 (N_19850,N_17044,N_18278);
or U19851 (N_19851,N_17880,N_16858);
nand U19852 (N_19852,N_16574,N_18084);
xor U19853 (N_19853,N_16757,N_16349);
nor U19854 (N_19854,N_18061,N_16539);
or U19855 (N_19855,N_16507,N_17251);
or U19856 (N_19856,N_15789,N_18633);
or U19857 (N_19857,N_18471,N_17456);
or U19858 (N_19858,N_17387,N_17530);
and U19859 (N_19859,N_16471,N_16056);
nor U19860 (N_19860,N_16706,N_18396);
or U19861 (N_19861,N_17280,N_16899);
or U19862 (N_19862,N_18682,N_17318);
and U19863 (N_19863,N_16130,N_16306);
and U19864 (N_19864,N_17093,N_17164);
or U19865 (N_19865,N_16150,N_17184);
nor U19866 (N_19866,N_17032,N_16256);
nand U19867 (N_19867,N_16317,N_18187);
and U19868 (N_19868,N_17813,N_17178);
nor U19869 (N_19869,N_16919,N_17113);
xor U19870 (N_19870,N_16684,N_16313);
and U19871 (N_19871,N_17657,N_18503);
and U19872 (N_19872,N_17734,N_17107);
nand U19873 (N_19873,N_17759,N_16586);
xor U19874 (N_19874,N_18000,N_18301);
xnor U19875 (N_19875,N_16227,N_16356);
xnor U19876 (N_19876,N_16651,N_17443);
nand U19877 (N_19877,N_15892,N_16841);
xnor U19878 (N_19878,N_17209,N_16261);
and U19879 (N_19879,N_17690,N_16670);
xnor U19880 (N_19880,N_16637,N_15842);
or U19881 (N_19881,N_17638,N_16511);
nor U19882 (N_19882,N_18671,N_16324);
and U19883 (N_19883,N_17893,N_18251);
nand U19884 (N_19884,N_18029,N_16120);
and U19885 (N_19885,N_16441,N_16907);
nor U19886 (N_19886,N_15936,N_17392);
or U19887 (N_19887,N_15647,N_18288);
or U19888 (N_19888,N_16249,N_17597);
nand U19889 (N_19889,N_18344,N_17137);
or U19890 (N_19890,N_17587,N_16928);
nand U19891 (N_19891,N_16367,N_16802);
nand U19892 (N_19892,N_18221,N_17400);
nand U19893 (N_19893,N_16560,N_18574);
nor U19894 (N_19894,N_16020,N_17596);
and U19895 (N_19895,N_16494,N_16730);
nand U19896 (N_19896,N_18564,N_16981);
nand U19897 (N_19897,N_17064,N_17494);
nand U19898 (N_19898,N_17049,N_16236);
or U19899 (N_19899,N_18609,N_18411);
nand U19900 (N_19900,N_16992,N_17931);
and U19901 (N_19901,N_15747,N_18171);
and U19902 (N_19902,N_16811,N_18066);
nand U19903 (N_19903,N_17777,N_18236);
nand U19904 (N_19904,N_17521,N_18593);
nor U19905 (N_19905,N_17883,N_16800);
or U19906 (N_19906,N_15822,N_17142);
xor U19907 (N_19907,N_17046,N_18348);
or U19908 (N_19908,N_17254,N_16951);
or U19909 (N_19909,N_16050,N_17742);
nand U19910 (N_19910,N_17129,N_16578);
nand U19911 (N_19911,N_16535,N_17047);
or U19912 (N_19912,N_18202,N_17095);
xnor U19913 (N_19913,N_17335,N_18022);
or U19914 (N_19914,N_16428,N_17102);
and U19915 (N_19915,N_17421,N_17243);
nor U19916 (N_19916,N_17384,N_16710);
and U19917 (N_19917,N_16258,N_17910);
and U19918 (N_19918,N_17998,N_17432);
and U19919 (N_19919,N_16335,N_17601);
nor U19920 (N_19920,N_18212,N_17364);
nor U19921 (N_19921,N_18645,N_18698);
nand U19922 (N_19922,N_16672,N_16922);
nor U19923 (N_19923,N_17969,N_16416);
and U19924 (N_19924,N_17401,N_15628);
nand U19925 (N_19925,N_16007,N_17793);
nand U19926 (N_19926,N_17592,N_18592);
nor U19927 (N_19927,N_18394,N_18245);
nand U19928 (N_19928,N_17236,N_18613);
xnor U19929 (N_19929,N_16242,N_18526);
or U19930 (N_19930,N_16224,N_16137);
or U19931 (N_19931,N_18231,N_16493);
nor U19932 (N_19932,N_16468,N_17239);
xnor U19933 (N_19933,N_17792,N_15885);
nand U19934 (N_19934,N_18461,N_16589);
nor U19935 (N_19935,N_18487,N_18359);
and U19936 (N_19936,N_17890,N_17344);
and U19937 (N_19937,N_17871,N_16689);
and U19938 (N_19938,N_16869,N_16521);
xnor U19939 (N_19939,N_18065,N_18738);
or U19940 (N_19940,N_17157,N_15629);
and U19941 (N_19941,N_18594,N_15681);
and U19942 (N_19942,N_16287,N_15990);
nor U19943 (N_19943,N_17100,N_18042);
xor U19944 (N_19944,N_15734,N_18393);
nand U19945 (N_19945,N_15840,N_15709);
nor U19946 (N_19946,N_16033,N_16403);
nor U19947 (N_19947,N_15773,N_15944);
nand U19948 (N_19948,N_16906,N_17774);
nand U19949 (N_19949,N_15760,N_16503);
xor U19950 (N_19950,N_18374,N_17776);
and U19951 (N_19951,N_16322,N_18279);
nand U19952 (N_19952,N_17073,N_16650);
nor U19953 (N_19953,N_18632,N_17989);
nor U19954 (N_19954,N_16579,N_17228);
or U19955 (N_19955,N_16844,N_17226);
or U19956 (N_19956,N_15918,N_17973);
or U19957 (N_19957,N_17159,N_16888);
and U19958 (N_19958,N_17656,N_15678);
and U19959 (N_19959,N_17002,N_17347);
or U19960 (N_19960,N_17017,N_16733);
or U19961 (N_19961,N_16250,N_15667);
nand U19962 (N_19962,N_16996,N_15811);
nand U19963 (N_19963,N_18188,N_16131);
or U19964 (N_19964,N_18369,N_18470);
xor U19965 (N_19965,N_15664,N_16253);
or U19966 (N_19966,N_15673,N_18198);
nand U19967 (N_19967,N_16517,N_16277);
or U19968 (N_19968,N_17492,N_16008);
and U19969 (N_19969,N_18442,N_16717);
xor U19970 (N_19970,N_16192,N_16464);
nand U19971 (N_19971,N_17416,N_16342);
nand U19972 (N_19972,N_15933,N_16932);
or U19973 (N_19973,N_15787,N_17300);
and U19974 (N_19974,N_16500,N_17297);
or U19975 (N_19975,N_15808,N_17565);
or U19976 (N_19976,N_16594,N_17153);
and U19977 (N_19977,N_16900,N_17150);
or U19978 (N_19978,N_17507,N_17849);
nor U19979 (N_19979,N_17009,N_16303);
nor U19980 (N_19980,N_17352,N_17838);
or U19981 (N_19981,N_18515,N_17489);
nor U19982 (N_19982,N_18152,N_17402);
nand U19983 (N_19983,N_15886,N_15974);
nor U19984 (N_19984,N_15694,N_15715);
xnor U19985 (N_19985,N_18346,N_18427);
or U19986 (N_19986,N_17848,N_18501);
nand U19987 (N_19987,N_16851,N_16839);
and U19988 (N_19988,N_15912,N_17595);
nor U19989 (N_19989,N_16531,N_16440);
nor U19990 (N_19990,N_16138,N_18256);
or U19991 (N_19991,N_15676,N_16515);
nand U19992 (N_19992,N_16260,N_17915);
or U19993 (N_19993,N_17561,N_16006);
nand U19994 (N_19994,N_17852,N_18373);
nand U19995 (N_19995,N_17874,N_16826);
and U19996 (N_19996,N_16972,N_16207);
nor U19997 (N_19997,N_16141,N_15903);
xnor U19998 (N_19998,N_16215,N_18258);
xnor U19999 (N_19999,N_17338,N_18585);
or U20000 (N_20000,N_16488,N_17963);
nand U20001 (N_20001,N_18576,N_17703);
or U20002 (N_20002,N_18353,N_18111);
or U20003 (N_20003,N_15721,N_15857);
xor U20004 (N_20004,N_17719,N_18291);
nand U20005 (N_20005,N_17077,N_15654);
xor U20006 (N_20006,N_16353,N_16654);
xor U20007 (N_20007,N_15827,N_17433);
nor U20008 (N_20008,N_16868,N_18142);
nand U20009 (N_20009,N_18717,N_18482);
nor U20010 (N_20010,N_18623,N_17033);
and U20011 (N_20011,N_16719,N_16038);
nand U20012 (N_20012,N_18332,N_18452);
nor U20013 (N_20013,N_17817,N_18120);
nand U20014 (N_20014,N_18260,N_18009);
nor U20015 (N_20015,N_17001,N_17738);
and U20016 (N_20016,N_17709,N_16551);
nor U20017 (N_20017,N_17373,N_18431);
nand U20018 (N_20018,N_18347,N_18382);
nand U20019 (N_20019,N_16177,N_17207);
nor U20020 (N_20020,N_17832,N_17950);
nand U20021 (N_20021,N_17935,N_17676);
and U20022 (N_20022,N_17324,N_15982);
nor U20023 (N_20023,N_18255,N_18201);
nor U20024 (N_20024,N_16423,N_17393);
and U20025 (N_20025,N_18271,N_15812);
nor U20026 (N_20026,N_17114,N_16053);
or U20027 (N_20027,N_18587,N_17637);
nand U20028 (N_20028,N_18134,N_18254);
or U20029 (N_20029,N_16119,N_18425);
nand U20030 (N_20030,N_17573,N_18234);
and U20031 (N_20031,N_17678,N_16764);
and U20032 (N_20032,N_16311,N_18575);
and U20033 (N_20033,N_15772,N_15915);
nand U20034 (N_20034,N_16747,N_15672);
nand U20035 (N_20035,N_16990,N_16235);
or U20036 (N_20036,N_18602,N_17736);
and U20037 (N_20037,N_17429,N_18103);
and U20038 (N_20038,N_16296,N_17085);
and U20039 (N_20039,N_17374,N_15922);
nor U20040 (N_20040,N_16937,N_17568);
nor U20041 (N_20041,N_17182,N_18530);
xnor U20042 (N_20042,N_17417,N_16135);
nor U20043 (N_20043,N_18552,N_17131);
and U20044 (N_20044,N_18590,N_16595);
and U20045 (N_20045,N_16762,N_18537);
nand U20046 (N_20046,N_17089,N_17547);
xor U20047 (N_20047,N_17309,N_17756);
and U20048 (N_20048,N_15750,N_16048);
xor U20049 (N_20049,N_16969,N_18338);
xnor U20050 (N_20050,N_16891,N_16086);
nor U20051 (N_20051,N_17909,N_16143);
nand U20052 (N_20052,N_16681,N_17370);
or U20053 (N_20053,N_16502,N_16190);
or U20054 (N_20054,N_17205,N_17697);
nand U20055 (N_20055,N_16970,N_16425);
or U20056 (N_20056,N_16699,N_18725);
and U20057 (N_20057,N_15697,N_17253);
or U20058 (N_20058,N_18728,N_18702);
and U20059 (N_20059,N_17612,N_17169);
nand U20060 (N_20060,N_16275,N_16708);
nand U20061 (N_20061,N_18265,N_16149);
nor U20062 (N_20062,N_16773,N_17272);
and U20063 (N_20063,N_18054,N_15908);
nor U20064 (N_20064,N_17673,N_17133);
or U20065 (N_20065,N_17074,N_15837);
and U20066 (N_20066,N_16761,N_16527);
xnor U20067 (N_20067,N_15799,N_16466);
or U20068 (N_20068,N_15963,N_17814);
or U20069 (N_20069,N_16401,N_16409);
nand U20070 (N_20070,N_18240,N_18580);
xor U20071 (N_20071,N_17960,N_17165);
xnor U20072 (N_20072,N_18144,N_17782);
or U20073 (N_20073,N_17369,N_17784);
nand U20074 (N_20074,N_16915,N_18259);
or U20075 (N_20075,N_15686,N_15640);
xnor U20076 (N_20076,N_17554,N_17683);
nand U20077 (N_20077,N_16200,N_17308);
or U20078 (N_20078,N_17829,N_15850);
or U20079 (N_20079,N_17146,N_15638);
xnor U20080 (N_20080,N_18551,N_18141);
or U20081 (N_20081,N_18410,N_16520);
and U20082 (N_20082,N_16237,N_16161);
nand U20083 (N_20083,N_16843,N_18241);
nor U20084 (N_20084,N_15931,N_16212);
and U20085 (N_20085,N_18064,N_16305);
nand U20086 (N_20086,N_17281,N_16604);
or U20087 (N_20087,N_18027,N_16084);
nand U20088 (N_20088,N_16262,N_18521);
nand U20089 (N_20089,N_16154,N_16750);
nand U20090 (N_20090,N_17119,N_16219);
nor U20091 (N_20091,N_17305,N_16128);
and U20092 (N_20092,N_17294,N_15769);
nand U20093 (N_20093,N_17917,N_18389);
or U20094 (N_20094,N_18116,N_16775);
nor U20095 (N_20095,N_18639,N_16147);
and U20096 (N_20096,N_16117,N_16572);
nand U20097 (N_20097,N_16347,N_18272);
nor U20098 (N_20098,N_18412,N_17922);
and U20099 (N_20099,N_17557,N_18719);
nand U20100 (N_20100,N_18371,N_18546);
nand U20101 (N_20101,N_17019,N_17720);
xnor U20102 (N_20102,N_17145,N_17332);
nor U20103 (N_20103,N_17903,N_17313);
nor U20104 (N_20104,N_16273,N_18360);
nor U20105 (N_20105,N_17563,N_16382);
and U20106 (N_20106,N_15731,N_16548);
or U20107 (N_20107,N_18137,N_16758);
nor U20108 (N_20108,N_17536,N_17535);
nor U20109 (N_20109,N_18333,N_18490);
nor U20110 (N_20110,N_17315,N_17351);
nand U20111 (N_20111,N_16645,N_15935);
or U20112 (N_20112,N_16623,N_15786);
or U20113 (N_20113,N_15952,N_18213);
nor U20114 (N_20114,N_15855,N_17603);
nand U20115 (N_20115,N_18030,N_18516);
or U20116 (N_20116,N_17474,N_16882);
or U20117 (N_20117,N_18599,N_16602);
or U20118 (N_20118,N_17975,N_16172);
or U20119 (N_20119,N_17746,N_17386);
xor U20120 (N_20120,N_17144,N_17763);
or U20121 (N_20121,N_16865,N_16600);
or U20122 (N_20122,N_17574,N_16765);
nand U20123 (N_20123,N_17514,N_16794);
or U20124 (N_20124,N_18636,N_17156);
nor U20125 (N_20125,N_16089,N_18319);
nand U20126 (N_20126,N_15849,N_16809);
nand U20127 (N_20127,N_17739,N_17528);
nand U20128 (N_20128,N_17555,N_16057);
or U20129 (N_20129,N_17576,N_17806);
and U20130 (N_20130,N_17608,N_16575);
and U20131 (N_20131,N_16698,N_16024);
and U20132 (N_20132,N_17532,N_17394);
or U20133 (N_20133,N_17823,N_18357);
and U20134 (N_20134,N_17055,N_18420);
nor U20135 (N_20135,N_17643,N_17938);
nand U20136 (N_20136,N_18208,N_18601);
nand U20137 (N_20137,N_15902,N_16950);
nand U20138 (N_20138,N_16487,N_15978);
or U20139 (N_20139,N_18432,N_16362);
nor U20140 (N_20140,N_17996,N_16853);
nand U20141 (N_20141,N_17267,N_16134);
nor U20142 (N_20142,N_16989,N_17258);
nand U20143 (N_20143,N_18244,N_18667);
xnor U20144 (N_20144,N_16380,N_18743);
nand U20145 (N_20145,N_15625,N_17250);
xor U20146 (N_20146,N_18217,N_17974);
nor U20147 (N_20147,N_15674,N_17326);
nor U20148 (N_20148,N_17343,N_16933);
nor U20149 (N_20149,N_17722,N_17787);
and U20150 (N_20150,N_18387,N_17447);
and U20151 (N_20151,N_17065,N_16729);
and U20152 (N_20152,N_15740,N_17646);
nor U20153 (N_20153,N_16686,N_17105);
nor U20154 (N_20154,N_17580,N_18684);
or U20155 (N_20155,N_16831,N_18458);
or U20156 (N_20156,N_18069,N_15766);
nor U20157 (N_20157,N_16847,N_16176);
and U20158 (N_20158,N_17141,N_17176);
nor U20159 (N_20159,N_17551,N_17469);
nand U20160 (N_20160,N_16427,N_17546);
and U20161 (N_20161,N_17628,N_18378);
nor U20162 (N_20162,N_15853,N_16113);
and U20163 (N_20163,N_17816,N_18617);
or U20164 (N_20164,N_16330,N_18041);
and U20165 (N_20165,N_16429,N_18618);
and U20166 (N_20166,N_16742,N_16547);
nor U20167 (N_20167,N_18117,N_16564);
and U20168 (N_20168,N_18584,N_15995);
nand U20169 (N_20169,N_16518,N_16642);
nand U20170 (N_20170,N_16299,N_16588);
or U20171 (N_20171,N_17740,N_16067);
and U20172 (N_20172,N_16596,N_17600);
nand U20173 (N_20173,N_18408,N_16846);
and U20174 (N_20174,N_17355,N_16526);
nor U20175 (N_20175,N_18207,N_17136);
nor U20176 (N_20176,N_15630,N_18493);
or U20177 (N_20177,N_18296,N_17864);
nor U20178 (N_20178,N_16018,N_18043);
and U20179 (N_20179,N_16213,N_16016);
and U20180 (N_20180,N_16772,N_16537);
nand U20181 (N_20181,N_15733,N_18635);
nand U20182 (N_20182,N_18223,N_16078);
or U20183 (N_20183,N_18091,N_16280);
or U20184 (N_20184,N_17765,N_16770);
and U20185 (N_20185,N_17642,N_15818);
xnor U20186 (N_20186,N_17360,N_16159);
or U20187 (N_20187,N_16540,N_16553);
or U20188 (N_20188,N_17488,N_15645);
or U20189 (N_20189,N_16715,N_17177);
nand U20190 (N_20190,N_15887,N_18459);
nand U20191 (N_20191,N_18003,N_18176);
nor U20192 (N_20192,N_16114,N_17115);
and U20193 (N_20193,N_17287,N_18316);
and U20194 (N_20194,N_16383,N_18318);
nor U20195 (N_20195,N_17834,N_16823);
xnor U20196 (N_20196,N_15735,N_17247);
nor U20197 (N_20197,N_15964,N_16068);
or U20198 (N_20198,N_17870,N_16100);
nand U20199 (N_20199,N_17071,N_15991);
and U20200 (N_20200,N_16052,N_15984);
nand U20201 (N_20201,N_16543,N_18428);
nand U20202 (N_20202,N_15955,N_17997);
nand U20203 (N_20203,N_17631,N_17544);
nand U20204 (N_20204,N_18687,N_17584);
nand U20205 (N_20205,N_16320,N_17781);
nor U20206 (N_20206,N_16587,N_17967);
and U20207 (N_20207,N_16205,N_18655);
or U20208 (N_20208,N_17964,N_15767);
xnor U20209 (N_20209,N_16767,N_16810);
and U20210 (N_20210,N_16728,N_17091);
or U20211 (N_20211,N_17288,N_16465);
nor U20212 (N_20212,N_16125,N_16449);
and U20213 (N_20213,N_15815,N_18563);
xor U20214 (N_20214,N_17124,N_15996);
and U20215 (N_20215,N_17937,N_17833);
nor U20216 (N_20216,N_16407,N_18732);
xnor U20217 (N_20217,N_15993,N_16074);
nor U20218 (N_20218,N_18572,N_17371);
nor U20219 (N_20219,N_18713,N_16044);
nand U20220 (N_20220,N_17509,N_17000);
or U20221 (N_20221,N_15701,N_16118);
nand U20222 (N_20222,N_17908,N_18211);
or U20223 (N_20223,N_16477,N_17901);
xor U20224 (N_20224,N_18072,N_17831);
and U20225 (N_20225,N_15774,N_16352);
and U20226 (N_20226,N_16676,N_18099);
xor U20227 (N_20227,N_17944,N_16995);
or U20228 (N_20228,N_17667,N_18638);
nor U20229 (N_20229,N_16265,N_15792);
nor U20230 (N_20230,N_18464,N_17186);
and U20231 (N_20231,N_16132,N_16302);
nand U20232 (N_20232,N_18653,N_16994);
xnor U20233 (N_20233,N_16195,N_18122);
or U20234 (N_20234,N_16004,N_16022);
and U20235 (N_20235,N_15924,N_18224);
or U20236 (N_20236,N_16439,N_16491);
or U20237 (N_20237,N_18476,N_16309);
nand U20238 (N_20238,N_16968,N_18596);
nand U20239 (N_20239,N_16359,N_17275);
and U20240 (N_20240,N_17066,N_17282);
nor U20241 (N_20241,N_16573,N_17620);
xor U20242 (N_20242,N_16045,N_16837);
and U20243 (N_20243,N_16315,N_15763);
and U20244 (N_20244,N_15770,N_15828);
xnor U20245 (N_20245,N_18562,N_18466);
or U20246 (N_20246,N_17248,N_17531);
nand U20247 (N_20247,N_18127,N_15810);
and U20248 (N_20248,N_16387,N_16075);
and U20249 (N_20249,N_18647,N_16486);
xnor U20250 (N_20250,N_15916,N_17516);
nor U20251 (N_20251,N_16960,N_16988);
and U20252 (N_20252,N_16571,N_15985);
or U20253 (N_20253,N_16103,N_17465);
nor U20254 (N_20254,N_18355,N_17438);
or U20255 (N_20255,N_18629,N_16495);
or U20256 (N_20256,N_16832,N_17869);
nor U20257 (N_20257,N_17337,N_16390);
nand U20258 (N_20258,N_17427,N_16849);
nor U20259 (N_20259,N_18615,N_16168);
or U20260 (N_20260,N_15758,N_16289);
nand U20261 (N_20261,N_18070,N_17092);
or U20262 (N_20262,N_16071,N_17050);
and U20263 (N_20263,N_16208,N_16855);
nor U20264 (N_20264,N_17732,N_18216);
and U20265 (N_20265,N_17225,N_17310);
nand U20266 (N_20266,N_16037,N_16415);
nor U20267 (N_20267,N_17618,N_17015);
xnor U20268 (N_20268,N_18478,N_18542);
nand U20269 (N_20269,N_16787,N_18167);
nand U20270 (N_20270,N_16099,N_17850);
nor U20271 (N_20271,N_17992,N_17362);
nand U20272 (N_20272,N_17654,N_17069);
and U20273 (N_20273,N_18313,N_16364);
nor U20274 (N_20274,N_16451,N_17701);
nor U20275 (N_20275,N_18285,N_17289);
nor U20276 (N_20276,N_15948,N_17270);
xnor U20277 (N_20277,N_17407,N_17772);
nand U20278 (N_20278,N_18535,N_18391);
nor U20279 (N_20279,N_16943,N_18155);
and U20280 (N_20280,N_17125,N_18083);
nor U20281 (N_20281,N_16140,N_16334);
nor U20282 (N_20282,N_18163,N_16777);
and U20283 (N_20283,N_15866,N_17246);
nor U20284 (N_20284,N_16690,N_18697);
and U20285 (N_20285,N_15632,N_17647);
nand U20286 (N_20286,N_18468,N_17914);
and U20287 (N_20287,N_17767,N_18349);
nor U20288 (N_20288,N_16939,N_16753);
or U20289 (N_20289,N_18644,N_17764);
and U20290 (N_20290,N_16827,N_15832);
and U20291 (N_20291,N_17662,N_18195);
nor U20292 (N_20292,N_16431,N_17839);
nor U20293 (N_20293,N_16136,N_17130);
or U20294 (N_20294,N_17197,N_17856);
or U20295 (N_20295,N_18436,N_17262);
or U20296 (N_20296,N_18721,N_17034);
xnor U20297 (N_20297,N_18712,N_18314);
or U20298 (N_20298,N_15829,N_18413);
or U20299 (N_20299,N_16611,N_18506);
and U20300 (N_20300,N_17390,N_15838);
nand U20301 (N_20301,N_18716,N_15744);
and U20302 (N_20302,N_16336,N_18345);
nor U20303 (N_20303,N_18399,N_17876);
and U20304 (N_20304,N_16840,N_17449);
or U20305 (N_20305,N_18559,N_16211);
or U20306 (N_20306,N_15994,N_15696);
and U20307 (N_20307,N_18415,N_16182);
nor U20308 (N_20308,N_15852,N_16926);
xor U20309 (N_20309,N_17290,N_15807);
nor U20310 (N_20310,N_16884,N_17936);
nor U20311 (N_20311,N_18145,N_16385);
or U20312 (N_20312,N_17610,N_16632);
nand U20313 (N_20313,N_17668,N_16473);
nand U20314 (N_20314,N_17121,N_17273);
and U20315 (N_20315,N_15721,N_16376);
nor U20316 (N_20316,N_16949,N_15652);
nand U20317 (N_20317,N_16740,N_17635);
and U20318 (N_20318,N_16948,N_16252);
nand U20319 (N_20319,N_18618,N_15712);
nand U20320 (N_20320,N_18700,N_17590);
nand U20321 (N_20321,N_17688,N_16004);
nor U20322 (N_20322,N_16460,N_17157);
and U20323 (N_20323,N_16501,N_15991);
nor U20324 (N_20324,N_17954,N_16897);
nand U20325 (N_20325,N_16632,N_15875);
and U20326 (N_20326,N_18235,N_17205);
and U20327 (N_20327,N_18444,N_17787);
nand U20328 (N_20328,N_16647,N_16915);
xor U20329 (N_20329,N_18429,N_17770);
xor U20330 (N_20330,N_17604,N_18656);
nand U20331 (N_20331,N_16984,N_17541);
and U20332 (N_20332,N_16421,N_17652);
or U20333 (N_20333,N_16368,N_16583);
and U20334 (N_20334,N_18192,N_16159);
and U20335 (N_20335,N_18741,N_18538);
nand U20336 (N_20336,N_16502,N_15927);
nor U20337 (N_20337,N_16285,N_16939);
or U20338 (N_20338,N_17193,N_16191);
and U20339 (N_20339,N_18295,N_15935);
nor U20340 (N_20340,N_18510,N_16412);
and U20341 (N_20341,N_16498,N_16426);
nand U20342 (N_20342,N_17918,N_18720);
and U20343 (N_20343,N_16594,N_18122);
xor U20344 (N_20344,N_18299,N_15725);
nand U20345 (N_20345,N_17272,N_17141);
and U20346 (N_20346,N_18556,N_16155);
nor U20347 (N_20347,N_16718,N_16035);
nand U20348 (N_20348,N_17885,N_16290);
xor U20349 (N_20349,N_16922,N_17776);
nand U20350 (N_20350,N_15801,N_17008);
nor U20351 (N_20351,N_15678,N_17841);
nand U20352 (N_20352,N_17600,N_16680);
or U20353 (N_20353,N_16847,N_17476);
nor U20354 (N_20354,N_18445,N_18437);
nand U20355 (N_20355,N_15778,N_15635);
or U20356 (N_20356,N_17878,N_17323);
nor U20357 (N_20357,N_18446,N_18694);
or U20358 (N_20358,N_16859,N_16001);
and U20359 (N_20359,N_18075,N_18329);
nand U20360 (N_20360,N_17896,N_16731);
xor U20361 (N_20361,N_15719,N_17746);
nand U20362 (N_20362,N_17174,N_17792);
nor U20363 (N_20363,N_17847,N_18399);
and U20364 (N_20364,N_17111,N_18158);
nor U20365 (N_20365,N_16962,N_18443);
and U20366 (N_20366,N_16836,N_17355);
nand U20367 (N_20367,N_17733,N_16719);
or U20368 (N_20368,N_18588,N_17990);
and U20369 (N_20369,N_15700,N_16265);
or U20370 (N_20370,N_18351,N_18057);
nand U20371 (N_20371,N_17487,N_17538);
or U20372 (N_20372,N_15727,N_17813);
or U20373 (N_20373,N_18631,N_16481);
xnor U20374 (N_20374,N_16226,N_17226);
or U20375 (N_20375,N_17809,N_16043);
nand U20376 (N_20376,N_18248,N_17001);
nor U20377 (N_20377,N_16887,N_16895);
and U20378 (N_20378,N_17942,N_17131);
nand U20379 (N_20379,N_17187,N_16979);
nand U20380 (N_20380,N_16678,N_17803);
and U20381 (N_20381,N_18205,N_15798);
nor U20382 (N_20382,N_17300,N_16941);
nand U20383 (N_20383,N_17635,N_16276);
or U20384 (N_20384,N_16784,N_18041);
and U20385 (N_20385,N_16842,N_17898);
nor U20386 (N_20386,N_15646,N_15881);
or U20387 (N_20387,N_18293,N_17261);
and U20388 (N_20388,N_18641,N_17640);
xnor U20389 (N_20389,N_17044,N_16358);
nand U20390 (N_20390,N_15762,N_18722);
and U20391 (N_20391,N_17406,N_18539);
nor U20392 (N_20392,N_15659,N_16995);
xnor U20393 (N_20393,N_15956,N_17928);
or U20394 (N_20394,N_17598,N_18747);
nand U20395 (N_20395,N_17274,N_17866);
nand U20396 (N_20396,N_17779,N_16940);
and U20397 (N_20397,N_18256,N_16462);
nor U20398 (N_20398,N_17166,N_16290);
and U20399 (N_20399,N_15922,N_15642);
nand U20400 (N_20400,N_17470,N_16588);
nand U20401 (N_20401,N_15650,N_17910);
nor U20402 (N_20402,N_15868,N_16944);
nor U20403 (N_20403,N_17363,N_17065);
xnor U20404 (N_20404,N_16706,N_16500);
or U20405 (N_20405,N_18231,N_15889);
xnor U20406 (N_20406,N_16458,N_16878);
or U20407 (N_20407,N_17689,N_18518);
xnor U20408 (N_20408,N_18332,N_15847);
or U20409 (N_20409,N_18438,N_15959);
nand U20410 (N_20410,N_18214,N_15844);
or U20411 (N_20411,N_18140,N_17139);
and U20412 (N_20412,N_17833,N_17259);
or U20413 (N_20413,N_18737,N_17071);
nor U20414 (N_20414,N_18264,N_17019);
or U20415 (N_20415,N_17468,N_18038);
or U20416 (N_20416,N_16642,N_17436);
nor U20417 (N_20417,N_18442,N_17893);
nor U20418 (N_20418,N_15797,N_17977);
nand U20419 (N_20419,N_16007,N_16767);
nand U20420 (N_20420,N_17041,N_16793);
or U20421 (N_20421,N_18579,N_15910);
nand U20422 (N_20422,N_18498,N_18467);
nor U20423 (N_20423,N_16787,N_17955);
and U20424 (N_20424,N_17420,N_15929);
xnor U20425 (N_20425,N_17911,N_17682);
and U20426 (N_20426,N_16282,N_18172);
nor U20427 (N_20427,N_16338,N_15794);
and U20428 (N_20428,N_16266,N_18739);
nand U20429 (N_20429,N_16350,N_17274);
nor U20430 (N_20430,N_16457,N_16245);
or U20431 (N_20431,N_17664,N_18336);
or U20432 (N_20432,N_17643,N_18155);
nor U20433 (N_20433,N_17001,N_17081);
nand U20434 (N_20434,N_18302,N_15780);
nand U20435 (N_20435,N_16076,N_17995);
nor U20436 (N_20436,N_16704,N_18062);
nand U20437 (N_20437,N_16938,N_16172);
xor U20438 (N_20438,N_18678,N_17723);
nor U20439 (N_20439,N_15771,N_17572);
or U20440 (N_20440,N_16344,N_17149);
nor U20441 (N_20441,N_16073,N_17502);
and U20442 (N_20442,N_16903,N_16179);
nand U20443 (N_20443,N_16033,N_16637);
and U20444 (N_20444,N_18713,N_18561);
nor U20445 (N_20445,N_17758,N_17246);
or U20446 (N_20446,N_16637,N_17452);
nor U20447 (N_20447,N_16944,N_16344);
nor U20448 (N_20448,N_16589,N_17680);
nand U20449 (N_20449,N_15690,N_18188);
or U20450 (N_20450,N_17726,N_18254);
and U20451 (N_20451,N_18648,N_16618);
nand U20452 (N_20452,N_17904,N_16242);
xnor U20453 (N_20453,N_17651,N_17104);
and U20454 (N_20454,N_18372,N_16824);
and U20455 (N_20455,N_18083,N_18212);
nand U20456 (N_20456,N_17293,N_16941);
nand U20457 (N_20457,N_17699,N_15902);
nor U20458 (N_20458,N_18695,N_15926);
nor U20459 (N_20459,N_17441,N_17115);
xor U20460 (N_20460,N_17110,N_17468);
nor U20461 (N_20461,N_16481,N_16347);
nand U20462 (N_20462,N_17447,N_16554);
nor U20463 (N_20463,N_16814,N_18609);
nand U20464 (N_20464,N_16558,N_16631);
nand U20465 (N_20465,N_17782,N_16684);
nor U20466 (N_20466,N_15976,N_17334);
nand U20467 (N_20467,N_16110,N_17393);
xnor U20468 (N_20468,N_18719,N_18005);
or U20469 (N_20469,N_18575,N_18352);
nor U20470 (N_20470,N_18713,N_18462);
nand U20471 (N_20471,N_16539,N_18418);
xor U20472 (N_20472,N_16114,N_16429);
nand U20473 (N_20473,N_17322,N_15672);
nor U20474 (N_20474,N_17690,N_15912);
nor U20475 (N_20475,N_16297,N_18490);
nand U20476 (N_20476,N_17035,N_18226);
and U20477 (N_20477,N_17689,N_18408);
or U20478 (N_20478,N_17212,N_17551);
nor U20479 (N_20479,N_15725,N_16257);
xnor U20480 (N_20480,N_17822,N_18693);
nand U20481 (N_20481,N_16481,N_16592);
and U20482 (N_20482,N_15852,N_17741);
nand U20483 (N_20483,N_18072,N_16093);
or U20484 (N_20484,N_15686,N_16310);
and U20485 (N_20485,N_15921,N_17886);
nand U20486 (N_20486,N_16152,N_18617);
or U20487 (N_20487,N_17227,N_17748);
and U20488 (N_20488,N_16425,N_17388);
nor U20489 (N_20489,N_18456,N_18241);
xnor U20490 (N_20490,N_16285,N_17966);
and U20491 (N_20491,N_16394,N_17511);
and U20492 (N_20492,N_17089,N_16601);
and U20493 (N_20493,N_16668,N_18170);
nand U20494 (N_20494,N_16627,N_17887);
nor U20495 (N_20495,N_18070,N_16037);
or U20496 (N_20496,N_18741,N_15982);
nand U20497 (N_20497,N_18120,N_16834);
and U20498 (N_20498,N_18635,N_18263);
nor U20499 (N_20499,N_16632,N_16825);
xor U20500 (N_20500,N_17823,N_16427);
nor U20501 (N_20501,N_18480,N_17814);
xnor U20502 (N_20502,N_15790,N_15797);
nand U20503 (N_20503,N_15963,N_16178);
nor U20504 (N_20504,N_16850,N_17992);
nand U20505 (N_20505,N_15807,N_17838);
xor U20506 (N_20506,N_17109,N_17836);
nor U20507 (N_20507,N_16351,N_18177);
nor U20508 (N_20508,N_15648,N_16519);
nand U20509 (N_20509,N_17501,N_17171);
nand U20510 (N_20510,N_16870,N_17057);
or U20511 (N_20511,N_16699,N_16405);
nor U20512 (N_20512,N_17376,N_18335);
xnor U20513 (N_20513,N_17469,N_16341);
or U20514 (N_20514,N_18174,N_17844);
or U20515 (N_20515,N_15829,N_16393);
nor U20516 (N_20516,N_18319,N_15973);
nand U20517 (N_20517,N_15865,N_15999);
and U20518 (N_20518,N_18183,N_16053);
and U20519 (N_20519,N_17290,N_16991);
and U20520 (N_20520,N_17802,N_18664);
xnor U20521 (N_20521,N_16121,N_18403);
xor U20522 (N_20522,N_17945,N_18191);
nand U20523 (N_20523,N_16696,N_16311);
or U20524 (N_20524,N_18612,N_18575);
nand U20525 (N_20525,N_17410,N_16942);
or U20526 (N_20526,N_18083,N_17697);
nand U20527 (N_20527,N_18402,N_17532);
xor U20528 (N_20528,N_18112,N_17446);
and U20529 (N_20529,N_16607,N_17363);
nor U20530 (N_20530,N_17752,N_18686);
or U20531 (N_20531,N_15998,N_16819);
and U20532 (N_20532,N_17289,N_16697);
nand U20533 (N_20533,N_18018,N_16587);
or U20534 (N_20534,N_17771,N_18417);
or U20535 (N_20535,N_16015,N_18330);
nand U20536 (N_20536,N_17392,N_16869);
xor U20537 (N_20537,N_16092,N_17744);
nand U20538 (N_20538,N_17736,N_15961);
and U20539 (N_20539,N_16880,N_16310);
or U20540 (N_20540,N_17637,N_17516);
and U20541 (N_20541,N_16807,N_17152);
xor U20542 (N_20542,N_18265,N_18323);
nand U20543 (N_20543,N_15695,N_17786);
nor U20544 (N_20544,N_17106,N_16236);
nand U20545 (N_20545,N_16853,N_18147);
or U20546 (N_20546,N_15647,N_16199);
and U20547 (N_20547,N_18394,N_16785);
nand U20548 (N_20548,N_17560,N_16376);
nand U20549 (N_20549,N_16215,N_16903);
nor U20550 (N_20550,N_16129,N_16968);
nor U20551 (N_20551,N_17325,N_17259);
nand U20552 (N_20552,N_17038,N_15797);
or U20553 (N_20553,N_17156,N_17708);
nand U20554 (N_20554,N_16890,N_17906);
or U20555 (N_20555,N_17613,N_15940);
nor U20556 (N_20556,N_17251,N_16941);
and U20557 (N_20557,N_18029,N_16722);
and U20558 (N_20558,N_17042,N_17311);
nor U20559 (N_20559,N_16766,N_16842);
and U20560 (N_20560,N_17266,N_16416);
nand U20561 (N_20561,N_16560,N_16874);
and U20562 (N_20562,N_15701,N_17852);
nand U20563 (N_20563,N_16341,N_16508);
and U20564 (N_20564,N_16788,N_17020);
nor U20565 (N_20565,N_17818,N_17743);
nand U20566 (N_20566,N_16027,N_18719);
nand U20567 (N_20567,N_16560,N_15764);
or U20568 (N_20568,N_16858,N_16309);
nor U20569 (N_20569,N_17290,N_17410);
and U20570 (N_20570,N_17733,N_18117);
or U20571 (N_20571,N_17429,N_16858);
or U20572 (N_20572,N_17254,N_18578);
xnor U20573 (N_20573,N_15815,N_17933);
nor U20574 (N_20574,N_17965,N_17330);
or U20575 (N_20575,N_16264,N_15850);
or U20576 (N_20576,N_15787,N_17779);
nor U20577 (N_20577,N_18376,N_16191);
and U20578 (N_20578,N_18066,N_18718);
and U20579 (N_20579,N_18330,N_17658);
and U20580 (N_20580,N_15953,N_17814);
nand U20581 (N_20581,N_16873,N_16742);
nor U20582 (N_20582,N_17680,N_17684);
and U20583 (N_20583,N_18247,N_17225);
and U20584 (N_20584,N_17054,N_17155);
or U20585 (N_20585,N_17212,N_18071);
or U20586 (N_20586,N_18379,N_17152);
xnor U20587 (N_20587,N_18234,N_17019);
xnor U20588 (N_20588,N_18095,N_15669);
xor U20589 (N_20589,N_18151,N_16748);
nand U20590 (N_20590,N_18419,N_15947);
and U20591 (N_20591,N_17211,N_17310);
or U20592 (N_20592,N_16633,N_17069);
nand U20593 (N_20593,N_17582,N_18574);
nor U20594 (N_20594,N_18113,N_18748);
nand U20595 (N_20595,N_17274,N_18069);
nor U20596 (N_20596,N_17755,N_18235);
nand U20597 (N_20597,N_17481,N_16207);
nor U20598 (N_20598,N_15644,N_17015);
or U20599 (N_20599,N_18546,N_18172);
nor U20600 (N_20600,N_18109,N_17649);
nor U20601 (N_20601,N_15852,N_17059);
and U20602 (N_20602,N_15728,N_15943);
nor U20603 (N_20603,N_18728,N_15837);
nor U20604 (N_20604,N_15846,N_17338);
or U20605 (N_20605,N_17794,N_17795);
xor U20606 (N_20606,N_18100,N_16435);
or U20607 (N_20607,N_18378,N_16559);
or U20608 (N_20608,N_18268,N_18319);
nor U20609 (N_20609,N_16435,N_16244);
or U20610 (N_20610,N_16868,N_17044);
and U20611 (N_20611,N_18004,N_17456);
nor U20612 (N_20612,N_17224,N_15899);
nor U20613 (N_20613,N_15871,N_17702);
nor U20614 (N_20614,N_18047,N_16739);
nor U20615 (N_20615,N_17152,N_17623);
nor U20616 (N_20616,N_17155,N_16181);
and U20617 (N_20617,N_16282,N_18694);
nand U20618 (N_20618,N_17396,N_18553);
nor U20619 (N_20619,N_16884,N_16995);
nand U20620 (N_20620,N_18335,N_18692);
and U20621 (N_20621,N_15924,N_17282);
and U20622 (N_20622,N_18519,N_17585);
xor U20623 (N_20623,N_16462,N_18561);
nand U20624 (N_20624,N_15959,N_18004);
and U20625 (N_20625,N_18491,N_15626);
or U20626 (N_20626,N_17786,N_16241);
nand U20627 (N_20627,N_17627,N_16880);
or U20628 (N_20628,N_18715,N_18237);
and U20629 (N_20629,N_17619,N_17764);
nor U20630 (N_20630,N_15803,N_17532);
or U20631 (N_20631,N_18050,N_16710);
nand U20632 (N_20632,N_17788,N_15938);
nor U20633 (N_20633,N_17641,N_18737);
and U20634 (N_20634,N_17179,N_16596);
nand U20635 (N_20635,N_16333,N_17010);
or U20636 (N_20636,N_17021,N_16870);
or U20637 (N_20637,N_18298,N_16555);
or U20638 (N_20638,N_16813,N_17770);
and U20639 (N_20639,N_16440,N_18508);
or U20640 (N_20640,N_16391,N_17884);
and U20641 (N_20641,N_17389,N_16284);
nand U20642 (N_20642,N_17774,N_18657);
and U20643 (N_20643,N_17842,N_17466);
or U20644 (N_20644,N_17317,N_15853);
nand U20645 (N_20645,N_16758,N_17025);
or U20646 (N_20646,N_18027,N_18507);
nor U20647 (N_20647,N_18538,N_18216);
or U20648 (N_20648,N_16671,N_16290);
nand U20649 (N_20649,N_17248,N_15659);
nor U20650 (N_20650,N_16270,N_18534);
nor U20651 (N_20651,N_17416,N_17254);
and U20652 (N_20652,N_16142,N_16507);
nand U20653 (N_20653,N_18359,N_18071);
nor U20654 (N_20654,N_16253,N_16255);
and U20655 (N_20655,N_16614,N_16219);
nor U20656 (N_20656,N_18168,N_18674);
and U20657 (N_20657,N_16516,N_16160);
and U20658 (N_20658,N_15773,N_17130);
or U20659 (N_20659,N_18063,N_18699);
or U20660 (N_20660,N_17119,N_18348);
xor U20661 (N_20661,N_16664,N_17525);
nand U20662 (N_20662,N_18544,N_16709);
nand U20663 (N_20663,N_16445,N_17760);
nor U20664 (N_20664,N_17770,N_17473);
and U20665 (N_20665,N_17904,N_16579);
nor U20666 (N_20666,N_16339,N_18392);
and U20667 (N_20667,N_17544,N_16634);
nor U20668 (N_20668,N_16174,N_16466);
nor U20669 (N_20669,N_17950,N_15675);
or U20670 (N_20670,N_15803,N_18490);
and U20671 (N_20671,N_17051,N_16302);
nand U20672 (N_20672,N_18188,N_17402);
or U20673 (N_20673,N_16768,N_15786);
and U20674 (N_20674,N_17295,N_16789);
nand U20675 (N_20675,N_15865,N_15868);
nor U20676 (N_20676,N_17482,N_18058);
nand U20677 (N_20677,N_18394,N_17081);
nand U20678 (N_20678,N_16831,N_18008);
and U20679 (N_20679,N_15948,N_18438);
or U20680 (N_20680,N_16128,N_17602);
nand U20681 (N_20681,N_17702,N_15921);
and U20682 (N_20682,N_17865,N_17366);
nor U20683 (N_20683,N_18603,N_16173);
or U20684 (N_20684,N_16148,N_18314);
and U20685 (N_20685,N_17514,N_18747);
nor U20686 (N_20686,N_15896,N_18054);
xnor U20687 (N_20687,N_15673,N_17209);
or U20688 (N_20688,N_18710,N_16783);
xor U20689 (N_20689,N_16549,N_17725);
and U20690 (N_20690,N_17107,N_16712);
nor U20691 (N_20691,N_15819,N_16781);
nand U20692 (N_20692,N_17809,N_17909);
nand U20693 (N_20693,N_18584,N_16344);
and U20694 (N_20694,N_17579,N_16615);
or U20695 (N_20695,N_15677,N_18282);
nor U20696 (N_20696,N_16406,N_15986);
nor U20697 (N_20697,N_17588,N_17947);
xnor U20698 (N_20698,N_17909,N_18615);
nand U20699 (N_20699,N_16175,N_16931);
nand U20700 (N_20700,N_16500,N_17284);
nand U20701 (N_20701,N_16314,N_16949);
nor U20702 (N_20702,N_17399,N_18603);
and U20703 (N_20703,N_16707,N_17467);
or U20704 (N_20704,N_17873,N_18309);
and U20705 (N_20705,N_17326,N_17805);
nor U20706 (N_20706,N_16601,N_17818);
nand U20707 (N_20707,N_16551,N_17815);
nand U20708 (N_20708,N_16926,N_16142);
nor U20709 (N_20709,N_15746,N_16805);
and U20710 (N_20710,N_18499,N_17583);
nand U20711 (N_20711,N_16512,N_16490);
nand U20712 (N_20712,N_17585,N_18200);
nor U20713 (N_20713,N_17115,N_16135);
nand U20714 (N_20714,N_16118,N_16390);
nor U20715 (N_20715,N_17738,N_18433);
or U20716 (N_20716,N_16269,N_17023);
or U20717 (N_20717,N_16305,N_18652);
nand U20718 (N_20718,N_15950,N_16090);
nand U20719 (N_20719,N_15799,N_18374);
nor U20720 (N_20720,N_17497,N_15991);
and U20721 (N_20721,N_16801,N_18245);
nand U20722 (N_20722,N_18395,N_16005);
and U20723 (N_20723,N_16810,N_17876);
and U20724 (N_20724,N_18328,N_16532);
nand U20725 (N_20725,N_18408,N_18358);
nor U20726 (N_20726,N_16171,N_16656);
or U20727 (N_20727,N_17518,N_17045);
nand U20728 (N_20728,N_18094,N_16417);
nand U20729 (N_20729,N_17978,N_18442);
nor U20730 (N_20730,N_17998,N_17658);
nand U20731 (N_20731,N_16249,N_16040);
nand U20732 (N_20732,N_15869,N_17935);
and U20733 (N_20733,N_16477,N_16472);
and U20734 (N_20734,N_16179,N_18299);
nand U20735 (N_20735,N_17527,N_17930);
or U20736 (N_20736,N_17632,N_17459);
and U20737 (N_20737,N_16330,N_17498);
and U20738 (N_20738,N_16659,N_15973);
and U20739 (N_20739,N_18251,N_17031);
and U20740 (N_20740,N_18081,N_17793);
and U20741 (N_20741,N_18016,N_16995);
nand U20742 (N_20742,N_16902,N_18654);
nand U20743 (N_20743,N_17288,N_16143);
nor U20744 (N_20744,N_17466,N_16109);
nor U20745 (N_20745,N_16028,N_18278);
nand U20746 (N_20746,N_17571,N_15727);
or U20747 (N_20747,N_16675,N_17353);
nand U20748 (N_20748,N_18356,N_17250);
and U20749 (N_20749,N_17810,N_17168);
xor U20750 (N_20750,N_18250,N_17945);
or U20751 (N_20751,N_17986,N_17061);
or U20752 (N_20752,N_17896,N_16920);
nor U20753 (N_20753,N_17253,N_18718);
or U20754 (N_20754,N_18715,N_15786);
nand U20755 (N_20755,N_17024,N_18587);
nor U20756 (N_20756,N_15718,N_16889);
and U20757 (N_20757,N_16180,N_18134);
or U20758 (N_20758,N_17688,N_18483);
nor U20759 (N_20759,N_17431,N_16905);
nor U20760 (N_20760,N_17425,N_17995);
and U20761 (N_20761,N_17539,N_15861);
nand U20762 (N_20762,N_17643,N_17257);
nand U20763 (N_20763,N_17699,N_15894);
nor U20764 (N_20764,N_18036,N_16476);
or U20765 (N_20765,N_17931,N_17758);
or U20766 (N_20766,N_17645,N_16671);
nor U20767 (N_20767,N_17804,N_16074);
or U20768 (N_20768,N_18401,N_18368);
or U20769 (N_20769,N_18590,N_16383);
xnor U20770 (N_20770,N_17325,N_16188);
nor U20771 (N_20771,N_17342,N_18077);
xnor U20772 (N_20772,N_18084,N_17479);
nand U20773 (N_20773,N_16735,N_18381);
nand U20774 (N_20774,N_15901,N_16042);
or U20775 (N_20775,N_17704,N_16792);
nand U20776 (N_20776,N_16418,N_16909);
or U20777 (N_20777,N_16942,N_17508);
and U20778 (N_20778,N_15872,N_15858);
nor U20779 (N_20779,N_15631,N_18080);
xnor U20780 (N_20780,N_16124,N_18093);
and U20781 (N_20781,N_17099,N_16927);
nor U20782 (N_20782,N_16986,N_17230);
or U20783 (N_20783,N_17407,N_17361);
nor U20784 (N_20784,N_17212,N_16051);
xor U20785 (N_20785,N_16716,N_16958);
or U20786 (N_20786,N_17050,N_16672);
and U20787 (N_20787,N_15790,N_18608);
or U20788 (N_20788,N_16475,N_15918);
nand U20789 (N_20789,N_17977,N_15897);
nor U20790 (N_20790,N_17572,N_18539);
or U20791 (N_20791,N_17386,N_17406);
nor U20792 (N_20792,N_16046,N_17899);
nor U20793 (N_20793,N_17103,N_18054);
or U20794 (N_20794,N_16061,N_17248);
and U20795 (N_20795,N_16691,N_17447);
or U20796 (N_20796,N_15821,N_16902);
and U20797 (N_20797,N_18732,N_16627);
nor U20798 (N_20798,N_18285,N_16047);
and U20799 (N_20799,N_16877,N_17651);
nor U20800 (N_20800,N_17056,N_18679);
xnor U20801 (N_20801,N_17099,N_17094);
nor U20802 (N_20802,N_18117,N_16942);
or U20803 (N_20803,N_18526,N_18453);
xnor U20804 (N_20804,N_16385,N_17353);
nor U20805 (N_20805,N_17712,N_18521);
or U20806 (N_20806,N_17024,N_16724);
or U20807 (N_20807,N_16227,N_18666);
and U20808 (N_20808,N_17504,N_17640);
nor U20809 (N_20809,N_16374,N_17006);
nor U20810 (N_20810,N_15627,N_17543);
nand U20811 (N_20811,N_17994,N_17920);
and U20812 (N_20812,N_16520,N_18665);
xor U20813 (N_20813,N_17158,N_16684);
and U20814 (N_20814,N_16915,N_16155);
nor U20815 (N_20815,N_16650,N_17990);
xor U20816 (N_20816,N_18086,N_16965);
xnor U20817 (N_20817,N_16094,N_16740);
or U20818 (N_20818,N_15693,N_18063);
or U20819 (N_20819,N_17073,N_15684);
nor U20820 (N_20820,N_18407,N_15864);
nor U20821 (N_20821,N_16256,N_16286);
xnor U20822 (N_20822,N_17924,N_16873);
and U20823 (N_20823,N_17262,N_16609);
or U20824 (N_20824,N_17624,N_17324);
and U20825 (N_20825,N_15674,N_16400);
nor U20826 (N_20826,N_17355,N_17426);
xor U20827 (N_20827,N_17890,N_16078);
or U20828 (N_20828,N_16268,N_15715);
or U20829 (N_20829,N_17679,N_17945);
and U20830 (N_20830,N_17433,N_16905);
or U20831 (N_20831,N_16831,N_17788);
nor U20832 (N_20832,N_18331,N_16294);
xnor U20833 (N_20833,N_17874,N_18181);
or U20834 (N_20834,N_18056,N_16163);
and U20835 (N_20835,N_16189,N_18420);
nand U20836 (N_20836,N_18299,N_16371);
and U20837 (N_20837,N_16871,N_15696);
or U20838 (N_20838,N_15983,N_16638);
and U20839 (N_20839,N_15687,N_18143);
and U20840 (N_20840,N_17616,N_16496);
nor U20841 (N_20841,N_15860,N_16225);
nand U20842 (N_20842,N_17706,N_15645);
or U20843 (N_20843,N_18148,N_18265);
nor U20844 (N_20844,N_18724,N_18217);
and U20845 (N_20845,N_18532,N_18684);
or U20846 (N_20846,N_18265,N_16881);
and U20847 (N_20847,N_16231,N_18504);
nor U20848 (N_20848,N_15875,N_16133);
nor U20849 (N_20849,N_18551,N_16547);
xnor U20850 (N_20850,N_17258,N_17637);
xnor U20851 (N_20851,N_16414,N_17875);
nand U20852 (N_20852,N_16884,N_17618);
or U20853 (N_20853,N_18357,N_18368);
nand U20854 (N_20854,N_16257,N_16752);
nand U20855 (N_20855,N_15960,N_18733);
or U20856 (N_20856,N_16501,N_18356);
nor U20857 (N_20857,N_18313,N_15909);
nor U20858 (N_20858,N_16043,N_15906);
nand U20859 (N_20859,N_16918,N_18585);
or U20860 (N_20860,N_15806,N_16578);
nor U20861 (N_20861,N_17624,N_15767);
nand U20862 (N_20862,N_17021,N_16235);
nor U20863 (N_20863,N_18449,N_15815);
nand U20864 (N_20864,N_17322,N_16983);
nor U20865 (N_20865,N_18400,N_15744);
and U20866 (N_20866,N_16300,N_17245);
nor U20867 (N_20867,N_18310,N_18341);
and U20868 (N_20868,N_18287,N_16267);
nor U20869 (N_20869,N_15732,N_16360);
nand U20870 (N_20870,N_18159,N_17020);
nand U20871 (N_20871,N_18276,N_15971);
or U20872 (N_20872,N_16882,N_17032);
nand U20873 (N_20873,N_16803,N_17974);
nor U20874 (N_20874,N_17174,N_16909);
nor U20875 (N_20875,N_16721,N_16539);
nor U20876 (N_20876,N_18594,N_17858);
xor U20877 (N_20877,N_17073,N_17038);
nand U20878 (N_20878,N_15874,N_16937);
nand U20879 (N_20879,N_17752,N_16675);
or U20880 (N_20880,N_17192,N_17627);
nand U20881 (N_20881,N_17521,N_17222);
or U20882 (N_20882,N_18139,N_17597);
and U20883 (N_20883,N_16993,N_18374);
nand U20884 (N_20884,N_16086,N_17340);
xor U20885 (N_20885,N_17733,N_16947);
and U20886 (N_20886,N_15752,N_17618);
and U20887 (N_20887,N_16764,N_16442);
or U20888 (N_20888,N_16030,N_16546);
or U20889 (N_20889,N_17880,N_15860);
and U20890 (N_20890,N_18112,N_15807);
nor U20891 (N_20891,N_17966,N_17894);
nor U20892 (N_20892,N_17904,N_16481);
or U20893 (N_20893,N_16854,N_17603);
xnor U20894 (N_20894,N_17421,N_17410);
or U20895 (N_20895,N_18515,N_17691);
nor U20896 (N_20896,N_16878,N_17482);
xor U20897 (N_20897,N_17110,N_17994);
nand U20898 (N_20898,N_18053,N_18322);
or U20899 (N_20899,N_16243,N_17667);
and U20900 (N_20900,N_17500,N_15859);
xor U20901 (N_20901,N_15743,N_18385);
and U20902 (N_20902,N_17576,N_15637);
nor U20903 (N_20903,N_16903,N_18128);
nor U20904 (N_20904,N_17840,N_16849);
and U20905 (N_20905,N_16671,N_18318);
and U20906 (N_20906,N_16685,N_16003);
nand U20907 (N_20907,N_17575,N_18023);
nand U20908 (N_20908,N_17946,N_15673);
nor U20909 (N_20909,N_15633,N_18590);
nor U20910 (N_20910,N_16995,N_17808);
and U20911 (N_20911,N_15633,N_18698);
and U20912 (N_20912,N_15787,N_17758);
nand U20913 (N_20913,N_18568,N_16367);
nand U20914 (N_20914,N_16869,N_17968);
nand U20915 (N_20915,N_16382,N_18288);
or U20916 (N_20916,N_17090,N_17403);
xor U20917 (N_20917,N_17719,N_18446);
or U20918 (N_20918,N_18436,N_15662);
nand U20919 (N_20919,N_16853,N_17426);
or U20920 (N_20920,N_17005,N_18726);
and U20921 (N_20921,N_17897,N_17061);
nor U20922 (N_20922,N_16760,N_16333);
nor U20923 (N_20923,N_16757,N_17490);
nand U20924 (N_20924,N_16069,N_17948);
or U20925 (N_20925,N_18308,N_16254);
nand U20926 (N_20926,N_16794,N_17164);
or U20927 (N_20927,N_16279,N_17456);
nor U20928 (N_20928,N_17992,N_17001);
and U20929 (N_20929,N_17837,N_16284);
nand U20930 (N_20930,N_15655,N_15738);
and U20931 (N_20931,N_18454,N_18159);
nand U20932 (N_20932,N_16364,N_17258);
and U20933 (N_20933,N_17442,N_16864);
and U20934 (N_20934,N_17931,N_17939);
and U20935 (N_20935,N_15848,N_18192);
nand U20936 (N_20936,N_16891,N_16508);
or U20937 (N_20937,N_18289,N_15648);
and U20938 (N_20938,N_16982,N_18337);
or U20939 (N_20939,N_18574,N_16434);
nand U20940 (N_20940,N_16024,N_18446);
nand U20941 (N_20941,N_18350,N_16113);
nand U20942 (N_20942,N_16959,N_18227);
nand U20943 (N_20943,N_18344,N_17580);
or U20944 (N_20944,N_17881,N_15749);
and U20945 (N_20945,N_18378,N_18691);
nand U20946 (N_20946,N_16138,N_16985);
xnor U20947 (N_20947,N_16375,N_15736);
or U20948 (N_20948,N_16838,N_17600);
nand U20949 (N_20949,N_15829,N_17265);
and U20950 (N_20950,N_16396,N_16982);
or U20951 (N_20951,N_16778,N_18194);
or U20952 (N_20952,N_16479,N_15667);
nor U20953 (N_20953,N_15628,N_17547);
or U20954 (N_20954,N_17083,N_16026);
and U20955 (N_20955,N_17914,N_18523);
nand U20956 (N_20956,N_18016,N_17108);
xor U20957 (N_20957,N_17739,N_16302);
or U20958 (N_20958,N_18563,N_18713);
and U20959 (N_20959,N_16400,N_16944);
and U20960 (N_20960,N_15761,N_16971);
nor U20961 (N_20961,N_15949,N_18522);
nor U20962 (N_20962,N_16430,N_16683);
nor U20963 (N_20963,N_15660,N_16053);
nand U20964 (N_20964,N_18169,N_17103);
nor U20965 (N_20965,N_16855,N_16867);
and U20966 (N_20966,N_18648,N_18527);
or U20967 (N_20967,N_16934,N_18485);
nor U20968 (N_20968,N_16064,N_16727);
and U20969 (N_20969,N_18082,N_18145);
nor U20970 (N_20970,N_17461,N_17846);
xor U20971 (N_20971,N_18565,N_17882);
nand U20972 (N_20972,N_17678,N_16696);
or U20973 (N_20973,N_17286,N_15685);
or U20974 (N_20974,N_15827,N_18227);
nand U20975 (N_20975,N_16649,N_16801);
nor U20976 (N_20976,N_17640,N_16397);
or U20977 (N_20977,N_16920,N_15664);
and U20978 (N_20978,N_18043,N_17226);
and U20979 (N_20979,N_16277,N_17291);
or U20980 (N_20980,N_17281,N_17267);
nand U20981 (N_20981,N_18202,N_15899);
and U20982 (N_20982,N_16319,N_16961);
and U20983 (N_20983,N_16036,N_17533);
or U20984 (N_20984,N_16435,N_17000);
nor U20985 (N_20985,N_16544,N_17975);
nor U20986 (N_20986,N_16385,N_16316);
and U20987 (N_20987,N_17724,N_16633);
xor U20988 (N_20988,N_17235,N_18722);
xor U20989 (N_20989,N_17317,N_16292);
or U20990 (N_20990,N_16508,N_15675);
and U20991 (N_20991,N_18135,N_18021);
or U20992 (N_20992,N_17014,N_18268);
nand U20993 (N_20993,N_16612,N_17000);
nor U20994 (N_20994,N_17325,N_18657);
xor U20995 (N_20995,N_18069,N_17712);
nand U20996 (N_20996,N_16559,N_16418);
nor U20997 (N_20997,N_18103,N_18247);
nor U20998 (N_20998,N_17967,N_18698);
nor U20999 (N_20999,N_17442,N_17621);
nand U21000 (N_21000,N_16487,N_18236);
and U21001 (N_21001,N_18034,N_18146);
nand U21002 (N_21002,N_16929,N_18650);
and U21003 (N_21003,N_17736,N_16098);
nand U21004 (N_21004,N_16641,N_17199);
or U21005 (N_21005,N_17900,N_17233);
or U21006 (N_21006,N_17593,N_16786);
nor U21007 (N_21007,N_16357,N_16428);
nor U21008 (N_21008,N_15829,N_17200);
or U21009 (N_21009,N_18083,N_16997);
xnor U21010 (N_21010,N_18051,N_18061);
nor U21011 (N_21011,N_17746,N_17100);
or U21012 (N_21012,N_17092,N_17409);
nor U21013 (N_21013,N_17720,N_16729);
or U21014 (N_21014,N_16889,N_17041);
nand U21015 (N_21015,N_18228,N_18561);
and U21016 (N_21016,N_16891,N_16935);
or U21017 (N_21017,N_16830,N_16735);
and U21018 (N_21018,N_16139,N_17678);
xnor U21019 (N_21019,N_17590,N_18643);
nand U21020 (N_21020,N_18532,N_16307);
nor U21021 (N_21021,N_18090,N_16308);
nor U21022 (N_21022,N_18194,N_18294);
and U21023 (N_21023,N_18577,N_16871);
and U21024 (N_21024,N_18284,N_18710);
nand U21025 (N_21025,N_18519,N_16496);
or U21026 (N_21026,N_16687,N_15811);
nor U21027 (N_21027,N_18030,N_17749);
xor U21028 (N_21028,N_16978,N_18528);
and U21029 (N_21029,N_16048,N_15895);
and U21030 (N_21030,N_17285,N_15813);
or U21031 (N_21031,N_16240,N_16237);
nand U21032 (N_21032,N_17335,N_17707);
nand U21033 (N_21033,N_16474,N_17763);
and U21034 (N_21034,N_16358,N_17707);
nand U21035 (N_21035,N_17572,N_15975);
or U21036 (N_21036,N_17308,N_18456);
and U21037 (N_21037,N_17074,N_15935);
nor U21038 (N_21038,N_18683,N_18694);
or U21039 (N_21039,N_17279,N_18366);
nand U21040 (N_21040,N_18191,N_15788);
nor U21041 (N_21041,N_15886,N_17944);
or U21042 (N_21042,N_16206,N_18575);
and U21043 (N_21043,N_17456,N_15854);
or U21044 (N_21044,N_16315,N_16647);
xnor U21045 (N_21045,N_17516,N_17737);
nand U21046 (N_21046,N_16238,N_16397);
and U21047 (N_21047,N_15692,N_18533);
nand U21048 (N_21048,N_17671,N_18623);
xnor U21049 (N_21049,N_16894,N_17793);
nand U21050 (N_21050,N_15937,N_17399);
nand U21051 (N_21051,N_15832,N_18302);
and U21052 (N_21052,N_15974,N_17445);
nor U21053 (N_21053,N_18493,N_15841);
nor U21054 (N_21054,N_15807,N_17951);
or U21055 (N_21055,N_18176,N_16772);
or U21056 (N_21056,N_18314,N_17446);
nor U21057 (N_21057,N_16034,N_17153);
xnor U21058 (N_21058,N_17583,N_18691);
and U21059 (N_21059,N_18717,N_17196);
and U21060 (N_21060,N_17894,N_17651);
and U21061 (N_21061,N_16343,N_17896);
nor U21062 (N_21062,N_15922,N_16576);
and U21063 (N_21063,N_17556,N_16356);
xnor U21064 (N_21064,N_18009,N_18571);
nor U21065 (N_21065,N_17595,N_15838);
nor U21066 (N_21066,N_15764,N_17405);
and U21067 (N_21067,N_16751,N_18668);
nor U21068 (N_21068,N_17799,N_16691);
and U21069 (N_21069,N_18472,N_17695);
nand U21070 (N_21070,N_15709,N_17502);
and U21071 (N_21071,N_17537,N_18683);
nand U21072 (N_21072,N_16302,N_18195);
xor U21073 (N_21073,N_18120,N_16587);
or U21074 (N_21074,N_15954,N_16515);
or U21075 (N_21075,N_17115,N_16023);
and U21076 (N_21076,N_18281,N_18286);
and U21077 (N_21077,N_17027,N_18462);
or U21078 (N_21078,N_18068,N_17714);
xor U21079 (N_21079,N_17183,N_17828);
nor U21080 (N_21080,N_17569,N_15687);
and U21081 (N_21081,N_17527,N_18288);
nor U21082 (N_21082,N_15640,N_17752);
nor U21083 (N_21083,N_17616,N_17001);
and U21084 (N_21084,N_18713,N_16771);
or U21085 (N_21085,N_18598,N_17394);
or U21086 (N_21086,N_15980,N_16119);
nor U21087 (N_21087,N_16002,N_18164);
nand U21088 (N_21088,N_17689,N_15977);
nor U21089 (N_21089,N_18259,N_18356);
or U21090 (N_21090,N_17877,N_15842);
nor U21091 (N_21091,N_17739,N_17126);
and U21092 (N_21092,N_16288,N_17316);
or U21093 (N_21093,N_16039,N_16522);
nor U21094 (N_21094,N_16392,N_16178);
nor U21095 (N_21095,N_16017,N_17876);
nor U21096 (N_21096,N_17143,N_17979);
and U21097 (N_21097,N_18111,N_17284);
and U21098 (N_21098,N_17688,N_18180);
nor U21099 (N_21099,N_17936,N_18496);
and U21100 (N_21100,N_18031,N_17594);
and U21101 (N_21101,N_18411,N_17049);
xnor U21102 (N_21102,N_17680,N_16716);
and U21103 (N_21103,N_18093,N_15735);
nor U21104 (N_21104,N_18193,N_18485);
nor U21105 (N_21105,N_18213,N_17519);
nand U21106 (N_21106,N_18237,N_16387);
and U21107 (N_21107,N_18190,N_17047);
nor U21108 (N_21108,N_16333,N_15786);
or U21109 (N_21109,N_18180,N_15643);
or U21110 (N_21110,N_16624,N_17515);
nand U21111 (N_21111,N_16838,N_16679);
or U21112 (N_21112,N_15729,N_18156);
or U21113 (N_21113,N_18270,N_15935);
nand U21114 (N_21114,N_18141,N_16515);
nand U21115 (N_21115,N_16920,N_18113);
xor U21116 (N_21116,N_16961,N_16562);
or U21117 (N_21117,N_16653,N_18079);
xor U21118 (N_21118,N_17296,N_16990);
or U21119 (N_21119,N_17536,N_16450);
nor U21120 (N_21120,N_18501,N_16380);
nor U21121 (N_21121,N_18124,N_18701);
and U21122 (N_21122,N_18378,N_18106);
and U21123 (N_21123,N_18029,N_16218);
and U21124 (N_21124,N_16643,N_16791);
nor U21125 (N_21125,N_15689,N_18364);
nand U21126 (N_21126,N_16649,N_16116);
and U21127 (N_21127,N_18728,N_18608);
nor U21128 (N_21128,N_16720,N_18169);
or U21129 (N_21129,N_16349,N_17556);
nor U21130 (N_21130,N_17450,N_16356);
nor U21131 (N_21131,N_18252,N_16588);
or U21132 (N_21132,N_17564,N_16453);
or U21133 (N_21133,N_17052,N_18083);
nor U21134 (N_21134,N_18032,N_16580);
nor U21135 (N_21135,N_16399,N_17734);
or U21136 (N_21136,N_18259,N_17914);
or U21137 (N_21137,N_16577,N_16005);
and U21138 (N_21138,N_18130,N_16136);
nand U21139 (N_21139,N_17364,N_16513);
or U21140 (N_21140,N_17502,N_18146);
nor U21141 (N_21141,N_18057,N_18543);
nand U21142 (N_21142,N_16611,N_18611);
xnor U21143 (N_21143,N_17350,N_16697);
and U21144 (N_21144,N_17379,N_17616);
nand U21145 (N_21145,N_15630,N_17816);
nor U21146 (N_21146,N_18226,N_15868);
xor U21147 (N_21147,N_16881,N_18355);
and U21148 (N_21148,N_17771,N_17197);
nor U21149 (N_21149,N_18308,N_17019);
nor U21150 (N_21150,N_16112,N_17534);
nand U21151 (N_21151,N_18742,N_15704);
nand U21152 (N_21152,N_18673,N_17013);
xnor U21153 (N_21153,N_17289,N_17557);
or U21154 (N_21154,N_15723,N_15858);
nand U21155 (N_21155,N_18401,N_16663);
xor U21156 (N_21156,N_18433,N_17053);
nand U21157 (N_21157,N_17974,N_17274);
or U21158 (N_21158,N_16423,N_17692);
and U21159 (N_21159,N_17700,N_16391);
and U21160 (N_21160,N_18429,N_16446);
nand U21161 (N_21161,N_16891,N_17130);
nand U21162 (N_21162,N_17909,N_17655);
nand U21163 (N_21163,N_17042,N_16345);
or U21164 (N_21164,N_17707,N_18275);
nor U21165 (N_21165,N_18556,N_16293);
nand U21166 (N_21166,N_16725,N_16601);
xnor U21167 (N_21167,N_16827,N_17245);
and U21168 (N_21168,N_18659,N_15706);
or U21169 (N_21169,N_16527,N_18068);
nor U21170 (N_21170,N_16047,N_17885);
nor U21171 (N_21171,N_16097,N_16215);
xnor U21172 (N_21172,N_17179,N_17855);
and U21173 (N_21173,N_15953,N_16985);
nor U21174 (N_21174,N_16725,N_15957);
and U21175 (N_21175,N_18354,N_17352);
or U21176 (N_21176,N_17076,N_17581);
nand U21177 (N_21177,N_17957,N_18233);
or U21178 (N_21178,N_17468,N_17636);
nand U21179 (N_21179,N_17416,N_16547);
or U21180 (N_21180,N_16437,N_17723);
or U21181 (N_21181,N_17926,N_15821);
nand U21182 (N_21182,N_16434,N_17931);
xnor U21183 (N_21183,N_18562,N_16288);
and U21184 (N_21184,N_16655,N_16464);
or U21185 (N_21185,N_18409,N_16282);
nor U21186 (N_21186,N_17899,N_18066);
or U21187 (N_21187,N_17421,N_18664);
and U21188 (N_21188,N_17452,N_16537);
and U21189 (N_21189,N_17140,N_18412);
nor U21190 (N_21190,N_16424,N_16428);
or U21191 (N_21191,N_18379,N_17891);
nand U21192 (N_21192,N_17637,N_17049);
and U21193 (N_21193,N_17783,N_17246);
nand U21194 (N_21194,N_16060,N_17837);
and U21195 (N_21195,N_17574,N_16028);
nor U21196 (N_21196,N_16153,N_18375);
or U21197 (N_21197,N_15803,N_17593);
and U21198 (N_21198,N_16441,N_15714);
xor U21199 (N_21199,N_16153,N_18230);
nor U21200 (N_21200,N_16382,N_15644);
and U21201 (N_21201,N_16117,N_18540);
and U21202 (N_21202,N_16577,N_15790);
nand U21203 (N_21203,N_16267,N_16859);
and U21204 (N_21204,N_17556,N_16514);
nor U21205 (N_21205,N_16536,N_18569);
or U21206 (N_21206,N_18230,N_16915);
xnor U21207 (N_21207,N_17384,N_16285);
nand U21208 (N_21208,N_15832,N_16128);
nor U21209 (N_21209,N_16153,N_17618);
and U21210 (N_21210,N_16932,N_16535);
and U21211 (N_21211,N_17914,N_18587);
nand U21212 (N_21212,N_18728,N_16076);
nand U21213 (N_21213,N_16866,N_16476);
nor U21214 (N_21214,N_18086,N_16259);
or U21215 (N_21215,N_18265,N_18351);
and U21216 (N_21216,N_15736,N_16454);
and U21217 (N_21217,N_15803,N_18669);
and U21218 (N_21218,N_17051,N_18491);
nor U21219 (N_21219,N_16803,N_16219);
and U21220 (N_21220,N_15971,N_18134);
xor U21221 (N_21221,N_16916,N_15928);
nand U21222 (N_21222,N_16374,N_16947);
nand U21223 (N_21223,N_17152,N_17853);
or U21224 (N_21224,N_17110,N_15796);
or U21225 (N_21225,N_18651,N_17131);
and U21226 (N_21226,N_16999,N_17107);
and U21227 (N_21227,N_16652,N_15850);
nor U21228 (N_21228,N_16807,N_18019);
and U21229 (N_21229,N_16511,N_17395);
or U21230 (N_21230,N_15745,N_15871);
and U21231 (N_21231,N_16482,N_17181);
nor U21232 (N_21232,N_17776,N_16926);
xor U21233 (N_21233,N_16477,N_18236);
nor U21234 (N_21234,N_18377,N_17812);
nand U21235 (N_21235,N_18022,N_16747);
xnor U21236 (N_21236,N_15795,N_17637);
or U21237 (N_21237,N_15822,N_18623);
or U21238 (N_21238,N_15649,N_17412);
or U21239 (N_21239,N_15697,N_16674);
or U21240 (N_21240,N_16272,N_17417);
nor U21241 (N_21241,N_16470,N_18418);
nor U21242 (N_21242,N_18137,N_15745);
nand U21243 (N_21243,N_18132,N_16574);
nor U21244 (N_21244,N_17466,N_17132);
nand U21245 (N_21245,N_16090,N_15660);
nand U21246 (N_21246,N_17705,N_17079);
nand U21247 (N_21247,N_15930,N_15992);
nor U21248 (N_21248,N_16486,N_16790);
or U21249 (N_21249,N_16433,N_17326);
nor U21250 (N_21250,N_17388,N_15783);
or U21251 (N_21251,N_15794,N_18492);
or U21252 (N_21252,N_15648,N_17956);
nand U21253 (N_21253,N_16892,N_16828);
nand U21254 (N_21254,N_18747,N_16043);
nand U21255 (N_21255,N_17674,N_17731);
and U21256 (N_21256,N_16226,N_16035);
xnor U21257 (N_21257,N_18383,N_18368);
nand U21258 (N_21258,N_17940,N_15738);
xnor U21259 (N_21259,N_16522,N_17583);
xor U21260 (N_21260,N_18460,N_17475);
nand U21261 (N_21261,N_17080,N_18555);
and U21262 (N_21262,N_16185,N_18337);
or U21263 (N_21263,N_18025,N_18679);
or U21264 (N_21264,N_16060,N_16220);
nor U21265 (N_21265,N_17557,N_18129);
nand U21266 (N_21266,N_15789,N_16452);
nor U21267 (N_21267,N_17983,N_18149);
nand U21268 (N_21268,N_16579,N_17198);
xnor U21269 (N_21269,N_16976,N_16721);
nand U21270 (N_21270,N_16097,N_16634);
nor U21271 (N_21271,N_17847,N_16863);
or U21272 (N_21272,N_15727,N_18417);
and U21273 (N_21273,N_17063,N_17024);
and U21274 (N_21274,N_18545,N_15899);
xnor U21275 (N_21275,N_16917,N_15688);
and U21276 (N_21276,N_18210,N_16421);
nor U21277 (N_21277,N_17129,N_17034);
nand U21278 (N_21278,N_16466,N_16259);
or U21279 (N_21279,N_18735,N_18480);
and U21280 (N_21280,N_17524,N_17948);
xor U21281 (N_21281,N_17215,N_15975);
or U21282 (N_21282,N_18430,N_17978);
nand U21283 (N_21283,N_15691,N_17512);
or U21284 (N_21284,N_18729,N_15948);
nand U21285 (N_21285,N_16869,N_16395);
and U21286 (N_21286,N_18512,N_16614);
and U21287 (N_21287,N_17063,N_18236);
xor U21288 (N_21288,N_17182,N_16611);
nand U21289 (N_21289,N_16476,N_16986);
xnor U21290 (N_21290,N_18471,N_16282);
xor U21291 (N_21291,N_17301,N_16554);
and U21292 (N_21292,N_16846,N_17055);
nor U21293 (N_21293,N_15886,N_17993);
xor U21294 (N_21294,N_17351,N_17641);
or U21295 (N_21295,N_16931,N_15990);
nand U21296 (N_21296,N_17371,N_18686);
xor U21297 (N_21297,N_17060,N_16862);
nor U21298 (N_21298,N_15900,N_17741);
nor U21299 (N_21299,N_17409,N_17890);
or U21300 (N_21300,N_15852,N_17914);
or U21301 (N_21301,N_17604,N_17019);
nand U21302 (N_21302,N_16597,N_15644);
nand U21303 (N_21303,N_16750,N_16870);
nor U21304 (N_21304,N_16593,N_16748);
xnor U21305 (N_21305,N_15688,N_18106);
xnor U21306 (N_21306,N_16035,N_15734);
xnor U21307 (N_21307,N_16219,N_16022);
nand U21308 (N_21308,N_17172,N_16403);
and U21309 (N_21309,N_16186,N_17135);
and U21310 (N_21310,N_16349,N_18709);
and U21311 (N_21311,N_18744,N_18409);
or U21312 (N_21312,N_16142,N_16957);
or U21313 (N_21313,N_18731,N_16924);
nor U21314 (N_21314,N_16462,N_18147);
nand U21315 (N_21315,N_17655,N_18551);
nand U21316 (N_21316,N_18236,N_16397);
nor U21317 (N_21317,N_16413,N_16274);
nor U21318 (N_21318,N_15884,N_16438);
nor U21319 (N_21319,N_16506,N_16312);
and U21320 (N_21320,N_15704,N_16470);
nor U21321 (N_21321,N_16114,N_17275);
or U21322 (N_21322,N_18204,N_17485);
xor U21323 (N_21323,N_16788,N_17475);
xor U21324 (N_21324,N_18068,N_15688);
nand U21325 (N_21325,N_17299,N_16687);
or U21326 (N_21326,N_18657,N_15939);
and U21327 (N_21327,N_17785,N_15648);
and U21328 (N_21328,N_18568,N_18584);
nand U21329 (N_21329,N_17699,N_16633);
or U21330 (N_21330,N_18488,N_16046);
xor U21331 (N_21331,N_15835,N_17779);
and U21332 (N_21332,N_15917,N_17727);
or U21333 (N_21333,N_17101,N_16776);
or U21334 (N_21334,N_18283,N_17787);
nor U21335 (N_21335,N_15934,N_16400);
nor U21336 (N_21336,N_18496,N_16105);
nor U21337 (N_21337,N_18670,N_17074);
nand U21338 (N_21338,N_16826,N_18328);
nand U21339 (N_21339,N_17775,N_18201);
xnor U21340 (N_21340,N_16391,N_17106);
or U21341 (N_21341,N_15956,N_16480);
or U21342 (N_21342,N_15743,N_18737);
nand U21343 (N_21343,N_16648,N_17397);
or U21344 (N_21344,N_16474,N_15929);
xnor U21345 (N_21345,N_16586,N_16768);
or U21346 (N_21346,N_16555,N_15757);
and U21347 (N_21347,N_17244,N_18162);
and U21348 (N_21348,N_16621,N_16027);
xnor U21349 (N_21349,N_15721,N_17711);
nand U21350 (N_21350,N_17184,N_18602);
or U21351 (N_21351,N_17367,N_16925);
xnor U21352 (N_21352,N_17742,N_17594);
nor U21353 (N_21353,N_18396,N_16618);
nand U21354 (N_21354,N_18423,N_16080);
nor U21355 (N_21355,N_18661,N_16459);
and U21356 (N_21356,N_18452,N_18359);
nand U21357 (N_21357,N_17975,N_18696);
nand U21358 (N_21358,N_18350,N_17010);
or U21359 (N_21359,N_18048,N_15693);
nand U21360 (N_21360,N_16127,N_16589);
nor U21361 (N_21361,N_18364,N_16051);
nand U21362 (N_21362,N_17799,N_18407);
nand U21363 (N_21363,N_17514,N_16247);
or U21364 (N_21364,N_17330,N_18063);
nand U21365 (N_21365,N_16395,N_16687);
xor U21366 (N_21366,N_16754,N_17298);
and U21367 (N_21367,N_17007,N_18416);
xnor U21368 (N_21368,N_17229,N_17615);
nor U21369 (N_21369,N_15664,N_18104);
nand U21370 (N_21370,N_16799,N_18314);
or U21371 (N_21371,N_15981,N_17248);
nand U21372 (N_21372,N_16034,N_15830);
or U21373 (N_21373,N_15983,N_18061);
and U21374 (N_21374,N_16766,N_16552);
xor U21375 (N_21375,N_17067,N_17461);
nand U21376 (N_21376,N_16819,N_17936);
nand U21377 (N_21377,N_17599,N_18362);
nor U21378 (N_21378,N_17209,N_17644);
nand U21379 (N_21379,N_18134,N_16843);
nor U21380 (N_21380,N_16910,N_16295);
or U21381 (N_21381,N_18596,N_18710);
or U21382 (N_21382,N_17495,N_18745);
or U21383 (N_21383,N_17349,N_16292);
or U21384 (N_21384,N_18547,N_15788);
nor U21385 (N_21385,N_15756,N_16148);
and U21386 (N_21386,N_17943,N_16834);
nand U21387 (N_21387,N_18372,N_16175);
nand U21388 (N_21388,N_17881,N_16395);
nor U21389 (N_21389,N_17341,N_16158);
nand U21390 (N_21390,N_17567,N_16896);
and U21391 (N_21391,N_15913,N_16798);
or U21392 (N_21392,N_17656,N_16930);
nand U21393 (N_21393,N_17220,N_18153);
or U21394 (N_21394,N_16316,N_17406);
nand U21395 (N_21395,N_18481,N_17583);
nor U21396 (N_21396,N_16149,N_16230);
nand U21397 (N_21397,N_16552,N_16936);
nand U21398 (N_21398,N_17218,N_17232);
and U21399 (N_21399,N_16493,N_17175);
and U21400 (N_21400,N_16635,N_16630);
nor U21401 (N_21401,N_17698,N_17676);
nand U21402 (N_21402,N_17621,N_16094);
nor U21403 (N_21403,N_17013,N_18066);
and U21404 (N_21404,N_16649,N_17182);
nand U21405 (N_21405,N_18738,N_18188);
or U21406 (N_21406,N_16112,N_17760);
and U21407 (N_21407,N_17831,N_17435);
and U21408 (N_21408,N_18672,N_18036);
nor U21409 (N_21409,N_16571,N_15790);
and U21410 (N_21410,N_17716,N_16532);
nor U21411 (N_21411,N_17615,N_17499);
or U21412 (N_21412,N_18027,N_17174);
nand U21413 (N_21413,N_17676,N_16604);
and U21414 (N_21414,N_16119,N_16668);
nor U21415 (N_21415,N_16593,N_15983);
or U21416 (N_21416,N_15677,N_17329);
nor U21417 (N_21417,N_16500,N_17073);
nand U21418 (N_21418,N_17308,N_18441);
xor U21419 (N_21419,N_16130,N_16799);
or U21420 (N_21420,N_16470,N_16902);
nand U21421 (N_21421,N_16407,N_17622);
and U21422 (N_21422,N_17638,N_16584);
nand U21423 (N_21423,N_18393,N_18525);
or U21424 (N_21424,N_18610,N_17439);
nor U21425 (N_21425,N_16656,N_17112);
or U21426 (N_21426,N_18518,N_15670);
or U21427 (N_21427,N_16357,N_17576);
xnor U21428 (N_21428,N_18253,N_16289);
nor U21429 (N_21429,N_17664,N_17404);
xor U21430 (N_21430,N_16067,N_15889);
nor U21431 (N_21431,N_15719,N_15935);
and U21432 (N_21432,N_17561,N_15633);
nand U21433 (N_21433,N_16989,N_18119);
nand U21434 (N_21434,N_16406,N_16753);
xnor U21435 (N_21435,N_16465,N_18363);
nand U21436 (N_21436,N_16056,N_16832);
nor U21437 (N_21437,N_18180,N_18663);
nor U21438 (N_21438,N_17923,N_18170);
nand U21439 (N_21439,N_17838,N_18430);
xnor U21440 (N_21440,N_16675,N_17403);
or U21441 (N_21441,N_17887,N_16323);
nor U21442 (N_21442,N_16236,N_16310);
or U21443 (N_21443,N_16270,N_17348);
or U21444 (N_21444,N_18277,N_17226);
nand U21445 (N_21445,N_16777,N_15674);
and U21446 (N_21446,N_16944,N_16859);
and U21447 (N_21447,N_17047,N_16920);
nor U21448 (N_21448,N_18468,N_18144);
nand U21449 (N_21449,N_17801,N_16293);
or U21450 (N_21450,N_17077,N_17477);
and U21451 (N_21451,N_17335,N_17464);
nor U21452 (N_21452,N_17215,N_16820);
nor U21453 (N_21453,N_16598,N_17213);
or U21454 (N_21454,N_18122,N_18000);
or U21455 (N_21455,N_18054,N_18728);
nand U21456 (N_21456,N_18524,N_16995);
nand U21457 (N_21457,N_18446,N_17309);
nor U21458 (N_21458,N_17021,N_16663);
and U21459 (N_21459,N_16958,N_18423);
xnor U21460 (N_21460,N_16615,N_18045);
or U21461 (N_21461,N_16930,N_16894);
nor U21462 (N_21462,N_17758,N_15912);
or U21463 (N_21463,N_17796,N_17143);
and U21464 (N_21464,N_17077,N_18246);
xor U21465 (N_21465,N_16345,N_17872);
nand U21466 (N_21466,N_17756,N_17246);
nand U21467 (N_21467,N_18149,N_17205);
nand U21468 (N_21468,N_17501,N_18526);
and U21469 (N_21469,N_17440,N_17936);
or U21470 (N_21470,N_17560,N_16113);
xnor U21471 (N_21471,N_16209,N_17893);
nand U21472 (N_21472,N_18457,N_18045);
and U21473 (N_21473,N_17347,N_18242);
and U21474 (N_21474,N_16851,N_17296);
nor U21475 (N_21475,N_17534,N_16475);
nor U21476 (N_21476,N_18507,N_17024);
and U21477 (N_21477,N_17370,N_18472);
or U21478 (N_21478,N_17297,N_18220);
nand U21479 (N_21479,N_17157,N_16766);
and U21480 (N_21480,N_18502,N_17796);
nand U21481 (N_21481,N_17891,N_17813);
nor U21482 (N_21482,N_17902,N_16759);
xor U21483 (N_21483,N_16514,N_18257);
nand U21484 (N_21484,N_15934,N_16692);
xor U21485 (N_21485,N_17465,N_17526);
or U21486 (N_21486,N_17364,N_15727);
nand U21487 (N_21487,N_17717,N_17423);
nand U21488 (N_21488,N_15698,N_18541);
or U21489 (N_21489,N_17540,N_18110);
and U21490 (N_21490,N_18675,N_18029);
and U21491 (N_21491,N_15800,N_18278);
nor U21492 (N_21492,N_18578,N_18392);
nand U21493 (N_21493,N_16239,N_16004);
xor U21494 (N_21494,N_16879,N_16037);
and U21495 (N_21495,N_16948,N_18185);
nor U21496 (N_21496,N_17204,N_16703);
xnor U21497 (N_21497,N_16373,N_17751);
and U21498 (N_21498,N_17052,N_17289);
nor U21499 (N_21499,N_17513,N_18486);
or U21500 (N_21500,N_17964,N_17247);
and U21501 (N_21501,N_17350,N_17629);
or U21502 (N_21502,N_16047,N_18701);
and U21503 (N_21503,N_16996,N_16040);
xor U21504 (N_21504,N_17697,N_18514);
nor U21505 (N_21505,N_17844,N_18461);
and U21506 (N_21506,N_15761,N_16755);
nor U21507 (N_21507,N_16917,N_17706);
and U21508 (N_21508,N_17232,N_18336);
nand U21509 (N_21509,N_16898,N_16641);
or U21510 (N_21510,N_15859,N_16861);
nand U21511 (N_21511,N_17379,N_17731);
xor U21512 (N_21512,N_16641,N_18724);
or U21513 (N_21513,N_18181,N_17277);
nand U21514 (N_21514,N_16677,N_17909);
nand U21515 (N_21515,N_18216,N_16915);
or U21516 (N_21516,N_16436,N_17488);
and U21517 (N_21517,N_16740,N_16340);
nand U21518 (N_21518,N_15743,N_17245);
or U21519 (N_21519,N_16987,N_16367);
nand U21520 (N_21520,N_17088,N_17563);
nor U21521 (N_21521,N_16969,N_15930);
nand U21522 (N_21522,N_17175,N_17126);
xnor U21523 (N_21523,N_17513,N_17017);
xor U21524 (N_21524,N_17967,N_15799);
nand U21525 (N_21525,N_15946,N_16792);
and U21526 (N_21526,N_16654,N_18121);
nand U21527 (N_21527,N_15905,N_16569);
or U21528 (N_21528,N_18187,N_17026);
or U21529 (N_21529,N_18217,N_16942);
or U21530 (N_21530,N_16283,N_17233);
or U21531 (N_21531,N_17049,N_18229);
nand U21532 (N_21532,N_17937,N_16383);
or U21533 (N_21533,N_16538,N_18214);
or U21534 (N_21534,N_17869,N_16524);
nor U21535 (N_21535,N_16494,N_16048);
xor U21536 (N_21536,N_17664,N_18604);
and U21537 (N_21537,N_17277,N_18145);
or U21538 (N_21538,N_17285,N_16909);
xnor U21539 (N_21539,N_16154,N_17847);
xor U21540 (N_21540,N_18586,N_15663);
nor U21541 (N_21541,N_17093,N_15751);
nor U21542 (N_21542,N_16725,N_16300);
and U21543 (N_21543,N_18541,N_18713);
or U21544 (N_21544,N_16343,N_18462);
xor U21545 (N_21545,N_16608,N_16784);
xnor U21546 (N_21546,N_18171,N_16720);
xnor U21547 (N_21547,N_16989,N_16198);
nor U21548 (N_21548,N_18631,N_18074);
or U21549 (N_21549,N_17734,N_18646);
nor U21550 (N_21550,N_16289,N_16223);
nor U21551 (N_21551,N_16289,N_15910);
nor U21552 (N_21552,N_16586,N_17629);
nand U21553 (N_21553,N_16354,N_16218);
or U21554 (N_21554,N_15863,N_18519);
nor U21555 (N_21555,N_17654,N_18712);
nor U21556 (N_21556,N_15747,N_17943);
nor U21557 (N_21557,N_18047,N_17797);
and U21558 (N_21558,N_17303,N_16775);
nor U21559 (N_21559,N_16692,N_16553);
and U21560 (N_21560,N_16188,N_18259);
nand U21561 (N_21561,N_16781,N_17510);
or U21562 (N_21562,N_17008,N_16203);
and U21563 (N_21563,N_16336,N_15775);
nor U21564 (N_21564,N_17570,N_16429);
nor U21565 (N_21565,N_18463,N_15902);
nor U21566 (N_21566,N_18492,N_17077);
nor U21567 (N_21567,N_16714,N_15970);
or U21568 (N_21568,N_17604,N_17736);
nor U21569 (N_21569,N_16342,N_16475);
and U21570 (N_21570,N_18067,N_15772);
nor U21571 (N_21571,N_16472,N_17046);
and U21572 (N_21572,N_18543,N_16486);
and U21573 (N_21573,N_16348,N_17429);
and U21574 (N_21574,N_17274,N_18501);
and U21575 (N_21575,N_18521,N_16350);
and U21576 (N_21576,N_17507,N_15902);
nor U21577 (N_21577,N_17867,N_18048);
or U21578 (N_21578,N_16128,N_18378);
and U21579 (N_21579,N_16585,N_18140);
nand U21580 (N_21580,N_18229,N_17556);
nor U21581 (N_21581,N_17591,N_15967);
nand U21582 (N_21582,N_18542,N_15986);
nand U21583 (N_21583,N_17027,N_18061);
and U21584 (N_21584,N_17030,N_17098);
nor U21585 (N_21585,N_16865,N_15940);
or U21586 (N_21586,N_17639,N_18106);
and U21587 (N_21587,N_18471,N_15974);
xnor U21588 (N_21588,N_16501,N_18508);
and U21589 (N_21589,N_18663,N_17628);
or U21590 (N_21590,N_17143,N_16665);
or U21591 (N_21591,N_18175,N_17574);
or U21592 (N_21592,N_18747,N_16081);
nor U21593 (N_21593,N_17152,N_16136);
and U21594 (N_21594,N_15749,N_18023);
nor U21595 (N_21595,N_18409,N_17641);
nand U21596 (N_21596,N_18433,N_17183);
and U21597 (N_21597,N_16376,N_15902);
nor U21598 (N_21598,N_16138,N_16699);
or U21599 (N_21599,N_16255,N_17428);
nor U21600 (N_21600,N_17221,N_18736);
nand U21601 (N_21601,N_18620,N_16028);
nor U21602 (N_21602,N_18294,N_15892);
nand U21603 (N_21603,N_16516,N_16735);
or U21604 (N_21604,N_15858,N_18404);
nand U21605 (N_21605,N_16303,N_16843);
nor U21606 (N_21606,N_17779,N_15984);
nor U21607 (N_21607,N_16700,N_15872);
and U21608 (N_21608,N_17067,N_18501);
nor U21609 (N_21609,N_16831,N_16310);
xnor U21610 (N_21610,N_17580,N_17180);
nand U21611 (N_21611,N_18267,N_17323);
or U21612 (N_21612,N_18375,N_18650);
and U21613 (N_21613,N_17567,N_16014);
and U21614 (N_21614,N_17018,N_16087);
and U21615 (N_21615,N_15648,N_18710);
nand U21616 (N_21616,N_15659,N_17309);
or U21617 (N_21617,N_16370,N_17236);
and U21618 (N_21618,N_18307,N_17938);
xor U21619 (N_21619,N_16376,N_17517);
xnor U21620 (N_21620,N_17377,N_17138);
xor U21621 (N_21621,N_16241,N_16107);
nor U21622 (N_21622,N_16478,N_18190);
and U21623 (N_21623,N_16616,N_17476);
or U21624 (N_21624,N_17124,N_17797);
or U21625 (N_21625,N_18618,N_16995);
or U21626 (N_21626,N_16212,N_16390);
or U21627 (N_21627,N_16002,N_18001);
nor U21628 (N_21628,N_15783,N_15732);
and U21629 (N_21629,N_15829,N_16752);
xor U21630 (N_21630,N_16080,N_16352);
nor U21631 (N_21631,N_16865,N_16055);
or U21632 (N_21632,N_17418,N_15676);
and U21633 (N_21633,N_18628,N_17412);
nor U21634 (N_21634,N_17732,N_16035);
or U21635 (N_21635,N_18448,N_17045);
nand U21636 (N_21636,N_17406,N_15875);
nor U21637 (N_21637,N_17472,N_17109);
xnor U21638 (N_21638,N_18703,N_16951);
and U21639 (N_21639,N_16557,N_17441);
and U21640 (N_21640,N_16017,N_18368);
xnor U21641 (N_21641,N_18389,N_17704);
nand U21642 (N_21642,N_17765,N_18722);
or U21643 (N_21643,N_16738,N_15933);
nor U21644 (N_21644,N_17873,N_16385);
and U21645 (N_21645,N_16230,N_18441);
nand U21646 (N_21646,N_17314,N_15811);
and U21647 (N_21647,N_17324,N_18471);
nand U21648 (N_21648,N_16222,N_17557);
nand U21649 (N_21649,N_17933,N_16776);
nor U21650 (N_21650,N_18261,N_17189);
nor U21651 (N_21651,N_17738,N_17462);
or U21652 (N_21652,N_17823,N_18290);
nand U21653 (N_21653,N_16112,N_18126);
nand U21654 (N_21654,N_16040,N_18137);
nor U21655 (N_21655,N_16003,N_17057);
nor U21656 (N_21656,N_15998,N_18685);
xor U21657 (N_21657,N_16478,N_17555);
nor U21658 (N_21658,N_16766,N_16229);
or U21659 (N_21659,N_18490,N_18498);
or U21660 (N_21660,N_17428,N_16179);
nand U21661 (N_21661,N_15776,N_17427);
nand U21662 (N_21662,N_17678,N_16343);
and U21663 (N_21663,N_17729,N_17894);
or U21664 (N_21664,N_16019,N_16222);
or U21665 (N_21665,N_17742,N_17191);
and U21666 (N_21666,N_15954,N_17358);
xnor U21667 (N_21667,N_17820,N_17861);
or U21668 (N_21668,N_16791,N_18549);
nand U21669 (N_21669,N_17678,N_16853);
xnor U21670 (N_21670,N_18684,N_16743);
and U21671 (N_21671,N_17768,N_16749);
nand U21672 (N_21672,N_18708,N_17539);
nand U21673 (N_21673,N_17741,N_17382);
or U21674 (N_21674,N_16211,N_17324);
nor U21675 (N_21675,N_18678,N_17966);
or U21676 (N_21676,N_17856,N_17328);
or U21677 (N_21677,N_17478,N_16711);
xnor U21678 (N_21678,N_15829,N_15866);
nor U21679 (N_21679,N_15805,N_17096);
and U21680 (N_21680,N_15659,N_16306);
nor U21681 (N_21681,N_15691,N_15870);
or U21682 (N_21682,N_18092,N_16866);
and U21683 (N_21683,N_17156,N_17825);
nor U21684 (N_21684,N_17003,N_16761);
nand U21685 (N_21685,N_18524,N_16949);
and U21686 (N_21686,N_18449,N_16076);
nor U21687 (N_21687,N_18112,N_18603);
nand U21688 (N_21688,N_17000,N_15743);
nor U21689 (N_21689,N_18109,N_16016);
nand U21690 (N_21690,N_16004,N_18076);
nand U21691 (N_21691,N_16210,N_17230);
or U21692 (N_21692,N_18558,N_18180);
nand U21693 (N_21693,N_17138,N_17953);
or U21694 (N_21694,N_18212,N_17060);
nor U21695 (N_21695,N_18679,N_18442);
xnor U21696 (N_21696,N_17082,N_18131);
nand U21697 (N_21697,N_16064,N_15713);
nor U21698 (N_21698,N_16543,N_15829);
nand U21699 (N_21699,N_17252,N_17875);
or U21700 (N_21700,N_16853,N_16085);
nand U21701 (N_21701,N_18452,N_16512);
nor U21702 (N_21702,N_15914,N_15718);
or U21703 (N_21703,N_15954,N_16132);
nand U21704 (N_21704,N_17893,N_17702);
xnor U21705 (N_21705,N_15775,N_17491);
xnor U21706 (N_21706,N_17318,N_15947);
nand U21707 (N_21707,N_17021,N_18749);
and U21708 (N_21708,N_18734,N_16504);
xor U21709 (N_21709,N_17767,N_17384);
and U21710 (N_21710,N_16744,N_18598);
nor U21711 (N_21711,N_16016,N_17716);
nand U21712 (N_21712,N_16135,N_17832);
nand U21713 (N_21713,N_16233,N_16976);
and U21714 (N_21714,N_16720,N_16911);
nor U21715 (N_21715,N_16677,N_16072);
and U21716 (N_21716,N_17201,N_16849);
and U21717 (N_21717,N_17511,N_15652);
or U21718 (N_21718,N_16389,N_17437);
nor U21719 (N_21719,N_18084,N_17217);
or U21720 (N_21720,N_16420,N_17218);
or U21721 (N_21721,N_15892,N_18553);
and U21722 (N_21722,N_16602,N_17877);
nand U21723 (N_21723,N_15629,N_17694);
xnor U21724 (N_21724,N_18181,N_17128);
or U21725 (N_21725,N_18624,N_18193);
or U21726 (N_21726,N_18455,N_16470);
nor U21727 (N_21727,N_17465,N_18104);
or U21728 (N_21728,N_18180,N_17477);
nand U21729 (N_21729,N_17745,N_16282);
and U21730 (N_21730,N_18692,N_16666);
nor U21731 (N_21731,N_16977,N_16563);
and U21732 (N_21732,N_17539,N_18740);
or U21733 (N_21733,N_15990,N_16440);
or U21734 (N_21734,N_17400,N_15703);
nand U21735 (N_21735,N_16365,N_16949);
xnor U21736 (N_21736,N_15981,N_16707);
nand U21737 (N_21737,N_17311,N_17703);
xnor U21738 (N_21738,N_17511,N_17709);
nor U21739 (N_21739,N_17018,N_17173);
and U21740 (N_21740,N_15992,N_18617);
nor U21741 (N_21741,N_17917,N_17090);
or U21742 (N_21742,N_17671,N_17528);
nand U21743 (N_21743,N_17606,N_17420);
and U21744 (N_21744,N_17490,N_16552);
and U21745 (N_21745,N_17938,N_16328);
nor U21746 (N_21746,N_18075,N_15935);
or U21747 (N_21747,N_17466,N_16987);
nor U21748 (N_21748,N_18693,N_15872);
and U21749 (N_21749,N_17503,N_16170);
nand U21750 (N_21750,N_15681,N_17448);
nand U21751 (N_21751,N_16832,N_16274);
or U21752 (N_21752,N_16541,N_18445);
or U21753 (N_21753,N_17539,N_15788);
nor U21754 (N_21754,N_17811,N_16123);
xor U21755 (N_21755,N_17115,N_17181);
and U21756 (N_21756,N_17193,N_16961);
nand U21757 (N_21757,N_17378,N_16144);
nand U21758 (N_21758,N_18716,N_17892);
nor U21759 (N_21759,N_16184,N_18383);
and U21760 (N_21760,N_16900,N_17549);
nor U21761 (N_21761,N_15934,N_16234);
nor U21762 (N_21762,N_15771,N_16976);
nand U21763 (N_21763,N_16494,N_18121);
nand U21764 (N_21764,N_18121,N_17456);
and U21765 (N_21765,N_16998,N_17666);
xnor U21766 (N_21766,N_15957,N_16603);
or U21767 (N_21767,N_18709,N_16078);
and U21768 (N_21768,N_17929,N_17065);
nand U21769 (N_21769,N_17694,N_16304);
nand U21770 (N_21770,N_16165,N_15929);
and U21771 (N_21771,N_17020,N_16536);
or U21772 (N_21772,N_17437,N_18633);
xor U21773 (N_21773,N_18267,N_15904);
and U21774 (N_21774,N_16842,N_16934);
nand U21775 (N_21775,N_17340,N_17088);
and U21776 (N_21776,N_17619,N_17520);
and U21777 (N_21777,N_15821,N_17274);
nand U21778 (N_21778,N_15701,N_17336);
nor U21779 (N_21779,N_16218,N_18393);
or U21780 (N_21780,N_16082,N_17160);
nor U21781 (N_21781,N_16523,N_17538);
and U21782 (N_21782,N_16046,N_17153);
or U21783 (N_21783,N_18644,N_16131);
xnor U21784 (N_21784,N_16010,N_17119);
and U21785 (N_21785,N_15753,N_16912);
nand U21786 (N_21786,N_17187,N_16056);
or U21787 (N_21787,N_18151,N_16313);
nor U21788 (N_21788,N_16896,N_18515);
nor U21789 (N_21789,N_17607,N_16830);
and U21790 (N_21790,N_18425,N_17234);
nand U21791 (N_21791,N_16349,N_18212);
nor U21792 (N_21792,N_16436,N_16098);
and U21793 (N_21793,N_17110,N_15671);
or U21794 (N_21794,N_16824,N_16682);
nand U21795 (N_21795,N_17770,N_16487);
and U21796 (N_21796,N_17097,N_15829);
nor U21797 (N_21797,N_18133,N_17658);
and U21798 (N_21798,N_18009,N_16409);
nor U21799 (N_21799,N_17661,N_17919);
xnor U21800 (N_21800,N_18043,N_18392);
or U21801 (N_21801,N_15771,N_17173);
or U21802 (N_21802,N_16842,N_16988);
xor U21803 (N_21803,N_17055,N_16286);
or U21804 (N_21804,N_17959,N_18450);
nand U21805 (N_21805,N_16299,N_17820);
or U21806 (N_21806,N_15820,N_16308);
or U21807 (N_21807,N_16059,N_16707);
or U21808 (N_21808,N_16494,N_17838);
nand U21809 (N_21809,N_16659,N_17638);
nand U21810 (N_21810,N_17489,N_15719);
or U21811 (N_21811,N_16007,N_18277);
nand U21812 (N_21812,N_18113,N_16852);
xor U21813 (N_21813,N_16838,N_17297);
nor U21814 (N_21814,N_17626,N_16216);
or U21815 (N_21815,N_16492,N_17690);
nand U21816 (N_21816,N_17177,N_16910);
or U21817 (N_21817,N_17771,N_17204);
or U21818 (N_21818,N_18639,N_17048);
nand U21819 (N_21819,N_16930,N_15646);
or U21820 (N_21820,N_17093,N_17751);
nand U21821 (N_21821,N_17868,N_17073);
or U21822 (N_21822,N_17506,N_17027);
and U21823 (N_21823,N_16285,N_17191);
or U21824 (N_21824,N_15803,N_16066);
nor U21825 (N_21825,N_17432,N_16794);
nand U21826 (N_21826,N_15795,N_16495);
nor U21827 (N_21827,N_17194,N_16925);
and U21828 (N_21828,N_18518,N_17869);
nand U21829 (N_21829,N_16104,N_17765);
nor U21830 (N_21830,N_16311,N_15803);
and U21831 (N_21831,N_16838,N_17916);
nor U21832 (N_21832,N_16146,N_17831);
nand U21833 (N_21833,N_16370,N_16631);
nor U21834 (N_21834,N_15798,N_17124);
nor U21835 (N_21835,N_17921,N_16221);
nor U21836 (N_21836,N_17697,N_16243);
or U21837 (N_21837,N_16503,N_15884);
or U21838 (N_21838,N_16542,N_17744);
and U21839 (N_21839,N_17251,N_17394);
xor U21840 (N_21840,N_18088,N_16372);
or U21841 (N_21841,N_16972,N_17098);
and U21842 (N_21842,N_16116,N_17121);
or U21843 (N_21843,N_15796,N_17188);
or U21844 (N_21844,N_17935,N_18353);
nand U21845 (N_21845,N_16105,N_18701);
and U21846 (N_21846,N_18456,N_17479);
and U21847 (N_21847,N_18221,N_18283);
or U21848 (N_21848,N_16245,N_16706);
xnor U21849 (N_21849,N_17767,N_16946);
and U21850 (N_21850,N_17642,N_16582);
nor U21851 (N_21851,N_18112,N_18090);
or U21852 (N_21852,N_16039,N_16260);
or U21853 (N_21853,N_18315,N_15849);
nor U21854 (N_21854,N_18631,N_17100);
and U21855 (N_21855,N_16517,N_15632);
nor U21856 (N_21856,N_17770,N_15951);
nor U21857 (N_21857,N_18111,N_18307);
nor U21858 (N_21858,N_17761,N_17141);
nor U21859 (N_21859,N_18087,N_16207);
nor U21860 (N_21860,N_17170,N_18462);
or U21861 (N_21861,N_17166,N_18616);
or U21862 (N_21862,N_17733,N_17769);
nor U21863 (N_21863,N_18421,N_16987);
and U21864 (N_21864,N_16676,N_16498);
nand U21865 (N_21865,N_18000,N_17324);
nor U21866 (N_21866,N_16902,N_17153);
xor U21867 (N_21867,N_16979,N_17815);
and U21868 (N_21868,N_17867,N_16844);
or U21869 (N_21869,N_16334,N_16393);
xnor U21870 (N_21870,N_18278,N_18409);
or U21871 (N_21871,N_16156,N_18481);
nor U21872 (N_21872,N_16273,N_16440);
nor U21873 (N_21873,N_16668,N_17747);
nand U21874 (N_21874,N_17819,N_17686);
or U21875 (N_21875,N_18803,N_21181);
or U21876 (N_21876,N_20694,N_19981);
nor U21877 (N_21877,N_19604,N_19398);
and U21878 (N_21878,N_18939,N_19381);
nand U21879 (N_21879,N_19690,N_20121);
or U21880 (N_21880,N_21463,N_21425);
nand U21881 (N_21881,N_19097,N_21050);
or U21882 (N_21882,N_19012,N_19758);
nor U21883 (N_21883,N_20253,N_19568);
and U21884 (N_21884,N_21360,N_18869);
nand U21885 (N_21885,N_20440,N_20296);
nor U21886 (N_21886,N_18875,N_19180);
or U21887 (N_21887,N_18752,N_21136);
nand U21888 (N_21888,N_20359,N_21279);
and U21889 (N_21889,N_19597,N_21631);
and U21890 (N_21890,N_20309,N_21722);
or U21891 (N_21891,N_20620,N_20517);
nand U21892 (N_21892,N_20918,N_21765);
nand U21893 (N_21893,N_20299,N_21156);
nand U21894 (N_21894,N_21025,N_20481);
nor U21895 (N_21895,N_18800,N_20449);
nor U21896 (N_21896,N_20738,N_20593);
xnor U21897 (N_21897,N_21599,N_20020);
or U21898 (N_21898,N_19327,N_19675);
or U21899 (N_21899,N_20109,N_19553);
nor U21900 (N_21900,N_18815,N_19799);
and U21901 (N_21901,N_18959,N_19533);
and U21902 (N_21902,N_20943,N_19020);
and U21903 (N_21903,N_21301,N_20644);
xnor U21904 (N_21904,N_19534,N_19850);
nor U21905 (N_21905,N_21310,N_19004);
xnor U21906 (N_21906,N_21217,N_21334);
xor U21907 (N_21907,N_20170,N_19696);
or U21908 (N_21908,N_21496,N_20342);
xor U21909 (N_21909,N_20500,N_21022);
nand U21910 (N_21910,N_20321,N_21501);
nand U21911 (N_21911,N_20165,N_20502);
nand U21912 (N_21912,N_20804,N_19703);
and U21913 (N_21913,N_18824,N_21677);
nand U21914 (N_21914,N_19495,N_19070);
and U21915 (N_21915,N_21013,N_21432);
nor U21916 (N_21916,N_20257,N_18776);
nor U21917 (N_21917,N_18955,N_20877);
nor U21918 (N_21918,N_20396,N_21758);
nand U21919 (N_21919,N_21570,N_20181);
or U21920 (N_21920,N_20624,N_20306);
nor U21921 (N_21921,N_19858,N_20975);
nor U21922 (N_21922,N_19793,N_21693);
or U21923 (N_21923,N_21093,N_18952);
and U21924 (N_21924,N_20681,N_19882);
and U21925 (N_21925,N_21158,N_20632);
xnor U21926 (N_21926,N_20643,N_18779);
nor U21927 (N_21927,N_20209,N_19844);
nand U21928 (N_21928,N_21518,N_18806);
and U21929 (N_21929,N_20154,N_21739);
nor U21930 (N_21930,N_19316,N_20808);
or U21931 (N_21931,N_20987,N_21733);
nand U21932 (N_21932,N_19454,N_19764);
nand U21933 (N_21933,N_20548,N_20035);
nor U21934 (N_21934,N_20001,N_21418);
and U21935 (N_21935,N_20485,N_20379);
nor U21936 (N_21936,N_20810,N_18837);
nand U21937 (N_21937,N_21014,N_19125);
nor U21938 (N_21938,N_19473,N_21191);
and U21939 (N_21939,N_21059,N_19985);
and U21940 (N_21940,N_20601,N_19284);
nor U21941 (N_21941,N_19252,N_21216);
or U21942 (N_21942,N_21430,N_19546);
and U21943 (N_21943,N_20460,N_19943);
or U21944 (N_21944,N_18798,N_20134);
and U21945 (N_21945,N_19245,N_20196);
xor U21946 (N_21946,N_20161,N_21340);
nor U21947 (N_21947,N_20639,N_20127);
nand U21948 (N_21948,N_20809,N_20085);
nor U21949 (N_21949,N_19267,N_21409);
nand U21950 (N_21950,N_20551,N_19126);
nand U21951 (N_21951,N_20111,N_20827);
or U21952 (N_21952,N_19967,N_21110);
nand U21953 (N_21953,N_18847,N_19328);
nand U21954 (N_21954,N_19140,N_19202);
nor U21955 (N_21955,N_18793,N_20026);
nand U21956 (N_21956,N_19156,N_19519);
nor U21957 (N_21957,N_19414,N_20673);
or U21958 (N_21958,N_21351,N_20842);
or U21959 (N_21959,N_21161,N_18820);
nor U21960 (N_21960,N_20276,N_21285);
xnor U21961 (N_21961,N_19053,N_20679);
or U21962 (N_21962,N_21659,N_20506);
nand U21963 (N_21963,N_19155,N_21610);
or U21964 (N_21964,N_19133,N_21069);
and U21965 (N_21965,N_20704,N_19806);
nand U21966 (N_21966,N_21778,N_19557);
and U21967 (N_21967,N_20578,N_20284);
xnor U21968 (N_21968,N_19132,N_19947);
xnor U21969 (N_21969,N_20378,N_18937);
nor U21970 (N_21970,N_20529,N_20742);
or U21971 (N_21971,N_20468,N_19246);
and U21972 (N_21972,N_20883,N_21754);
or U21973 (N_21973,N_19596,N_21336);
and U21974 (N_21974,N_18769,N_19626);
xor U21975 (N_21975,N_19410,N_20915);
and U21976 (N_21976,N_21005,N_21445);
xnor U21977 (N_21977,N_19804,N_19294);
nor U21978 (N_21978,N_19095,N_19725);
nor U21979 (N_21979,N_19777,N_20408);
nand U21980 (N_21980,N_18948,N_20323);
or U21981 (N_21981,N_21800,N_19067);
or U21982 (N_21982,N_21099,N_19279);
or U21983 (N_21983,N_19489,N_18942);
and U21984 (N_21984,N_21332,N_19555);
or U21985 (N_21985,N_19667,N_21745);
and U21986 (N_21986,N_21811,N_19408);
nand U21987 (N_21987,N_20508,N_18980);
or U21988 (N_21988,N_18788,N_19442);
and U21989 (N_21989,N_20988,N_21202);
xnor U21990 (N_21990,N_19605,N_19818);
or U21991 (N_21991,N_21578,N_21150);
nand U21992 (N_21992,N_21535,N_19382);
nor U21993 (N_21993,N_20743,N_21166);
nor U21994 (N_21994,N_19479,N_18977);
nor U21995 (N_21995,N_19162,N_19203);
nand U21996 (N_21996,N_21474,N_19647);
nand U21997 (N_21997,N_20903,N_20017);
nor U21998 (N_21998,N_20982,N_19213);
and U21999 (N_21999,N_21092,N_20854);
or U22000 (N_22000,N_21412,N_18960);
nand U22001 (N_22001,N_20554,N_21117);
or U22002 (N_22002,N_21625,N_20893);
and U22003 (N_22003,N_21580,N_19571);
nor U22004 (N_22004,N_19700,N_21483);
nand U22005 (N_22005,N_18920,N_18817);
nor U22006 (N_22006,N_20172,N_21742);
nand U22007 (N_22007,N_21818,N_20352);
xor U22008 (N_22008,N_20814,N_20906);
nand U22009 (N_22009,N_21807,N_19364);
nand U22010 (N_22010,N_21539,N_18970);
nand U22011 (N_22011,N_20431,N_21658);
and U22012 (N_22012,N_19225,N_20032);
or U22013 (N_22013,N_19201,N_19324);
nand U22014 (N_22014,N_20243,N_20163);
xor U22015 (N_22015,N_19431,N_20845);
and U22016 (N_22016,N_20876,N_20919);
or U22017 (N_22017,N_19288,N_19503);
nor U22018 (N_22018,N_19021,N_20687);
or U22019 (N_22019,N_21715,N_21169);
and U22020 (N_22020,N_20217,N_21195);
nor U22021 (N_22021,N_21065,N_19472);
xor U22022 (N_22022,N_20092,N_19405);
or U22023 (N_22023,N_21521,N_21495);
nand U22024 (N_22024,N_19109,N_21172);
and U22025 (N_22025,N_21121,N_19194);
nor U22026 (N_22026,N_20737,N_20900);
and U22027 (N_22027,N_20182,N_19154);
and U22028 (N_22028,N_19720,N_19560);
nor U22029 (N_22029,N_18968,N_21176);
nand U22030 (N_22030,N_19247,N_21643);
or U22031 (N_22031,N_19529,N_20291);
xor U22032 (N_22032,N_19061,N_18765);
nand U22033 (N_22033,N_20778,N_19144);
or U22034 (N_22034,N_20776,N_21324);
nand U22035 (N_22035,N_21633,N_18927);
or U22036 (N_22036,N_21615,N_19035);
xor U22037 (N_22037,N_20953,N_21687);
nand U22038 (N_22038,N_21583,N_19307);
or U22039 (N_22039,N_21477,N_19449);
or U22040 (N_22040,N_18963,N_19130);
or U22041 (N_22041,N_18854,N_20968);
xnor U22042 (N_22042,N_19153,N_19009);
nor U22043 (N_22043,N_20774,N_19370);
nand U22044 (N_22044,N_19372,N_21300);
or U22045 (N_22045,N_21469,N_20447);
nor U22046 (N_22046,N_18768,N_19358);
nand U22047 (N_22047,N_20666,N_20806);
and U22048 (N_22048,N_20357,N_20247);
xor U22049 (N_22049,N_21740,N_20912);
nor U22050 (N_22050,N_21016,N_21287);
and U22051 (N_22051,N_21009,N_21572);
and U22052 (N_22052,N_21037,N_21170);
nor U22053 (N_22053,N_19150,N_19709);
nor U22054 (N_22054,N_19893,N_20494);
nand U22055 (N_22055,N_20269,N_19927);
nand U22056 (N_22056,N_21002,N_21874);
nor U22057 (N_22057,N_20822,N_20581);
xor U22058 (N_22058,N_21288,N_20852);
or U22059 (N_22059,N_19903,N_21263);
or U22060 (N_22060,N_19822,N_19045);
nand U22061 (N_22061,N_20803,N_21138);
nand U22062 (N_22062,N_21188,N_20555);
nor U22063 (N_22063,N_20612,N_18792);
or U22064 (N_22064,N_21563,N_19369);
nand U22065 (N_22065,N_19664,N_19896);
and U22066 (N_22066,N_19309,N_21604);
or U22067 (N_22067,N_19206,N_20722);
or U22068 (N_22068,N_20927,N_21489);
nor U22069 (N_22069,N_18915,N_20627);
nand U22070 (N_22070,N_20300,N_20800);
and U22071 (N_22071,N_21204,N_21760);
nor U22072 (N_22072,N_18925,N_18995);
nor U22073 (N_22073,N_19867,N_21321);
nor U22074 (N_22074,N_21787,N_19627);
xnor U22075 (N_22075,N_20277,N_21338);
and U22076 (N_22076,N_21080,N_21061);
nor U22077 (N_22077,N_19505,N_21676);
nor U22078 (N_22078,N_20415,N_20260);
nor U22079 (N_22079,N_20335,N_18751);
nor U22080 (N_22080,N_19355,N_20333);
and U22081 (N_22081,N_19010,N_19456);
nor U22082 (N_22082,N_21809,N_20273);
and U22083 (N_22083,N_21319,N_20663);
nand U22084 (N_22084,N_21226,N_19524);
or U22085 (N_22085,N_21784,N_21690);
nor U22086 (N_22086,N_19025,N_20599);
or U22087 (N_22087,N_19030,N_21648);
nand U22088 (N_22088,N_19447,N_20347);
nor U22089 (N_22089,N_19727,N_19969);
nor U22090 (N_22090,N_19752,N_21184);
and U22091 (N_22091,N_21675,N_18958);
nor U22092 (N_22092,N_21804,N_19468);
nor U22093 (N_22093,N_21323,N_18954);
or U22094 (N_22094,N_21264,N_20685);
nor U22095 (N_22095,N_19390,N_20167);
nand U22096 (N_22096,N_21476,N_19165);
and U22097 (N_22097,N_20931,N_20048);
nand U22098 (N_22098,N_19464,N_20713);
nand U22099 (N_22099,N_19393,N_20414);
or U22100 (N_22100,N_19019,N_20527);
nor U22101 (N_22101,N_20563,N_19276);
or U22102 (N_22102,N_19746,N_21764);
xnor U22103 (N_22103,N_21045,N_19453);
or U22104 (N_22104,N_19711,N_19926);
xnor U22105 (N_22105,N_19513,N_21389);
or U22106 (N_22106,N_20138,N_18918);
or U22107 (N_22107,N_20073,N_19601);
and U22108 (N_22108,N_20311,N_21040);
and U22109 (N_22109,N_20049,N_20629);
nor U22110 (N_22110,N_21330,N_19600);
and U22111 (N_22111,N_21845,N_19821);
or U22112 (N_22112,N_19710,N_21327);
and U22113 (N_22113,N_21577,N_21132);
and U22114 (N_22114,N_20084,N_20761);
nor U22115 (N_22115,N_20202,N_20010);
nor U22116 (N_22116,N_19418,N_20326);
and U22117 (N_22117,N_19875,N_20360);
nor U22118 (N_22118,N_19535,N_21420);
nand U22119 (N_22119,N_19808,N_19840);
or U22120 (N_22120,N_19041,N_19643);
and U22121 (N_22121,N_19353,N_20298);
or U22122 (N_22122,N_19892,N_21183);
xnor U22123 (N_22123,N_19129,N_19987);
xor U22124 (N_22124,N_20823,N_19744);
nand U22125 (N_22125,N_21507,N_21637);
and U22126 (N_22126,N_20794,N_20861);
nor U22127 (N_22127,N_18883,N_21020);
nand U22128 (N_22128,N_19006,N_21433);
xnor U22129 (N_22129,N_20755,N_20495);
and U22130 (N_22130,N_20866,N_21666);
or U22131 (N_22131,N_20549,N_18951);
and U22132 (N_22132,N_21095,N_21545);
or U22133 (N_22133,N_20426,N_20319);
nor U22134 (N_22134,N_20331,N_20746);
or U22135 (N_22135,N_19598,N_20797);
xnor U22136 (N_22136,N_21066,N_20956);
or U22137 (N_22137,N_18829,N_21417);
nand U22138 (N_22138,N_19565,N_19787);
or U22139 (N_22139,N_19116,N_19174);
nor U22140 (N_22140,N_19959,N_21052);
and U22141 (N_22141,N_21556,N_19929);
and U22142 (N_22142,N_21791,N_21510);
or U22143 (N_22143,N_21243,N_18848);
nor U22144 (N_22144,N_20795,N_20130);
and U22145 (N_22145,N_20546,N_19491);
nand U22146 (N_22146,N_20516,N_20984);
and U22147 (N_22147,N_19567,N_21528);
nand U22148 (N_22148,N_19421,N_19237);
or U22149 (N_22149,N_19072,N_19948);
nand U22150 (N_22150,N_20853,N_21317);
or U22151 (N_22151,N_20902,N_21581);
and U22152 (N_22152,N_20290,N_19005);
or U22153 (N_22153,N_18997,N_20981);
nor U22154 (N_22154,N_20420,N_21182);
or U22155 (N_22155,N_20976,N_18865);
and U22156 (N_22156,N_21437,N_20540);
nand U22157 (N_22157,N_19602,N_20701);
nor U22158 (N_22158,N_20552,N_20507);
or U22159 (N_22159,N_19029,N_21485);
nand U22160 (N_22160,N_21326,N_21311);
nor U22161 (N_22161,N_19766,N_21214);
or U22162 (N_22162,N_21617,N_21361);
and U22163 (N_22163,N_20421,N_21869);
or U22164 (N_22164,N_21542,N_19349);
nor U22165 (N_22165,N_19320,N_20436);
nor U22166 (N_22166,N_19389,N_19363);
nor U22167 (N_22167,N_19343,N_19909);
nor U22168 (N_22168,N_18879,N_18907);
and U22169 (N_22169,N_21297,N_18984);
or U22170 (N_22170,N_21753,N_18860);
nand U22171 (N_22171,N_18876,N_20524);
nor U22172 (N_22172,N_20771,N_20171);
or U22173 (N_22173,N_20169,N_21159);
or U22174 (N_22174,N_21124,N_21442);
and U22175 (N_22175,N_19815,N_19993);
xor U22176 (N_22176,N_20236,N_21139);
nor U22177 (N_22177,N_21678,N_20242);
nand U22178 (N_22178,N_19348,N_20404);
or U22179 (N_22179,N_18809,N_20097);
xor U22180 (N_22180,N_20263,N_19190);
or U22181 (N_22181,N_21224,N_20938);
or U22182 (N_22182,N_20535,N_19526);
or U22183 (N_22183,N_19217,N_21431);
and U22184 (N_22184,N_20648,N_19558);
nor U22185 (N_22185,N_19119,N_21377);
nand U22186 (N_22186,N_19078,N_20005);
nor U22187 (N_22187,N_18914,N_21465);
xor U22188 (N_22188,N_19107,N_19439);
xnor U22189 (N_22189,N_19516,N_21587);
nor U22190 (N_22190,N_20185,N_21685);
or U22191 (N_22191,N_19285,N_20446);
nand U22192 (N_22192,N_20232,N_21509);
xor U22193 (N_22193,N_21428,N_21815);
and U22194 (N_22194,N_21702,N_19606);
or U22195 (N_22195,N_20231,N_20219);
nor U22196 (N_22196,N_20302,N_19114);
or U22197 (N_22197,N_19197,N_20106);
nand U22198 (N_22198,N_20952,N_20840);
nor U22199 (N_22199,N_21736,N_20641);
and U22200 (N_22200,N_21048,N_19876);
xor U22201 (N_22201,N_19232,N_20394);
xor U22202 (N_22202,N_19674,N_21266);
nor U22203 (N_22203,N_20891,N_21337);
or U22204 (N_22204,N_19055,N_20683);
nor U22205 (N_22205,N_20820,N_21567);
and U22206 (N_22206,N_21375,N_19617);
or U22207 (N_22207,N_20646,N_20634);
or U22208 (N_22208,N_21605,N_19427);
nand U22209 (N_22209,N_18943,N_20056);
and U22210 (N_22210,N_20621,N_20098);
nor U22211 (N_22211,N_18982,N_19968);
or U22212 (N_22212,N_20882,N_21211);
xor U22213 (N_22213,N_19152,N_19158);
nand U22214 (N_22214,N_19795,N_20412);
or U22215 (N_22215,N_21547,N_19322);
and U22216 (N_22216,N_20286,N_21459);
nor U22217 (N_22217,N_21096,N_18789);
or U22218 (N_22218,N_19792,N_21741);
nand U22219 (N_22219,N_19460,N_20002);
and U22220 (N_22220,N_21656,N_20509);
and U22221 (N_22221,N_21466,N_20004);
nand U22222 (N_22222,N_18807,N_20239);
and U22223 (N_22223,N_20235,N_21088);
nor U22224 (N_22224,N_19120,N_21616);
or U22225 (N_22225,N_20076,N_18753);
nand U22226 (N_22226,N_19919,N_20583);
nor U22227 (N_22227,N_20762,N_20884);
or U22228 (N_22228,N_21388,N_20285);
xor U22229 (N_22229,N_19687,N_19488);
and U22230 (N_22230,N_19612,N_20234);
and U22231 (N_22231,N_18972,N_21399);
or U22232 (N_22232,N_20177,N_20836);
and U22233 (N_22233,N_21557,N_21651);
xor U22234 (N_22234,N_21363,N_19031);
and U22235 (N_22235,N_19028,N_19255);
or U22236 (N_22236,N_21426,N_21628);
nor U22237 (N_22237,N_20969,N_20011);
nor U22238 (N_22238,N_20758,N_20736);
nand U22239 (N_22239,N_19734,N_20417);
nor U22240 (N_22240,N_19699,N_20033);
nor U22241 (N_22241,N_21108,N_19229);
and U22242 (N_22242,N_19113,N_18922);
and U22243 (N_22243,N_19798,N_21180);
or U22244 (N_22244,N_21667,N_21582);
nand U22245 (N_22245,N_21055,N_21374);
or U22246 (N_22246,N_19013,N_19333);
and U22247 (N_22247,N_20208,N_20675);
nor U22248 (N_22248,N_20512,N_18756);
nand U22249 (N_22249,N_18873,N_20728);
nand U22250 (N_22250,N_20091,N_20099);
or U22251 (N_22251,N_19728,N_20457);
or U22252 (N_22252,N_21186,N_18901);
nor U22253 (N_22253,N_18762,N_21554);
and U22254 (N_22254,N_18899,N_19058);
nand U22255 (N_22255,N_21700,N_19856);
and U22256 (N_22256,N_20199,N_20081);
or U22257 (N_22257,N_20513,N_21021);
nand U22258 (N_22258,N_19362,N_18826);
nand U22259 (N_22259,N_19345,N_20467);
or U22260 (N_22260,N_18992,N_19921);
nand U22261 (N_22261,N_19550,N_19216);
nand U22262 (N_22262,N_19480,N_20278);
nand U22263 (N_22263,N_20329,N_19003);
and U22264 (N_22264,N_19931,N_19088);
nand U22265 (N_22265,N_20668,N_19536);
nor U22266 (N_22266,N_21209,N_18956);
nand U22267 (N_22267,N_20933,N_19962);
nor U22268 (N_22268,N_19658,N_21320);
nand U22269 (N_22269,N_19471,N_21592);
nand U22270 (N_22270,N_20935,N_19951);
xor U22271 (N_22271,N_19040,N_19251);
xor U22272 (N_22272,N_20233,N_21562);
nand U22273 (N_22273,N_20454,N_19419);
nand U22274 (N_22274,N_20433,N_20107);
nand U22275 (N_22275,N_21705,N_20445);
xnor U22276 (N_22276,N_19737,N_21561);
or U22277 (N_22277,N_18814,N_21104);
nor U22278 (N_22278,N_20542,N_19134);
nor U22279 (N_22279,N_20006,N_20661);
and U22280 (N_22280,N_21611,N_21242);
nand U22281 (N_22281,N_20672,N_19494);
or U22282 (N_22282,N_21795,N_21467);
and U22283 (N_22283,N_18813,N_21732);
nor U22284 (N_22284,N_20047,N_19254);
nor U22285 (N_22285,N_20148,N_21039);
or U22286 (N_22286,N_19071,N_19124);
or U22287 (N_22287,N_18771,N_20784);
nor U22288 (N_22288,N_21590,N_20395);
xnor U22289 (N_22289,N_18851,N_21857);
or U22290 (N_22290,N_21316,N_18857);
nor U22291 (N_22291,N_19625,N_21298);
nand U22292 (N_22292,N_19809,N_20580);
or U22293 (N_22293,N_20030,N_20730);
nor U22294 (N_22294,N_19064,N_21642);
or U22295 (N_22295,N_19610,N_19044);
and U22296 (N_22296,N_19729,N_20218);
xor U22297 (N_22297,N_20305,N_18766);
xnor U22298 (N_22298,N_20294,N_19430);
and U22299 (N_22299,N_19677,N_19917);
nand U22300 (N_22300,N_20280,N_20287);
nand U22301 (N_22301,N_19650,N_21262);
nand U22302 (N_22302,N_21499,N_19960);
nand U22303 (N_22303,N_21373,N_21109);
nor U22304 (N_22304,N_19691,N_21506);
or U22305 (N_22305,N_19634,N_20455);
or U22306 (N_22306,N_19399,N_19540);
and U22307 (N_22307,N_18993,N_19995);
nor U22308 (N_22308,N_19790,N_20409);
xnor U22309 (N_22309,N_20860,N_19918);
and U22310 (N_22310,N_19038,N_20137);
nor U22311 (N_22311,N_21470,N_20929);
and U22312 (N_22312,N_19498,N_20867);
or U22313 (N_22313,N_18791,N_19397);
or U22314 (N_22314,N_19577,N_19544);
and U22315 (N_22315,N_19847,N_20203);
nor U22316 (N_22316,N_20832,N_21516);
nand U22317 (N_22317,N_19891,N_19539);
and U22318 (N_22318,N_20965,N_19905);
or U22319 (N_22319,N_20979,N_21566);
xnor U22320 (N_22320,N_21488,N_21386);
nor U22321 (N_22321,N_19683,N_21073);
nor U22322 (N_22322,N_19811,N_18944);
nand U22323 (N_22323,N_19853,N_21047);
and U22324 (N_22324,N_19308,N_20103);
or U22325 (N_22325,N_21291,N_20413);
nand U22326 (N_22326,N_19765,N_19378);
xnor U22327 (N_22327,N_21423,N_20080);
xor U22328 (N_22328,N_19256,N_20895);
and U22329 (N_22329,N_21457,N_20256);
and U22330 (N_22330,N_18988,N_18834);
nand U22331 (N_22331,N_18892,N_19230);
nor U22332 (N_22332,N_21801,N_19476);
and U22333 (N_22333,N_20270,N_21089);
or U22334 (N_22334,N_19936,N_20688);
nand U22335 (N_22335,N_19672,N_21460);
nor U22336 (N_22336,N_21768,N_21387);
or U22337 (N_22337,N_21662,N_19807);
nor U22338 (N_22338,N_20693,N_20514);
and U22339 (N_22339,N_18750,N_19933);
and U22340 (N_22340,N_19365,N_21709);
and U22341 (N_22341,N_21255,N_20961);
or U22342 (N_22342,N_19924,N_21011);
nor U22343 (N_22343,N_21820,N_19749);
nor U22344 (N_22344,N_21714,N_20957);
or U22345 (N_22345,N_18867,N_21012);
or U22346 (N_22346,N_21484,N_21663);
or U22347 (N_22347,N_19066,N_19296);
nand U22348 (N_22348,N_21620,N_19313);
xor U22349 (N_22349,N_19240,N_20619);
or U22350 (N_22350,N_20924,N_19830);
or U22351 (N_22351,N_21290,N_20677);
and U22352 (N_22352,N_18906,N_19923);
nand U22353 (N_22353,N_19863,N_20411);
and U22354 (N_22354,N_21726,N_20754);
and U22355 (N_22355,N_21381,N_20392);
nand U22356 (N_22356,N_21230,N_21372);
or U22357 (N_22357,N_21725,N_20125);
xor U22358 (N_22358,N_20928,N_19930);
nand U22359 (N_22359,N_19827,N_20427);
and U22360 (N_22360,N_21559,N_21223);
and U22361 (N_22361,N_20591,N_21036);
nand U22362 (N_22362,N_21771,N_18773);
or U22363 (N_22363,N_18767,N_20102);
or U22364 (N_22364,N_19406,N_20532);
and U22365 (N_22365,N_19289,N_18833);
nor U22366 (N_22366,N_19236,N_18830);
or U22367 (N_22367,N_19100,N_18872);
and U22368 (N_22368,N_21835,N_18933);
nand U22369 (N_22369,N_20139,N_19226);
xnor U22370 (N_22370,N_19175,N_19087);
or U22371 (N_22371,N_20096,N_20650);
nor U22372 (N_22372,N_21142,N_21537);
or U22373 (N_22373,N_20916,N_20123);
nand U22374 (N_22374,N_20977,N_20786);
nand U22375 (N_22375,N_19351,N_20131);
nand U22376 (N_22376,N_20012,N_21411);
or U22377 (N_22377,N_20301,N_21404);
or U22378 (N_22378,N_20633,N_20948);
nand U22379 (N_22379,N_19848,N_21086);
xnor U22380 (N_22380,N_20482,N_20921);
nor U22381 (N_22381,N_20147,N_19956);
nor U22382 (N_22382,N_19426,N_20946);
nor U22383 (N_22383,N_21382,N_21212);
nor U22384 (N_22384,N_21006,N_19299);
nor U22385 (N_22385,N_21862,N_20369);
and U22386 (N_22386,N_19051,N_20497);
or U22387 (N_22387,N_20843,N_19205);
nand U22388 (N_22388,N_19657,N_20279);
or U22389 (N_22389,N_19172,N_19511);
and U22390 (N_22390,N_20371,N_21679);
and U22391 (N_22391,N_21806,N_19177);
nor U22392 (N_22392,N_19527,N_20885);
or U22393 (N_22393,N_19545,N_20837);
nand U22394 (N_22394,N_19486,N_21817);
xor U22395 (N_22395,N_19591,N_21356);
nand U22396 (N_22396,N_20536,N_19586);
nand U22397 (N_22397,N_21640,N_18973);
or U22398 (N_22398,N_20429,N_20074);
or U22399 (N_22399,N_20223,N_20934);
nand U22400 (N_22400,N_19975,N_20989);
nor U22401 (N_22401,N_20873,N_20610);
xnor U22402 (N_22402,N_21538,N_20588);
and U22403 (N_22403,N_20267,N_19323);
nand U22404 (N_22404,N_21295,N_19263);
xor U22405 (N_22405,N_20225,N_19954);
xnor U22406 (N_22406,N_20191,N_21257);
nand U22407 (N_22407,N_18778,N_21129);
or U22408 (N_22408,N_20707,N_20733);
or U22409 (N_22409,N_20625,N_20700);
nand U22410 (N_22410,N_21201,N_18947);
nand U22411 (N_22411,N_21260,N_20732);
nor U22412 (N_22412,N_20892,N_21222);
nor U22413 (N_22413,N_21357,N_18930);
nand U22414 (N_22414,N_21552,N_19857);
nand U22415 (N_22415,N_21464,N_20558);
nand U22416 (N_22416,N_18775,N_19235);
or U22417 (N_22417,N_21534,N_19171);
xor U22418 (N_22418,N_21077,N_19339);
or U22419 (N_22419,N_21473,N_18821);
xor U22420 (N_22420,N_19089,N_21293);
or U22421 (N_22421,N_19692,N_20734);
or U22422 (N_22422,N_18924,N_19748);
nor U22423 (N_22423,N_20990,N_19668);
and U22424 (N_22424,N_19306,N_21500);
nor U22425 (N_22425,N_19761,N_20164);
nor U22426 (N_22426,N_21174,N_21478);
and U22427 (N_22427,N_21276,N_20040);
xor U22428 (N_22428,N_19566,N_21823);
xnor U22429 (N_22429,N_19779,N_21849);
nor U22430 (N_22430,N_19290,N_19594);
and U22431 (N_22431,N_18975,N_20325);
and U22432 (N_22432,N_18831,N_20197);
or U22433 (N_22433,N_20955,N_20553);
nand U22434 (N_22434,N_21249,N_19027);
and U22435 (N_22435,N_20520,N_20871);
or U22436 (N_22436,N_20462,N_19395);
or U22437 (N_22437,N_21712,N_21122);
nor U22438 (N_22438,N_20483,N_19481);
nand U22439 (N_22439,N_19271,N_21250);
nor U22440 (N_22440,N_20024,N_19781);
nand U22441 (N_22441,N_18796,N_20192);
nand U22442 (N_22442,N_20972,N_20567);
and U22443 (N_22443,N_19122,N_19118);
nand U22444 (N_22444,N_19671,N_19992);
and U22445 (N_22445,N_20490,N_20505);
nand U22446 (N_22446,N_21543,N_20013);
or U22447 (N_22447,N_20766,N_21299);
nor U22448 (N_22448,N_19257,N_19483);
nor U22449 (N_22449,N_19278,N_21403);
or U22450 (N_22450,N_19706,N_20416);
and U22451 (N_22451,N_18878,N_20652);
nor U22452 (N_22452,N_21342,N_21160);
nand U22453 (N_22453,N_21821,N_20116);
nand U22454 (N_22454,N_21352,N_21256);
nand U22455 (N_22455,N_21408,N_21789);
or U22456 (N_22456,N_19445,N_20828);
nor U22457 (N_22457,N_19743,N_19817);
xnor U22458 (N_22458,N_20992,N_20207);
or U22459 (N_22459,N_20367,N_21555);
nor U22460 (N_22460,N_19448,N_19778);
and U22461 (N_22461,N_19776,N_20067);
nor U22462 (N_22462,N_18964,N_21851);
nor U22463 (N_22463,N_18974,N_21167);
and U22464 (N_22464,N_21595,N_21008);
nand U22465 (N_22465,N_20941,N_21586);
and U22466 (N_22466,N_19945,N_18912);
nor U22467 (N_22467,N_19110,N_21051);
nor U22468 (N_22468,N_20135,N_19514);
nor U22469 (N_22469,N_20055,N_19356);
nor U22470 (N_22470,N_19074,N_20802);
and U22471 (N_22471,N_20783,N_19832);
and U22472 (N_22472,N_21824,N_19907);
nand U22473 (N_22473,N_21118,N_21720);
and U22474 (N_22474,N_19648,N_20503);
and U22475 (N_22475,N_20834,N_20105);
nor U22476 (N_22476,N_21208,N_19062);
nand U22477 (N_22477,N_21187,N_19241);
nor U22478 (N_22478,N_19715,N_20258);
nand U22479 (N_22479,N_21626,N_21145);
nor U22480 (N_22480,N_21271,N_21103);
xnor U22481 (N_22481,N_19249,N_20706);
or U22482 (N_22482,N_21629,N_19446);
nor U22483 (N_22483,N_18900,N_19127);
nand U22484 (N_22484,N_21834,N_18990);
nor U22485 (N_22485,N_20573,N_20274);
and U22486 (N_22486,N_19531,N_19797);
and U22487 (N_22487,N_19239,N_19898);
and U22488 (N_22488,N_19772,N_20117);
nor U22489 (N_22489,N_19723,N_21415);
and U22490 (N_22490,N_20949,N_21019);
and U22491 (N_22491,N_21826,N_21533);
or U22492 (N_22492,N_19970,N_19906);
and U22493 (N_22493,N_19002,N_19060);
or U22494 (N_22494,N_19443,N_19988);
xnor U22495 (N_22495,N_18799,N_20456);
nor U22496 (N_22496,N_19467,N_19024);
nor U22497 (N_22497,N_21522,N_19504);
or U22498 (N_22498,N_20194,N_19855);
or U22499 (N_22499,N_20077,N_18812);
nor U22500 (N_22500,N_21196,N_20970);
nand U22501 (N_22501,N_20721,N_21704);
nand U22502 (N_22502,N_18889,N_21102);
or U22503 (N_22503,N_21031,N_18953);
and U22504 (N_22504,N_19913,N_21618);
nor U22505 (N_22505,N_20140,N_20424);
nand U22506 (N_22506,N_21517,N_20855);
and U22507 (N_22507,N_20361,N_18790);
or U22508 (N_22508,N_19769,N_20993);
or U22509 (N_22509,N_21441,N_20264);
xnor U22510 (N_22510,N_20534,N_18763);
or U22511 (N_22511,N_21636,N_20533);
nor U22512 (N_22512,N_21402,N_19137);
and U22513 (N_22513,N_21328,N_20708);
nand U22514 (N_22514,N_20389,N_20151);
nor U22515 (N_22515,N_20757,N_21452);
or U22516 (N_22516,N_19938,N_19187);
or U22517 (N_22517,N_20691,N_20078);
and U22518 (N_22518,N_20348,N_21168);
or U22519 (N_22519,N_21770,N_21461);
nand U22520 (N_22520,N_18887,N_19705);
nand U22521 (N_22521,N_19678,N_20739);
nor U22522 (N_22522,N_20577,N_20910);
or U22523 (N_22523,N_21788,N_20724);
or U22524 (N_22524,N_20759,N_18885);
or U22525 (N_22525,N_19317,N_19050);
nand U22526 (N_22526,N_19157,N_19682);
xnor U22527 (N_22527,N_20660,N_19774);
nor U22528 (N_22528,N_21383,N_20126);
xor U22529 (N_22529,N_20215,N_20387);
nor U22530 (N_22530,N_18921,N_19195);
nor U22531 (N_22531,N_21866,N_19654);
or U22532 (N_22532,N_19694,N_21245);
xor U22533 (N_22533,N_21221,N_18819);
nor U22534 (N_22534,N_20113,N_21863);
and U22535 (N_22535,N_21085,N_19275);
nor U22536 (N_22536,N_20531,N_20519);
and U22537 (N_22537,N_19730,N_21270);
or U22538 (N_22538,N_20959,N_19063);
and U22539 (N_22539,N_20680,N_20149);
or U22540 (N_22540,N_21392,N_20166);
nor U22541 (N_22541,N_21035,N_20966);
nand U22542 (N_22542,N_20914,N_20362);
nor U22543 (N_22543,N_20623,N_20930);
nand U22544 (N_22544,N_20393,N_21588);
nand U22545 (N_22545,N_20595,N_21248);
and U22546 (N_22546,N_19388,N_21710);
and U22547 (N_22547,N_20665,N_19176);
xnor U22548 (N_22548,N_21125,N_20418);
nand U22549 (N_22549,N_21668,N_20603);
and U22550 (N_22550,N_20705,N_20478);
or U22551 (N_22551,N_21724,N_21623);
and U22552 (N_22552,N_20162,N_19211);
or U22553 (N_22553,N_21691,N_19963);
nor U22554 (N_22554,N_20332,N_18774);
or U22555 (N_22555,N_19911,N_19016);
or U22556 (N_22556,N_20526,N_21149);
or U22557 (N_22557,N_20390,N_21378);
nand U22558 (N_22558,N_20477,N_21773);
xnor U22559 (N_22559,N_21746,N_20386);
and U22560 (N_22560,N_20909,N_19816);
and U22561 (N_22561,N_20377,N_19966);
xnor U22562 (N_22562,N_20464,N_19735);
xor U22563 (N_22563,N_21007,N_21173);
nor U22564 (N_22564,N_18877,N_20571);
nand U22565 (N_22565,N_21068,N_19826);
or U22566 (N_22566,N_20168,N_20695);
or U22567 (N_22567,N_19042,N_21274);
nor U22568 (N_22568,N_21630,N_21371);
xor U22569 (N_22569,N_21070,N_19525);
and U22570 (N_22570,N_20061,N_21540);
and U22571 (N_22571,N_18858,N_20925);
nand U22572 (N_22572,N_19344,N_20770);
or U22573 (N_22573,N_19888,N_18757);
nand U22574 (N_22574,N_20604,N_21280);
and U22575 (N_22575,N_19588,N_19872);
nor U22576 (N_22576,N_19361,N_18781);
and U22577 (N_22577,N_20053,N_19470);
nand U22578 (N_22578,N_18810,N_20590);
nand U22579 (N_22579,N_21776,N_21769);
and U22580 (N_22580,N_20340,N_20031);
nand U22581 (N_22581,N_19338,N_19302);
or U22582 (N_22582,N_20330,N_20510);
and U22583 (N_22583,N_20110,N_19904);
or U22584 (N_22584,N_20570,N_20341);
nor U22585 (N_22585,N_21832,N_21689);
nor U22586 (N_22586,N_19043,N_19452);
and U22587 (N_22587,N_21672,N_19101);
or U22588 (N_22588,N_19075,N_21344);
or U22589 (N_22589,N_21434,N_20725);
nor U22590 (N_22590,N_19554,N_20851);
nor U22591 (N_22591,N_19587,N_20718);
and U22592 (N_22592,N_20384,N_20198);
nor U22593 (N_22593,N_21728,N_20338);
xnor U22594 (N_22594,N_18828,N_20865);
or U22595 (N_22595,N_19796,N_20385);
and U22596 (N_22596,N_21719,N_19139);
or U22597 (N_22597,N_19620,N_19712);
xnor U22598 (N_22598,N_19736,N_20289);
xnor U22599 (N_22599,N_19852,N_19173);
or U22600 (N_22600,N_21251,N_20801);
xnor U22601 (N_22601,N_19704,N_19552);
xor U22602 (N_22602,N_19726,N_21737);
or U22603 (N_22603,N_19656,N_20252);
nor U22604 (N_22604,N_19583,N_21283);
or U22605 (N_22605,N_19767,N_20423);
xnor U22606 (N_22606,N_21304,N_19582);
and U22607 (N_22607,N_21797,N_20997);
nand U22608 (N_22608,N_21254,N_19958);
nand U22609 (N_22609,N_19391,N_20674);
nor U22610 (N_22610,N_20484,N_20537);
and U22611 (N_22611,N_21438,N_21646);
nand U22612 (N_22612,N_19141,N_20696);
nand U22613 (N_22613,N_21796,N_19082);
nor U22614 (N_22614,N_20187,N_20796);
nand U22615 (N_22615,N_21652,N_20451);
nor U22616 (N_22616,N_21692,N_19652);
nand U22617 (N_22617,N_19999,N_19741);
xor U22618 (N_22618,N_19819,N_18882);
and U22619 (N_22619,N_20383,N_20750);
or U22620 (N_22620,N_18855,N_21775);
xnor U22621 (N_22621,N_21369,N_20962);
nor U22622 (N_22622,N_20474,N_19300);
nor U22623 (N_22623,N_21614,N_20498);
nand U22624 (N_22624,N_20281,N_21101);
and U22625 (N_22625,N_18863,N_21529);
xnor U22626 (N_22626,N_19637,N_21842);
or U22627 (N_22627,N_21861,N_19523);
or U22628 (N_22628,N_20336,N_19614);
nand U22629 (N_22629,N_20093,N_21090);
nor U22630 (N_22630,N_19559,N_21598);
nand U22631 (N_22631,N_20881,N_21046);
and U22632 (N_22632,N_21030,N_20714);
or U22633 (N_22633,N_21641,N_20744);
and U22634 (N_22634,N_21569,N_19572);
nor U22635 (N_22635,N_20283,N_19584);
xor U22636 (N_22636,N_19222,N_18870);
nor U22637 (N_22637,N_21503,N_20849);
and U22638 (N_22638,N_19592,N_19629);
or U22639 (N_22639,N_19360,N_20785);
nand U22640 (N_22640,N_19713,N_20115);
nand U22641 (N_22641,N_21841,N_19059);
and U22642 (N_22642,N_20450,N_18804);
and U22643 (N_22643,N_18908,N_20087);
nand U22644 (N_22644,N_21207,N_20238);
nand U22645 (N_22645,N_20419,N_20479);
nor U22646 (N_22646,N_21738,N_19780);
nor U22647 (N_22647,N_20402,N_19068);
nor U22648 (N_22648,N_20726,N_20631);
and U22649 (N_22649,N_19396,N_21205);
nor U22650 (N_22650,N_21015,N_20339);
xnor U22651 (N_22651,N_19258,N_18909);
and U22652 (N_22652,N_20582,N_19092);
xor U22653 (N_22653,N_21727,N_19820);
and U22654 (N_22654,N_20991,N_20150);
and U22655 (N_22655,N_20986,N_21860);
nor U22656 (N_22656,N_19312,N_20136);
xor U22657 (N_22657,N_19429,N_19547);
nor U22658 (N_22658,N_20435,N_19802);
and U22659 (N_22659,N_20821,N_21424);
and U22660 (N_22660,N_20453,N_19466);
or U22661 (N_22661,N_21443,N_18782);
or U22662 (N_22662,N_21471,N_19207);
nor U22663 (N_22663,N_20874,N_19618);
or U22664 (N_22664,N_21296,N_20574);
and U22665 (N_22665,N_20141,N_21854);
nor U22666 (N_22666,N_19653,N_20844);
nand U22667 (N_22667,N_21695,N_21364);
and U22668 (N_22668,N_19091,N_19651);
and U22669 (N_22669,N_20717,N_19649);
nand U22670 (N_22670,N_18881,N_21153);
nor U22671 (N_22671,N_21370,N_21657);
nand U22672 (N_22672,N_19394,N_19805);
xnor U22673 (N_22673,N_21157,N_20391);
nand U22674 (N_22674,N_18890,N_21038);
nand U22675 (N_22675,N_20936,N_18903);
or U22676 (N_22676,N_19221,N_19662);
and U22677 (N_22677,N_21127,N_20568);
nand U22678 (N_22678,N_18961,N_19794);
and U22679 (N_22679,N_18957,N_20444);
nor U22680 (N_22680,N_20790,N_19384);
and U22681 (N_22681,N_19739,N_21227);
or U22682 (N_22682,N_20857,N_19889);
nand U22683 (N_22683,N_21843,N_21435);
and U22684 (N_22684,N_21723,N_19838);
and U22685 (N_22685,N_20833,N_19457);
or U22686 (N_22686,N_18965,N_20101);
and U22687 (N_22687,N_19842,N_19094);
nand U22688 (N_22688,N_20014,N_19233);
nand U22689 (N_22689,N_19693,N_19166);
nand U22690 (N_22690,N_21579,N_21143);
nor U22691 (N_22691,N_19812,N_20054);
nor U22692 (N_22692,N_21120,N_18935);
or U22693 (N_22693,N_21401,N_20222);
and U22694 (N_22694,N_20373,N_20939);
and U22695 (N_22695,N_21458,N_21790);
nor U22696 (N_22696,N_19846,N_21225);
and U22697 (N_22697,N_19920,N_19996);
nor U22698 (N_22698,N_20124,N_21619);
xnor U22699 (N_22699,N_21472,N_21353);
xnor U22700 (N_22700,N_21318,N_21721);
nand U22701 (N_22701,N_18926,N_19944);
and U22702 (N_22702,N_19714,N_19093);
and U22703 (N_22703,N_20355,N_20259);
nor U22704 (N_22704,N_21491,N_20587);
and U22705 (N_22705,N_21743,N_21343);
and U22706 (N_22706,N_20316,N_21779);
nand U22707 (N_22707,N_20070,N_19775);
nor U22708 (N_22708,N_19666,N_18981);
nand U22709 (N_22709,N_18895,N_20476);
or U22710 (N_22710,N_19864,N_20050);
and U22711 (N_22711,N_19458,N_19900);
xnor U22712 (N_22712,N_20251,N_20923);
nor U22713 (N_22713,N_20817,N_19352);
xnor U22714 (N_22714,N_21833,N_19751);
xor U22715 (N_22715,N_19575,N_20351);
nor U22716 (N_22716,N_19803,N_21067);
or U22717 (N_22717,N_20607,N_20859);
xor U22718 (N_22718,N_19056,N_19849);
and U22719 (N_22719,N_19274,N_19178);
and U22720 (N_22720,N_21203,N_19104);
nor U22721 (N_22721,N_21144,N_19701);
or U22722 (N_22722,N_19484,N_20597);
and U22723 (N_22723,N_21839,N_19789);
nand U22724 (N_22724,N_20152,N_20647);
nor U22725 (N_22725,N_20372,N_20839);
nor U22726 (N_22726,N_20716,N_19814);
and U22727 (N_22727,N_21277,N_21783);
nor U22728 (N_22728,N_21694,N_21376);
and U22729 (N_22729,N_21278,N_19638);
nand U22730 (N_22730,N_21141,N_21044);
or U22731 (N_22731,N_20594,N_20178);
nor U22732 (N_22732,N_20037,N_20886);
or U22733 (N_22733,N_21349,N_19301);
nand U22734 (N_22734,N_21855,N_19433);
nand U22735 (N_22735,N_21131,N_21645);
or U22736 (N_22736,N_20942,N_19702);
and U22737 (N_22737,N_19159,N_21750);
nand U22738 (N_22738,N_20100,N_19782);
nand U22739 (N_22739,N_20220,N_20153);
nor U22740 (N_22740,N_21341,N_19542);
and U22741 (N_22741,N_21812,N_21384);
xnor U22742 (N_22742,N_20062,N_19444);
nand U22743 (N_22743,N_20007,N_21060);
xor U22744 (N_22744,N_20789,N_20848);
nand U22745 (N_22745,N_20904,N_21234);
xor U22746 (N_22746,N_21550,N_19015);
nand U22747 (N_22747,N_21856,N_20042);
and U22748 (N_22748,N_19490,N_19350);
and U22749 (N_22749,N_19196,N_21275);
and U22750 (N_22750,N_19635,N_21647);
xnor U22751 (N_22751,N_21140,N_21634);
nand U22752 (N_22752,N_19599,N_19371);
nor U22753 (N_22753,N_20768,N_20272);
nand U22754 (N_22754,N_19576,N_19955);
nand U22755 (N_22755,N_19564,N_21215);
nand U22756 (N_22756,N_20345,N_20428);
and U22757 (N_22757,N_20541,N_20227);
nand U22758 (N_22758,N_18919,N_18931);
or U22759 (N_22759,N_21236,N_18971);
or U22760 (N_22760,N_21265,N_20617);
or U22761 (N_22761,N_20995,N_20288);
nor U22762 (N_22762,N_20133,N_21063);
nand U22763 (N_22763,N_19506,N_21847);
xnor U22764 (N_22764,N_19425,N_20328);
and U22765 (N_22765,N_19054,N_21130);
or U22766 (N_22766,N_19259,N_19983);
or U22767 (N_22767,N_20388,N_21508);
nand U22768 (N_22768,N_18845,N_21218);
or U22769 (N_22769,N_19319,N_21147);
or U22770 (N_22770,N_21660,N_21701);
nor U22771 (N_22771,N_19624,N_20618);
nor U22772 (N_22772,N_20064,N_20664);
or U22773 (N_22773,N_20144,N_21154);
and U22774 (N_22774,N_20868,N_20913);
and U22775 (N_22775,N_20229,N_20547);
or U22776 (N_22776,N_19437,N_20818);
or U22777 (N_22777,N_19184,N_20856);
nor U22778 (N_22778,N_21708,N_21444);
or U22779 (N_22779,N_21808,N_20132);
and U22780 (N_22780,N_21071,N_20205);
and U22781 (N_22781,N_20066,N_18818);
or U22782 (N_22782,N_21368,N_18976);
xnor U22783 (N_22783,N_21683,N_20015);
xor U22784 (N_22784,N_20947,N_21192);
or U22785 (N_22785,N_21447,N_19182);
or U22786 (N_22786,N_19633,N_21644);
nor U22787 (N_22787,N_19147,N_20188);
and U22788 (N_22788,N_19537,N_21269);
or U22789 (N_22789,N_18772,N_20826);
or U22790 (N_22790,N_20983,N_21439);
xor U22791 (N_22791,N_19916,N_21003);
nand U22792 (N_22792,N_18898,N_20812);
or U22793 (N_22793,N_19902,N_20523);
and U22794 (N_22794,N_20221,N_21305);
xnor U22795 (N_22795,N_18794,N_20753);
nor U22796 (N_22796,N_21075,N_20815);
or U22797 (N_22797,N_21751,N_20830);
nor U22798 (N_22798,N_20626,N_20926);
or U22799 (N_22799,N_19167,N_19641);
and U22800 (N_22800,N_19084,N_21419);
xnor U22801 (N_22801,N_19434,N_19894);
nand U22802 (N_22802,N_19989,N_20616);
and U22803 (N_22803,N_20058,N_19543);
nor U22804 (N_22804,N_21347,N_21390);
nand U22805 (N_22805,N_19117,N_19990);
nor U22806 (N_22806,N_21115,N_21451);
or U22807 (N_22807,N_21624,N_19556);
nor U22808 (N_22808,N_20438,N_20611);
or U22809 (N_22809,N_19722,N_19784);
nor U22810 (N_22810,N_19138,N_19270);
xnor U22811 (N_22811,N_19688,N_20813);
or U22812 (N_22812,N_20317,N_19961);
xor U22813 (N_22813,N_21571,N_21653);
nor U22814 (N_22814,N_21654,N_21358);
nor U22815 (N_22815,N_18989,N_19630);
or U22816 (N_22816,N_18759,N_20690);
and U22817 (N_22817,N_19515,N_21837);
nand U22818 (N_22818,N_21486,N_21024);
nor U22819 (N_22819,N_20448,N_21766);
and U22820 (N_22820,N_20798,N_21175);
and U22821 (N_22821,N_19801,N_20888);
nand U22822 (N_22822,N_19199,N_20569);
and U22823 (N_22823,N_19756,N_20337);
nor U22824 (N_22824,N_19763,N_21134);
nand U22825 (N_22825,N_20237,N_21128);
nor U22826 (N_22826,N_19561,N_21852);
or U22827 (N_22827,N_19914,N_19681);
or U22828 (N_22828,N_19310,N_20556);
nand U22829 (N_22829,N_19994,N_21238);
or U22830 (N_22830,N_20592,N_21831);
and U22831 (N_22831,N_21544,N_19859);
and U22832 (N_22832,N_20312,N_19883);
nand U22833 (N_22833,N_19478,N_18844);
or U22834 (N_22834,N_20403,N_20266);
or U22835 (N_22835,N_18805,N_19500);
or U22836 (N_22836,N_21688,N_20937);
nand U22837 (N_22837,N_19507,N_20304);
and U22838 (N_22838,N_18985,N_19487);
or U22839 (N_22839,N_20008,N_20028);
and U22840 (N_22840,N_20441,N_19409);
or U22841 (N_22841,N_19788,N_19164);
xnor U22842 (N_22842,N_20082,N_20715);
and U22843 (N_22843,N_18825,N_21850);
and U22844 (N_22844,N_18886,N_20994);
or U22845 (N_22845,N_19870,N_19932);
and U22846 (N_22846,N_19485,N_20896);
or U22847 (N_22847,N_20343,N_19357);
and U22848 (N_22848,N_19359,N_19385);
and U22849 (N_22849,N_21468,N_20712);
nor U22850 (N_22850,N_20767,N_19950);
and U22851 (N_22851,N_20747,N_20905);
nand U22852 (N_22852,N_19023,N_20698);
nand U22853 (N_22853,N_20667,N_19168);
nor U22854 (N_22854,N_19839,N_19603);
xnor U22855 (N_22855,N_21482,N_19977);
and U22856 (N_22856,N_21492,N_21001);
nand U22857 (N_22857,N_21532,N_20346);
and U22858 (N_22858,N_21840,N_18835);
nor U22859 (N_22859,N_20201,N_21608);
nand U22860 (N_22860,N_21531,N_21414);
nand U22861 (N_22861,N_19655,N_21116);
nor U22862 (N_22862,N_19595,N_21872);
nor U22863 (N_22863,N_18780,N_21761);
nor U22864 (N_22864,N_21600,N_19014);
nor U22865 (N_22865,N_20249,N_21237);
or U22866 (N_22866,N_19387,N_20586);
nor U22867 (N_22867,N_21098,N_20676);
nand U22868 (N_22868,N_21100,N_21028);
and U22869 (N_22869,N_19183,N_20944);
nand U22870 (N_22870,N_19880,N_21126);
nor U22871 (N_22871,N_21339,N_20773);
xnor U22872 (N_22872,N_21546,N_21042);
nand U22873 (N_22873,N_21429,N_19644);
xor U22874 (N_22874,N_20657,N_19277);
or U22875 (N_22875,N_19493,N_20752);
nor U22876 (N_22876,N_21462,N_21232);
and U22877 (N_22877,N_20781,N_19972);
or U22878 (N_22878,N_20211,N_18983);
nand U22879 (N_22879,N_19204,N_20470);
xor U22880 (N_22880,N_21713,N_21380);
xnor U22881 (N_22881,N_20729,N_20907);
xnor U22882 (N_22882,N_20999,N_21830);
nor U22883 (N_22883,N_21220,N_20963);
nor U22884 (N_22884,N_20176,N_19851);
xor U22885 (N_22885,N_21706,N_19745);
and U22886 (N_22886,N_21548,N_20282);
nand U22887 (N_22887,N_21699,N_19033);
and U22888 (N_22888,N_19342,N_19619);
and U22889 (N_22889,N_21056,N_21057);
nand U22890 (N_22890,N_20320,N_21497);
xor U22891 (N_22891,N_19615,N_21367);
nand U22892 (N_22892,N_20120,N_19768);
nand U22893 (N_22893,N_18929,N_20562);
xnor U22894 (N_22894,N_21346,N_19499);
or U22895 (N_22895,N_20723,N_21155);
nor U22896 (N_22896,N_20642,N_19402);
or U22897 (N_22897,N_21524,N_21574);
or U22898 (N_22898,N_18864,N_21609);
xor U22899 (N_22899,N_20019,N_21774);
xor U22900 (N_22900,N_21043,N_20075);
nor U22901 (N_22901,N_19106,N_20405);
nor U22902 (N_22902,N_20370,N_20475);
nor U22903 (N_22903,N_20173,N_21785);
nor U22904 (N_22904,N_19915,N_20945);
and U22905 (N_22905,N_18802,N_19336);
nor U22906 (N_22906,N_18850,N_20879);
nand U22907 (N_22907,N_21199,N_19897);
and U22908 (N_22908,N_21078,N_20561);
xnor U22909 (N_22909,N_20465,N_19304);
nand U22910 (N_22910,N_20213,N_19331);
xor U22911 (N_22911,N_20160,N_20230);
and U22912 (N_22912,N_19076,N_21819);
nor U22913 (N_22913,N_19080,N_19136);
nor U22914 (N_22914,N_21680,N_21512);
or U22915 (N_22915,N_21853,N_19551);
nor U22916 (N_22916,N_20069,N_19791);
nor U22917 (N_22917,N_20684,N_19874);
or U22918 (N_22918,N_20656,N_19272);
nor U22919 (N_22919,N_21825,N_20838);
nand U22920 (N_22920,N_20059,N_21193);
xnor U22921 (N_22921,N_21200,N_21481);
xnor U22922 (N_22922,N_21671,N_19411);
nor U22923 (N_22923,N_19253,N_21292);
nand U22924 (N_22924,N_20564,N_19569);
nand U22925 (N_22925,N_19135,N_20088);
nand U22926 (N_22926,N_18923,N_19841);
nor U22927 (N_22927,N_21558,N_18816);
or U22928 (N_22928,N_19099,N_20023);
and U22929 (N_22929,N_20608,N_20089);
or U22930 (N_22930,N_19908,N_20374);
or U22931 (N_22931,N_20292,N_19432);
and U22932 (N_22932,N_21606,N_20057);
and U22933 (N_22933,N_20114,N_20442);
nand U22934 (N_22934,N_20072,N_19757);
xnor U22935 (N_22935,N_20246,N_20572);
or U22936 (N_22936,N_20193,N_21494);
or U22937 (N_22937,N_20271,N_20824);
xnor U22938 (N_22938,N_21859,N_21197);
nand U22939 (N_22939,N_19979,N_20740);
nor U22940 (N_22940,N_19632,N_20775);
or U22941 (N_22941,N_18938,N_20763);
nand U22942 (N_22942,N_18842,N_19148);
and U22943 (N_22943,N_21597,N_20655);
or U22944 (N_22944,N_19708,N_19039);
or U22945 (N_22945,N_18862,N_19034);
and U22946 (N_22946,N_21247,N_21798);
nand U22947 (N_22947,N_21072,N_19474);
nand U22948 (N_22948,N_18940,N_18786);
or U22949 (N_22949,N_20958,N_20609);
nor U22950 (N_22950,N_21772,N_19008);
and U22951 (N_22951,N_19760,N_21306);
or U22952 (N_22952,N_18795,N_19669);
or U22953 (N_22953,N_19719,N_21454);
and U22954 (N_22954,N_19562,N_21406);
or U22955 (N_22955,N_21514,N_20980);
nor U22956 (N_22956,N_19242,N_19198);
nand U22957 (N_22957,N_19860,N_19834);
or U22958 (N_22958,N_21252,N_21198);
nand U22959 (N_22959,N_21749,N_21594);
nor U22960 (N_22960,N_19262,N_20142);
or U22961 (N_22961,N_21793,N_20887);
xnor U22962 (N_22962,N_18979,N_21844);
nor U22963 (N_22963,N_21627,N_21246);
or U22964 (N_22964,N_19146,N_18941);
or U22965 (N_22965,N_21734,N_20122);
xnor U22966 (N_22966,N_21716,N_20709);
and U22967 (N_22967,N_20265,N_20364);
or U22968 (N_22968,N_21632,N_19368);
or U22969 (N_22969,N_18770,N_18871);
nor U22970 (N_22970,N_20911,N_19001);
nand U22971 (N_22971,N_19522,N_21397);
or U22972 (N_22972,N_19170,N_20897);
nor U22973 (N_22973,N_18836,N_19079);
nor U22974 (N_22974,N_21703,N_19502);
nor U22975 (N_22975,N_19477,N_21707);
and U22976 (N_22976,N_18962,N_20322);
or U22977 (N_22977,N_20525,N_21239);
nor U22978 (N_22978,N_20112,N_19465);
nor U22979 (N_22979,N_19496,N_20731);
and U22980 (N_22980,N_18894,N_21325);
nor U22981 (N_22981,N_20027,N_20071);
nand U22982 (N_22982,N_20649,N_21487);
nand U22983 (N_22983,N_19698,N_20985);
nand U22984 (N_22984,N_19836,N_20353);
nor U22985 (N_22985,N_19878,N_21805);
or U22986 (N_22986,N_19949,N_21829);
and U22987 (N_22987,N_21350,N_21113);
or U22988 (N_22988,N_19215,N_19639);
nand U22989 (N_22989,N_20344,N_20579);
or U22990 (N_22990,N_20443,N_19046);
nor U22991 (N_22991,N_18888,N_20086);
or U22992 (N_22992,N_20469,N_20407);
nor U22993 (N_22993,N_20241,N_20504);
nand U22994 (N_22994,N_20295,N_19689);
nand U22995 (N_22995,N_21560,N_20406);
nor U22996 (N_22996,N_19305,N_20602);
or U22997 (N_22997,N_20720,N_19912);
nand U22998 (N_22998,N_19011,N_19679);
and U22999 (N_22999,N_18758,N_20787);
and U23000 (N_23000,N_21449,N_20769);
and U23001 (N_23001,N_20862,N_21858);
and U23002 (N_23002,N_19685,N_19837);
and U23003 (N_23003,N_19971,N_21613);
and U23004 (N_23004,N_21267,N_21074);
xnor U23005 (N_23005,N_19895,N_20901);
nor U23006 (N_23006,N_19281,N_20399);
or U23007 (N_23007,N_18897,N_20458);
and U23008 (N_23008,N_20434,N_21490);
nor U23009 (N_23009,N_21405,N_20670);
nand U23010 (N_23010,N_21241,N_19753);
nor U23011 (N_23011,N_18823,N_20518);
or U23012 (N_23012,N_20636,N_20422);
nand U23013 (N_23013,N_21612,N_18808);
nor U23014 (N_23014,N_21711,N_21673);
nand U23015 (N_23015,N_18911,N_20268);
or U23016 (N_23016,N_20605,N_20245);
nor U23017 (N_23017,N_20682,N_19510);
xnor U23018 (N_23018,N_20128,N_19697);
nor U23019 (N_23019,N_21273,N_19590);
nor U23020 (N_23020,N_19877,N_21244);
and U23021 (N_23021,N_20354,N_21762);
and U23022 (N_23022,N_19622,N_19991);
or U23023 (N_23023,N_21004,N_21450);
nand U23024 (N_23024,N_20560,N_20045);
or U23025 (N_23025,N_20043,N_19661);
nand U23026 (N_23026,N_20158,N_18801);
xor U23027 (N_23027,N_19742,N_19833);
and U23028 (N_23028,N_20466,N_21171);
or U23029 (N_23029,N_20825,N_21289);
or U23030 (N_23030,N_18994,N_19145);
nor U23031 (N_23031,N_21698,N_20307);
or U23032 (N_23032,N_20792,N_20799);
or U23033 (N_23033,N_20459,N_19354);
and U23034 (N_23034,N_21268,N_21272);
nand U23035 (N_23035,N_21584,N_21747);
xor U23036 (N_23036,N_19407,N_21054);
and U23037 (N_23037,N_19581,N_20777);
and U23038 (N_23038,N_21194,N_19998);
or U23039 (N_23039,N_21034,N_19048);
or U23040 (N_23040,N_20829,N_20974);
nor U23041 (N_23041,N_19738,N_19191);
nand U23042 (N_23042,N_19018,N_19461);
nor U23043 (N_23043,N_19330,N_21049);
and U23044 (N_23044,N_21729,N_21752);
xnor U23045 (N_23045,N_19492,N_19283);
xor U23046 (N_23046,N_19026,N_19280);
nor U23047 (N_23047,N_20226,N_19549);
or U23048 (N_23048,N_19321,N_18949);
nor U23049 (N_23049,N_19022,N_18868);
and U23050 (N_23050,N_20908,N_21794);
xnor U23051 (N_23051,N_19450,N_19828);
and U23052 (N_23052,N_18902,N_21697);
or U23053 (N_23053,N_19081,N_21573);
and U23054 (N_23054,N_20375,N_18967);
nand U23055 (N_23055,N_19593,N_18832);
or U23056 (N_23056,N_19282,N_20538);
nor U23057 (N_23057,N_19436,N_19825);
nand U23058 (N_23058,N_20240,N_19111);
nand U23059 (N_23059,N_21137,N_20869);
and U23060 (N_23060,N_20889,N_20356);
nor U23061 (N_23061,N_21686,N_19438);
nand U23062 (N_23062,N_21836,N_19403);
or U23063 (N_23063,N_21650,N_21593);
or U23064 (N_23064,N_20671,N_20917);
or U23065 (N_23065,N_19532,N_21799);
nand U23066 (N_23066,N_21568,N_21670);
or U23067 (N_23067,N_19508,N_19973);
and U23068 (N_23068,N_21151,N_19223);
and U23069 (N_23069,N_19530,N_19451);
nand U23070 (N_23070,N_20314,N_21394);
or U23071 (N_23071,N_20692,N_19747);
nand U23072 (N_23072,N_19640,N_18853);
nor U23073 (N_23073,N_21087,N_19731);
and U23074 (N_23074,N_20598,N_21777);
nand U23075 (N_23075,N_20000,N_21229);
nand U23076 (N_23076,N_20334,N_19528);
nand U23077 (N_23077,N_19380,N_20297);
nand U23078 (N_23078,N_18783,N_18934);
and U23079 (N_23079,N_19098,N_21827);
nand U23080 (N_23080,N_21041,N_20539);
or U23081 (N_23081,N_20036,N_18755);
or U23082 (N_23082,N_20363,N_19810);
or U23083 (N_23083,N_19298,N_20846);
nor U23084 (N_23084,N_20932,N_19631);
and U23085 (N_23085,N_20606,N_19228);
nor U23086 (N_23086,N_21307,N_19935);
or U23087 (N_23087,N_21165,N_20003);
nand U23088 (N_23088,N_20628,N_20156);
or U23089 (N_23089,N_19073,N_21162);
or U23090 (N_23090,N_18880,N_20183);
or U23091 (N_23091,N_20318,N_21062);
and U23092 (N_23092,N_21359,N_19623);
or U23093 (N_23093,N_20119,N_19417);
nor U23094 (N_23094,N_19160,N_19260);
and U23095 (N_23095,N_18764,N_19227);
xor U23096 (N_23096,N_18913,N_19754);
nand U23097 (N_23097,N_21591,N_19188);
xor U23098 (N_23098,N_20878,N_20366);
nor U23099 (N_23099,N_21755,N_19268);
or U23100 (N_23100,N_19142,N_21133);
nor U23101 (N_23101,N_20250,N_21308);
and U23102 (N_23102,N_20973,N_18760);
nor U23103 (N_23103,N_19563,N_19108);
and U23104 (N_23104,N_19269,N_20174);
nand U23105 (N_23105,N_21029,N_21258);
xor U23106 (N_23106,N_19783,N_20041);
nor U23107 (N_23107,N_20492,N_18838);
nand U23108 (N_23108,N_19718,N_21603);
xor U23109 (N_23109,N_21231,N_20044);
or U23110 (N_23110,N_18999,N_20425);
xnor U23111 (N_23111,N_21314,N_18852);
or U23112 (N_23112,N_19940,N_19585);
nand U23113 (N_23113,N_20473,N_20184);
nor U23114 (N_23114,N_19210,N_19412);
nand U23115 (N_23115,N_19469,N_19952);
nand U23116 (N_23116,N_20397,N_19314);
xnor U23117 (N_23117,N_21553,N_21455);
or U23118 (N_23118,N_18893,N_20922);
nor U23119 (N_23119,N_21146,N_21767);
or U23120 (N_23120,N_20228,N_20180);
xor U23121 (N_23121,N_21526,N_20596);
nor U23122 (N_23122,N_21440,N_20254);
nand U23123 (N_23123,N_19244,N_21398);
nor U23124 (N_23124,N_19037,N_19248);
nor U23125 (N_23125,N_20950,N_18841);
and U23126 (N_23126,N_20157,N_19318);
and U23127 (N_23127,N_20016,N_19383);
and U23128 (N_23128,N_20864,N_19112);
nor U23129 (N_23129,N_19415,N_20711);
nand U23130 (N_23130,N_19570,N_19986);
nand U23131 (N_23131,N_21185,N_19861);
xnor U23132 (N_23132,N_21718,N_21097);
and U23133 (N_23133,N_19400,N_20960);
nand U23134 (N_23134,N_21219,N_20293);
and U23135 (N_23135,N_20212,N_19036);
xnor U23136 (N_23136,N_20095,N_18874);
and U23137 (N_23137,N_20600,N_19341);
and U23138 (N_23138,N_20491,N_21865);
and U23139 (N_23139,N_19401,N_20793);
nand U23140 (N_23140,N_18840,N_20489);
or U23141 (N_23141,N_19965,N_19939);
nand U23142 (N_23142,N_19663,N_21504);
nand U23143 (N_23143,N_19234,N_19243);
or U23144 (N_23144,N_19642,N_20630);
or U23145 (N_23145,N_20068,N_19209);
nor U23146 (N_23146,N_18811,N_19750);
xor U23147 (N_23147,N_20760,N_19684);
nand U23148 (N_23148,N_21870,N_19311);
or U23149 (N_23149,N_19934,N_21601);
nand U23150 (N_23150,N_21094,N_18936);
or U23151 (N_23151,N_20576,N_21410);
nand U23152 (N_23152,N_20480,N_20654);
nand U23153 (N_23153,N_19976,N_19941);
or U23154 (N_23154,N_21081,N_21366);
xor U23155 (N_23155,N_18910,N_19375);
nand U23156 (N_23156,N_19416,N_20039);
xnor U23157 (N_23157,N_19192,N_21802);
nand U23158 (N_23158,N_21119,N_21228);
nor U23159 (N_23159,N_20565,N_19367);
nor U23160 (N_23160,N_21748,N_19910);
and U23161 (N_23161,N_20735,N_20145);
nor U23162 (N_23162,N_19771,N_20376);
and U23163 (N_23163,N_20034,N_21079);
or U23164 (N_23164,N_21333,N_19161);
and U23165 (N_23165,N_19925,N_19266);
or U23166 (N_23166,N_19000,N_19901);
nor U23167 (N_23167,N_19574,N_19974);
or U23168 (N_23168,N_21446,N_20381);
nand U23169 (N_23169,N_20559,N_21407);
nor U23170 (N_23170,N_19422,N_20051);
and U23171 (N_23171,N_19957,N_21513);
nand U23172 (N_23172,N_21240,N_19785);
xnor U23173 (N_23173,N_20175,N_20719);
nor U23174 (N_23174,N_21493,N_21033);
and U23175 (N_23175,N_19090,N_19676);
nor U23176 (N_23176,N_20756,N_20009);
nor U23177 (N_23177,N_19660,N_19169);
nor U23178 (N_23178,N_20368,N_20544);
xnor U23179 (N_23179,N_21027,N_20622);
nand U23180 (N_23180,N_21622,N_19813);
or U23181 (N_23181,N_18784,N_21782);
or U23182 (N_23182,N_21822,N_19086);
and U23183 (N_23183,N_20614,N_20400);
or U23184 (N_23184,N_18785,N_21864);
nand U23185 (N_23185,N_21781,N_21456);
and U23186 (N_23186,N_20589,N_20038);
nand U23187 (N_23187,N_19686,N_18849);
nor U23188 (N_23188,N_20206,N_19424);
or U23189 (N_23189,N_20108,N_21813);
or U23190 (N_23190,N_18996,N_19325);
or U23191 (N_23191,N_20584,N_20303);
and U23192 (N_23192,N_19611,N_21322);
and U23193 (N_23193,N_20262,N_19501);
nand U23194 (N_23194,N_19121,N_19845);
nand U23195 (N_23195,N_21585,N_19609);
and U23196 (N_23196,N_20214,N_19659);
nand U23197 (N_23197,N_19007,N_19580);
and U23198 (N_23198,N_19373,N_21421);
nand U23199 (N_23199,N_19250,N_21064);
nand U23200 (N_23200,N_21527,N_19326);
nand U23201 (N_23201,N_20637,N_19047);
nand U23202 (N_23202,N_21177,N_20496);
xnor U23203 (N_23203,N_20566,N_21076);
nor U23204 (N_23204,N_19303,N_21635);
nor U23205 (N_23205,N_19346,N_19548);
or U23206 (N_23206,N_19366,N_19866);
nor U23207 (N_23207,N_20699,N_21511);
and U23208 (N_23208,N_20488,N_18991);
nor U23209 (N_23209,N_20349,N_19287);
nand U23210 (N_23210,N_21365,N_20835);
or U23211 (N_23211,N_20850,N_20653);
nor U23212 (N_23212,N_19717,N_21846);
and U23213 (N_23213,N_21810,N_21523);
nand U23214 (N_23214,N_20788,N_21520);
nand U23215 (N_23215,N_20748,N_19512);
nand U23216 (N_23216,N_19297,N_20880);
nor U23217 (N_23217,N_19964,N_19193);
nor U23218 (N_23218,N_21393,N_19123);
nor U23219 (N_23219,N_19065,N_19131);
nor U23220 (N_23220,N_21210,N_21763);
or U23221 (N_23221,N_19721,N_19869);
and U23222 (N_23222,N_20204,N_19759);
nand U23223 (N_23223,N_19497,N_21313);
and U23224 (N_23224,N_19520,N_20710);
nand U23225 (N_23225,N_19428,N_20046);
nand U23226 (N_23226,N_19862,N_19128);
nand U23227 (N_23227,N_20779,N_20638);
xnor U23228 (N_23228,N_19829,N_20382);
and U23229 (N_23229,N_19578,N_19873);
nor U23230 (N_23230,N_21602,N_21848);
nor U23231 (N_23231,N_19423,N_21759);
and U23232 (N_23232,N_21565,N_19261);
nor U23233 (N_23233,N_20380,N_21479);
nor U23234 (N_23234,N_19335,N_19329);
or U23235 (N_23235,N_21541,N_20764);
or U23236 (N_23236,N_21284,N_20613);
and U23237 (N_23237,N_19238,N_21735);
nor U23238 (N_23238,N_18998,N_19835);
and U23239 (N_23239,N_20898,N_19212);
and U23240 (N_23240,N_21253,N_19334);
nor U23241 (N_23241,N_20635,N_20678);
nor U23242 (N_23242,N_21355,N_18945);
nor U23243 (N_23243,N_19608,N_21576);
nor U23244 (N_23244,N_20021,N_21084);
nor U23245 (N_23245,N_18846,N_20486);
or U23246 (N_23246,N_21649,N_20063);
and U23247 (N_23247,N_21017,N_20315);
nand U23248 (N_23248,N_21422,N_19332);
and U23249 (N_23249,N_20324,N_18891);
and U23250 (N_23250,N_21661,N_21436);
nand U23251 (N_23251,N_21621,N_21286);
nor U23252 (N_23252,N_21786,N_20702);
nand U23253 (N_23253,N_19208,N_21235);
nand U23254 (N_23254,N_21498,N_21838);
nor U23255 (N_23255,N_20018,N_19636);
or U23256 (N_23256,N_21018,N_20689);
nand U23257 (N_23257,N_20261,N_18797);
nand U23258 (N_23258,N_20430,N_18966);
and U23259 (N_23259,N_19102,N_21163);
nor U23260 (N_23260,N_18928,N_21281);
and U23261 (N_23261,N_21549,N_19224);
xor U23262 (N_23262,N_20772,N_21259);
nand U23263 (N_23263,N_20749,N_20437);
and U23264 (N_23264,N_20858,N_19286);
nand U23265 (N_23265,N_20872,N_20920);
or U23266 (N_23266,N_19573,N_19613);
or U23267 (N_23267,N_19085,N_21329);
or U23268 (N_23268,N_20439,N_20511);
nor U23269 (N_23269,N_21744,N_18987);
and U23270 (N_23270,N_21792,N_19455);
and U23271 (N_23271,N_21756,N_21354);
or U23272 (N_23272,N_19463,N_21607);
nand U23273 (N_23273,N_20461,N_20971);
or U23274 (N_23274,N_21515,N_20870);
nand U23275 (N_23275,N_19200,N_20200);
and U23276 (N_23276,N_20255,N_20585);
nand U23277 (N_23277,N_21639,N_21575);
nand U23278 (N_23278,N_18978,N_20195);
nand U23279 (N_23279,N_20805,N_19899);
nand U23280 (N_23280,N_18787,N_21135);
or U23281 (N_23281,N_19273,N_19953);
nor U23282 (N_23282,N_20398,N_19032);
nand U23283 (N_23283,N_19770,N_21731);
and U23284 (N_23284,N_19762,N_19997);
nor U23285 (N_23285,N_21525,N_20327);
nor U23286 (N_23286,N_21867,N_19978);
nand U23287 (N_23287,N_21164,N_20819);
nor U23288 (N_23288,N_21282,N_20210);
or U23289 (N_23289,N_19379,N_21505);
and U23290 (N_23290,N_21111,N_21427);
or U23291 (N_23291,N_19854,N_21475);
nor U23292 (N_23292,N_19509,N_18777);
nor U23293 (N_23293,N_19115,N_20452);
nand U23294 (N_23294,N_19946,N_20894);
nor U23295 (N_23295,N_19984,N_20847);
nand U23296 (N_23296,N_19293,N_20501);
and U23297 (N_23297,N_19186,N_20155);
and U23298 (N_23298,N_19404,N_20493);
nand U23299 (N_23299,N_21400,N_21696);
or U23300 (N_23300,N_21480,N_20807);
nand U23301 (N_23301,N_19017,N_20248);
or U23302 (N_23302,N_18986,N_19214);
xor U23303 (N_23303,N_19823,N_19843);
and U23304 (N_23304,N_19149,N_21309);
xnor U23305 (N_23305,N_19218,N_20471);
or U23306 (N_23306,N_21026,N_19680);
or U23307 (N_23307,N_19420,N_19052);
nand U23308 (N_23308,N_18969,N_20515);
nor U23309 (N_23309,N_20244,N_20651);
nand U23310 (N_23310,N_20765,N_19374);
or U23311 (N_23311,N_19482,N_20967);
or U23312 (N_23312,N_19083,N_21413);
and U23313 (N_23313,N_21757,N_19231);
nand U23314 (N_23314,N_19386,N_20522);
and U23315 (N_23315,N_20432,N_21335);
or U23316 (N_23316,N_18861,N_19340);
nand U23317 (N_23317,N_19441,N_19096);
and U23318 (N_23318,N_21107,N_21682);
xor U23319 (N_23319,N_18916,N_18950);
xnor U23320 (N_23320,N_21303,N_18932);
nand U23321 (N_23321,N_19143,N_20940);
nor U23322 (N_23322,N_20186,N_18843);
nand U23323 (N_23323,N_21730,N_20052);
nor U23324 (N_23324,N_21530,N_20550);
nor U23325 (N_23325,N_18839,N_19179);
nand U23326 (N_23326,N_21053,N_20487);
nand U23327 (N_23327,N_21416,N_19646);
and U23328 (N_23328,N_19982,N_21780);
nand U23329 (N_23329,N_20118,N_19377);
xnor U23330 (N_23330,N_21152,N_20659);
nand U23331 (N_23331,N_19291,N_19518);
nor U23332 (N_23332,N_19928,N_19645);
or U23333 (N_23333,N_21551,N_19885);
or U23334 (N_23334,N_19220,N_20022);
or U23335 (N_23335,N_19475,N_20472);
nor U23336 (N_23336,N_18856,N_20129);
and U23337 (N_23337,N_19589,N_19163);
and U23338 (N_23338,N_20727,N_18884);
nor U23339 (N_23339,N_21873,N_21396);
nor U23340 (N_23340,N_20697,N_19392);
and U23341 (N_23341,N_21312,N_19376);
nor U23342 (N_23342,N_20545,N_20159);
nand U23343 (N_23343,N_21655,N_19865);
and U23344 (N_23344,N_20662,N_21091);
or U23345 (N_23345,N_19103,N_19732);
or U23346 (N_23346,N_19673,N_21638);
or U23347 (N_23347,N_20410,N_18754);
nand U23348 (N_23348,N_18905,N_21536);
and U23349 (N_23349,N_20899,N_20350);
nand U23350 (N_23350,N_20615,N_19459);
xnor U23351 (N_23351,N_21502,N_20358);
nor U23352 (N_23352,N_19665,N_20831);
and U23353 (N_23353,N_20686,N_20094);
nor U23354 (N_23354,N_21814,N_19189);
nor U23355 (N_23355,N_20811,N_21348);
nand U23356 (N_23356,N_19887,N_18917);
and U23357 (N_23357,N_19937,N_21315);
nand U23358 (N_23358,N_19980,N_19740);
and U23359 (N_23359,N_19315,N_21082);
and U23360 (N_23360,N_20528,N_19755);
or U23361 (N_23361,N_19824,N_20791);
nor U23362 (N_23362,N_19695,N_21391);
nand U23363 (N_23363,N_20998,N_19670);
nand U23364 (N_23364,N_20065,N_20745);
or U23365 (N_23365,N_19773,N_19942);
or U23366 (N_23366,N_19831,N_18822);
or U23367 (N_23367,N_21448,N_20090);
and U23368 (N_23368,N_20401,N_20025);
nor U23369 (N_23369,N_21190,N_19049);
or U23370 (N_23370,N_19871,N_20816);
nor U23371 (N_23371,N_19077,N_21302);
nand U23372 (N_23372,N_21294,N_21105);
or U23373 (N_23373,N_21674,N_19462);
or U23374 (N_23374,N_19541,N_21114);
and U23375 (N_23375,N_21519,N_21058);
nand U23376 (N_23376,N_19616,N_19440);
and U23377 (N_23377,N_21665,N_21453);
or U23378 (N_23378,N_20189,N_20645);
nor U23379 (N_23379,N_20863,N_20313);
nand U23380 (N_23380,N_21331,N_21083);
or U23381 (N_23381,N_21385,N_19265);
and U23382 (N_23382,N_20463,N_18904);
nand U23383 (N_23383,N_18866,N_19347);
xnor U23384 (N_23384,N_19922,N_21681);
nor U23385 (N_23385,N_20521,N_20658);
or U23386 (N_23386,N_21564,N_21664);
nand U23387 (N_23387,N_21148,N_20669);
and U23388 (N_23388,N_20951,N_21395);
nand U23389 (N_23389,N_21112,N_19517);
or U23390 (N_23390,N_20365,N_21589);
nor U23391 (N_23391,N_20029,N_19607);
nor U23392 (N_23392,N_19886,N_18859);
and U23393 (N_23393,N_21379,N_18946);
xnor U23394 (N_23394,N_18761,N_21871);
nand U23395 (N_23395,N_20741,N_20703);
nand U23396 (N_23396,N_21596,N_21189);
nor U23397 (N_23397,N_21669,N_21106);
or U23398 (N_23398,N_20104,N_19724);
xor U23399 (N_23399,N_20780,N_20557);
and U23400 (N_23400,N_20216,N_21684);
or U23401 (N_23401,N_19538,N_19628);
nand U23402 (N_23402,N_20751,N_20179);
and U23403 (N_23403,N_19707,N_21345);
or U23404 (N_23404,N_21868,N_19881);
xor U23405 (N_23405,N_19733,N_20964);
or U23406 (N_23406,N_18896,N_21233);
or U23407 (N_23407,N_21032,N_20996);
nand U23408 (N_23408,N_20143,N_21010);
and U23409 (N_23409,N_20146,N_20083);
or U23410 (N_23410,N_19435,N_19521);
and U23411 (N_23411,N_20841,N_19181);
xor U23412 (N_23412,N_19890,N_19716);
nor U23413 (N_23413,N_19579,N_19151);
and U23414 (N_23414,N_21816,N_19069);
nand U23415 (N_23415,N_21362,N_21213);
nor U23416 (N_23416,N_19057,N_19786);
or U23417 (N_23417,N_21717,N_21179);
and U23418 (N_23418,N_19264,N_19868);
and U23419 (N_23419,N_19337,N_20310);
nor U23420 (N_23420,N_19413,N_21261);
nand U23421 (N_23421,N_21178,N_20275);
nand U23422 (N_23422,N_20640,N_21123);
xnor U23423 (N_23423,N_20543,N_20224);
and U23424 (N_23424,N_21000,N_20060);
or U23425 (N_23425,N_20190,N_20954);
nand U23426 (N_23426,N_20308,N_21023);
nor U23427 (N_23427,N_20782,N_19621);
xnor U23428 (N_23428,N_19884,N_19879);
nor U23429 (N_23429,N_20499,N_18827);
and U23430 (N_23430,N_21803,N_19295);
nand U23431 (N_23431,N_20978,N_20875);
and U23432 (N_23432,N_19800,N_20079);
nor U23433 (N_23433,N_20575,N_19219);
nor U23434 (N_23434,N_19185,N_21206);
xor U23435 (N_23435,N_19292,N_19105);
and U23436 (N_23436,N_20890,N_21828);
and U23437 (N_23437,N_20530,N_21560);
and U23438 (N_23438,N_20386,N_19020);
nand U23439 (N_23439,N_18947,N_20415);
and U23440 (N_23440,N_20317,N_20679);
nor U23441 (N_23441,N_19170,N_20124);
or U23442 (N_23442,N_20650,N_21066);
nand U23443 (N_23443,N_19639,N_20660);
nor U23444 (N_23444,N_21027,N_21454);
or U23445 (N_23445,N_19317,N_21121);
xnor U23446 (N_23446,N_20334,N_20712);
or U23447 (N_23447,N_19885,N_20325);
or U23448 (N_23448,N_19453,N_19725);
xnor U23449 (N_23449,N_18811,N_21848);
nor U23450 (N_23450,N_19175,N_21450);
or U23451 (N_23451,N_19654,N_20129);
and U23452 (N_23452,N_19788,N_19139);
nor U23453 (N_23453,N_20955,N_20082);
nor U23454 (N_23454,N_19663,N_21704);
and U23455 (N_23455,N_21101,N_21185);
nor U23456 (N_23456,N_20658,N_21710);
and U23457 (N_23457,N_20084,N_19508);
or U23458 (N_23458,N_20135,N_19352);
or U23459 (N_23459,N_20856,N_19146);
nor U23460 (N_23460,N_21775,N_20668);
nor U23461 (N_23461,N_18787,N_21151);
nor U23462 (N_23462,N_20367,N_21162);
xnor U23463 (N_23463,N_19399,N_21153);
and U23464 (N_23464,N_19019,N_20551);
nand U23465 (N_23465,N_21316,N_18818);
and U23466 (N_23466,N_18818,N_20956);
or U23467 (N_23467,N_20717,N_20276);
nor U23468 (N_23468,N_19559,N_19100);
nor U23469 (N_23469,N_19901,N_20322);
and U23470 (N_23470,N_18837,N_21675);
and U23471 (N_23471,N_19965,N_19446);
xor U23472 (N_23472,N_21604,N_20276);
xor U23473 (N_23473,N_20315,N_21525);
nand U23474 (N_23474,N_20907,N_20856);
nand U23475 (N_23475,N_19421,N_20528);
and U23476 (N_23476,N_18752,N_19387);
and U23477 (N_23477,N_21598,N_19498);
nand U23478 (N_23478,N_19806,N_18896);
xnor U23479 (N_23479,N_19371,N_20245);
nor U23480 (N_23480,N_20607,N_21405);
nand U23481 (N_23481,N_19119,N_21147);
or U23482 (N_23482,N_21590,N_19928);
and U23483 (N_23483,N_20270,N_19549);
xor U23484 (N_23484,N_21569,N_20065);
nand U23485 (N_23485,N_19875,N_20298);
nor U23486 (N_23486,N_19288,N_21106);
nand U23487 (N_23487,N_20761,N_21582);
nand U23488 (N_23488,N_19228,N_20277);
xor U23489 (N_23489,N_21313,N_21739);
nand U23490 (N_23490,N_19340,N_19739);
nor U23491 (N_23491,N_21694,N_18758);
nor U23492 (N_23492,N_20711,N_21535);
nor U23493 (N_23493,N_21817,N_19191);
or U23494 (N_23494,N_19581,N_20065);
and U23495 (N_23495,N_20241,N_21211);
and U23496 (N_23496,N_18804,N_20568);
nor U23497 (N_23497,N_21595,N_20700);
nand U23498 (N_23498,N_18765,N_20688);
nand U23499 (N_23499,N_19234,N_19015);
and U23500 (N_23500,N_19022,N_21634);
xor U23501 (N_23501,N_19167,N_20913);
xor U23502 (N_23502,N_21628,N_21699);
nand U23503 (N_23503,N_20194,N_21568);
or U23504 (N_23504,N_19975,N_20604);
nand U23505 (N_23505,N_19432,N_19859);
and U23506 (N_23506,N_20831,N_19035);
nor U23507 (N_23507,N_19594,N_19694);
or U23508 (N_23508,N_20441,N_21718);
or U23509 (N_23509,N_19915,N_21359);
nor U23510 (N_23510,N_20126,N_19641);
nor U23511 (N_23511,N_20718,N_19152);
and U23512 (N_23512,N_21622,N_21308);
or U23513 (N_23513,N_20089,N_19890);
xor U23514 (N_23514,N_19104,N_18795);
nand U23515 (N_23515,N_20039,N_19237);
or U23516 (N_23516,N_21805,N_19262);
and U23517 (N_23517,N_19959,N_20362);
nand U23518 (N_23518,N_18914,N_21660);
nor U23519 (N_23519,N_19283,N_21056);
nor U23520 (N_23520,N_19573,N_18830);
or U23521 (N_23521,N_20518,N_21699);
and U23522 (N_23522,N_20594,N_20853);
nor U23523 (N_23523,N_18847,N_21133);
or U23524 (N_23524,N_19109,N_18939);
nand U23525 (N_23525,N_20141,N_21175);
nor U23526 (N_23526,N_18868,N_19359);
xnor U23527 (N_23527,N_21476,N_20077);
or U23528 (N_23528,N_19830,N_19920);
or U23529 (N_23529,N_20376,N_20009);
and U23530 (N_23530,N_19552,N_20810);
nor U23531 (N_23531,N_20504,N_20467);
nor U23532 (N_23532,N_21231,N_19342);
or U23533 (N_23533,N_20461,N_19179);
nor U23534 (N_23534,N_19215,N_19465);
and U23535 (N_23535,N_20269,N_20530);
or U23536 (N_23536,N_21413,N_18949);
and U23537 (N_23537,N_20979,N_21806);
or U23538 (N_23538,N_21631,N_20845);
or U23539 (N_23539,N_20273,N_18851);
or U23540 (N_23540,N_20111,N_20769);
nand U23541 (N_23541,N_19217,N_19895);
xnor U23542 (N_23542,N_19678,N_20751);
nand U23543 (N_23543,N_19686,N_20061);
xnor U23544 (N_23544,N_20177,N_20990);
nor U23545 (N_23545,N_19604,N_21422);
nand U23546 (N_23546,N_21517,N_19507);
nor U23547 (N_23547,N_18840,N_19625);
nor U23548 (N_23548,N_20045,N_18998);
nor U23549 (N_23549,N_21566,N_20840);
and U23550 (N_23550,N_21385,N_20876);
and U23551 (N_23551,N_21716,N_21815);
and U23552 (N_23552,N_21820,N_19423);
and U23553 (N_23553,N_19216,N_21583);
nor U23554 (N_23554,N_19488,N_20685);
or U23555 (N_23555,N_19760,N_21516);
and U23556 (N_23556,N_19474,N_19059);
and U23557 (N_23557,N_19847,N_20319);
and U23558 (N_23558,N_18918,N_19096);
nor U23559 (N_23559,N_19990,N_21053);
xor U23560 (N_23560,N_20264,N_19636);
and U23561 (N_23561,N_19271,N_20833);
or U23562 (N_23562,N_20779,N_21251);
xnor U23563 (N_23563,N_20762,N_19529);
nand U23564 (N_23564,N_19099,N_19544);
or U23565 (N_23565,N_19380,N_18825);
or U23566 (N_23566,N_21836,N_20949);
nor U23567 (N_23567,N_21676,N_19944);
nand U23568 (N_23568,N_19618,N_21127);
and U23569 (N_23569,N_20156,N_20670);
or U23570 (N_23570,N_19599,N_20256);
nor U23571 (N_23571,N_19613,N_19598);
xor U23572 (N_23572,N_19691,N_19386);
nand U23573 (N_23573,N_19916,N_21578);
nand U23574 (N_23574,N_21853,N_20585);
and U23575 (N_23575,N_21848,N_20484);
nor U23576 (N_23576,N_21007,N_19070);
nor U23577 (N_23577,N_20141,N_19151);
nand U23578 (N_23578,N_21631,N_21042);
nand U23579 (N_23579,N_19158,N_20671);
nand U23580 (N_23580,N_21518,N_19491);
nand U23581 (N_23581,N_20964,N_19877);
or U23582 (N_23582,N_20630,N_19404);
xor U23583 (N_23583,N_21447,N_19249);
nor U23584 (N_23584,N_20548,N_21787);
xor U23585 (N_23585,N_20711,N_19078);
nand U23586 (N_23586,N_20348,N_21413);
nand U23587 (N_23587,N_21404,N_19562);
and U23588 (N_23588,N_21679,N_18860);
and U23589 (N_23589,N_19549,N_20330);
and U23590 (N_23590,N_21802,N_20730);
and U23591 (N_23591,N_20648,N_19539);
nand U23592 (N_23592,N_20735,N_19487);
nand U23593 (N_23593,N_21683,N_18936);
nor U23594 (N_23594,N_20225,N_21016);
nand U23595 (N_23595,N_18847,N_19540);
nand U23596 (N_23596,N_20224,N_19510);
nand U23597 (N_23597,N_19881,N_20783);
and U23598 (N_23598,N_19447,N_19781);
or U23599 (N_23599,N_21364,N_19946);
nor U23600 (N_23600,N_19763,N_20627);
and U23601 (N_23601,N_20034,N_20092);
nand U23602 (N_23602,N_20160,N_21865);
nor U23603 (N_23603,N_21663,N_18973);
and U23604 (N_23604,N_20212,N_21130);
and U23605 (N_23605,N_21255,N_20982);
and U23606 (N_23606,N_19607,N_20636);
nand U23607 (N_23607,N_20703,N_20861);
or U23608 (N_23608,N_20795,N_19641);
nand U23609 (N_23609,N_20159,N_19284);
or U23610 (N_23610,N_19912,N_21190);
nand U23611 (N_23611,N_21648,N_20703);
xnor U23612 (N_23612,N_19482,N_21124);
nor U23613 (N_23613,N_19674,N_19815);
nand U23614 (N_23614,N_20935,N_21054);
nor U23615 (N_23615,N_19875,N_21768);
or U23616 (N_23616,N_21136,N_19632);
or U23617 (N_23617,N_20342,N_21023);
nand U23618 (N_23618,N_18993,N_19386);
nor U23619 (N_23619,N_19432,N_21079);
and U23620 (N_23620,N_20549,N_19552);
or U23621 (N_23621,N_21143,N_20656);
nand U23622 (N_23622,N_21849,N_19122);
xnor U23623 (N_23623,N_19882,N_19173);
xnor U23624 (N_23624,N_21581,N_21428);
nand U23625 (N_23625,N_21416,N_21159);
or U23626 (N_23626,N_19467,N_19595);
nand U23627 (N_23627,N_19252,N_21414);
xnor U23628 (N_23628,N_19832,N_19631);
and U23629 (N_23629,N_21432,N_20387);
or U23630 (N_23630,N_19016,N_20211);
nor U23631 (N_23631,N_19374,N_21619);
or U23632 (N_23632,N_18895,N_21238);
nor U23633 (N_23633,N_19165,N_20186);
and U23634 (N_23634,N_19221,N_19176);
and U23635 (N_23635,N_20444,N_21568);
and U23636 (N_23636,N_20643,N_19283);
nor U23637 (N_23637,N_20267,N_21724);
xnor U23638 (N_23638,N_19804,N_20146);
nand U23639 (N_23639,N_20927,N_21337);
nor U23640 (N_23640,N_20450,N_21817);
or U23641 (N_23641,N_21654,N_20932);
and U23642 (N_23642,N_21381,N_19393);
nor U23643 (N_23643,N_19583,N_20195);
and U23644 (N_23644,N_20652,N_20641);
or U23645 (N_23645,N_21632,N_21801);
and U23646 (N_23646,N_20123,N_19331);
and U23647 (N_23647,N_19593,N_18899);
or U23648 (N_23648,N_20041,N_19005);
and U23649 (N_23649,N_21270,N_20954);
nor U23650 (N_23650,N_20459,N_20541);
or U23651 (N_23651,N_21696,N_20364);
nor U23652 (N_23652,N_21424,N_19076);
nor U23653 (N_23653,N_19102,N_20705);
and U23654 (N_23654,N_20017,N_21754);
and U23655 (N_23655,N_19577,N_19279);
nor U23656 (N_23656,N_20134,N_21420);
nor U23657 (N_23657,N_21283,N_20939);
and U23658 (N_23658,N_19576,N_20734);
nor U23659 (N_23659,N_20631,N_19169);
nand U23660 (N_23660,N_19958,N_21840);
and U23661 (N_23661,N_19042,N_20385);
nor U23662 (N_23662,N_20054,N_20592);
nand U23663 (N_23663,N_20230,N_20481);
xor U23664 (N_23664,N_20600,N_18993);
or U23665 (N_23665,N_19700,N_19693);
nor U23666 (N_23666,N_20539,N_20331);
or U23667 (N_23667,N_19986,N_19834);
nand U23668 (N_23668,N_20468,N_20401);
or U23669 (N_23669,N_21807,N_19502);
xnor U23670 (N_23670,N_21254,N_20539);
or U23671 (N_23671,N_20873,N_20393);
and U23672 (N_23672,N_18928,N_19816);
and U23673 (N_23673,N_19751,N_19528);
or U23674 (N_23674,N_20219,N_19141);
nor U23675 (N_23675,N_20478,N_21386);
or U23676 (N_23676,N_21403,N_20981);
or U23677 (N_23677,N_18862,N_19456);
nand U23678 (N_23678,N_21042,N_19737);
nand U23679 (N_23679,N_20507,N_21752);
nand U23680 (N_23680,N_21391,N_20220);
nor U23681 (N_23681,N_21258,N_19564);
nand U23682 (N_23682,N_21862,N_19082);
nand U23683 (N_23683,N_21386,N_20836);
or U23684 (N_23684,N_18941,N_19565);
or U23685 (N_23685,N_20486,N_19957);
or U23686 (N_23686,N_18752,N_21558);
nor U23687 (N_23687,N_21376,N_21165);
and U23688 (N_23688,N_18770,N_18801);
xor U23689 (N_23689,N_19715,N_19992);
nand U23690 (N_23690,N_21354,N_19347);
nand U23691 (N_23691,N_19219,N_21632);
and U23692 (N_23692,N_20070,N_19535);
xor U23693 (N_23693,N_20467,N_21182);
nor U23694 (N_23694,N_18828,N_19971);
nand U23695 (N_23695,N_21273,N_21563);
nor U23696 (N_23696,N_18970,N_21390);
nor U23697 (N_23697,N_19661,N_20069);
xor U23698 (N_23698,N_20623,N_21792);
nand U23699 (N_23699,N_20559,N_20677);
or U23700 (N_23700,N_20437,N_19348);
xnor U23701 (N_23701,N_18871,N_18863);
nand U23702 (N_23702,N_19089,N_21859);
nor U23703 (N_23703,N_21856,N_20530);
nor U23704 (N_23704,N_21733,N_20101);
xor U23705 (N_23705,N_20995,N_20273);
and U23706 (N_23706,N_21380,N_21772);
nor U23707 (N_23707,N_21803,N_19474);
and U23708 (N_23708,N_21870,N_20264);
nor U23709 (N_23709,N_19594,N_18794);
nor U23710 (N_23710,N_20622,N_21364);
or U23711 (N_23711,N_20959,N_18840);
or U23712 (N_23712,N_20793,N_18811);
nand U23713 (N_23713,N_21371,N_21786);
and U23714 (N_23714,N_21769,N_19396);
and U23715 (N_23715,N_19295,N_19692);
and U23716 (N_23716,N_20230,N_20073);
nand U23717 (N_23717,N_18754,N_20826);
or U23718 (N_23718,N_21686,N_18780);
nand U23719 (N_23719,N_19486,N_21395);
and U23720 (N_23720,N_20473,N_20437);
nor U23721 (N_23721,N_19101,N_19078);
nor U23722 (N_23722,N_21008,N_19050);
and U23723 (N_23723,N_19779,N_21552);
xnor U23724 (N_23724,N_20642,N_21785);
nor U23725 (N_23725,N_21291,N_20445);
and U23726 (N_23726,N_19967,N_20682);
nand U23727 (N_23727,N_19983,N_21073);
xor U23728 (N_23728,N_20237,N_19401);
xnor U23729 (N_23729,N_20593,N_20920);
and U23730 (N_23730,N_19731,N_19614);
nor U23731 (N_23731,N_21390,N_19306);
nor U23732 (N_23732,N_21054,N_20780);
nor U23733 (N_23733,N_19516,N_20588);
nor U23734 (N_23734,N_19387,N_19002);
nand U23735 (N_23735,N_20423,N_19080);
or U23736 (N_23736,N_21401,N_21566);
and U23737 (N_23737,N_20374,N_19249);
or U23738 (N_23738,N_19532,N_20985);
or U23739 (N_23739,N_20195,N_20920);
nand U23740 (N_23740,N_19444,N_19595);
nor U23741 (N_23741,N_19463,N_19918);
nand U23742 (N_23742,N_21034,N_19489);
or U23743 (N_23743,N_20563,N_21371);
nand U23744 (N_23744,N_21744,N_19310);
nor U23745 (N_23745,N_21439,N_19601);
xnor U23746 (N_23746,N_21553,N_19428);
nor U23747 (N_23747,N_18848,N_19027);
and U23748 (N_23748,N_21410,N_21393);
nor U23749 (N_23749,N_18879,N_19702);
and U23750 (N_23750,N_20694,N_20328);
nor U23751 (N_23751,N_19675,N_20420);
nand U23752 (N_23752,N_21462,N_21540);
nor U23753 (N_23753,N_18835,N_20269);
or U23754 (N_23754,N_19915,N_20968);
nor U23755 (N_23755,N_21779,N_20555);
and U23756 (N_23756,N_19701,N_18937);
and U23757 (N_23757,N_19375,N_19514);
or U23758 (N_23758,N_19655,N_19735);
or U23759 (N_23759,N_18767,N_21245);
nor U23760 (N_23760,N_20354,N_18799);
nor U23761 (N_23761,N_20163,N_20992);
nor U23762 (N_23762,N_20461,N_20763);
and U23763 (N_23763,N_19786,N_19579);
and U23764 (N_23764,N_20826,N_20528);
or U23765 (N_23765,N_20496,N_20269);
nor U23766 (N_23766,N_21635,N_21761);
nand U23767 (N_23767,N_20918,N_21737);
and U23768 (N_23768,N_21778,N_21012);
nor U23769 (N_23769,N_20002,N_21540);
nand U23770 (N_23770,N_21252,N_19520);
xor U23771 (N_23771,N_19929,N_20464);
nand U23772 (N_23772,N_19902,N_20354);
or U23773 (N_23773,N_20593,N_21436);
nand U23774 (N_23774,N_19863,N_20216);
xnor U23775 (N_23775,N_20862,N_19595);
or U23776 (N_23776,N_20120,N_20024);
or U23777 (N_23777,N_20964,N_18834);
and U23778 (N_23778,N_20448,N_20724);
nor U23779 (N_23779,N_19200,N_20010);
nor U23780 (N_23780,N_20132,N_19601);
or U23781 (N_23781,N_18780,N_21752);
and U23782 (N_23782,N_20975,N_20665);
and U23783 (N_23783,N_20178,N_21209);
and U23784 (N_23784,N_21384,N_18985);
nand U23785 (N_23785,N_19011,N_21737);
nor U23786 (N_23786,N_19966,N_18890);
nand U23787 (N_23787,N_20845,N_19744);
or U23788 (N_23788,N_19535,N_20245);
or U23789 (N_23789,N_19056,N_19785);
or U23790 (N_23790,N_20527,N_20358);
nand U23791 (N_23791,N_21600,N_18786);
or U23792 (N_23792,N_20068,N_20818);
nor U23793 (N_23793,N_20351,N_20182);
nor U23794 (N_23794,N_20252,N_20680);
nand U23795 (N_23795,N_20476,N_21403);
nor U23796 (N_23796,N_19962,N_19948);
nand U23797 (N_23797,N_19715,N_21479);
nor U23798 (N_23798,N_19081,N_20637);
and U23799 (N_23799,N_19802,N_18810);
nor U23800 (N_23800,N_21371,N_19337);
or U23801 (N_23801,N_20975,N_19683);
and U23802 (N_23802,N_20724,N_20646);
or U23803 (N_23803,N_21731,N_18759);
nor U23804 (N_23804,N_20836,N_21329);
nor U23805 (N_23805,N_20475,N_21016);
and U23806 (N_23806,N_21054,N_21559);
nor U23807 (N_23807,N_19937,N_18752);
or U23808 (N_23808,N_19987,N_18905);
and U23809 (N_23809,N_20671,N_19635);
xnor U23810 (N_23810,N_21630,N_18788);
and U23811 (N_23811,N_21297,N_19973);
or U23812 (N_23812,N_21850,N_20190);
or U23813 (N_23813,N_21623,N_19035);
nor U23814 (N_23814,N_21147,N_20136);
nand U23815 (N_23815,N_20590,N_21251);
nand U23816 (N_23816,N_20066,N_20804);
nor U23817 (N_23817,N_19058,N_21313);
and U23818 (N_23818,N_20060,N_20124);
nor U23819 (N_23819,N_18991,N_19958);
and U23820 (N_23820,N_19140,N_20115);
or U23821 (N_23821,N_19774,N_19582);
nand U23822 (N_23822,N_21350,N_21396);
or U23823 (N_23823,N_20842,N_19191);
xor U23824 (N_23824,N_20790,N_20805);
nor U23825 (N_23825,N_19206,N_20169);
xnor U23826 (N_23826,N_21135,N_20771);
and U23827 (N_23827,N_19574,N_19503);
nand U23828 (N_23828,N_20192,N_19993);
nand U23829 (N_23829,N_19204,N_20779);
and U23830 (N_23830,N_21642,N_18928);
nor U23831 (N_23831,N_20364,N_20531);
nor U23832 (N_23832,N_19371,N_19480);
nor U23833 (N_23833,N_20019,N_21405);
and U23834 (N_23834,N_19284,N_19293);
xor U23835 (N_23835,N_19271,N_21467);
and U23836 (N_23836,N_19736,N_19478);
and U23837 (N_23837,N_20213,N_19178);
nand U23838 (N_23838,N_20811,N_20631);
nor U23839 (N_23839,N_21382,N_21677);
nand U23840 (N_23840,N_20918,N_20741);
nor U23841 (N_23841,N_19861,N_21459);
nor U23842 (N_23842,N_19707,N_20430);
xor U23843 (N_23843,N_19753,N_19297);
or U23844 (N_23844,N_20632,N_21138);
nand U23845 (N_23845,N_21000,N_19974);
and U23846 (N_23846,N_19250,N_21593);
nor U23847 (N_23847,N_20433,N_19308);
nor U23848 (N_23848,N_20903,N_19020);
nand U23849 (N_23849,N_18812,N_19240);
and U23850 (N_23850,N_19061,N_20832);
nand U23851 (N_23851,N_19965,N_20296);
xnor U23852 (N_23852,N_19780,N_20359);
nor U23853 (N_23853,N_19567,N_18751);
or U23854 (N_23854,N_20998,N_19861);
or U23855 (N_23855,N_19016,N_19455);
nor U23856 (N_23856,N_19820,N_21535);
nand U23857 (N_23857,N_21753,N_20115);
nor U23858 (N_23858,N_19951,N_21092);
xnor U23859 (N_23859,N_19561,N_19269);
or U23860 (N_23860,N_19164,N_18870);
nor U23861 (N_23861,N_19615,N_21550);
nand U23862 (N_23862,N_21148,N_19362);
and U23863 (N_23863,N_20352,N_19226);
nand U23864 (N_23864,N_20376,N_19401);
or U23865 (N_23865,N_20751,N_20225);
nand U23866 (N_23866,N_19861,N_20699);
nor U23867 (N_23867,N_18909,N_19241);
nor U23868 (N_23868,N_20386,N_18915);
and U23869 (N_23869,N_20962,N_19857);
nor U23870 (N_23870,N_20537,N_21602);
nand U23871 (N_23871,N_19666,N_20935);
nor U23872 (N_23872,N_20213,N_20416);
or U23873 (N_23873,N_20319,N_18932);
nor U23874 (N_23874,N_21849,N_20483);
nand U23875 (N_23875,N_19367,N_20609);
nor U23876 (N_23876,N_21036,N_21840);
or U23877 (N_23877,N_19873,N_21699);
xnor U23878 (N_23878,N_20823,N_21737);
or U23879 (N_23879,N_21506,N_21416);
xor U23880 (N_23880,N_21485,N_20732);
nor U23881 (N_23881,N_19593,N_19681);
or U23882 (N_23882,N_20213,N_18760);
or U23883 (N_23883,N_19912,N_20194);
nand U23884 (N_23884,N_20648,N_21685);
nand U23885 (N_23885,N_18776,N_19062);
xnor U23886 (N_23886,N_21157,N_20625);
nand U23887 (N_23887,N_20755,N_19303);
nand U23888 (N_23888,N_19757,N_21189);
nand U23889 (N_23889,N_20951,N_19181);
or U23890 (N_23890,N_20620,N_19203);
nor U23891 (N_23891,N_21638,N_19708);
or U23892 (N_23892,N_20136,N_21831);
nor U23893 (N_23893,N_21792,N_21560);
nor U23894 (N_23894,N_21103,N_21848);
nor U23895 (N_23895,N_20523,N_19200);
and U23896 (N_23896,N_19407,N_21278);
nor U23897 (N_23897,N_21647,N_21737);
nand U23898 (N_23898,N_19393,N_21357);
and U23899 (N_23899,N_20132,N_20028);
and U23900 (N_23900,N_20027,N_19328);
nor U23901 (N_23901,N_20951,N_20826);
nor U23902 (N_23902,N_18873,N_18893);
nor U23903 (N_23903,N_18979,N_21262);
or U23904 (N_23904,N_21833,N_19471);
nor U23905 (N_23905,N_20795,N_19110);
nand U23906 (N_23906,N_20854,N_21078);
nand U23907 (N_23907,N_19346,N_20864);
and U23908 (N_23908,N_19812,N_21832);
or U23909 (N_23909,N_20385,N_20944);
and U23910 (N_23910,N_20888,N_20686);
and U23911 (N_23911,N_19204,N_19818);
nand U23912 (N_23912,N_20009,N_20062);
or U23913 (N_23913,N_19122,N_19119);
nor U23914 (N_23914,N_21678,N_20926);
nand U23915 (N_23915,N_19327,N_21353);
nand U23916 (N_23916,N_21869,N_20936);
and U23917 (N_23917,N_19464,N_20462);
or U23918 (N_23918,N_20700,N_19223);
nand U23919 (N_23919,N_21054,N_18819);
and U23920 (N_23920,N_18883,N_20959);
nand U23921 (N_23921,N_19319,N_21727);
xnor U23922 (N_23922,N_21669,N_19040);
and U23923 (N_23923,N_21174,N_19275);
nor U23924 (N_23924,N_21429,N_20752);
xor U23925 (N_23925,N_19061,N_19835);
and U23926 (N_23926,N_20361,N_20699);
nor U23927 (N_23927,N_21211,N_19391);
and U23928 (N_23928,N_20287,N_19184);
and U23929 (N_23929,N_20706,N_21695);
nor U23930 (N_23930,N_21013,N_21689);
or U23931 (N_23931,N_19625,N_20798);
and U23932 (N_23932,N_21485,N_18924);
nor U23933 (N_23933,N_19795,N_20176);
and U23934 (N_23934,N_20259,N_19658);
nand U23935 (N_23935,N_20893,N_21815);
nand U23936 (N_23936,N_20665,N_21379);
nor U23937 (N_23937,N_18969,N_19244);
nand U23938 (N_23938,N_20105,N_20999);
or U23939 (N_23939,N_19598,N_19673);
nand U23940 (N_23940,N_20668,N_20446);
nand U23941 (N_23941,N_20387,N_20536);
nand U23942 (N_23942,N_19036,N_19166);
or U23943 (N_23943,N_21779,N_21023);
nor U23944 (N_23944,N_21658,N_20902);
nand U23945 (N_23945,N_19701,N_18845);
and U23946 (N_23946,N_20894,N_21181);
or U23947 (N_23947,N_20473,N_19967);
nor U23948 (N_23948,N_21351,N_20068);
and U23949 (N_23949,N_21632,N_18944);
nand U23950 (N_23950,N_19640,N_19334);
nor U23951 (N_23951,N_20056,N_21807);
nor U23952 (N_23952,N_21412,N_18809);
nand U23953 (N_23953,N_18832,N_21753);
nand U23954 (N_23954,N_20587,N_20047);
or U23955 (N_23955,N_21072,N_18993);
nand U23956 (N_23956,N_18823,N_20868);
and U23957 (N_23957,N_19723,N_19057);
nor U23958 (N_23958,N_20541,N_20246);
nor U23959 (N_23959,N_19722,N_20042);
xor U23960 (N_23960,N_19567,N_20114);
xor U23961 (N_23961,N_20992,N_20072);
nor U23962 (N_23962,N_21702,N_18973);
or U23963 (N_23963,N_19559,N_19343);
nand U23964 (N_23964,N_20707,N_20295);
nor U23965 (N_23965,N_19407,N_20561);
or U23966 (N_23966,N_18796,N_18913);
nand U23967 (N_23967,N_20613,N_19330);
nor U23968 (N_23968,N_19149,N_20350);
and U23969 (N_23969,N_19644,N_21591);
or U23970 (N_23970,N_20491,N_19506);
or U23971 (N_23971,N_20179,N_19963);
nor U23972 (N_23972,N_20906,N_20324);
or U23973 (N_23973,N_20649,N_19038);
nor U23974 (N_23974,N_21297,N_19751);
nor U23975 (N_23975,N_21000,N_19664);
and U23976 (N_23976,N_19549,N_19301);
xnor U23977 (N_23977,N_20361,N_19775);
and U23978 (N_23978,N_19993,N_21630);
or U23979 (N_23979,N_21177,N_19484);
nand U23980 (N_23980,N_20796,N_20817);
and U23981 (N_23981,N_20458,N_20996);
or U23982 (N_23982,N_19673,N_18869);
or U23983 (N_23983,N_20501,N_19882);
nor U23984 (N_23984,N_21405,N_19578);
and U23985 (N_23985,N_21084,N_19374);
or U23986 (N_23986,N_19409,N_20732);
or U23987 (N_23987,N_18824,N_19338);
or U23988 (N_23988,N_20552,N_21521);
and U23989 (N_23989,N_20191,N_20668);
and U23990 (N_23990,N_21340,N_20211);
nor U23991 (N_23991,N_21615,N_21167);
and U23992 (N_23992,N_20074,N_21167);
or U23993 (N_23993,N_20439,N_20072);
and U23994 (N_23994,N_18799,N_19278);
nor U23995 (N_23995,N_21432,N_19872);
and U23996 (N_23996,N_19095,N_21336);
nor U23997 (N_23997,N_20973,N_21060);
and U23998 (N_23998,N_20881,N_20950);
and U23999 (N_23999,N_19067,N_21765);
and U24000 (N_24000,N_20634,N_21453);
nor U24001 (N_24001,N_21779,N_19617);
and U24002 (N_24002,N_19857,N_21215);
nand U24003 (N_24003,N_21210,N_20769);
nor U24004 (N_24004,N_19175,N_21334);
nor U24005 (N_24005,N_19982,N_18989);
or U24006 (N_24006,N_18973,N_19223);
xor U24007 (N_24007,N_18869,N_20164);
or U24008 (N_24008,N_20292,N_21217);
xor U24009 (N_24009,N_20988,N_21655);
nand U24010 (N_24010,N_21213,N_21365);
or U24011 (N_24011,N_19663,N_21020);
nand U24012 (N_24012,N_18792,N_19123);
or U24013 (N_24013,N_21306,N_20974);
or U24014 (N_24014,N_20877,N_19137);
xor U24015 (N_24015,N_20917,N_20562);
xnor U24016 (N_24016,N_21311,N_18807);
nor U24017 (N_24017,N_20373,N_19978);
or U24018 (N_24018,N_19206,N_20059);
and U24019 (N_24019,N_19471,N_19308);
nor U24020 (N_24020,N_21577,N_21556);
nor U24021 (N_24021,N_21036,N_20653);
nor U24022 (N_24022,N_19641,N_20055);
and U24023 (N_24023,N_19952,N_20834);
xor U24024 (N_24024,N_18884,N_21591);
xnor U24025 (N_24025,N_18949,N_20665);
xor U24026 (N_24026,N_19756,N_19257);
nand U24027 (N_24027,N_19539,N_21367);
nor U24028 (N_24028,N_18841,N_18923);
or U24029 (N_24029,N_19692,N_19763);
and U24030 (N_24030,N_18991,N_20655);
xnor U24031 (N_24031,N_20458,N_18751);
or U24032 (N_24032,N_21014,N_20774);
and U24033 (N_24033,N_21532,N_21190);
and U24034 (N_24034,N_21255,N_18849);
xnor U24035 (N_24035,N_20984,N_19627);
and U24036 (N_24036,N_21632,N_19716);
nand U24037 (N_24037,N_20902,N_21289);
and U24038 (N_24038,N_20650,N_21451);
or U24039 (N_24039,N_19027,N_19622);
xor U24040 (N_24040,N_21747,N_21576);
or U24041 (N_24041,N_20790,N_19446);
nor U24042 (N_24042,N_19950,N_19100);
nand U24043 (N_24043,N_20721,N_20888);
xor U24044 (N_24044,N_20852,N_20967);
and U24045 (N_24045,N_20814,N_20050);
and U24046 (N_24046,N_20646,N_19353);
nand U24047 (N_24047,N_21297,N_19536);
and U24048 (N_24048,N_18782,N_21169);
xnor U24049 (N_24049,N_19495,N_20402);
and U24050 (N_24050,N_21290,N_18993);
nand U24051 (N_24051,N_19430,N_20621);
and U24052 (N_24052,N_21664,N_19887);
nand U24053 (N_24053,N_20052,N_21276);
nand U24054 (N_24054,N_19614,N_21075);
or U24055 (N_24055,N_21664,N_20946);
nor U24056 (N_24056,N_21220,N_20836);
and U24057 (N_24057,N_20662,N_19127);
nand U24058 (N_24058,N_21459,N_20943);
or U24059 (N_24059,N_18969,N_19308);
nor U24060 (N_24060,N_20354,N_21856);
nand U24061 (N_24061,N_21069,N_19793);
or U24062 (N_24062,N_19864,N_19780);
xor U24063 (N_24063,N_21208,N_20537);
and U24064 (N_24064,N_21218,N_20552);
nand U24065 (N_24065,N_19505,N_21377);
and U24066 (N_24066,N_20003,N_19238);
or U24067 (N_24067,N_19271,N_20455);
nor U24068 (N_24068,N_21041,N_19602);
nor U24069 (N_24069,N_19674,N_20710);
and U24070 (N_24070,N_19527,N_19874);
and U24071 (N_24071,N_21837,N_19876);
and U24072 (N_24072,N_21543,N_19111);
nor U24073 (N_24073,N_19505,N_21719);
and U24074 (N_24074,N_21362,N_19828);
nand U24075 (N_24075,N_19103,N_21804);
and U24076 (N_24076,N_20852,N_20486);
and U24077 (N_24077,N_21621,N_19539);
and U24078 (N_24078,N_21210,N_18762);
or U24079 (N_24079,N_19798,N_19004);
or U24080 (N_24080,N_18960,N_19171);
and U24081 (N_24081,N_19403,N_20905);
nor U24082 (N_24082,N_21407,N_21729);
and U24083 (N_24083,N_21440,N_19557);
and U24084 (N_24084,N_20345,N_19619);
nand U24085 (N_24085,N_21045,N_20185);
or U24086 (N_24086,N_21859,N_18993);
or U24087 (N_24087,N_19148,N_21706);
or U24088 (N_24088,N_19199,N_20431);
or U24089 (N_24089,N_20845,N_20125);
or U24090 (N_24090,N_21766,N_19873);
nand U24091 (N_24091,N_20671,N_21309);
and U24092 (N_24092,N_19700,N_21779);
or U24093 (N_24093,N_20952,N_20148);
and U24094 (N_24094,N_21568,N_18757);
nand U24095 (N_24095,N_20449,N_18904);
or U24096 (N_24096,N_20602,N_21436);
xor U24097 (N_24097,N_20090,N_20056);
nand U24098 (N_24098,N_19057,N_20567);
nand U24099 (N_24099,N_18818,N_20866);
and U24100 (N_24100,N_19976,N_19514);
and U24101 (N_24101,N_18833,N_18927);
or U24102 (N_24102,N_19792,N_21598);
nor U24103 (N_24103,N_19743,N_19704);
or U24104 (N_24104,N_21751,N_19126);
nor U24105 (N_24105,N_20406,N_19515);
nor U24106 (N_24106,N_21532,N_19602);
or U24107 (N_24107,N_19340,N_19899);
or U24108 (N_24108,N_19957,N_21041);
xnor U24109 (N_24109,N_21838,N_21220);
nor U24110 (N_24110,N_20502,N_20120);
nand U24111 (N_24111,N_21298,N_19624);
nor U24112 (N_24112,N_20071,N_21077);
nor U24113 (N_24113,N_20493,N_20122);
xor U24114 (N_24114,N_21759,N_19297);
xnor U24115 (N_24115,N_19529,N_18767);
xor U24116 (N_24116,N_20333,N_19596);
or U24117 (N_24117,N_21238,N_19008);
nand U24118 (N_24118,N_21756,N_19867);
nor U24119 (N_24119,N_20381,N_20179);
and U24120 (N_24120,N_21541,N_20307);
nand U24121 (N_24121,N_20100,N_20855);
or U24122 (N_24122,N_19300,N_19481);
nor U24123 (N_24123,N_20758,N_21525);
nor U24124 (N_24124,N_18930,N_20557);
or U24125 (N_24125,N_21679,N_21217);
nor U24126 (N_24126,N_19071,N_21827);
and U24127 (N_24127,N_21672,N_21814);
and U24128 (N_24128,N_20916,N_19068);
nor U24129 (N_24129,N_21595,N_20635);
or U24130 (N_24130,N_21703,N_20857);
nor U24131 (N_24131,N_21094,N_21480);
nand U24132 (N_24132,N_19052,N_21457);
nand U24133 (N_24133,N_20396,N_21801);
nand U24134 (N_24134,N_20283,N_21468);
nand U24135 (N_24135,N_21846,N_21369);
xnor U24136 (N_24136,N_20332,N_19390);
nand U24137 (N_24137,N_20225,N_21827);
or U24138 (N_24138,N_21686,N_21335);
and U24139 (N_24139,N_20667,N_21872);
nor U24140 (N_24140,N_20839,N_19916);
or U24141 (N_24141,N_20831,N_19774);
nand U24142 (N_24142,N_18809,N_20653);
xnor U24143 (N_24143,N_18921,N_20484);
xnor U24144 (N_24144,N_19525,N_20272);
and U24145 (N_24145,N_18912,N_20926);
nand U24146 (N_24146,N_21418,N_19477);
or U24147 (N_24147,N_19049,N_20108);
nor U24148 (N_24148,N_20576,N_20374);
nand U24149 (N_24149,N_21024,N_20971);
xnor U24150 (N_24150,N_21274,N_19075);
or U24151 (N_24151,N_21756,N_19403);
nor U24152 (N_24152,N_18851,N_20693);
nor U24153 (N_24153,N_19416,N_21480);
and U24154 (N_24154,N_20203,N_21163);
nand U24155 (N_24155,N_21423,N_19422);
nand U24156 (N_24156,N_19216,N_19495);
or U24157 (N_24157,N_19866,N_21561);
xor U24158 (N_24158,N_19405,N_21312);
and U24159 (N_24159,N_21240,N_21552);
xnor U24160 (N_24160,N_20013,N_20899);
nor U24161 (N_24161,N_20028,N_19938);
xor U24162 (N_24162,N_20321,N_20842);
nand U24163 (N_24163,N_20321,N_20658);
or U24164 (N_24164,N_21116,N_19253);
and U24165 (N_24165,N_20599,N_20134);
nor U24166 (N_24166,N_21069,N_19720);
xor U24167 (N_24167,N_19699,N_21505);
and U24168 (N_24168,N_18830,N_18777);
and U24169 (N_24169,N_21605,N_18771);
xor U24170 (N_24170,N_21627,N_20684);
and U24171 (N_24171,N_20932,N_20960);
nand U24172 (N_24172,N_20368,N_19926);
nand U24173 (N_24173,N_20235,N_18910);
and U24174 (N_24174,N_20904,N_19104);
nor U24175 (N_24175,N_19311,N_21709);
or U24176 (N_24176,N_21859,N_19983);
or U24177 (N_24177,N_19488,N_20569);
nand U24178 (N_24178,N_18776,N_20162);
nor U24179 (N_24179,N_18775,N_21248);
and U24180 (N_24180,N_20384,N_19136);
or U24181 (N_24181,N_21294,N_19293);
xor U24182 (N_24182,N_20666,N_18909);
and U24183 (N_24183,N_20586,N_20022);
nor U24184 (N_24184,N_19338,N_21805);
or U24185 (N_24185,N_21666,N_20645);
and U24186 (N_24186,N_18896,N_19290);
or U24187 (N_24187,N_19106,N_20485);
nand U24188 (N_24188,N_18828,N_20737);
or U24189 (N_24189,N_20572,N_20809);
xor U24190 (N_24190,N_20276,N_20700);
and U24191 (N_24191,N_21354,N_19264);
nor U24192 (N_24192,N_21309,N_19474);
nand U24193 (N_24193,N_20208,N_21734);
nand U24194 (N_24194,N_21377,N_20026);
nor U24195 (N_24195,N_21385,N_20487);
or U24196 (N_24196,N_19623,N_20551);
xnor U24197 (N_24197,N_18831,N_19881);
xor U24198 (N_24198,N_20273,N_19365);
nand U24199 (N_24199,N_21341,N_19209);
or U24200 (N_24200,N_20417,N_21761);
nor U24201 (N_24201,N_21202,N_21540);
nor U24202 (N_24202,N_21401,N_21605);
and U24203 (N_24203,N_20311,N_19065);
nand U24204 (N_24204,N_20437,N_20994);
nor U24205 (N_24205,N_20183,N_21844);
or U24206 (N_24206,N_20694,N_19203);
or U24207 (N_24207,N_21762,N_19009);
nor U24208 (N_24208,N_21317,N_21795);
and U24209 (N_24209,N_19082,N_20232);
nor U24210 (N_24210,N_20926,N_21405);
xor U24211 (N_24211,N_20060,N_21242);
and U24212 (N_24212,N_18757,N_18882);
and U24213 (N_24213,N_20624,N_19410);
or U24214 (N_24214,N_20488,N_20826);
nor U24215 (N_24215,N_20050,N_20226);
xnor U24216 (N_24216,N_20575,N_19131);
nor U24217 (N_24217,N_19503,N_20351);
nor U24218 (N_24218,N_21612,N_20569);
and U24219 (N_24219,N_21422,N_20668);
and U24220 (N_24220,N_19942,N_21622);
nor U24221 (N_24221,N_20352,N_20822);
and U24222 (N_24222,N_19790,N_19202);
xor U24223 (N_24223,N_19178,N_21675);
nand U24224 (N_24224,N_21857,N_19435);
nor U24225 (N_24225,N_20958,N_21350);
nand U24226 (N_24226,N_20798,N_20310);
or U24227 (N_24227,N_21727,N_20196);
and U24228 (N_24228,N_20478,N_18972);
and U24229 (N_24229,N_20952,N_21217);
nor U24230 (N_24230,N_19722,N_21460);
and U24231 (N_24231,N_20167,N_21389);
or U24232 (N_24232,N_19422,N_20468);
nor U24233 (N_24233,N_19806,N_20672);
nand U24234 (N_24234,N_20962,N_21272);
nand U24235 (N_24235,N_21055,N_20344);
nand U24236 (N_24236,N_19217,N_19398);
nor U24237 (N_24237,N_19625,N_21734);
or U24238 (N_24238,N_20416,N_21795);
and U24239 (N_24239,N_19907,N_19552);
and U24240 (N_24240,N_18995,N_19156);
nand U24241 (N_24241,N_20980,N_21692);
or U24242 (N_24242,N_19927,N_21798);
or U24243 (N_24243,N_21725,N_19298);
nand U24244 (N_24244,N_19867,N_20599);
nor U24245 (N_24245,N_20655,N_19448);
xor U24246 (N_24246,N_20950,N_21439);
nand U24247 (N_24247,N_19546,N_20262);
nand U24248 (N_24248,N_20597,N_19464);
or U24249 (N_24249,N_21013,N_19235);
nor U24250 (N_24250,N_20955,N_19098);
or U24251 (N_24251,N_19221,N_21065);
and U24252 (N_24252,N_20813,N_19395);
or U24253 (N_24253,N_19440,N_20013);
and U24254 (N_24254,N_21555,N_20216);
or U24255 (N_24255,N_21706,N_21334);
or U24256 (N_24256,N_20596,N_21354);
xor U24257 (N_24257,N_19793,N_20546);
nand U24258 (N_24258,N_18826,N_20842);
nor U24259 (N_24259,N_21148,N_20301);
xor U24260 (N_24260,N_20881,N_19391);
and U24261 (N_24261,N_21013,N_20471);
xnor U24262 (N_24262,N_18770,N_19456);
and U24263 (N_24263,N_20401,N_18859);
or U24264 (N_24264,N_21585,N_19643);
and U24265 (N_24265,N_19060,N_20957);
xor U24266 (N_24266,N_21236,N_20158);
nand U24267 (N_24267,N_20518,N_19916);
and U24268 (N_24268,N_21621,N_21035);
and U24269 (N_24269,N_19516,N_20004);
or U24270 (N_24270,N_18993,N_18906);
nor U24271 (N_24271,N_19456,N_21048);
nand U24272 (N_24272,N_20305,N_20104);
or U24273 (N_24273,N_21394,N_19289);
and U24274 (N_24274,N_20308,N_19594);
nor U24275 (N_24275,N_19981,N_20741);
and U24276 (N_24276,N_20809,N_21069);
nand U24277 (N_24277,N_21671,N_21571);
nor U24278 (N_24278,N_19447,N_19723);
nor U24279 (N_24279,N_20141,N_19374);
or U24280 (N_24280,N_20340,N_21061);
xnor U24281 (N_24281,N_19863,N_20039);
nand U24282 (N_24282,N_21027,N_19032);
and U24283 (N_24283,N_21012,N_19813);
nor U24284 (N_24284,N_21677,N_19118);
and U24285 (N_24285,N_20887,N_19455);
xor U24286 (N_24286,N_19857,N_20722);
nand U24287 (N_24287,N_19227,N_20816);
and U24288 (N_24288,N_20727,N_21336);
xor U24289 (N_24289,N_19173,N_19769);
nand U24290 (N_24290,N_20153,N_21033);
and U24291 (N_24291,N_19428,N_21139);
and U24292 (N_24292,N_20956,N_19052);
nor U24293 (N_24293,N_20312,N_19383);
nor U24294 (N_24294,N_20365,N_21567);
nor U24295 (N_24295,N_19185,N_18880);
and U24296 (N_24296,N_19154,N_21719);
nand U24297 (N_24297,N_21273,N_21232);
or U24298 (N_24298,N_19104,N_19702);
nand U24299 (N_24299,N_20355,N_21109);
nor U24300 (N_24300,N_21339,N_19661);
or U24301 (N_24301,N_21303,N_19870);
xnor U24302 (N_24302,N_19233,N_19936);
nand U24303 (N_24303,N_18779,N_19471);
and U24304 (N_24304,N_20960,N_20933);
nor U24305 (N_24305,N_21280,N_19758);
or U24306 (N_24306,N_21248,N_21192);
nand U24307 (N_24307,N_19573,N_18753);
nand U24308 (N_24308,N_21749,N_19846);
or U24309 (N_24309,N_20471,N_20220);
and U24310 (N_24310,N_21393,N_19573);
nand U24311 (N_24311,N_21063,N_20636);
or U24312 (N_24312,N_21704,N_20335);
or U24313 (N_24313,N_19322,N_18969);
and U24314 (N_24314,N_20757,N_20631);
nor U24315 (N_24315,N_20204,N_19945);
xor U24316 (N_24316,N_20305,N_21596);
nand U24317 (N_24317,N_19116,N_20637);
and U24318 (N_24318,N_19535,N_21369);
nor U24319 (N_24319,N_20275,N_21580);
and U24320 (N_24320,N_21327,N_18981);
nor U24321 (N_24321,N_19931,N_18802);
and U24322 (N_24322,N_21231,N_19354);
nor U24323 (N_24323,N_19864,N_19945);
nand U24324 (N_24324,N_18833,N_20019);
or U24325 (N_24325,N_21220,N_19460);
nand U24326 (N_24326,N_19379,N_19684);
and U24327 (N_24327,N_20956,N_21808);
and U24328 (N_24328,N_19407,N_20752);
nand U24329 (N_24329,N_19754,N_19889);
nand U24330 (N_24330,N_18900,N_19046);
nand U24331 (N_24331,N_19309,N_21326);
or U24332 (N_24332,N_19297,N_20418);
nor U24333 (N_24333,N_21808,N_19327);
or U24334 (N_24334,N_20873,N_20587);
nor U24335 (N_24335,N_20387,N_20749);
and U24336 (N_24336,N_21422,N_19770);
and U24337 (N_24337,N_20487,N_19489);
or U24338 (N_24338,N_20184,N_21279);
or U24339 (N_24339,N_20569,N_18834);
and U24340 (N_24340,N_21139,N_20894);
xnor U24341 (N_24341,N_19480,N_20692);
nor U24342 (N_24342,N_19714,N_19834);
and U24343 (N_24343,N_20646,N_20315);
nor U24344 (N_24344,N_18802,N_19765);
nor U24345 (N_24345,N_19164,N_19038);
or U24346 (N_24346,N_21625,N_19715);
or U24347 (N_24347,N_20830,N_20113);
xor U24348 (N_24348,N_20791,N_21153);
and U24349 (N_24349,N_21234,N_20958);
nand U24350 (N_24350,N_21229,N_20922);
xor U24351 (N_24351,N_19785,N_19223);
nor U24352 (N_24352,N_19599,N_21629);
or U24353 (N_24353,N_19685,N_19771);
or U24354 (N_24354,N_20646,N_21682);
nor U24355 (N_24355,N_18972,N_20346);
and U24356 (N_24356,N_20186,N_20507);
xor U24357 (N_24357,N_21785,N_21517);
xor U24358 (N_24358,N_19048,N_20952);
nor U24359 (N_24359,N_21844,N_20567);
xor U24360 (N_24360,N_21286,N_20116);
nand U24361 (N_24361,N_19958,N_20448);
nor U24362 (N_24362,N_19111,N_19637);
or U24363 (N_24363,N_19824,N_20611);
nand U24364 (N_24364,N_19847,N_20905);
nor U24365 (N_24365,N_19041,N_18916);
nand U24366 (N_24366,N_20262,N_18969);
nand U24367 (N_24367,N_21792,N_19760);
and U24368 (N_24368,N_18889,N_18866);
or U24369 (N_24369,N_19859,N_20505);
nor U24370 (N_24370,N_19052,N_20544);
nor U24371 (N_24371,N_21278,N_20885);
or U24372 (N_24372,N_20189,N_20036);
nor U24373 (N_24373,N_20478,N_20474);
nand U24374 (N_24374,N_21342,N_19931);
nand U24375 (N_24375,N_21098,N_20527);
nand U24376 (N_24376,N_20048,N_21482);
nor U24377 (N_24377,N_19672,N_20998);
nor U24378 (N_24378,N_21731,N_21638);
or U24379 (N_24379,N_21634,N_20119);
nand U24380 (N_24380,N_21568,N_19806);
or U24381 (N_24381,N_20513,N_18823);
or U24382 (N_24382,N_19481,N_20398);
nand U24383 (N_24383,N_20122,N_21804);
or U24384 (N_24384,N_19274,N_19083);
nand U24385 (N_24385,N_20195,N_20983);
nor U24386 (N_24386,N_20566,N_19617);
or U24387 (N_24387,N_21784,N_19468);
nand U24388 (N_24388,N_19186,N_20458);
or U24389 (N_24389,N_20031,N_20767);
xor U24390 (N_24390,N_21353,N_19869);
and U24391 (N_24391,N_21448,N_21299);
and U24392 (N_24392,N_19321,N_19013);
xnor U24393 (N_24393,N_20869,N_21678);
or U24394 (N_24394,N_18877,N_21356);
or U24395 (N_24395,N_21255,N_20129);
and U24396 (N_24396,N_20987,N_19189);
nand U24397 (N_24397,N_21496,N_19705);
nor U24398 (N_24398,N_20526,N_20609);
or U24399 (N_24399,N_21687,N_19144);
and U24400 (N_24400,N_19979,N_21816);
and U24401 (N_24401,N_19978,N_21464);
nor U24402 (N_24402,N_21210,N_21843);
xnor U24403 (N_24403,N_19348,N_19999);
or U24404 (N_24404,N_19739,N_19313);
or U24405 (N_24405,N_21684,N_20437);
and U24406 (N_24406,N_19213,N_20926);
nand U24407 (N_24407,N_20933,N_21849);
nor U24408 (N_24408,N_19943,N_19419);
nand U24409 (N_24409,N_21131,N_19120);
nor U24410 (N_24410,N_20409,N_20359);
nor U24411 (N_24411,N_21081,N_20151);
and U24412 (N_24412,N_21204,N_19082);
and U24413 (N_24413,N_19532,N_20827);
nand U24414 (N_24414,N_21437,N_19543);
nor U24415 (N_24415,N_19015,N_19266);
xor U24416 (N_24416,N_18965,N_19513);
nand U24417 (N_24417,N_20320,N_19789);
nand U24418 (N_24418,N_19313,N_21640);
nand U24419 (N_24419,N_20166,N_19818);
and U24420 (N_24420,N_19860,N_18877);
nand U24421 (N_24421,N_20958,N_19420);
or U24422 (N_24422,N_21713,N_20153);
nor U24423 (N_24423,N_19371,N_19158);
and U24424 (N_24424,N_21666,N_21632);
xor U24425 (N_24425,N_19164,N_20822);
nand U24426 (N_24426,N_21790,N_21260);
nand U24427 (N_24427,N_19233,N_19485);
xor U24428 (N_24428,N_20700,N_19603);
nor U24429 (N_24429,N_19311,N_21129);
nor U24430 (N_24430,N_21362,N_20497);
nor U24431 (N_24431,N_20779,N_21734);
and U24432 (N_24432,N_18906,N_21320);
and U24433 (N_24433,N_20502,N_21868);
nand U24434 (N_24434,N_19339,N_19472);
nand U24435 (N_24435,N_19093,N_19878);
and U24436 (N_24436,N_21598,N_19202);
xnor U24437 (N_24437,N_21298,N_20647);
nand U24438 (N_24438,N_21658,N_21254);
nor U24439 (N_24439,N_20171,N_19123);
or U24440 (N_24440,N_20740,N_19608);
nand U24441 (N_24441,N_21443,N_21850);
nand U24442 (N_24442,N_20365,N_19217);
or U24443 (N_24443,N_19395,N_19044);
nand U24444 (N_24444,N_21804,N_19235);
xnor U24445 (N_24445,N_18996,N_19921);
xor U24446 (N_24446,N_19966,N_19589);
nor U24447 (N_24447,N_21228,N_19196);
nor U24448 (N_24448,N_21026,N_18935);
and U24449 (N_24449,N_21060,N_18782);
nand U24450 (N_24450,N_19512,N_21369);
and U24451 (N_24451,N_19083,N_19335);
nor U24452 (N_24452,N_20699,N_21456);
nand U24453 (N_24453,N_20394,N_20334);
xor U24454 (N_24454,N_20673,N_18987);
nand U24455 (N_24455,N_21058,N_19763);
and U24456 (N_24456,N_21634,N_19992);
nor U24457 (N_24457,N_19479,N_21276);
and U24458 (N_24458,N_20859,N_18945);
nor U24459 (N_24459,N_19265,N_19195);
and U24460 (N_24460,N_20677,N_21240);
and U24461 (N_24461,N_21293,N_20200);
and U24462 (N_24462,N_19622,N_19041);
nor U24463 (N_24463,N_20090,N_21006);
and U24464 (N_24464,N_19883,N_20776);
nand U24465 (N_24465,N_18910,N_20193);
and U24466 (N_24466,N_19446,N_19318);
or U24467 (N_24467,N_20377,N_19527);
and U24468 (N_24468,N_21120,N_19242);
xor U24469 (N_24469,N_20514,N_19584);
or U24470 (N_24470,N_19763,N_21048);
nor U24471 (N_24471,N_21607,N_20562);
nor U24472 (N_24472,N_21450,N_21131);
or U24473 (N_24473,N_20220,N_19081);
or U24474 (N_24474,N_21483,N_20755);
and U24475 (N_24475,N_19607,N_21322);
and U24476 (N_24476,N_20191,N_20462);
and U24477 (N_24477,N_21119,N_19217);
or U24478 (N_24478,N_21410,N_20016);
nor U24479 (N_24479,N_19294,N_21019);
nand U24480 (N_24480,N_18988,N_19568);
nor U24481 (N_24481,N_19101,N_21702);
and U24482 (N_24482,N_18766,N_20912);
and U24483 (N_24483,N_20162,N_21836);
nor U24484 (N_24484,N_21546,N_18799);
and U24485 (N_24485,N_18886,N_19099);
nand U24486 (N_24486,N_21066,N_20402);
nand U24487 (N_24487,N_19955,N_19501);
nor U24488 (N_24488,N_18879,N_19475);
nand U24489 (N_24489,N_20219,N_19481);
nand U24490 (N_24490,N_19061,N_20177);
nand U24491 (N_24491,N_18974,N_19269);
xnor U24492 (N_24492,N_20331,N_19459);
or U24493 (N_24493,N_19688,N_18840);
nand U24494 (N_24494,N_21546,N_20842);
or U24495 (N_24495,N_20977,N_19493);
or U24496 (N_24496,N_20816,N_19497);
nand U24497 (N_24497,N_19348,N_20894);
or U24498 (N_24498,N_18875,N_20834);
and U24499 (N_24499,N_20662,N_21848);
or U24500 (N_24500,N_19673,N_20013);
or U24501 (N_24501,N_19684,N_19202);
nor U24502 (N_24502,N_19145,N_18967);
nor U24503 (N_24503,N_21713,N_19977);
or U24504 (N_24504,N_20889,N_19965);
xor U24505 (N_24505,N_21185,N_19200);
nor U24506 (N_24506,N_21689,N_20577);
and U24507 (N_24507,N_18843,N_18973);
or U24508 (N_24508,N_19513,N_20545);
and U24509 (N_24509,N_18929,N_20557);
xor U24510 (N_24510,N_21303,N_20315);
or U24511 (N_24511,N_20919,N_20982);
and U24512 (N_24512,N_20444,N_19034);
xor U24513 (N_24513,N_20084,N_20836);
and U24514 (N_24514,N_19684,N_19358);
nand U24515 (N_24515,N_19407,N_19220);
nand U24516 (N_24516,N_21807,N_20915);
nor U24517 (N_24517,N_20590,N_21278);
nand U24518 (N_24518,N_20625,N_21630);
or U24519 (N_24519,N_21789,N_19729);
nand U24520 (N_24520,N_20772,N_20830);
nor U24521 (N_24521,N_20055,N_20740);
and U24522 (N_24522,N_19849,N_20753);
and U24523 (N_24523,N_20529,N_20762);
xnor U24524 (N_24524,N_19100,N_20059);
xor U24525 (N_24525,N_18926,N_21088);
and U24526 (N_24526,N_18975,N_19779);
nand U24527 (N_24527,N_21057,N_19104);
xnor U24528 (N_24528,N_20080,N_20152);
nor U24529 (N_24529,N_20619,N_20989);
nor U24530 (N_24530,N_18922,N_19479);
nor U24531 (N_24531,N_20025,N_19730);
or U24532 (N_24532,N_20579,N_20948);
xor U24533 (N_24533,N_21552,N_19558);
nor U24534 (N_24534,N_20521,N_19671);
xor U24535 (N_24535,N_19800,N_18880);
nand U24536 (N_24536,N_20839,N_20431);
nor U24537 (N_24537,N_21527,N_19026);
or U24538 (N_24538,N_18874,N_21580);
nand U24539 (N_24539,N_21637,N_20170);
or U24540 (N_24540,N_19847,N_21460);
or U24541 (N_24541,N_21314,N_19296);
or U24542 (N_24542,N_19925,N_21744);
and U24543 (N_24543,N_20687,N_20901);
nor U24544 (N_24544,N_20321,N_20169);
and U24545 (N_24545,N_19260,N_20519);
nand U24546 (N_24546,N_21089,N_20308);
nand U24547 (N_24547,N_21038,N_21433);
nand U24548 (N_24548,N_20232,N_21495);
nor U24549 (N_24549,N_20836,N_18940);
xor U24550 (N_24550,N_19664,N_18900);
and U24551 (N_24551,N_21808,N_20961);
nor U24552 (N_24552,N_21304,N_19466);
nand U24553 (N_24553,N_21008,N_20647);
or U24554 (N_24554,N_21111,N_19532);
nor U24555 (N_24555,N_21312,N_19705);
and U24556 (N_24556,N_21686,N_19769);
xor U24557 (N_24557,N_20881,N_19917);
or U24558 (N_24558,N_21279,N_21068);
xnor U24559 (N_24559,N_20278,N_19317);
and U24560 (N_24560,N_21042,N_19076);
or U24561 (N_24561,N_19208,N_19137);
and U24562 (N_24562,N_20720,N_21806);
or U24563 (N_24563,N_19451,N_21479);
and U24564 (N_24564,N_20622,N_19105);
and U24565 (N_24565,N_20169,N_19976);
nor U24566 (N_24566,N_20663,N_19402);
or U24567 (N_24567,N_18904,N_19707);
nand U24568 (N_24568,N_20596,N_20797);
and U24569 (N_24569,N_21460,N_19637);
nor U24570 (N_24570,N_19598,N_20995);
and U24571 (N_24571,N_19436,N_20546);
xor U24572 (N_24572,N_21512,N_20446);
or U24573 (N_24573,N_21714,N_21291);
xnor U24574 (N_24574,N_19123,N_20343);
nand U24575 (N_24575,N_18839,N_20833);
and U24576 (N_24576,N_19307,N_21462);
nand U24577 (N_24577,N_21169,N_19192);
nand U24578 (N_24578,N_18912,N_20196);
xnor U24579 (N_24579,N_21250,N_21410);
nor U24580 (N_24580,N_20734,N_19329);
nor U24581 (N_24581,N_20562,N_21565);
and U24582 (N_24582,N_20859,N_19761);
or U24583 (N_24583,N_19561,N_19346);
nor U24584 (N_24584,N_20767,N_20474);
nand U24585 (N_24585,N_19946,N_19610);
xor U24586 (N_24586,N_20902,N_19626);
and U24587 (N_24587,N_21491,N_19721);
or U24588 (N_24588,N_19280,N_19184);
or U24589 (N_24589,N_19294,N_21771);
or U24590 (N_24590,N_19326,N_21630);
or U24591 (N_24591,N_19471,N_21388);
or U24592 (N_24592,N_21386,N_20165);
and U24593 (N_24593,N_19321,N_18836);
nor U24594 (N_24594,N_19037,N_18837);
xor U24595 (N_24595,N_21524,N_19411);
and U24596 (N_24596,N_21420,N_21339);
nand U24597 (N_24597,N_20056,N_19064);
or U24598 (N_24598,N_21714,N_19587);
or U24599 (N_24599,N_20032,N_18965);
xnor U24600 (N_24600,N_20884,N_20097);
and U24601 (N_24601,N_21522,N_20879);
nor U24602 (N_24602,N_20006,N_20204);
or U24603 (N_24603,N_20980,N_19781);
and U24604 (N_24604,N_20165,N_19853);
and U24605 (N_24605,N_18761,N_21428);
and U24606 (N_24606,N_19140,N_20907);
nand U24607 (N_24607,N_20511,N_18770);
or U24608 (N_24608,N_19285,N_21005);
nor U24609 (N_24609,N_18899,N_19768);
or U24610 (N_24610,N_20569,N_21576);
nand U24611 (N_24611,N_18763,N_20589);
xor U24612 (N_24612,N_19995,N_21333);
nand U24613 (N_24613,N_21451,N_19142);
or U24614 (N_24614,N_19052,N_21400);
and U24615 (N_24615,N_19197,N_21405);
and U24616 (N_24616,N_19479,N_21174);
nand U24617 (N_24617,N_19707,N_21792);
nand U24618 (N_24618,N_18991,N_20226);
nor U24619 (N_24619,N_21741,N_19754);
and U24620 (N_24620,N_20350,N_18846);
or U24621 (N_24621,N_19273,N_20567);
nor U24622 (N_24622,N_19319,N_19484);
nor U24623 (N_24623,N_21801,N_19827);
nand U24624 (N_24624,N_20264,N_20734);
nand U24625 (N_24625,N_20516,N_20373);
nor U24626 (N_24626,N_21263,N_18834);
or U24627 (N_24627,N_21799,N_20541);
xor U24628 (N_24628,N_20073,N_18992);
nor U24629 (N_24629,N_19928,N_19159);
nand U24630 (N_24630,N_19098,N_19055);
or U24631 (N_24631,N_19594,N_19932);
nand U24632 (N_24632,N_19069,N_20031);
or U24633 (N_24633,N_20454,N_19246);
nand U24634 (N_24634,N_21569,N_19645);
xnor U24635 (N_24635,N_20506,N_21530);
or U24636 (N_24636,N_19744,N_20817);
nor U24637 (N_24637,N_21522,N_20542);
and U24638 (N_24638,N_18903,N_20114);
and U24639 (N_24639,N_19612,N_18859);
nor U24640 (N_24640,N_20664,N_19626);
or U24641 (N_24641,N_19527,N_20281);
nor U24642 (N_24642,N_21538,N_19412);
or U24643 (N_24643,N_20050,N_19719);
nor U24644 (N_24644,N_21209,N_19213);
nand U24645 (N_24645,N_19381,N_20158);
or U24646 (N_24646,N_21110,N_19437);
and U24647 (N_24647,N_20800,N_20982);
nand U24648 (N_24648,N_20565,N_19383);
nor U24649 (N_24649,N_21801,N_19082);
or U24650 (N_24650,N_19158,N_19207);
or U24651 (N_24651,N_19512,N_21073);
and U24652 (N_24652,N_19990,N_20160);
or U24653 (N_24653,N_19348,N_21033);
nand U24654 (N_24654,N_19581,N_20464);
and U24655 (N_24655,N_21629,N_21098);
or U24656 (N_24656,N_20682,N_19946);
nor U24657 (N_24657,N_21812,N_19086);
or U24658 (N_24658,N_20024,N_20309);
nor U24659 (N_24659,N_21309,N_21407);
nor U24660 (N_24660,N_19107,N_21381);
nor U24661 (N_24661,N_19534,N_21033);
nor U24662 (N_24662,N_20228,N_20616);
or U24663 (N_24663,N_19334,N_21666);
nor U24664 (N_24664,N_21329,N_20488);
xnor U24665 (N_24665,N_21856,N_19772);
and U24666 (N_24666,N_21034,N_18954);
or U24667 (N_24667,N_19928,N_20101);
nor U24668 (N_24668,N_19879,N_19898);
and U24669 (N_24669,N_21632,N_21327);
and U24670 (N_24670,N_19819,N_20670);
nor U24671 (N_24671,N_21702,N_20529);
nand U24672 (N_24672,N_19463,N_21087);
or U24673 (N_24673,N_20451,N_20410);
xnor U24674 (N_24674,N_21423,N_19651);
nand U24675 (N_24675,N_20550,N_20118);
xnor U24676 (N_24676,N_20877,N_19245);
and U24677 (N_24677,N_18944,N_19935);
or U24678 (N_24678,N_19122,N_19363);
nand U24679 (N_24679,N_20197,N_20015);
xnor U24680 (N_24680,N_19306,N_19226);
nor U24681 (N_24681,N_19362,N_20121);
nand U24682 (N_24682,N_19504,N_21230);
nand U24683 (N_24683,N_20051,N_20941);
nand U24684 (N_24684,N_21659,N_21712);
nor U24685 (N_24685,N_21591,N_21007);
and U24686 (N_24686,N_19701,N_20146);
xor U24687 (N_24687,N_18972,N_19667);
or U24688 (N_24688,N_21231,N_21816);
and U24689 (N_24689,N_19993,N_18860);
or U24690 (N_24690,N_20278,N_19077);
xor U24691 (N_24691,N_19925,N_20532);
nor U24692 (N_24692,N_20481,N_21288);
and U24693 (N_24693,N_21201,N_21459);
or U24694 (N_24694,N_21306,N_21012);
or U24695 (N_24695,N_19505,N_19803);
nand U24696 (N_24696,N_19757,N_20618);
and U24697 (N_24697,N_19732,N_21248);
nor U24698 (N_24698,N_20575,N_21580);
and U24699 (N_24699,N_20411,N_20679);
or U24700 (N_24700,N_19645,N_19452);
xnor U24701 (N_24701,N_19511,N_19424);
or U24702 (N_24702,N_20261,N_19374);
nor U24703 (N_24703,N_21671,N_19520);
nor U24704 (N_24704,N_21380,N_21317);
nand U24705 (N_24705,N_19929,N_21256);
or U24706 (N_24706,N_20427,N_20996);
and U24707 (N_24707,N_20846,N_20083);
or U24708 (N_24708,N_20185,N_21065);
nor U24709 (N_24709,N_20788,N_20744);
nand U24710 (N_24710,N_19017,N_20315);
and U24711 (N_24711,N_19634,N_19171);
nand U24712 (N_24712,N_21126,N_19472);
nand U24713 (N_24713,N_20384,N_21681);
nor U24714 (N_24714,N_21830,N_21530);
nor U24715 (N_24715,N_21170,N_19789);
and U24716 (N_24716,N_21190,N_21088);
and U24717 (N_24717,N_19542,N_21292);
and U24718 (N_24718,N_21459,N_20875);
nand U24719 (N_24719,N_20078,N_19435);
nor U24720 (N_24720,N_19399,N_20431);
nand U24721 (N_24721,N_19512,N_19167);
and U24722 (N_24722,N_19973,N_19232);
or U24723 (N_24723,N_21041,N_19037);
xnor U24724 (N_24724,N_21499,N_21496);
and U24725 (N_24725,N_19889,N_21247);
nor U24726 (N_24726,N_21621,N_20514);
or U24727 (N_24727,N_19547,N_21197);
xnor U24728 (N_24728,N_21152,N_21664);
nor U24729 (N_24729,N_18790,N_21733);
nor U24730 (N_24730,N_21490,N_20780);
or U24731 (N_24731,N_19030,N_20705);
or U24732 (N_24732,N_21823,N_18800);
or U24733 (N_24733,N_21119,N_21664);
or U24734 (N_24734,N_20680,N_21477);
and U24735 (N_24735,N_18861,N_21274);
xor U24736 (N_24736,N_20445,N_20732);
or U24737 (N_24737,N_20540,N_19781);
nand U24738 (N_24738,N_21450,N_21165);
or U24739 (N_24739,N_20919,N_20722);
and U24740 (N_24740,N_19267,N_20842);
or U24741 (N_24741,N_18965,N_21585);
or U24742 (N_24742,N_19133,N_18944);
nor U24743 (N_24743,N_19942,N_19801);
nand U24744 (N_24744,N_19912,N_19866);
or U24745 (N_24745,N_20872,N_21336);
or U24746 (N_24746,N_19567,N_20364);
and U24747 (N_24747,N_19810,N_20998);
nor U24748 (N_24748,N_21543,N_20787);
nor U24749 (N_24749,N_20435,N_20749);
or U24750 (N_24750,N_19851,N_19201);
nand U24751 (N_24751,N_21333,N_20437);
and U24752 (N_24752,N_19110,N_20979);
nor U24753 (N_24753,N_19256,N_21794);
or U24754 (N_24754,N_20987,N_21332);
nor U24755 (N_24755,N_20214,N_21724);
and U24756 (N_24756,N_20577,N_20300);
nor U24757 (N_24757,N_21595,N_19248);
nand U24758 (N_24758,N_21592,N_20948);
nor U24759 (N_24759,N_20788,N_18801);
xor U24760 (N_24760,N_19267,N_19650);
xnor U24761 (N_24761,N_21625,N_19448);
or U24762 (N_24762,N_19526,N_19165);
nor U24763 (N_24763,N_21447,N_18972);
nand U24764 (N_24764,N_20488,N_20874);
and U24765 (N_24765,N_20517,N_20839);
or U24766 (N_24766,N_20391,N_21248);
and U24767 (N_24767,N_21394,N_19689);
nor U24768 (N_24768,N_21832,N_21650);
nor U24769 (N_24769,N_19898,N_19958);
or U24770 (N_24770,N_19664,N_18945);
xor U24771 (N_24771,N_19107,N_21643);
or U24772 (N_24772,N_20513,N_20709);
or U24773 (N_24773,N_20853,N_19747);
and U24774 (N_24774,N_21594,N_18837);
and U24775 (N_24775,N_19162,N_21217);
nor U24776 (N_24776,N_21838,N_21247);
or U24777 (N_24777,N_21504,N_21527);
nand U24778 (N_24778,N_20750,N_19026);
nand U24779 (N_24779,N_20359,N_21796);
and U24780 (N_24780,N_19399,N_18936);
xnor U24781 (N_24781,N_18776,N_19450);
and U24782 (N_24782,N_19753,N_19135);
xor U24783 (N_24783,N_21182,N_21262);
nor U24784 (N_24784,N_21182,N_21791);
nand U24785 (N_24785,N_20887,N_19490);
and U24786 (N_24786,N_21770,N_21274);
nor U24787 (N_24787,N_20032,N_21052);
nand U24788 (N_24788,N_19769,N_20985);
and U24789 (N_24789,N_20990,N_20806);
nor U24790 (N_24790,N_20185,N_19923);
nand U24791 (N_24791,N_19376,N_20321);
nor U24792 (N_24792,N_21148,N_19853);
or U24793 (N_24793,N_20149,N_19975);
and U24794 (N_24794,N_20211,N_21296);
nand U24795 (N_24795,N_21684,N_20785);
and U24796 (N_24796,N_20470,N_19241);
and U24797 (N_24797,N_21267,N_21620);
nand U24798 (N_24798,N_19111,N_19221);
or U24799 (N_24799,N_21692,N_20963);
or U24800 (N_24800,N_21083,N_21474);
nand U24801 (N_24801,N_20708,N_19422);
nand U24802 (N_24802,N_19374,N_19420);
and U24803 (N_24803,N_19266,N_19574);
nand U24804 (N_24804,N_19535,N_20509);
nor U24805 (N_24805,N_18975,N_19930);
and U24806 (N_24806,N_18927,N_19540);
nor U24807 (N_24807,N_19870,N_19392);
nor U24808 (N_24808,N_21744,N_21312);
nor U24809 (N_24809,N_19972,N_21831);
or U24810 (N_24810,N_21782,N_19003);
or U24811 (N_24811,N_21784,N_21671);
or U24812 (N_24812,N_21506,N_21718);
nor U24813 (N_24813,N_21799,N_21702);
xor U24814 (N_24814,N_20586,N_21135);
nand U24815 (N_24815,N_20506,N_20089);
and U24816 (N_24816,N_19087,N_21176);
or U24817 (N_24817,N_19675,N_20323);
nand U24818 (N_24818,N_18843,N_21750);
and U24819 (N_24819,N_19337,N_20121);
and U24820 (N_24820,N_19944,N_19847);
nor U24821 (N_24821,N_18757,N_18836);
and U24822 (N_24822,N_20235,N_19894);
or U24823 (N_24823,N_20330,N_19937);
nor U24824 (N_24824,N_20426,N_19064);
nand U24825 (N_24825,N_19759,N_18842);
nor U24826 (N_24826,N_21495,N_21343);
or U24827 (N_24827,N_21786,N_21683);
nor U24828 (N_24828,N_20950,N_20545);
nor U24829 (N_24829,N_19094,N_20904);
and U24830 (N_24830,N_18905,N_21446);
nor U24831 (N_24831,N_19169,N_21320);
xnor U24832 (N_24832,N_21282,N_21865);
and U24833 (N_24833,N_20314,N_20486);
nand U24834 (N_24834,N_19842,N_19916);
xor U24835 (N_24835,N_21769,N_20083);
nand U24836 (N_24836,N_19470,N_21212);
xor U24837 (N_24837,N_19116,N_19389);
or U24838 (N_24838,N_21198,N_21091);
nor U24839 (N_24839,N_21003,N_20239);
and U24840 (N_24840,N_20047,N_19210);
and U24841 (N_24841,N_21222,N_19177);
nand U24842 (N_24842,N_19676,N_20702);
and U24843 (N_24843,N_21529,N_21278);
xnor U24844 (N_24844,N_20725,N_19271);
and U24845 (N_24845,N_18901,N_21332);
xor U24846 (N_24846,N_21375,N_20886);
and U24847 (N_24847,N_21075,N_21444);
and U24848 (N_24848,N_20192,N_19229);
or U24849 (N_24849,N_21732,N_20410);
and U24850 (N_24850,N_20846,N_18927);
nor U24851 (N_24851,N_21158,N_19085);
nor U24852 (N_24852,N_19839,N_19579);
nor U24853 (N_24853,N_20539,N_19709);
and U24854 (N_24854,N_21165,N_19329);
or U24855 (N_24855,N_21043,N_19024);
or U24856 (N_24856,N_19989,N_21211);
nand U24857 (N_24857,N_21838,N_19254);
or U24858 (N_24858,N_20450,N_21651);
nand U24859 (N_24859,N_18995,N_21758);
nor U24860 (N_24860,N_20832,N_20988);
nand U24861 (N_24861,N_20449,N_19046);
nor U24862 (N_24862,N_18865,N_21266);
nor U24863 (N_24863,N_21863,N_21618);
nand U24864 (N_24864,N_19115,N_21541);
nor U24865 (N_24865,N_20286,N_18957);
nor U24866 (N_24866,N_21497,N_21362);
and U24867 (N_24867,N_21755,N_20666);
and U24868 (N_24868,N_21088,N_18879);
nand U24869 (N_24869,N_21838,N_20935);
nor U24870 (N_24870,N_20359,N_20122);
xor U24871 (N_24871,N_19040,N_19565);
nor U24872 (N_24872,N_20041,N_20701);
or U24873 (N_24873,N_21300,N_20583);
nand U24874 (N_24874,N_21666,N_18953);
or U24875 (N_24875,N_19121,N_21556);
xnor U24876 (N_24876,N_21662,N_19496);
xor U24877 (N_24877,N_20487,N_20313);
xor U24878 (N_24878,N_20973,N_19860);
xnor U24879 (N_24879,N_19256,N_20979);
or U24880 (N_24880,N_20508,N_21291);
and U24881 (N_24881,N_20423,N_20529);
and U24882 (N_24882,N_20768,N_21374);
nor U24883 (N_24883,N_21188,N_20834);
and U24884 (N_24884,N_19200,N_20973);
nand U24885 (N_24885,N_19768,N_20620);
nand U24886 (N_24886,N_21310,N_21824);
nor U24887 (N_24887,N_20240,N_21378);
nand U24888 (N_24888,N_20698,N_20597);
or U24889 (N_24889,N_19958,N_19500);
nor U24890 (N_24890,N_18959,N_21768);
or U24891 (N_24891,N_19030,N_20233);
and U24892 (N_24892,N_20006,N_21792);
and U24893 (N_24893,N_18872,N_21046);
or U24894 (N_24894,N_21377,N_20808);
xnor U24895 (N_24895,N_20802,N_21781);
or U24896 (N_24896,N_19468,N_19571);
and U24897 (N_24897,N_21640,N_19104);
nand U24898 (N_24898,N_21468,N_20833);
xnor U24899 (N_24899,N_19485,N_20129);
nand U24900 (N_24900,N_20231,N_19006);
and U24901 (N_24901,N_21031,N_21189);
and U24902 (N_24902,N_18845,N_20742);
or U24903 (N_24903,N_21693,N_21539);
or U24904 (N_24904,N_20493,N_18769);
xnor U24905 (N_24905,N_20280,N_20454);
nor U24906 (N_24906,N_20153,N_21587);
xnor U24907 (N_24907,N_19210,N_20382);
and U24908 (N_24908,N_21142,N_20883);
or U24909 (N_24909,N_20310,N_19341);
and U24910 (N_24910,N_19883,N_19656);
and U24911 (N_24911,N_20540,N_19908);
nand U24912 (N_24912,N_18916,N_19021);
nor U24913 (N_24913,N_21353,N_20356);
xor U24914 (N_24914,N_19482,N_20182);
or U24915 (N_24915,N_19070,N_20532);
and U24916 (N_24916,N_20717,N_21675);
and U24917 (N_24917,N_20149,N_21302);
nand U24918 (N_24918,N_20628,N_20824);
xnor U24919 (N_24919,N_20682,N_20545);
nor U24920 (N_24920,N_20798,N_19532);
nor U24921 (N_24921,N_20482,N_21305);
nor U24922 (N_24922,N_21466,N_19356);
and U24923 (N_24923,N_20581,N_20551);
and U24924 (N_24924,N_19312,N_21608);
nor U24925 (N_24925,N_19301,N_20693);
nor U24926 (N_24926,N_21816,N_19811);
nor U24927 (N_24927,N_19681,N_21188);
nand U24928 (N_24928,N_21160,N_20377);
or U24929 (N_24929,N_20228,N_20747);
nand U24930 (N_24930,N_19638,N_20965);
nand U24931 (N_24931,N_20554,N_20606);
and U24932 (N_24932,N_19002,N_19976);
nand U24933 (N_24933,N_19885,N_20394);
or U24934 (N_24934,N_19226,N_20288);
and U24935 (N_24935,N_19350,N_20327);
xor U24936 (N_24936,N_18764,N_19460);
and U24937 (N_24937,N_19966,N_19518);
nor U24938 (N_24938,N_21183,N_19966);
or U24939 (N_24939,N_20873,N_21098);
nor U24940 (N_24940,N_19130,N_19444);
and U24941 (N_24941,N_19689,N_21796);
xnor U24942 (N_24942,N_18883,N_19904);
nor U24943 (N_24943,N_19934,N_20416);
xnor U24944 (N_24944,N_20229,N_21556);
or U24945 (N_24945,N_21097,N_19587);
nand U24946 (N_24946,N_20513,N_18767);
nor U24947 (N_24947,N_21383,N_21169);
or U24948 (N_24948,N_19438,N_19405);
nor U24949 (N_24949,N_19419,N_19973);
xnor U24950 (N_24950,N_20739,N_19956);
and U24951 (N_24951,N_21852,N_20835);
nor U24952 (N_24952,N_19121,N_20016);
and U24953 (N_24953,N_21620,N_19797);
and U24954 (N_24954,N_21705,N_20918);
nand U24955 (N_24955,N_21556,N_20115);
nand U24956 (N_24956,N_21234,N_20745);
nand U24957 (N_24957,N_21263,N_19939);
xnor U24958 (N_24958,N_21504,N_21592);
or U24959 (N_24959,N_19988,N_18764);
nor U24960 (N_24960,N_18825,N_19317);
nand U24961 (N_24961,N_19633,N_20063);
nor U24962 (N_24962,N_21705,N_18833);
nor U24963 (N_24963,N_19370,N_19265);
and U24964 (N_24964,N_18825,N_19576);
and U24965 (N_24965,N_21376,N_21195);
and U24966 (N_24966,N_20040,N_19037);
nand U24967 (N_24967,N_19645,N_21587);
nand U24968 (N_24968,N_21815,N_19586);
nand U24969 (N_24969,N_20096,N_20341);
and U24970 (N_24970,N_19623,N_19019);
nor U24971 (N_24971,N_21831,N_19060);
xor U24972 (N_24972,N_21039,N_18983);
and U24973 (N_24973,N_21263,N_20579);
or U24974 (N_24974,N_21537,N_20512);
or U24975 (N_24975,N_21642,N_19574);
nand U24976 (N_24976,N_19970,N_18788);
nor U24977 (N_24977,N_20401,N_18761);
nand U24978 (N_24978,N_19404,N_19961);
nand U24979 (N_24979,N_21665,N_21305);
nor U24980 (N_24980,N_19327,N_18807);
xnor U24981 (N_24981,N_20663,N_19394);
nor U24982 (N_24982,N_18854,N_19877);
nand U24983 (N_24983,N_18838,N_20600);
or U24984 (N_24984,N_20761,N_20686);
nand U24985 (N_24985,N_21164,N_20820);
nor U24986 (N_24986,N_20493,N_19396);
and U24987 (N_24987,N_21490,N_19556);
xor U24988 (N_24988,N_20258,N_19565);
xnor U24989 (N_24989,N_21540,N_21145);
and U24990 (N_24990,N_21318,N_20533);
or U24991 (N_24991,N_20803,N_21161);
and U24992 (N_24992,N_19157,N_21713);
nor U24993 (N_24993,N_19387,N_19947);
or U24994 (N_24994,N_20461,N_19688);
and U24995 (N_24995,N_19859,N_21559);
or U24996 (N_24996,N_21607,N_21062);
and U24997 (N_24997,N_19305,N_21100);
nand U24998 (N_24998,N_21548,N_21820);
xor U24999 (N_24999,N_20748,N_21206);
nand UO_0 (O_0,N_22011,N_23644);
nor UO_1 (O_1,N_24336,N_24567);
xnor UO_2 (O_2,N_24579,N_24597);
or UO_3 (O_3,N_24231,N_23910);
or UO_4 (O_4,N_24834,N_24887);
xnor UO_5 (O_5,N_24990,N_24046);
or UO_6 (O_6,N_23436,N_23716);
nand UO_7 (O_7,N_21962,N_22523);
nand UO_8 (O_8,N_24234,N_24487);
nor UO_9 (O_9,N_24413,N_24528);
and UO_10 (O_10,N_23685,N_23623);
nand UO_11 (O_11,N_24871,N_23162);
or UO_12 (O_12,N_23834,N_23509);
or UO_13 (O_13,N_22764,N_23246);
nand UO_14 (O_14,N_22905,N_24242);
xnor UO_15 (O_15,N_22375,N_24859);
xor UO_16 (O_16,N_23747,N_22411);
or UO_17 (O_17,N_23840,N_22837);
nor UO_18 (O_18,N_24893,N_24237);
nor UO_19 (O_19,N_23822,N_24310);
nand UO_20 (O_20,N_22821,N_21951);
nor UO_21 (O_21,N_22360,N_21933);
or UO_22 (O_22,N_22270,N_24441);
and UO_23 (O_23,N_24855,N_22164);
nand UO_24 (O_24,N_24468,N_24308);
or UO_25 (O_25,N_24381,N_24081);
nor UO_26 (O_26,N_23109,N_23356);
nand UO_27 (O_27,N_24062,N_24130);
or UO_28 (O_28,N_23132,N_21955);
nand UO_29 (O_29,N_24992,N_23468);
and UO_30 (O_30,N_22145,N_23239);
nor UO_31 (O_31,N_22428,N_21969);
nor UO_32 (O_32,N_24374,N_22777);
and UO_33 (O_33,N_22845,N_23758);
nand UO_34 (O_34,N_24019,N_23961);
xor UO_35 (O_35,N_21876,N_22887);
nor UO_36 (O_36,N_22756,N_23086);
nand UO_37 (O_37,N_24017,N_23633);
nand UO_38 (O_38,N_22820,N_24030);
nor UO_39 (O_39,N_23382,N_22989);
nand UO_40 (O_40,N_24809,N_23430);
nand UO_41 (O_41,N_22708,N_22617);
xor UO_42 (O_42,N_24171,N_22319);
nor UO_43 (O_43,N_23155,N_22878);
or UO_44 (O_44,N_22851,N_23577);
or UO_45 (O_45,N_23981,N_24865);
and UO_46 (O_46,N_22746,N_23069);
nor UO_47 (O_47,N_22479,N_23434);
nor UO_48 (O_48,N_24087,N_22947);
or UO_49 (O_49,N_24266,N_22180);
nand UO_50 (O_50,N_24535,N_23927);
nand UO_51 (O_51,N_22147,N_24458);
or UO_52 (O_52,N_24942,N_22805);
nand UO_53 (O_53,N_24898,N_23256);
nor UO_54 (O_54,N_23091,N_22298);
or UO_55 (O_55,N_22836,N_22912);
and UO_56 (O_56,N_23121,N_22525);
nor UO_57 (O_57,N_24802,N_24657);
or UO_58 (O_58,N_22748,N_23049);
and UO_59 (O_59,N_23932,N_24335);
nor UO_60 (O_60,N_22467,N_24720);
or UO_61 (O_61,N_23003,N_24581);
nor UO_62 (O_62,N_24074,N_22075);
nand UO_63 (O_63,N_23228,N_24502);
nor UO_64 (O_64,N_22597,N_22028);
or UO_65 (O_65,N_23360,N_24377);
nor UO_66 (O_66,N_23540,N_22719);
nor UO_67 (O_67,N_23147,N_23576);
xor UO_68 (O_68,N_23921,N_22323);
nor UO_69 (O_69,N_24268,N_23782);
nor UO_70 (O_70,N_23322,N_23774);
nor UO_71 (O_71,N_22600,N_22291);
nand UO_72 (O_72,N_23887,N_24155);
nand UO_73 (O_73,N_23939,N_22302);
nor UO_74 (O_74,N_23108,N_22731);
nand UO_75 (O_75,N_22050,N_22220);
and UO_76 (O_76,N_24613,N_22561);
and UO_77 (O_77,N_24034,N_22374);
xnor UO_78 (O_78,N_23559,N_24544);
or UO_79 (O_79,N_24550,N_24967);
xnor UO_80 (O_80,N_23672,N_22181);
nand UO_81 (O_81,N_24211,N_23312);
or UO_82 (O_82,N_22348,N_23843);
nand UO_83 (O_83,N_22615,N_24519);
and UO_84 (O_84,N_24571,N_22645);
nand UO_85 (O_85,N_23815,N_24209);
or UO_86 (O_86,N_24445,N_24626);
and UO_87 (O_87,N_24921,N_22642);
or UO_88 (O_88,N_23301,N_24257);
or UO_89 (O_89,N_24862,N_22384);
nand UO_90 (O_90,N_23207,N_22172);
nand UO_91 (O_91,N_22728,N_23235);
and UO_92 (O_92,N_23022,N_22659);
nand UO_93 (O_93,N_22857,N_24463);
nor UO_94 (O_94,N_24486,N_23488);
nor UO_95 (O_95,N_23861,N_24765);
or UO_96 (O_96,N_22214,N_22663);
nand UO_97 (O_97,N_22967,N_22611);
xnor UO_98 (O_98,N_22796,N_23056);
nand UO_99 (O_99,N_23988,N_24392);
nand UO_100 (O_100,N_24700,N_24603);
nand UO_101 (O_101,N_24606,N_23689);
nand UO_102 (O_102,N_22937,N_23309);
and UO_103 (O_103,N_21924,N_24818);
and UO_104 (O_104,N_23190,N_22039);
nor UO_105 (O_105,N_24806,N_24988);
and UO_106 (O_106,N_22566,N_22883);
nor UO_107 (O_107,N_24610,N_22520);
nor UO_108 (O_108,N_24536,N_22077);
or UO_109 (O_109,N_24545,N_24972);
or UO_110 (O_110,N_23691,N_22779);
nor UO_111 (O_111,N_23524,N_23817);
and UO_112 (O_112,N_22688,N_24584);
and UO_113 (O_113,N_23094,N_22787);
nor UO_114 (O_114,N_23006,N_22677);
nor UO_115 (O_115,N_22282,N_22193);
xnor UO_116 (O_116,N_23637,N_23619);
xor UO_117 (O_117,N_24848,N_24338);
and UO_118 (O_118,N_21967,N_23385);
xnor UO_119 (O_119,N_24330,N_22293);
xor UO_120 (O_120,N_24758,N_21917);
and UO_121 (O_121,N_23127,N_24852);
nor UO_122 (O_122,N_23258,N_23138);
nand UO_123 (O_123,N_22662,N_22927);
xnor UO_124 (O_124,N_23500,N_22024);
nand UO_125 (O_125,N_23076,N_24555);
nor UO_126 (O_126,N_21894,N_22350);
nor UO_127 (O_127,N_22007,N_22473);
nand UO_128 (O_128,N_22186,N_24140);
nor UO_129 (O_129,N_22847,N_24616);
nor UO_130 (O_130,N_23037,N_24115);
xor UO_131 (O_131,N_24451,N_24228);
or UO_132 (O_132,N_22591,N_24741);
nor UO_133 (O_133,N_24396,N_24345);
nand UO_134 (O_134,N_23184,N_22464);
nand UO_135 (O_135,N_24284,N_24838);
nand UO_136 (O_136,N_22227,N_24901);
and UO_137 (O_137,N_24585,N_22266);
and UO_138 (O_138,N_22674,N_22130);
and UO_139 (O_139,N_23561,N_24215);
or UO_140 (O_140,N_23053,N_24247);
xnor UO_141 (O_141,N_22246,N_23484);
nand UO_142 (O_142,N_23123,N_22741);
nand UO_143 (O_143,N_22735,N_22896);
and UO_144 (O_144,N_22827,N_22529);
nand UO_145 (O_145,N_24051,N_24191);
and UO_146 (O_146,N_24977,N_24746);
nor UO_147 (O_147,N_23522,N_24684);
nor UO_148 (O_148,N_23656,N_23451);
nor UO_149 (O_149,N_24431,N_22084);
nand UO_150 (O_150,N_23553,N_23113);
nand UO_151 (O_151,N_24269,N_24334);
xor UO_152 (O_152,N_21954,N_22672);
or UO_153 (O_153,N_23057,N_24238);
or UO_154 (O_154,N_24154,N_23174);
and UO_155 (O_155,N_24000,N_24744);
nor UO_156 (O_156,N_23205,N_22786);
nor UO_157 (O_157,N_23894,N_22049);
nor UO_158 (O_158,N_24880,N_24542);
nand UO_159 (O_159,N_22290,N_22966);
and UO_160 (O_160,N_23377,N_22539);
nand UO_161 (O_161,N_24907,N_23471);
or UO_162 (O_162,N_22650,N_22134);
nor UO_163 (O_163,N_22461,N_22415);
nand UO_164 (O_164,N_24937,N_23501);
nor UO_165 (O_165,N_23967,N_24240);
and UO_166 (O_166,N_24905,N_22682);
nand UO_167 (O_167,N_22492,N_23379);
nor UO_168 (O_168,N_24936,N_24889);
and UO_169 (O_169,N_24391,N_23265);
nor UO_170 (O_170,N_22144,N_23420);
and UO_171 (O_171,N_24742,N_23450);
nor UO_172 (O_172,N_24143,N_22613);
nand UO_173 (O_173,N_22973,N_22341);
xnor UO_174 (O_174,N_22920,N_23178);
nand UO_175 (O_175,N_24134,N_23852);
or UO_176 (O_176,N_22229,N_24687);
or UO_177 (O_177,N_23418,N_24319);
nand UO_178 (O_178,N_22352,N_23329);
nand UO_179 (O_179,N_22556,N_22151);
or UO_180 (O_180,N_23415,N_24221);
nand UO_181 (O_181,N_22578,N_23074);
nand UO_182 (O_182,N_21975,N_24229);
and UO_183 (O_183,N_24452,N_21880);
and UO_184 (O_184,N_23550,N_22954);
or UO_185 (O_185,N_22394,N_22140);
or UO_186 (O_186,N_23581,N_23290);
xor UO_187 (O_187,N_24253,N_24389);
nor UO_188 (O_188,N_24104,N_23659);
nand UO_189 (O_189,N_22053,N_21949);
nor UO_190 (O_190,N_23135,N_24235);
xor UO_191 (O_191,N_24232,N_22286);
nor UO_192 (O_192,N_24110,N_22074);
nor UO_193 (O_193,N_22793,N_24218);
nand UO_194 (O_194,N_21971,N_22109);
or UO_195 (O_195,N_24931,N_22505);
nand UO_196 (O_196,N_23762,N_22113);
nor UO_197 (O_197,N_22970,N_22395);
xnor UO_198 (O_198,N_23958,N_23532);
and UO_199 (O_199,N_24342,N_22045);
or UO_200 (O_200,N_24149,N_24696);
nand UO_201 (O_201,N_22378,N_22508);
or UO_202 (O_202,N_23586,N_24690);
nor UO_203 (O_203,N_22019,N_24819);
nand UO_204 (O_204,N_22054,N_24174);
and UO_205 (O_205,N_24794,N_23497);
nor UO_206 (O_206,N_23118,N_22648);
or UO_207 (O_207,N_22644,N_22958);
nand UO_208 (O_208,N_24350,N_24793);
nand UO_209 (O_209,N_22906,N_23442);
nand UO_210 (O_210,N_24303,N_24680);
xor UO_211 (O_211,N_24801,N_22183);
nor UO_212 (O_212,N_22148,N_22435);
nand UO_213 (O_213,N_23820,N_23611);
or UO_214 (O_214,N_22828,N_22824);
or UO_215 (O_215,N_24093,N_23479);
or UO_216 (O_216,N_23739,N_22006);
nand UO_217 (O_217,N_22807,N_23064);
and UO_218 (O_218,N_23573,N_22044);
xnor UO_219 (O_219,N_24673,N_24222);
or UO_220 (O_220,N_22998,N_24612);
and UO_221 (O_221,N_22752,N_24077);
nand UO_222 (O_222,N_24733,N_22038);
and UO_223 (O_223,N_24394,N_23938);
xor UO_224 (O_224,N_24586,N_24157);
nand UO_225 (O_225,N_22097,N_22660);
nand UO_226 (O_226,N_24332,N_22440);
nand UO_227 (O_227,N_23759,N_22632);
nor UO_228 (O_228,N_24025,N_24653);
nor UO_229 (O_229,N_22441,N_22722);
or UO_230 (O_230,N_24895,N_23681);
nor UO_231 (O_231,N_21878,N_23182);
nor UO_232 (O_232,N_22577,N_23321);
nand UO_233 (O_233,N_22487,N_24840);
nor UO_234 (O_234,N_22707,N_22198);
nor UO_235 (O_235,N_24991,N_23307);
nor UO_236 (O_236,N_23279,N_22297);
nor UO_237 (O_237,N_22488,N_22060);
nand UO_238 (O_238,N_24493,N_23039);
and UO_239 (O_239,N_23883,N_21963);
or UO_240 (O_240,N_23917,N_22726);
or UO_241 (O_241,N_24210,N_23324);
nor UO_242 (O_242,N_23068,N_23499);
nor UO_243 (O_243,N_24291,N_24861);
nor UO_244 (O_244,N_22939,N_24122);
xor UO_245 (O_245,N_24812,N_22849);
nand UO_246 (O_246,N_22742,N_21960);
nor UO_247 (O_247,N_22736,N_23605);
nand UO_248 (O_248,N_22507,N_21926);
and UO_249 (O_249,N_21911,N_22965);
or UO_250 (O_250,N_23911,N_22629);
and UO_251 (O_251,N_24023,N_22718);
and UO_252 (O_252,N_23206,N_22607);
nand UO_253 (O_253,N_23195,N_24691);
and UO_254 (O_254,N_21928,N_24633);
nor UO_255 (O_255,N_24123,N_24792);
nand UO_256 (O_256,N_23261,N_21906);
nand UO_257 (O_257,N_24343,N_24828);
xnor UO_258 (O_258,N_24915,N_23873);
nand UO_259 (O_259,N_24164,N_24710);
and UO_260 (O_260,N_22397,N_22749);
or UO_261 (O_261,N_22775,N_24021);
nand UO_262 (O_262,N_24817,N_23350);
or UO_263 (O_263,N_23160,N_22163);
and UO_264 (O_264,N_23765,N_21980);
nand UO_265 (O_265,N_24899,N_24418);
nand UO_266 (O_266,N_23300,N_22103);
or UO_267 (O_267,N_23598,N_24436);
and UO_268 (O_268,N_24661,N_24196);
xnor UO_269 (O_269,N_22637,N_23240);
nor UO_270 (O_270,N_22098,N_21939);
nor UO_271 (O_271,N_24922,N_24595);
nand UO_272 (O_272,N_23084,N_23720);
xnor UO_273 (O_273,N_22889,N_24572);
xnor UO_274 (O_274,N_23862,N_22313);
and UO_275 (O_275,N_23931,N_24485);
and UO_276 (O_276,N_23083,N_23714);
and UO_277 (O_277,N_24704,N_23713);
xor UO_278 (O_278,N_22800,N_24011);
nor UO_279 (O_279,N_22080,N_22862);
and UO_280 (O_280,N_22940,N_24444);
or UO_281 (O_281,N_24668,N_21922);
or UO_282 (O_282,N_22021,N_23455);
or UO_283 (O_283,N_24379,N_24026);
or UO_284 (O_284,N_24024,N_23342);
xnor UO_285 (O_285,N_23915,N_24146);
nand UO_286 (O_286,N_23390,N_22686);
xnor UO_287 (O_287,N_22499,N_22733);
nand UO_288 (O_288,N_22223,N_22537);
or UO_289 (O_289,N_24040,N_22991);
nor UO_290 (O_290,N_23472,N_22706);
or UO_291 (O_291,N_23165,N_22961);
xnor UO_292 (O_292,N_22171,N_21990);
nand UO_293 (O_293,N_23133,N_24596);
or UO_294 (O_294,N_22831,N_23715);
nand UO_295 (O_295,N_23443,N_23475);
or UO_296 (O_296,N_22919,N_24782);
or UO_297 (O_297,N_22249,N_22226);
and UO_298 (O_298,N_24609,N_24730);
nand UO_299 (O_299,N_22734,N_23845);
nor UO_300 (O_300,N_22612,N_22225);
and UO_301 (O_301,N_23569,N_22359);
or UO_302 (O_302,N_23166,N_24872);
nand UO_303 (O_303,N_22243,N_24968);
or UO_304 (O_304,N_23146,N_24490);
and UO_305 (O_305,N_24096,N_24402);
nand UO_306 (O_306,N_24594,N_21957);
nand UO_307 (O_307,N_24461,N_23051);
xor UO_308 (O_308,N_22610,N_23215);
and UO_309 (O_309,N_24701,N_23869);
or UO_310 (O_310,N_22609,N_24035);
and UO_311 (O_311,N_24136,N_22913);
nand UO_312 (O_312,N_23802,N_22085);
and UO_313 (O_313,N_23250,N_23730);
and UO_314 (O_314,N_22004,N_23337);
nand UO_315 (O_315,N_23331,N_22729);
and UO_316 (O_316,N_24286,N_24190);
and UO_317 (O_317,N_21945,N_22311);
nand UO_318 (O_318,N_24446,N_23340);
nor UO_319 (O_319,N_21921,N_24152);
xnor UO_320 (O_320,N_24217,N_23687);
or UO_321 (O_321,N_24472,N_22801);
nand UO_322 (O_322,N_22550,N_23947);
and UO_323 (O_323,N_24158,N_24719);
nand UO_324 (O_324,N_22468,N_24280);
nand UO_325 (O_325,N_24662,N_24843);
nand UO_326 (O_326,N_23694,N_23679);
and UO_327 (O_327,N_23814,N_24534);
nand UO_328 (O_328,N_24422,N_23989);
or UO_329 (O_329,N_23630,N_24849);
nand UO_330 (O_330,N_23233,N_23936);
nor UO_331 (O_331,N_22278,N_22195);
nor UO_332 (O_332,N_23303,N_24230);
or UO_333 (O_333,N_23226,N_24156);
nand UO_334 (O_334,N_22056,N_22964);
nand UO_335 (O_335,N_24781,N_22868);
or UO_336 (O_336,N_22622,N_23131);
nor UO_337 (O_337,N_23800,N_23372);
nor UO_338 (O_338,N_22304,N_24560);
nand UO_339 (O_339,N_22251,N_24999);
nor UO_340 (O_340,N_23529,N_23618);
nand UO_341 (O_341,N_22437,N_24067);
nand UO_342 (O_342,N_22673,N_23650);
or UO_343 (O_343,N_24941,N_22497);
or UO_344 (O_344,N_23425,N_24857);
and UO_345 (O_345,N_23027,N_23589);
nand UO_346 (O_346,N_22414,N_24750);
nor UO_347 (O_347,N_22699,N_24114);
or UO_348 (O_348,N_23139,N_24649);
or UO_349 (O_349,N_23191,N_23032);
xnor UO_350 (O_350,N_23404,N_23567);
nand UO_351 (O_351,N_23962,N_22299);
or UO_352 (O_352,N_23036,N_24900);
and UO_353 (O_353,N_22396,N_23120);
nand UO_354 (O_354,N_22274,N_23310);
and UO_355 (O_355,N_24362,N_23722);
and UO_356 (O_356,N_23327,N_23217);
nor UO_357 (O_357,N_24370,N_24489);
nor UO_358 (O_358,N_22649,N_23317);
or UO_359 (O_359,N_22239,N_22369);
or UO_360 (O_360,N_22176,N_24405);
nor UO_361 (O_361,N_22541,N_23386);
xor UO_362 (O_362,N_22003,N_23588);
and UO_363 (O_363,N_21927,N_22325);
nor UO_364 (O_364,N_23628,N_22772);
xor UO_365 (O_365,N_23695,N_23624);
nand UO_366 (O_366,N_23399,N_22854);
or UO_367 (O_367,N_21958,N_21987);
nor UO_368 (O_368,N_24983,N_23394);
nand UO_369 (O_369,N_23103,N_24356);
nand UO_370 (O_370,N_24103,N_23009);
or UO_371 (O_371,N_22009,N_24996);
xnor UO_372 (O_372,N_24403,N_21937);
and UO_373 (O_373,N_23507,N_24955);
nand UO_374 (O_374,N_24307,N_24706);
and UO_375 (O_375,N_24213,N_23908);
nor UO_376 (O_376,N_21976,N_24902);
nor UO_377 (O_377,N_23371,N_23014);
and UO_378 (O_378,N_23306,N_21999);
and UO_379 (O_379,N_23643,N_23859);
or UO_380 (O_380,N_22386,N_22197);
nand UO_381 (O_381,N_23987,N_22261);
nand UO_382 (O_382,N_22565,N_22101);
nand UO_383 (O_383,N_24762,N_24602);
and UO_384 (O_384,N_23073,N_23208);
nand UO_385 (O_385,N_22480,N_22408);
or UO_386 (O_386,N_22231,N_22549);
nand UO_387 (O_387,N_23535,N_22737);
or UO_388 (O_388,N_23159,N_24961);
nand UO_389 (O_389,N_22554,N_24789);
and UO_390 (O_390,N_22212,N_24117);
or UO_391 (O_391,N_22112,N_23737);
or UO_392 (O_392,N_24060,N_23106);
or UO_393 (O_393,N_22562,N_22242);
nand UO_394 (O_394,N_23515,N_24978);
nand UO_395 (O_395,N_21905,N_24482);
or UO_396 (O_396,N_23362,N_24951);
and UO_397 (O_397,N_22139,N_21988);
nor UO_398 (O_398,N_22013,N_24283);
and UO_399 (O_399,N_24301,N_23531);
or UO_400 (O_400,N_23960,N_23344);
nand UO_401 (O_401,N_23848,N_22546);
nand UO_402 (O_402,N_23993,N_24499);
and UO_403 (O_403,N_22806,N_22988);
nand UO_404 (O_404,N_24462,N_23140);
nand UO_405 (O_405,N_22483,N_23419);
nor UO_406 (O_406,N_24787,N_23851);
and UO_407 (O_407,N_23245,N_24755);
and UO_408 (O_408,N_24292,N_23366);
and UO_409 (O_409,N_23710,N_24929);
and UO_410 (O_410,N_23411,N_23287);
xor UO_411 (O_411,N_24775,N_23920);
nand UO_412 (O_412,N_22608,N_23042);
nand UO_413 (O_413,N_22856,N_23330);
xor UO_414 (O_414,N_24749,N_22335);
nand UO_415 (O_415,N_24904,N_22391);
or UO_416 (O_416,N_21950,N_23760);
or UO_417 (O_417,N_24650,N_24644);
and UO_418 (O_418,N_24611,N_22711);
or UO_419 (O_419,N_22863,N_23842);
and UO_420 (O_420,N_23836,N_23732);
and UO_421 (O_421,N_24360,N_22956);
nand UO_422 (O_422,N_22938,N_24496);
nand UO_423 (O_423,N_23568,N_23065);
and UO_424 (O_424,N_24648,N_24264);
or UO_425 (O_425,N_22292,N_22143);
xnor UO_426 (O_426,N_23899,N_23614);
nor UO_427 (O_427,N_24008,N_22982);
nor UO_428 (O_428,N_23526,N_23487);
xor UO_429 (O_429,N_24767,N_24016);
nor UO_430 (O_430,N_23518,N_22758);
nand UO_431 (O_431,N_23895,N_23652);
nand UO_432 (O_432,N_24070,N_22853);
nand UO_433 (O_433,N_24722,N_22587);
or UO_434 (O_434,N_24717,N_23089);
nand UO_435 (O_435,N_22633,N_23119);
or UO_436 (O_436,N_24548,N_23653);
nand UO_437 (O_437,N_22126,N_24005);
or UO_438 (O_438,N_23128,N_24768);
nand UO_439 (O_439,N_23383,N_21965);
nor UO_440 (O_440,N_24688,N_23516);
nor UO_441 (O_441,N_23878,N_24491);
nand UO_442 (O_442,N_23092,N_21974);
nor UO_443 (O_443,N_23352,N_23703);
or UO_444 (O_444,N_24290,N_24891);
or UO_445 (O_445,N_22190,N_21943);
nor UO_446 (O_446,N_24655,N_23122);
xor UO_447 (O_447,N_22058,N_24090);
nor UO_448 (O_448,N_24388,N_24289);
and UO_449 (O_449,N_24304,N_22349);
or UO_450 (O_450,N_23244,N_21895);
or UO_451 (O_451,N_22570,N_24300);
nand UO_452 (O_452,N_24830,N_24415);
nor UO_453 (O_453,N_22926,N_23945);
or UO_454 (O_454,N_22679,N_24224);
nor UO_455 (O_455,N_22738,N_24642);
nor UO_456 (O_456,N_24979,N_22819);
and UO_457 (O_457,N_22027,N_24677);
and UO_458 (O_458,N_24826,N_24565);
and UO_459 (O_459,N_23474,N_22064);
nor UO_460 (O_460,N_24364,N_24440);
or UO_461 (O_461,N_22055,N_24348);
and UO_462 (O_462,N_22710,N_23426);
and UO_463 (O_463,N_24770,N_23816);
nand UO_464 (O_464,N_23634,N_22205);
or UO_465 (O_465,N_22517,N_24888);
nor UO_466 (O_466,N_24393,N_24091);
nand UO_467 (O_467,N_23696,N_22848);
and UO_468 (O_468,N_24325,N_24363);
xor UO_469 (O_469,N_23682,N_24724);
or UO_470 (O_470,N_22560,N_23562);
and UO_471 (O_471,N_22066,N_23761);
or UO_472 (O_472,N_22052,N_24800);
or UO_473 (O_473,N_24698,N_24438);
xor UO_474 (O_474,N_22388,N_23163);
and UO_475 (O_475,N_22252,N_23098);
and UO_476 (O_476,N_23546,N_23054);
or UO_477 (O_477,N_22122,N_22656);
nor UO_478 (O_478,N_23863,N_24417);
and UO_479 (O_479,N_24531,N_24219);
or UO_480 (O_480,N_24557,N_23173);
nand UO_481 (O_481,N_23361,N_23222);
nand UO_482 (O_482,N_23683,N_23251);
nor UO_483 (O_483,N_22675,N_24745);
xnor UO_484 (O_484,N_23158,N_22153);
nor UO_485 (O_485,N_24095,N_24250);
nand UO_486 (O_486,N_24271,N_22209);
nand UO_487 (O_487,N_23583,N_23566);
and UO_488 (O_488,N_23595,N_22953);
nor UO_489 (O_489,N_24854,N_22502);
or UO_490 (O_490,N_24876,N_23414);
nand UO_491 (O_491,N_22888,N_24837);
nor UO_492 (O_492,N_22002,N_23176);
nor UO_493 (O_493,N_23354,N_24678);
nand UO_494 (O_494,N_22766,N_24404);
nor UO_495 (O_495,N_24294,N_23050);
and UO_496 (O_496,N_22757,N_23698);
nor UO_497 (O_497,N_22977,N_22639);
or UO_498 (O_498,N_21994,N_23647);
nor UO_499 (O_499,N_22141,N_23460);
nand UO_500 (O_500,N_22543,N_23775);
or UO_501 (O_501,N_23607,N_24637);
and UO_502 (O_502,N_23552,N_24950);
and UO_503 (O_503,N_23170,N_22745);
nor UO_504 (O_504,N_22201,N_23323);
or UO_505 (O_505,N_24246,N_24708);
nand UO_506 (O_506,N_24197,N_23667);
nand UO_507 (O_507,N_23104,N_22385);
nand UO_508 (O_508,N_22783,N_23757);
nor UO_509 (O_509,N_24697,N_23482);
nor UO_510 (O_510,N_22364,N_22850);
nor UO_511 (O_511,N_22192,N_22340);
xnor UO_512 (O_512,N_24537,N_24359);
nand UO_513 (O_513,N_22469,N_23444);
or UO_514 (O_514,N_21920,N_23130);
and UO_515 (O_515,N_22356,N_22264);
and UO_516 (O_516,N_24395,N_22713);
xnor UO_517 (O_517,N_23786,N_23844);
or UO_518 (O_518,N_22690,N_23070);
and UO_519 (O_519,N_24168,N_23891);
or UO_520 (O_520,N_22199,N_24845);
and UO_521 (O_521,N_24761,N_23900);
or UO_522 (O_522,N_23437,N_23789);
nand UO_523 (O_523,N_22312,N_24810);
xor UO_524 (O_524,N_23857,N_21995);
and UO_525 (O_525,N_22876,N_23403);
nor UO_526 (O_526,N_24501,N_23270);
or UO_527 (O_527,N_24368,N_23992);
or UO_528 (O_528,N_24656,N_24600);
or UO_529 (O_529,N_24339,N_24408);
or UO_530 (O_530,N_22018,N_22630);
or UO_531 (O_531,N_22761,N_22747);
and UO_532 (O_532,N_22767,N_22476);
or UO_533 (O_533,N_23755,N_22361);
xor UO_534 (O_534,N_23890,N_22925);
nand UO_535 (O_535,N_22516,N_23072);
or UO_536 (O_536,N_23314,N_22986);
nand UO_537 (O_537,N_22259,N_24667);
or UO_538 (O_538,N_23734,N_23071);
and UO_539 (O_539,N_24779,N_23870);
and UO_540 (O_540,N_22874,N_23242);
or UO_541 (O_541,N_22972,N_22640);
nand UO_542 (O_542,N_22125,N_22247);
xor UO_543 (O_543,N_21925,N_22115);
and UO_544 (O_544,N_22771,N_22338);
and UO_545 (O_545,N_24175,N_23082);
or UO_546 (O_546,N_22890,N_24663);
nor UO_547 (O_547,N_22753,N_22347);
nor UO_548 (O_548,N_24409,N_22185);
and UO_549 (O_549,N_24387,N_24514);
and UO_550 (O_550,N_24740,N_24055);
xnor UO_551 (O_551,N_23726,N_23214);
or UO_552 (O_552,N_24299,N_24851);
and UO_553 (O_553,N_23519,N_22132);
nor UO_554 (O_554,N_23295,N_22160);
nand UO_555 (O_555,N_22284,N_23678);
nand UO_556 (O_556,N_24167,N_22908);
nand UO_557 (O_557,N_22111,N_21897);
nand UO_558 (O_558,N_23364,N_23697);
xor UO_559 (O_559,N_22031,N_23373);
and UO_560 (O_560,N_22794,N_24142);
xor UO_561 (O_561,N_23884,N_23249);
or UO_562 (O_562,N_24913,N_23416);
or UO_563 (O_563,N_24313,N_22826);
or UO_564 (O_564,N_24317,N_24320);
or UO_565 (O_565,N_23807,N_23541);
and UO_566 (O_566,N_22023,N_24957);
or UO_567 (O_567,N_22217,N_24966);
nor UO_568 (O_568,N_24315,N_22416);
and UO_569 (O_569,N_22237,N_23012);
nand UO_570 (O_570,N_23609,N_24689);
nand UO_571 (O_571,N_24116,N_22701);
xor UO_572 (O_572,N_21942,N_22449);
xor UO_573 (O_573,N_22995,N_24881);
nor UO_574 (O_574,N_22563,N_23658);
nand UO_575 (O_575,N_22162,N_22465);
nand UO_576 (O_576,N_23302,N_22020);
and UO_577 (O_577,N_24166,N_23943);
xnor UO_578 (O_578,N_22750,N_24419);
and UO_579 (O_579,N_22484,N_24207);
and UO_580 (O_580,N_22294,N_24448);
or UO_581 (O_581,N_23276,N_24976);
and UO_582 (O_582,N_22337,N_23610);
and UO_583 (O_583,N_23804,N_22526);
nor UO_584 (O_584,N_22929,N_22393);
nand UO_585 (O_585,N_23728,N_23902);
nand UO_586 (O_586,N_23473,N_23912);
nand UO_587 (O_587,N_24427,N_22255);
xor UO_588 (O_588,N_24188,N_22166);
and UO_589 (O_589,N_23771,N_24367);
nand UO_590 (O_590,N_22451,N_23368);
nand UO_591 (O_591,N_24523,N_23978);
and UO_592 (O_592,N_23821,N_23335);
nor UO_593 (O_593,N_24144,N_24475);
and UO_594 (O_594,N_24912,N_24552);
nor UO_595 (O_595,N_23741,N_23751);
and UO_596 (O_596,N_23596,N_22512);
nand UO_597 (O_597,N_24150,N_24721);
or UO_598 (O_598,N_24088,N_24302);
and UO_599 (O_599,N_24260,N_24270);
nor UO_600 (O_600,N_22263,N_22308);
and UO_601 (O_601,N_23431,N_24263);
and UO_602 (O_602,N_22230,N_22285);
xor UO_603 (O_603,N_23286,N_23353);
xnor UO_604 (O_604,N_23044,N_23066);
or UO_605 (O_605,N_23389,N_23591);
or UO_606 (O_606,N_23028,N_22533);
or UO_607 (O_607,N_23427,N_22515);
xnor UO_608 (O_608,N_23828,N_23880);
nand UO_609 (O_609,N_21889,N_23477);
and UO_610 (O_610,N_22695,N_23781);
nand UO_611 (O_611,N_22138,N_22839);
xnor UO_612 (O_612,N_24956,N_22877);
and UO_613 (O_613,N_22833,N_23102);
or UO_614 (O_614,N_23795,N_22029);
nor UO_615 (O_615,N_23785,N_22945);
and UO_616 (O_616,N_24566,N_24316);
nor UO_617 (O_617,N_23554,N_23955);
or UO_618 (O_618,N_24037,N_24153);
nor UO_619 (O_619,N_22789,N_23923);
or UO_620 (O_620,N_24033,N_23401);
and UO_621 (O_621,N_23305,N_22893);
or UO_622 (O_622,N_22689,N_23801);
xor UO_623 (O_623,N_24699,N_23391);
and UO_624 (O_624,N_22918,N_22008);
and UO_625 (O_625,N_23793,N_24635);
and UO_626 (O_626,N_24193,N_24084);
nand UO_627 (O_627,N_23168,N_24686);
and UO_628 (O_628,N_24997,N_23584);
nor UO_629 (O_629,N_22643,N_23005);
nand UO_630 (O_630,N_23230,N_24883);
nand UO_631 (O_631,N_23615,N_22202);
nand UO_632 (O_632,N_23575,N_24546);
nor UO_633 (O_633,N_24054,N_24480);
nand UO_634 (O_634,N_22530,N_21996);
nor UO_635 (O_635,N_24549,N_24541);
or UO_636 (O_636,N_23349,N_24974);
and UO_637 (O_637,N_24520,N_24752);
and UO_638 (O_638,N_23060,N_22079);
nand UO_639 (O_639,N_23972,N_23429);
or UO_640 (O_640,N_22169,N_24647);
nor UO_641 (O_641,N_23274,N_24474);
and UO_642 (O_642,N_22346,N_22802);
and UO_643 (O_643,N_24305,N_23202);
and UO_644 (O_644,N_24827,N_21898);
or UO_645 (O_645,N_23810,N_24910);
nor UO_646 (O_646,N_24753,N_23966);
nand UO_647 (O_647,N_22191,N_22534);
nor UO_648 (O_648,N_23711,N_23448);
and UO_649 (O_649,N_24058,N_22812);
nand UO_650 (O_650,N_23956,N_23684);
or UO_651 (O_651,N_24989,N_21956);
xor UO_652 (O_652,N_22089,N_24672);
and UO_653 (O_653,N_21892,N_24715);
xnor UO_654 (O_654,N_22712,N_23153);
or UO_655 (O_655,N_24998,N_23151);
and UO_656 (O_656,N_22557,N_24593);
or UO_657 (O_657,N_24517,N_23152);
nand UO_658 (O_658,N_24399,N_22167);
nand UO_659 (O_659,N_23664,N_22732);
or UO_660 (O_660,N_23078,N_23918);
and UO_661 (O_661,N_21948,N_24492);
nand UO_662 (O_662,N_23105,N_24601);
nand UO_663 (O_663,N_24214,N_24428);
or UO_664 (O_664,N_21981,N_23913);
and UO_665 (O_665,N_22474,N_24986);
nand UO_666 (O_666,N_24666,N_23975);
nand UO_667 (O_667,N_24926,N_21993);
xor UO_668 (O_668,N_22458,N_23809);
nor UO_669 (O_669,N_22310,N_22322);
nand UO_670 (O_670,N_23985,N_24412);
xnor UO_671 (O_671,N_24780,N_23928);
and UO_672 (O_672,N_23196,N_22280);
nor UO_673 (O_673,N_24592,N_22762);
nor UO_674 (O_674,N_24694,N_22616);
nor UO_675 (O_675,N_24729,N_22620);
and UO_676 (O_676,N_23204,N_22065);
or UO_677 (O_677,N_24098,N_24220);
xnor UO_678 (O_678,N_22324,N_24614);
nor UO_679 (O_679,N_24705,N_22303);
or UO_680 (O_680,N_24113,N_23642);
nor UO_681 (O_681,N_24120,N_22133);
or UO_682 (O_682,N_24473,N_23101);
nor UO_683 (O_683,N_22981,N_22426);
xnor UO_684 (O_684,N_22365,N_22383);
and UO_685 (O_685,N_23538,N_24524);
or UO_686 (O_686,N_22447,N_22326);
nor UO_687 (O_687,N_24119,N_22715);
nand UO_688 (O_688,N_24530,N_24012);
and UO_689 (O_689,N_23579,N_22117);
nor UO_690 (O_690,N_22493,N_22048);
and UO_691 (O_691,N_24846,N_24351);
nor UO_692 (O_692,N_24867,N_22067);
nand UO_693 (O_693,N_22879,N_22866);
or UO_694 (O_694,N_23602,N_22107);
and UO_695 (O_695,N_24879,N_24112);
nand UO_696 (O_696,N_22524,N_23746);
nor UO_697 (O_697,N_23129,N_24411);
or UO_698 (O_698,N_24366,N_24869);
or UO_699 (O_699,N_23971,N_22135);
or UO_700 (O_700,N_22182,N_22078);
nor UO_701 (O_701,N_22317,N_24760);
nor UO_702 (O_702,N_23660,N_24599);
and UO_703 (O_703,N_23234,N_22852);
or UO_704 (O_704,N_22072,N_22471);
or UO_705 (O_705,N_22575,N_22368);
nor UO_706 (O_706,N_22880,N_22454);
nand UO_707 (O_707,N_23000,N_23423);
nand UO_708 (O_708,N_23875,N_22692);
and UO_709 (O_709,N_22327,N_22475);
or UO_710 (O_710,N_23736,N_24275);
nor UO_711 (O_711,N_23087,N_21877);
and UO_712 (O_712,N_22624,N_22379);
nor UO_713 (O_713,N_22720,N_23052);
and UO_714 (O_714,N_23351,N_22683);
or UO_715 (O_715,N_24790,N_24897);
or UO_716 (O_716,N_23058,N_24709);
xor UO_717 (O_717,N_24454,N_24788);
nand UO_718 (O_718,N_24738,N_22559);
or UO_719 (O_719,N_22985,N_24340);
xnor UO_720 (O_720,N_23381,N_23916);
xnor UO_721 (O_721,N_23413,N_23824);
nand UO_722 (O_722,N_23282,N_23047);
xor UO_723 (O_723,N_22037,N_23026);
and UO_724 (O_724,N_24450,N_23100);
nand UO_725 (O_725,N_23002,N_23970);
xnor UO_726 (O_726,N_22288,N_22859);
nand UO_727 (O_727,N_24028,N_22096);
and UO_728 (O_728,N_24798,N_23141);
nand UO_729 (O_729,N_21979,N_24829);
and UO_730 (O_730,N_24503,N_22840);
or UO_731 (O_731,N_23629,N_23662);
nor UO_732 (O_732,N_21884,N_22207);
or UO_733 (O_733,N_23384,N_22861);
xnor UO_734 (O_734,N_23849,N_24433);
and UO_735 (O_735,N_24437,N_24975);
and UO_736 (O_736,N_22792,N_22922);
and UO_737 (O_737,N_23485,N_22636);
and UO_738 (O_738,N_24932,N_24182);
or UO_739 (O_739,N_24163,N_24131);
xnor UO_740 (O_740,N_24886,N_22932);
nor UO_741 (O_741,N_24401,N_23409);
nor UO_742 (O_742,N_23243,N_23493);
and UO_743 (O_743,N_24086,N_23081);
or UO_744 (O_744,N_22705,N_24556);
nand UO_745 (O_745,N_23269,N_22962);
nand UO_746 (O_746,N_24406,N_23877);
or UO_747 (O_747,N_22944,N_23527);
or UO_748 (O_748,N_23735,N_24126);
nor UO_749 (O_749,N_24097,N_22443);
nand UO_750 (O_750,N_22087,N_22948);
xnor UO_751 (O_751,N_23896,N_22928);
and UO_752 (O_752,N_24162,N_24309);
nor UO_753 (O_753,N_24604,N_23187);
nor UO_754 (O_754,N_23783,N_22960);
or UO_755 (O_755,N_23458,N_21941);
and UO_756 (O_756,N_22882,N_23740);
and UO_757 (O_757,N_22522,N_23547);
nor UO_758 (O_758,N_23557,N_22581);
nand UO_759 (O_759,N_22646,N_23267);
and UO_760 (O_760,N_24916,N_22795);
or UO_761 (O_761,N_24285,N_22872);
or UO_762 (O_762,N_24919,N_24858);
or UO_763 (O_763,N_23536,N_23367);
and UO_764 (O_764,N_23799,N_22030);
or UO_765 (O_765,N_23930,N_22498);
or UO_766 (O_766,N_23879,N_23161);
or UO_767 (O_767,N_22258,N_22987);
and UO_768 (O_768,N_23210,N_22398);
nand UO_769 (O_769,N_23560,N_24878);
and UO_770 (O_770,N_23021,N_23582);
or UO_771 (O_771,N_24080,N_23453);
or UO_772 (O_772,N_22099,N_23537);
xor UO_773 (O_773,N_22455,N_23750);
nand UO_774 (O_774,N_24695,N_24106);
nand UO_775 (O_775,N_24179,N_22418);
nor UO_776 (O_776,N_22614,N_22664);
or UO_777 (O_777,N_24518,N_24773);
or UO_778 (O_778,N_22090,N_22320);
nor UO_779 (O_779,N_22818,N_22495);
and UO_780 (O_780,N_22552,N_24841);
xor UO_781 (O_781,N_22015,N_22569);
or UO_782 (O_782,N_24727,N_24962);
nand UO_783 (O_783,N_23212,N_24564);
nor UO_784 (O_784,N_24620,N_22511);
nand UO_785 (O_785,N_22924,N_23417);
or UO_786 (O_786,N_23045,N_22403);
nand UO_787 (O_787,N_23565,N_23742);
and UO_788 (O_788,N_23316,N_21940);
nor UO_789 (O_789,N_22331,N_23649);
nand UO_790 (O_790,N_22042,N_22277);
nor UO_791 (O_791,N_22685,N_23483);
nand UO_792 (O_792,N_22946,N_22838);
nor UO_793 (O_793,N_24497,N_22892);
or UO_794 (O_794,N_22528,N_23223);
or UO_795 (O_795,N_23999,N_24692);
nand UO_796 (O_796,N_22670,N_24607);
and UO_797 (O_797,N_22619,N_22061);
or UO_798 (O_798,N_24526,N_24276);
nand UO_799 (O_799,N_23023,N_22158);
nand UO_800 (O_800,N_23017,N_23898);
or UO_801 (O_801,N_24508,N_22694);
xor UO_802 (O_802,N_23494,N_23973);
and UO_803 (O_803,N_22477,N_23639);
nor UO_804 (O_804,N_22187,N_24823);
nand UO_805 (O_805,N_23661,N_24227);
nand UO_806 (O_806,N_23788,N_23892);
nor UO_807 (O_807,N_24842,N_22564);
nor UO_808 (O_808,N_21992,N_24894);
and UO_809 (O_809,N_24132,N_23640);
nor UO_810 (O_810,N_24397,N_22963);
and UO_811 (O_811,N_24873,N_22071);
nor UO_812 (O_812,N_22309,N_23200);
or UO_813 (O_813,N_23991,N_24447);
or UO_814 (O_814,N_22224,N_23358);
or UO_815 (O_815,N_22921,N_23754);
and UO_816 (O_816,N_23855,N_23646);
or UO_817 (O_817,N_23142,N_22903);
and UO_818 (O_818,N_22235,N_22997);
and UO_819 (O_819,N_24466,N_22248);
and UO_820 (O_820,N_22835,N_22943);
nand UO_821 (O_821,N_21918,N_23941);
or UO_822 (O_822,N_24265,N_24273);
or UO_823 (O_823,N_22001,N_22161);
nor UO_824 (O_824,N_21900,N_23199);
xnor UO_825 (O_825,N_23797,N_22971);
nor UO_826 (O_826,N_24971,N_21883);
nand UO_827 (O_827,N_23339,N_23397);
and UO_828 (O_828,N_22823,N_23203);
nand UO_829 (O_829,N_22241,N_22257);
nand UO_830 (O_830,N_23463,N_23038);
or UO_831 (O_831,N_24748,N_21890);
xnor UO_832 (O_832,N_23556,N_24836);
nand UO_833 (O_833,N_24206,N_22785);
or UO_834 (O_834,N_23040,N_23853);
nand UO_835 (O_835,N_22897,N_23764);
nor UO_836 (O_836,N_23169,N_24844);
nand UO_837 (O_837,N_22716,N_23019);
or UO_838 (O_838,N_22404,N_22353);
xnor UO_839 (O_839,N_24954,N_23124);
or UO_840 (O_840,N_23925,N_24032);
or UO_841 (O_841,N_23271,N_24036);
or UO_842 (O_842,N_23974,N_22822);
or UO_843 (O_843,N_22102,N_24459);
nand UO_844 (O_844,N_24646,N_24712);
or UO_845 (O_845,N_23183,N_22816);
or UO_846 (O_846,N_22496,N_24772);
nand UO_847 (O_847,N_23829,N_22433);
nor UO_848 (O_848,N_22626,N_22025);
or UO_849 (O_849,N_24065,N_24498);
nor UO_850 (O_850,N_21931,N_24928);
xnor UO_851 (O_851,N_23172,N_22236);
or UO_852 (O_852,N_22544,N_22506);
or UO_853 (O_853,N_23008,N_23291);
and UO_854 (O_854,N_23357,N_24481);
or UO_855 (O_855,N_24043,N_23984);
nor UO_856 (O_856,N_24510,N_23937);
or UO_857 (O_857,N_24958,N_23294);
and UO_858 (O_858,N_23268,N_22121);
and UO_859 (O_859,N_23723,N_23259);
and UO_860 (O_860,N_22316,N_23995);
nand UO_861 (O_861,N_24151,N_22073);
and UO_862 (O_862,N_24833,N_24183);
or UO_863 (O_863,N_24737,N_24416);
or UO_864 (O_864,N_22572,N_23705);
and UO_865 (O_865,N_24262,N_23749);
and UO_866 (O_866,N_24766,N_23440);
or UO_867 (O_867,N_23355,N_22532);
xor UO_868 (O_868,N_24177,N_23665);
nand UO_869 (O_869,N_22366,N_23865);
nor UO_870 (O_870,N_24776,N_22265);
nand UO_871 (O_871,N_23940,N_22124);
xnor UO_872 (O_872,N_23593,N_21938);
or UO_873 (O_873,N_24344,N_24049);
or UO_874 (O_874,N_22470,N_23293);
and UO_875 (O_875,N_23115,N_23763);
and UO_876 (O_876,N_24439,N_22430);
and UO_877 (O_877,N_24638,N_23263);
or UO_878 (O_878,N_24892,N_22486);
or UO_879 (O_879,N_22407,N_24639);
nor UO_880 (O_880,N_23635,N_22653);
nor UO_881 (O_881,N_24981,N_24509);
xor UO_882 (O_882,N_22466,N_23114);
nand UO_883 (O_883,N_24914,N_22760);
nand UO_884 (O_884,N_24532,N_24799);
xnor UO_885 (O_885,N_24365,N_22189);
and UO_886 (O_886,N_24007,N_24636);
and UO_887 (O_887,N_23504,N_21934);
or UO_888 (O_888,N_23025,N_23702);
nor UO_889 (O_889,N_22438,N_22931);
nor UO_890 (O_890,N_24476,N_23563);
and UO_891 (O_891,N_24608,N_22864);
nor UO_892 (O_892,N_24430,N_24835);
nor UO_893 (O_893,N_22881,N_22358);
nand UO_894 (O_894,N_23369,N_23606);
xnor UO_895 (O_895,N_23289,N_22262);
and UO_896 (O_896,N_22036,N_24629);
xor UO_897 (O_897,N_22051,N_22923);
nand UO_898 (O_898,N_24674,N_23011);
nor UO_899 (O_899,N_23674,N_23055);
nor UO_900 (O_900,N_24953,N_22041);
nand UO_901 (O_901,N_23313,N_23530);
nand UO_902 (O_902,N_24133,N_24890);
nand UO_903 (O_903,N_23061,N_23496);
xor UO_904 (O_904,N_22152,N_23673);
xor UO_905 (O_905,N_23534,N_22016);
nor UO_906 (O_906,N_23523,N_24425);
nor UO_907 (O_907,N_24318,N_22788);
nand UO_908 (O_908,N_22228,N_23926);
or UO_909 (O_909,N_23502,N_24908);
nand UO_910 (O_910,N_24627,N_21986);
nor UO_911 (O_911,N_24582,N_23676);
or UO_912 (O_912,N_23398,N_24641);
and UO_913 (O_913,N_24443,N_23819);
and UO_914 (O_914,N_24774,N_22769);
nand UO_915 (O_915,N_22941,N_24732);
nand UO_916 (O_916,N_22104,N_22419);
xor UO_917 (O_917,N_22427,N_24124);
nand UO_918 (O_918,N_24625,N_22593);
xor UO_919 (O_919,N_24298,N_24314);
and UO_920 (O_920,N_24652,N_24778);
and UO_921 (O_921,N_23185,N_23671);
or UO_922 (O_922,N_22781,N_22123);
or UO_923 (O_923,N_24102,N_24529);
xor UO_924 (O_924,N_24631,N_22307);
nand UO_925 (O_925,N_22628,N_23976);
and UO_926 (O_926,N_23858,N_22233);
or UO_927 (O_927,N_22417,N_24354);
nand UO_928 (O_928,N_23492,N_22780);
and UO_929 (O_929,N_23677,N_24052);
nand UO_930 (O_930,N_23167,N_23097);
and UO_931 (O_931,N_23508,N_22032);
or UO_932 (O_932,N_23218,N_24038);
nand UO_933 (O_933,N_23278,N_24288);
and UO_934 (O_934,N_22188,N_23847);
or UO_935 (O_935,N_23262,N_21923);
or UO_936 (O_936,N_24076,N_24059);
or UO_937 (O_937,N_22588,N_24516);
nand UO_938 (O_938,N_24660,N_23048);
nor UO_939 (O_939,N_22213,N_23830);
nand UO_940 (O_940,N_24756,N_23638);
and UO_941 (O_941,N_23134,N_24328);
nand UO_942 (O_942,N_23213,N_23348);
or UO_943 (O_943,N_22975,N_24651);
or UO_944 (O_944,N_23542,N_22842);
or UO_945 (O_945,N_24147,N_24118);
nand UO_946 (O_946,N_24066,N_23838);
nor UO_947 (O_947,N_23211,N_24643);
nand UO_948 (O_948,N_23445,N_23248);
and UO_949 (O_949,N_23315,N_22318);
or UO_950 (O_950,N_22791,N_22910);
xor UO_951 (O_951,N_22724,N_22798);
xor UO_952 (O_952,N_23175,N_24039);
nand UO_953 (O_953,N_24875,N_22315);
or UO_954 (O_954,N_22333,N_24337);
nor UO_955 (O_955,N_22667,N_23319);
and UO_956 (O_956,N_23446,N_23548);
xnor UO_957 (O_957,N_22033,N_23533);
or UO_958 (O_958,N_24831,N_23919);
or UO_959 (O_959,N_24906,N_24202);
or UO_960 (O_960,N_21968,N_23935);
and UO_961 (O_961,N_24071,N_22131);
and UO_962 (O_962,N_23675,N_21915);
or UO_963 (O_963,N_23990,N_23654);
and UO_964 (O_964,N_23221,N_22576);
nand UO_965 (O_965,N_22902,N_22159);
and UO_966 (O_966,N_22585,N_24948);
nand UO_967 (O_967,N_24369,N_22173);
nor UO_968 (O_968,N_22996,N_23965);
nand UO_969 (O_969,N_24832,N_23148);
or UO_970 (O_970,N_22332,N_22300);
nor UO_971 (O_971,N_22494,N_24079);
or UO_972 (O_972,N_22177,N_22094);
or UO_973 (O_973,N_23209,N_23837);
nor UO_974 (O_974,N_22873,N_21901);
nand UO_975 (O_975,N_24045,N_22272);
xnor UO_976 (O_976,N_22432,N_24515);
nor UO_977 (O_977,N_24815,N_22717);
or UO_978 (O_978,N_23934,N_24850);
and UO_979 (O_979,N_22489,N_24312);
or UO_980 (O_980,N_22095,N_23592);
or UO_981 (O_981,N_23603,N_22116);
nand UO_982 (O_982,N_22504,N_22057);
and UO_983 (O_983,N_21929,N_24973);
nor UO_984 (O_984,N_23277,N_24321);
xor UO_985 (O_985,N_24681,N_22146);
or UO_986 (O_986,N_24807,N_23622);
nand UO_987 (O_987,N_24985,N_23909);
nand UO_988 (O_988,N_24769,N_23668);
or UO_989 (O_989,N_24683,N_23954);
nand UO_990 (O_990,N_24181,N_23388);
nand UO_991 (O_991,N_21978,N_23464);
and UO_992 (O_992,N_23881,N_23145);
nand UO_993 (O_993,N_22935,N_23254);
and UO_994 (O_994,N_23343,N_22603);
and UO_995 (O_995,N_23570,N_23778);
nor UO_996 (O_996,N_24353,N_23435);
xnor UO_997 (O_997,N_23551,N_23882);
and UO_998 (O_998,N_24824,N_23296);
nand UO_999 (O_999,N_22829,N_22355);
and UO_1000 (O_1000,N_24771,N_24010);
nor UO_1001 (O_1001,N_21881,N_23299);
nand UO_1002 (O_1002,N_23708,N_22082);
nand UO_1003 (O_1003,N_23457,N_24669);
and UO_1004 (O_1004,N_22260,N_23365);
and UO_1005 (O_1005,N_23669,N_23827);
nand UO_1006 (O_1006,N_23461,N_22093);
or UO_1007 (O_1007,N_22413,N_23798);
xnor UO_1008 (O_1008,N_22768,N_23498);
xor UO_1009 (O_1009,N_23590,N_22509);
and UO_1010 (O_1010,N_22178,N_22681);
nor UO_1011 (O_1011,N_22334,N_23983);
xnor UO_1012 (O_1012,N_23247,N_23986);
nand UO_1013 (O_1013,N_22363,N_21991);
nand UO_1014 (O_1014,N_22070,N_22436);
nor UO_1015 (O_1015,N_23601,N_23874);
xnor UO_1016 (O_1016,N_22703,N_22105);
xor UO_1017 (O_1017,N_24658,N_24736);
nor UO_1018 (O_1018,N_24398,N_22527);
and UO_1019 (O_1019,N_22551,N_22271);
or UO_1020 (O_1020,N_23001,N_23015);
nand UO_1021 (O_1021,N_24107,N_22655);
or UO_1022 (O_1022,N_24424,N_24868);
nand UO_1023 (O_1023,N_23856,N_22119);
and UO_1024 (O_1024,N_22647,N_22869);
nor UO_1025 (O_1025,N_24751,N_22448);
or UO_1026 (O_1026,N_23201,N_24376);
or UO_1027 (O_1027,N_22573,N_22797);
and UO_1028 (O_1028,N_22330,N_22170);
nand UO_1029 (O_1029,N_22203,N_21909);
and UO_1030 (O_1030,N_24559,N_24380);
and UO_1031 (O_1031,N_24161,N_23766);
or UO_1032 (O_1032,N_23555,N_22380);
nor UO_1033 (O_1033,N_24212,N_23621);
or UO_1034 (O_1034,N_22452,N_24022);
nor UO_1035 (O_1035,N_24654,N_24574);
nand UO_1036 (O_1036,N_23380,N_24243);
xor UO_1037 (O_1037,N_24189,N_23264);
and UO_1038 (O_1038,N_23745,N_22809);
or UO_1039 (O_1039,N_23868,N_24575);
nand UO_1040 (O_1040,N_24141,N_23359);
xor UO_1041 (O_1041,N_23224,N_24420);
nand UO_1042 (O_1042,N_22218,N_24075);
nand UO_1043 (O_1043,N_24903,N_23099);
and UO_1044 (O_1044,N_23030,N_23564);
xor UO_1045 (O_1045,N_23998,N_23636);
and UO_1046 (O_1046,N_24429,N_24471);
and UO_1047 (O_1047,N_23831,N_24538);
nand UO_1048 (O_1048,N_22917,N_23034);
and UO_1049 (O_1049,N_22446,N_21885);
and UO_1050 (O_1050,N_22245,N_24186);
or UO_1051 (O_1051,N_24505,N_22086);
nor UO_1052 (O_1052,N_21904,N_23116);
nor UO_1053 (O_1053,N_23818,N_23893);
and UO_1054 (O_1054,N_23670,N_22759);
or UO_1055 (O_1055,N_22638,N_24279);
nand UO_1056 (O_1056,N_23558,N_22598);
nand UO_1057 (O_1057,N_23769,N_24129);
or UO_1058 (O_1058,N_22950,N_22855);
xnor UO_1059 (O_1059,N_24791,N_24553);
nor UO_1060 (O_1060,N_22328,N_22875);
and UO_1061 (O_1061,N_23231,N_24723);
nand UO_1062 (O_1062,N_24617,N_23510);
nand UO_1063 (O_1063,N_23752,N_24679);
and UO_1064 (O_1064,N_23866,N_22727);
or UO_1065 (O_1065,N_22547,N_22371);
or UO_1066 (O_1066,N_23864,N_22040);
nand UO_1067 (O_1067,N_22372,N_22755);
nand UO_1068 (O_1068,N_24013,N_23336);
xnor UO_1069 (O_1069,N_22567,N_22244);
or UO_1070 (O_1070,N_22604,N_22491);
xnor UO_1071 (O_1071,N_24469,N_23171);
xnor UO_1072 (O_1072,N_24184,N_24199);
nand UO_1073 (O_1073,N_23503,N_22936);
or UO_1074 (O_1074,N_23393,N_22344);
and UO_1075 (O_1075,N_23232,N_22730);
xnor UO_1076 (O_1076,N_21887,N_23004);
or UO_1077 (O_1077,N_24002,N_22580);
nor UO_1078 (O_1078,N_23608,N_23318);
nand UO_1079 (O_1079,N_22157,N_22399);
nand UO_1080 (O_1080,N_24960,N_24874);
or UO_1081 (O_1081,N_22618,N_24522);
nand UO_1082 (O_1082,N_24057,N_22952);
and UO_1083 (O_1083,N_24331,N_24747);
nand UO_1084 (O_1084,N_24233,N_23823);
nor UO_1085 (O_1085,N_23273,N_24127);
or UO_1086 (O_1086,N_24053,N_22283);
nor UO_1087 (O_1087,N_23345,N_24665);
xnor UO_1088 (O_1088,N_23075,N_24825);
and UO_1089 (O_1089,N_21899,N_22114);
or UO_1090 (O_1090,N_24252,N_24573);
nand UO_1091 (O_1091,N_24371,N_23090);
and UO_1092 (O_1092,N_24245,N_23812);
or UO_1093 (O_1093,N_23549,N_23651);
or UO_1094 (O_1094,N_22510,N_23035);
nand UO_1095 (O_1095,N_23197,N_24495);
nor UO_1096 (O_1096,N_24588,N_23545);
nor UO_1097 (O_1097,N_22012,N_24707);
nand UO_1098 (O_1098,N_22814,N_22900);
nor UO_1099 (O_1099,N_24964,N_23311);
nor UO_1100 (O_1100,N_23476,N_24346);
nand UO_1101 (O_1101,N_22165,N_24676);
and UO_1102 (O_1102,N_23625,N_22933);
nand UO_1103 (O_1103,N_22811,N_24078);
nor UO_1104 (O_1104,N_24877,N_24814);
and UO_1105 (O_1105,N_23994,N_23525);
and UO_1106 (O_1106,N_23517,N_24216);
xor UO_1107 (O_1107,N_22959,N_24372);
or UO_1108 (O_1108,N_22582,N_22778);
and UO_1109 (O_1109,N_23253,N_24094);
nand UO_1110 (O_1110,N_24675,N_22179);
nand UO_1111 (O_1111,N_23236,N_24583);
nor UO_1112 (O_1112,N_22276,N_22651);
or UO_1113 (O_1113,N_22721,N_22702);
xor UO_1114 (O_1114,N_23860,N_23452);
nand UO_1115 (O_1115,N_23370,N_24554);
and UO_1116 (O_1116,N_23304,N_23901);
nand UO_1117 (O_1117,N_23257,N_24347);
nand UO_1118 (O_1118,N_22150,N_22744);
nor UO_1119 (O_1119,N_22142,N_22482);
and UO_1120 (O_1120,N_23738,N_23188);
or UO_1121 (O_1121,N_22295,N_23229);
nor UO_1122 (O_1122,N_24925,N_23627);
nor UO_1123 (O_1123,N_24909,N_23680);
nor UO_1124 (O_1124,N_24159,N_24711);
and UO_1125 (O_1125,N_24959,N_22373);
and UO_1126 (O_1126,N_24731,N_23376);
nor UO_1127 (O_1127,N_24165,N_24031);
nor UO_1128 (O_1128,N_22657,N_22751);
or UO_1129 (O_1129,N_23275,N_22763);
and UO_1130 (O_1130,N_24200,N_24521);
nand UO_1131 (O_1131,N_24050,N_23977);
nor UO_1132 (O_1132,N_22083,N_22765);
nand UO_1133 (O_1133,N_22595,N_24410);
or UO_1134 (O_1134,N_21952,N_22658);
nand UO_1135 (O_1135,N_24563,N_24896);
nand UO_1136 (O_1136,N_24170,N_24225);
or UO_1137 (O_1137,N_24064,N_22680);
nor UO_1138 (O_1138,N_23712,N_22208);
nor UO_1139 (O_1139,N_23753,N_24804);
and UO_1140 (O_1140,N_23024,N_23238);
or UO_1141 (O_1141,N_23717,N_22904);
xnor UO_1142 (O_1142,N_22420,N_22754);
nor UO_1143 (O_1143,N_24820,N_23933);
or UO_1144 (O_1144,N_24725,N_24101);
nor UO_1145 (O_1145,N_23950,N_23907);
or UO_1146 (O_1146,N_24180,N_23666);
and UO_1147 (O_1147,N_23422,N_22206);
nor UO_1148 (O_1148,N_24382,N_22934);
or UO_1149 (O_1149,N_22422,N_24917);
and UO_1150 (O_1150,N_24373,N_24796);
or UO_1151 (O_1151,N_23010,N_22389);
and UO_1152 (O_1152,N_23428,N_22623);
nand UO_1153 (O_1153,N_23079,N_23117);
and UO_1154 (O_1154,N_24255,N_24864);
nand UO_1155 (O_1155,N_22909,N_22860);
or UO_1156 (O_1156,N_23969,N_23407);
nand UO_1157 (O_1157,N_22059,N_24970);
or UO_1158 (O_1158,N_23041,N_22696);
nor UO_1159 (O_1159,N_23406,N_22536);
nor UO_1160 (O_1160,N_24125,N_23886);
nor UO_1161 (O_1161,N_22005,N_22976);
and UO_1162 (O_1162,N_23744,N_23095);
and UO_1163 (O_1163,N_23721,N_22574);
nand UO_1164 (O_1164,N_22485,N_23952);
nor UO_1165 (O_1165,N_22062,N_22503);
xor UO_1166 (O_1166,N_23470,N_21985);
nor UO_1167 (O_1167,N_22669,N_24083);
or UO_1168 (O_1168,N_24137,N_23832);
or UO_1169 (O_1169,N_24477,N_24576);
nand UO_1170 (O_1170,N_22046,N_23626);
nor UO_1171 (O_1171,N_23835,N_24258);
nor UO_1172 (O_1172,N_23284,N_24640);
or UO_1173 (O_1173,N_23466,N_23029);
nor UO_1174 (O_1174,N_23164,N_24685);
and UO_1175 (O_1175,N_23421,N_22671);
and UO_1176 (O_1176,N_23805,N_23587);
and UO_1177 (O_1177,N_21959,N_24488);
nor UO_1178 (O_1178,N_22571,N_24352);
or UO_1179 (O_1179,N_23885,N_23572);
nand UO_1180 (O_1180,N_24426,N_24984);
or UO_1181 (O_1181,N_24527,N_21998);
and UO_1182 (O_1182,N_22200,N_24805);
nand UO_1183 (O_1183,N_24241,N_22951);
xnor UO_1184 (O_1184,N_22590,N_24944);
or UO_1185 (O_1185,N_24407,N_22799);
xor UO_1186 (O_1186,N_22267,N_21907);
nor UO_1187 (O_1187,N_23181,N_22661);
nand UO_1188 (O_1188,N_24702,N_24783);
nor UO_1189 (O_1189,N_22412,N_22010);
or UO_1190 (O_1190,N_23663,N_24870);
nand UO_1191 (O_1191,N_23107,N_24580);
nand UO_1192 (O_1192,N_24201,N_23520);
or UO_1193 (O_1193,N_24821,N_22184);
or UO_1194 (O_1194,N_23400,N_22993);
and UO_1195 (O_1195,N_22453,N_24484);
nor UO_1196 (O_1196,N_24716,N_22627);
nand UO_1197 (O_1197,N_22602,N_23363);
or UO_1198 (O_1198,N_22289,N_22709);
nor UO_1199 (O_1199,N_23489,N_24384);
nand UO_1200 (O_1200,N_22668,N_22434);
and UO_1201 (O_1201,N_24918,N_22456);
and UO_1202 (O_1202,N_23252,N_22583);
nor UO_1203 (O_1203,N_21944,N_22542);
nor UO_1204 (O_1204,N_22782,N_22376);
nand UO_1205 (O_1205,N_22460,N_24866);
nand UO_1206 (O_1206,N_24068,N_24598);
nor UO_1207 (O_1207,N_23914,N_24759);
nand UO_1208 (O_1208,N_24296,N_23544);
and UO_1209 (O_1209,N_22770,N_23018);
or UO_1210 (O_1210,N_22519,N_22354);
nand UO_1211 (O_1211,N_22942,N_22254);
nand UO_1212 (O_1212,N_23088,N_24927);
or UO_1213 (O_1213,N_23571,N_22275);
xnor UO_1214 (O_1214,N_23062,N_22601);
and UO_1215 (O_1215,N_23424,N_24464);
nand UO_1216 (O_1216,N_21913,N_24839);
xor UO_1217 (O_1217,N_23718,N_22034);
nor UO_1218 (O_1218,N_24329,N_23904);
nand UO_1219 (O_1219,N_21908,N_24853);
nor UO_1220 (O_1220,N_24539,N_24816);
and UO_1221 (O_1221,N_22957,N_24435);
nor UO_1222 (O_1222,N_24223,N_24500);
and UO_1223 (O_1223,N_22631,N_22081);
xor UO_1224 (O_1224,N_24587,N_24108);
nand UO_1225 (O_1225,N_24085,N_22253);
or UO_1226 (O_1226,N_23016,N_23889);
or UO_1227 (O_1227,N_24282,N_22400);
nor UO_1228 (O_1228,N_24003,N_23924);
nand UO_1229 (O_1229,N_22535,N_22342);
nand UO_1230 (O_1230,N_22803,N_24483);
or UO_1231 (O_1231,N_22870,N_23792);
nor UO_1232 (O_1232,N_22584,N_23441);
nor UO_1233 (O_1233,N_22625,N_22704);
nor UO_1234 (O_1234,N_24390,N_23727);
nand UO_1235 (O_1235,N_22980,N_22834);
nor UO_1236 (O_1236,N_24947,N_24763);
and UO_1237 (O_1237,N_22825,N_24295);
nor UO_1238 (O_1238,N_23241,N_24176);
xnor UO_1239 (O_1239,N_23031,N_24287);
nor UO_1240 (O_1240,N_22678,N_23077);
xnor UO_1241 (O_1241,N_22599,N_23410);
and UO_1242 (O_1242,N_24847,N_22314);
or UO_1243 (O_1243,N_21983,N_21970);
nor UO_1244 (O_1244,N_22268,N_22886);
nand UO_1245 (O_1245,N_24943,N_22621);
or UO_1246 (O_1246,N_24621,N_24195);
or UO_1247 (O_1247,N_23180,N_21947);
nor UO_1248 (O_1248,N_22450,N_22287);
or UO_1249 (O_1249,N_24924,N_23285);
nor UO_1250 (O_1250,N_24455,N_22867);
nand UO_1251 (O_1251,N_24808,N_22665);
nor UO_1252 (O_1252,N_22634,N_24204);
nand UO_1253 (O_1253,N_22339,N_23433);
and UO_1254 (O_1254,N_23980,N_23996);
or UO_1255 (O_1255,N_24811,N_23454);
and UO_1256 (O_1256,N_23375,N_22017);
xnor UO_1257 (O_1257,N_24994,N_24047);
nor UO_1258 (O_1258,N_22885,N_24645);
nor UO_1259 (O_1259,N_23465,N_22871);
xor UO_1260 (O_1260,N_23481,N_24965);
and UO_1261 (O_1261,N_24670,N_22901);
xnor UO_1262 (O_1262,N_23903,N_23085);
nor UO_1263 (O_1263,N_23111,N_24465);
xor UO_1264 (O_1264,N_22992,N_23020);
nand UO_1265 (O_1265,N_24293,N_23825);
nand UO_1266 (O_1266,N_22221,N_24735);
or UO_1267 (O_1267,N_23219,N_22994);
nand UO_1268 (O_1268,N_24272,N_23768);
nand UO_1269 (O_1269,N_22444,N_23288);
and UO_1270 (O_1270,N_24226,N_24073);
nor UO_1271 (O_1271,N_24856,N_23707);
or UO_1272 (O_1272,N_23266,N_24187);
nand UO_1273 (O_1273,N_21903,N_22830);
or UO_1274 (O_1274,N_24513,N_22401);
or UO_1275 (O_1275,N_24361,N_24558);
nor UO_1276 (O_1276,N_24442,N_21930);
nand UO_1277 (O_1277,N_22128,N_24099);
or UO_1278 (O_1278,N_24009,N_24739);
nor UO_1279 (O_1279,N_22043,N_24764);
nor UO_1280 (O_1280,N_22687,N_24044);
and UO_1281 (O_1281,N_21932,N_24457);
nor UO_1282 (O_1282,N_24048,N_22990);
or UO_1283 (O_1283,N_24027,N_24533);
or UO_1284 (O_1284,N_23942,N_22739);
xnor UO_1285 (O_1285,N_24277,N_23641);
or UO_1286 (O_1286,N_22969,N_24267);
and UO_1287 (O_1287,N_22329,N_22127);
xnor UO_1288 (O_1288,N_24323,N_23796);
and UO_1289 (O_1289,N_24069,N_23780);
or UO_1290 (O_1290,N_24949,N_23704);
and UO_1291 (O_1291,N_22204,N_24386);
nor UO_1292 (O_1292,N_24591,N_24072);
and UO_1293 (O_1293,N_22429,N_24934);
and UO_1294 (O_1294,N_22377,N_24139);
and UO_1295 (O_1295,N_23395,N_22979);
nor UO_1296 (O_1296,N_24203,N_22714);
and UO_1297 (O_1297,N_24138,N_22301);
nand UO_1298 (O_1298,N_23688,N_24333);
or UO_1299 (O_1299,N_24414,N_23144);
and UO_1300 (O_1300,N_23949,N_24623);
and UO_1301 (O_1301,N_23787,N_22279);
nor UO_1302 (O_1302,N_23013,N_22250);
nor UO_1303 (O_1303,N_22120,N_22999);
nor UO_1304 (O_1304,N_23216,N_23599);
and UO_1305 (O_1305,N_21953,N_24194);
and UO_1306 (O_1306,N_24460,N_22219);
and UO_1307 (O_1307,N_24121,N_24169);
nor UO_1308 (O_1308,N_23325,N_22652);
or UO_1309 (O_1309,N_23699,N_24507);
xor UO_1310 (O_1310,N_24322,N_24281);
and UO_1311 (O_1311,N_23225,N_22154);
xor UO_1312 (O_1312,N_22463,N_22306);
or UO_1313 (O_1313,N_24920,N_22457);
xnor UO_1314 (O_1314,N_24249,N_23193);
nand UO_1315 (O_1315,N_23332,N_24777);
and UO_1316 (O_1316,N_23811,N_23612);
or UO_1317 (O_1317,N_24004,N_23272);
nor UO_1318 (O_1318,N_23462,N_22156);
and UO_1319 (O_1319,N_21973,N_22445);
nor UO_1320 (O_1320,N_24453,N_23790);
or UO_1321 (O_1321,N_23543,N_24128);
or UO_1322 (O_1322,N_24615,N_22091);
or UO_1323 (O_1323,N_22676,N_22693);
xnor UO_1324 (O_1324,N_22776,N_22281);
nand UO_1325 (O_1325,N_23794,N_24145);
nor UO_1326 (O_1326,N_22392,N_22424);
or UO_1327 (O_1327,N_23600,N_22915);
nand UO_1328 (O_1328,N_22808,N_23347);
or UO_1329 (O_1329,N_24884,N_22518);
and UO_1330 (O_1330,N_23341,N_23192);
nor UO_1331 (O_1331,N_23645,N_23968);
nand UO_1332 (O_1332,N_23574,N_23096);
or UO_1333 (O_1333,N_23080,N_21910);
xor UO_1334 (O_1334,N_23876,N_24935);
or UO_1335 (O_1335,N_22137,N_24980);
nor UO_1336 (O_1336,N_22478,N_24236);
and UO_1337 (O_1337,N_23063,N_23149);
nand UO_1338 (O_1338,N_23438,N_24111);
and UO_1339 (O_1339,N_24562,N_22336);
xor UO_1340 (O_1340,N_23447,N_23959);
or UO_1341 (O_1341,N_23743,N_24693);
and UO_1342 (O_1342,N_24178,N_23260);
nor UO_1343 (O_1343,N_24173,N_22296);
nor UO_1344 (O_1344,N_24605,N_24743);
xor UO_1345 (O_1345,N_23997,N_22222);
and UO_1346 (O_1346,N_23408,N_22194);
nand UO_1347 (O_1347,N_22817,N_23872);
nand UO_1348 (O_1348,N_23506,N_24995);
nand UO_1349 (O_1349,N_24400,N_22149);
nand UO_1350 (O_1350,N_23772,N_24274);
and UO_1351 (O_1351,N_23725,N_23655);
or UO_1352 (O_1352,N_23922,N_23396);
nor UO_1353 (O_1353,N_23093,N_22367);
nor UO_1354 (O_1354,N_23724,N_21879);
and UO_1355 (O_1355,N_22063,N_22841);
and UO_1356 (O_1356,N_22846,N_21891);
nor UO_1357 (O_1357,N_23486,N_22069);
and UO_1358 (O_1358,N_22211,N_23326);
nand UO_1359 (O_1359,N_22579,N_23616);
or UO_1360 (O_1360,N_24946,N_24256);
and UO_1361 (O_1361,N_23432,N_22810);
and UO_1362 (O_1362,N_24100,N_22382);
nor UO_1363 (O_1363,N_24547,N_24378);
nand UO_1364 (O_1364,N_23469,N_23846);
nor UO_1365 (O_1365,N_24251,N_23528);
nand UO_1366 (O_1366,N_23867,N_23951);
or UO_1367 (O_1367,N_23033,N_24785);
or UO_1368 (O_1368,N_23594,N_24987);
xor UO_1369 (O_1369,N_24561,N_24795);
nand UO_1370 (O_1370,N_23513,N_24940);
and UO_1371 (O_1371,N_22804,N_23136);
xor UO_1372 (O_1372,N_23459,N_23604);
nor UO_1373 (O_1373,N_22844,N_22700);
nand UO_1374 (O_1374,N_22514,N_21914);
or UO_1375 (O_1375,N_21984,N_22472);
or UO_1376 (O_1376,N_24006,N_23580);
nor UO_1377 (O_1377,N_22978,N_23467);
nand UO_1378 (O_1378,N_22402,N_24628);
nand UO_1379 (O_1379,N_23776,N_23126);
or UO_1380 (O_1380,N_23521,N_23491);
nand UO_1381 (O_1381,N_24056,N_22558);
and UO_1382 (O_1382,N_22531,N_23511);
and UO_1383 (O_1383,N_22813,N_24261);
nand UO_1384 (O_1384,N_23826,N_23701);
and UO_1385 (O_1385,N_24860,N_23813);
nor UO_1386 (O_1386,N_22790,N_24421);
or UO_1387 (O_1387,N_24969,N_22100);
nor UO_1388 (O_1388,N_22555,N_22362);
nor UO_1389 (O_1389,N_23154,N_23439);
xnor UO_1390 (O_1390,N_21961,N_24713);
and UO_1391 (O_1391,N_22911,N_24797);
nand UO_1392 (O_1392,N_22635,N_24664);
nor UO_1393 (O_1393,N_24470,N_23194);
and UO_1394 (O_1394,N_24239,N_22442);
nand UO_1395 (O_1395,N_21893,N_21896);
and UO_1396 (O_1396,N_24192,N_24029);
or UO_1397 (O_1397,N_24160,N_23632);
nand UO_1398 (O_1398,N_23979,N_23283);
nand UO_1399 (O_1399,N_22974,N_24001);
xor UO_1400 (O_1400,N_23512,N_22387);
or UO_1401 (O_1401,N_22092,N_23905);
nand UO_1402 (O_1402,N_22666,N_24244);
nor UO_1403 (O_1403,N_22654,N_22606);
or UO_1404 (O_1404,N_22022,N_24923);
nor UO_1405 (O_1405,N_24619,N_22907);
or UO_1406 (O_1406,N_22955,N_21989);
or UO_1407 (O_1407,N_22343,N_24624);
nor UO_1408 (O_1408,N_21888,N_22381);
xor UO_1409 (O_1409,N_23700,N_24467);
nor UO_1410 (O_1410,N_22215,N_24383);
nand UO_1411 (O_1411,N_24822,N_22589);
nand UO_1412 (O_1412,N_23731,N_23402);
and UO_1413 (O_1413,N_24568,N_24930);
or UO_1414 (O_1414,N_24063,N_22076);
nor UO_1415 (O_1415,N_23833,N_23387);
and UO_1416 (O_1416,N_24570,N_22899);
and UO_1417 (O_1417,N_22110,N_21935);
nand UO_1418 (O_1418,N_22439,N_23220);
nand UO_1419 (O_1419,N_22592,N_22238);
nand UO_1420 (O_1420,N_24630,N_23748);
and UO_1421 (O_1421,N_24714,N_23297);
and UO_1422 (O_1422,N_22210,N_22513);
nand UO_1423 (O_1423,N_24590,N_24939);
nor UO_1424 (O_1424,N_24341,N_23112);
nand UO_1425 (O_1425,N_23143,N_22129);
and UO_1426 (O_1426,N_22891,N_22174);
and UO_1427 (O_1427,N_22500,N_24208);
xor UO_1428 (O_1428,N_23770,N_23392);
and UO_1429 (O_1429,N_22594,N_23706);
or UO_1430 (O_1430,N_24254,N_24634);
or UO_1431 (O_1431,N_22501,N_23803);
and UO_1432 (O_1432,N_23779,N_23620);
and UO_1433 (O_1433,N_23150,N_22175);
nor UO_1434 (O_1434,N_24734,N_24092);
and UO_1435 (O_1435,N_23043,N_23480);
nor UO_1436 (O_1436,N_24938,N_24015);
and UO_1437 (O_1437,N_24349,N_22743);
or UO_1438 (O_1438,N_22815,N_22605);
nand UO_1439 (O_1439,N_22884,N_24355);
and UO_1440 (O_1440,N_22895,N_24423);
xnor UO_1441 (O_1441,N_24297,N_22425);
nand UO_1442 (O_1442,N_22521,N_21966);
nand UO_1443 (O_1443,N_23729,N_22321);
nor UO_1444 (O_1444,N_23505,N_22784);
and UO_1445 (O_1445,N_22968,N_24358);
and UO_1446 (O_1446,N_24456,N_24185);
nor UO_1447 (O_1447,N_23328,N_24803);
nor UO_1448 (O_1448,N_22553,N_22725);
or UO_1449 (O_1449,N_23179,N_24506);
and UO_1450 (O_1450,N_24982,N_24945);
or UO_1451 (O_1451,N_24882,N_24434);
or UO_1452 (O_1452,N_23137,N_23929);
xor UO_1453 (O_1453,N_23539,N_24018);
or UO_1454 (O_1454,N_23709,N_24248);
xnor UO_1455 (O_1455,N_22273,N_23773);
nand UO_1456 (O_1456,N_22490,N_24326);
and UO_1457 (O_1457,N_24061,N_23767);
xnor UO_1458 (O_1458,N_24432,N_24933);
nor UO_1459 (O_1459,N_24993,N_24728);
nand UO_1460 (O_1460,N_23125,N_22232);
or UO_1461 (O_1461,N_24311,N_23157);
nand UO_1462 (O_1462,N_24479,N_21919);
nor UO_1463 (O_1463,N_24726,N_24682);
or UO_1464 (O_1464,N_23059,N_21982);
and UO_1465 (O_1465,N_23046,N_23690);
nand UO_1466 (O_1466,N_21936,N_23957);
and UO_1467 (O_1467,N_24042,N_24105);
xnor UO_1468 (O_1468,N_21916,N_23906);
nor UO_1469 (O_1469,N_22047,N_23854);
xnor UO_1470 (O_1470,N_22168,N_23585);
nand UO_1471 (O_1471,N_23850,N_24478);
nor UO_1472 (O_1472,N_23841,N_22723);
or UO_1473 (O_1473,N_22540,N_24041);
nor UO_1474 (O_1474,N_23490,N_23334);
nand UO_1475 (O_1475,N_24703,N_22390);
nand UO_1476 (O_1476,N_23280,N_22894);
nand UO_1477 (O_1477,N_24449,N_22548);
nand UO_1478 (O_1478,N_24205,N_21882);
nor UO_1479 (O_1479,N_22155,N_23198);
nand UO_1480 (O_1480,N_22930,N_24885);
nor UO_1481 (O_1481,N_22421,N_21946);
nand UO_1482 (O_1482,N_22216,N_24494);
and UO_1483 (O_1483,N_22740,N_22406);
xor UO_1484 (O_1484,N_22234,N_23156);
xnor UO_1485 (O_1485,N_23378,N_22118);
xnor UO_1486 (O_1486,N_23964,N_23227);
or UO_1487 (O_1487,N_21972,N_23613);
nand UO_1488 (O_1488,N_24632,N_23963);
nand UO_1489 (O_1489,N_24375,N_24135);
and UO_1490 (O_1490,N_23067,N_22462);
and UO_1491 (O_1491,N_22984,N_22423);
nand UO_1492 (O_1492,N_22088,N_23308);
nor UO_1493 (O_1493,N_24784,N_24172);
or UO_1494 (O_1494,N_23733,N_23186);
nand UO_1495 (O_1495,N_21875,N_22269);
nor UO_1496 (O_1496,N_22684,N_24278);
or UO_1497 (O_1497,N_23756,N_23449);
or UO_1498 (O_1498,N_23456,N_22949);
nor UO_1499 (O_1499,N_22431,N_23784);
and UO_1500 (O_1500,N_24911,N_24589);
nor UO_1501 (O_1501,N_23189,N_23888);
and UO_1502 (O_1502,N_21886,N_21912);
nor UO_1503 (O_1503,N_23298,N_22256);
or UO_1504 (O_1504,N_21977,N_23808);
or UO_1505 (O_1505,N_24109,N_23692);
nand UO_1506 (O_1506,N_24512,N_22898);
and UO_1507 (O_1507,N_23777,N_22858);
and UO_1508 (O_1508,N_23578,N_23495);
nand UO_1509 (O_1509,N_23657,N_24577);
nand UO_1510 (O_1510,N_21997,N_22698);
or UO_1511 (O_1511,N_22691,N_24324);
or UO_1512 (O_1512,N_22108,N_22410);
and UO_1513 (O_1513,N_23478,N_24578);
nand UO_1514 (O_1514,N_23953,N_22983);
and UO_1515 (O_1515,N_22773,N_24020);
nand UO_1516 (O_1516,N_23374,N_24863);
and UO_1517 (O_1517,N_23110,N_23281);
or UO_1518 (O_1518,N_23237,N_24569);
or UO_1519 (O_1519,N_22586,N_23871);
and UO_1520 (O_1520,N_23791,N_22035);
nor UO_1521 (O_1521,N_23007,N_23719);
xor UO_1522 (O_1522,N_24198,N_22914);
nor UO_1523 (O_1523,N_23944,N_22370);
or UO_1524 (O_1524,N_22832,N_22697);
nand UO_1525 (O_1525,N_24718,N_23897);
nor UO_1526 (O_1526,N_22641,N_22305);
xnor UO_1527 (O_1527,N_24082,N_23686);
xnor UO_1528 (O_1528,N_23412,N_22357);
and UO_1529 (O_1529,N_23514,N_22196);
nand UO_1530 (O_1530,N_22916,N_24148);
and UO_1531 (O_1531,N_24671,N_24385);
and UO_1532 (O_1532,N_23982,N_24551);
nand UO_1533 (O_1533,N_22409,N_23177);
nand UO_1534 (O_1534,N_23405,N_24504);
or UO_1535 (O_1535,N_24786,N_22568);
or UO_1536 (O_1536,N_22136,N_23597);
nor UO_1537 (O_1537,N_24754,N_24306);
nor UO_1538 (O_1538,N_22000,N_24659);
and UO_1539 (O_1539,N_24327,N_23320);
xnor UO_1540 (O_1540,N_22345,N_24963);
xor UO_1541 (O_1541,N_24813,N_22106);
or UO_1542 (O_1542,N_22596,N_22843);
or UO_1543 (O_1543,N_23617,N_24543);
nor UO_1544 (O_1544,N_23839,N_22351);
xor UO_1545 (O_1545,N_24525,N_23333);
and UO_1546 (O_1546,N_22068,N_24622);
or UO_1547 (O_1547,N_22865,N_24618);
and UO_1548 (O_1548,N_23292,N_22014);
nand UO_1549 (O_1549,N_23806,N_24540);
and UO_1550 (O_1550,N_22481,N_22240);
nor UO_1551 (O_1551,N_22538,N_24511);
or UO_1552 (O_1552,N_24952,N_24757);
nor UO_1553 (O_1553,N_24014,N_22405);
nor UO_1554 (O_1554,N_23631,N_22459);
nor UO_1555 (O_1555,N_23338,N_22026);
or UO_1556 (O_1556,N_23946,N_23648);
nor UO_1557 (O_1557,N_23693,N_23255);
and UO_1558 (O_1558,N_24357,N_23948);
nor UO_1559 (O_1559,N_21964,N_24089);
and UO_1560 (O_1560,N_23346,N_22545);
nor UO_1561 (O_1561,N_24259,N_22774);
nand UO_1562 (O_1562,N_21902,N_22379);
and UO_1563 (O_1563,N_24596,N_24385);
and UO_1564 (O_1564,N_22191,N_22550);
nor UO_1565 (O_1565,N_22396,N_22186);
nor UO_1566 (O_1566,N_23920,N_24429);
or UO_1567 (O_1567,N_22019,N_22405);
xnor UO_1568 (O_1568,N_24635,N_24067);
and UO_1569 (O_1569,N_24392,N_23113);
or UO_1570 (O_1570,N_22917,N_24848);
nor UO_1571 (O_1571,N_24887,N_22535);
and UO_1572 (O_1572,N_23257,N_23068);
and UO_1573 (O_1573,N_22806,N_22877);
nand UO_1574 (O_1574,N_24860,N_21912);
or UO_1575 (O_1575,N_24362,N_22468);
nand UO_1576 (O_1576,N_24787,N_22087);
and UO_1577 (O_1577,N_22032,N_23890);
nand UO_1578 (O_1578,N_22248,N_23457);
xor UO_1579 (O_1579,N_24559,N_24585);
or UO_1580 (O_1580,N_24141,N_24401);
and UO_1581 (O_1581,N_23059,N_23082);
nand UO_1582 (O_1582,N_22286,N_22322);
nor UO_1583 (O_1583,N_24435,N_24934);
or UO_1584 (O_1584,N_22133,N_22063);
and UO_1585 (O_1585,N_22437,N_23842);
nor UO_1586 (O_1586,N_23244,N_22381);
xor UO_1587 (O_1587,N_24121,N_23535);
nand UO_1588 (O_1588,N_22003,N_22785);
or UO_1589 (O_1589,N_24488,N_23603);
nand UO_1590 (O_1590,N_22478,N_24369);
or UO_1591 (O_1591,N_24385,N_24152);
nor UO_1592 (O_1592,N_22417,N_22653);
and UO_1593 (O_1593,N_23317,N_24215);
and UO_1594 (O_1594,N_24656,N_21890);
or UO_1595 (O_1595,N_22738,N_24546);
or UO_1596 (O_1596,N_22523,N_24990);
nand UO_1597 (O_1597,N_22773,N_23590);
nor UO_1598 (O_1598,N_23762,N_24915);
or UO_1599 (O_1599,N_24878,N_22886);
nor UO_1600 (O_1600,N_22162,N_23028);
and UO_1601 (O_1601,N_23891,N_22252);
nand UO_1602 (O_1602,N_23807,N_23662);
nor UO_1603 (O_1603,N_22592,N_22729);
or UO_1604 (O_1604,N_22769,N_23533);
and UO_1605 (O_1605,N_24841,N_24993);
nor UO_1606 (O_1606,N_22752,N_21999);
xor UO_1607 (O_1607,N_22136,N_24275);
nand UO_1608 (O_1608,N_22515,N_24370);
nor UO_1609 (O_1609,N_24341,N_22611);
xor UO_1610 (O_1610,N_24197,N_22192);
or UO_1611 (O_1611,N_22720,N_24186);
xor UO_1612 (O_1612,N_22168,N_22074);
and UO_1613 (O_1613,N_21891,N_23260);
nand UO_1614 (O_1614,N_23401,N_23394);
nand UO_1615 (O_1615,N_22746,N_22284);
and UO_1616 (O_1616,N_24896,N_23773);
or UO_1617 (O_1617,N_22981,N_24911);
nand UO_1618 (O_1618,N_23231,N_24437);
or UO_1619 (O_1619,N_24239,N_22662);
nor UO_1620 (O_1620,N_23508,N_24313);
nand UO_1621 (O_1621,N_24205,N_24068);
or UO_1622 (O_1622,N_23812,N_24608);
nand UO_1623 (O_1623,N_22600,N_24906);
and UO_1624 (O_1624,N_21887,N_24147);
and UO_1625 (O_1625,N_24288,N_22475);
or UO_1626 (O_1626,N_23979,N_24029);
nand UO_1627 (O_1627,N_22516,N_23784);
or UO_1628 (O_1628,N_22645,N_22852);
nand UO_1629 (O_1629,N_23448,N_24509);
and UO_1630 (O_1630,N_23650,N_23137);
nor UO_1631 (O_1631,N_22564,N_22785);
or UO_1632 (O_1632,N_22936,N_22213);
xnor UO_1633 (O_1633,N_22952,N_23950);
or UO_1634 (O_1634,N_24096,N_22897);
or UO_1635 (O_1635,N_22792,N_22286);
or UO_1636 (O_1636,N_23029,N_22361);
nand UO_1637 (O_1637,N_23834,N_23966);
nand UO_1638 (O_1638,N_24942,N_23914);
nor UO_1639 (O_1639,N_24259,N_23429);
and UO_1640 (O_1640,N_22735,N_22790);
and UO_1641 (O_1641,N_23689,N_22860);
nor UO_1642 (O_1642,N_22065,N_22979);
nor UO_1643 (O_1643,N_24884,N_21969);
nor UO_1644 (O_1644,N_23303,N_24303);
and UO_1645 (O_1645,N_24562,N_24310);
xnor UO_1646 (O_1646,N_22498,N_23494);
nor UO_1647 (O_1647,N_24556,N_23894);
or UO_1648 (O_1648,N_23916,N_22390);
nor UO_1649 (O_1649,N_24690,N_23802);
and UO_1650 (O_1650,N_23129,N_22451);
or UO_1651 (O_1651,N_24355,N_24457);
nor UO_1652 (O_1652,N_23244,N_24358);
and UO_1653 (O_1653,N_22978,N_22607);
or UO_1654 (O_1654,N_22775,N_24538);
or UO_1655 (O_1655,N_23944,N_24729);
and UO_1656 (O_1656,N_22648,N_23424);
nand UO_1657 (O_1657,N_24550,N_24912);
nor UO_1658 (O_1658,N_23991,N_22793);
and UO_1659 (O_1659,N_22660,N_23378);
or UO_1660 (O_1660,N_23548,N_24879);
and UO_1661 (O_1661,N_22967,N_21913);
nor UO_1662 (O_1662,N_21996,N_23761);
nand UO_1663 (O_1663,N_23531,N_23662);
and UO_1664 (O_1664,N_22783,N_24443);
and UO_1665 (O_1665,N_22192,N_24030);
or UO_1666 (O_1666,N_23214,N_23854);
xor UO_1667 (O_1667,N_22802,N_22842);
nor UO_1668 (O_1668,N_24795,N_23043);
nor UO_1669 (O_1669,N_24852,N_21906);
and UO_1670 (O_1670,N_23954,N_24523);
or UO_1671 (O_1671,N_23026,N_23367);
or UO_1672 (O_1672,N_23126,N_24149);
or UO_1673 (O_1673,N_21945,N_22791);
or UO_1674 (O_1674,N_21920,N_22870);
nand UO_1675 (O_1675,N_23594,N_24274);
nand UO_1676 (O_1676,N_22614,N_24770);
nand UO_1677 (O_1677,N_24621,N_22344);
and UO_1678 (O_1678,N_22998,N_24966);
and UO_1679 (O_1679,N_22179,N_22711);
nor UO_1680 (O_1680,N_23545,N_24896);
or UO_1681 (O_1681,N_22149,N_24976);
nor UO_1682 (O_1682,N_24425,N_23594);
nor UO_1683 (O_1683,N_24947,N_22629);
or UO_1684 (O_1684,N_23774,N_22611);
and UO_1685 (O_1685,N_23206,N_24542);
nor UO_1686 (O_1686,N_22953,N_22877);
nor UO_1687 (O_1687,N_24926,N_22363);
nand UO_1688 (O_1688,N_24499,N_22449);
nand UO_1689 (O_1689,N_24094,N_24590);
xnor UO_1690 (O_1690,N_22791,N_22303);
nand UO_1691 (O_1691,N_22699,N_23066);
and UO_1692 (O_1692,N_24018,N_23862);
or UO_1693 (O_1693,N_23306,N_23384);
nor UO_1694 (O_1694,N_24594,N_22600);
and UO_1695 (O_1695,N_23106,N_24713);
nor UO_1696 (O_1696,N_23733,N_23383);
and UO_1697 (O_1697,N_23024,N_23837);
or UO_1698 (O_1698,N_22930,N_22881);
and UO_1699 (O_1699,N_23548,N_22331);
or UO_1700 (O_1700,N_23570,N_23237);
xnor UO_1701 (O_1701,N_24430,N_24810);
xnor UO_1702 (O_1702,N_21936,N_23704);
nand UO_1703 (O_1703,N_24957,N_23349);
nor UO_1704 (O_1704,N_22748,N_22003);
nor UO_1705 (O_1705,N_24157,N_24292);
nor UO_1706 (O_1706,N_22444,N_24361);
and UO_1707 (O_1707,N_24271,N_22022);
or UO_1708 (O_1708,N_21971,N_24386);
or UO_1709 (O_1709,N_23274,N_24441);
or UO_1710 (O_1710,N_23887,N_23639);
or UO_1711 (O_1711,N_24064,N_22206);
nand UO_1712 (O_1712,N_22473,N_24985);
or UO_1713 (O_1713,N_23803,N_23346);
nand UO_1714 (O_1714,N_23240,N_23977);
xnor UO_1715 (O_1715,N_22471,N_23997);
nand UO_1716 (O_1716,N_23679,N_22610);
nand UO_1717 (O_1717,N_23683,N_24990);
and UO_1718 (O_1718,N_22259,N_24674);
and UO_1719 (O_1719,N_24392,N_22982);
and UO_1720 (O_1720,N_23191,N_23883);
or UO_1721 (O_1721,N_23835,N_22956);
nor UO_1722 (O_1722,N_22498,N_24057);
nor UO_1723 (O_1723,N_22125,N_24895);
xor UO_1724 (O_1724,N_24751,N_23374);
and UO_1725 (O_1725,N_24347,N_22345);
nand UO_1726 (O_1726,N_24488,N_23143);
nand UO_1727 (O_1727,N_22233,N_24336);
nor UO_1728 (O_1728,N_22434,N_22412);
or UO_1729 (O_1729,N_24896,N_23750);
nor UO_1730 (O_1730,N_23395,N_23153);
nor UO_1731 (O_1731,N_23861,N_22255);
nand UO_1732 (O_1732,N_23244,N_22851);
nor UO_1733 (O_1733,N_22578,N_21940);
nand UO_1734 (O_1734,N_24143,N_23727);
and UO_1735 (O_1735,N_23129,N_23265);
and UO_1736 (O_1736,N_24205,N_24329);
or UO_1737 (O_1737,N_24503,N_24589);
nand UO_1738 (O_1738,N_22737,N_24852);
nand UO_1739 (O_1739,N_24821,N_22496);
nand UO_1740 (O_1740,N_24560,N_21931);
nand UO_1741 (O_1741,N_23275,N_22531);
nor UO_1742 (O_1742,N_24242,N_24969);
nand UO_1743 (O_1743,N_24018,N_22866);
and UO_1744 (O_1744,N_23620,N_22489);
and UO_1745 (O_1745,N_23127,N_23452);
or UO_1746 (O_1746,N_24786,N_22077);
or UO_1747 (O_1747,N_21895,N_24806);
nand UO_1748 (O_1748,N_24821,N_24956);
nor UO_1749 (O_1749,N_22177,N_24092);
nor UO_1750 (O_1750,N_24389,N_22527);
nor UO_1751 (O_1751,N_24800,N_24732);
xor UO_1752 (O_1752,N_22965,N_22073);
nand UO_1753 (O_1753,N_22802,N_22039);
xnor UO_1754 (O_1754,N_23335,N_23683);
xnor UO_1755 (O_1755,N_24924,N_24560);
or UO_1756 (O_1756,N_23156,N_23061);
nor UO_1757 (O_1757,N_22353,N_23074);
or UO_1758 (O_1758,N_24465,N_22599);
and UO_1759 (O_1759,N_23868,N_22459);
or UO_1760 (O_1760,N_23516,N_23278);
or UO_1761 (O_1761,N_22661,N_23003);
or UO_1762 (O_1762,N_23232,N_22320);
nand UO_1763 (O_1763,N_22900,N_23120);
or UO_1764 (O_1764,N_23188,N_24285);
nand UO_1765 (O_1765,N_21919,N_22642);
nor UO_1766 (O_1766,N_24573,N_23751);
xnor UO_1767 (O_1767,N_23272,N_22782);
nand UO_1768 (O_1768,N_24617,N_23519);
or UO_1769 (O_1769,N_23360,N_22156);
and UO_1770 (O_1770,N_22180,N_24754);
nand UO_1771 (O_1771,N_22066,N_23707);
nor UO_1772 (O_1772,N_22383,N_22727);
and UO_1773 (O_1773,N_24050,N_23216);
or UO_1774 (O_1774,N_23121,N_22118);
and UO_1775 (O_1775,N_23018,N_22609);
nor UO_1776 (O_1776,N_23362,N_22600);
nand UO_1777 (O_1777,N_23961,N_22828);
nand UO_1778 (O_1778,N_24170,N_23564);
or UO_1779 (O_1779,N_23201,N_24200);
or UO_1780 (O_1780,N_22868,N_23418);
nor UO_1781 (O_1781,N_24751,N_24439);
xor UO_1782 (O_1782,N_21880,N_22911);
and UO_1783 (O_1783,N_23115,N_23205);
nor UO_1784 (O_1784,N_24752,N_23228);
or UO_1785 (O_1785,N_24747,N_23622);
nand UO_1786 (O_1786,N_23282,N_23417);
nand UO_1787 (O_1787,N_21995,N_22118);
nor UO_1788 (O_1788,N_24939,N_21949);
and UO_1789 (O_1789,N_22099,N_22872);
nor UO_1790 (O_1790,N_24445,N_22257);
or UO_1791 (O_1791,N_23219,N_23297);
nand UO_1792 (O_1792,N_22445,N_22618);
nand UO_1793 (O_1793,N_22959,N_23370);
or UO_1794 (O_1794,N_24178,N_24538);
or UO_1795 (O_1795,N_22220,N_24621);
or UO_1796 (O_1796,N_24027,N_24684);
and UO_1797 (O_1797,N_24280,N_21896);
xnor UO_1798 (O_1798,N_23715,N_24767);
nand UO_1799 (O_1799,N_24834,N_22565);
xor UO_1800 (O_1800,N_22059,N_24777);
nand UO_1801 (O_1801,N_22118,N_22753);
or UO_1802 (O_1802,N_24628,N_24476);
nand UO_1803 (O_1803,N_22898,N_22495);
and UO_1804 (O_1804,N_22699,N_23672);
nor UO_1805 (O_1805,N_24225,N_22231);
nor UO_1806 (O_1806,N_22694,N_22872);
nor UO_1807 (O_1807,N_22625,N_23353);
nor UO_1808 (O_1808,N_24872,N_24328);
or UO_1809 (O_1809,N_24181,N_22280);
and UO_1810 (O_1810,N_23268,N_24313);
and UO_1811 (O_1811,N_23574,N_22942);
nand UO_1812 (O_1812,N_22254,N_24057);
nor UO_1813 (O_1813,N_22913,N_23870);
xor UO_1814 (O_1814,N_22967,N_23288);
and UO_1815 (O_1815,N_21926,N_24830);
or UO_1816 (O_1816,N_22696,N_24289);
and UO_1817 (O_1817,N_24737,N_24632);
nand UO_1818 (O_1818,N_23354,N_24843);
xor UO_1819 (O_1819,N_22498,N_22245);
and UO_1820 (O_1820,N_22197,N_22878);
nand UO_1821 (O_1821,N_24337,N_22180);
or UO_1822 (O_1822,N_24586,N_22186);
nand UO_1823 (O_1823,N_22500,N_24992);
nor UO_1824 (O_1824,N_24730,N_22965);
or UO_1825 (O_1825,N_22785,N_24558);
nand UO_1826 (O_1826,N_23846,N_23589);
xnor UO_1827 (O_1827,N_24603,N_23844);
and UO_1828 (O_1828,N_22040,N_23515);
nand UO_1829 (O_1829,N_22387,N_24771);
nor UO_1830 (O_1830,N_23705,N_22452);
nand UO_1831 (O_1831,N_24158,N_24647);
xor UO_1832 (O_1832,N_23044,N_23255);
or UO_1833 (O_1833,N_23762,N_22891);
xnor UO_1834 (O_1834,N_23979,N_23943);
or UO_1835 (O_1835,N_23152,N_24450);
or UO_1836 (O_1836,N_23756,N_24379);
xor UO_1837 (O_1837,N_23752,N_23318);
or UO_1838 (O_1838,N_23363,N_24810);
or UO_1839 (O_1839,N_24510,N_24797);
nor UO_1840 (O_1840,N_24655,N_23201);
nor UO_1841 (O_1841,N_22294,N_23823);
and UO_1842 (O_1842,N_24302,N_23154);
nand UO_1843 (O_1843,N_24294,N_23668);
or UO_1844 (O_1844,N_22715,N_22777);
and UO_1845 (O_1845,N_22421,N_24074);
or UO_1846 (O_1846,N_23342,N_22005);
nand UO_1847 (O_1847,N_23525,N_22014);
xnor UO_1848 (O_1848,N_21927,N_21887);
nand UO_1849 (O_1849,N_24126,N_22416);
nand UO_1850 (O_1850,N_23580,N_24019);
nor UO_1851 (O_1851,N_22440,N_22357);
or UO_1852 (O_1852,N_24755,N_23049);
or UO_1853 (O_1853,N_22519,N_22166);
xor UO_1854 (O_1854,N_22328,N_22290);
nand UO_1855 (O_1855,N_24734,N_24323);
nor UO_1856 (O_1856,N_22093,N_22327);
or UO_1857 (O_1857,N_24247,N_24827);
or UO_1858 (O_1858,N_23940,N_24764);
or UO_1859 (O_1859,N_23286,N_21977);
nor UO_1860 (O_1860,N_24924,N_23417);
or UO_1861 (O_1861,N_24967,N_22952);
xor UO_1862 (O_1862,N_22958,N_22661);
and UO_1863 (O_1863,N_22971,N_24730);
or UO_1864 (O_1864,N_21959,N_23845);
nor UO_1865 (O_1865,N_24352,N_24783);
xnor UO_1866 (O_1866,N_22065,N_23590);
or UO_1867 (O_1867,N_24229,N_23322);
nor UO_1868 (O_1868,N_22387,N_23830);
nor UO_1869 (O_1869,N_22209,N_23857);
xnor UO_1870 (O_1870,N_22167,N_22877);
nor UO_1871 (O_1871,N_23541,N_24808);
nand UO_1872 (O_1872,N_23474,N_21992);
nand UO_1873 (O_1873,N_23006,N_23417);
and UO_1874 (O_1874,N_22074,N_21936);
xnor UO_1875 (O_1875,N_22072,N_24688);
xnor UO_1876 (O_1876,N_23464,N_23886);
nor UO_1877 (O_1877,N_23399,N_22483);
or UO_1878 (O_1878,N_22373,N_21886);
nand UO_1879 (O_1879,N_23551,N_22205);
and UO_1880 (O_1880,N_23022,N_23153);
or UO_1881 (O_1881,N_24413,N_24991);
nand UO_1882 (O_1882,N_24617,N_24814);
nor UO_1883 (O_1883,N_22965,N_22842);
xnor UO_1884 (O_1884,N_24921,N_22198);
or UO_1885 (O_1885,N_24265,N_24456);
xor UO_1886 (O_1886,N_24597,N_23363);
nand UO_1887 (O_1887,N_23596,N_24657);
nor UO_1888 (O_1888,N_23686,N_23786);
xor UO_1889 (O_1889,N_23862,N_24651);
nor UO_1890 (O_1890,N_24068,N_23799);
nand UO_1891 (O_1891,N_22938,N_24523);
or UO_1892 (O_1892,N_22238,N_22141);
nand UO_1893 (O_1893,N_22151,N_23872);
and UO_1894 (O_1894,N_23751,N_22979);
and UO_1895 (O_1895,N_24145,N_23692);
nor UO_1896 (O_1896,N_23628,N_22063);
or UO_1897 (O_1897,N_24971,N_22606);
nor UO_1898 (O_1898,N_24942,N_22603);
nor UO_1899 (O_1899,N_21989,N_24299);
xnor UO_1900 (O_1900,N_23502,N_23802);
or UO_1901 (O_1901,N_24147,N_24470);
or UO_1902 (O_1902,N_23064,N_23699);
nor UO_1903 (O_1903,N_23545,N_23108);
or UO_1904 (O_1904,N_23001,N_23290);
or UO_1905 (O_1905,N_23918,N_24218);
xnor UO_1906 (O_1906,N_22877,N_24284);
and UO_1907 (O_1907,N_22882,N_22943);
xnor UO_1908 (O_1908,N_22266,N_23792);
nor UO_1909 (O_1909,N_21882,N_22362);
xnor UO_1910 (O_1910,N_22811,N_22213);
nand UO_1911 (O_1911,N_24401,N_24308);
and UO_1912 (O_1912,N_24963,N_22485);
or UO_1913 (O_1913,N_24512,N_22757);
and UO_1914 (O_1914,N_24760,N_24208);
nor UO_1915 (O_1915,N_23359,N_22773);
nand UO_1916 (O_1916,N_23278,N_21955);
or UO_1917 (O_1917,N_24705,N_24440);
nand UO_1918 (O_1918,N_22467,N_22602);
nor UO_1919 (O_1919,N_23154,N_24535);
or UO_1920 (O_1920,N_23808,N_24688);
xnor UO_1921 (O_1921,N_24406,N_24798);
and UO_1922 (O_1922,N_24645,N_22558);
nor UO_1923 (O_1923,N_22052,N_24275);
and UO_1924 (O_1924,N_22900,N_23629);
nor UO_1925 (O_1925,N_22336,N_24250);
nand UO_1926 (O_1926,N_23667,N_24672);
nor UO_1927 (O_1927,N_23071,N_22425);
nor UO_1928 (O_1928,N_24640,N_23414);
and UO_1929 (O_1929,N_24715,N_23079);
nand UO_1930 (O_1930,N_23052,N_23469);
or UO_1931 (O_1931,N_23909,N_22983);
and UO_1932 (O_1932,N_22580,N_23990);
and UO_1933 (O_1933,N_22974,N_24533);
or UO_1934 (O_1934,N_24264,N_22658);
and UO_1935 (O_1935,N_24819,N_24418);
nor UO_1936 (O_1936,N_23771,N_23343);
and UO_1937 (O_1937,N_23982,N_22091);
xnor UO_1938 (O_1938,N_23510,N_24178);
nor UO_1939 (O_1939,N_21993,N_24179);
nor UO_1940 (O_1940,N_24661,N_24891);
nand UO_1941 (O_1941,N_22317,N_24670);
nand UO_1942 (O_1942,N_23738,N_24048);
and UO_1943 (O_1943,N_22221,N_24428);
xnor UO_1944 (O_1944,N_22290,N_23931);
and UO_1945 (O_1945,N_23937,N_23169);
or UO_1946 (O_1946,N_23088,N_22001);
or UO_1947 (O_1947,N_21940,N_22652);
nand UO_1948 (O_1948,N_24752,N_24918);
nor UO_1949 (O_1949,N_23890,N_23710);
nor UO_1950 (O_1950,N_23457,N_24607);
and UO_1951 (O_1951,N_23708,N_24079);
or UO_1952 (O_1952,N_23672,N_22806);
nand UO_1953 (O_1953,N_22772,N_22735);
xor UO_1954 (O_1954,N_24281,N_22319);
nor UO_1955 (O_1955,N_24290,N_22412);
nor UO_1956 (O_1956,N_23637,N_22518);
or UO_1957 (O_1957,N_22182,N_22586);
xor UO_1958 (O_1958,N_22985,N_23117);
or UO_1959 (O_1959,N_24002,N_24569);
and UO_1960 (O_1960,N_24527,N_23563);
nor UO_1961 (O_1961,N_22193,N_21998);
and UO_1962 (O_1962,N_24341,N_24639);
nand UO_1963 (O_1963,N_24348,N_24763);
nand UO_1964 (O_1964,N_23594,N_22905);
or UO_1965 (O_1965,N_24796,N_21954);
and UO_1966 (O_1966,N_22404,N_24837);
or UO_1967 (O_1967,N_24865,N_24034);
or UO_1968 (O_1968,N_24279,N_22337);
nor UO_1969 (O_1969,N_22897,N_24641);
nor UO_1970 (O_1970,N_23194,N_24103);
nor UO_1971 (O_1971,N_23080,N_24272);
nand UO_1972 (O_1972,N_24963,N_24849);
and UO_1973 (O_1973,N_23205,N_23437);
and UO_1974 (O_1974,N_24105,N_23222);
or UO_1975 (O_1975,N_23363,N_22826);
xor UO_1976 (O_1976,N_23087,N_24018);
nand UO_1977 (O_1977,N_23483,N_23916);
nor UO_1978 (O_1978,N_24602,N_23218);
nand UO_1979 (O_1979,N_23163,N_22759);
nor UO_1980 (O_1980,N_24012,N_23474);
nand UO_1981 (O_1981,N_21917,N_22895);
nor UO_1982 (O_1982,N_23074,N_22313);
or UO_1983 (O_1983,N_22439,N_23374);
nand UO_1984 (O_1984,N_23172,N_23588);
xnor UO_1985 (O_1985,N_23943,N_21945);
nand UO_1986 (O_1986,N_22113,N_22821);
and UO_1987 (O_1987,N_23386,N_24758);
and UO_1988 (O_1988,N_22817,N_23991);
and UO_1989 (O_1989,N_24712,N_23750);
and UO_1990 (O_1990,N_24949,N_22502);
nand UO_1991 (O_1991,N_23655,N_22704);
and UO_1992 (O_1992,N_23068,N_24309);
and UO_1993 (O_1993,N_24400,N_24780);
or UO_1994 (O_1994,N_23664,N_21959);
nand UO_1995 (O_1995,N_23524,N_22991);
or UO_1996 (O_1996,N_22778,N_24283);
and UO_1997 (O_1997,N_22904,N_23500);
nor UO_1998 (O_1998,N_23447,N_21965);
nor UO_1999 (O_1999,N_22632,N_21889);
nand UO_2000 (O_2000,N_23095,N_23283);
nor UO_2001 (O_2001,N_22948,N_23939);
nor UO_2002 (O_2002,N_24833,N_24648);
nand UO_2003 (O_2003,N_22989,N_24169);
or UO_2004 (O_2004,N_24059,N_22915);
or UO_2005 (O_2005,N_24004,N_22136);
nor UO_2006 (O_2006,N_24442,N_24684);
nor UO_2007 (O_2007,N_22394,N_21895);
nor UO_2008 (O_2008,N_22735,N_22870);
nor UO_2009 (O_2009,N_22742,N_24302);
and UO_2010 (O_2010,N_23605,N_23930);
or UO_2011 (O_2011,N_24841,N_22497);
and UO_2012 (O_2012,N_24071,N_23916);
and UO_2013 (O_2013,N_23865,N_22436);
nand UO_2014 (O_2014,N_21900,N_22360);
nor UO_2015 (O_2015,N_22441,N_24558);
nor UO_2016 (O_2016,N_24008,N_23344);
and UO_2017 (O_2017,N_24793,N_23494);
nand UO_2018 (O_2018,N_24962,N_23631);
nor UO_2019 (O_2019,N_22739,N_23049);
nor UO_2020 (O_2020,N_22647,N_24881);
and UO_2021 (O_2021,N_23176,N_22665);
or UO_2022 (O_2022,N_22939,N_23681);
nor UO_2023 (O_2023,N_24376,N_22570);
xor UO_2024 (O_2024,N_23594,N_22657);
and UO_2025 (O_2025,N_22643,N_23916);
or UO_2026 (O_2026,N_22239,N_24417);
or UO_2027 (O_2027,N_23357,N_24147);
or UO_2028 (O_2028,N_23079,N_22948);
nand UO_2029 (O_2029,N_23274,N_23640);
nand UO_2030 (O_2030,N_22192,N_22734);
xor UO_2031 (O_2031,N_22841,N_23275);
nor UO_2032 (O_2032,N_22948,N_24876);
and UO_2033 (O_2033,N_23489,N_23399);
nand UO_2034 (O_2034,N_22281,N_23922);
nand UO_2035 (O_2035,N_23777,N_22302);
and UO_2036 (O_2036,N_22923,N_23917);
or UO_2037 (O_2037,N_22845,N_23893);
and UO_2038 (O_2038,N_23670,N_22736);
nand UO_2039 (O_2039,N_22174,N_23191);
or UO_2040 (O_2040,N_23661,N_24957);
or UO_2041 (O_2041,N_24106,N_24943);
nand UO_2042 (O_2042,N_23944,N_24156);
xor UO_2043 (O_2043,N_23242,N_23003);
or UO_2044 (O_2044,N_22088,N_24226);
and UO_2045 (O_2045,N_21994,N_22745);
nand UO_2046 (O_2046,N_24353,N_24177);
or UO_2047 (O_2047,N_23077,N_21926);
nand UO_2048 (O_2048,N_23954,N_23138);
nand UO_2049 (O_2049,N_21948,N_24411);
or UO_2050 (O_2050,N_22003,N_23267);
or UO_2051 (O_2051,N_22824,N_23532);
and UO_2052 (O_2052,N_24096,N_22433);
xor UO_2053 (O_2053,N_23241,N_24903);
and UO_2054 (O_2054,N_24459,N_22939);
and UO_2055 (O_2055,N_23927,N_24628);
xor UO_2056 (O_2056,N_23867,N_23025);
or UO_2057 (O_2057,N_24576,N_23329);
nand UO_2058 (O_2058,N_22402,N_23890);
nor UO_2059 (O_2059,N_21959,N_21955);
nor UO_2060 (O_2060,N_23159,N_22044);
and UO_2061 (O_2061,N_23134,N_22635);
or UO_2062 (O_2062,N_22536,N_24523);
and UO_2063 (O_2063,N_22723,N_22066);
and UO_2064 (O_2064,N_23764,N_23010);
or UO_2065 (O_2065,N_22414,N_24669);
and UO_2066 (O_2066,N_23894,N_22805);
nand UO_2067 (O_2067,N_22661,N_24958);
nand UO_2068 (O_2068,N_23784,N_23412);
and UO_2069 (O_2069,N_24022,N_24393);
or UO_2070 (O_2070,N_24970,N_24053);
or UO_2071 (O_2071,N_24537,N_23878);
nor UO_2072 (O_2072,N_23350,N_24340);
or UO_2073 (O_2073,N_24764,N_23763);
or UO_2074 (O_2074,N_22657,N_22382);
nor UO_2075 (O_2075,N_22995,N_24180);
xor UO_2076 (O_2076,N_22989,N_23154);
and UO_2077 (O_2077,N_23404,N_22095);
nand UO_2078 (O_2078,N_22439,N_24485);
or UO_2079 (O_2079,N_23657,N_24311);
and UO_2080 (O_2080,N_23519,N_22081);
nand UO_2081 (O_2081,N_24107,N_23407);
nor UO_2082 (O_2082,N_23683,N_23134);
nor UO_2083 (O_2083,N_22624,N_23366);
nor UO_2084 (O_2084,N_23216,N_23158);
and UO_2085 (O_2085,N_22324,N_22118);
nor UO_2086 (O_2086,N_23062,N_23331);
and UO_2087 (O_2087,N_24179,N_22662);
nand UO_2088 (O_2088,N_23645,N_22917);
or UO_2089 (O_2089,N_23931,N_24174);
nand UO_2090 (O_2090,N_23017,N_23651);
nand UO_2091 (O_2091,N_22227,N_22279);
nor UO_2092 (O_2092,N_23363,N_23380);
nor UO_2093 (O_2093,N_23738,N_23198);
and UO_2094 (O_2094,N_22990,N_22178);
and UO_2095 (O_2095,N_22688,N_23327);
xnor UO_2096 (O_2096,N_24259,N_24806);
or UO_2097 (O_2097,N_22030,N_23991);
or UO_2098 (O_2098,N_22047,N_22819);
xnor UO_2099 (O_2099,N_23314,N_22919);
nand UO_2100 (O_2100,N_23370,N_22128);
nor UO_2101 (O_2101,N_24144,N_22921);
or UO_2102 (O_2102,N_22718,N_23282);
nand UO_2103 (O_2103,N_23782,N_23582);
nor UO_2104 (O_2104,N_23176,N_24253);
nor UO_2105 (O_2105,N_22439,N_23623);
xnor UO_2106 (O_2106,N_23336,N_22732);
or UO_2107 (O_2107,N_23309,N_23171);
nor UO_2108 (O_2108,N_22965,N_22490);
and UO_2109 (O_2109,N_24473,N_23484);
and UO_2110 (O_2110,N_22040,N_22870);
nor UO_2111 (O_2111,N_24072,N_22638);
nand UO_2112 (O_2112,N_24172,N_22948);
nand UO_2113 (O_2113,N_24063,N_22528);
or UO_2114 (O_2114,N_22664,N_24456);
xnor UO_2115 (O_2115,N_24531,N_23013);
nor UO_2116 (O_2116,N_24418,N_23708);
xor UO_2117 (O_2117,N_23464,N_22987);
nor UO_2118 (O_2118,N_24539,N_24577);
xnor UO_2119 (O_2119,N_24210,N_23115);
nor UO_2120 (O_2120,N_24624,N_24969);
nor UO_2121 (O_2121,N_24198,N_24621);
or UO_2122 (O_2122,N_23235,N_22368);
or UO_2123 (O_2123,N_23653,N_23872);
or UO_2124 (O_2124,N_23393,N_24557);
and UO_2125 (O_2125,N_23688,N_23266);
nor UO_2126 (O_2126,N_24140,N_22213);
nor UO_2127 (O_2127,N_24661,N_23699);
nor UO_2128 (O_2128,N_23678,N_24017);
or UO_2129 (O_2129,N_24741,N_22216);
and UO_2130 (O_2130,N_23849,N_23478);
nor UO_2131 (O_2131,N_22707,N_22784);
xor UO_2132 (O_2132,N_23901,N_22872);
nand UO_2133 (O_2133,N_21878,N_23160);
nor UO_2134 (O_2134,N_23187,N_22957);
nand UO_2135 (O_2135,N_24995,N_23557);
nand UO_2136 (O_2136,N_23830,N_22989);
and UO_2137 (O_2137,N_22758,N_23987);
or UO_2138 (O_2138,N_24835,N_24358);
or UO_2139 (O_2139,N_22283,N_24379);
xor UO_2140 (O_2140,N_24935,N_22161);
or UO_2141 (O_2141,N_22611,N_24769);
and UO_2142 (O_2142,N_23614,N_24120);
and UO_2143 (O_2143,N_24870,N_22962);
xor UO_2144 (O_2144,N_22411,N_24773);
nand UO_2145 (O_2145,N_23805,N_22064);
xor UO_2146 (O_2146,N_22918,N_22216);
nor UO_2147 (O_2147,N_23987,N_23824);
and UO_2148 (O_2148,N_24882,N_23468);
nand UO_2149 (O_2149,N_22512,N_24910);
or UO_2150 (O_2150,N_24723,N_22990);
and UO_2151 (O_2151,N_23985,N_24637);
and UO_2152 (O_2152,N_22807,N_22598);
nor UO_2153 (O_2153,N_23740,N_23357);
or UO_2154 (O_2154,N_23406,N_22364);
or UO_2155 (O_2155,N_23976,N_22372);
or UO_2156 (O_2156,N_22290,N_22253);
and UO_2157 (O_2157,N_22219,N_22708);
or UO_2158 (O_2158,N_24443,N_23124);
or UO_2159 (O_2159,N_23932,N_23280);
and UO_2160 (O_2160,N_22632,N_22513);
and UO_2161 (O_2161,N_24935,N_24086);
xor UO_2162 (O_2162,N_23856,N_22922);
or UO_2163 (O_2163,N_22776,N_22333);
nor UO_2164 (O_2164,N_22342,N_24118);
nand UO_2165 (O_2165,N_23357,N_22795);
or UO_2166 (O_2166,N_23534,N_23749);
xnor UO_2167 (O_2167,N_23229,N_22453);
and UO_2168 (O_2168,N_24480,N_23205);
and UO_2169 (O_2169,N_24747,N_24697);
nand UO_2170 (O_2170,N_23988,N_24349);
or UO_2171 (O_2171,N_24478,N_23354);
nand UO_2172 (O_2172,N_24489,N_23019);
nand UO_2173 (O_2173,N_24828,N_21966);
xnor UO_2174 (O_2174,N_24666,N_24835);
and UO_2175 (O_2175,N_24779,N_21941);
and UO_2176 (O_2176,N_22147,N_23000);
nor UO_2177 (O_2177,N_24447,N_23602);
nor UO_2178 (O_2178,N_24499,N_23488);
and UO_2179 (O_2179,N_24030,N_24813);
and UO_2180 (O_2180,N_23499,N_23155);
xnor UO_2181 (O_2181,N_22487,N_22024);
or UO_2182 (O_2182,N_23764,N_23633);
nor UO_2183 (O_2183,N_21884,N_23406);
nor UO_2184 (O_2184,N_22692,N_24687);
nor UO_2185 (O_2185,N_23231,N_23201);
nand UO_2186 (O_2186,N_24717,N_22647);
or UO_2187 (O_2187,N_22073,N_24907);
and UO_2188 (O_2188,N_23185,N_23839);
nand UO_2189 (O_2189,N_23503,N_23948);
nor UO_2190 (O_2190,N_23891,N_22503);
xor UO_2191 (O_2191,N_24757,N_24379);
and UO_2192 (O_2192,N_22076,N_22973);
or UO_2193 (O_2193,N_24964,N_23957);
and UO_2194 (O_2194,N_24563,N_24153);
xnor UO_2195 (O_2195,N_24594,N_23431);
or UO_2196 (O_2196,N_24586,N_24091);
nor UO_2197 (O_2197,N_24915,N_22441);
nor UO_2198 (O_2198,N_23899,N_22312);
and UO_2199 (O_2199,N_24743,N_24507);
and UO_2200 (O_2200,N_24114,N_22940);
nor UO_2201 (O_2201,N_24962,N_23744);
and UO_2202 (O_2202,N_23814,N_24163);
or UO_2203 (O_2203,N_24711,N_24997);
nand UO_2204 (O_2204,N_23279,N_23284);
or UO_2205 (O_2205,N_23788,N_22314);
and UO_2206 (O_2206,N_22418,N_23728);
and UO_2207 (O_2207,N_22743,N_22999);
xor UO_2208 (O_2208,N_22324,N_23939);
or UO_2209 (O_2209,N_22291,N_22850);
and UO_2210 (O_2210,N_21935,N_24805);
and UO_2211 (O_2211,N_22273,N_24625);
xor UO_2212 (O_2212,N_24686,N_22361);
nor UO_2213 (O_2213,N_22763,N_23462);
and UO_2214 (O_2214,N_22025,N_24327);
and UO_2215 (O_2215,N_24595,N_23737);
nand UO_2216 (O_2216,N_23276,N_23327);
nand UO_2217 (O_2217,N_24874,N_23947);
and UO_2218 (O_2218,N_24961,N_24301);
or UO_2219 (O_2219,N_24962,N_24800);
xnor UO_2220 (O_2220,N_23505,N_24334);
and UO_2221 (O_2221,N_23358,N_23719);
and UO_2222 (O_2222,N_24086,N_24605);
or UO_2223 (O_2223,N_24105,N_24325);
nor UO_2224 (O_2224,N_22420,N_23081);
or UO_2225 (O_2225,N_22665,N_24019);
xor UO_2226 (O_2226,N_21995,N_24228);
nor UO_2227 (O_2227,N_22245,N_24936);
or UO_2228 (O_2228,N_22215,N_24801);
and UO_2229 (O_2229,N_24606,N_22952);
xor UO_2230 (O_2230,N_22401,N_23968);
or UO_2231 (O_2231,N_22412,N_22937);
nor UO_2232 (O_2232,N_23108,N_23982);
and UO_2233 (O_2233,N_24211,N_24954);
xor UO_2234 (O_2234,N_22536,N_24121);
nor UO_2235 (O_2235,N_24020,N_23027);
nand UO_2236 (O_2236,N_24730,N_24690);
and UO_2237 (O_2237,N_22824,N_23743);
nand UO_2238 (O_2238,N_24734,N_24542);
nor UO_2239 (O_2239,N_22838,N_24820);
or UO_2240 (O_2240,N_22391,N_24594);
nor UO_2241 (O_2241,N_24887,N_22040);
nand UO_2242 (O_2242,N_22921,N_22375);
nand UO_2243 (O_2243,N_21963,N_22458);
and UO_2244 (O_2244,N_22024,N_22777);
nor UO_2245 (O_2245,N_22018,N_22871);
and UO_2246 (O_2246,N_23326,N_24063);
nor UO_2247 (O_2247,N_22580,N_24290);
and UO_2248 (O_2248,N_24757,N_23982);
and UO_2249 (O_2249,N_24692,N_22814);
xor UO_2250 (O_2250,N_24176,N_22207);
or UO_2251 (O_2251,N_24562,N_23828);
nand UO_2252 (O_2252,N_23516,N_24469);
nand UO_2253 (O_2253,N_22845,N_23556);
xor UO_2254 (O_2254,N_22067,N_23101);
nor UO_2255 (O_2255,N_23372,N_24897);
nor UO_2256 (O_2256,N_22993,N_24966);
or UO_2257 (O_2257,N_23449,N_22258);
and UO_2258 (O_2258,N_24001,N_23087);
nor UO_2259 (O_2259,N_24930,N_23142);
and UO_2260 (O_2260,N_24042,N_24119);
and UO_2261 (O_2261,N_23217,N_22724);
nand UO_2262 (O_2262,N_24634,N_22096);
nor UO_2263 (O_2263,N_24905,N_23912);
nand UO_2264 (O_2264,N_22095,N_22064);
nand UO_2265 (O_2265,N_22595,N_23267);
or UO_2266 (O_2266,N_22154,N_22570);
nand UO_2267 (O_2267,N_23891,N_22282);
nor UO_2268 (O_2268,N_22199,N_24538);
and UO_2269 (O_2269,N_23606,N_23708);
nor UO_2270 (O_2270,N_24181,N_24753);
or UO_2271 (O_2271,N_23804,N_23344);
or UO_2272 (O_2272,N_22415,N_24142);
nand UO_2273 (O_2273,N_23444,N_24000);
xor UO_2274 (O_2274,N_24814,N_23423);
nor UO_2275 (O_2275,N_22797,N_24136);
or UO_2276 (O_2276,N_24044,N_24166);
nand UO_2277 (O_2277,N_23512,N_24854);
and UO_2278 (O_2278,N_24372,N_24296);
nand UO_2279 (O_2279,N_23016,N_23915);
xor UO_2280 (O_2280,N_24203,N_22050);
and UO_2281 (O_2281,N_22978,N_21965);
nand UO_2282 (O_2282,N_23312,N_23166);
nand UO_2283 (O_2283,N_23655,N_22586);
nand UO_2284 (O_2284,N_24211,N_22111);
nor UO_2285 (O_2285,N_24213,N_22127);
or UO_2286 (O_2286,N_24470,N_22107);
or UO_2287 (O_2287,N_24441,N_24734);
nor UO_2288 (O_2288,N_24468,N_23607);
nand UO_2289 (O_2289,N_22283,N_24336);
or UO_2290 (O_2290,N_24245,N_24039);
or UO_2291 (O_2291,N_23258,N_22667);
xnor UO_2292 (O_2292,N_23685,N_22048);
and UO_2293 (O_2293,N_23607,N_24733);
nand UO_2294 (O_2294,N_23962,N_22931);
or UO_2295 (O_2295,N_23363,N_23522);
nor UO_2296 (O_2296,N_23468,N_24950);
and UO_2297 (O_2297,N_22526,N_23464);
nor UO_2298 (O_2298,N_23657,N_24777);
or UO_2299 (O_2299,N_24677,N_22565);
nand UO_2300 (O_2300,N_24059,N_23132);
and UO_2301 (O_2301,N_21968,N_22317);
and UO_2302 (O_2302,N_22197,N_21957);
nand UO_2303 (O_2303,N_22644,N_23844);
or UO_2304 (O_2304,N_21983,N_23143);
and UO_2305 (O_2305,N_23345,N_24980);
and UO_2306 (O_2306,N_22851,N_23467);
nand UO_2307 (O_2307,N_22992,N_22201);
or UO_2308 (O_2308,N_22775,N_24991);
nand UO_2309 (O_2309,N_23925,N_21948);
nor UO_2310 (O_2310,N_24193,N_23633);
and UO_2311 (O_2311,N_24089,N_24111);
nor UO_2312 (O_2312,N_23930,N_22664);
or UO_2313 (O_2313,N_22650,N_22789);
nor UO_2314 (O_2314,N_22837,N_23569);
and UO_2315 (O_2315,N_23783,N_24397);
xor UO_2316 (O_2316,N_23360,N_23486);
or UO_2317 (O_2317,N_22583,N_24531);
nand UO_2318 (O_2318,N_24175,N_24063);
nor UO_2319 (O_2319,N_24172,N_22589);
or UO_2320 (O_2320,N_22282,N_23404);
and UO_2321 (O_2321,N_21919,N_23943);
nand UO_2322 (O_2322,N_23413,N_23631);
and UO_2323 (O_2323,N_24539,N_24685);
and UO_2324 (O_2324,N_22590,N_24065);
nand UO_2325 (O_2325,N_24917,N_23648);
nor UO_2326 (O_2326,N_23456,N_22443);
nor UO_2327 (O_2327,N_24823,N_24380);
or UO_2328 (O_2328,N_23235,N_22388);
or UO_2329 (O_2329,N_23848,N_24099);
nor UO_2330 (O_2330,N_22759,N_22524);
nor UO_2331 (O_2331,N_23415,N_24882);
or UO_2332 (O_2332,N_22614,N_22789);
and UO_2333 (O_2333,N_23323,N_24141);
and UO_2334 (O_2334,N_23739,N_24832);
xor UO_2335 (O_2335,N_24369,N_24704);
nor UO_2336 (O_2336,N_22483,N_22738);
nor UO_2337 (O_2337,N_22911,N_24078);
and UO_2338 (O_2338,N_22675,N_24339);
or UO_2339 (O_2339,N_22689,N_22719);
nor UO_2340 (O_2340,N_23661,N_24520);
and UO_2341 (O_2341,N_22721,N_23469);
nand UO_2342 (O_2342,N_24445,N_24800);
nand UO_2343 (O_2343,N_22108,N_22741);
or UO_2344 (O_2344,N_23841,N_24100);
xor UO_2345 (O_2345,N_23292,N_24370);
nand UO_2346 (O_2346,N_23693,N_24585);
or UO_2347 (O_2347,N_22559,N_24207);
xnor UO_2348 (O_2348,N_24225,N_23252);
nor UO_2349 (O_2349,N_24186,N_24577);
nand UO_2350 (O_2350,N_24141,N_23141);
or UO_2351 (O_2351,N_22153,N_23682);
or UO_2352 (O_2352,N_24932,N_24635);
nor UO_2353 (O_2353,N_24077,N_22424);
nor UO_2354 (O_2354,N_22350,N_22890);
and UO_2355 (O_2355,N_23932,N_21909);
nand UO_2356 (O_2356,N_22799,N_21946);
and UO_2357 (O_2357,N_23145,N_23857);
and UO_2358 (O_2358,N_22146,N_21906);
nand UO_2359 (O_2359,N_23593,N_23354);
xor UO_2360 (O_2360,N_22949,N_23651);
or UO_2361 (O_2361,N_23531,N_23732);
or UO_2362 (O_2362,N_22014,N_22063);
and UO_2363 (O_2363,N_22100,N_24398);
and UO_2364 (O_2364,N_22242,N_22129);
and UO_2365 (O_2365,N_24855,N_21897);
nor UO_2366 (O_2366,N_23839,N_22266);
nor UO_2367 (O_2367,N_23169,N_23636);
xor UO_2368 (O_2368,N_24950,N_22187);
nand UO_2369 (O_2369,N_23566,N_24427);
or UO_2370 (O_2370,N_23346,N_22671);
nor UO_2371 (O_2371,N_22176,N_24375);
nor UO_2372 (O_2372,N_24827,N_22287);
nor UO_2373 (O_2373,N_22831,N_24566);
and UO_2374 (O_2374,N_23487,N_22583);
nand UO_2375 (O_2375,N_23835,N_22152);
and UO_2376 (O_2376,N_22716,N_24912);
nand UO_2377 (O_2377,N_23239,N_24398);
nor UO_2378 (O_2378,N_23343,N_22744);
and UO_2379 (O_2379,N_23551,N_23496);
nand UO_2380 (O_2380,N_23880,N_22407);
and UO_2381 (O_2381,N_24338,N_24601);
and UO_2382 (O_2382,N_24628,N_22222);
or UO_2383 (O_2383,N_23831,N_21984);
nor UO_2384 (O_2384,N_24061,N_22779);
nor UO_2385 (O_2385,N_23762,N_23922);
and UO_2386 (O_2386,N_23111,N_23155);
or UO_2387 (O_2387,N_24624,N_21975);
nand UO_2388 (O_2388,N_24446,N_24351);
nand UO_2389 (O_2389,N_22168,N_22678);
nand UO_2390 (O_2390,N_22276,N_22315);
nor UO_2391 (O_2391,N_22141,N_23163);
nand UO_2392 (O_2392,N_23359,N_22719);
or UO_2393 (O_2393,N_23547,N_23090);
and UO_2394 (O_2394,N_24785,N_23080);
and UO_2395 (O_2395,N_23449,N_23544);
nor UO_2396 (O_2396,N_24295,N_24394);
and UO_2397 (O_2397,N_23943,N_22132);
nor UO_2398 (O_2398,N_24516,N_22767);
xnor UO_2399 (O_2399,N_21968,N_22970);
or UO_2400 (O_2400,N_22321,N_23817);
or UO_2401 (O_2401,N_22973,N_23265);
and UO_2402 (O_2402,N_22086,N_23868);
and UO_2403 (O_2403,N_24438,N_23087);
and UO_2404 (O_2404,N_23428,N_24179);
xor UO_2405 (O_2405,N_22942,N_24668);
and UO_2406 (O_2406,N_23328,N_23497);
nand UO_2407 (O_2407,N_23526,N_23884);
and UO_2408 (O_2408,N_24271,N_23143);
and UO_2409 (O_2409,N_22696,N_23368);
nand UO_2410 (O_2410,N_23843,N_23202);
and UO_2411 (O_2411,N_24426,N_24732);
xnor UO_2412 (O_2412,N_23068,N_22548);
or UO_2413 (O_2413,N_24129,N_23907);
nand UO_2414 (O_2414,N_22426,N_23570);
xor UO_2415 (O_2415,N_23328,N_22015);
and UO_2416 (O_2416,N_22871,N_22714);
or UO_2417 (O_2417,N_22095,N_22486);
and UO_2418 (O_2418,N_22669,N_23319);
nor UO_2419 (O_2419,N_23287,N_23256);
and UO_2420 (O_2420,N_24351,N_21907);
nand UO_2421 (O_2421,N_22397,N_24398);
or UO_2422 (O_2422,N_23171,N_24999);
nand UO_2423 (O_2423,N_21929,N_24608);
xor UO_2424 (O_2424,N_23632,N_23591);
and UO_2425 (O_2425,N_22091,N_24857);
and UO_2426 (O_2426,N_23770,N_24075);
and UO_2427 (O_2427,N_23236,N_23674);
nand UO_2428 (O_2428,N_23362,N_24028);
nand UO_2429 (O_2429,N_24851,N_23205);
nand UO_2430 (O_2430,N_21940,N_23973);
xnor UO_2431 (O_2431,N_22551,N_24318);
or UO_2432 (O_2432,N_23742,N_24376);
nand UO_2433 (O_2433,N_21972,N_23792);
and UO_2434 (O_2434,N_23578,N_22162);
or UO_2435 (O_2435,N_23310,N_23588);
nand UO_2436 (O_2436,N_23171,N_24988);
nand UO_2437 (O_2437,N_24908,N_23649);
or UO_2438 (O_2438,N_23414,N_22719);
nor UO_2439 (O_2439,N_24310,N_22161);
nor UO_2440 (O_2440,N_23156,N_24749);
xor UO_2441 (O_2441,N_23259,N_23073);
and UO_2442 (O_2442,N_24421,N_24400);
xor UO_2443 (O_2443,N_24034,N_24864);
xor UO_2444 (O_2444,N_22225,N_24588);
and UO_2445 (O_2445,N_24150,N_22020);
or UO_2446 (O_2446,N_24222,N_24980);
and UO_2447 (O_2447,N_23276,N_22981);
or UO_2448 (O_2448,N_23772,N_23553);
and UO_2449 (O_2449,N_23869,N_22941);
nand UO_2450 (O_2450,N_23613,N_23699);
xnor UO_2451 (O_2451,N_24270,N_22752);
nor UO_2452 (O_2452,N_23560,N_22325);
nor UO_2453 (O_2453,N_24273,N_22009);
and UO_2454 (O_2454,N_22559,N_22934);
xor UO_2455 (O_2455,N_24154,N_23580);
nor UO_2456 (O_2456,N_23004,N_22900);
xor UO_2457 (O_2457,N_22921,N_22440);
nor UO_2458 (O_2458,N_24641,N_23199);
nand UO_2459 (O_2459,N_24196,N_24884);
or UO_2460 (O_2460,N_22754,N_24296);
or UO_2461 (O_2461,N_21905,N_23298);
xnor UO_2462 (O_2462,N_24245,N_22154);
nand UO_2463 (O_2463,N_23089,N_22582);
nand UO_2464 (O_2464,N_22995,N_24733);
and UO_2465 (O_2465,N_24254,N_24734);
nor UO_2466 (O_2466,N_22698,N_24856);
xnor UO_2467 (O_2467,N_24113,N_22100);
and UO_2468 (O_2468,N_21895,N_23533);
nand UO_2469 (O_2469,N_24207,N_21926);
or UO_2470 (O_2470,N_22302,N_24132);
or UO_2471 (O_2471,N_22584,N_24872);
nor UO_2472 (O_2472,N_22167,N_23302);
nand UO_2473 (O_2473,N_22061,N_21939);
and UO_2474 (O_2474,N_24208,N_24018);
nand UO_2475 (O_2475,N_22087,N_22396);
nand UO_2476 (O_2476,N_21907,N_22695);
or UO_2477 (O_2477,N_22123,N_24595);
or UO_2478 (O_2478,N_23954,N_23071);
or UO_2479 (O_2479,N_24394,N_22958);
nand UO_2480 (O_2480,N_23293,N_24232);
xor UO_2481 (O_2481,N_24592,N_22317);
nor UO_2482 (O_2482,N_23721,N_22852);
nand UO_2483 (O_2483,N_22105,N_24547);
and UO_2484 (O_2484,N_24998,N_22699);
or UO_2485 (O_2485,N_23658,N_24813);
or UO_2486 (O_2486,N_24606,N_22561);
nand UO_2487 (O_2487,N_23675,N_24663);
or UO_2488 (O_2488,N_22487,N_24365);
nand UO_2489 (O_2489,N_24481,N_22208);
nor UO_2490 (O_2490,N_24948,N_23923);
or UO_2491 (O_2491,N_22866,N_24338);
or UO_2492 (O_2492,N_24409,N_24322);
and UO_2493 (O_2493,N_23022,N_24559);
or UO_2494 (O_2494,N_24595,N_24123);
and UO_2495 (O_2495,N_24308,N_22823);
nand UO_2496 (O_2496,N_23906,N_23031);
or UO_2497 (O_2497,N_22328,N_23522);
nor UO_2498 (O_2498,N_23095,N_24651);
nor UO_2499 (O_2499,N_23822,N_24590);
or UO_2500 (O_2500,N_22795,N_24473);
or UO_2501 (O_2501,N_22149,N_23840);
xnor UO_2502 (O_2502,N_24239,N_24167);
nor UO_2503 (O_2503,N_24793,N_24457);
or UO_2504 (O_2504,N_22762,N_22881);
and UO_2505 (O_2505,N_23408,N_23736);
nor UO_2506 (O_2506,N_22556,N_22671);
nor UO_2507 (O_2507,N_23014,N_23354);
nor UO_2508 (O_2508,N_23501,N_22242);
nor UO_2509 (O_2509,N_24575,N_24183);
or UO_2510 (O_2510,N_22571,N_23293);
nor UO_2511 (O_2511,N_22657,N_24037);
or UO_2512 (O_2512,N_22914,N_24201);
nor UO_2513 (O_2513,N_24769,N_21979);
nand UO_2514 (O_2514,N_22264,N_24535);
and UO_2515 (O_2515,N_22023,N_24091);
or UO_2516 (O_2516,N_24824,N_23330);
nand UO_2517 (O_2517,N_24673,N_23461);
and UO_2518 (O_2518,N_23374,N_22377);
nand UO_2519 (O_2519,N_21930,N_22266);
or UO_2520 (O_2520,N_22352,N_24893);
or UO_2521 (O_2521,N_22155,N_24342);
nand UO_2522 (O_2522,N_22067,N_23610);
nor UO_2523 (O_2523,N_22337,N_22858);
or UO_2524 (O_2524,N_24207,N_23103);
nand UO_2525 (O_2525,N_23080,N_21914);
nand UO_2526 (O_2526,N_23213,N_24611);
or UO_2527 (O_2527,N_23895,N_24901);
xor UO_2528 (O_2528,N_24104,N_24815);
or UO_2529 (O_2529,N_22546,N_23059);
or UO_2530 (O_2530,N_22395,N_23907);
nor UO_2531 (O_2531,N_23846,N_23038);
nor UO_2532 (O_2532,N_23678,N_23560);
and UO_2533 (O_2533,N_22646,N_22976);
and UO_2534 (O_2534,N_24905,N_24792);
nand UO_2535 (O_2535,N_22180,N_22423);
and UO_2536 (O_2536,N_23938,N_24766);
or UO_2537 (O_2537,N_22536,N_24213);
nor UO_2538 (O_2538,N_23697,N_22476);
nor UO_2539 (O_2539,N_22925,N_22334);
or UO_2540 (O_2540,N_24662,N_24995);
or UO_2541 (O_2541,N_24924,N_23731);
nand UO_2542 (O_2542,N_24558,N_24893);
nand UO_2543 (O_2543,N_24478,N_24672);
or UO_2544 (O_2544,N_23996,N_23271);
nor UO_2545 (O_2545,N_22484,N_23257);
nor UO_2546 (O_2546,N_22232,N_24827);
or UO_2547 (O_2547,N_24812,N_22712);
nand UO_2548 (O_2548,N_23821,N_22514);
nand UO_2549 (O_2549,N_22422,N_24479);
xnor UO_2550 (O_2550,N_24435,N_22404);
or UO_2551 (O_2551,N_24816,N_22284);
or UO_2552 (O_2552,N_23245,N_22948);
nor UO_2553 (O_2553,N_22233,N_24514);
nand UO_2554 (O_2554,N_22038,N_23281);
nand UO_2555 (O_2555,N_23110,N_24763);
nand UO_2556 (O_2556,N_24095,N_24419);
and UO_2557 (O_2557,N_24199,N_22217);
and UO_2558 (O_2558,N_24047,N_23853);
nand UO_2559 (O_2559,N_24429,N_22028);
and UO_2560 (O_2560,N_23270,N_24248);
nand UO_2561 (O_2561,N_22800,N_24316);
or UO_2562 (O_2562,N_22398,N_23847);
nor UO_2563 (O_2563,N_23866,N_22323);
and UO_2564 (O_2564,N_24754,N_23525);
or UO_2565 (O_2565,N_24165,N_22998);
or UO_2566 (O_2566,N_22480,N_22855);
nor UO_2567 (O_2567,N_22173,N_23812);
nor UO_2568 (O_2568,N_22704,N_22014);
or UO_2569 (O_2569,N_23280,N_23700);
or UO_2570 (O_2570,N_22947,N_22966);
and UO_2571 (O_2571,N_22580,N_23685);
nor UO_2572 (O_2572,N_22987,N_24928);
xnor UO_2573 (O_2573,N_22166,N_22122);
nor UO_2574 (O_2574,N_22184,N_22862);
or UO_2575 (O_2575,N_22305,N_23847);
and UO_2576 (O_2576,N_24604,N_23135);
and UO_2577 (O_2577,N_23148,N_24677);
nand UO_2578 (O_2578,N_22143,N_23678);
and UO_2579 (O_2579,N_23157,N_22072);
nor UO_2580 (O_2580,N_21999,N_24785);
nor UO_2581 (O_2581,N_23441,N_22507);
nand UO_2582 (O_2582,N_22064,N_24780);
and UO_2583 (O_2583,N_22501,N_23089);
nor UO_2584 (O_2584,N_23588,N_24044);
xor UO_2585 (O_2585,N_22040,N_23287);
nand UO_2586 (O_2586,N_22573,N_23751);
or UO_2587 (O_2587,N_22121,N_22649);
and UO_2588 (O_2588,N_23905,N_24820);
nand UO_2589 (O_2589,N_24385,N_23171);
and UO_2590 (O_2590,N_23711,N_24980);
xor UO_2591 (O_2591,N_24641,N_24211);
or UO_2592 (O_2592,N_23259,N_22556);
xor UO_2593 (O_2593,N_23683,N_24296);
xnor UO_2594 (O_2594,N_22018,N_22724);
and UO_2595 (O_2595,N_22156,N_23275);
nand UO_2596 (O_2596,N_22212,N_24819);
or UO_2597 (O_2597,N_24820,N_22603);
and UO_2598 (O_2598,N_24684,N_21882);
nor UO_2599 (O_2599,N_22459,N_22977);
and UO_2600 (O_2600,N_24562,N_22523);
or UO_2601 (O_2601,N_24475,N_24587);
or UO_2602 (O_2602,N_22286,N_23049);
nand UO_2603 (O_2603,N_22741,N_24573);
or UO_2604 (O_2604,N_23921,N_23746);
nand UO_2605 (O_2605,N_24653,N_24135);
nand UO_2606 (O_2606,N_21876,N_23172);
and UO_2607 (O_2607,N_22256,N_24806);
nand UO_2608 (O_2608,N_24708,N_24007);
or UO_2609 (O_2609,N_21905,N_24127);
nand UO_2610 (O_2610,N_24749,N_24316);
and UO_2611 (O_2611,N_24159,N_24659);
or UO_2612 (O_2612,N_22828,N_23672);
nand UO_2613 (O_2613,N_24078,N_24540);
and UO_2614 (O_2614,N_23069,N_22131);
and UO_2615 (O_2615,N_24449,N_21906);
nand UO_2616 (O_2616,N_24253,N_22913);
nand UO_2617 (O_2617,N_24447,N_24366);
or UO_2618 (O_2618,N_24428,N_23982);
nor UO_2619 (O_2619,N_22652,N_22062);
nor UO_2620 (O_2620,N_23207,N_24282);
or UO_2621 (O_2621,N_23993,N_23510);
nor UO_2622 (O_2622,N_22759,N_24760);
or UO_2623 (O_2623,N_21940,N_23137);
xnor UO_2624 (O_2624,N_22607,N_21963);
nor UO_2625 (O_2625,N_22196,N_23533);
nor UO_2626 (O_2626,N_23261,N_24627);
and UO_2627 (O_2627,N_23011,N_21959);
and UO_2628 (O_2628,N_24769,N_23240);
and UO_2629 (O_2629,N_24228,N_22404);
and UO_2630 (O_2630,N_22490,N_22940);
nor UO_2631 (O_2631,N_24518,N_23369);
nor UO_2632 (O_2632,N_24090,N_23078);
nand UO_2633 (O_2633,N_22251,N_24216);
xnor UO_2634 (O_2634,N_23195,N_24038);
or UO_2635 (O_2635,N_24167,N_23944);
or UO_2636 (O_2636,N_22864,N_23678);
and UO_2637 (O_2637,N_23280,N_23334);
nor UO_2638 (O_2638,N_24241,N_22419);
nand UO_2639 (O_2639,N_23147,N_23953);
nand UO_2640 (O_2640,N_22380,N_22229);
nand UO_2641 (O_2641,N_23451,N_23396);
xnor UO_2642 (O_2642,N_22909,N_22027);
or UO_2643 (O_2643,N_24790,N_24158);
xnor UO_2644 (O_2644,N_22176,N_23062);
and UO_2645 (O_2645,N_24232,N_22393);
xnor UO_2646 (O_2646,N_22986,N_24099);
nand UO_2647 (O_2647,N_23406,N_22520);
nand UO_2648 (O_2648,N_22201,N_23393);
nor UO_2649 (O_2649,N_23521,N_23162);
nor UO_2650 (O_2650,N_23043,N_23466);
nand UO_2651 (O_2651,N_24753,N_24955);
nand UO_2652 (O_2652,N_22718,N_23013);
or UO_2653 (O_2653,N_22853,N_23616);
nor UO_2654 (O_2654,N_24352,N_23855);
or UO_2655 (O_2655,N_24780,N_22169);
nand UO_2656 (O_2656,N_23200,N_24776);
nand UO_2657 (O_2657,N_22946,N_24444);
xnor UO_2658 (O_2658,N_22882,N_22890);
xnor UO_2659 (O_2659,N_24184,N_22782);
or UO_2660 (O_2660,N_22712,N_24973);
nor UO_2661 (O_2661,N_22207,N_22462);
and UO_2662 (O_2662,N_24511,N_22519);
nand UO_2663 (O_2663,N_22151,N_24336);
nand UO_2664 (O_2664,N_24706,N_22486);
nor UO_2665 (O_2665,N_24316,N_24600);
and UO_2666 (O_2666,N_22027,N_24682);
nand UO_2667 (O_2667,N_23730,N_24291);
and UO_2668 (O_2668,N_24104,N_23003);
nand UO_2669 (O_2669,N_23076,N_22698);
or UO_2670 (O_2670,N_24569,N_23368);
and UO_2671 (O_2671,N_24049,N_23938);
or UO_2672 (O_2672,N_22322,N_22095);
nor UO_2673 (O_2673,N_23597,N_22127);
or UO_2674 (O_2674,N_22335,N_21885);
and UO_2675 (O_2675,N_21958,N_23111);
nor UO_2676 (O_2676,N_24362,N_23531);
nand UO_2677 (O_2677,N_24152,N_24310);
nand UO_2678 (O_2678,N_23582,N_23144);
nand UO_2679 (O_2679,N_24451,N_22215);
and UO_2680 (O_2680,N_24525,N_23995);
xnor UO_2681 (O_2681,N_24370,N_23019);
or UO_2682 (O_2682,N_24110,N_21911);
or UO_2683 (O_2683,N_22858,N_23370);
nor UO_2684 (O_2684,N_23737,N_24229);
nand UO_2685 (O_2685,N_22207,N_24260);
or UO_2686 (O_2686,N_23896,N_22107);
nand UO_2687 (O_2687,N_23279,N_22589);
nand UO_2688 (O_2688,N_22381,N_24430);
nand UO_2689 (O_2689,N_24927,N_23680);
and UO_2690 (O_2690,N_22568,N_24257);
nand UO_2691 (O_2691,N_23061,N_21919);
and UO_2692 (O_2692,N_24667,N_22041);
nand UO_2693 (O_2693,N_24486,N_24740);
nand UO_2694 (O_2694,N_23973,N_23955);
xnor UO_2695 (O_2695,N_23950,N_23367);
nor UO_2696 (O_2696,N_22973,N_24660);
or UO_2697 (O_2697,N_23769,N_23083);
nor UO_2698 (O_2698,N_24568,N_22938);
or UO_2699 (O_2699,N_22890,N_23975);
nor UO_2700 (O_2700,N_24779,N_23528);
or UO_2701 (O_2701,N_23490,N_24309);
and UO_2702 (O_2702,N_22409,N_23809);
nand UO_2703 (O_2703,N_23076,N_23074);
or UO_2704 (O_2704,N_24825,N_23623);
nand UO_2705 (O_2705,N_22033,N_22288);
nand UO_2706 (O_2706,N_24777,N_24215);
nor UO_2707 (O_2707,N_24642,N_23798);
and UO_2708 (O_2708,N_23246,N_24203);
and UO_2709 (O_2709,N_22812,N_23812);
and UO_2710 (O_2710,N_22830,N_24499);
or UO_2711 (O_2711,N_23458,N_22778);
nand UO_2712 (O_2712,N_24652,N_22262);
or UO_2713 (O_2713,N_22765,N_22457);
or UO_2714 (O_2714,N_24692,N_22453);
and UO_2715 (O_2715,N_23184,N_22087);
and UO_2716 (O_2716,N_22901,N_22527);
or UO_2717 (O_2717,N_24965,N_24272);
nor UO_2718 (O_2718,N_24865,N_22689);
and UO_2719 (O_2719,N_22133,N_24267);
or UO_2720 (O_2720,N_22770,N_24269);
xor UO_2721 (O_2721,N_24172,N_23983);
nor UO_2722 (O_2722,N_24211,N_24091);
or UO_2723 (O_2723,N_22048,N_23971);
nand UO_2724 (O_2724,N_22968,N_23516);
nand UO_2725 (O_2725,N_23001,N_22537);
nor UO_2726 (O_2726,N_24935,N_23656);
and UO_2727 (O_2727,N_22823,N_22529);
xor UO_2728 (O_2728,N_22452,N_22526);
and UO_2729 (O_2729,N_23394,N_22330);
xnor UO_2730 (O_2730,N_22286,N_22023);
nand UO_2731 (O_2731,N_23835,N_24021);
xnor UO_2732 (O_2732,N_23955,N_23950);
nand UO_2733 (O_2733,N_24114,N_23370);
or UO_2734 (O_2734,N_22356,N_22063);
and UO_2735 (O_2735,N_23074,N_22767);
xor UO_2736 (O_2736,N_21894,N_24440);
xor UO_2737 (O_2737,N_22144,N_23404);
nor UO_2738 (O_2738,N_22647,N_23833);
or UO_2739 (O_2739,N_21981,N_24690);
xnor UO_2740 (O_2740,N_23838,N_24595);
and UO_2741 (O_2741,N_24468,N_24260);
xnor UO_2742 (O_2742,N_24603,N_22537);
nor UO_2743 (O_2743,N_22245,N_24772);
or UO_2744 (O_2744,N_22473,N_22792);
or UO_2745 (O_2745,N_24196,N_23102);
xor UO_2746 (O_2746,N_23970,N_23281);
and UO_2747 (O_2747,N_23125,N_23041);
nand UO_2748 (O_2748,N_24581,N_22927);
xnor UO_2749 (O_2749,N_23161,N_22653);
nand UO_2750 (O_2750,N_23460,N_22099);
or UO_2751 (O_2751,N_23631,N_22429);
and UO_2752 (O_2752,N_23879,N_22617);
or UO_2753 (O_2753,N_23038,N_24557);
xor UO_2754 (O_2754,N_23900,N_23864);
nand UO_2755 (O_2755,N_22425,N_22192);
xnor UO_2756 (O_2756,N_24846,N_22664);
nor UO_2757 (O_2757,N_22208,N_24841);
nand UO_2758 (O_2758,N_22886,N_24329);
nor UO_2759 (O_2759,N_22478,N_22071);
nor UO_2760 (O_2760,N_23877,N_24319);
and UO_2761 (O_2761,N_23926,N_24257);
and UO_2762 (O_2762,N_23041,N_22906);
nand UO_2763 (O_2763,N_22658,N_22581);
nor UO_2764 (O_2764,N_24293,N_23865);
nand UO_2765 (O_2765,N_22044,N_24405);
nand UO_2766 (O_2766,N_23897,N_22576);
nor UO_2767 (O_2767,N_24666,N_23392);
nor UO_2768 (O_2768,N_22640,N_24608);
nand UO_2769 (O_2769,N_24844,N_24496);
xnor UO_2770 (O_2770,N_24190,N_24480);
or UO_2771 (O_2771,N_22380,N_22545);
or UO_2772 (O_2772,N_22920,N_22332);
and UO_2773 (O_2773,N_24646,N_23934);
xnor UO_2774 (O_2774,N_24032,N_22675);
or UO_2775 (O_2775,N_22685,N_24453);
nand UO_2776 (O_2776,N_23024,N_22304);
or UO_2777 (O_2777,N_24485,N_24710);
nor UO_2778 (O_2778,N_21943,N_24285);
and UO_2779 (O_2779,N_22108,N_21963);
nor UO_2780 (O_2780,N_24382,N_22670);
and UO_2781 (O_2781,N_24724,N_24886);
xor UO_2782 (O_2782,N_23936,N_24537);
and UO_2783 (O_2783,N_24726,N_23800);
and UO_2784 (O_2784,N_24659,N_22558);
or UO_2785 (O_2785,N_23471,N_22464);
nand UO_2786 (O_2786,N_23053,N_23190);
and UO_2787 (O_2787,N_23543,N_22626);
nor UO_2788 (O_2788,N_24459,N_24645);
or UO_2789 (O_2789,N_24396,N_22412);
or UO_2790 (O_2790,N_22763,N_24895);
xor UO_2791 (O_2791,N_24952,N_22268);
or UO_2792 (O_2792,N_23874,N_23370);
nand UO_2793 (O_2793,N_24901,N_24576);
nor UO_2794 (O_2794,N_22969,N_22854);
and UO_2795 (O_2795,N_23909,N_22597);
and UO_2796 (O_2796,N_22967,N_23630);
nor UO_2797 (O_2797,N_24847,N_23464);
or UO_2798 (O_2798,N_23442,N_23986);
nand UO_2799 (O_2799,N_22911,N_24656);
and UO_2800 (O_2800,N_24470,N_23889);
nor UO_2801 (O_2801,N_24655,N_21986);
and UO_2802 (O_2802,N_22893,N_23922);
and UO_2803 (O_2803,N_22954,N_24631);
or UO_2804 (O_2804,N_24439,N_23786);
nor UO_2805 (O_2805,N_24726,N_22544);
xor UO_2806 (O_2806,N_23167,N_22959);
and UO_2807 (O_2807,N_23605,N_22661);
and UO_2808 (O_2808,N_24724,N_22639);
xor UO_2809 (O_2809,N_21934,N_23272);
or UO_2810 (O_2810,N_24678,N_23193);
nor UO_2811 (O_2811,N_24016,N_22769);
or UO_2812 (O_2812,N_24036,N_22400);
nor UO_2813 (O_2813,N_23883,N_22357);
nor UO_2814 (O_2814,N_23461,N_24093);
and UO_2815 (O_2815,N_24519,N_24538);
or UO_2816 (O_2816,N_23721,N_22669);
or UO_2817 (O_2817,N_23915,N_24115);
nand UO_2818 (O_2818,N_23042,N_22198);
or UO_2819 (O_2819,N_24713,N_22363);
and UO_2820 (O_2820,N_24130,N_23810);
and UO_2821 (O_2821,N_22788,N_22558);
nand UO_2822 (O_2822,N_22356,N_22499);
nor UO_2823 (O_2823,N_23101,N_24676);
or UO_2824 (O_2824,N_24259,N_23271);
nand UO_2825 (O_2825,N_22103,N_24356);
nor UO_2826 (O_2826,N_22226,N_24033);
nor UO_2827 (O_2827,N_22943,N_23374);
nor UO_2828 (O_2828,N_23733,N_23247);
nand UO_2829 (O_2829,N_23616,N_22361);
nand UO_2830 (O_2830,N_23022,N_22905);
nor UO_2831 (O_2831,N_24361,N_22276);
xor UO_2832 (O_2832,N_23350,N_24061);
nor UO_2833 (O_2833,N_23330,N_22526);
or UO_2834 (O_2834,N_22953,N_23497);
or UO_2835 (O_2835,N_23838,N_22842);
or UO_2836 (O_2836,N_23515,N_22418);
and UO_2837 (O_2837,N_22525,N_22677);
nor UO_2838 (O_2838,N_23484,N_22305);
nand UO_2839 (O_2839,N_22936,N_24852);
nand UO_2840 (O_2840,N_22830,N_23558);
nand UO_2841 (O_2841,N_23076,N_23345);
and UO_2842 (O_2842,N_24292,N_23294);
nand UO_2843 (O_2843,N_24829,N_24358);
nor UO_2844 (O_2844,N_23646,N_22252);
nand UO_2845 (O_2845,N_24056,N_24635);
or UO_2846 (O_2846,N_22820,N_22888);
and UO_2847 (O_2847,N_22965,N_23156);
and UO_2848 (O_2848,N_23995,N_22821);
and UO_2849 (O_2849,N_24115,N_22731);
nor UO_2850 (O_2850,N_24341,N_23139);
or UO_2851 (O_2851,N_23177,N_23993);
nor UO_2852 (O_2852,N_21967,N_23259);
and UO_2853 (O_2853,N_23771,N_24090);
and UO_2854 (O_2854,N_23025,N_24290);
and UO_2855 (O_2855,N_24181,N_24518);
xor UO_2856 (O_2856,N_22495,N_21959);
nor UO_2857 (O_2857,N_23182,N_22152);
xor UO_2858 (O_2858,N_24993,N_24374);
nor UO_2859 (O_2859,N_24443,N_24832);
nand UO_2860 (O_2860,N_24316,N_23294);
xnor UO_2861 (O_2861,N_24302,N_24602);
and UO_2862 (O_2862,N_24140,N_22266);
xnor UO_2863 (O_2863,N_24654,N_24327);
or UO_2864 (O_2864,N_23697,N_24530);
or UO_2865 (O_2865,N_24116,N_23100);
or UO_2866 (O_2866,N_23436,N_22557);
nor UO_2867 (O_2867,N_23431,N_23467);
nor UO_2868 (O_2868,N_22292,N_22571);
and UO_2869 (O_2869,N_24422,N_24483);
and UO_2870 (O_2870,N_23955,N_22454);
nor UO_2871 (O_2871,N_23214,N_24898);
nor UO_2872 (O_2872,N_24906,N_22451);
xnor UO_2873 (O_2873,N_22394,N_22849);
xor UO_2874 (O_2874,N_24747,N_22717);
nand UO_2875 (O_2875,N_24787,N_23536);
or UO_2876 (O_2876,N_23777,N_24905);
and UO_2877 (O_2877,N_23409,N_23188);
nand UO_2878 (O_2878,N_22860,N_23651);
and UO_2879 (O_2879,N_22577,N_22745);
xor UO_2880 (O_2880,N_24120,N_22851);
and UO_2881 (O_2881,N_23029,N_22776);
xor UO_2882 (O_2882,N_23826,N_22150);
and UO_2883 (O_2883,N_23288,N_24636);
nor UO_2884 (O_2884,N_24488,N_22432);
nor UO_2885 (O_2885,N_22058,N_24384);
and UO_2886 (O_2886,N_23244,N_24036);
or UO_2887 (O_2887,N_23986,N_24477);
and UO_2888 (O_2888,N_24380,N_24618);
or UO_2889 (O_2889,N_23462,N_24134);
nor UO_2890 (O_2890,N_24214,N_23549);
nand UO_2891 (O_2891,N_24661,N_23779);
nor UO_2892 (O_2892,N_23492,N_22707);
nor UO_2893 (O_2893,N_22426,N_22221);
or UO_2894 (O_2894,N_22288,N_23095);
or UO_2895 (O_2895,N_24193,N_23694);
nand UO_2896 (O_2896,N_22757,N_22193);
nor UO_2897 (O_2897,N_23069,N_22720);
nand UO_2898 (O_2898,N_23994,N_23211);
nor UO_2899 (O_2899,N_23219,N_22802);
nor UO_2900 (O_2900,N_23064,N_24005);
or UO_2901 (O_2901,N_24517,N_24395);
and UO_2902 (O_2902,N_22534,N_23900);
or UO_2903 (O_2903,N_22134,N_24935);
or UO_2904 (O_2904,N_24201,N_22578);
and UO_2905 (O_2905,N_24290,N_22540);
or UO_2906 (O_2906,N_24235,N_24878);
and UO_2907 (O_2907,N_22937,N_23752);
and UO_2908 (O_2908,N_22049,N_23079);
xnor UO_2909 (O_2909,N_22760,N_24742);
nor UO_2910 (O_2910,N_22539,N_24172);
nor UO_2911 (O_2911,N_24402,N_22291);
nand UO_2912 (O_2912,N_24572,N_22696);
or UO_2913 (O_2913,N_22198,N_23317);
xnor UO_2914 (O_2914,N_21908,N_24801);
nand UO_2915 (O_2915,N_22685,N_24015);
nand UO_2916 (O_2916,N_23035,N_23982);
or UO_2917 (O_2917,N_22419,N_23404);
nand UO_2918 (O_2918,N_22979,N_23817);
nand UO_2919 (O_2919,N_22388,N_24208);
nand UO_2920 (O_2920,N_24743,N_23969);
nor UO_2921 (O_2921,N_24373,N_23533);
or UO_2922 (O_2922,N_23792,N_24917);
nand UO_2923 (O_2923,N_22580,N_24333);
or UO_2924 (O_2924,N_22448,N_23510);
nor UO_2925 (O_2925,N_21994,N_24765);
or UO_2926 (O_2926,N_24574,N_22172);
nor UO_2927 (O_2927,N_23170,N_22418);
or UO_2928 (O_2928,N_22249,N_22058);
or UO_2929 (O_2929,N_24700,N_24382);
xnor UO_2930 (O_2930,N_22731,N_22359);
or UO_2931 (O_2931,N_23939,N_23178);
nand UO_2932 (O_2932,N_24389,N_24600);
or UO_2933 (O_2933,N_23148,N_21950);
nand UO_2934 (O_2934,N_23547,N_23422);
nor UO_2935 (O_2935,N_24949,N_23883);
nor UO_2936 (O_2936,N_22025,N_22335);
or UO_2937 (O_2937,N_23394,N_23986);
nor UO_2938 (O_2938,N_23501,N_24098);
or UO_2939 (O_2939,N_22192,N_23257);
nor UO_2940 (O_2940,N_24653,N_24040);
or UO_2941 (O_2941,N_22713,N_24107);
and UO_2942 (O_2942,N_24169,N_22850);
nand UO_2943 (O_2943,N_22495,N_22976);
nor UO_2944 (O_2944,N_24629,N_22478);
nor UO_2945 (O_2945,N_22345,N_22679);
nand UO_2946 (O_2946,N_22947,N_22118);
nand UO_2947 (O_2947,N_22179,N_23595);
or UO_2948 (O_2948,N_22417,N_24129);
or UO_2949 (O_2949,N_22780,N_22655);
or UO_2950 (O_2950,N_23056,N_23260);
nor UO_2951 (O_2951,N_24266,N_22389);
and UO_2952 (O_2952,N_23429,N_23364);
xnor UO_2953 (O_2953,N_23671,N_22020);
or UO_2954 (O_2954,N_23862,N_24857);
nor UO_2955 (O_2955,N_24139,N_24598);
xor UO_2956 (O_2956,N_23538,N_23048);
or UO_2957 (O_2957,N_23664,N_23525);
or UO_2958 (O_2958,N_23600,N_24664);
and UO_2959 (O_2959,N_23237,N_23035);
nor UO_2960 (O_2960,N_23006,N_22923);
nand UO_2961 (O_2961,N_22548,N_21969);
xor UO_2962 (O_2962,N_23389,N_24751);
xor UO_2963 (O_2963,N_24676,N_22581);
or UO_2964 (O_2964,N_22793,N_24519);
nor UO_2965 (O_2965,N_24259,N_23855);
and UO_2966 (O_2966,N_22302,N_23394);
nor UO_2967 (O_2967,N_22617,N_22268);
and UO_2968 (O_2968,N_24483,N_23981);
nor UO_2969 (O_2969,N_24897,N_21895);
and UO_2970 (O_2970,N_24170,N_23035);
and UO_2971 (O_2971,N_21959,N_22600);
nand UO_2972 (O_2972,N_22127,N_23606);
and UO_2973 (O_2973,N_24462,N_22544);
xnor UO_2974 (O_2974,N_22730,N_24094);
nor UO_2975 (O_2975,N_23024,N_22488);
nand UO_2976 (O_2976,N_23613,N_22782);
and UO_2977 (O_2977,N_23870,N_24604);
and UO_2978 (O_2978,N_24879,N_23137);
nand UO_2979 (O_2979,N_24832,N_24867);
nor UO_2980 (O_2980,N_23388,N_23669);
nor UO_2981 (O_2981,N_22822,N_22703);
and UO_2982 (O_2982,N_24443,N_22065);
nor UO_2983 (O_2983,N_23230,N_24439);
or UO_2984 (O_2984,N_22727,N_24046);
or UO_2985 (O_2985,N_22530,N_24416);
xor UO_2986 (O_2986,N_23938,N_23212);
nand UO_2987 (O_2987,N_23660,N_23164);
and UO_2988 (O_2988,N_22253,N_24399);
and UO_2989 (O_2989,N_23600,N_23405);
nand UO_2990 (O_2990,N_23926,N_24038);
xnor UO_2991 (O_2991,N_24735,N_24822);
nand UO_2992 (O_2992,N_24854,N_23444);
nor UO_2993 (O_2993,N_23054,N_23409);
and UO_2994 (O_2994,N_22135,N_24268);
nor UO_2995 (O_2995,N_22572,N_24566);
or UO_2996 (O_2996,N_24598,N_24303);
nand UO_2997 (O_2997,N_23784,N_22434);
and UO_2998 (O_2998,N_24477,N_23598);
nor UO_2999 (O_2999,N_24697,N_22004);
endmodule