module basic_2500_25000_3000_5_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1411,In_2058);
nor U1 (N_1,In_450,In_1700);
or U2 (N_2,In_704,In_413);
nor U3 (N_3,In_1882,In_344);
nor U4 (N_4,In_756,In_2296);
or U5 (N_5,In_460,In_1526);
xnor U6 (N_6,In_1704,In_707);
nor U7 (N_7,In_1253,In_1810);
nand U8 (N_8,In_1190,In_1494);
or U9 (N_9,In_741,In_865);
xor U10 (N_10,In_1500,In_2235);
or U11 (N_11,In_1866,In_5);
xnor U12 (N_12,In_28,In_1556);
and U13 (N_13,In_1375,In_1309);
nor U14 (N_14,In_877,In_404);
or U15 (N_15,In_2242,In_899);
or U16 (N_16,In_1199,In_1127);
or U17 (N_17,In_576,In_579);
and U18 (N_18,In_212,In_302);
and U19 (N_19,In_1907,In_2199);
nor U20 (N_20,In_112,In_128);
nand U21 (N_21,In_1489,In_2366);
nand U22 (N_22,In_1240,In_306);
nand U23 (N_23,In_407,In_1481);
nand U24 (N_24,In_2267,In_233);
or U25 (N_25,In_1705,In_674);
nor U26 (N_26,In_292,In_816);
or U27 (N_27,In_2153,In_263);
nand U28 (N_28,In_2364,In_13);
or U29 (N_29,In_2196,In_1543);
and U30 (N_30,In_879,In_626);
nand U31 (N_31,In_1498,In_2100);
nand U32 (N_32,In_2405,In_716);
and U33 (N_33,In_1044,In_1069);
or U34 (N_34,In_571,In_2390);
nand U35 (N_35,In_804,In_36);
or U36 (N_36,In_1809,In_914);
nor U37 (N_37,In_1643,In_1008);
nand U38 (N_38,In_922,In_1848);
nand U39 (N_39,In_1460,In_1890);
xnor U40 (N_40,In_102,In_2461);
and U41 (N_41,In_157,In_2229);
or U42 (N_42,In_1263,In_1847);
and U43 (N_43,In_1875,In_1785);
nor U44 (N_44,In_1086,In_1400);
nand U45 (N_45,In_1287,In_2457);
nand U46 (N_46,In_1145,In_875);
and U47 (N_47,In_313,In_377);
xor U48 (N_48,In_1657,In_791);
nand U49 (N_49,In_1827,In_1153);
nor U50 (N_50,In_1037,In_949);
nand U51 (N_51,In_621,In_1858);
or U52 (N_52,In_2142,In_1738);
and U53 (N_53,In_1349,In_1800);
or U54 (N_54,In_1773,In_170);
and U55 (N_55,In_1404,In_2228);
xnor U56 (N_56,In_316,In_2059);
nand U57 (N_57,In_1169,In_2175);
nor U58 (N_58,In_1225,In_1049);
nor U59 (N_59,In_1530,In_57);
or U60 (N_60,In_662,In_146);
or U61 (N_61,In_902,In_1805);
or U62 (N_62,In_758,In_1916);
or U63 (N_63,In_518,In_2474);
and U64 (N_64,In_1832,In_1947);
or U65 (N_65,In_2408,In_1651);
or U66 (N_66,In_98,In_2038);
nand U67 (N_67,In_893,In_1293);
or U68 (N_68,In_1139,In_1811);
and U69 (N_69,In_582,In_2265);
nand U70 (N_70,In_2037,In_1621);
nand U71 (N_71,In_779,In_1959);
nand U72 (N_72,In_2389,In_2429);
nor U73 (N_73,In_2083,In_1568);
or U74 (N_74,In_2039,In_1041);
and U75 (N_75,In_2013,In_2383);
and U76 (N_76,In_1697,In_1024);
or U77 (N_77,In_417,In_2092);
xnor U78 (N_78,In_1908,In_1217);
nor U79 (N_79,In_1173,In_1960);
or U80 (N_80,In_960,In_1103);
nand U81 (N_81,In_2171,In_551);
nor U82 (N_82,In_507,In_288);
and U83 (N_83,In_1678,In_1874);
nand U84 (N_84,In_947,In_371);
or U85 (N_85,In_1633,In_1906);
nand U86 (N_86,In_863,In_19);
nand U87 (N_87,In_1516,In_132);
and U88 (N_88,In_2041,In_1646);
nand U89 (N_89,In_1572,In_437);
nand U90 (N_90,In_1424,In_1446);
or U91 (N_91,In_1248,In_1979);
nor U92 (N_92,In_1609,In_1383);
or U93 (N_93,In_750,In_352);
and U94 (N_94,In_712,In_1444);
nor U95 (N_95,In_355,In_2019);
and U96 (N_96,In_1904,In_1788);
xnor U97 (N_97,In_1414,In_362);
xor U98 (N_98,In_2317,In_1687);
and U99 (N_99,In_933,In_408);
xnor U100 (N_100,In_1204,In_732);
or U101 (N_101,In_1186,In_1701);
or U102 (N_102,In_347,In_1155);
and U103 (N_103,In_121,In_1246);
xnor U104 (N_104,In_249,In_841);
and U105 (N_105,In_443,In_1455);
xnor U106 (N_106,In_1611,In_2146);
or U107 (N_107,In_1459,In_1698);
nand U108 (N_108,In_1891,In_2177);
nor U109 (N_109,In_1470,In_2414);
or U110 (N_110,In_1073,In_1294);
and U111 (N_111,In_673,In_106);
nor U112 (N_112,In_220,In_2481);
nand U113 (N_113,In_1421,In_1883);
and U114 (N_114,In_1903,In_929);
nor U115 (N_115,In_1931,In_1967);
and U116 (N_116,In_2201,In_1275);
nor U117 (N_117,In_62,In_1946);
or U118 (N_118,In_1072,In_2376);
and U119 (N_119,In_1365,In_1971);
or U120 (N_120,In_300,In_1117);
and U121 (N_121,In_583,In_1791);
and U122 (N_122,In_1793,In_1571);
nand U123 (N_123,In_1055,In_1822);
and U124 (N_124,In_1099,In_1438);
nand U125 (N_125,In_1221,In_2469);
and U126 (N_126,In_1047,In_1540);
xnor U127 (N_127,In_1005,In_1084);
and U128 (N_128,In_1867,In_801);
or U129 (N_129,In_2157,In_1815);
nor U130 (N_130,In_1708,In_1951);
or U131 (N_131,In_2277,In_410);
xor U132 (N_132,In_764,In_494);
xor U133 (N_133,In_993,In_2378);
nand U134 (N_134,In_1723,In_755);
nor U135 (N_135,In_2188,In_130);
nor U136 (N_136,In_314,In_787);
nand U137 (N_137,In_1770,In_1237);
nand U138 (N_138,In_2377,In_980);
nand U139 (N_139,In_1080,In_612);
nand U140 (N_140,In_2118,In_2096);
nand U141 (N_141,In_322,In_3);
or U142 (N_142,In_452,In_2238);
nand U143 (N_143,In_1388,In_620);
and U144 (N_144,In_1988,In_427);
xor U145 (N_145,In_984,In_2154);
nor U146 (N_146,In_881,In_2491);
or U147 (N_147,In_399,In_70);
or U148 (N_148,In_80,In_340);
and U149 (N_149,In_1000,In_825);
and U150 (N_150,In_645,In_2221);
or U151 (N_151,In_796,In_1549);
or U152 (N_152,In_1391,In_891);
nand U153 (N_153,In_1046,In_1012);
nand U154 (N_154,In_2093,In_651);
nor U155 (N_155,In_2424,In_2126);
nor U156 (N_156,In_2033,In_1652);
nand U157 (N_157,In_2324,In_1417);
nand U158 (N_158,In_2095,In_930);
nor U159 (N_159,In_1566,In_1197);
nor U160 (N_160,In_2163,In_1545);
and U161 (N_161,In_374,In_545);
nand U162 (N_162,In_1667,In_574);
nor U163 (N_163,In_2478,In_1283);
nand U164 (N_164,In_2453,In_2187);
nand U165 (N_165,In_2403,In_1504);
and U166 (N_166,In_393,In_1022);
xnor U167 (N_167,In_990,In_1838);
xnor U168 (N_168,In_2328,In_1081);
and U169 (N_169,In_1288,In_231);
nor U170 (N_170,In_2371,In_1653);
nand U171 (N_171,In_2288,In_2050);
or U172 (N_172,In_1096,In_1920);
or U173 (N_173,In_92,In_222);
and U174 (N_174,In_1168,In_15);
or U175 (N_175,In_1050,In_1250);
and U176 (N_176,In_21,In_2011);
xnor U177 (N_177,In_2073,In_108);
nor U178 (N_178,In_1662,In_1614);
xnor U179 (N_179,In_861,In_2477);
or U180 (N_180,In_466,In_46);
nor U181 (N_181,In_2003,In_96);
xor U182 (N_182,In_859,In_189);
xnor U183 (N_183,In_1062,In_1772);
or U184 (N_184,In_800,In_2111);
nand U185 (N_185,In_1813,In_822);
or U186 (N_186,In_2483,In_1974);
nand U187 (N_187,In_1991,In_118);
and U188 (N_188,In_2295,In_857);
xor U189 (N_189,In_2244,In_1843);
and U190 (N_190,In_2005,In_2079);
nor U191 (N_191,In_2113,In_2393);
nand U192 (N_192,In_356,In_549);
and U193 (N_193,In_1059,In_1987);
nand U194 (N_194,In_2460,In_686);
nand U195 (N_195,In_752,In_2070);
or U196 (N_196,In_584,In_1745);
nor U197 (N_197,In_1681,In_2203);
xor U198 (N_198,In_1669,In_2140);
nand U199 (N_199,In_2313,In_2074);
nor U200 (N_200,In_1527,In_987);
nand U201 (N_201,In_1380,In_2386);
and U202 (N_202,In_1921,In_1165);
nand U203 (N_203,In_2125,In_2127);
or U204 (N_204,In_1606,In_1851);
or U205 (N_205,In_25,In_196);
and U206 (N_206,In_1006,In_522);
or U207 (N_207,In_2042,In_762);
or U208 (N_208,In_1660,In_1803);
and U209 (N_209,In_2489,In_2485);
or U210 (N_210,In_163,In_1241);
nand U211 (N_211,In_766,In_597);
nand U212 (N_212,In_634,In_1267);
nand U213 (N_213,In_1277,In_958);
or U214 (N_214,In_1258,In_1247);
nor U215 (N_215,In_2078,In_640);
or U216 (N_216,In_2261,In_1854);
nor U217 (N_217,In_2048,In_2069);
and U218 (N_218,In_2433,In_2446);
and U219 (N_219,In_595,In_2129);
xor U220 (N_220,In_1136,In_1881);
nand U221 (N_221,In_363,In_324);
xnor U222 (N_222,In_649,In_2448);
nor U223 (N_223,In_1079,In_1483);
nand U224 (N_224,In_653,In_1842);
nand U225 (N_225,In_1475,In_2466);
and U226 (N_226,In_1964,In_2475);
nand U227 (N_227,In_412,In_126);
or U228 (N_228,In_820,In_892);
or U229 (N_229,In_191,In_1725);
nand U230 (N_230,In_400,In_2077);
nand U231 (N_231,In_1496,In_525);
or U232 (N_232,In_166,In_911);
nor U233 (N_233,In_1422,In_424);
nor U234 (N_234,In_100,In_1397);
nand U235 (N_235,In_244,In_124);
nor U236 (N_236,In_1354,In_1271);
nor U237 (N_237,In_216,In_1392);
and U238 (N_238,In_71,In_725);
or U239 (N_239,In_1410,In_1943);
and U240 (N_240,In_229,In_623);
or U241 (N_241,In_438,In_2174);
or U242 (N_242,In_1473,In_1063);
and U243 (N_243,In_1347,In_1913);
nor U244 (N_244,In_659,In_1990);
xor U245 (N_245,In_2028,In_2391);
or U246 (N_246,In_1185,In_1739);
and U247 (N_247,In_546,In_1597);
and U248 (N_248,In_617,In_1213);
nand U249 (N_249,In_966,In_1747);
xnor U250 (N_250,In_1023,In_591);
or U251 (N_251,In_2076,In_1781);
nand U252 (N_252,In_678,In_160);
or U253 (N_253,In_2331,In_768);
or U254 (N_254,In_1799,In_670);
xnor U255 (N_255,In_1887,In_1447);
nor U256 (N_256,In_461,In_1761);
or U257 (N_257,In_839,In_786);
or U258 (N_258,In_1149,In_543);
xor U259 (N_259,In_565,In_1176);
nand U260 (N_260,In_33,In_1450);
nand U261 (N_261,In_2200,In_1039);
or U262 (N_262,In_1366,In_468);
xor U263 (N_263,In_2394,In_480);
or U264 (N_264,In_473,In_981);
nand U265 (N_265,In_22,In_1111);
and U266 (N_266,In_2392,In_1715);
xor U267 (N_267,In_1521,In_137);
nor U268 (N_268,In_2418,In_1860);
and U269 (N_269,In_533,In_116);
and U270 (N_270,In_2164,In_1939);
and U271 (N_271,In_2495,In_2071);
nor U272 (N_272,In_2266,In_1020);
xor U273 (N_273,In_1311,In_2349);
nand U274 (N_274,In_1409,In_593);
or U275 (N_275,In_1290,In_599);
or U276 (N_276,In_2099,In_378);
nand U277 (N_277,In_1488,In_150);
and U278 (N_278,In_323,In_1709);
or U279 (N_279,In_589,In_269);
nand U280 (N_280,In_1721,In_1192);
xnor U281 (N_281,In_873,In_75);
and U282 (N_282,In_2497,In_1735);
or U283 (N_283,In_304,In_1817);
nor U284 (N_284,In_763,In_996);
xor U285 (N_285,In_199,In_1299);
nand U286 (N_286,In_293,In_742);
and U287 (N_287,In_1742,In_299);
and U288 (N_288,In_421,In_1120);
or U289 (N_289,In_2442,In_1930);
or U290 (N_290,In_2316,In_1905);
nor U291 (N_291,In_896,In_813);
xor U292 (N_292,In_1323,In_1028);
and U293 (N_293,In_1075,In_2462);
and U294 (N_294,In_259,In_1528);
or U295 (N_295,In_88,In_1749);
or U296 (N_296,In_1638,In_2252);
xor U297 (N_297,In_122,In_1087);
nand U298 (N_298,In_1717,In_1485);
or U299 (N_299,In_1324,In_1257);
nand U300 (N_300,In_1352,In_226);
or U301 (N_301,In_1702,In_1302);
xnor U302 (N_302,In_44,In_1398);
nor U303 (N_303,In_349,In_1802);
nand U304 (N_304,In_925,In_775);
and U305 (N_305,In_17,In_217);
and U306 (N_306,In_1327,In_1463);
and U307 (N_307,In_2212,In_552);
xnor U308 (N_308,In_1834,In_1682);
nor U309 (N_309,In_2130,In_1477);
nand U310 (N_310,In_2152,In_1506);
and U311 (N_311,In_1367,In_824);
nor U312 (N_312,In_1910,In_602);
and U313 (N_313,In_78,In_1112);
and U314 (N_314,In_2415,In_1448);
nand U315 (N_315,In_72,In_928);
nor U316 (N_316,In_447,In_1515);
nor U317 (N_317,In_713,In_275);
or U318 (N_318,In_1379,In_1840);
xor U319 (N_319,In_2087,In_1816);
xnor U320 (N_320,In_1591,In_2009);
nand U321 (N_321,In_1401,In_2309);
or U322 (N_322,In_353,In_2344);
nand U323 (N_323,In_2305,In_140);
nor U324 (N_324,In_245,In_2421);
nand U325 (N_325,In_1592,In_2339);
and U326 (N_326,In_1849,In_1292);
and U327 (N_327,In_1178,In_702);
nor U328 (N_328,In_1406,In_253);
nor U329 (N_329,In_982,In_272);
and U330 (N_330,In_335,In_1989);
xnor U331 (N_331,In_167,In_328);
nor U332 (N_332,In_1694,In_303);
and U333 (N_333,In_1403,In_1035);
nor U334 (N_334,In_992,In_1599);
and U335 (N_335,In_1360,In_611);
or U336 (N_336,In_773,In_1937);
xnor U337 (N_337,In_708,In_1466);
and U338 (N_338,In_476,In_1334);
and U339 (N_339,In_37,In_2131);
and U340 (N_340,In_370,In_1227);
nor U341 (N_341,In_345,In_2214);
nand U342 (N_342,In_2427,In_1465);
and U343 (N_343,In_2490,In_1886);
nor U344 (N_344,In_1808,In_359);
nor U345 (N_345,In_920,In_828);
or U346 (N_346,In_1452,In_1707);
or U347 (N_347,In_1868,In_793);
or U348 (N_348,In_1985,In_1582);
nor U349 (N_349,In_1172,In_1656);
xnor U350 (N_350,In_711,In_1272);
or U351 (N_351,In_842,In_1513);
nand U352 (N_352,In_321,In_557);
xnor U353 (N_353,In_474,In_1839);
nand U354 (N_354,In_405,In_529);
nor U355 (N_355,In_1436,In_320);
or U356 (N_356,In_1115,In_1699);
nand U357 (N_357,In_1342,In_1612);
and U358 (N_358,In_843,In_1231);
and U359 (N_359,In_829,In_1353);
xnor U360 (N_360,In_1390,In_504);
nand U361 (N_361,In_93,In_1297);
xor U362 (N_362,In_1680,In_1563);
and U363 (N_363,In_1376,In_1659);
and U364 (N_364,In_650,In_2271);
xor U365 (N_365,In_213,In_778);
and U366 (N_366,In_32,In_1986);
xnor U367 (N_367,In_1018,In_1420);
or U368 (N_368,In_700,In_561);
and U369 (N_369,In_2167,In_2144);
nand U370 (N_370,In_42,In_580);
nand U371 (N_371,In_182,In_117);
nand U372 (N_372,In_1100,In_1546);
xor U373 (N_373,In_1983,In_1285);
and U374 (N_374,In_1266,In_2206);
nor U375 (N_375,In_1203,In_684);
or U376 (N_376,In_1507,In_1378);
nor U377 (N_377,In_2239,In_1647);
and U378 (N_378,In_1917,In_740);
nor U379 (N_379,In_680,In_722);
nor U380 (N_380,In_2444,In_1544);
or U381 (N_381,In_2148,In_1357);
nand U382 (N_382,In_1596,In_605);
nor U383 (N_383,In_1892,In_156);
nand U384 (N_384,In_2124,In_995);
nor U385 (N_385,In_2255,In_1620);
xor U386 (N_386,In_569,In_1751);
nand U387 (N_387,In_2101,In_596);
and U388 (N_388,In_1377,In_777);
nand U389 (N_389,In_310,In_1083);
nor U390 (N_390,In_530,In_1567);
and U391 (N_391,In_2186,In_127);
and U392 (N_392,In_848,In_811);
xor U393 (N_393,In_1634,In_1273);
and U394 (N_394,In_2089,In_45);
or U395 (N_395,In_2227,In_479);
and U396 (N_396,In_2346,In_1013);
nor U397 (N_397,In_202,In_637);
xor U398 (N_398,In_1181,In_181);
nand U399 (N_399,In_1101,In_221);
and U400 (N_400,In_1131,In_1141);
nor U401 (N_401,In_1233,In_63);
nand U402 (N_402,In_587,In_658);
nand U403 (N_403,In_433,In_878);
xnor U404 (N_404,In_481,In_721);
nor U405 (N_405,In_1286,In_368);
xnor U406 (N_406,In_2236,In_1753);
xnor U407 (N_407,In_2417,In_2117);
and U408 (N_408,In_2343,In_588);
or U409 (N_409,In_1889,In_469);
xnor U410 (N_410,In_586,In_1955);
and U411 (N_411,In_301,In_581);
nand U412 (N_412,In_1262,In_343);
nand U413 (N_413,In_1748,In_1108);
and U414 (N_414,In_1278,In_1956);
or U415 (N_415,In_553,In_1763);
nor U416 (N_416,In_1664,In_1689);
or U417 (N_417,In_1641,In_2425);
or U418 (N_418,In_1994,In_1161);
xor U419 (N_419,In_120,In_2456);
nor U420 (N_420,In_615,In_1551);
or U421 (N_421,In_2381,In_532);
or U422 (N_422,In_754,In_175);
and U423 (N_423,In_74,In_1274);
or U424 (N_424,In_904,In_1457);
nand U425 (N_425,In_1661,In_1301);
nand U426 (N_426,In_2254,In_197);
nor U427 (N_427,In_1160,In_698);
nor U428 (N_428,In_2159,In_386);
xnor U429 (N_429,In_446,In_1045);
nor U430 (N_430,In_523,In_205);
xor U431 (N_431,In_2122,In_2396);
and U432 (N_432,In_190,In_592);
nor U433 (N_433,In_155,In_1026);
nand U434 (N_434,In_1997,In_1512);
nand U435 (N_435,In_333,In_1195);
and U436 (N_436,In_1432,In_1758);
and U437 (N_437,In_2043,In_1518);
or U438 (N_438,In_1415,In_2385);
or U439 (N_439,In_1663,In_2054);
nand U440 (N_440,In_1553,In_1893);
and U441 (N_441,In_1603,In_1928);
or U442 (N_442,In_1322,In_414);
xor U443 (N_443,In_1533,In_2097);
nand U444 (N_444,In_1236,In_2367);
and U445 (N_445,In_657,In_1109);
nor U446 (N_446,In_1374,In_1878);
nor U447 (N_447,In_2247,In_1268);
or U448 (N_448,In_1590,In_977);
nand U449 (N_449,In_1501,In_2310);
xor U450 (N_450,In_2323,In_2270);
xnor U451 (N_451,In_1066,In_724);
nor U452 (N_452,In_578,In_1784);
nor U453 (N_453,In_517,In_2289);
and U454 (N_454,In_1071,In_51);
xnor U455 (N_455,In_897,In_1674);
xor U456 (N_456,In_429,In_1980);
nand U457 (N_457,In_1829,In_2325);
and U458 (N_458,In_968,In_1065);
nand U459 (N_459,In_1778,In_2493);
nand U460 (N_460,In_864,In_153);
or U461 (N_461,In_910,In_1757);
or U462 (N_462,In_2134,In_2185);
or U463 (N_463,In_998,In_1831);
or U464 (N_464,In_465,In_2220);
nor U465 (N_465,In_2222,In_944);
or U466 (N_466,In_1695,In_805);
xnor U467 (N_467,In_745,In_2435);
xor U468 (N_468,In_2399,In_2213);
nor U469 (N_469,In_2355,In_43);
nor U470 (N_470,In_2436,In_2193);
nand U471 (N_471,In_1156,In_1317);
or U472 (N_472,In_2018,In_885);
and U473 (N_473,In_56,In_81);
and U474 (N_474,In_236,In_723);
xnor U475 (N_475,In_1325,In_2025);
nand U476 (N_476,In_1525,In_2350);
or U477 (N_477,In_90,In_261);
xnor U478 (N_478,In_798,In_308);
xnor U479 (N_479,In_206,In_2158);
nor U480 (N_480,In_1593,In_366);
nor U481 (N_481,In_854,In_2368);
or U482 (N_482,In_431,In_2307);
or U483 (N_483,In_161,In_1077);
or U484 (N_484,In_751,In_139);
and U485 (N_485,In_2075,In_2285);
or U486 (N_486,In_1295,In_6);
xor U487 (N_487,In_230,In_270);
xnor U488 (N_488,In_1394,In_2291);
nand U489 (N_489,In_2432,In_1002);
nand U490 (N_490,In_1595,In_607);
or U491 (N_491,In_1794,In_2308);
nor U492 (N_492,In_1522,In_1497);
or U493 (N_493,In_1925,In_105);
or U494 (N_494,In_979,In_2135);
or U495 (N_495,In_66,In_2387);
and U496 (N_496,In_2063,In_1355);
nand U497 (N_497,In_188,In_2401);
nand U498 (N_498,In_671,In_1484);
or U499 (N_499,In_883,In_1058);
and U500 (N_500,In_1205,In_2443);
and U501 (N_501,In_281,In_554);
and U502 (N_502,In_1345,In_2176);
and U503 (N_503,In_224,In_458);
xor U504 (N_504,In_1003,In_1942);
xor U505 (N_505,In_2428,In_731);
nor U506 (N_506,In_2149,In_1416);
and U507 (N_507,In_871,In_869);
nor U508 (N_508,In_1613,In_2216);
and U509 (N_509,In_1885,In_1057);
xnor U510 (N_510,In_1637,In_60);
nor U511 (N_511,In_989,In_2298);
nand U512 (N_512,In_627,In_1855);
or U513 (N_513,In_1836,In_1922);
or U514 (N_514,In_860,In_2114);
nor U515 (N_515,In_403,In_179);
nor U516 (N_516,In_1509,In_1439);
nor U517 (N_517,In_309,In_1395);
xor U518 (N_518,In_939,In_67);
xnor U519 (N_519,In_247,In_1629);
or U520 (N_520,In_1321,In_512);
nor U521 (N_521,In_2061,In_1147);
nor U522 (N_522,In_1179,In_1537);
or U523 (N_523,In_12,In_2333);
and U524 (N_524,In_1102,In_1534);
and U525 (N_525,In_2249,In_1706);
nor U526 (N_526,In_952,In_2494);
nand U527 (N_527,In_1636,In_1193);
nor U528 (N_528,In_398,In_1965);
and U529 (N_529,In_257,In_1232);
or U530 (N_530,In_1146,In_943);
or U531 (N_531,In_242,In_1766);
and U532 (N_532,In_2106,In_2312);
nor U533 (N_533,In_886,In_2332);
and U534 (N_534,In_1671,In_959);
nor U535 (N_535,In_1625,In_1780);
and U536 (N_536,In_1070,In_1038);
xnor U537 (N_537,In_1399,In_192);
nor U538 (N_538,In_903,In_397);
xnor U539 (N_539,In_1618,In_1110);
and U540 (N_540,In_1648,In_706);
nand U541 (N_541,In_890,In_2303);
nand U542 (N_542,In_462,In_681);
nor U543 (N_543,In_567,In_1932);
nand U544 (N_544,In_214,In_1196);
nor U545 (N_545,In_1710,In_1873);
or U546 (N_546,In_2015,In_287);
and U547 (N_547,In_2210,In_2006);
and U548 (N_548,In_456,In_683);
xnor U549 (N_549,In_1269,In_1339);
xor U550 (N_550,In_1152,In_1654);
or U551 (N_551,In_174,In_1790);
nand U552 (N_552,In_1209,In_538);
nor U553 (N_553,In_2225,In_1116);
and U554 (N_554,In_351,In_2055);
nor U555 (N_555,In_2172,In_1030);
nor U556 (N_556,In_1622,In_830);
nand U557 (N_557,In_1783,In_1759);
nor U558 (N_558,In_639,In_2360);
xnor U559 (N_559,In_2022,In_1557);
nand U560 (N_560,In_646,In_1245);
nand U561 (N_561,In_61,In_84);
or U562 (N_562,In_1467,In_1604);
and U563 (N_563,In_2029,In_1076);
xor U564 (N_564,In_738,In_1754);
xor U565 (N_565,In_537,In_1740);
xnor U566 (N_566,In_2180,In_383);
nor U567 (N_567,In_2147,In_2208);
and U568 (N_568,In_1769,In_1996);
or U569 (N_569,In_1220,In_1594);
or U570 (N_570,In_1589,In_2351);
or U571 (N_571,In_380,In_138);
nand U572 (N_572,In_874,In_1480);
xnor U573 (N_573,In_1021,In_1777);
xor U574 (N_574,In_2231,In_564);
nor U575 (N_575,In_280,In_1216);
or U576 (N_576,In_95,In_1993);
or U577 (N_577,In_496,In_1348);
and U578 (N_578,In_1623,In_912);
xor U579 (N_579,In_159,In_2281);
or U580 (N_580,In_1341,In_1054);
nand U581 (N_581,In_1975,In_2358);
nor U582 (N_582,In_638,In_1555);
nand U583 (N_583,In_1163,In_635);
nor U584 (N_584,In_2045,In_1775);
nor U585 (N_585,In_967,In_1315);
and U586 (N_586,In_1313,In_660);
and U587 (N_587,In_136,In_1871);
nand U588 (N_588,In_2151,In_2240);
and U589 (N_589,In_82,In_1060);
nand U590 (N_590,In_2141,In_1126);
nor U591 (N_591,In_425,In_1476);
or U592 (N_592,In_1413,In_855);
nor U593 (N_593,In_2260,In_265);
nand U594 (N_594,In_50,In_1091);
xnor U595 (N_595,In_1043,In_2470);
xnor U596 (N_596,In_194,In_2353);
nand U597 (N_597,In_1536,In_331);
or U598 (N_598,In_1356,In_248);
nor U599 (N_599,In_2487,In_1732);
or U600 (N_600,In_125,In_743);
nand U601 (N_601,In_204,In_382);
or U602 (N_602,In_511,In_2098);
nand U603 (N_603,In_923,In_85);
and U604 (N_604,In_1692,In_1135);
nand U605 (N_605,In_1106,In_2123);
nand U606 (N_606,In_817,In_285);
and U607 (N_607,In_760,In_1159);
nand U608 (N_608,In_1482,In_379);
nor U609 (N_609,In_1212,In_1679);
xnor U610 (N_610,In_264,In_2060);
xor U611 (N_611,In_2384,In_2411);
or U612 (N_612,In_83,In_185);
xor U613 (N_613,In_158,In_2463);
nor U614 (N_614,In_485,In_2430);
xnor U615 (N_615,In_880,In_935);
or U616 (N_616,In_629,In_1923);
and U617 (N_617,In_336,In_709);
or U618 (N_618,In_243,In_260);
or U619 (N_619,In_2459,In_2088);
nand U620 (N_620,In_195,In_1412);
xnor U621 (N_621,In_1737,In_2091);
nand U622 (N_622,In_327,In_1564);
or U623 (N_623,In_2363,In_2287);
xor U624 (N_624,In_459,In_2192);
nand U625 (N_625,In_1449,In_296);
nand U626 (N_626,In_536,In_2388);
nand U627 (N_627,In_1559,In_2482);
nor U628 (N_628,In_1626,In_1550);
and U629 (N_629,In_1952,In_631);
xor U630 (N_630,In_1547,In_1255);
or U631 (N_631,In_625,In_1495);
xnor U632 (N_632,In_2110,In_1862);
nand U633 (N_633,In_311,In_1015);
and U634 (N_634,In_436,In_1132);
or U635 (N_635,In_1469,In_2027);
or U636 (N_636,In_1598,In_815);
nand U637 (N_637,In_853,In_759);
xor U638 (N_638,In_267,In_570);
or U639 (N_639,In_1092,In_426);
and U640 (N_640,In_1142,In_1981);
or U641 (N_641,In_2062,In_2374);
nand U642 (N_642,In_2105,In_326);
xor U643 (N_643,In_164,In_2282);
nor U644 (N_644,In_2286,In_2189);
nand U645 (N_645,In_556,In_2440);
nand U646 (N_646,In_2280,In_2000);
nor U647 (N_647,In_1686,In_2);
and U648 (N_648,In_1499,In_664);
xor U649 (N_649,In_1427,In_965);
and U650 (N_650,In_2334,In_2036);
or U651 (N_651,In_970,In_974);
and U652 (N_652,In_1014,In_1787);
nand U653 (N_653,In_703,In_332);
and U654 (N_654,In_887,In_273);
or U655 (N_655,In_1655,In_2357);
or U656 (N_656,In_1260,In_388);
nand U657 (N_657,In_1472,In_614);
or U658 (N_658,In_2292,In_346);
xnor U659 (N_659,In_152,In_516);
and U660 (N_660,In_113,In_2329);
and U661 (N_661,In_2416,In_1458);
or U662 (N_662,In_894,In_1175);
nand U663 (N_663,In_2365,In_1558);
and U664 (N_664,In_2452,In_271);
or U665 (N_665,In_610,In_1426);
nor U666 (N_666,In_2207,In_2166);
or U667 (N_667,In_99,In_1337);
nand U668 (N_668,In_1456,In_1306);
nor U669 (N_669,In_603,In_500);
nor U670 (N_670,In_1097,In_1927);
nand U671 (N_671,In_16,In_1121);
xnor U672 (N_672,In_1768,In_1381);
nor U673 (N_673,In_1284,In_1605);
or U674 (N_674,In_2311,In_223);
nor U675 (N_675,In_1453,In_402);
nor U676 (N_676,In_1343,In_1093);
nor U677 (N_677,In_598,In_1486);
and U678 (N_678,In_1818,In_1896);
nor U679 (N_679,In_1252,In_0);
or U680 (N_680,In_836,In_938);
xnor U681 (N_681,In_1256,In_616);
nand U682 (N_682,In_2471,In_515);
xnor U683 (N_683,In_2107,In_1650);
xnor U684 (N_684,In_797,In_357);
and U685 (N_685,In_2090,In_808);
and U686 (N_686,In_1333,In_2184);
xor U687 (N_687,In_973,In_1542);
or U688 (N_688,In_2081,In_1688);
nor U689 (N_689,In_2215,In_2115);
and U690 (N_690,In_2356,In_632);
or U691 (N_691,In_1428,In_1082);
nand U692 (N_692,In_2085,In_1649);
xnor U693 (N_693,In_1814,In_2336);
nand U694 (N_694,In_394,In_2066);
xnor U695 (N_695,In_2498,In_688);
xnor U696 (N_696,In_1580,In_656);
xnor U697 (N_697,In_685,In_905);
nand U698 (N_698,In_1856,In_390);
or U699 (N_699,In_444,In_774);
or U700 (N_700,In_1167,In_2173);
nand U701 (N_701,In_2315,In_1451);
and U702 (N_702,In_2318,In_341);
and U703 (N_703,In_1462,In_1776);
xor U704 (N_704,In_1396,In_1510);
and U705 (N_705,In_643,In_2064);
and U706 (N_706,In_1369,In_1329);
and U707 (N_707,In_279,In_1191);
nand U708 (N_708,In_696,In_1307);
nor U709 (N_709,In_1418,In_1251);
nor U710 (N_710,In_1870,In_1051);
or U711 (N_711,In_1812,In_1264);
and U712 (N_712,In_558,In_2275);
and U713 (N_713,In_171,In_1548);
xnor U714 (N_714,In_477,In_1201);
or U715 (N_715,In_1902,In_1405);
xnor U716 (N_716,In_812,In_420);
nand U717 (N_717,In_1491,In_373);
nor U718 (N_718,In_945,In_719);
xor U719 (N_719,In_1644,In_1249);
nand U720 (N_720,In_1880,In_1140);
xor U721 (N_721,In_365,In_1950);
xnor U722 (N_722,In_844,In_1958);
nor U723 (N_723,In_64,In_434);
nand U724 (N_724,In_1561,In_2072);
and U725 (N_725,In_2031,In_1143);
xnor U726 (N_726,In_168,In_1616);
nand U727 (N_727,In_1230,In_502);
and U728 (N_728,In_1279,In_482);
or U729 (N_729,In_1177,In_489);
nand U730 (N_730,In_2293,In_521);
and U731 (N_731,In_1579,In_988);
and U732 (N_732,In_1969,In_868);
nor U733 (N_733,In_765,In_2273);
or U734 (N_734,In_2301,In_1852);
nor U735 (N_735,In_94,In_409);
nor U736 (N_736,In_1801,In_2297);
or U737 (N_737,In_2084,In_1578);
nand U738 (N_738,In_601,In_1628);
nor U739 (N_739,In_720,In_2341);
xor U740 (N_740,In_802,In_675);
and U741 (N_741,In_1305,In_232);
nor U742 (N_742,In_2250,In_1119);
and U743 (N_743,In_789,In_2001);
nor U744 (N_744,In_1876,In_361);
or U745 (N_745,In_2195,In_2165);
xor U746 (N_746,In_2080,In_1011);
and U747 (N_747,In_1954,In_1085);
nor U748 (N_748,In_7,In_889);
and U749 (N_749,In_2181,In_187);
and U750 (N_750,In_503,In_1957);
nand U751 (N_751,In_2473,In_534);
nand U752 (N_752,In_1642,In_1034);
or U753 (N_753,In_177,In_1774);
nand U754 (N_754,In_1541,In_1133);
xor U755 (N_755,In_1304,In_198);
and U756 (N_756,In_1128,In_419);
nand U757 (N_757,In_757,In_814);
xnor U758 (N_758,In_364,In_767);
or U759 (N_759,In_1061,In_1207);
and U760 (N_760,In_1713,In_1373);
and U761 (N_761,In_1727,In_430);
or U762 (N_762,In_568,In_535);
and U763 (N_763,In_1435,In_2294);
xor U764 (N_764,In_2337,In_1210);
xor U765 (N_765,In_1915,In_73);
xor U766 (N_766,In_2467,In_104);
or U767 (N_767,In_2409,In_1632);
xor U768 (N_768,In_154,In_487);
or U769 (N_769,In_2268,In_1926);
nand U770 (N_770,In_728,In_1731);
nor U771 (N_771,In_484,In_832);
nor U772 (N_772,In_672,In_1479);
xor U773 (N_773,In_338,In_445);
or U774 (N_774,In_312,In_1254);
nand U775 (N_775,In_2455,In_133);
nand U776 (N_776,In_1819,In_1004);
nand U777 (N_777,In_1853,In_490);
nor U778 (N_778,In_1382,In_1042);
or U779 (N_779,In_946,In_2402);
nor U780 (N_780,In_1935,In_449);
nor U781 (N_781,In_1107,In_1123);
xnor U782 (N_782,In_866,In_1270);
or U783 (N_783,In_550,In_667);
and U784 (N_784,In_1171,In_734);
nand U785 (N_785,In_337,In_2103);
xor U786 (N_786,In_2082,In_964);
nand U787 (N_787,In_55,In_2302);
xor U788 (N_788,In_491,In_2338);
nor U789 (N_789,In_2419,In_951);
xnor U790 (N_790,In_548,In_307);
xor U791 (N_791,In_560,In_771);
or U792 (N_792,In_1344,In_1863);
xor U793 (N_793,In_2051,In_499);
or U794 (N_794,In_1529,In_1741);
or U795 (N_795,In_1570,In_2256);
and U796 (N_796,In_23,In_749);
and U797 (N_797,In_514,In_747);
xor U798 (N_798,In_1792,In_89);
and U799 (N_799,In_225,In_1431);
nand U800 (N_800,In_1425,In_1430);
and U801 (N_801,In_2304,In_210);
or U802 (N_802,In_668,In_2162);
xor U803 (N_803,In_2237,In_234);
nor U804 (N_804,In_2209,In_348);
nand U805 (N_805,In_1690,In_2253);
and U806 (N_806,In_58,In_1806);
nand U807 (N_807,In_692,In_1992);
and U808 (N_808,In_1338,In_1508);
or U809 (N_809,In_2211,In_145);
xor U810 (N_810,In_358,In_647);
xnor U811 (N_811,In_1976,In_1074);
xor U812 (N_812,In_957,In_2034);
and U813 (N_813,In_218,In_1973);
nor U814 (N_814,In_726,In_2035);
xnor U815 (N_815,In_2259,In_547);
xor U816 (N_816,In_453,In_1712);
and U817 (N_817,In_2410,In_1877);
and U818 (N_818,In_1408,In_276);
nand U819 (N_819,In_68,In_1869);
nand U820 (N_820,In_2191,In_1764);
xor U821 (N_821,In_1782,In_628);
nand U822 (N_822,In_415,In_526);
nor U823 (N_823,In_785,In_1936);
xor U824 (N_824,In_1734,In_18);
nor U825 (N_825,In_566,In_1068);
nor U826 (N_826,In_663,In_29);
and U827 (N_827,In_2057,In_2102);
xor U828 (N_828,In_1532,In_1531);
nor U829 (N_829,In_666,In_1474);
or U830 (N_830,In_983,In_1978);
or U831 (N_831,In_442,In_239);
xor U832 (N_832,In_1296,In_14);
nor U833 (N_833,In_2370,In_1821);
or U834 (N_834,In_2040,In_401);
or U835 (N_835,In_941,In_927);
and U836 (N_836,In_1691,In_385);
nor U837 (N_837,In_2128,In_2161);
xor U838 (N_838,In_2279,In_1461);
nand U839 (N_839,In_208,In_1335);
and U840 (N_840,In_2423,In_1441);
or U841 (N_841,In_618,In_1303);
or U842 (N_842,In_2008,In_1823);
and U843 (N_843,In_1067,In_1361);
xor U844 (N_844,In_2137,In_1610);
xor U845 (N_845,In_2046,In_701);
xnor U846 (N_846,In_369,In_342);
xor U847 (N_847,In_2007,In_2380);
xor U848 (N_848,In_143,In_147);
or U849 (N_849,In_1492,In_1238);
nor U850 (N_850,In_1223,In_2116);
xnor U851 (N_851,In_613,In_1511);
and U852 (N_852,In_2359,In_1385);
or U853 (N_853,In_744,In_2119);
or U854 (N_854,In_1864,In_1402);
or U855 (N_855,In_478,In_918);
nand U856 (N_856,In_375,In_852);
and U857 (N_857,In_40,In_391);
nand U858 (N_858,In_2169,In_186);
xor U859 (N_859,In_2439,In_954);
or U860 (N_860,In_1586,In_1350);
nand U861 (N_861,In_1025,In_1900);
xor U862 (N_862,In_510,In_1666);
and U863 (N_863,In_389,In_268);
and U864 (N_864,In_1844,In_1319);
and U865 (N_865,In_1235,In_2021);
nand U866 (N_866,In_1517,In_1901);
and U867 (N_867,In_2369,In_1114);
or U868 (N_868,In_2283,In_590);
nand U869 (N_869,In_1953,In_934);
xor U870 (N_870,In_821,In_2065);
xor U871 (N_871,In_609,In_513);
or U872 (N_872,In_2204,In_1585);
or U873 (N_873,In_1861,In_2434);
xnor U874 (N_874,In_1228,In_360);
nand U875 (N_875,In_572,In_1797);
and U876 (N_876,In_1089,In_876);
and U877 (N_877,In_950,In_803);
nor U878 (N_878,In_1804,In_1970);
and U879 (N_879,In_1575,In_2340);
xnor U880 (N_880,In_1144,In_1833);
nand U881 (N_881,In_4,In_1328);
and U882 (N_882,In_227,In_1961);
xnor U883 (N_883,In_1711,In_255);
and U884 (N_884,In_1031,In_1944);
and U885 (N_885,In_2373,In_783);
and U886 (N_886,In_241,In_178);
and U887 (N_887,In_1300,In_2322);
or U888 (N_888,In_2217,In_1372);
or U889 (N_889,In_2112,In_1442);
nor U890 (N_890,In_2016,In_493);
and U891 (N_891,In_455,In_1919);
xnor U892 (N_892,In_1029,In_418);
and U893 (N_893,In_2150,In_772);
or U894 (N_894,In_1948,In_2413);
nor U895 (N_895,In_49,In_1234);
and U896 (N_896,In_544,In_475);
and U897 (N_897,In_2284,In_1724);
and U898 (N_898,In_109,In_907);
nand U899 (N_899,In_1539,In_114);
nor U900 (N_900,In_806,In_238);
nor U901 (N_901,In_792,In_1577);
nor U902 (N_902,In_52,In_644);
nor U903 (N_903,In_2183,In_41);
or U904 (N_904,In_1716,In_851);
and U905 (N_905,In_823,In_169);
xor U906 (N_906,In_2246,In_1982);
xor U907 (N_907,In_2138,In_1677);
and U908 (N_908,In_1733,In_2190);
xor U909 (N_909,In_739,In_2182);
or U910 (N_910,In_807,In_142);
and U911 (N_911,In_2020,In_1576);
and U912 (N_912,In_2030,In_619);
xor U913 (N_913,In_1113,In_207);
xor U914 (N_914,In_294,In_1364);
or U915 (N_915,In_788,In_1909);
or U916 (N_916,In_2407,In_1166);
nand U917 (N_917,In_2342,In_1226);
nor U918 (N_918,In_677,In_1503);
or U919 (N_919,In_1588,In_1587);
and U920 (N_920,In_737,In_2395);
or U921 (N_921,In_27,In_2053);
xor U922 (N_922,In_2472,In_2262);
and U923 (N_923,In_882,In_180);
nor U924 (N_924,In_682,In_1850);
and U925 (N_925,In_2219,In_931);
nor U926 (N_926,In_20,In_395);
xor U927 (N_927,In_129,In_454);
nor U928 (N_928,In_1314,In_2326);
and U929 (N_929,In_648,In_1972);
or U930 (N_930,In_2449,In_1924);
xor U931 (N_931,In_940,In_1182);
xor U932 (N_932,In_838,In_2278);
and U933 (N_933,In_994,In_1857);
or U934 (N_934,In_291,In_483);
nor U935 (N_935,In_1796,In_283);
or U936 (N_936,In_520,In_1019);
xor U937 (N_937,In_506,In_856);
or U938 (N_938,In_1215,In_528);
nand U939 (N_939,In_1490,In_2108);
and U940 (N_940,In_1048,In_2404);
xor U941 (N_941,In_209,In_123);
or U942 (N_942,In_915,In_2347);
xor U943 (N_943,In_942,In_508);
nand U944 (N_944,In_111,In_470);
or U945 (N_945,In_1214,In_330);
xor U946 (N_946,In_1312,In_1726);
xnor U947 (N_947,In_898,In_325);
nor U948 (N_948,In_2178,In_641);
xor U949 (N_949,In_1326,In_2263);
and U950 (N_950,In_1998,In_661);
or U951 (N_951,In_1719,In_999);
xor U952 (N_952,In_1583,In_2230);
and U953 (N_953,In_1310,In_1407);
or U954 (N_954,In_790,In_246);
nor U955 (N_955,In_2014,In_2450);
nand U956 (N_956,In_79,In_1560);
or U957 (N_957,In_1514,In_286);
or U958 (N_958,In_1897,In_1798);
and U959 (N_959,In_1368,In_1703);
nand U960 (N_960,In_1265,In_1524);
or U961 (N_961,In_2314,In_1938);
nor U962 (N_962,In_2170,In_334);
nor U963 (N_963,In_1828,In_962);
xor U964 (N_964,In_695,In_1371);
and U965 (N_965,In_1846,In_1281);
xnor U966 (N_966,In_2032,In_416);
or U967 (N_967,In_2362,In_1098);
nand U968 (N_968,In_1929,In_562);
and U969 (N_969,In_1624,In_2321);
nor U970 (N_970,In_2012,In_1162);
nand U971 (N_971,In_467,In_2431);
and U972 (N_972,In_1242,In_827);
xor U973 (N_973,In_274,In_2133);
nand U974 (N_974,In_1440,In_1779);
xnor U975 (N_975,In_8,In_2348);
nand U976 (N_976,In_679,In_1899);
or U977 (N_977,In_1148,In_1502);
or U978 (N_978,In_486,In_2412);
nor U979 (N_979,In_2067,In_519);
and U980 (N_980,In_654,In_141);
nor U981 (N_981,In_1183,In_1911);
or U982 (N_982,In_1194,In_784);
or U983 (N_983,In_1478,In_1351);
xor U984 (N_984,In_1825,In_1468);
and U985 (N_985,In_1820,In_809);
xor U986 (N_986,In_1090,In_1138);
nor U987 (N_987,In_630,In_1918);
or U988 (N_988,In_1645,In_542);
or U989 (N_989,In_636,In_1150);
and U990 (N_990,In_727,In_406);
nor U991 (N_991,In_1052,In_1665);
nor U992 (N_992,In_173,In_969);
nand U993 (N_993,In_228,In_669);
nor U994 (N_994,In_329,In_600);
or U995 (N_995,In_622,In_901);
nand U996 (N_996,In_381,In_39);
xor U997 (N_997,In_2441,In_144);
and U998 (N_998,In_746,In_2017);
or U999 (N_999,In_30,In_1016);
or U1000 (N_1000,In_1617,In_1894);
xor U1001 (N_1001,In_53,In_1750);
or U1002 (N_1002,In_219,In_826);
or U1003 (N_1003,In_1276,In_2145);
and U1004 (N_1004,In_2136,In_1718);
nor U1005 (N_1005,In_505,In_909);
or U1006 (N_1006,In_563,In_463);
or U1007 (N_1007,In_2352,In_1040);
or U1008 (N_1008,In_2465,In_847);
xor U1009 (N_1009,In_972,In_2476);
nor U1010 (N_1010,In_846,In_1771);
nor U1011 (N_1011,In_2438,In_833);
xor U1012 (N_1012,In_1443,In_834);
xnor U1013 (N_1013,In_110,In_200);
or U1014 (N_1014,In_1730,In_151);
xor U1015 (N_1015,In_604,In_714);
nand U1016 (N_1016,In_2155,In_1211);
xnor U1017 (N_1017,In_392,In_252);
nand U1018 (N_1018,In_376,In_1673);
and U1019 (N_1019,In_2382,In_921);
nor U1020 (N_1020,In_2479,In_1);
nand U1021 (N_1021,In_1826,In_1229);
nand U1022 (N_1022,In_282,In_2168);
nor U1023 (N_1023,In_888,In_730);
or U1024 (N_1024,In_1720,In_2445);
or U1025 (N_1025,In_975,In_733);
nand U1026 (N_1026,In_1056,In_2243);
nand U1027 (N_1027,In_1362,In_870);
xor U1028 (N_1028,In_1746,In_1184);
and U1029 (N_1029,In_1670,In_2320);
xnor U1030 (N_1030,In_11,In_1683);
and U1031 (N_1031,In_162,In_963);
and U1032 (N_1032,In_2026,In_1187);
nor U1033 (N_1033,In_251,In_235);
or U1034 (N_1034,In_770,In_262);
xnor U1035 (N_1035,In_913,In_2226);
nor U1036 (N_1036,In_2406,In_917);
xor U1037 (N_1037,In_2024,In_908);
nand U1038 (N_1038,In_1736,In_2197);
xor U1039 (N_1039,In_350,In_1898);
and U1040 (N_1040,In_1684,In_1884);
nor U1041 (N_1041,In_1280,In_172);
or U1042 (N_1042,In_2132,In_991);
and U1043 (N_1043,In_1569,In_1554);
nor U1044 (N_1044,In_2458,In_2422);
or U1045 (N_1045,In_2496,In_2056);
nor U1046 (N_1046,In_1845,In_718);
or U1047 (N_1047,In_575,In_539);
or U1048 (N_1048,In_710,In_1180);
and U1049 (N_1049,In_2002,In_2044);
nand U1050 (N_1050,In_165,In_193);
nand U1051 (N_1051,In_69,In_119);
and U1052 (N_1052,In_432,In_2468);
xor U1053 (N_1053,In_986,In_1693);
nor U1054 (N_1054,In_1007,In_585);
or U1055 (N_1055,In_642,In_2306);
or U1056 (N_1056,In_1243,In_1487);
nor U1057 (N_1057,In_97,In_633);
nor U1058 (N_1058,In_753,In_2319);
nand U1059 (N_1059,In_183,In_1523);
xor U1060 (N_1060,In_237,In_1157);
nor U1061 (N_1061,In_54,In_367);
nand U1062 (N_1062,In_776,In_559);
or U1063 (N_1063,In_1129,In_65);
nand U1064 (N_1064,In_985,In_1581);
nand U1065 (N_1065,In_1158,In_1188);
nand U1066 (N_1066,In_2464,In_735);
nor U1067 (N_1067,In_1244,In_440);
nand U1068 (N_1068,In_1968,In_9);
xnor U1069 (N_1069,In_2488,In_149);
xnor U1070 (N_1070,In_387,In_1888);
nor U1071 (N_1071,In_540,In_441);
nor U1072 (N_1072,In_978,In_916);
xnor U1073 (N_1073,In_691,In_1118);
xor U1074 (N_1074,In_1189,In_1786);
and U1075 (N_1075,In_1454,In_1602);
nand U1076 (N_1076,In_1389,In_1386);
and U1077 (N_1077,In_1332,In_464);
nor U1078 (N_1078,In_872,In_1320);
nor U1079 (N_1079,In_87,In_2205);
and U1080 (N_1080,In_926,In_254);
or U1081 (N_1081,In_495,In_448);
nand U1082 (N_1082,In_1001,In_531);
nor U1083 (N_1083,In_2484,In_1914);
nand U1084 (N_1084,In_240,In_884);
xor U1085 (N_1085,In_936,In_1835);
nand U1086 (N_1086,In_1464,In_1222);
xor U1087 (N_1087,In_250,In_266);
nor U1088 (N_1088,In_1949,In_524);
and U1089 (N_1089,In_1017,In_1760);
nor U1090 (N_1090,In_2139,In_573);
nor U1091 (N_1091,In_1200,In_1239);
nand U1092 (N_1092,In_1675,In_900);
or U1093 (N_1093,In_1094,In_845);
xor U1094 (N_1094,In_1743,In_1130);
or U1095 (N_1095,In_1493,In_2245);
and U1096 (N_1096,In_34,In_976);
and U1097 (N_1097,In_1933,In_2400);
nand U1098 (N_1098,In_2437,In_1600);
or U1099 (N_1099,In_2218,In_1627);
nand U1100 (N_1100,In_103,In_971);
nor U1101 (N_1101,In_298,In_1359);
xor U1102 (N_1102,In_1879,In_10);
and U1103 (N_1103,In_1316,In_256);
and U1104 (N_1104,In_782,In_59);
and U1105 (N_1105,In_2109,In_1088);
or U1106 (N_1106,In_961,In_1154);
xor U1107 (N_1107,In_1824,In_1137);
nand U1108 (N_1108,In_48,In_203);
or U1109 (N_1109,In_1318,In_2234);
or U1110 (N_1110,In_694,In_1298);
xor U1111 (N_1111,In_2179,In_2202);
and U1112 (N_1112,In_2258,In_201);
or U1113 (N_1113,In_2454,In_1945);
or U1114 (N_1114,In_715,In_471);
nand U1115 (N_1115,In_2194,In_1807);
xor U1116 (N_1116,In_2272,In_1009);
xor U1117 (N_1117,In_1505,In_1423);
or U1118 (N_1118,In_1535,In_451);
xnor U1119 (N_1119,In_148,In_354);
or U1120 (N_1120,In_818,In_953);
or U1121 (N_1121,In_47,In_2257);
nor U1122 (N_1122,In_1164,In_1308);
and U1123 (N_1123,In_77,In_2379);
or U1124 (N_1124,In_835,In_1053);
and U1125 (N_1125,In_608,In_319);
or U1126 (N_1126,In_1125,In_2345);
and U1127 (N_1127,In_315,In_318);
nor U1128 (N_1128,In_1433,In_1358);
xnor U1129 (N_1129,In_1562,In_2420);
or U1130 (N_1130,In_2198,In_2068);
or U1131 (N_1131,In_1429,In_837);
and U1132 (N_1132,In_2398,In_1755);
nor U1133 (N_1133,In_422,In_1966);
and U1134 (N_1134,In_457,In_780);
and U1135 (N_1135,In_1714,In_289);
and U1136 (N_1136,In_1865,In_748);
and U1137 (N_1137,In_1995,In_2010);
and U1138 (N_1138,In_1912,In_624);
and U1139 (N_1139,In_91,In_1206);
nor U1140 (N_1140,In_2299,In_2451);
xor U1141 (N_1141,In_2120,In_1752);
nand U1142 (N_1142,In_1584,In_1756);
xor U1143 (N_1143,In_1370,In_2143);
nand U1144 (N_1144,In_2094,In_184);
nand U1145 (N_1145,In_1685,In_76);
nor U1146 (N_1146,In_1762,In_372);
and U1147 (N_1147,In_1419,In_1291);
xnor U1148 (N_1148,In_1336,In_1722);
nor U1149 (N_1149,In_652,In_2300);
and U1150 (N_1150,In_1601,In_948);
or U1151 (N_1151,In_1384,In_1387);
xnor U1152 (N_1152,In_794,In_284);
or U1153 (N_1153,In_497,In_1640);
nor U1154 (N_1154,In_1331,In_858);
and U1155 (N_1155,In_1941,In_2104);
xnor U1156 (N_1156,In_435,In_1170);
xnor U1157 (N_1157,In_997,In_577);
or U1158 (N_1158,In_1259,In_1434);
nor U1159 (N_1159,In_2426,In_862);
xor U1160 (N_1160,In_411,In_1202);
and U1161 (N_1161,In_2447,In_1520);
or U1162 (N_1162,In_135,In_215);
and U1163 (N_1163,In_428,In_1630);
xnor U1164 (N_1164,In_1134,In_795);
or U1165 (N_1165,In_2047,In_924);
or U1166 (N_1166,In_2004,In_1830);
or U1167 (N_1167,In_1289,In_1744);
nand U1168 (N_1168,In_472,In_2232);
xnor U1169 (N_1169,In_729,In_1218);
nor U1170 (N_1170,In_1340,In_2224);
xor U1171 (N_1171,In_1934,In_555);
xnor U1172 (N_1172,In_1608,In_86);
nand U1173 (N_1173,In_687,In_849);
and U1174 (N_1174,In_339,In_2499);
or U1175 (N_1175,In_1795,In_1224);
xnor U1176 (N_1176,In_1363,In_278);
nand U1177 (N_1177,In_2397,In_769);
nor U1178 (N_1178,In_1696,In_1538);
nor U1179 (N_1179,In_2264,In_1728);
nand U1180 (N_1180,In_423,In_297);
xor U1181 (N_1181,In_840,In_850);
or U1182 (N_1182,In_2086,In_736);
nor U1183 (N_1183,In_1124,In_2492);
xor U1184 (N_1184,In_492,In_1767);
xor U1185 (N_1185,In_1032,In_2361);
and U1186 (N_1186,In_2486,In_1033);
or U1187 (N_1187,In_541,In_932);
nor U1188 (N_1188,In_689,In_1445);
and U1189 (N_1189,In_761,In_895);
or U1190 (N_1190,In_35,In_1330);
nor U1191 (N_1191,In_1174,In_131);
nor U1192 (N_1192,In_937,In_1984);
xnor U1193 (N_1193,In_38,In_1208);
or U1194 (N_1194,In_2049,In_1064);
and U1195 (N_1195,In_2269,In_501);
or U1196 (N_1196,In_1282,In_31);
nor U1197 (N_1197,In_810,In_509);
or U1198 (N_1198,In_1895,In_1765);
xnor U1199 (N_1199,In_1977,In_2375);
xor U1200 (N_1200,In_305,In_697);
nand U1201 (N_1201,In_439,In_799);
and U1202 (N_1202,In_655,In_1036);
nor U1203 (N_1203,In_1027,In_699);
nand U1204 (N_1204,In_2327,In_2335);
nand U1205 (N_1205,In_1635,In_1607);
nor U1206 (N_1206,In_258,In_290);
nand U1207 (N_1207,In_690,In_107);
and U1208 (N_1208,In_1729,In_676);
nand U1209 (N_1209,In_831,In_1552);
and U1210 (N_1210,In_819,In_384);
or U1211 (N_1211,In_115,In_24);
nor U1212 (N_1212,In_781,In_1631);
xor U1213 (N_1213,In_1619,In_594);
or U1214 (N_1214,In_1346,In_134);
nand U1215 (N_1215,In_1963,In_1437);
xnor U1216 (N_1216,In_1574,In_1962);
or U1217 (N_1217,In_211,In_277);
nor U1218 (N_1218,In_1940,In_1095);
nor U1219 (N_1219,In_1639,In_1078);
nand U1220 (N_1220,In_717,In_1872);
nand U1221 (N_1221,In_2354,In_1859);
and U1222 (N_1222,In_2274,In_955);
xor U1223 (N_1223,In_1393,In_2330);
xnor U1224 (N_1224,In_396,In_1010);
xnor U1225 (N_1225,In_101,In_919);
nor U1226 (N_1226,In_527,In_2233);
nand U1227 (N_1227,In_693,In_2290);
xnor U1228 (N_1228,In_498,In_2156);
and U1229 (N_1229,In_1999,In_906);
or U1230 (N_1230,In_2241,In_1519);
nand U1231 (N_1231,In_1672,In_2372);
nand U1232 (N_1232,In_1837,In_1676);
xor U1233 (N_1233,In_295,In_1565);
or U1234 (N_1234,In_1122,In_606);
nand U1235 (N_1235,In_2121,In_2248);
and U1236 (N_1236,In_1668,In_705);
or U1237 (N_1237,In_1615,In_26);
or U1238 (N_1238,In_488,In_1789);
and U1239 (N_1239,In_1471,In_1658);
xnor U1240 (N_1240,In_317,In_1261);
nor U1241 (N_1241,In_2023,In_176);
nand U1242 (N_1242,In_2160,In_1104);
nor U1243 (N_1243,In_2276,In_867);
nand U1244 (N_1244,In_665,In_1151);
or U1245 (N_1245,In_1198,In_956);
nand U1246 (N_1246,In_2052,In_2480);
and U1247 (N_1247,In_1219,In_1573);
nor U1248 (N_1248,In_2251,In_1841);
or U1249 (N_1249,In_1105,In_2223);
and U1250 (N_1250,In_1123,In_1965);
nor U1251 (N_1251,In_836,In_504);
or U1252 (N_1252,In_1765,In_145);
nand U1253 (N_1253,In_1979,In_890);
or U1254 (N_1254,In_1222,In_1774);
or U1255 (N_1255,In_1023,In_2140);
nand U1256 (N_1256,In_523,In_1642);
xor U1257 (N_1257,In_667,In_528);
or U1258 (N_1258,In_1638,In_731);
and U1259 (N_1259,In_110,In_1593);
and U1260 (N_1260,In_736,In_730);
or U1261 (N_1261,In_810,In_1090);
nand U1262 (N_1262,In_1238,In_2195);
and U1263 (N_1263,In_824,In_2244);
and U1264 (N_1264,In_2293,In_2023);
nand U1265 (N_1265,In_1909,In_1874);
nand U1266 (N_1266,In_583,In_220);
nand U1267 (N_1267,In_1503,In_1641);
nor U1268 (N_1268,In_1509,In_647);
or U1269 (N_1269,In_1119,In_2490);
nand U1270 (N_1270,In_860,In_1321);
nor U1271 (N_1271,In_353,In_1601);
or U1272 (N_1272,In_1291,In_2280);
xnor U1273 (N_1273,In_829,In_2440);
or U1274 (N_1274,In_813,In_871);
or U1275 (N_1275,In_2157,In_1174);
nor U1276 (N_1276,In_732,In_1856);
xor U1277 (N_1277,In_713,In_2293);
nor U1278 (N_1278,In_937,In_2009);
xor U1279 (N_1279,In_1198,In_820);
xnor U1280 (N_1280,In_555,In_487);
nand U1281 (N_1281,In_2288,In_1859);
nand U1282 (N_1282,In_1813,In_2110);
or U1283 (N_1283,In_419,In_1676);
nor U1284 (N_1284,In_2191,In_298);
or U1285 (N_1285,In_1849,In_534);
nor U1286 (N_1286,In_2063,In_2402);
or U1287 (N_1287,In_919,In_2337);
nand U1288 (N_1288,In_2486,In_1985);
nand U1289 (N_1289,In_156,In_1168);
or U1290 (N_1290,In_1732,In_343);
xnor U1291 (N_1291,In_1148,In_1958);
xor U1292 (N_1292,In_2028,In_1030);
nand U1293 (N_1293,In_1642,In_773);
nand U1294 (N_1294,In_939,In_1577);
or U1295 (N_1295,In_1128,In_2363);
nor U1296 (N_1296,In_562,In_2236);
xor U1297 (N_1297,In_1736,In_182);
nor U1298 (N_1298,In_566,In_449);
and U1299 (N_1299,In_609,In_704);
xnor U1300 (N_1300,In_1784,In_2192);
xor U1301 (N_1301,In_2196,In_1542);
or U1302 (N_1302,In_2460,In_606);
xor U1303 (N_1303,In_496,In_1971);
nor U1304 (N_1304,In_53,In_987);
nor U1305 (N_1305,In_1121,In_2011);
xnor U1306 (N_1306,In_2115,In_136);
nand U1307 (N_1307,In_2085,In_2431);
and U1308 (N_1308,In_1547,In_1917);
nand U1309 (N_1309,In_1241,In_1941);
and U1310 (N_1310,In_2002,In_2152);
or U1311 (N_1311,In_15,In_2367);
nand U1312 (N_1312,In_1255,In_130);
nor U1313 (N_1313,In_983,In_532);
nand U1314 (N_1314,In_211,In_968);
nor U1315 (N_1315,In_1164,In_1066);
xor U1316 (N_1316,In_2111,In_1974);
xnor U1317 (N_1317,In_1938,In_169);
nand U1318 (N_1318,In_2081,In_1725);
nand U1319 (N_1319,In_2126,In_2371);
xnor U1320 (N_1320,In_220,In_2302);
or U1321 (N_1321,In_1158,In_1589);
nor U1322 (N_1322,In_888,In_1133);
nand U1323 (N_1323,In_1647,In_1563);
or U1324 (N_1324,In_51,In_139);
nand U1325 (N_1325,In_1181,In_1292);
nand U1326 (N_1326,In_1631,In_11);
xor U1327 (N_1327,In_255,In_477);
or U1328 (N_1328,In_361,In_897);
and U1329 (N_1329,In_1696,In_411);
or U1330 (N_1330,In_2033,In_878);
xnor U1331 (N_1331,In_1185,In_1763);
nand U1332 (N_1332,In_1934,In_1401);
xor U1333 (N_1333,In_1784,In_256);
xor U1334 (N_1334,In_503,In_1961);
and U1335 (N_1335,In_2220,In_688);
nand U1336 (N_1336,In_1424,In_1734);
nand U1337 (N_1337,In_1479,In_2339);
nor U1338 (N_1338,In_255,In_1977);
xor U1339 (N_1339,In_696,In_917);
and U1340 (N_1340,In_1838,In_1141);
xnor U1341 (N_1341,In_2388,In_1865);
nor U1342 (N_1342,In_1853,In_14);
or U1343 (N_1343,In_1756,In_604);
and U1344 (N_1344,In_1221,In_1147);
or U1345 (N_1345,In_1813,In_2324);
and U1346 (N_1346,In_1023,In_2303);
or U1347 (N_1347,In_1042,In_2123);
xnor U1348 (N_1348,In_570,In_1300);
nand U1349 (N_1349,In_365,In_1687);
nand U1350 (N_1350,In_1109,In_1517);
and U1351 (N_1351,In_1881,In_34);
or U1352 (N_1352,In_440,In_1778);
nor U1353 (N_1353,In_1958,In_53);
nand U1354 (N_1354,In_2463,In_84);
and U1355 (N_1355,In_591,In_2489);
or U1356 (N_1356,In_1574,In_1649);
nand U1357 (N_1357,In_449,In_1901);
and U1358 (N_1358,In_2281,In_275);
nand U1359 (N_1359,In_2075,In_266);
or U1360 (N_1360,In_1653,In_1487);
or U1361 (N_1361,In_151,In_2125);
and U1362 (N_1362,In_1385,In_82);
or U1363 (N_1363,In_938,In_1435);
nor U1364 (N_1364,In_431,In_2447);
xor U1365 (N_1365,In_2360,In_1564);
nor U1366 (N_1366,In_917,In_1447);
nand U1367 (N_1367,In_983,In_282);
or U1368 (N_1368,In_1437,In_1770);
xnor U1369 (N_1369,In_2140,In_2481);
nand U1370 (N_1370,In_990,In_2233);
nor U1371 (N_1371,In_2320,In_1055);
nand U1372 (N_1372,In_202,In_2397);
and U1373 (N_1373,In_2220,In_1123);
xor U1374 (N_1374,In_636,In_452);
and U1375 (N_1375,In_95,In_2214);
nand U1376 (N_1376,In_300,In_113);
and U1377 (N_1377,In_702,In_2122);
and U1378 (N_1378,In_2347,In_302);
or U1379 (N_1379,In_1371,In_1317);
nand U1380 (N_1380,In_1169,In_1644);
xor U1381 (N_1381,In_256,In_503);
nand U1382 (N_1382,In_2258,In_1550);
nand U1383 (N_1383,In_1839,In_430);
and U1384 (N_1384,In_221,In_1175);
xnor U1385 (N_1385,In_2003,In_814);
and U1386 (N_1386,In_928,In_1745);
nor U1387 (N_1387,In_942,In_1582);
or U1388 (N_1388,In_2040,In_2212);
nor U1389 (N_1389,In_1580,In_2165);
nand U1390 (N_1390,In_2118,In_286);
nand U1391 (N_1391,In_450,In_700);
nand U1392 (N_1392,In_362,In_2208);
and U1393 (N_1393,In_2286,In_1616);
xnor U1394 (N_1394,In_1535,In_52);
nor U1395 (N_1395,In_918,In_1297);
xor U1396 (N_1396,In_813,In_983);
xnor U1397 (N_1397,In_1111,In_49);
or U1398 (N_1398,In_1658,In_45);
or U1399 (N_1399,In_1067,In_2175);
xor U1400 (N_1400,In_1987,In_191);
xnor U1401 (N_1401,In_835,In_2237);
xor U1402 (N_1402,In_1631,In_1442);
and U1403 (N_1403,In_1409,In_1899);
nand U1404 (N_1404,In_908,In_2448);
or U1405 (N_1405,In_2199,In_632);
or U1406 (N_1406,In_754,In_5);
and U1407 (N_1407,In_735,In_846);
xor U1408 (N_1408,In_1434,In_942);
nor U1409 (N_1409,In_2274,In_578);
and U1410 (N_1410,In_1844,In_472);
nand U1411 (N_1411,In_241,In_679);
nand U1412 (N_1412,In_23,In_619);
xor U1413 (N_1413,In_1166,In_1556);
xnor U1414 (N_1414,In_379,In_2480);
nand U1415 (N_1415,In_1216,In_1498);
nor U1416 (N_1416,In_2106,In_474);
or U1417 (N_1417,In_1602,In_591);
nand U1418 (N_1418,In_129,In_1800);
and U1419 (N_1419,In_1980,In_1915);
nor U1420 (N_1420,In_629,In_1885);
and U1421 (N_1421,In_318,In_594);
nor U1422 (N_1422,In_2122,In_111);
xnor U1423 (N_1423,In_635,In_2476);
nor U1424 (N_1424,In_509,In_1939);
or U1425 (N_1425,In_2069,In_2155);
xnor U1426 (N_1426,In_2471,In_411);
and U1427 (N_1427,In_910,In_351);
nand U1428 (N_1428,In_235,In_496);
and U1429 (N_1429,In_1506,In_1838);
or U1430 (N_1430,In_1037,In_1277);
nand U1431 (N_1431,In_1716,In_2046);
or U1432 (N_1432,In_406,In_1217);
xnor U1433 (N_1433,In_2404,In_1806);
xor U1434 (N_1434,In_66,In_2328);
nor U1435 (N_1435,In_316,In_2171);
xnor U1436 (N_1436,In_409,In_688);
or U1437 (N_1437,In_1304,In_2432);
nand U1438 (N_1438,In_979,In_1147);
nor U1439 (N_1439,In_1457,In_1128);
and U1440 (N_1440,In_403,In_1797);
or U1441 (N_1441,In_1088,In_651);
nor U1442 (N_1442,In_147,In_190);
or U1443 (N_1443,In_1979,In_2048);
nand U1444 (N_1444,In_519,In_1603);
or U1445 (N_1445,In_2092,In_320);
nor U1446 (N_1446,In_217,In_485);
nand U1447 (N_1447,In_458,In_1434);
and U1448 (N_1448,In_1460,In_969);
nand U1449 (N_1449,In_1116,In_2021);
or U1450 (N_1450,In_408,In_769);
and U1451 (N_1451,In_1297,In_811);
or U1452 (N_1452,In_2154,In_315);
nand U1453 (N_1453,In_209,In_2133);
or U1454 (N_1454,In_1329,In_1738);
nor U1455 (N_1455,In_2495,In_2487);
and U1456 (N_1456,In_359,In_2165);
and U1457 (N_1457,In_865,In_2374);
nand U1458 (N_1458,In_329,In_2491);
nor U1459 (N_1459,In_1663,In_43);
nand U1460 (N_1460,In_1313,In_995);
nand U1461 (N_1461,In_840,In_1393);
xnor U1462 (N_1462,In_257,In_2160);
or U1463 (N_1463,In_771,In_1313);
nor U1464 (N_1464,In_2142,In_746);
xor U1465 (N_1465,In_1807,In_1836);
nor U1466 (N_1466,In_1950,In_867);
nor U1467 (N_1467,In_976,In_630);
xnor U1468 (N_1468,In_1033,In_1635);
nor U1469 (N_1469,In_1857,In_1695);
nor U1470 (N_1470,In_1883,In_952);
and U1471 (N_1471,In_515,In_351);
xnor U1472 (N_1472,In_1793,In_233);
and U1473 (N_1473,In_2392,In_2404);
or U1474 (N_1474,In_361,In_786);
or U1475 (N_1475,In_475,In_604);
and U1476 (N_1476,In_1314,In_256);
nor U1477 (N_1477,In_1122,In_2095);
or U1478 (N_1478,In_1261,In_328);
or U1479 (N_1479,In_2167,In_2370);
and U1480 (N_1480,In_2275,In_359);
or U1481 (N_1481,In_746,In_997);
nand U1482 (N_1482,In_2313,In_1957);
nor U1483 (N_1483,In_863,In_952);
or U1484 (N_1484,In_1448,In_626);
nor U1485 (N_1485,In_1957,In_1090);
or U1486 (N_1486,In_1668,In_2367);
and U1487 (N_1487,In_1957,In_157);
nand U1488 (N_1488,In_899,In_2182);
nand U1489 (N_1489,In_832,In_1005);
and U1490 (N_1490,In_662,In_1312);
or U1491 (N_1491,In_1848,In_1425);
xnor U1492 (N_1492,In_940,In_2474);
and U1493 (N_1493,In_712,In_826);
or U1494 (N_1494,In_1768,In_47);
xor U1495 (N_1495,In_1512,In_10);
nand U1496 (N_1496,In_650,In_1557);
nor U1497 (N_1497,In_865,In_1057);
and U1498 (N_1498,In_606,In_957);
nand U1499 (N_1499,In_538,In_510);
or U1500 (N_1500,In_484,In_1785);
and U1501 (N_1501,In_230,In_934);
and U1502 (N_1502,In_205,In_1522);
or U1503 (N_1503,In_1449,In_2405);
nor U1504 (N_1504,In_2166,In_12);
or U1505 (N_1505,In_2107,In_2222);
nand U1506 (N_1506,In_2269,In_2241);
or U1507 (N_1507,In_1648,In_854);
or U1508 (N_1508,In_2045,In_1696);
nor U1509 (N_1509,In_556,In_1038);
nand U1510 (N_1510,In_1676,In_726);
nor U1511 (N_1511,In_1295,In_1407);
xnor U1512 (N_1512,In_219,In_598);
nor U1513 (N_1513,In_1061,In_90);
xnor U1514 (N_1514,In_1776,In_2313);
nor U1515 (N_1515,In_1424,In_429);
nand U1516 (N_1516,In_1096,In_1372);
xnor U1517 (N_1517,In_1343,In_1163);
xor U1518 (N_1518,In_367,In_1937);
nand U1519 (N_1519,In_2318,In_1132);
nand U1520 (N_1520,In_2468,In_2419);
nor U1521 (N_1521,In_1407,In_469);
and U1522 (N_1522,In_2372,In_2009);
and U1523 (N_1523,In_1487,In_1443);
nand U1524 (N_1524,In_1348,In_2244);
xor U1525 (N_1525,In_2267,In_2487);
nand U1526 (N_1526,In_704,In_1283);
xor U1527 (N_1527,In_709,In_2317);
and U1528 (N_1528,In_1013,In_2294);
nand U1529 (N_1529,In_1218,In_1331);
or U1530 (N_1530,In_2466,In_1266);
nand U1531 (N_1531,In_1113,In_830);
nand U1532 (N_1532,In_750,In_2206);
nand U1533 (N_1533,In_2071,In_2219);
xor U1534 (N_1534,In_1131,In_1963);
nor U1535 (N_1535,In_1685,In_104);
and U1536 (N_1536,In_2472,In_801);
or U1537 (N_1537,In_556,In_533);
or U1538 (N_1538,In_2308,In_60);
or U1539 (N_1539,In_1223,In_416);
and U1540 (N_1540,In_235,In_1644);
and U1541 (N_1541,In_2255,In_631);
and U1542 (N_1542,In_658,In_713);
nand U1543 (N_1543,In_1511,In_1142);
and U1544 (N_1544,In_1222,In_836);
or U1545 (N_1545,In_1388,In_1953);
xnor U1546 (N_1546,In_2197,In_1516);
nor U1547 (N_1547,In_1980,In_1227);
nor U1548 (N_1548,In_482,In_1018);
nand U1549 (N_1549,In_2349,In_1988);
xnor U1550 (N_1550,In_1875,In_1445);
nand U1551 (N_1551,In_1412,In_132);
nor U1552 (N_1552,In_813,In_1407);
or U1553 (N_1553,In_1265,In_1126);
and U1554 (N_1554,In_776,In_598);
and U1555 (N_1555,In_1062,In_1077);
and U1556 (N_1556,In_1113,In_1776);
or U1557 (N_1557,In_2442,In_1780);
and U1558 (N_1558,In_1998,In_692);
or U1559 (N_1559,In_2458,In_380);
xnor U1560 (N_1560,In_2004,In_2108);
and U1561 (N_1561,In_1540,In_329);
or U1562 (N_1562,In_301,In_1752);
xor U1563 (N_1563,In_192,In_1919);
or U1564 (N_1564,In_1951,In_1138);
nor U1565 (N_1565,In_767,In_902);
nor U1566 (N_1566,In_1905,In_12);
or U1567 (N_1567,In_80,In_2080);
nand U1568 (N_1568,In_433,In_825);
nor U1569 (N_1569,In_452,In_547);
nor U1570 (N_1570,In_2422,In_2063);
xnor U1571 (N_1571,In_623,In_1396);
or U1572 (N_1572,In_1463,In_905);
nor U1573 (N_1573,In_928,In_1911);
xnor U1574 (N_1574,In_1319,In_2025);
or U1575 (N_1575,In_47,In_142);
or U1576 (N_1576,In_1142,In_809);
nor U1577 (N_1577,In_1338,In_867);
or U1578 (N_1578,In_2067,In_1231);
xnor U1579 (N_1579,In_1663,In_391);
nand U1580 (N_1580,In_2257,In_852);
nand U1581 (N_1581,In_1869,In_644);
and U1582 (N_1582,In_2281,In_1310);
or U1583 (N_1583,In_114,In_175);
xnor U1584 (N_1584,In_963,In_2358);
xor U1585 (N_1585,In_1977,In_566);
and U1586 (N_1586,In_2207,In_2030);
nand U1587 (N_1587,In_1460,In_149);
xnor U1588 (N_1588,In_2020,In_1478);
xor U1589 (N_1589,In_1804,In_1325);
nor U1590 (N_1590,In_2180,In_973);
and U1591 (N_1591,In_1174,In_733);
nor U1592 (N_1592,In_711,In_2031);
and U1593 (N_1593,In_1619,In_506);
nor U1594 (N_1594,In_206,In_1180);
and U1595 (N_1595,In_1904,In_1189);
or U1596 (N_1596,In_1238,In_1647);
nand U1597 (N_1597,In_1712,In_550);
or U1598 (N_1598,In_2405,In_1664);
and U1599 (N_1599,In_1009,In_2351);
or U1600 (N_1600,In_665,In_30);
nand U1601 (N_1601,In_1680,In_151);
nor U1602 (N_1602,In_237,In_1225);
nor U1603 (N_1603,In_581,In_833);
nand U1604 (N_1604,In_2364,In_1091);
xnor U1605 (N_1605,In_746,In_2203);
nand U1606 (N_1606,In_209,In_744);
xor U1607 (N_1607,In_671,In_1169);
nand U1608 (N_1608,In_2357,In_277);
and U1609 (N_1609,In_2320,In_1418);
xnor U1610 (N_1610,In_1186,In_920);
and U1611 (N_1611,In_2059,In_694);
nand U1612 (N_1612,In_1819,In_1312);
xnor U1613 (N_1613,In_956,In_1274);
nor U1614 (N_1614,In_1840,In_1875);
nand U1615 (N_1615,In_2250,In_650);
and U1616 (N_1616,In_410,In_797);
and U1617 (N_1617,In_1483,In_657);
nand U1618 (N_1618,In_189,In_1141);
nand U1619 (N_1619,In_1081,In_322);
and U1620 (N_1620,In_1362,In_809);
nor U1621 (N_1621,In_2306,In_2169);
nand U1622 (N_1622,In_692,In_616);
nand U1623 (N_1623,In_707,In_224);
nand U1624 (N_1624,In_2464,In_981);
xnor U1625 (N_1625,In_1630,In_2095);
nand U1626 (N_1626,In_1987,In_2211);
nand U1627 (N_1627,In_1394,In_283);
nor U1628 (N_1628,In_2143,In_106);
xor U1629 (N_1629,In_2069,In_2370);
nand U1630 (N_1630,In_1374,In_1275);
xnor U1631 (N_1631,In_298,In_90);
nor U1632 (N_1632,In_909,In_867);
and U1633 (N_1633,In_1342,In_1186);
nor U1634 (N_1634,In_922,In_1968);
nor U1635 (N_1635,In_2290,In_2204);
nand U1636 (N_1636,In_584,In_2008);
and U1637 (N_1637,In_2243,In_2373);
nand U1638 (N_1638,In_1144,In_567);
nand U1639 (N_1639,In_1907,In_1161);
or U1640 (N_1640,In_2419,In_1448);
nor U1641 (N_1641,In_2175,In_1937);
or U1642 (N_1642,In_1568,In_603);
or U1643 (N_1643,In_789,In_1986);
nor U1644 (N_1644,In_2469,In_2392);
and U1645 (N_1645,In_694,In_157);
and U1646 (N_1646,In_481,In_781);
xor U1647 (N_1647,In_1229,In_1626);
or U1648 (N_1648,In_2066,In_1702);
nand U1649 (N_1649,In_1908,In_129);
or U1650 (N_1650,In_2095,In_1678);
or U1651 (N_1651,In_2120,In_1386);
nand U1652 (N_1652,In_2158,In_2263);
and U1653 (N_1653,In_1562,In_36);
and U1654 (N_1654,In_1944,In_2254);
xor U1655 (N_1655,In_504,In_1245);
or U1656 (N_1656,In_729,In_1545);
and U1657 (N_1657,In_398,In_1385);
xnor U1658 (N_1658,In_1614,In_629);
nand U1659 (N_1659,In_1418,In_2136);
xnor U1660 (N_1660,In_39,In_2183);
xor U1661 (N_1661,In_321,In_911);
nor U1662 (N_1662,In_1719,In_1121);
and U1663 (N_1663,In_899,In_1681);
nand U1664 (N_1664,In_1249,In_810);
nor U1665 (N_1665,In_889,In_1139);
or U1666 (N_1666,In_1652,In_1901);
xor U1667 (N_1667,In_2117,In_401);
nand U1668 (N_1668,In_1850,In_11);
or U1669 (N_1669,In_368,In_1060);
or U1670 (N_1670,In_271,In_73);
or U1671 (N_1671,In_610,In_1201);
nand U1672 (N_1672,In_1114,In_1693);
nand U1673 (N_1673,In_2228,In_954);
and U1674 (N_1674,In_1986,In_88);
or U1675 (N_1675,In_2405,In_2311);
nand U1676 (N_1676,In_1384,In_1415);
and U1677 (N_1677,In_1932,In_2350);
or U1678 (N_1678,In_1959,In_1059);
xnor U1679 (N_1679,In_659,In_1102);
or U1680 (N_1680,In_1669,In_1315);
and U1681 (N_1681,In_1947,In_1531);
nor U1682 (N_1682,In_1567,In_1842);
nor U1683 (N_1683,In_763,In_1883);
xnor U1684 (N_1684,In_1623,In_1154);
xor U1685 (N_1685,In_267,In_471);
or U1686 (N_1686,In_588,In_2128);
or U1687 (N_1687,In_2047,In_1691);
or U1688 (N_1688,In_1520,In_1597);
xnor U1689 (N_1689,In_466,In_800);
or U1690 (N_1690,In_1876,In_742);
nand U1691 (N_1691,In_304,In_1589);
xnor U1692 (N_1692,In_1308,In_918);
or U1693 (N_1693,In_547,In_2329);
xnor U1694 (N_1694,In_944,In_593);
xor U1695 (N_1695,In_1316,In_360);
xor U1696 (N_1696,In_80,In_570);
nand U1697 (N_1697,In_1157,In_1219);
and U1698 (N_1698,In_1360,In_951);
and U1699 (N_1699,In_15,In_1063);
or U1700 (N_1700,In_1027,In_1792);
xor U1701 (N_1701,In_1830,In_212);
xnor U1702 (N_1702,In_1750,In_1512);
xnor U1703 (N_1703,In_1244,In_1586);
nor U1704 (N_1704,In_1740,In_2161);
xnor U1705 (N_1705,In_1882,In_1903);
xor U1706 (N_1706,In_488,In_1513);
xnor U1707 (N_1707,In_2036,In_2421);
nand U1708 (N_1708,In_1730,In_1403);
or U1709 (N_1709,In_2454,In_651);
or U1710 (N_1710,In_202,In_2152);
nand U1711 (N_1711,In_1787,In_2400);
nor U1712 (N_1712,In_2,In_1764);
and U1713 (N_1713,In_831,In_2178);
xor U1714 (N_1714,In_167,In_2354);
nor U1715 (N_1715,In_728,In_136);
nor U1716 (N_1716,In_347,In_1946);
or U1717 (N_1717,In_1442,In_426);
nand U1718 (N_1718,In_1529,In_1173);
or U1719 (N_1719,In_456,In_2339);
and U1720 (N_1720,In_2421,In_336);
nor U1721 (N_1721,In_1965,In_2074);
nor U1722 (N_1722,In_2468,In_371);
nor U1723 (N_1723,In_2383,In_1449);
and U1724 (N_1724,In_4,In_924);
nor U1725 (N_1725,In_1403,In_2059);
or U1726 (N_1726,In_243,In_970);
xor U1727 (N_1727,In_288,In_977);
nor U1728 (N_1728,In_919,In_2492);
nand U1729 (N_1729,In_2387,In_1578);
nand U1730 (N_1730,In_437,In_1600);
nor U1731 (N_1731,In_114,In_1824);
and U1732 (N_1732,In_2244,In_2495);
nand U1733 (N_1733,In_329,In_998);
and U1734 (N_1734,In_1322,In_856);
or U1735 (N_1735,In_2423,In_256);
nor U1736 (N_1736,In_571,In_1559);
nand U1737 (N_1737,In_1226,In_1746);
nor U1738 (N_1738,In_2122,In_2013);
nand U1739 (N_1739,In_1061,In_375);
or U1740 (N_1740,In_861,In_1444);
nor U1741 (N_1741,In_30,In_1279);
nand U1742 (N_1742,In_2494,In_2091);
nor U1743 (N_1743,In_635,In_1364);
nor U1744 (N_1744,In_2275,In_2112);
or U1745 (N_1745,In_646,In_221);
or U1746 (N_1746,In_1015,In_61);
xnor U1747 (N_1747,In_1555,In_1958);
and U1748 (N_1748,In_714,In_2230);
nor U1749 (N_1749,In_1680,In_2179);
and U1750 (N_1750,In_745,In_633);
nand U1751 (N_1751,In_56,In_436);
xor U1752 (N_1752,In_136,In_421);
and U1753 (N_1753,In_2001,In_1180);
xor U1754 (N_1754,In_731,In_411);
nor U1755 (N_1755,In_1231,In_22);
or U1756 (N_1756,In_2068,In_46);
nand U1757 (N_1757,In_2106,In_2098);
nand U1758 (N_1758,In_1348,In_1671);
nand U1759 (N_1759,In_713,In_1322);
and U1760 (N_1760,In_1536,In_1455);
and U1761 (N_1761,In_2296,In_1129);
nand U1762 (N_1762,In_1728,In_1131);
and U1763 (N_1763,In_1622,In_1808);
and U1764 (N_1764,In_1562,In_2010);
or U1765 (N_1765,In_1908,In_1761);
xnor U1766 (N_1766,In_1244,In_1150);
or U1767 (N_1767,In_737,In_2112);
nand U1768 (N_1768,In_233,In_2486);
nor U1769 (N_1769,In_488,In_319);
xnor U1770 (N_1770,In_1508,In_2349);
xnor U1771 (N_1771,In_819,In_1948);
or U1772 (N_1772,In_537,In_205);
nand U1773 (N_1773,In_697,In_1564);
or U1774 (N_1774,In_1151,In_1225);
xor U1775 (N_1775,In_1490,In_1827);
or U1776 (N_1776,In_1168,In_1677);
nand U1777 (N_1777,In_1269,In_2055);
nor U1778 (N_1778,In_471,In_887);
nor U1779 (N_1779,In_1002,In_522);
nand U1780 (N_1780,In_1970,In_2485);
and U1781 (N_1781,In_1977,In_1132);
xnor U1782 (N_1782,In_408,In_1505);
xor U1783 (N_1783,In_210,In_607);
or U1784 (N_1784,In_67,In_2189);
or U1785 (N_1785,In_972,In_1538);
nand U1786 (N_1786,In_683,In_1990);
or U1787 (N_1787,In_940,In_418);
xor U1788 (N_1788,In_1207,In_2328);
xnor U1789 (N_1789,In_1019,In_994);
or U1790 (N_1790,In_1656,In_703);
and U1791 (N_1791,In_753,In_2460);
nand U1792 (N_1792,In_959,In_738);
and U1793 (N_1793,In_1168,In_1645);
xor U1794 (N_1794,In_364,In_1516);
nor U1795 (N_1795,In_244,In_1665);
and U1796 (N_1796,In_2122,In_2499);
nand U1797 (N_1797,In_2020,In_163);
and U1798 (N_1798,In_362,In_519);
nand U1799 (N_1799,In_840,In_1299);
nand U1800 (N_1800,In_1899,In_2143);
nor U1801 (N_1801,In_1920,In_1040);
or U1802 (N_1802,In_1063,In_121);
xor U1803 (N_1803,In_1069,In_216);
or U1804 (N_1804,In_2132,In_2342);
and U1805 (N_1805,In_1581,In_1870);
or U1806 (N_1806,In_1788,In_1563);
nand U1807 (N_1807,In_508,In_2465);
nand U1808 (N_1808,In_116,In_2209);
xnor U1809 (N_1809,In_558,In_372);
and U1810 (N_1810,In_2362,In_582);
and U1811 (N_1811,In_1583,In_1414);
nor U1812 (N_1812,In_1382,In_761);
nand U1813 (N_1813,In_893,In_1869);
xor U1814 (N_1814,In_1829,In_912);
xor U1815 (N_1815,In_1877,In_1147);
and U1816 (N_1816,In_164,In_2335);
and U1817 (N_1817,In_2209,In_1837);
nor U1818 (N_1818,In_771,In_455);
and U1819 (N_1819,In_910,In_2321);
xnor U1820 (N_1820,In_426,In_1608);
or U1821 (N_1821,In_839,In_1770);
xor U1822 (N_1822,In_114,In_1175);
and U1823 (N_1823,In_598,In_1322);
nor U1824 (N_1824,In_144,In_91);
nor U1825 (N_1825,In_1716,In_1288);
or U1826 (N_1826,In_545,In_1511);
and U1827 (N_1827,In_626,In_120);
nor U1828 (N_1828,In_1592,In_1621);
nor U1829 (N_1829,In_471,In_811);
nor U1830 (N_1830,In_256,In_1285);
nand U1831 (N_1831,In_188,In_1972);
and U1832 (N_1832,In_225,In_1252);
nor U1833 (N_1833,In_1695,In_23);
nand U1834 (N_1834,In_529,In_2236);
and U1835 (N_1835,In_1908,In_1161);
nand U1836 (N_1836,In_1730,In_798);
nand U1837 (N_1837,In_2269,In_471);
nor U1838 (N_1838,In_54,In_224);
nor U1839 (N_1839,In_1856,In_1886);
and U1840 (N_1840,In_1925,In_864);
or U1841 (N_1841,In_1939,In_535);
and U1842 (N_1842,In_184,In_764);
nor U1843 (N_1843,In_304,In_2207);
and U1844 (N_1844,In_230,In_1990);
xnor U1845 (N_1845,In_1799,In_1901);
xnor U1846 (N_1846,In_341,In_2284);
or U1847 (N_1847,In_2300,In_2264);
nor U1848 (N_1848,In_1111,In_1736);
nand U1849 (N_1849,In_1826,In_2016);
nor U1850 (N_1850,In_2363,In_1234);
and U1851 (N_1851,In_101,In_938);
xor U1852 (N_1852,In_2206,In_2229);
nor U1853 (N_1853,In_1162,In_482);
and U1854 (N_1854,In_1,In_1970);
nand U1855 (N_1855,In_635,In_851);
and U1856 (N_1856,In_1830,In_513);
nor U1857 (N_1857,In_795,In_1946);
nand U1858 (N_1858,In_598,In_1304);
or U1859 (N_1859,In_327,In_1439);
nor U1860 (N_1860,In_199,In_1418);
nand U1861 (N_1861,In_2478,In_283);
xor U1862 (N_1862,In_287,In_1558);
and U1863 (N_1863,In_1873,In_1099);
nor U1864 (N_1864,In_2389,In_91);
xnor U1865 (N_1865,In_324,In_958);
xnor U1866 (N_1866,In_2152,In_402);
and U1867 (N_1867,In_2084,In_1820);
and U1868 (N_1868,In_2160,In_2374);
xnor U1869 (N_1869,In_834,In_2359);
xor U1870 (N_1870,In_2275,In_1884);
or U1871 (N_1871,In_1710,In_322);
xnor U1872 (N_1872,In_56,In_2035);
or U1873 (N_1873,In_1551,In_969);
xnor U1874 (N_1874,In_394,In_249);
or U1875 (N_1875,In_228,In_2033);
nor U1876 (N_1876,In_2137,In_1561);
nand U1877 (N_1877,In_1956,In_827);
nor U1878 (N_1878,In_2180,In_1165);
xor U1879 (N_1879,In_11,In_1182);
and U1880 (N_1880,In_134,In_1446);
and U1881 (N_1881,In_1818,In_265);
xor U1882 (N_1882,In_262,In_523);
nand U1883 (N_1883,In_1040,In_1019);
or U1884 (N_1884,In_2048,In_1076);
nand U1885 (N_1885,In_1917,In_2341);
and U1886 (N_1886,In_1234,In_1469);
nor U1887 (N_1887,In_647,In_2332);
xor U1888 (N_1888,In_1756,In_1399);
or U1889 (N_1889,In_1678,In_659);
nor U1890 (N_1890,In_1276,In_667);
nand U1891 (N_1891,In_851,In_426);
xnor U1892 (N_1892,In_180,In_985);
xor U1893 (N_1893,In_1323,In_2490);
or U1894 (N_1894,In_2373,In_388);
nand U1895 (N_1895,In_1652,In_245);
nor U1896 (N_1896,In_382,In_2230);
nor U1897 (N_1897,In_1936,In_441);
nor U1898 (N_1898,In_1306,In_2220);
nor U1899 (N_1899,In_2426,In_1674);
nor U1900 (N_1900,In_842,In_2495);
nor U1901 (N_1901,In_2411,In_1403);
and U1902 (N_1902,In_2061,In_385);
nand U1903 (N_1903,In_368,In_225);
or U1904 (N_1904,In_317,In_963);
nor U1905 (N_1905,In_2101,In_1963);
nor U1906 (N_1906,In_1677,In_1183);
xor U1907 (N_1907,In_2324,In_1104);
nand U1908 (N_1908,In_482,In_2288);
xnor U1909 (N_1909,In_935,In_784);
nand U1910 (N_1910,In_1902,In_288);
nor U1911 (N_1911,In_1308,In_296);
nand U1912 (N_1912,In_60,In_1060);
nor U1913 (N_1913,In_926,In_1385);
or U1914 (N_1914,In_2231,In_1325);
or U1915 (N_1915,In_2194,In_2332);
nand U1916 (N_1916,In_98,In_1233);
and U1917 (N_1917,In_1980,In_1689);
and U1918 (N_1918,In_2429,In_1485);
and U1919 (N_1919,In_1615,In_1360);
and U1920 (N_1920,In_2481,In_2209);
nand U1921 (N_1921,In_1160,In_1526);
and U1922 (N_1922,In_958,In_562);
or U1923 (N_1923,In_1998,In_2025);
or U1924 (N_1924,In_1845,In_2440);
xor U1925 (N_1925,In_2033,In_2445);
and U1926 (N_1926,In_1916,In_2247);
nor U1927 (N_1927,In_501,In_724);
nand U1928 (N_1928,In_1803,In_2260);
nor U1929 (N_1929,In_1869,In_2072);
nand U1930 (N_1930,In_1421,In_1543);
nor U1931 (N_1931,In_409,In_1340);
nand U1932 (N_1932,In_1720,In_959);
xnor U1933 (N_1933,In_1042,In_1062);
nand U1934 (N_1934,In_1678,In_1616);
and U1935 (N_1935,In_388,In_380);
and U1936 (N_1936,In_20,In_1853);
nor U1937 (N_1937,In_300,In_631);
and U1938 (N_1938,In_110,In_155);
nand U1939 (N_1939,In_1304,In_2376);
or U1940 (N_1940,In_376,In_1440);
nor U1941 (N_1941,In_1838,In_1724);
or U1942 (N_1942,In_2115,In_877);
nand U1943 (N_1943,In_2123,In_2267);
nor U1944 (N_1944,In_161,In_2343);
or U1945 (N_1945,In_1651,In_1226);
nand U1946 (N_1946,In_2389,In_1683);
nor U1947 (N_1947,In_1074,In_1481);
and U1948 (N_1948,In_682,In_1375);
or U1949 (N_1949,In_1186,In_2467);
xnor U1950 (N_1950,In_1869,In_2282);
and U1951 (N_1951,In_306,In_1815);
xnor U1952 (N_1952,In_1985,In_565);
nand U1953 (N_1953,In_2346,In_278);
xnor U1954 (N_1954,In_567,In_555);
or U1955 (N_1955,In_1846,In_1573);
xor U1956 (N_1956,In_1099,In_2076);
xnor U1957 (N_1957,In_948,In_646);
nand U1958 (N_1958,In_159,In_2031);
xnor U1959 (N_1959,In_966,In_56);
or U1960 (N_1960,In_142,In_1129);
nor U1961 (N_1961,In_144,In_1247);
xnor U1962 (N_1962,In_866,In_2014);
nor U1963 (N_1963,In_1836,In_1963);
or U1964 (N_1964,In_1272,In_2280);
or U1965 (N_1965,In_1390,In_1750);
nor U1966 (N_1966,In_1738,In_111);
xnor U1967 (N_1967,In_2381,In_492);
or U1968 (N_1968,In_1728,In_597);
and U1969 (N_1969,In_94,In_1827);
and U1970 (N_1970,In_1728,In_1403);
and U1971 (N_1971,In_1566,In_1792);
xor U1972 (N_1972,In_370,In_2133);
nor U1973 (N_1973,In_808,In_2072);
nor U1974 (N_1974,In_1147,In_744);
nand U1975 (N_1975,In_1300,In_385);
nor U1976 (N_1976,In_89,In_49);
or U1977 (N_1977,In_1621,In_2109);
xor U1978 (N_1978,In_1728,In_2310);
nor U1979 (N_1979,In_890,In_10);
or U1980 (N_1980,In_234,In_2012);
nand U1981 (N_1981,In_463,In_993);
nor U1982 (N_1982,In_244,In_1423);
and U1983 (N_1983,In_1477,In_773);
nor U1984 (N_1984,In_470,In_270);
nand U1985 (N_1985,In_65,In_662);
nor U1986 (N_1986,In_952,In_942);
nand U1987 (N_1987,In_1343,In_1395);
nor U1988 (N_1988,In_2274,In_1731);
or U1989 (N_1989,In_838,In_2396);
xnor U1990 (N_1990,In_348,In_1684);
xnor U1991 (N_1991,In_1672,In_1324);
nor U1992 (N_1992,In_1858,In_2104);
or U1993 (N_1993,In_229,In_1159);
and U1994 (N_1994,In_1764,In_1987);
nand U1995 (N_1995,In_1784,In_16);
xnor U1996 (N_1996,In_35,In_1160);
or U1997 (N_1997,In_630,In_1460);
nor U1998 (N_1998,In_1579,In_2414);
xnor U1999 (N_1999,In_1630,In_407);
xor U2000 (N_2000,In_389,In_656);
xnor U2001 (N_2001,In_1453,In_1792);
and U2002 (N_2002,In_931,In_313);
nor U2003 (N_2003,In_1083,In_767);
and U2004 (N_2004,In_713,In_950);
or U2005 (N_2005,In_477,In_1150);
nor U2006 (N_2006,In_1128,In_2362);
xnor U2007 (N_2007,In_1043,In_953);
nor U2008 (N_2008,In_48,In_1629);
nor U2009 (N_2009,In_294,In_181);
nor U2010 (N_2010,In_15,In_1274);
xor U2011 (N_2011,In_1423,In_1938);
nand U2012 (N_2012,In_1334,In_2012);
and U2013 (N_2013,In_1615,In_960);
xnor U2014 (N_2014,In_1701,In_160);
nor U2015 (N_2015,In_648,In_295);
or U2016 (N_2016,In_296,In_1065);
nand U2017 (N_2017,In_1450,In_2426);
nand U2018 (N_2018,In_2131,In_972);
xnor U2019 (N_2019,In_2163,In_855);
nand U2020 (N_2020,In_1094,In_280);
nand U2021 (N_2021,In_384,In_1136);
and U2022 (N_2022,In_2367,In_753);
and U2023 (N_2023,In_1954,In_1253);
or U2024 (N_2024,In_2413,In_313);
nand U2025 (N_2025,In_1030,In_1587);
or U2026 (N_2026,In_2098,In_290);
nor U2027 (N_2027,In_1325,In_224);
nand U2028 (N_2028,In_581,In_2343);
and U2029 (N_2029,In_2069,In_613);
and U2030 (N_2030,In_109,In_349);
nand U2031 (N_2031,In_1300,In_771);
and U2032 (N_2032,In_1072,In_869);
xor U2033 (N_2033,In_31,In_1197);
nor U2034 (N_2034,In_1803,In_387);
and U2035 (N_2035,In_1876,In_1559);
and U2036 (N_2036,In_1110,In_139);
or U2037 (N_2037,In_1545,In_1899);
and U2038 (N_2038,In_1215,In_1967);
or U2039 (N_2039,In_948,In_123);
xor U2040 (N_2040,In_2134,In_357);
or U2041 (N_2041,In_1160,In_251);
or U2042 (N_2042,In_1502,In_488);
nand U2043 (N_2043,In_2101,In_2390);
nor U2044 (N_2044,In_1693,In_1940);
nor U2045 (N_2045,In_1925,In_733);
nand U2046 (N_2046,In_1076,In_476);
nor U2047 (N_2047,In_918,In_391);
and U2048 (N_2048,In_1913,In_1145);
or U2049 (N_2049,In_165,In_213);
nand U2050 (N_2050,In_1838,In_50);
and U2051 (N_2051,In_347,In_1414);
or U2052 (N_2052,In_640,In_2341);
or U2053 (N_2053,In_2384,In_2253);
nor U2054 (N_2054,In_114,In_1302);
and U2055 (N_2055,In_2152,In_82);
nand U2056 (N_2056,In_694,In_1200);
or U2057 (N_2057,In_789,In_39);
nand U2058 (N_2058,In_2376,In_469);
and U2059 (N_2059,In_1882,In_150);
xnor U2060 (N_2060,In_1139,In_2227);
and U2061 (N_2061,In_1683,In_1198);
nor U2062 (N_2062,In_581,In_508);
xnor U2063 (N_2063,In_126,In_2237);
nor U2064 (N_2064,In_1693,In_1373);
or U2065 (N_2065,In_321,In_1592);
nand U2066 (N_2066,In_429,In_1853);
nor U2067 (N_2067,In_145,In_2441);
nand U2068 (N_2068,In_27,In_2152);
and U2069 (N_2069,In_2367,In_1066);
xor U2070 (N_2070,In_1097,In_1860);
nand U2071 (N_2071,In_150,In_1469);
and U2072 (N_2072,In_0,In_1152);
or U2073 (N_2073,In_2069,In_1993);
nor U2074 (N_2074,In_828,In_1040);
or U2075 (N_2075,In_822,In_483);
nand U2076 (N_2076,In_560,In_2472);
or U2077 (N_2077,In_2121,In_1115);
nor U2078 (N_2078,In_685,In_337);
or U2079 (N_2079,In_1624,In_1993);
and U2080 (N_2080,In_1292,In_24);
nor U2081 (N_2081,In_544,In_242);
xnor U2082 (N_2082,In_1233,In_683);
and U2083 (N_2083,In_574,In_2445);
nand U2084 (N_2084,In_1623,In_415);
nand U2085 (N_2085,In_2258,In_1378);
nand U2086 (N_2086,In_2431,In_946);
or U2087 (N_2087,In_606,In_2190);
nor U2088 (N_2088,In_2421,In_1662);
and U2089 (N_2089,In_544,In_290);
or U2090 (N_2090,In_3,In_325);
nor U2091 (N_2091,In_1355,In_68);
and U2092 (N_2092,In_740,In_73);
xor U2093 (N_2093,In_2057,In_1648);
xor U2094 (N_2094,In_130,In_649);
nand U2095 (N_2095,In_382,In_1716);
and U2096 (N_2096,In_1500,In_313);
xor U2097 (N_2097,In_284,In_185);
xnor U2098 (N_2098,In_1550,In_1544);
nor U2099 (N_2099,In_544,In_1345);
nor U2100 (N_2100,In_1323,In_27);
nor U2101 (N_2101,In_734,In_426);
and U2102 (N_2102,In_954,In_1853);
nor U2103 (N_2103,In_1681,In_1391);
and U2104 (N_2104,In_1295,In_954);
xor U2105 (N_2105,In_2474,In_1318);
or U2106 (N_2106,In_274,In_908);
and U2107 (N_2107,In_1404,In_655);
or U2108 (N_2108,In_0,In_1473);
nor U2109 (N_2109,In_1014,In_2144);
nor U2110 (N_2110,In_36,In_486);
nand U2111 (N_2111,In_243,In_1862);
or U2112 (N_2112,In_704,In_1725);
xor U2113 (N_2113,In_853,In_746);
and U2114 (N_2114,In_1678,In_1789);
and U2115 (N_2115,In_1332,In_106);
or U2116 (N_2116,In_1229,In_804);
or U2117 (N_2117,In_329,In_2449);
or U2118 (N_2118,In_1227,In_1194);
nand U2119 (N_2119,In_200,In_256);
or U2120 (N_2120,In_684,In_1418);
nor U2121 (N_2121,In_833,In_2157);
xnor U2122 (N_2122,In_1400,In_707);
xor U2123 (N_2123,In_630,In_1512);
or U2124 (N_2124,In_1353,In_1101);
nand U2125 (N_2125,In_787,In_1343);
xnor U2126 (N_2126,In_2382,In_2268);
xnor U2127 (N_2127,In_25,In_1072);
and U2128 (N_2128,In_1301,In_395);
nor U2129 (N_2129,In_987,In_66);
nor U2130 (N_2130,In_1444,In_1827);
nand U2131 (N_2131,In_586,In_1157);
nor U2132 (N_2132,In_854,In_637);
xnor U2133 (N_2133,In_2333,In_710);
nand U2134 (N_2134,In_1122,In_943);
and U2135 (N_2135,In_2224,In_1264);
xnor U2136 (N_2136,In_1041,In_719);
nand U2137 (N_2137,In_1959,In_602);
or U2138 (N_2138,In_343,In_937);
and U2139 (N_2139,In_489,In_2221);
nor U2140 (N_2140,In_125,In_908);
nor U2141 (N_2141,In_361,In_852);
or U2142 (N_2142,In_246,In_351);
xnor U2143 (N_2143,In_1811,In_1487);
or U2144 (N_2144,In_587,In_882);
xor U2145 (N_2145,In_1776,In_1893);
xnor U2146 (N_2146,In_2230,In_479);
and U2147 (N_2147,In_1929,In_2477);
nor U2148 (N_2148,In_786,In_985);
xnor U2149 (N_2149,In_493,In_2337);
xor U2150 (N_2150,In_1878,In_197);
xnor U2151 (N_2151,In_297,In_1830);
and U2152 (N_2152,In_1175,In_1004);
xor U2153 (N_2153,In_1901,In_667);
and U2154 (N_2154,In_1838,In_553);
and U2155 (N_2155,In_1873,In_2408);
nor U2156 (N_2156,In_1685,In_1972);
and U2157 (N_2157,In_1090,In_142);
nor U2158 (N_2158,In_187,In_295);
or U2159 (N_2159,In_357,In_1626);
or U2160 (N_2160,In_1031,In_721);
nor U2161 (N_2161,In_2309,In_508);
nor U2162 (N_2162,In_1378,In_1764);
xor U2163 (N_2163,In_1339,In_2474);
nor U2164 (N_2164,In_832,In_1534);
xor U2165 (N_2165,In_1673,In_2186);
nor U2166 (N_2166,In_2488,In_2396);
nor U2167 (N_2167,In_968,In_1385);
and U2168 (N_2168,In_1503,In_2360);
or U2169 (N_2169,In_1814,In_688);
nor U2170 (N_2170,In_1882,In_2267);
nor U2171 (N_2171,In_1665,In_1883);
nor U2172 (N_2172,In_2470,In_690);
or U2173 (N_2173,In_1641,In_965);
nand U2174 (N_2174,In_2401,In_2245);
and U2175 (N_2175,In_2147,In_926);
nand U2176 (N_2176,In_388,In_918);
nor U2177 (N_2177,In_1213,In_1931);
nor U2178 (N_2178,In_1708,In_7);
nand U2179 (N_2179,In_1165,In_601);
nand U2180 (N_2180,In_1496,In_2255);
xor U2181 (N_2181,In_2483,In_2129);
nor U2182 (N_2182,In_1359,In_1875);
xor U2183 (N_2183,In_322,In_1577);
nor U2184 (N_2184,In_1305,In_1382);
nand U2185 (N_2185,In_994,In_811);
nor U2186 (N_2186,In_1907,In_5);
xor U2187 (N_2187,In_866,In_888);
and U2188 (N_2188,In_723,In_608);
nor U2189 (N_2189,In_16,In_1381);
xnor U2190 (N_2190,In_589,In_1353);
nor U2191 (N_2191,In_1902,In_1565);
nand U2192 (N_2192,In_1420,In_1234);
nor U2193 (N_2193,In_373,In_859);
nor U2194 (N_2194,In_1794,In_1238);
nor U2195 (N_2195,In_171,In_2141);
nor U2196 (N_2196,In_398,In_1728);
nor U2197 (N_2197,In_2370,In_2468);
and U2198 (N_2198,In_2101,In_825);
nand U2199 (N_2199,In_1425,In_133);
or U2200 (N_2200,In_822,In_440);
and U2201 (N_2201,In_2256,In_1621);
and U2202 (N_2202,In_594,In_2043);
or U2203 (N_2203,In_32,In_287);
or U2204 (N_2204,In_591,In_1795);
nor U2205 (N_2205,In_103,In_87);
and U2206 (N_2206,In_2284,In_1397);
or U2207 (N_2207,In_1082,In_1378);
xor U2208 (N_2208,In_582,In_1759);
and U2209 (N_2209,In_2492,In_1538);
and U2210 (N_2210,In_589,In_2470);
or U2211 (N_2211,In_1104,In_1518);
xor U2212 (N_2212,In_2485,In_1502);
nor U2213 (N_2213,In_639,In_1690);
and U2214 (N_2214,In_537,In_325);
or U2215 (N_2215,In_2341,In_306);
nor U2216 (N_2216,In_1826,In_2224);
nor U2217 (N_2217,In_2216,In_1174);
nor U2218 (N_2218,In_2080,In_1565);
xnor U2219 (N_2219,In_643,In_1715);
xor U2220 (N_2220,In_1102,In_2071);
nand U2221 (N_2221,In_727,In_917);
nand U2222 (N_2222,In_207,In_482);
xnor U2223 (N_2223,In_914,In_42);
and U2224 (N_2224,In_597,In_1107);
nor U2225 (N_2225,In_817,In_750);
nand U2226 (N_2226,In_1698,In_538);
and U2227 (N_2227,In_523,In_2088);
and U2228 (N_2228,In_2172,In_1624);
nand U2229 (N_2229,In_2187,In_778);
nor U2230 (N_2230,In_1597,In_671);
or U2231 (N_2231,In_1555,In_989);
or U2232 (N_2232,In_2418,In_1052);
nand U2233 (N_2233,In_1081,In_159);
xor U2234 (N_2234,In_2263,In_271);
and U2235 (N_2235,In_687,In_1693);
or U2236 (N_2236,In_1161,In_46);
and U2237 (N_2237,In_314,In_2362);
xnor U2238 (N_2238,In_943,In_1086);
and U2239 (N_2239,In_2391,In_304);
nand U2240 (N_2240,In_422,In_1659);
xor U2241 (N_2241,In_2427,In_2170);
and U2242 (N_2242,In_914,In_537);
xnor U2243 (N_2243,In_208,In_420);
nor U2244 (N_2244,In_2182,In_1888);
xnor U2245 (N_2245,In_1224,In_1717);
nor U2246 (N_2246,In_1594,In_1779);
and U2247 (N_2247,In_1231,In_2325);
and U2248 (N_2248,In_799,In_788);
nand U2249 (N_2249,In_1261,In_1525);
or U2250 (N_2250,In_745,In_985);
nor U2251 (N_2251,In_1646,In_0);
xnor U2252 (N_2252,In_865,In_1177);
and U2253 (N_2253,In_2173,In_1913);
xor U2254 (N_2254,In_507,In_1019);
and U2255 (N_2255,In_111,In_2284);
and U2256 (N_2256,In_349,In_1870);
or U2257 (N_2257,In_2229,In_672);
nand U2258 (N_2258,In_2344,In_1271);
or U2259 (N_2259,In_896,In_2041);
and U2260 (N_2260,In_1824,In_784);
and U2261 (N_2261,In_2242,In_2209);
xnor U2262 (N_2262,In_780,In_1428);
nor U2263 (N_2263,In_2064,In_2441);
xor U2264 (N_2264,In_123,In_2054);
xnor U2265 (N_2265,In_739,In_1865);
xnor U2266 (N_2266,In_590,In_1980);
or U2267 (N_2267,In_2411,In_2222);
nor U2268 (N_2268,In_2306,In_1196);
nor U2269 (N_2269,In_1274,In_1494);
xor U2270 (N_2270,In_1045,In_38);
or U2271 (N_2271,In_651,In_1953);
or U2272 (N_2272,In_1448,In_2175);
or U2273 (N_2273,In_876,In_2000);
nand U2274 (N_2274,In_1789,In_1125);
xnor U2275 (N_2275,In_2111,In_2081);
nor U2276 (N_2276,In_410,In_1621);
and U2277 (N_2277,In_787,In_1313);
and U2278 (N_2278,In_234,In_2066);
and U2279 (N_2279,In_1211,In_763);
xor U2280 (N_2280,In_1793,In_1756);
or U2281 (N_2281,In_1503,In_916);
or U2282 (N_2282,In_1890,In_1355);
nand U2283 (N_2283,In_500,In_1568);
nand U2284 (N_2284,In_802,In_2104);
nand U2285 (N_2285,In_2018,In_1584);
nor U2286 (N_2286,In_1789,In_50);
nand U2287 (N_2287,In_595,In_1941);
nor U2288 (N_2288,In_1379,In_196);
or U2289 (N_2289,In_1221,In_1233);
nand U2290 (N_2290,In_1415,In_2415);
nand U2291 (N_2291,In_1239,In_981);
xor U2292 (N_2292,In_1989,In_1708);
nand U2293 (N_2293,In_1898,In_2261);
xnor U2294 (N_2294,In_1705,In_498);
or U2295 (N_2295,In_2239,In_707);
or U2296 (N_2296,In_608,In_1337);
nor U2297 (N_2297,In_10,In_1944);
and U2298 (N_2298,In_862,In_2075);
nand U2299 (N_2299,In_1476,In_1923);
and U2300 (N_2300,In_669,In_1381);
xnor U2301 (N_2301,In_650,In_265);
xor U2302 (N_2302,In_2454,In_50);
xor U2303 (N_2303,In_1975,In_1827);
nand U2304 (N_2304,In_1767,In_2340);
nand U2305 (N_2305,In_453,In_1420);
nand U2306 (N_2306,In_1486,In_1313);
or U2307 (N_2307,In_2380,In_1962);
or U2308 (N_2308,In_2410,In_385);
and U2309 (N_2309,In_2041,In_515);
nor U2310 (N_2310,In_2492,In_909);
nor U2311 (N_2311,In_1366,In_1212);
or U2312 (N_2312,In_2455,In_2118);
nand U2313 (N_2313,In_2333,In_1126);
and U2314 (N_2314,In_385,In_711);
and U2315 (N_2315,In_810,In_563);
nand U2316 (N_2316,In_216,In_1109);
and U2317 (N_2317,In_2099,In_239);
xnor U2318 (N_2318,In_802,In_2255);
nand U2319 (N_2319,In_1564,In_309);
and U2320 (N_2320,In_755,In_940);
xnor U2321 (N_2321,In_1317,In_1292);
nand U2322 (N_2322,In_226,In_1975);
and U2323 (N_2323,In_75,In_97);
or U2324 (N_2324,In_903,In_574);
xnor U2325 (N_2325,In_1223,In_54);
xnor U2326 (N_2326,In_1843,In_880);
xor U2327 (N_2327,In_1985,In_1427);
or U2328 (N_2328,In_1464,In_1587);
nor U2329 (N_2329,In_277,In_612);
and U2330 (N_2330,In_1345,In_1453);
or U2331 (N_2331,In_470,In_496);
xnor U2332 (N_2332,In_1386,In_1065);
nand U2333 (N_2333,In_1177,In_1117);
or U2334 (N_2334,In_55,In_831);
or U2335 (N_2335,In_242,In_1314);
nor U2336 (N_2336,In_1796,In_165);
nor U2337 (N_2337,In_2244,In_1807);
or U2338 (N_2338,In_2482,In_866);
nor U2339 (N_2339,In_904,In_1460);
and U2340 (N_2340,In_2423,In_2268);
nand U2341 (N_2341,In_1640,In_1742);
xnor U2342 (N_2342,In_134,In_1931);
nor U2343 (N_2343,In_2347,In_168);
nand U2344 (N_2344,In_1185,In_1753);
nand U2345 (N_2345,In_829,In_1431);
nand U2346 (N_2346,In_2081,In_1313);
or U2347 (N_2347,In_1714,In_814);
nor U2348 (N_2348,In_1404,In_1360);
nor U2349 (N_2349,In_667,In_895);
or U2350 (N_2350,In_2467,In_1475);
nor U2351 (N_2351,In_355,In_1185);
and U2352 (N_2352,In_216,In_415);
nor U2353 (N_2353,In_2222,In_1279);
xor U2354 (N_2354,In_1809,In_1112);
nand U2355 (N_2355,In_333,In_1969);
and U2356 (N_2356,In_961,In_622);
and U2357 (N_2357,In_907,In_750);
or U2358 (N_2358,In_1022,In_578);
nor U2359 (N_2359,In_1121,In_1809);
nand U2360 (N_2360,In_2332,In_231);
and U2361 (N_2361,In_1079,In_1822);
nand U2362 (N_2362,In_1493,In_1314);
nand U2363 (N_2363,In_281,In_494);
and U2364 (N_2364,In_284,In_252);
nand U2365 (N_2365,In_1689,In_1432);
nor U2366 (N_2366,In_1503,In_1302);
or U2367 (N_2367,In_256,In_1347);
nand U2368 (N_2368,In_1114,In_2291);
and U2369 (N_2369,In_1090,In_1532);
nand U2370 (N_2370,In_1736,In_2405);
or U2371 (N_2371,In_92,In_94);
nand U2372 (N_2372,In_1419,In_1494);
nor U2373 (N_2373,In_879,In_831);
nand U2374 (N_2374,In_846,In_1937);
nand U2375 (N_2375,In_1731,In_1067);
or U2376 (N_2376,In_1917,In_874);
nor U2377 (N_2377,In_5,In_486);
or U2378 (N_2378,In_1657,In_1936);
xnor U2379 (N_2379,In_1437,In_404);
nor U2380 (N_2380,In_1621,In_221);
nand U2381 (N_2381,In_1146,In_328);
nand U2382 (N_2382,In_371,In_2029);
or U2383 (N_2383,In_125,In_1158);
nor U2384 (N_2384,In_2030,In_824);
or U2385 (N_2385,In_1116,In_150);
xnor U2386 (N_2386,In_893,In_608);
nor U2387 (N_2387,In_703,In_195);
and U2388 (N_2388,In_1086,In_1793);
nand U2389 (N_2389,In_293,In_419);
or U2390 (N_2390,In_25,In_221);
nor U2391 (N_2391,In_136,In_2246);
xnor U2392 (N_2392,In_1279,In_2188);
nand U2393 (N_2393,In_828,In_1312);
and U2394 (N_2394,In_849,In_2116);
nor U2395 (N_2395,In_1414,In_1257);
or U2396 (N_2396,In_2044,In_1144);
xnor U2397 (N_2397,In_1246,In_2250);
and U2398 (N_2398,In_1420,In_2476);
xnor U2399 (N_2399,In_795,In_1611);
nand U2400 (N_2400,In_1759,In_899);
xor U2401 (N_2401,In_364,In_2328);
xor U2402 (N_2402,In_397,In_205);
xor U2403 (N_2403,In_1846,In_946);
nand U2404 (N_2404,In_1484,In_1907);
nor U2405 (N_2405,In_1206,In_1173);
and U2406 (N_2406,In_1453,In_2384);
or U2407 (N_2407,In_806,In_1753);
xor U2408 (N_2408,In_2489,In_806);
nor U2409 (N_2409,In_600,In_300);
or U2410 (N_2410,In_1940,In_637);
xnor U2411 (N_2411,In_449,In_2119);
nor U2412 (N_2412,In_1659,In_1145);
xor U2413 (N_2413,In_619,In_1031);
xor U2414 (N_2414,In_1518,In_2196);
or U2415 (N_2415,In_2491,In_1024);
nor U2416 (N_2416,In_1532,In_2393);
and U2417 (N_2417,In_921,In_360);
and U2418 (N_2418,In_2045,In_188);
nand U2419 (N_2419,In_2021,In_1705);
nor U2420 (N_2420,In_1358,In_2071);
nor U2421 (N_2421,In_1633,In_1459);
xor U2422 (N_2422,In_1716,In_2005);
and U2423 (N_2423,In_645,In_1811);
nor U2424 (N_2424,In_1542,In_998);
and U2425 (N_2425,In_451,In_519);
and U2426 (N_2426,In_1862,In_1658);
nand U2427 (N_2427,In_1602,In_1204);
nand U2428 (N_2428,In_990,In_157);
nand U2429 (N_2429,In_15,In_1892);
and U2430 (N_2430,In_985,In_929);
nor U2431 (N_2431,In_1694,In_1086);
nor U2432 (N_2432,In_1417,In_66);
nor U2433 (N_2433,In_2449,In_1831);
or U2434 (N_2434,In_1875,In_1062);
and U2435 (N_2435,In_2394,In_1113);
and U2436 (N_2436,In_285,In_2433);
or U2437 (N_2437,In_785,In_1596);
or U2438 (N_2438,In_1360,In_932);
and U2439 (N_2439,In_1701,In_1450);
nand U2440 (N_2440,In_828,In_1416);
xnor U2441 (N_2441,In_1929,In_547);
nand U2442 (N_2442,In_887,In_930);
nand U2443 (N_2443,In_0,In_1578);
nor U2444 (N_2444,In_156,In_1399);
xor U2445 (N_2445,In_1343,In_117);
nor U2446 (N_2446,In_57,In_1515);
or U2447 (N_2447,In_1849,In_1465);
nor U2448 (N_2448,In_284,In_868);
or U2449 (N_2449,In_885,In_1831);
xnor U2450 (N_2450,In_2092,In_323);
nor U2451 (N_2451,In_1636,In_1492);
nand U2452 (N_2452,In_689,In_117);
and U2453 (N_2453,In_525,In_93);
and U2454 (N_2454,In_402,In_189);
xnor U2455 (N_2455,In_1761,In_281);
nand U2456 (N_2456,In_596,In_724);
or U2457 (N_2457,In_1448,In_1200);
nor U2458 (N_2458,In_1490,In_2126);
nor U2459 (N_2459,In_1650,In_374);
or U2460 (N_2460,In_1372,In_542);
or U2461 (N_2461,In_2118,In_1918);
nor U2462 (N_2462,In_2284,In_356);
and U2463 (N_2463,In_1012,In_610);
xor U2464 (N_2464,In_132,In_587);
and U2465 (N_2465,In_1571,In_519);
or U2466 (N_2466,In_999,In_1231);
nand U2467 (N_2467,In_1424,In_1843);
or U2468 (N_2468,In_2111,In_1594);
nand U2469 (N_2469,In_1738,In_815);
nor U2470 (N_2470,In_2415,In_1435);
and U2471 (N_2471,In_1050,In_678);
nor U2472 (N_2472,In_1964,In_808);
or U2473 (N_2473,In_568,In_2430);
xnor U2474 (N_2474,In_548,In_1046);
or U2475 (N_2475,In_1751,In_1974);
and U2476 (N_2476,In_2294,In_1520);
or U2477 (N_2477,In_1194,In_1836);
nand U2478 (N_2478,In_672,In_230);
and U2479 (N_2479,In_2485,In_104);
nor U2480 (N_2480,In_2447,In_1685);
xor U2481 (N_2481,In_2154,In_2243);
or U2482 (N_2482,In_6,In_213);
and U2483 (N_2483,In_1067,In_1334);
xnor U2484 (N_2484,In_15,In_1875);
or U2485 (N_2485,In_1949,In_1921);
and U2486 (N_2486,In_2106,In_2177);
nor U2487 (N_2487,In_631,In_1282);
and U2488 (N_2488,In_704,In_1555);
nor U2489 (N_2489,In_1523,In_1432);
nand U2490 (N_2490,In_1254,In_2455);
nand U2491 (N_2491,In_631,In_1312);
or U2492 (N_2492,In_1085,In_1971);
and U2493 (N_2493,In_1842,In_414);
xor U2494 (N_2494,In_757,In_1408);
xor U2495 (N_2495,In_393,In_2469);
or U2496 (N_2496,In_1979,In_278);
xnor U2497 (N_2497,In_112,In_1242);
and U2498 (N_2498,In_791,In_2472);
and U2499 (N_2499,In_1466,In_798);
or U2500 (N_2500,In_1098,In_843);
nor U2501 (N_2501,In_1647,In_2194);
xnor U2502 (N_2502,In_101,In_790);
and U2503 (N_2503,In_681,In_957);
and U2504 (N_2504,In_722,In_76);
or U2505 (N_2505,In_2313,In_1661);
xnor U2506 (N_2506,In_285,In_380);
nor U2507 (N_2507,In_265,In_910);
xor U2508 (N_2508,In_1872,In_1397);
or U2509 (N_2509,In_2329,In_2386);
and U2510 (N_2510,In_1027,In_308);
or U2511 (N_2511,In_1745,In_1380);
or U2512 (N_2512,In_1253,In_95);
or U2513 (N_2513,In_533,In_1358);
nor U2514 (N_2514,In_2366,In_671);
nand U2515 (N_2515,In_591,In_1284);
nand U2516 (N_2516,In_2451,In_130);
nor U2517 (N_2517,In_1159,In_783);
xor U2518 (N_2518,In_1802,In_1570);
or U2519 (N_2519,In_2066,In_1092);
or U2520 (N_2520,In_1872,In_576);
nor U2521 (N_2521,In_2424,In_394);
and U2522 (N_2522,In_1674,In_1436);
nand U2523 (N_2523,In_2171,In_1164);
and U2524 (N_2524,In_614,In_2241);
xnor U2525 (N_2525,In_2059,In_481);
xnor U2526 (N_2526,In_371,In_2073);
and U2527 (N_2527,In_1996,In_90);
or U2528 (N_2528,In_2430,In_277);
or U2529 (N_2529,In_68,In_2408);
nor U2530 (N_2530,In_1708,In_1376);
xnor U2531 (N_2531,In_2113,In_1190);
nand U2532 (N_2532,In_2428,In_276);
xor U2533 (N_2533,In_1934,In_1493);
nand U2534 (N_2534,In_473,In_1012);
xor U2535 (N_2535,In_497,In_1527);
nand U2536 (N_2536,In_1885,In_1286);
and U2537 (N_2537,In_1439,In_1945);
and U2538 (N_2538,In_9,In_1693);
xnor U2539 (N_2539,In_1926,In_1648);
or U2540 (N_2540,In_160,In_52);
nor U2541 (N_2541,In_1065,In_819);
nor U2542 (N_2542,In_2290,In_1095);
xnor U2543 (N_2543,In_1853,In_769);
nand U2544 (N_2544,In_1674,In_1926);
nor U2545 (N_2545,In_758,In_2386);
nor U2546 (N_2546,In_1842,In_520);
nor U2547 (N_2547,In_1045,In_1537);
and U2548 (N_2548,In_2485,In_2177);
and U2549 (N_2549,In_224,In_931);
or U2550 (N_2550,In_2405,In_2168);
nand U2551 (N_2551,In_2349,In_1614);
xor U2552 (N_2552,In_112,In_1871);
nor U2553 (N_2553,In_591,In_481);
nand U2554 (N_2554,In_1942,In_1437);
nand U2555 (N_2555,In_1305,In_966);
or U2556 (N_2556,In_1047,In_1813);
and U2557 (N_2557,In_544,In_2127);
nor U2558 (N_2558,In_2085,In_792);
or U2559 (N_2559,In_1977,In_2256);
xnor U2560 (N_2560,In_693,In_1038);
or U2561 (N_2561,In_373,In_802);
nand U2562 (N_2562,In_355,In_1330);
and U2563 (N_2563,In_1670,In_411);
nor U2564 (N_2564,In_529,In_1457);
and U2565 (N_2565,In_2231,In_2341);
nand U2566 (N_2566,In_66,In_746);
or U2567 (N_2567,In_1288,In_1764);
xor U2568 (N_2568,In_1106,In_2111);
or U2569 (N_2569,In_1410,In_138);
nand U2570 (N_2570,In_1691,In_544);
nand U2571 (N_2571,In_2240,In_1259);
xor U2572 (N_2572,In_1120,In_732);
or U2573 (N_2573,In_569,In_1087);
or U2574 (N_2574,In_1002,In_396);
and U2575 (N_2575,In_2230,In_101);
nor U2576 (N_2576,In_427,In_1357);
xnor U2577 (N_2577,In_108,In_1007);
nand U2578 (N_2578,In_740,In_362);
nor U2579 (N_2579,In_69,In_61);
nand U2580 (N_2580,In_451,In_1465);
xnor U2581 (N_2581,In_2061,In_1051);
nand U2582 (N_2582,In_2356,In_914);
nand U2583 (N_2583,In_116,In_281);
xor U2584 (N_2584,In_855,In_808);
nor U2585 (N_2585,In_626,In_2411);
or U2586 (N_2586,In_2234,In_2112);
nor U2587 (N_2587,In_2271,In_1483);
xnor U2588 (N_2588,In_1824,In_148);
nand U2589 (N_2589,In_1528,In_2475);
nand U2590 (N_2590,In_641,In_2470);
nand U2591 (N_2591,In_1728,In_2347);
xnor U2592 (N_2592,In_2418,In_2008);
nor U2593 (N_2593,In_2438,In_77);
and U2594 (N_2594,In_954,In_1351);
xnor U2595 (N_2595,In_1989,In_667);
or U2596 (N_2596,In_2382,In_2458);
nand U2597 (N_2597,In_1795,In_1880);
or U2598 (N_2598,In_1432,In_639);
xnor U2599 (N_2599,In_365,In_1120);
and U2600 (N_2600,In_1832,In_841);
nand U2601 (N_2601,In_1490,In_956);
nand U2602 (N_2602,In_1485,In_1476);
xor U2603 (N_2603,In_190,In_1113);
xor U2604 (N_2604,In_1801,In_831);
xor U2605 (N_2605,In_650,In_980);
or U2606 (N_2606,In_1344,In_1662);
nand U2607 (N_2607,In_2030,In_1691);
and U2608 (N_2608,In_1082,In_93);
nand U2609 (N_2609,In_18,In_2067);
and U2610 (N_2610,In_2363,In_2103);
and U2611 (N_2611,In_994,In_498);
nor U2612 (N_2612,In_1954,In_1417);
xor U2613 (N_2613,In_458,In_740);
xnor U2614 (N_2614,In_2221,In_741);
nand U2615 (N_2615,In_34,In_1865);
or U2616 (N_2616,In_707,In_2041);
nand U2617 (N_2617,In_1896,In_1827);
xnor U2618 (N_2618,In_357,In_82);
and U2619 (N_2619,In_1628,In_1572);
nand U2620 (N_2620,In_2417,In_221);
xor U2621 (N_2621,In_1896,In_565);
and U2622 (N_2622,In_2111,In_847);
nor U2623 (N_2623,In_1308,In_753);
or U2624 (N_2624,In_679,In_2392);
nor U2625 (N_2625,In_1744,In_2120);
nand U2626 (N_2626,In_1291,In_1992);
nand U2627 (N_2627,In_1727,In_254);
nand U2628 (N_2628,In_1439,In_1813);
and U2629 (N_2629,In_338,In_1856);
nor U2630 (N_2630,In_940,In_1544);
and U2631 (N_2631,In_792,In_628);
nand U2632 (N_2632,In_203,In_1150);
or U2633 (N_2633,In_322,In_880);
nor U2634 (N_2634,In_583,In_264);
and U2635 (N_2635,In_368,In_369);
nand U2636 (N_2636,In_45,In_389);
xnor U2637 (N_2637,In_745,In_1515);
and U2638 (N_2638,In_164,In_1488);
xor U2639 (N_2639,In_381,In_2344);
xnor U2640 (N_2640,In_2251,In_1343);
xnor U2641 (N_2641,In_1919,In_176);
nand U2642 (N_2642,In_1506,In_2034);
nor U2643 (N_2643,In_1484,In_916);
xor U2644 (N_2644,In_1381,In_1486);
nor U2645 (N_2645,In_541,In_45);
and U2646 (N_2646,In_1712,In_1323);
and U2647 (N_2647,In_601,In_576);
nor U2648 (N_2648,In_1411,In_1524);
xor U2649 (N_2649,In_2329,In_390);
nand U2650 (N_2650,In_2189,In_1142);
and U2651 (N_2651,In_464,In_2155);
nor U2652 (N_2652,In_2202,In_1487);
nor U2653 (N_2653,In_575,In_464);
nor U2654 (N_2654,In_958,In_1924);
and U2655 (N_2655,In_1008,In_2242);
nor U2656 (N_2656,In_1745,In_1462);
or U2657 (N_2657,In_738,In_2087);
and U2658 (N_2658,In_543,In_1210);
and U2659 (N_2659,In_598,In_628);
nor U2660 (N_2660,In_520,In_361);
and U2661 (N_2661,In_577,In_2167);
and U2662 (N_2662,In_2416,In_152);
or U2663 (N_2663,In_2084,In_2232);
xnor U2664 (N_2664,In_1232,In_1703);
and U2665 (N_2665,In_1104,In_2444);
or U2666 (N_2666,In_345,In_999);
nor U2667 (N_2667,In_2044,In_1847);
nand U2668 (N_2668,In_1725,In_2431);
nand U2669 (N_2669,In_1791,In_2125);
nand U2670 (N_2670,In_1562,In_1994);
xnor U2671 (N_2671,In_1364,In_2405);
nand U2672 (N_2672,In_2233,In_221);
xnor U2673 (N_2673,In_2048,In_2068);
xnor U2674 (N_2674,In_2284,In_1171);
or U2675 (N_2675,In_550,In_1547);
xnor U2676 (N_2676,In_923,In_2066);
nand U2677 (N_2677,In_92,In_752);
nor U2678 (N_2678,In_115,In_738);
xor U2679 (N_2679,In_1886,In_50);
or U2680 (N_2680,In_2131,In_1579);
nor U2681 (N_2681,In_360,In_783);
nor U2682 (N_2682,In_1646,In_479);
nand U2683 (N_2683,In_754,In_1246);
or U2684 (N_2684,In_1675,In_1524);
or U2685 (N_2685,In_1409,In_194);
xnor U2686 (N_2686,In_1310,In_246);
and U2687 (N_2687,In_898,In_1012);
xor U2688 (N_2688,In_1119,In_1985);
nor U2689 (N_2689,In_627,In_759);
nor U2690 (N_2690,In_2037,In_1357);
xnor U2691 (N_2691,In_971,In_989);
nor U2692 (N_2692,In_2175,In_1225);
or U2693 (N_2693,In_172,In_2260);
or U2694 (N_2694,In_1032,In_1812);
and U2695 (N_2695,In_441,In_724);
xor U2696 (N_2696,In_925,In_25);
nor U2697 (N_2697,In_875,In_1156);
xor U2698 (N_2698,In_607,In_1120);
and U2699 (N_2699,In_1156,In_1840);
xor U2700 (N_2700,In_901,In_1406);
and U2701 (N_2701,In_997,In_1007);
nor U2702 (N_2702,In_1594,In_2255);
and U2703 (N_2703,In_1717,In_2338);
and U2704 (N_2704,In_382,In_2162);
nor U2705 (N_2705,In_254,In_2206);
xnor U2706 (N_2706,In_900,In_991);
nand U2707 (N_2707,In_160,In_1268);
xor U2708 (N_2708,In_450,In_1104);
nor U2709 (N_2709,In_23,In_1911);
nor U2710 (N_2710,In_2051,In_1830);
and U2711 (N_2711,In_252,In_793);
xor U2712 (N_2712,In_733,In_1248);
or U2713 (N_2713,In_555,In_364);
nor U2714 (N_2714,In_1389,In_1578);
xor U2715 (N_2715,In_2061,In_522);
xnor U2716 (N_2716,In_785,In_236);
nand U2717 (N_2717,In_2147,In_260);
nand U2718 (N_2718,In_61,In_211);
or U2719 (N_2719,In_1953,In_419);
nor U2720 (N_2720,In_2363,In_1227);
nor U2721 (N_2721,In_1095,In_23);
nand U2722 (N_2722,In_2261,In_1817);
or U2723 (N_2723,In_68,In_2209);
nor U2724 (N_2724,In_1816,In_1149);
or U2725 (N_2725,In_2082,In_1642);
nor U2726 (N_2726,In_390,In_239);
nand U2727 (N_2727,In_883,In_1301);
and U2728 (N_2728,In_695,In_1475);
or U2729 (N_2729,In_1185,In_1036);
and U2730 (N_2730,In_2338,In_212);
nor U2731 (N_2731,In_2084,In_1619);
nand U2732 (N_2732,In_312,In_313);
and U2733 (N_2733,In_611,In_1650);
and U2734 (N_2734,In_268,In_863);
xnor U2735 (N_2735,In_1116,In_517);
nand U2736 (N_2736,In_1497,In_851);
nor U2737 (N_2737,In_94,In_1480);
and U2738 (N_2738,In_1700,In_508);
nor U2739 (N_2739,In_617,In_174);
nand U2740 (N_2740,In_1245,In_508);
nor U2741 (N_2741,In_1334,In_450);
nor U2742 (N_2742,In_341,In_205);
nand U2743 (N_2743,In_1500,In_1565);
and U2744 (N_2744,In_542,In_488);
or U2745 (N_2745,In_595,In_1225);
nor U2746 (N_2746,In_972,In_1308);
xnor U2747 (N_2747,In_1446,In_2437);
nor U2748 (N_2748,In_1959,In_30);
nand U2749 (N_2749,In_2314,In_538);
xor U2750 (N_2750,In_126,In_419);
or U2751 (N_2751,In_77,In_1641);
nor U2752 (N_2752,In_1299,In_365);
or U2753 (N_2753,In_2437,In_278);
or U2754 (N_2754,In_1343,In_1578);
and U2755 (N_2755,In_682,In_147);
or U2756 (N_2756,In_1400,In_1634);
nor U2757 (N_2757,In_885,In_1963);
nor U2758 (N_2758,In_1696,In_1013);
xor U2759 (N_2759,In_1833,In_1436);
or U2760 (N_2760,In_257,In_2390);
nor U2761 (N_2761,In_1068,In_966);
nor U2762 (N_2762,In_85,In_2332);
and U2763 (N_2763,In_955,In_1509);
nand U2764 (N_2764,In_1223,In_505);
nand U2765 (N_2765,In_799,In_1343);
xnor U2766 (N_2766,In_2418,In_1698);
nor U2767 (N_2767,In_2302,In_837);
or U2768 (N_2768,In_106,In_1261);
nand U2769 (N_2769,In_633,In_2372);
or U2770 (N_2770,In_1811,In_2079);
or U2771 (N_2771,In_1994,In_116);
nand U2772 (N_2772,In_171,In_1778);
or U2773 (N_2773,In_428,In_2343);
or U2774 (N_2774,In_260,In_1714);
nand U2775 (N_2775,In_1798,In_1725);
xnor U2776 (N_2776,In_1833,In_2081);
xor U2777 (N_2777,In_1252,In_165);
nor U2778 (N_2778,In_271,In_1917);
and U2779 (N_2779,In_1898,In_2401);
and U2780 (N_2780,In_426,In_881);
xnor U2781 (N_2781,In_1349,In_882);
nand U2782 (N_2782,In_2320,In_2470);
and U2783 (N_2783,In_2009,In_1991);
and U2784 (N_2784,In_277,In_2105);
and U2785 (N_2785,In_17,In_186);
or U2786 (N_2786,In_985,In_176);
and U2787 (N_2787,In_2146,In_871);
xnor U2788 (N_2788,In_810,In_1525);
or U2789 (N_2789,In_1861,In_1919);
and U2790 (N_2790,In_1441,In_679);
nor U2791 (N_2791,In_2261,In_743);
or U2792 (N_2792,In_514,In_1461);
nand U2793 (N_2793,In_2361,In_292);
and U2794 (N_2794,In_2459,In_2351);
nor U2795 (N_2795,In_466,In_1080);
and U2796 (N_2796,In_1316,In_591);
nor U2797 (N_2797,In_1277,In_411);
xor U2798 (N_2798,In_2340,In_1654);
and U2799 (N_2799,In_794,In_1205);
or U2800 (N_2800,In_418,In_975);
xnor U2801 (N_2801,In_2211,In_2073);
xnor U2802 (N_2802,In_594,In_1171);
nand U2803 (N_2803,In_2486,In_1309);
and U2804 (N_2804,In_1427,In_146);
nor U2805 (N_2805,In_1098,In_1185);
nor U2806 (N_2806,In_2111,In_1558);
nand U2807 (N_2807,In_1482,In_1539);
xnor U2808 (N_2808,In_2265,In_2279);
and U2809 (N_2809,In_1788,In_11);
xor U2810 (N_2810,In_805,In_634);
and U2811 (N_2811,In_1624,In_720);
or U2812 (N_2812,In_590,In_713);
nor U2813 (N_2813,In_543,In_1882);
or U2814 (N_2814,In_178,In_2145);
or U2815 (N_2815,In_1559,In_1632);
nor U2816 (N_2816,In_928,In_1837);
or U2817 (N_2817,In_1236,In_87);
and U2818 (N_2818,In_278,In_1666);
nor U2819 (N_2819,In_2089,In_70);
nor U2820 (N_2820,In_2197,In_587);
and U2821 (N_2821,In_2305,In_983);
xnor U2822 (N_2822,In_479,In_369);
or U2823 (N_2823,In_834,In_398);
nand U2824 (N_2824,In_1716,In_1043);
xnor U2825 (N_2825,In_1758,In_1031);
nor U2826 (N_2826,In_332,In_614);
nor U2827 (N_2827,In_1828,In_2443);
and U2828 (N_2828,In_1078,In_504);
nor U2829 (N_2829,In_1155,In_2005);
nand U2830 (N_2830,In_1618,In_552);
nand U2831 (N_2831,In_1409,In_961);
nand U2832 (N_2832,In_1906,In_618);
xnor U2833 (N_2833,In_1737,In_1214);
and U2834 (N_2834,In_2336,In_1136);
nor U2835 (N_2835,In_2193,In_141);
xor U2836 (N_2836,In_1785,In_1624);
nor U2837 (N_2837,In_765,In_1746);
and U2838 (N_2838,In_438,In_2350);
nand U2839 (N_2839,In_1271,In_1181);
xor U2840 (N_2840,In_1674,In_954);
xor U2841 (N_2841,In_2234,In_1051);
or U2842 (N_2842,In_568,In_2267);
or U2843 (N_2843,In_1361,In_237);
nand U2844 (N_2844,In_2105,In_1776);
and U2845 (N_2845,In_2040,In_617);
and U2846 (N_2846,In_1526,In_573);
nand U2847 (N_2847,In_375,In_2484);
or U2848 (N_2848,In_976,In_1618);
nor U2849 (N_2849,In_717,In_791);
nand U2850 (N_2850,In_150,In_1492);
or U2851 (N_2851,In_787,In_2420);
or U2852 (N_2852,In_2284,In_2224);
or U2853 (N_2853,In_2199,In_1023);
xnor U2854 (N_2854,In_2300,In_1826);
nand U2855 (N_2855,In_905,In_1731);
xnor U2856 (N_2856,In_1430,In_2371);
nor U2857 (N_2857,In_1244,In_482);
or U2858 (N_2858,In_1237,In_1870);
and U2859 (N_2859,In_401,In_321);
nand U2860 (N_2860,In_7,In_1239);
xnor U2861 (N_2861,In_26,In_803);
nand U2862 (N_2862,In_1521,In_2259);
and U2863 (N_2863,In_2284,In_1368);
xor U2864 (N_2864,In_1693,In_1194);
and U2865 (N_2865,In_799,In_1422);
nand U2866 (N_2866,In_191,In_1299);
or U2867 (N_2867,In_57,In_1982);
nand U2868 (N_2868,In_168,In_473);
or U2869 (N_2869,In_220,In_1416);
nand U2870 (N_2870,In_118,In_2298);
nor U2871 (N_2871,In_2113,In_172);
and U2872 (N_2872,In_1237,In_589);
nand U2873 (N_2873,In_1418,In_893);
xnor U2874 (N_2874,In_2045,In_1169);
nor U2875 (N_2875,In_369,In_2398);
and U2876 (N_2876,In_363,In_252);
xnor U2877 (N_2877,In_1684,In_1845);
nand U2878 (N_2878,In_243,In_1303);
xor U2879 (N_2879,In_1076,In_2377);
nor U2880 (N_2880,In_455,In_2165);
and U2881 (N_2881,In_1864,In_360);
nand U2882 (N_2882,In_1485,In_650);
xor U2883 (N_2883,In_1117,In_592);
xnor U2884 (N_2884,In_2376,In_1628);
and U2885 (N_2885,In_1946,In_2024);
and U2886 (N_2886,In_1743,In_1404);
and U2887 (N_2887,In_298,In_812);
and U2888 (N_2888,In_216,In_1574);
or U2889 (N_2889,In_395,In_2295);
and U2890 (N_2890,In_1465,In_1847);
xnor U2891 (N_2891,In_373,In_615);
xor U2892 (N_2892,In_405,In_2204);
nor U2893 (N_2893,In_1417,In_2418);
and U2894 (N_2894,In_500,In_1705);
nor U2895 (N_2895,In_1316,In_1765);
and U2896 (N_2896,In_117,In_1775);
or U2897 (N_2897,In_1567,In_1488);
or U2898 (N_2898,In_2202,In_1750);
nor U2899 (N_2899,In_122,In_355);
or U2900 (N_2900,In_1157,In_1053);
nor U2901 (N_2901,In_919,In_2462);
nor U2902 (N_2902,In_1741,In_1102);
or U2903 (N_2903,In_480,In_2226);
nand U2904 (N_2904,In_782,In_2238);
nor U2905 (N_2905,In_2363,In_301);
or U2906 (N_2906,In_2074,In_1125);
and U2907 (N_2907,In_1862,In_697);
and U2908 (N_2908,In_700,In_433);
or U2909 (N_2909,In_2122,In_727);
and U2910 (N_2910,In_507,In_2386);
nand U2911 (N_2911,In_572,In_662);
xnor U2912 (N_2912,In_881,In_1152);
xnor U2913 (N_2913,In_2271,In_1);
and U2914 (N_2914,In_2488,In_1886);
and U2915 (N_2915,In_542,In_1814);
xor U2916 (N_2916,In_1548,In_424);
nor U2917 (N_2917,In_1231,In_2468);
nor U2918 (N_2918,In_1209,In_954);
xnor U2919 (N_2919,In_1087,In_1662);
nor U2920 (N_2920,In_2345,In_1415);
xor U2921 (N_2921,In_1191,In_1842);
xnor U2922 (N_2922,In_1383,In_1733);
nand U2923 (N_2923,In_123,In_1801);
and U2924 (N_2924,In_723,In_2097);
nand U2925 (N_2925,In_1992,In_489);
nand U2926 (N_2926,In_657,In_2179);
and U2927 (N_2927,In_302,In_933);
nand U2928 (N_2928,In_1711,In_1211);
and U2929 (N_2929,In_1668,In_852);
and U2930 (N_2930,In_320,In_1029);
or U2931 (N_2931,In_2129,In_1878);
nor U2932 (N_2932,In_438,In_2394);
xor U2933 (N_2933,In_1043,In_1767);
xor U2934 (N_2934,In_2177,In_1889);
and U2935 (N_2935,In_1098,In_377);
or U2936 (N_2936,In_529,In_2111);
nand U2937 (N_2937,In_399,In_1861);
xor U2938 (N_2938,In_941,In_3);
and U2939 (N_2939,In_62,In_2347);
nor U2940 (N_2940,In_1130,In_2298);
or U2941 (N_2941,In_1552,In_200);
nand U2942 (N_2942,In_545,In_2440);
nand U2943 (N_2943,In_1625,In_1830);
xnor U2944 (N_2944,In_75,In_1431);
nor U2945 (N_2945,In_387,In_906);
and U2946 (N_2946,In_383,In_46);
and U2947 (N_2947,In_251,In_1800);
nor U2948 (N_2948,In_1056,In_1441);
and U2949 (N_2949,In_2388,In_1255);
and U2950 (N_2950,In_497,In_1158);
or U2951 (N_2951,In_2274,In_182);
nand U2952 (N_2952,In_2281,In_2449);
xnor U2953 (N_2953,In_2316,In_1411);
and U2954 (N_2954,In_1901,In_2397);
nor U2955 (N_2955,In_2453,In_1146);
and U2956 (N_2956,In_997,In_275);
or U2957 (N_2957,In_2312,In_1190);
nand U2958 (N_2958,In_141,In_1501);
or U2959 (N_2959,In_711,In_1729);
nor U2960 (N_2960,In_567,In_655);
nand U2961 (N_2961,In_227,In_1119);
or U2962 (N_2962,In_154,In_964);
nor U2963 (N_2963,In_1994,In_2256);
nor U2964 (N_2964,In_1172,In_668);
xnor U2965 (N_2965,In_2485,In_1429);
xnor U2966 (N_2966,In_450,In_798);
and U2967 (N_2967,In_31,In_369);
nor U2968 (N_2968,In_1863,In_996);
xor U2969 (N_2969,In_1626,In_2359);
or U2970 (N_2970,In_472,In_2236);
xnor U2971 (N_2971,In_2175,In_1273);
nor U2972 (N_2972,In_333,In_133);
or U2973 (N_2973,In_1309,In_2328);
or U2974 (N_2974,In_720,In_1369);
nand U2975 (N_2975,In_1765,In_2354);
or U2976 (N_2976,In_1142,In_2367);
or U2977 (N_2977,In_1803,In_1588);
nand U2978 (N_2978,In_1586,In_125);
xnor U2979 (N_2979,In_716,In_2241);
or U2980 (N_2980,In_139,In_1670);
xor U2981 (N_2981,In_1849,In_154);
nand U2982 (N_2982,In_2176,In_1850);
and U2983 (N_2983,In_1105,In_166);
nor U2984 (N_2984,In_2381,In_69);
nor U2985 (N_2985,In_1583,In_1938);
or U2986 (N_2986,In_788,In_601);
nor U2987 (N_2987,In_1129,In_834);
nor U2988 (N_2988,In_464,In_1418);
or U2989 (N_2989,In_1906,In_82);
xor U2990 (N_2990,In_772,In_1670);
and U2991 (N_2991,In_345,In_867);
nand U2992 (N_2992,In_1073,In_479);
xor U2993 (N_2993,In_446,In_730);
or U2994 (N_2994,In_767,In_895);
and U2995 (N_2995,In_1732,In_1729);
or U2996 (N_2996,In_1936,In_1297);
nand U2997 (N_2997,In_1839,In_1943);
xnor U2998 (N_2998,In_1412,In_1158);
or U2999 (N_2999,In_1250,In_1696);
or U3000 (N_3000,In_104,In_1164);
and U3001 (N_3001,In_937,In_142);
xor U3002 (N_3002,In_2263,In_828);
nand U3003 (N_3003,In_1635,In_1317);
nand U3004 (N_3004,In_405,In_925);
and U3005 (N_3005,In_2257,In_1909);
nand U3006 (N_3006,In_1404,In_1912);
and U3007 (N_3007,In_2104,In_169);
and U3008 (N_3008,In_1518,In_984);
nand U3009 (N_3009,In_2067,In_1226);
xnor U3010 (N_3010,In_2440,In_1127);
xnor U3011 (N_3011,In_2190,In_972);
and U3012 (N_3012,In_778,In_534);
or U3013 (N_3013,In_2044,In_2475);
or U3014 (N_3014,In_236,In_628);
nand U3015 (N_3015,In_2446,In_1768);
or U3016 (N_3016,In_1518,In_1368);
xor U3017 (N_3017,In_1961,In_157);
and U3018 (N_3018,In_1117,In_891);
or U3019 (N_3019,In_1565,In_2161);
nand U3020 (N_3020,In_111,In_1317);
or U3021 (N_3021,In_700,In_1084);
xnor U3022 (N_3022,In_1539,In_970);
or U3023 (N_3023,In_770,In_499);
xnor U3024 (N_3024,In_671,In_966);
and U3025 (N_3025,In_906,In_1582);
xor U3026 (N_3026,In_395,In_1348);
or U3027 (N_3027,In_462,In_855);
or U3028 (N_3028,In_142,In_710);
nor U3029 (N_3029,In_671,In_569);
or U3030 (N_3030,In_2414,In_646);
or U3031 (N_3031,In_1383,In_2068);
or U3032 (N_3032,In_187,In_398);
nand U3033 (N_3033,In_424,In_1732);
xnor U3034 (N_3034,In_282,In_306);
nand U3035 (N_3035,In_1578,In_834);
nor U3036 (N_3036,In_792,In_846);
nor U3037 (N_3037,In_2337,In_1852);
xnor U3038 (N_3038,In_5,In_1694);
xor U3039 (N_3039,In_1517,In_2124);
or U3040 (N_3040,In_77,In_1475);
or U3041 (N_3041,In_2399,In_1511);
nor U3042 (N_3042,In_206,In_433);
nor U3043 (N_3043,In_1122,In_143);
and U3044 (N_3044,In_47,In_340);
xnor U3045 (N_3045,In_2249,In_1631);
xor U3046 (N_3046,In_2263,In_1690);
nor U3047 (N_3047,In_769,In_2284);
and U3048 (N_3048,In_579,In_2225);
nor U3049 (N_3049,In_1468,In_485);
nand U3050 (N_3050,In_1441,In_1924);
nand U3051 (N_3051,In_242,In_1508);
nand U3052 (N_3052,In_1145,In_858);
nand U3053 (N_3053,In_1414,In_1355);
nor U3054 (N_3054,In_467,In_1301);
nor U3055 (N_3055,In_1987,In_993);
and U3056 (N_3056,In_1197,In_1092);
nor U3057 (N_3057,In_2172,In_2009);
nor U3058 (N_3058,In_1716,In_912);
nand U3059 (N_3059,In_225,In_1927);
nand U3060 (N_3060,In_1240,In_2142);
or U3061 (N_3061,In_178,In_1679);
xor U3062 (N_3062,In_1693,In_707);
nand U3063 (N_3063,In_347,In_2278);
xor U3064 (N_3064,In_581,In_1619);
xor U3065 (N_3065,In_1305,In_605);
xnor U3066 (N_3066,In_887,In_855);
and U3067 (N_3067,In_1386,In_39);
nor U3068 (N_3068,In_1258,In_1137);
nor U3069 (N_3069,In_863,In_1395);
nand U3070 (N_3070,In_2371,In_835);
xor U3071 (N_3071,In_637,In_1141);
and U3072 (N_3072,In_1692,In_1560);
nand U3073 (N_3073,In_1420,In_958);
or U3074 (N_3074,In_2099,In_1293);
or U3075 (N_3075,In_220,In_902);
or U3076 (N_3076,In_2051,In_2027);
nor U3077 (N_3077,In_1649,In_1589);
nand U3078 (N_3078,In_560,In_2269);
nor U3079 (N_3079,In_664,In_577);
and U3080 (N_3080,In_1722,In_1027);
and U3081 (N_3081,In_1159,In_487);
xnor U3082 (N_3082,In_220,In_1077);
and U3083 (N_3083,In_1709,In_2418);
nor U3084 (N_3084,In_2358,In_876);
nand U3085 (N_3085,In_793,In_2302);
nor U3086 (N_3086,In_1911,In_130);
nor U3087 (N_3087,In_880,In_1095);
or U3088 (N_3088,In_1629,In_838);
xor U3089 (N_3089,In_16,In_1474);
or U3090 (N_3090,In_2124,In_776);
and U3091 (N_3091,In_1934,In_152);
or U3092 (N_3092,In_248,In_1920);
and U3093 (N_3093,In_1134,In_622);
nand U3094 (N_3094,In_190,In_794);
nand U3095 (N_3095,In_1763,In_1431);
nand U3096 (N_3096,In_2089,In_1068);
nand U3097 (N_3097,In_867,In_1516);
or U3098 (N_3098,In_1274,In_1060);
nor U3099 (N_3099,In_2434,In_1546);
and U3100 (N_3100,In_1040,In_2005);
nor U3101 (N_3101,In_1505,In_1009);
nor U3102 (N_3102,In_621,In_2012);
xor U3103 (N_3103,In_1852,In_927);
and U3104 (N_3104,In_1252,In_127);
xor U3105 (N_3105,In_1667,In_81);
xor U3106 (N_3106,In_1800,In_2342);
xor U3107 (N_3107,In_2128,In_1324);
and U3108 (N_3108,In_205,In_936);
and U3109 (N_3109,In_187,In_682);
and U3110 (N_3110,In_709,In_749);
or U3111 (N_3111,In_2088,In_2328);
or U3112 (N_3112,In_1453,In_955);
nand U3113 (N_3113,In_675,In_1386);
nor U3114 (N_3114,In_2192,In_1457);
xor U3115 (N_3115,In_1850,In_104);
and U3116 (N_3116,In_370,In_1971);
nor U3117 (N_3117,In_1230,In_1411);
nand U3118 (N_3118,In_617,In_867);
and U3119 (N_3119,In_1607,In_1338);
nor U3120 (N_3120,In_1320,In_1737);
and U3121 (N_3121,In_2079,In_124);
xor U3122 (N_3122,In_2213,In_340);
xor U3123 (N_3123,In_906,In_2225);
xor U3124 (N_3124,In_2201,In_928);
nor U3125 (N_3125,In_1502,In_2144);
xnor U3126 (N_3126,In_752,In_105);
nand U3127 (N_3127,In_2445,In_2142);
nand U3128 (N_3128,In_327,In_109);
nand U3129 (N_3129,In_325,In_1183);
nor U3130 (N_3130,In_433,In_1987);
nand U3131 (N_3131,In_148,In_1264);
and U3132 (N_3132,In_2088,In_1864);
nand U3133 (N_3133,In_1188,In_298);
and U3134 (N_3134,In_618,In_675);
nor U3135 (N_3135,In_1156,In_843);
and U3136 (N_3136,In_2083,In_528);
nand U3137 (N_3137,In_1105,In_1698);
or U3138 (N_3138,In_1082,In_1710);
or U3139 (N_3139,In_1500,In_1010);
xor U3140 (N_3140,In_1214,In_295);
or U3141 (N_3141,In_1414,In_761);
or U3142 (N_3142,In_1721,In_1481);
nor U3143 (N_3143,In_832,In_2477);
and U3144 (N_3144,In_984,In_1118);
or U3145 (N_3145,In_14,In_726);
xnor U3146 (N_3146,In_1141,In_49);
and U3147 (N_3147,In_360,In_1539);
nand U3148 (N_3148,In_1414,In_355);
nor U3149 (N_3149,In_692,In_204);
or U3150 (N_3150,In_602,In_2363);
or U3151 (N_3151,In_1261,In_140);
nor U3152 (N_3152,In_2196,In_589);
nor U3153 (N_3153,In_2439,In_758);
and U3154 (N_3154,In_63,In_2401);
or U3155 (N_3155,In_1751,In_480);
or U3156 (N_3156,In_265,In_603);
and U3157 (N_3157,In_1798,In_1815);
nand U3158 (N_3158,In_1257,In_1737);
xor U3159 (N_3159,In_2324,In_1496);
xnor U3160 (N_3160,In_240,In_290);
nand U3161 (N_3161,In_948,In_1875);
nand U3162 (N_3162,In_1728,In_545);
and U3163 (N_3163,In_1736,In_1040);
or U3164 (N_3164,In_2239,In_188);
and U3165 (N_3165,In_988,In_1357);
nand U3166 (N_3166,In_548,In_2227);
xor U3167 (N_3167,In_1923,In_2093);
nand U3168 (N_3168,In_2336,In_2330);
and U3169 (N_3169,In_1244,In_559);
or U3170 (N_3170,In_1904,In_2150);
nand U3171 (N_3171,In_2299,In_730);
nand U3172 (N_3172,In_86,In_1322);
nand U3173 (N_3173,In_207,In_1147);
or U3174 (N_3174,In_857,In_815);
nor U3175 (N_3175,In_2208,In_2213);
xor U3176 (N_3176,In_520,In_1763);
or U3177 (N_3177,In_659,In_986);
nor U3178 (N_3178,In_1921,In_905);
or U3179 (N_3179,In_58,In_1955);
nand U3180 (N_3180,In_1335,In_560);
nand U3181 (N_3181,In_114,In_1481);
nor U3182 (N_3182,In_683,In_134);
nand U3183 (N_3183,In_1526,In_2062);
nand U3184 (N_3184,In_440,In_1309);
nor U3185 (N_3185,In_1418,In_128);
or U3186 (N_3186,In_624,In_785);
and U3187 (N_3187,In_1359,In_1363);
and U3188 (N_3188,In_340,In_468);
nor U3189 (N_3189,In_78,In_1321);
nor U3190 (N_3190,In_1714,In_2128);
xor U3191 (N_3191,In_1354,In_2282);
or U3192 (N_3192,In_1015,In_1167);
and U3193 (N_3193,In_1627,In_1588);
nand U3194 (N_3194,In_718,In_1691);
nand U3195 (N_3195,In_737,In_295);
nor U3196 (N_3196,In_2497,In_384);
xor U3197 (N_3197,In_890,In_1944);
nand U3198 (N_3198,In_697,In_2289);
nand U3199 (N_3199,In_1671,In_1592);
xnor U3200 (N_3200,In_1619,In_1042);
and U3201 (N_3201,In_2476,In_164);
nand U3202 (N_3202,In_320,In_71);
or U3203 (N_3203,In_1157,In_774);
or U3204 (N_3204,In_2313,In_1711);
and U3205 (N_3205,In_1379,In_2201);
xnor U3206 (N_3206,In_655,In_890);
nand U3207 (N_3207,In_277,In_640);
and U3208 (N_3208,In_1298,In_2357);
xor U3209 (N_3209,In_1673,In_2381);
and U3210 (N_3210,In_2340,In_1702);
nor U3211 (N_3211,In_966,In_1362);
or U3212 (N_3212,In_1822,In_2052);
xnor U3213 (N_3213,In_1534,In_1655);
and U3214 (N_3214,In_1229,In_2124);
nand U3215 (N_3215,In_725,In_1422);
nand U3216 (N_3216,In_774,In_560);
or U3217 (N_3217,In_2369,In_1300);
and U3218 (N_3218,In_299,In_637);
nor U3219 (N_3219,In_246,In_624);
nand U3220 (N_3220,In_2050,In_2376);
or U3221 (N_3221,In_88,In_1409);
or U3222 (N_3222,In_2020,In_1125);
xor U3223 (N_3223,In_1097,In_2036);
xor U3224 (N_3224,In_1851,In_44);
nor U3225 (N_3225,In_1568,In_34);
and U3226 (N_3226,In_2172,In_1415);
and U3227 (N_3227,In_1155,In_393);
nand U3228 (N_3228,In_218,In_1494);
and U3229 (N_3229,In_2445,In_1264);
nand U3230 (N_3230,In_918,In_115);
and U3231 (N_3231,In_1510,In_181);
or U3232 (N_3232,In_349,In_1010);
nor U3233 (N_3233,In_223,In_312);
or U3234 (N_3234,In_1733,In_1468);
or U3235 (N_3235,In_2383,In_1533);
or U3236 (N_3236,In_2213,In_1527);
xnor U3237 (N_3237,In_1694,In_2243);
and U3238 (N_3238,In_408,In_2275);
or U3239 (N_3239,In_1107,In_1310);
nor U3240 (N_3240,In_1517,In_1482);
and U3241 (N_3241,In_404,In_788);
nand U3242 (N_3242,In_1073,In_198);
xnor U3243 (N_3243,In_1145,In_1412);
and U3244 (N_3244,In_2444,In_1954);
and U3245 (N_3245,In_2311,In_662);
nor U3246 (N_3246,In_1365,In_163);
nor U3247 (N_3247,In_113,In_561);
or U3248 (N_3248,In_2227,In_1984);
nand U3249 (N_3249,In_399,In_2050);
or U3250 (N_3250,In_1323,In_120);
xor U3251 (N_3251,In_1155,In_1);
or U3252 (N_3252,In_1682,In_1945);
nand U3253 (N_3253,In_246,In_23);
xor U3254 (N_3254,In_703,In_993);
nand U3255 (N_3255,In_636,In_840);
nand U3256 (N_3256,In_139,In_2152);
nand U3257 (N_3257,In_750,In_2303);
nand U3258 (N_3258,In_1486,In_1472);
xor U3259 (N_3259,In_2215,In_233);
nor U3260 (N_3260,In_97,In_1546);
and U3261 (N_3261,In_513,In_2158);
and U3262 (N_3262,In_549,In_277);
nand U3263 (N_3263,In_344,In_1381);
nor U3264 (N_3264,In_2243,In_2226);
nand U3265 (N_3265,In_1466,In_1002);
nand U3266 (N_3266,In_2218,In_742);
nor U3267 (N_3267,In_2182,In_918);
or U3268 (N_3268,In_1003,In_2306);
and U3269 (N_3269,In_985,In_1128);
and U3270 (N_3270,In_1669,In_232);
or U3271 (N_3271,In_406,In_252);
nand U3272 (N_3272,In_1873,In_2045);
nand U3273 (N_3273,In_1212,In_674);
or U3274 (N_3274,In_1334,In_1507);
nand U3275 (N_3275,In_166,In_795);
and U3276 (N_3276,In_480,In_1395);
and U3277 (N_3277,In_2110,In_1716);
nor U3278 (N_3278,In_837,In_60);
xnor U3279 (N_3279,In_1980,In_251);
or U3280 (N_3280,In_2424,In_1337);
and U3281 (N_3281,In_983,In_1903);
and U3282 (N_3282,In_2061,In_46);
nor U3283 (N_3283,In_1596,In_70);
or U3284 (N_3284,In_902,In_1034);
xnor U3285 (N_3285,In_2454,In_1024);
nor U3286 (N_3286,In_960,In_480);
xor U3287 (N_3287,In_977,In_1181);
xor U3288 (N_3288,In_1828,In_2224);
xor U3289 (N_3289,In_1396,In_430);
nand U3290 (N_3290,In_18,In_1115);
nand U3291 (N_3291,In_1307,In_1618);
nand U3292 (N_3292,In_2117,In_2075);
nor U3293 (N_3293,In_2005,In_488);
nor U3294 (N_3294,In_598,In_2316);
xnor U3295 (N_3295,In_2364,In_1803);
nor U3296 (N_3296,In_642,In_1618);
or U3297 (N_3297,In_1136,In_2462);
nor U3298 (N_3298,In_1765,In_492);
nor U3299 (N_3299,In_143,In_514);
xnor U3300 (N_3300,In_536,In_2155);
xnor U3301 (N_3301,In_1283,In_1990);
xnor U3302 (N_3302,In_1522,In_632);
or U3303 (N_3303,In_950,In_1764);
or U3304 (N_3304,In_1593,In_2411);
nor U3305 (N_3305,In_2038,In_2445);
nor U3306 (N_3306,In_2483,In_2220);
nand U3307 (N_3307,In_666,In_2478);
or U3308 (N_3308,In_2230,In_1521);
nor U3309 (N_3309,In_1689,In_221);
xor U3310 (N_3310,In_115,In_1108);
and U3311 (N_3311,In_2399,In_144);
or U3312 (N_3312,In_2007,In_2420);
nor U3313 (N_3313,In_411,In_720);
xor U3314 (N_3314,In_1195,In_2188);
and U3315 (N_3315,In_2272,In_1069);
nor U3316 (N_3316,In_508,In_2014);
and U3317 (N_3317,In_2234,In_1702);
and U3318 (N_3318,In_943,In_1734);
and U3319 (N_3319,In_1164,In_1041);
nand U3320 (N_3320,In_251,In_2338);
nand U3321 (N_3321,In_1287,In_78);
or U3322 (N_3322,In_792,In_28);
nor U3323 (N_3323,In_170,In_509);
nor U3324 (N_3324,In_300,In_1758);
xor U3325 (N_3325,In_1932,In_1685);
xor U3326 (N_3326,In_1446,In_2251);
xnor U3327 (N_3327,In_270,In_793);
xnor U3328 (N_3328,In_1807,In_2342);
nand U3329 (N_3329,In_1662,In_1177);
xnor U3330 (N_3330,In_437,In_801);
xnor U3331 (N_3331,In_677,In_126);
nor U3332 (N_3332,In_2038,In_1558);
nor U3333 (N_3333,In_2075,In_475);
nor U3334 (N_3334,In_1444,In_175);
nor U3335 (N_3335,In_569,In_1937);
and U3336 (N_3336,In_399,In_311);
or U3337 (N_3337,In_413,In_1150);
nand U3338 (N_3338,In_151,In_1779);
or U3339 (N_3339,In_2143,In_1504);
and U3340 (N_3340,In_1237,In_1825);
nor U3341 (N_3341,In_1314,In_1222);
and U3342 (N_3342,In_528,In_1280);
and U3343 (N_3343,In_1704,In_147);
and U3344 (N_3344,In_1936,In_1432);
or U3345 (N_3345,In_367,In_1536);
xor U3346 (N_3346,In_1349,In_1375);
or U3347 (N_3347,In_1466,In_670);
or U3348 (N_3348,In_102,In_1939);
xnor U3349 (N_3349,In_2002,In_1897);
nand U3350 (N_3350,In_2468,In_1596);
nand U3351 (N_3351,In_883,In_317);
and U3352 (N_3352,In_1255,In_1466);
nor U3353 (N_3353,In_506,In_1138);
nor U3354 (N_3354,In_931,In_1132);
nor U3355 (N_3355,In_1531,In_394);
and U3356 (N_3356,In_198,In_1887);
and U3357 (N_3357,In_2140,In_1904);
or U3358 (N_3358,In_355,In_1387);
nor U3359 (N_3359,In_2047,In_2199);
nor U3360 (N_3360,In_1358,In_2391);
and U3361 (N_3361,In_1390,In_581);
nor U3362 (N_3362,In_525,In_307);
xnor U3363 (N_3363,In_1337,In_729);
and U3364 (N_3364,In_2263,In_636);
and U3365 (N_3365,In_878,In_1721);
nand U3366 (N_3366,In_806,In_864);
and U3367 (N_3367,In_307,In_1350);
xnor U3368 (N_3368,In_659,In_583);
xor U3369 (N_3369,In_497,In_100);
nand U3370 (N_3370,In_610,In_1496);
and U3371 (N_3371,In_955,In_1868);
nor U3372 (N_3372,In_1452,In_2202);
and U3373 (N_3373,In_863,In_140);
xnor U3374 (N_3374,In_259,In_2169);
nand U3375 (N_3375,In_2327,In_2090);
nand U3376 (N_3376,In_2063,In_604);
nor U3377 (N_3377,In_1736,In_1784);
nor U3378 (N_3378,In_980,In_2410);
nor U3379 (N_3379,In_1823,In_1845);
nor U3380 (N_3380,In_161,In_2308);
and U3381 (N_3381,In_2371,In_1975);
or U3382 (N_3382,In_1821,In_1337);
and U3383 (N_3383,In_1473,In_234);
xor U3384 (N_3384,In_1281,In_1355);
nand U3385 (N_3385,In_2373,In_483);
nand U3386 (N_3386,In_681,In_2459);
xnor U3387 (N_3387,In_1501,In_974);
nor U3388 (N_3388,In_527,In_99);
xor U3389 (N_3389,In_697,In_681);
or U3390 (N_3390,In_95,In_626);
and U3391 (N_3391,In_564,In_88);
or U3392 (N_3392,In_833,In_728);
and U3393 (N_3393,In_915,In_48);
xnor U3394 (N_3394,In_34,In_1908);
and U3395 (N_3395,In_200,In_1609);
or U3396 (N_3396,In_2252,In_1175);
or U3397 (N_3397,In_1726,In_715);
nor U3398 (N_3398,In_152,In_1283);
and U3399 (N_3399,In_834,In_1197);
xor U3400 (N_3400,In_645,In_648);
xor U3401 (N_3401,In_924,In_573);
xnor U3402 (N_3402,In_235,In_1660);
xor U3403 (N_3403,In_233,In_2037);
or U3404 (N_3404,In_1391,In_1445);
nor U3405 (N_3405,In_2120,In_635);
xor U3406 (N_3406,In_2247,In_1407);
xnor U3407 (N_3407,In_470,In_2016);
nand U3408 (N_3408,In_60,In_770);
or U3409 (N_3409,In_1625,In_2155);
nand U3410 (N_3410,In_516,In_1861);
nand U3411 (N_3411,In_1416,In_2311);
nor U3412 (N_3412,In_1894,In_770);
nand U3413 (N_3413,In_729,In_792);
nand U3414 (N_3414,In_192,In_2251);
nand U3415 (N_3415,In_347,In_2401);
and U3416 (N_3416,In_2254,In_1941);
and U3417 (N_3417,In_541,In_1448);
xor U3418 (N_3418,In_1003,In_776);
xnor U3419 (N_3419,In_281,In_210);
or U3420 (N_3420,In_477,In_1487);
or U3421 (N_3421,In_677,In_601);
xnor U3422 (N_3422,In_239,In_2200);
nor U3423 (N_3423,In_1494,In_647);
and U3424 (N_3424,In_1862,In_1680);
xor U3425 (N_3425,In_1602,In_1735);
nor U3426 (N_3426,In_2441,In_1534);
nand U3427 (N_3427,In_2265,In_53);
xnor U3428 (N_3428,In_986,In_798);
or U3429 (N_3429,In_2001,In_2195);
nand U3430 (N_3430,In_1267,In_2161);
xnor U3431 (N_3431,In_1579,In_975);
or U3432 (N_3432,In_574,In_2239);
nand U3433 (N_3433,In_1175,In_439);
and U3434 (N_3434,In_2227,In_590);
or U3435 (N_3435,In_948,In_77);
or U3436 (N_3436,In_2488,In_1524);
nand U3437 (N_3437,In_101,In_1724);
nand U3438 (N_3438,In_1890,In_628);
and U3439 (N_3439,In_480,In_1413);
nand U3440 (N_3440,In_44,In_2320);
xor U3441 (N_3441,In_1641,In_2001);
or U3442 (N_3442,In_2401,In_1397);
xor U3443 (N_3443,In_1750,In_781);
or U3444 (N_3444,In_64,In_1792);
xnor U3445 (N_3445,In_2111,In_1992);
and U3446 (N_3446,In_1816,In_288);
nand U3447 (N_3447,In_1047,In_1272);
and U3448 (N_3448,In_304,In_854);
xor U3449 (N_3449,In_157,In_1069);
or U3450 (N_3450,In_1757,In_1210);
xor U3451 (N_3451,In_2135,In_1806);
and U3452 (N_3452,In_1167,In_1118);
nor U3453 (N_3453,In_737,In_1826);
xnor U3454 (N_3454,In_667,In_200);
nor U3455 (N_3455,In_1382,In_2446);
xnor U3456 (N_3456,In_1624,In_1486);
nand U3457 (N_3457,In_769,In_183);
or U3458 (N_3458,In_762,In_2281);
nor U3459 (N_3459,In_1679,In_310);
nor U3460 (N_3460,In_1315,In_1394);
nand U3461 (N_3461,In_2219,In_406);
nand U3462 (N_3462,In_727,In_974);
nand U3463 (N_3463,In_1213,In_1501);
xnor U3464 (N_3464,In_423,In_271);
nand U3465 (N_3465,In_2362,In_1327);
or U3466 (N_3466,In_846,In_1982);
nand U3467 (N_3467,In_516,In_1358);
xnor U3468 (N_3468,In_455,In_1674);
xor U3469 (N_3469,In_1786,In_971);
and U3470 (N_3470,In_1775,In_1546);
and U3471 (N_3471,In_905,In_9);
nor U3472 (N_3472,In_2282,In_577);
nor U3473 (N_3473,In_480,In_1261);
or U3474 (N_3474,In_2222,In_1972);
and U3475 (N_3475,In_817,In_533);
nand U3476 (N_3476,In_1509,In_1390);
nand U3477 (N_3477,In_1462,In_588);
nand U3478 (N_3478,In_2202,In_1868);
or U3479 (N_3479,In_854,In_2438);
xor U3480 (N_3480,In_1544,In_1392);
and U3481 (N_3481,In_329,In_97);
or U3482 (N_3482,In_2201,In_1266);
nor U3483 (N_3483,In_459,In_631);
xnor U3484 (N_3484,In_483,In_1406);
nor U3485 (N_3485,In_666,In_1684);
xor U3486 (N_3486,In_725,In_1287);
nand U3487 (N_3487,In_1761,In_1327);
nor U3488 (N_3488,In_2321,In_402);
and U3489 (N_3489,In_2157,In_660);
nor U3490 (N_3490,In_2473,In_1247);
or U3491 (N_3491,In_2481,In_1048);
xnor U3492 (N_3492,In_577,In_1494);
or U3493 (N_3493,In_377,In_50);
nand U3494 (N_3494,In_2264,In_2014);
or U3495 (N_3495,In_1398,In_1059);
or U3496 (N_3496,In_1471,In_49);
nor U3497 (N_3497,In_1137,In_1059);
nor U3498 (N_3498,In_4,In_2027);
and U3499 (N_3499,In_566,In_646);
xnor U3500 (N_3500,In_908,In_1592);
nand U3501 (N_3501,In_1026,In_1231);
nand U3502 (N_3502,In_133,In_461);
nor U3503 (N_3503,In_1168,In_1146);
nor U3504 (N_3504,In_2041,In_832);
nor U3505 (N_3505,In_197,In_1337);
nor U3506 (N_3506,In_737,In_200);
or U3507 (N_3507,In_1423,In_2291);
nor U3508 (N_3508,In_998,In_1307);
nor U3509 (N_3509,In_1812,In_1023);
or U3510 (N_3510,In_324,In_1856);
or U3511 (N_3511,In_1397,In_249);
or U3512 (N_3512,In_1053,In_1278);
and U3513 (N_3513,In_128,In_2124);
xor U3514 (N_3514,In_1640,In_844);
and U3515 (N_3515,In_2402,In_1909);
xnor U3516 (N_3516,In_843,In_124);
and U3517 (N_3517,In_2381,In_1525);
nand U3518 (N_3518,In_2354,In_1739);
and U3519 (N_3519,In_892,In_709);
nand U3520 (N_3520,In_1951,In_1327);
and U3521 (N_3521,In_1575,In_354);
nand U3522 (N_3522,In_1858,In_2220);
and U3523 (N_3523,In_477,In_64);
or U3524 (N_3524,In_2157,In_2145);
xnor U3525 (N_3525,In_2365,In_1470);
nor U3526 (N_3526,In_1611,In_1915);
xor U3527 (N_3527,In_331,In_1418);
or U3528 (N_3528,In_420,In_1686);
and U3529 (N_3529,In_694,In_274);
and U3530 (N_3530,In_1228,In_1382);
or U3531 (N_3531,In_1563,In_2458);
and U3532 (N_3532,In_614,In_2434);
xnor U3533 (N_3533,In_1330,In_1502);
or U3534 (N_3534,In_1730,In_1913);
nand U3535 (N_3535,In_1112,In_2266);
or U3536 (N_3536,In_1470,In_207);
xnor U3537 (N_3537,In_1838,In_258);
nor U3538 (N_3538,In_1086,In_2174);
and U3539 (N_3539,In_1862,In_1697);
or U3540 (N_3540,In_1035,In_460);
nor U3541 (N_3541,In_2274,In_2075);
nor U3542 (N_3542,In_2293,In_1423);
or U3543 (N_3543,In_1772,In_78);
or U3544 (N_3544,In_857,In_110);
and U3545 (N_3545,In_503,In_1293);
nor U3546 (N_3546,In_1320,In_1174);
xnor U3547 (N_3547,In_2232,In_2247);
or U3548 (N_3548,In_1531,In_1256);
xnor U3549 (N_3549,In_168,In_1254);
xor U3550 (N_3550,In_26,In_2262);
and U3551 (N_3551,In_2206,In_32);
and U3552 (N_3552,In_2121,In_2014);
nor U3553 (N_3553,In_716,In_1244);
nand U3554 (N_3554,In_52,In_2433);
or U3555 (N_3555,In_1740,In_1079);
or U3556 (N_3556,In_109,In_1136);
nand U3557 (N_3557,In_726,In_2473);
and U3558 (N_3558,In_214,In_1799);
nand U3559 (N_3559,In_890,In_100);
xnor U3560 (N_3560,In_735,In_2033);
nand U3561 (N_3561,In_2340,In_2466);
or U3562 (N_3562,In_288,In_736);
nor U3563 (N_3563,In_1299,In_745);
nor U3564 (N_3564,In_554,In_2133);
or U3565 (N_3565,In_2118,In_1902);
and U3566 (N_3566,In_1151,In_2004);
or U3567 (N_3567,In_36,In_2288);
nor U3568 (N_3568,In_1494,In_140);
or U3569 (N_3569,In_1843,In_27);
xor U3570 (N_3570,In_1671,In_377);
nand U3571 (N_3571,In_732,In_233);
or U3572 (N_3572,In_29,In_1645);
or U3573 (N_3573,In_1252,In_1839);
xor U3574 (N_3574,In_289,In_1468);
nor U3575 (N_3575,In_887,In_91);
nand U3576 (N_3576,In_22,In_1989);
nand U3577 (N_3577,In_1589,In_1058);
nand U3578 (N_3578,In_1160,In_1355);
or U3579 (N_3579,In_1988,In_543);
nand U3580 (N_3580,In_2277,In_1073);
nor U3581 (N_3581,In_1654,In_600);
or U3582 (N_3582,In_1541,In_551);
nor U3583 (N_3583,In_1973,In_2302);
xor U3584 (N_3584,In_726,In_269);
and U3585 (N_3585,In_38,In_2021);
or U3586 (N_3586,In_1409,In_290);
and U3587 (N_3587,In_1668,In_1747);
nor U3588 (N_3588,In_141,In_1885);
nor U3589 (N_3589,In_1898,In_1);
nor U3590 (N_3590,In_1828,In_2113);
and U3591 (N_3591,In_277,In_330);
or U3592 (N_3592,In_1012,In_308);
nor U3593 (N_3593,In_1052,In_1530);
xnor U3594 (N_3594,In_2331,In_2137);
xor U3595 (N_3595,In_1358,In_1851);
nor U3596 (N_3596,In_1410,In_810);
xnor U3597 (N_3597,In_2053,In_553);
xor U3598 (N_3598,In_1326,In_49);
or U3599 (N_3599,In_524,In_174);
or U3600 (N_3600,In_14,In_1968);
or U3601 (N_3601,In_178,In_600);
xnor U3602 (N_3602,In_1533,In_1628);
or U3603 (N_3603,In_48,In_671);
or U3604 (N_3604,In_567,In_1937);
nand U3605 (N_3605,In_1160,In_241);
xnor U3606 (N_3606,In_429,In_2250);
or U3607 (N_3607,In_1826,In_571);
or U3608 (N_3608,In_452,In_370);
and U3609 (N_3609,In_1075,In_785);
nand U3610 (N_3610,In_150,In_107);
nor U3611 (N_3611,In_178,In_2179);
xnor U3612 (N_3612,In_1477,In_1833);
xor U3613 (N_3613,In_280,In_152);
nor U3614 (N_3614,In_133,In_1542);
and U3615 (N_3615,In_2168,In_350);
nand U3616 (N_3616,In_889,In_1512);
nand U3617 (N_3617,In_497,In_1331);
or U3618 (N_3618,In_960,In_716);
xnor U3619 (N_3619,In_2303,In_1085);
or U3620 (N_3620,In_507,In_390);
nand U3621 (N_3621,In_1669,In_1752);
xnor U3622 (N_3622,In_2203,In_1749);
and U3623 (N_3623,In_136,In_1732);
nand U3624 (N_3624,In_753,In_97);
nand U3625 (N_3625,In_2477,In_1029);
nor U3626 (N_3626,In_101,In_2293);
nor U3627 (N_3627,In_2127,In_976);
and U3628 (N_3628,In_914,In_1056);
nand U3629 (N_3629,In_1309,In_2419);
nand U3630 (N_3630,In_1558,In_1322);
nand U3631 (N_3631,In_2100,In_1074);
xnor U3632 (N_3632,In_149,In_1804);
nor U3633 (N_3633,In_904,In_75);
nor U3634 (N_3634,In_1162,In_11);
or U3635 (N_3635,In_1402,In_1265);
nor U3636 (N_3636,In_2403,In_385);
nand U3637 (N_3637,In_1199,In_2092);
or U3638 (N_3638,In_2494,In_1582);
nand U3639 (N_3639,In_283,In_2054);
and U3640 (N_3640,In_1401,In_1758);
or U3641 (N_3641,In_591,In_2188);
and U3642 (N_3642,In_2291,In_2262);
nand U3643 (N_3643,In_831,In_2476);
xnor U3644 (N_3644,In_495,In_1318);
and U3645 (N_3645,In_1544,In_1453);
xnor U3646 (N_3646,In_1277,In_1088);
nand U3647 (N_3647,In_2152,In_1310);
and U3648 (N_3648,In_2323,In_1909);
or U3649 (N_3649,In_374,In_1274);
xnor U3650 (N_3650,In_1932,In_1968);
nand U3651 (N_3651,In_966,In_1561);
nor U3652 (N_3652,In_1395,In_1449);
nor U3653 (N_3653,In_1213,In_463);
xor U3654 (N_3654,In_1214,In_2180);
xor U3655 (N_3655,In_2434,In_949);
nor U3656 (N_3656,In_2270,In_945);
and U3657 (N_3657,In_506,In_1705);
and U3658 (N_3658,In_991,In_1841);
or U3659 (N_3659,In_411,In_2101);
or U3660 (N_3660,In_2249,In_301);
nor U3661 (N_3661,In_2173,In_978);
and U3662 (N_3662,In_584,In_958);
nand U3663 (N_3663,In_2228,In_2261);
nand U3664 (N_3664,In_1712,In_352);
and U3665 (N_3665,In_863,In_424);
and U3666 (N_3666,In_8,In_1567);
nor U3667 (N_3667,In_542,In_165);
xor U3668 (N_3668,In_2448,In_1559);
or U3669 (N_3669,In_1589,In_1525);
nand U3670 (N_3670,In_600,In_2238);
nand U3671 (N_3671,In_115,In_1954);
and U3672 (N_3672,In_471,In_8);
xnor U3673 (N_3673,In_1258,In_570);
or U3674 (N_3674,In_2364,In_1458);
xor U3675 (N_3675,In_1268,In_268);
nor U3676 (N_3676,In_133,In_217);
and U3677 (N_3677,In_1520,In_392);
or U3678 (N_3678,In_1266,In_745);
or U3679 (N_3679,In_271,In_1017);
or U3680 (N_3680,In_82,In_434);
and U3681 (N_3681,In_1794,In_432);
xor U3682 (N_3682,In_2260,In_959);
and U3683 (N_3683,In_1332,In_1742);
nor U3684 (N_3684,In_840,In_2147);
nand U3685 (N_3685,In_1968,In_813);
nor U3686 (N_3686,In_41,In_2367);
nor U3687 (N_3687,In_387,In_305);
and U3688 (N_3688,In_2170,In_790);
xnor U3689 (N_3689,In_232,In_86);
or U3690 (N_3690,In_1850,In_1970);
or U3691 (N_3691,In_96,In_428);
and U3692 (N_3692,In_2204,In_1971);
or U3693 (N_3693,In_645,In_535);
and U3694 (N_3694,In_2388,In_1828);
or U3695 (N_3695,In_457,In_1834);
nand U3696 (N_3696,In_2089,In_1066);
nor U3697 (N_3697,In_1653,In_19);
nor U3698 (N_3698,In_1543,In_122);
and U3699 (N_3699,In_97,In_2424);
and U3700 (N_3700,In_411,In_630);
and U3701 (N_3701,In_1296,In_1265);
and U3702 (N_3702,In_1162,In_2217);
and U3703 (N_3703,In_1680,In_1442);
nand U3704 (N_3704,In_276,In_2275);
xnor U3705 (N_3705,In_1800,In_1039);
nor U3706 (N_3706,In_996,In_1239);
and U3707 (N_3707,In_125,In_2437);
nor U3708 (N_3708,In_2316,In_799);
xnor U3709 (N_3709,In_1033,In_1281);
nand U3710 (N_3710,In_199,In_1829);
nand U3711 (N_3711,In_980,In_1446);
nand U3712 (N_3712,In_2115,In_53);
nor U3713 (N_3713,In_412,In_2462);
nand U3714 (N_3714,In_1505,In_1326);
xnor U3715 (N_3715,In_60,In_556);
and U3716 (N_3716,In_171,In_571);
nor U3717 (N_3717,In_2084,In_1189);
nand U3718 (N_3718,In_1875,In_1463);
nand U3719 (N_3719,In_733,In_357);
nor U3720 (N_3720,In_583,In_1342);
and U3721 (N_3721,In_1905,In_506);
nor U3722 (N_3722,In_458,In_2086);
xnor U3723 (N_3723,In_1467,In_1614);
and U3724 (N_3724,In_1977,In_2015);
or U3725 (N_3725,In_2456,In_1279);
xnor U3726 (N_3726,In_690,In_1889);
and U3727 (N_3727,In_1031,In_850);
and U3728 (N_3728,In_873,In_1470);
nor U3729 (N_3729,In_818,In_1118);
or U3730 (N_3730,In_2316,In_1189);
xnor U3731 (N_3731,In_1752,In_13);
nor U3732 (N_3732,In_1624,In_1032);
nand U3733 (N_3733,In_1177,In_964);
nand U3734 (N_3734,In_1020,In_2449);
or U3735 (N_3735,In_1561,In_1417);
nor U3736 (N_3736,In_2106,In_2068);
nand U3737 (N_3737,In_970,In_884);
nor U3738 (N_3738,In_30,In_1593);
or U3739 (N_3739,In_2193,In_1218);
or U3740 (N_3740,In_2202,In_1241);
and U3741 (N_3741,In_1919,In_1337);
xor U3742 (N_3742,In_2196,In_299);
nand U3743 (N_3743,In_804,In_2096);
xnor U3744 (N_3744,In_1566,In_1319);
xnor U3745 (N_3745,In_511,In_1235);
xor U3746 (N_3746,In_2121,In_57);
xor U3747 (N_3747,In_491,In_525);
xnor U3748 (N_3748,In_700,In_2392);
or U3749 (N_3749,In_11,In_1795);
nor U3750 (N_3750,In_345,In_947);
nor U3751 (N_3751,In_651,In_654);
or U3752 (N_3752,In_1117,In_805);
nor U3753 (N_3753,In_103,In_1017);
xnor U3754 (N_3754,In_317,In_810);
or U3755 (N_3755,In_938,In_277);
or U3756 (N_3756,In_1375,In_1658);
xnor U3757 (N_3757,In_245,In_159);
and U3758 (N_3758,In_248,In_1994);
or U3759 (N_3759,In_1283,In_2135);
or U3760 (N_3760,In_1828,In_2166);
or U3761 (N_3761,In_1914,In_2322);
and U3762 (N_3762,In_621,In_102);
or U3763 (N_3763,In_110,In_1930);
nor U3764 (N_3764,In_1589,In_517);
or U3765 (N_3765,In_1659,In_183);
nand U3766 (N_3766,In_117,In_2411);
nor U3767 (N_3767,In_662,In_330);
nand U3768 (N_3768,In_1180,In_2480);
nand U3769 (N_3769,In_1675,In_361);
xnor U3770 (N_3770,In_991,In_1306);
or U3771 (N_3771,In_1349,In_1009);
or U3772 (N_3772,In_166,In_2309);
or U3773 (N_3773,In_2424,In_1601);
or U3774 (N_3774,In_463,In_2128);
and U3775 (N_3775,In_499,In_2408);
and U3776 (N_3776,In_2128,In_724);
or U3777 (N_3777,In_504,In_1721);
xnor U3778 (N_3778,In_468,In_1106);
and U3779 (N_3779,In_1444,In_2251);
or U3780 (N_3780,In_2173,In_1468);
nor U3781 (N_3781,In_50,In_2034);
xor U3782 (N_3782,In_33,In_1356);
nor U3783 (N_3783,In_1917,In_1960);
or U3784 (N_3784,In_747,In_4);
nor U3785 (N_3785,In_153,In_1293);
nand U3786 (N_3786,In_2276,In_824);
or U3787 (N_3787,In_35,In_1102);
xor U3788 (N_3788,In_2318,In_579);
and U3789 (N_3789,In_210,In_833);
nor U3790 (N_3790,In_233,In_707);
nor U3791 (N_3791,In_130,In_962);
and U3792 (N_3792,In_679,In_1519);
or U3793 (N_3793,In_127,In_1167);
nor U3794 (N_3794,In_176,In_1536);
or U3795 (N_3795,In_1171,In_1489);
and U3796 (N_3796,In_91,In_844);
nand U3797 (N_3797,In_1551,In_1121);
or U3798 (N_3798,In_2324,In_1405);
nand U3799 (N_3799,In_1481,In_468);
xor U3800 (N_3800,In_454,In_2198);
nand U3801 (N_3801,In_267,In_185);
nand U3802 (N_3802,In_1450,In_1508);
xor U3803 (N_3803,In_1710,In_1192);
or U3804 (N_3804,In_888,In_96);
and U3805 (N_3805,In_785,In_2014);
xor U3806 (N_3806,In_1690,In_493);
and U3807 (N_3807,In_2316,In_1054);
nor U3808 (N_3808,In_2116,In_1676);
nand U3809 (N_3809,In_1935,In_2194);
xor U3810 (N_3810,In_2074,In_1938);
nor U3811 (N_3811,In_386,In_1357);
or U3812 (N_3812,In_26,In_1309);
and U3813 (N_3813,In_2282,In_22);
or U3814 (N_3814,In_1129,In_431);
nor U3815 (N_3815,In_1028,In_2204);
xnor U3816 (N_3816,In_1165,In_1898);
and U3817 (N_3817,In_1736,In_1151);
xor U3818 (N_3818,In_18,In_2190);
and U3819 (N_3819,In_1897,In_104);
nor U3820 (N_3820,In_1511,In_153);
nand U3821 (N_3821,In_1956,In_1591);
and U3822 (N_3822,In_519,In_474);
xor U3823 (N_3823,In_2402,In_1773);
and U3824 (N_3824,In_1793,In_696);
or U3825 (N_3825,In_1306,In_873);
and U3826 (N_3826,In_1260,In_1511);
nand U3827 (N_3827,In_1860,In_2084);
nor U3828 (N_3828,In_2280,In_1953);
and U3829 (N_3829,In_1483,In_1882);
or U3830 (N_3830,In_2294,In_459);
and U3831 (N_3831,In_2062,In_2180);
nor U3832 (N_3832,In_1747,In_238);
xor U3833 (N_3833,In_2195,In_2172);
nor U3834 (N_3834,In_696,In_2479);
and U3835 (N_3835,In_1084,In_285);
nor U3836 (N_3836,In_1088,In_2171);
and U3837 (N_3837,In_30,In_1299);
nand U3838 (N_3838,In_1120,In_1997);
and U3839 (N_3839,In_1691,In_1519);
or U3840 (N_3840,In_400,In_15);
nor U3841 (N_3841,In_773,In_11);
nor U3842 (N_3842,In_1594,In_1754);
or U3843 (N_3843,In_409,In_886);
and U3844 (N_3844,In_1055,In_1137);
nand U3845 (N_3845,In_227,In_1821);
or U3846 (N_3846,In_556,In_2261);
and U3847 (N_3847,In_2390,In_1100);
xor U3848 (N_3848,In_1958,In_1629);
and U3849 (N_3849,In_347,In_436);
and U3850 (N_3850,In_1998,In_1380);
and U3851 (N_3851,In_1475,In_969);
nor U3852 (N_3852,In_1743,In_2063);
and U3853 (N_3853,In_183,In_1873);
or U3854 (N_3854,In_1859,In_774);
xor U3855 (N_3855,In_1798,In_1285);
and U3856 (N_3856,In_202,In_1516);
nor U3857 (N_3857,In_808,In_1025);
xor U3858 (N_3858,In_9,In_266);
nor U3859 (N_3859,In_1465,In_1675);
nor U3860 (N_3860,In_1593,In_1800);
or U3861 (N_3861,In_1396,In_1321);
nor U3862 (N_3862,In_1765,In_1950);
nor U3863 (N_3863,In_2271,In_42);
xor U3864 (N_3864,In_1314,In_1161);
or U3865 (N_3865,In_30,In_1381);
xor U3866 (N_3866,In_629,In_79);
nor U3867 (N_3867,In_89,In_675);
nand U3868 (N_3868,In_1504,In_316);
and U3869 (N_3869,In_240,In_2428);
nor U3870 (N_3870,In_380,In_126);
or U3871 (N_3871,In_1344,In_2446);
and U3872 (N_3872,In_934,In_596);
nand U3873 (N_3873,In_1633,In_1153);
nand U3874 (N_3874,In_1554,In_2336);
nor U3875 (N_3875,In_1276,In_1912);
or U3876 (N_3876,In_2376,In_1536);
nand U3877 (N_3877,In_1215,In_1827);
xnor U3878 (N_3878,In_2086,In_0);
xnor U3879 (N_3879,In_900,In_1371);
nand U3880 (N_3880,In_966,In_1964);
xnor U3881 (N_3881,In_1919,In_727);
xnor U3882 (N_3882,In_631,In_126);
or U3883 (N_3883,In_140,In_2475);
nand U3884 (N_3884,In_552,In_324);
xnor U3885 (N_3885,In_246,In_1562);
xnor U3886 (N_3886,In_1002,In_242);
and U3887 (N_3887,In_2429,In_2402);
or U3888 (N_3888,In_52,In_2000);
nor U3889 (N_3889,In_242,In_2184);
or U3890 (N_3890,In_261,In_1898);
or U3891 (N_3891,In_591,In_1386);
xnor U3892 (N_3892,In_2455,In_1817);
or U3893 (N_3893,In_566,In_2071);
nor U3894 (N_3894,In_2007,In_2418);
nor U3895 (N_3895,In_2262,In_1186);
nor U3896 (N_3896,In_992,In_770);
and U3897 (N_3897,In_1313,In_357);
nor U3898 (N_3898,In_350,In_432);
xnor U3899 (N_3899,In_1144,In_572);
and U3900 (N_3900,In_426,In_129);
xor U3901 (N_3901,In_942,In_970);
nor U3902 (N_3902,In_1725,In_2054);
nand U3903 (N_3903,In_557,In_2118);
and U3904 (N_3904,In_1635,In_586);
or U3905 (N_3905,In_349,In_220);
nor U3906 (N_3906,In_1710,In_1440);
xnor U3907 (N_3907,In_741,In_425);
or U3908 (N_3908,In_2181,In_1303);
and U3909 (N_3909,In_732,In_1474);
xor U3910 (N_3910,In_786,In_5);
or U3911 (N_3911,In_1534,In_1230);
or U3912 (N_3912,In_1480,In_1582);
nand U3913 (N_3913,In_2082,In_2133);
nand U3914 (N_3914,In_2493,In_734);
nor U3915 (N_3915,In_2094,In_1116);
or U3916 (N_3916,In_1779,In_2399);
or U3917 (N_3917,In_286,In_1247);
nor U3918 (N_3918,In_1886,In_1459);
nand U3919 (N_3919,In_1501,In_1002);
or U3920 (N_3920,In_1179,In_482);
xnor U3921 (N_3921,In_2469,In_134);
and U3922 (N_3922,In_289,In_1734);
nor U3923 (N_3923,In_513,In_1293);
and U3924 (N_3924,In_2378,In_275);
nor U3925 (N_3925,In_909,In_2361);
and U3926 (N_3926,In_1369,In_543);
xor U3927 (N_3927,In_2001,In_2015);
nor U3928 (N_3928,In_1345,In_1639);
nor U3929 (N_3929,In_1462,In_175);
nor U3930 (N_3930,In_408,In_1302);
or U3931 (N_3931,In_1552,In_2448);
nand U3932 (N_3932,In_943,In_2237);
or U3933 (N_3933,In_1173,In_2289);
and U3934 (N_3934,In_972,In_2274);
xor U3935 (N_3935,In_1262,In_1310);
or U3936 (N_3936,In_2226,In_1538);
xnor U3937 (N_3937,In_748,In_1032);
and U3938 (N_3938,In_2108,In_1744);
and U3939 (N_3939,In_1074,In_1836);
or U3940 (N_3940,In_1794,In_638);
and U3941 (N_3941,In_1969,In_1598);
and U3942 (N_3942,In_251,In_457);
xnor U3943 (N_3943,In_1137,In_2399);
nor U3944 (N_3944,In_1137,In_2122);
xor U3945 (N_3945,In_1822,In_2209);
nand U3946 (N_3946,In_2106,In_1210);
and U3947 (N_3947,In_708,In_243);
nand U3948 (N_3948,In_440,In_1585);
or U3949 (N_3949,In_746,In_1862);
xor U3950 (N_3950,In_682,In_2401);
or U3951 (N_3951,In_532,In_946);
xor U3952 (N_3952,In_532,In_1535);
or U3953 (N_3953,In_2364,In_410);
xnor U3954 (N_3954,In_2414,In_751);
nand U3955 (N_3955,In_2077,In_298);
or U3956 (N_3956,In_1618,In_2356);
and U3957 (N_3957,In_1582,In_1344);
xnor U3958 (N_3958,In_1505,In_174);
xnor U3959 (N_3959,In_2012,In_1933);
xor U3960 (N_3960,In_1344,In_1782);
and U3961 (N_3961,In_2290,In_1287);
or U3962 (N_3962,In_589,In_1833);
nor U3963 (N_3963,In_1468,In_2480);
and U3964 (N_3964,In_1422,In_1402);
and U3965 (N_3965,In_1507,In_436);
xor U3966 (N_3966,In_1937,In_560);
nor U3967 (N_3967,In_1216,In_591);
nand U3968 (N_3968,In_1641,In_950);
nand U3969 (N_3969,In_1801,In_2476);
xnor U3970 (N_3970,In_897,In_403);
and U3971 (N_3971,In_1735,In_1301);
nor U3972 (N_3972,In_386,In_883);
xor U3973 (N_3973,In_874,In_376);
and U3974 (N_3974,In_1028,In_1220);
xnor U3975 (N_3975,In_2387,In_1691);
or U3976 (N_3976,In_1207,In_411);
nand U3977 (N_3977,In_478,In_2222);
nor U3978 (N_3978,In_662,In_440);
nand U3979 (N_3979,In_1957,In_2242);
nand U3980 (N_3980,In_2409,In_947);
xnor U3981 (N_3981,In_2162,In_433);
xor U3982 (N_3982,In_2455,In_977);
nor U3983 (N_3983,In_272,In_2206);
xnor U3984 (N_3984,In_1880,In_152);
nand U3985 (N_3985,In_1673,In_1141);
and U3986 (N_3986,In_230,In_2220);
or U3987 (N_3987,In_116,In_1895);
or U3988 (N_3988,In_1921,In_1711);
and U3989 (N_3989,In_595,In_1358);
nand U3990 (N_3990,In_1218,In_1758);
or U3991 (N_3991,In_285,In_986);
and U3992 (N_3992,In_213,In_1431);
nand U3993 (N_3993,In_1911,In_926);
nor U3994 (N_3994,In_195,In_2485);
or U3995 (N_3995,In_904,In_1224);
and U3996 (N_3996,In_699,In_1094);
or U3997 (N_3997,In_1683,In_1912);
nand U3998 (N_3998,In_256,In_2448);
nand U3999 (N_3999,In_2313,In_2029);
nor U4000 (N_4000,In_1712,In_2055);
and U4001 (N_4001,In_1325,In_0);
xor U4002 (N_4002,In_606,In_2393);
or U4003 (N_4003,In_221,In_1232);
and U4004 (N_4004,In_2361,In_201);
and U4005 (N_4005,In_475,In_527);
xnor U4006 (N_4006,In_1192,In_514);
nor U4007 (N_4007,In_113,In_963);
and U4008 (N_4008,In_617,In_1464);
nand U4009 (N_4009,In_308,In_1864);
xor U4010 (N_4010,In_2112,In_336);
nand U4011 (N_4011,In_1539,In_1643);
xnor U4012 (N_4012,In_2288,In_2271);
or U4013 (N_4013,In_2200,In_2096);
and U4014 (N_4014,In_1715,In_541);
nand U4015 (N_4015,In_683,In_789);
nand U4016 (N_4016,In_2236,In_751);
nand U4017 (N_4017,In_1373,In_1282);
nor U4018 (N_4018,In_2202,In_253);
xnor U4019 (N_4019,In_2464,In_2407);
nand U4020 (N_4020,In_1758,In_2407);
xnor U4021 (N_4021,In_1527,In_212);
and U4022 (N_4022,In_2301,In_952);
nand U4023 (N_4023,In_301,In_1970);
xnor U4024 (N_4024,In_1278,In_1670);
nand U4025 (N_4025,In_364,In_1004);
nand U4026 (N_4026,In_788,In_1175);
xor U4027 (N_4027,In_828,In_1490);
nor U4028 (N_4028,In_2205,In_572);
and U4029 (N_4029,In_2168,In_145);
nor U4030 (N_4030,In_1891,In_1548);
xnor U4031 (N_4031,In_2232,In_448);
nor U4032 (N_4032,In_2368,In_516);
and U4033 (N_4033,In_1458,In_391);
xor U4034 (N_4034,In_1464,In_1923);
nand U4035 (N_4035,In_184,In_643);
or U4036 (N_4036,In_382,In_1943);
xnor U4037 (N_4037,In_1149,In_262);
xor U4038 (N_4038,In_2104,In_2342);
nor U4039 (N_4039,In_519,In_423);
xnor U4040 (N_4040,In_1713,In_1732);
nand U4041 (N_4041,In_868,In_2101);
nand U4042 (N_4042,In_77,In_1084);
nand U4043 (N_4043,In_458,In_1987);
xor U4044 (N_4044,In_264,In_2276);
xor U4045 (N_4045,In_1906,In_1454);
xor U4046 (N_4046,In_2116,In_1389);
xor U4047 (N_4047,In_57,In_1245);
or U4048 (N_4048,In_438,In_2327);
xor U4049 (N_4049,In_1395,In_1909);
and U4050 (N_4050,In_835,In_2342);
nand U4051 (N_4051,In_1503,In_1525);
and U4052 (N_4052,In_223,In_649);
xnor U4053 (N_4053,In_2261,In_78);
or U4054 (N_4054,In_325,In_919);
and U4055 (N_4055,In_276,In_2483);
and U4056 (N_4056,In_723,In_2067);
nor U4057 (N_4057,In_53,In_1752);
and U4058 (N_4058,In_612,In_801);
nand U4059 (N_4059,In_2428,In_1257);
or U4060 (N_4060,In_1455,In_1773);
or U4061 (N_4061,In_1090,In_2462);
or U4062 (N_4062,In_1813,In_1258);
xnor U4063 (N_4063,In_1467,In_521);
and U4064 (N_4064,In_202,In_216);
nor U4065 (N_4065,In_2404,In_1561);
and U4066 (N_4066,In_1373,In_370);
and U4067 (N_4067,In_835,In_2307);
nor U4068 (N_4068,In_1074,In_541);
nor U4069 (N_4069,In_1065,In_2288);
nand U4070 (N_4070,In_1733,In_1719);
or U4071 (N_4071,In_439,In_2227);
or U4072 (N_4072,In_954,In_1114);
or U4073 (N_4073,In_522,In_1174);
nor U4074 (N_4074,In_205,In_1417);
nor U4075 (N_4075,In_1222,In_278);
nor U4076 (N_4076,In_2115,In_326);
nand U4077 (N_4077,In_1168,In_2094);
nand U4078 (N_4078,In_2365,In_1834);
and U4079 (N_4079,In_1956,In_2303);
xnor U4080 (N_4080,In_214,In_2256);
nor U4081 (N_4081,In_826,In_831);
nand U4082 (N_4082,In_2096,In_114);
nor U4083 (N_4083,In_2009,In_2342);
nor U4084 (N_4084,In_1886,In_1676);
and U4085 (N_4085,In_391,In_8);
nand U4086 (N_4086,In_445,In_1836);
or U4087 (N_4087,In_888,In_636);
nand U4088 (N_4088,In_2465,In_333);
nor U4089 (N_4089,In_1088,In_1865);
nand U4090 (N_4090,In_528,In_1445);
or U4091 (N_4091,In_171,In_1013);
or U4092 (N_4092,In_907,In_1372);
or U4093 (N_4093,In_465,In_1659);
xor U4094 (N_4094,In_2041,In_1465);
or U4095 (N_4095,In_1355,In_1006);
xnor U4096 (N_4096,In_913,In_1202);
and U4097 (N_4097,In_2350,In_1889);
nand U4098 (N_4098,In_1784,In_2268);
nor U4099 (N_4099,In_2043,In_1487);
nand U4100 (N_4100,In_541,In_2383);
and U4101 (N_4101,In_1738,In_163);
xor U4102 (N_4102,In_1684,In_2355);
nand U4103 (N_4103,In_2288,In_732);
xor U4104 (N_4104,In_1588,In_756);
nand U4105 (N_4105,In_1924,In_1317);
nand U4106 (N_4106,In_1561,In_590);
or U4107 (N_4107,In_1865,In_2410);
xnor U4108 (N_4108,In_124,In_566);
nor U4109 (N_4109,In_2485,In_1967);
nor U4110 (N_4110,In_398,In_1271);
nand U4111 (N_4111,In_2352,In_1740);
nor U4112 (N_4112,In_2182,In_2456);
xnor U4113 (N_4113,In_2344,In_355);
or U4114 (N_4114,In_1357,In_2031);
and U4115 (N_4115,In_530,In_536);
xor U4116 (N_4116,In_229,In_2390);
or U4117 (N_4117,In_1640,In_1199);
nand U4118 (N_4118,In_1995,In_855);
xor U4119 (N_4119,In_700,In_960);
xnor U4120 (N_4120,In_178,In_1308);
nor U4121 (N_4121,In_1433,In_1854);
nor U4122 (N_4122,In_28,In_1903);
nand U4123 (N_4123,In_138,In_1010);
nor U4124 (N_4124,In_251,In_1535);
nand U4125 (N_4125,In_2224,In_486);
nand U4126 (N_4126,In_148,In_1895);
or U4127 (N_4127,In_2134,In_3);
or U4128 (N_4128,In_486,In_522);
nor U4129 (N_4129,In_594,In_1152);
nand U4130 (N_4130,In_108,In_76);
xor U4131 (N_4131,In_2041,In_2191);
or U4132 (N_4132,In_2471,In_2186);
xnor U4133 (N_4133,In_1319,In_1738);
nand U4134 (N_4134,In_765,In_445);
or U4135 (N_4135,In_1110,In_1104);
xnor U4136 (N_4136,In_2493,In_1761);
nor U4137 (N_4137,In_585,In_883);
or U4138 (N_4138,In_267,In_1773);
and U4139 (N_4139,In_1297,In_1482);
nor U4140 (N_4140,In_94,In_2465);
xor U4141 (N_4141,In_1532,In_2444);
or U4142 (N_4142,In_131,In_88);
xnor U4143 (N_4143,In_2204,In_485);
nand U4144 (N_4144,In_2034,In_678);
xnor U4145 (N_4145,In_1166,In_971);
nand U4146 (N_4146,In_1112,In_2218);
xor U4147 (N_4147,In_808,In_1904);
xor U4148 (N_4148,In_673,In_1343);
nor U4149 (N_4149,In_1698,In_174);
or U4150 (N_4150,In_1485,In_219);
nor U4151 (N_4151,In_2191,In_1894);
nand U4152 (N_4152,In_2247,In_604);
xnor U4153 (N_4153,In_1323,In_1141);
xor U4154 (N_4154,In_2053,In_1904);
nand U4155 (N_4155,In_2416,In_62);
nor U4156 (N_4156,In_2134,In_44);
nor U4157 (N_4157,In_161,In_1984);
and U4158 (N_4158,In_1106,In_1751);
nand U4159 (N_4159,In_1534,In_1713);
or U4160 (N_4160,In_1491,In_1956);
nand U4161 (N_4161,In_2262,In_1447);
or U4162 (N_4162,In_963,In_110);
nand U4163 (N_4163,In_656,In_582);
nand U4164 (N_4164,In_1165,In_2462);
xnor U4165 (N_4165,In_1725,In_1067);
nand U4166 (N_4166,In_1297,In_1887);
xnor U4167 (N_4167,In_1403,In_2359);
and U4168 (N_4168,In_1175,In_920);
xnor U4169 (N_4169,In_516,In_2261);
and U4170 (N_4170,In_2161,In_252);
and U4171 (N_4171,In_153,In_383);
nand U4172 (N_4172,In_2234,In_1560);
xor U4173 (N_4173,In_666,In_1387);
or U4174 (N_4174,In_1552,In_2439);
nor U4175 (N_4175,In_282,In_2077);
nand U4176 (N_4176,In_553,In_2043);
and U4177 (N_4177,In_1237,In_989);
and U4178 (N_4178,In_2326,In_1632);
xnor U4179 (N_4179,In_121,In_1196);
and U4180 (N_4180,In_1502,In_1183);
xnor U4181 (N_4181,In_1246,In_715);
and U4182 (N_4182,In_1614,In_93);
nor U4183 (N_4183,In_2397,In_1400);
and U4184 (N_4184,In_2446,In_1762);
nor U4185 (N_4185,In_206,In_1105);
or U4186 (N_4186,In_628,In_724);
and U4187 (N_4187,In_348,In_329);
nand U4188 (N_4188,In_2296,In_926);
nor U4189 (N_4189,In_1209,In_1384);
and U4190 (N_4190,In_133,In_1848);
xnor U4191 (N_4191,In_2277,In_1643);
and U4192 (N_4192,In_2343,In_301);
and U4193 (N_4193,In_1377,In_211);
or U4194 (N_4194,In_1530,In_1851);
and U4195 (N_4195,In_1928,In_2265);
and U4196 (N_4196,In_571,In_829);
nand U4197 (N_4197,In_827,In_1848);
nand U4198 (N_4198,In_893,In_1606);
or U4199 (N_4199,In_2395,In_13);
or U4200 (N_4200,In_246,In_2314);
nand U4201 (N_4201,In_736,In_2246);
or U4202 (N_4202,In_1309,In_1243);
or U4203 (N_4203,In_564,In_1142);
nand U4204 (N_4204,In_1074,In_643);
nor U4205 (N_4205,In_1452,In_269);
and U4206 (N_4206,In_934,In_1210);
nand U4207 (N_4207,In_1364,In_2075);
nor U4208 (N_4208,In_2146,In_2356);
nor U4209 (N_4209,In_1560,In_749);
nor U4210 (N_4210,In_1642,In_597);
and U4211 (N_4211,In_732,In_2289);
xor U4212 (N_4212,In_2420,In_1489);
xor U4213 (N_4213,In_112,In_1696);
xor U4214 (N_4214,In_2420,In_1804);
xor U4215 (N_4215,In_1285,In_516);
nand U4216 (N_4216,In_1517,In_1420);
nand U4217 (N_4217,In_2424,In_2252);
nor U4218 (N_4218,In_2007,In_2170);
xnor U4219 (N_4219,In_1994,In_476);
and U4220 (N_4220,In_924,In_841);
and U4221 (N_4221,In_670,In_2321);
and U4222 (N_4222,In_1337,In_1024);
or U4223 (N_4223,In_1668,In_2089);
or U4224 (N_4224,In_2195,In_5);
nor U4225 (N_4225,In_1534,In_1951);
or U4226 (N_4226,In_1379,In_857);
xnor U4227 (N_4227,In_71,In_1545);
nand U4228 (N_4228,In_421,In_531);
nor U4229 (N_4229,In_1061,In_943);
and U4230 (N_4230,In_2359,In_645);
xnor U4231 (N_4231,In_2177,In_1842);
and U4232 (N_4232,In_272,In_803);
xor U4233 (N_4233,In_1949,In_1547);
nor U4234 (N_4234,In_2028,In_283);
and U4235 (N_4235,In_1224,In_1768);
nor U4236 (N_4236,In_1544,In_874);
and U4237 (N_4237,In_2261,In_1561);
nor U4238 (N_4238,In_2087,In_1865);
xor U4239 (N_4239,In_1397,In_1347);
xor U4240 (N_4240,In_2124,In_2460);
nor U4241 (N_4241,In_2395,In_2186);
or U4242 (N_4242,In_1441,In_2313);
or U4243 (N_4243,In_1328,In_2257);
nand U4244 (N_4244,In_2146,In_2227);
or U4245 (N_4245,In_2298,In_1739);
and U4246 (N_4246,In_798,In_39);
xnor U4247 (N_4247,In_14,In_920);
nor U4248 (N_4248,In_2190,In_520);
or U4249 (N_4249,In_141,In_2355);
and U4250 (N_4250,In_1949,In_580);
nand U4251 (N_4251,In_524,In_2388);
nand U4252 (N_4252,In_1972,In_783);
and U4253 (N_4253,In_19,In_558);
nand U4254 (N_4254,In_1291,In_1223);
or U4255 (N_4255,In_1856,In_52);
nand U4256 (N_4256,In_1829,In_2114);
xor U4257 (N_4257,In_543,In_47);
or U4258 (N_4258,In_1747,In_360);
nor U4259 (N_4259,In_1063,In_306);
xnor U4260 (N_4260,In_1425,In_692);
nand U4261 (N_4261,In_2425,In_2166);
nor U4262 (N_4262,In_867,In_1601);
and U4263 (N_4263,In_1136,In_537);
xor U4264 (N_4264,In_1199,In_281);
nor U4265 (N_4265,In_1724,In_1567);
or U4266 (N_4266,In_2106,In_297);
or U4267 (N_4267,In_1403,In_1575);
or U4268 (N_4268,In_1500,In_1116);
or U4269 (N_4269,In_0,In_2063);
xnor U4270 (N_4270,In_2077,In_1569);
xnor U4271 (N_4271,In_135,In_2324);
or U4272 (N_4272,In_457,In_2067);
and U4273 (N_4273,In_2298,In_2480);
xor U4274 (N_4274,In_838,In_2041);
xnor U4275 (N_4275,In_1901,In_1272);
xnor U4276 (N_4276,In_564,In_1468);
nor U4277 (N_4277,In_1534,In_823);
nand U4278 (N_4278,In_108,In_6);
and U4279 (N_4279,In_1373,In_259);
nor U4280 (N_4280,In_552,In_278);
nand U4281 (N_4281,In_2375,In_1556);
nand U4282 (N_4282,In_1256,In_874);
and U4283 (N_4283,In_1083,In_2376);
or U4284 (N_4284,In_1375,In_791);
or U4285 (N_4285,In_13,In_1298);
or U4286 (N_4286,In_260,In_565);
nor U4287 (N_4287,In_959,In_2310);
or U4288 (N_4288,In_239,In_500);
xnor U4289 (N_4289,In_733,In_1851);
nand U4290 (N_4290,In_2142,In_1411);
xnor U4291 (N_4291,In_1808,In_2259);
and U4292 (N_4292,In_801,In_2486);
nand U4293 (N_4293,In_1613,In_1952);
xor U4294 (N_4294,In_1161,In_1993);
xnor U4295 (N_4295,In_1412,In_2107);
xnor U4296 (N_4296,In_1326,In_1174);
xor U4297 (N_4297,In_360,In_728);
xnor U4298 (N_4298,In_465,In_1100);
and U4299 (N_4299,In_1419,In_2440);
and U4300 (N_4300,In_1228,In_778);
nor U4301 (N_4301,In_1785,In_1578);
or U4302 (N_4302,In_945,In_664);
and U4303 (N_4303,In_1565,In_350);
or U4304 (N_4304,In_1898,In_1416);
nor U4305 (N_4305,In_1704,In_1439);
nor U4306 (N_4306,In_1709,In_2388);
xor U4307 (N_4307,In_1087,In_315);
xnor U4308 (N_4308,In_400,In_1635);
and U4309 (N_4309,In_707,In_308);
and U4310 (N_4310,In_2372,In_388);
or U4311 (N_4311,In_1111,In_532);
and U4312 (N_4312,In_1679,In_130);
nor U4313 (N_4313,In_1926,In_1509);
and U4314 (N_4314,In_205,In_1343);
nor U4315 (N_4315,In_1981,In_1404);
and U4316 (N_4316,In_1754,In_2486);
nand U4317 (N_4317,In_1482,In_1213);
nand U4318 (N_4318,In_1293,In_1308);
nor U4319 (N_4319,In_864,In_1771);
nor U4320 (N_4320,In_253,In_2447);
and U4321 (N_4321,In_1423,In_236);
xor U4322 (N_4322,In_190,In_1709);
xor U4323 (N_4323,In_1790,In_2154);
nor U4324 (N_4324,In_1744,In_1032);
xor U4325 (N_4325,In_1688,In_1934);
nand U4326 (N_4326,In_2338,In_771);
nor U4327 (N_4327,In_23,In_662);
and U4328 (N_4328,In_528,In_1063);
and U4329 (N_4329,In_1952,In_2015);
xor U4330 (N_4330,In_1793,In_1272);
nor U4331 (N_4331,In_1768,In_147);
nand U4332 (N_4332,In_1041,In_1599);
or U4333 (N_4333,In_2180,In_611);
and U4334 (N_4334,In_1573,In_1065);
nand U4335 (N_4335,In_1297,In_90);
nand U4336 (N_4336,In_1654,In_888);
xnor U4337 (N_4337,In_237,In_2136);
nor U4338 (N_4338,In_1871,In_1856);
xnor U4339 (N_4339,In_2314,In_1925);
nand U4340 (N_4340,In_1702,In_2112);
and U4341 (N_4341,In_8,In_2471);
or U4342 (N_4342,In_2176,In_1130);
or U4343 (N_4343,In_549,In_413);
and U4344 (N_4344,In_308,In_617);
xor U4345 (N_4345,In_1010,In_136);
nand U4346 (N_4346,In_1141,In_1147);
xor U4347 (N_4347,In_1924,In_1475);
xnor U4348 (N_4348,In_2189,In_2452);
and U4349 (N_4349,In_1349,In_2151);
nor U4350 (N_4350,In_0,In_2429);
or U4351 (N_4351,In_974,In_2159);
nand U4352 (N_4352,In_195,In_1725);
nand U4353 (N_4353,In_964,In_329);
nor U4354 (N_4354,In_711,In_953);
nand U4355 (N_4355,In_875,In_1631);
nor U4356 (N_4356,In_1423,In_2262);
nand U4357 (N_4357,In_2322,In_2022);
nand U4358 (N_4358,In_2404,In_2380);
xnor U4359 (N_4359,In_2144,In_2475);
and U4360 (N_4360,In_945,In_1939);
xnor U4361 (N_4361,In_1653,In_1493);
nand U4362 (N_4362,In_2175,In_1096);
or U4363 (N_4363,In_430,In_895);
and U4364 (N_4364,In_529,In_474);
and U4365 (N_4365,In_1680,In_986);
nand U4366 (N_4366,In_1263,In_1253);
and U4367 (N_4367,In_818,In_1249);
nand U4368 (N_4368,In_285,In_308);
xnor U4369 (N_4369,In_949,In_2307);
nand U4370 (N_4370,In_2156,In_269);
nor U4371 (N_4371,In_22,In_1345);
nand U4372 (N_4372,In_1459,In_710);
or U4373 (N_4373,In_1525,In_883);
nor U4374 (N_4374,In_2455,In_1834);
xor U4375 (N_4375,In_847,In_1399);
nand U4376 (N_4376,In_1352,In_2455);
or U4377 (N_4377,In_459,In_1746);
nor U4378 (N_4378,In_1653,In_5);
nor U4379 (N_4379,In_566,In_1797);
or U4380 (N_4380,In_863,In_1913);
nand U4381 (N_4381,In_2133,In_1418);
or U4382 (N_4382,In_2368,In_1856);
xor U4383 (N_4383,In_577,In_1896);
nor U4384 (N_4384,In_2423,In_448);
and U4385 (N_4385,In_2168,In_449);
nand U4386 (N_4386,In_2440,In_689);
or U4387 (N_4387,In_1304,In_1389);
nand U4388 (N_4388,In_547,In_6);
xor U4389 (N_4389,In_2402,In_1595);
or U4390 (N_4390,In_898,In_1145);
xor U4391 (N_4391,In_1389,In_1404);
nand U4392 (N_4392,In_1544,In_722);
and U4393 (N_4393,In_1769,In_69);
or U4394 (N_4394,In_1752,In_2303);
or U4395 (N_4395,In_1203,In_2113);
xnor U4396 (N_4396,In_2301,In_1356);
nor U4397 (N_4397,In_2004,In_2116);
xnor U4398 (N_4398,In_59,In_880);
nor U4399 (N_4399,In_65,In_1038);
xor U4400 (N_4400,In_57,In_426);
nand U4401 (N_4401,In_440,In_323);
xnor U4402 (N_4402,In_1576,In_2149);
nand U4403 (N_4403,In_251,In_1881);
nor U4404 (N_4404,In_1950,In_1229);
xor U4405 (N_4405,In_983,In_2061);
nor U4406 (N_4406,In_1938,In_2292);
nand U4407 (N_4407,In_2382,In_2280);
xor U4408 (N_4408,In_1309,In_515);
or U4409 (N_4409,In_715,In_379);
xor U4410 (N_4410,In_436,In_408);
nor U4411 (N_4411,In_1312,In_2452);
and U4412 (N_4412,In_2047,In_1337);
xor U4413 (N_4413,In_912,In_551);
nand U4414 (N_4414,In_1646,In_188);
xnor U4415 (N_4415,In_1948,In_615);
nor U4416 (N_4416,In_1657,In_251);
xor U4417 (N_4417,In_2361,In_880);
nand U4418 (N_4418,In_967,In_2329);
nand U4419 (N_4419,In_1365,In_1881);
nand U4420 (N_4420,In_175,In_744);
xor U4421 (N_4421,In_1558,In_1411);
nand U4422 (N_4422,In_488,In_794);
or U4423 (N_4423,In_1812,In_1188);
nand U4424 (N_4424,In_2103,In_1326);
or U4425 (N_4425,In_1979,In_2047);
nand U4426 (N_4426,In_1846,In_2298);
and U4427 (N_4427,In_1811,In_1633);
nor U4428 (N_4428,In_844,In_2355);
nand U4429 (N_4429,In_2148,In_2165);
xor U4430 (N_4430,In_977,In_2200);
nand U4431 (N_4431,In_915,In_2135);
nor U4432 (N_4432,In_1643,In_1028);
xor U4433 (N_4433,In_141,In_1195);
or U4434 (N_4434,In_1577,In_2157);
or U4435 (N_4435,In_2453,In_1812);
nor U4436 (N_4436,In_1539,In_140);
nand U4437 (N_4437,In_677,In_87);
or U4438 (N_4438,In_560,In_520);
and U4439 (N_4439,In_62,In_1021);
nor U4440 (N_4440,In_1513,In_2462);
or U4441 (N_4441,In_1985,In_2413);
nand U4442 (N_4442,In_325,In_2157);
nor U4443 (N_4443,In_1862,In_2485);
xor U4444 (N_4444,In_960,In_2463);
nand U4445 (N_4445,In_2181,In_273);
and U4446 (N_4446,In_2193,In_2373);
xor U4447 (N_4447,In_2127,In_1967);
nand U4448 (N_4448,In_523,In_2190);
nor U4449 (N_4449,In_1500,In_931);
xnor U4450 (N_4450,In_1175,In_1205);
xnor U4451 (N_4451,In_1691,In_1247);
or U4452 (N_4452,In_364,In_883);
nor U4453 (N_4453,In_998,In_2161);
nand U4454 (N_4454,In_1355,In_2225);
nand U4455 (N_4455,In_2479,In_1100);
nand U4456 (N_4456,In_2301,In_684);
xnor U4457 (N_4457,In_1122,In_1757);
nand U4458 (N_4458,In_1947,In_477);
or U4459 (N_4459,In_1910,In_2218);
nor U4460 (N_4460,In_479,In_1253);
nand U4461 (N_4461,In_651,In_110);
nor U4462 (N_4462,In_2468,In_1871);
and U4463 (N_4463,In_110,In_1566);
nor U4464 (N_4464,In_1129,In_1231);
nand U4465 (N_4465,In_574,In_2439);
or U4466 (N_4466,In_623,In_1629);
nand U4467 (N_4467,In_1068,In_372);
nand U4468 (N_4468,In_139,In_895);
or U4469 (N_4469,In_1996,In_1120);
nor U4470 (N_4470,In_1642,In_1142);
nor U4471 (N_4471,In_1398,In_1216);
nor U4472 (N_4472,In_297,In_284);
or U4473 (N_4473,In_2360,In_592);
nand U4474 (N_4474,In_1548,In_569);
and U4475 (N_4475,In_1277,In_1247);
nand U4476 (N_4476,In_2146,In_644);
xnor U4477 (N_4477,In_169,In_157);
and U4478 (N_4478,In_1286,In_953);
or U4479 (N_4479,In_1629,In_2100);
or U4480 (N_4480,In_1427,In_903);
nand U4481 (N_4481,In_1886,In_1820);
or U4482 (N_4482,In_423,In_1594);
or U4483 (N_4483,In_1569,In_381);
or U4484 (N_4484,In_72,In_1203);
xnor U4485 (N_4485,In_1894,In_554);
nand U4486 (N_4486,In_7,In_244);
xor U4487 (N_4487,In_424,In_2273);
nor U4488 (N_4488,In_1885,In_1596);
nor U4489 (N_4489,In_1290,In_226);
nor U4490 (N_4490,In_2264,In_384);
or U4491 (N_4491,In_126,In_545);
or U4492 (N_4492,In_64,In_1424);
and U4493 (N_4493,In_2160,In_1714);
nand U4494 (N_4494,In_711,In_1258);
nand U4495 (N_4495,In_823,In_792);
xnor U4496 (N_4496,In_1589,In_69);
and U4497 (N_4497,In_43,In_1580);
nor U4498 (N_4498,In_911,In_248);
and U4499 (N_4499,In_2074,In_2358);
xnor U4500 (N_4500,In_1423,In_1317);
nor U4501 (N_4501,In_1465,In_1219);
nand U4502 (N_4502,In_1019,In_2283);
and U4503 (N_4503,In_2019,In_1174);
nand U4504 (N_4504,In_906,In_1967);
and U4505 (N_4505,In_962,In_674);
xnor U4506 (N_4506,In_2089,In_1620);
nor U4507 (N_4507,In_623,In_2341);
and U4508 (N_4508,In_387,In_789);
nand U4509 (N_4509,In_1676,In_2222);
and U4510 (N_4510,In_796,In_552);
nand U4511 (N_4511,In_790,In_145);
and U4512 (N_4512,In_1059,In_2493);
nand U4513 (N_4513,In_1159,In_2233);
nand U4514 (N_4514,In_2463,In_1146);
nand U4515 (N_4515,In_1344,In_262);
nand U4516 (N_4516,In_1521,In_819);
nand U4517 (N_4517,In_773,In_2187);
nor U4518 (N_4518,In_382,In_694);
or U4519 (N_4519,In_927,In_1315);
or U4520 (N_4520,In_164,In_457);
xnor U4521 (N_4521,In_2189,In_1128);
xor U4522 (N_4522,In_440,In_28);
or U4523 (N_4523,In_1900,In_312);
or U4524 (N_4524,In_1937,In_2000);
nor U4525 (N_4525,In_917,In_698);
nor U4526 (N_4526,In_878,In_1734);
nor U4527 (N_4527,In_246,In_114);
nand U4528 (N_4528,In_1224,In_720);
nand U4529 (N_4529,In_2464,In_1489);
nand U4530 (N_4530,In_94,In_95);
nand U4531 (N_4531,In_1928,In_1322);
and U4532 (N_4532,In_939,In_1001);
or U4533 (N_4533,In_310,In_1980);
nand U4534 (N_4534,In_2375,In_1409);
or U4535 (N_4535,In_13,In_1448);
xnor U4536 (N_4536,In_1434,In_633);
or U4537 (N_4537,In_1231,In_2317);
nand U4538 (N_4538,In_1159,In_1677);
nor U4539 (N_4539,In_1765,In_475);
xor U4540 (N_4540,In_2004,In_843);
nor U4541 (N_4541,In_231,In_2220);
xnor U4542 (N_4542,In_2469,In_252);
nand U4543 (N_4543,In_676,In_190);
xnor U4544 (N_4544,In_2368,In_2058);
xnor U4545 (N_4545,In_1438,In_355);
and U4546 (N_4546,In_1251,In_2005);
or U4547 (N_4547,In_416,In_2089);
nor U4548 (N_4548,In_2486,In_37);
and U4549 (N_4549,In_1917,In_758);
nor U4550 (N_4550,In_942,In_241);
nand U4551 (N_4551,In_627,In_370);
or U4552 (N_4552,In_2004,In_1783);
and U4553 (N_4553,In_715,In_1145);
or U4554 (N_4554,In_1764,In_1959);
nor U4555 (N_4555,In_1771,In_2039);
nor U4556 (N_4556,In_1574,In_1973);
nand U4557 (N_4557,In_2284,In_677);
nand U4558 (N_4558,In_743,In_354);
nor U4559 (N_4559,In_2373,In_1392);
and U4560 (N_4560,In_451,In_567);
and U4561 (N_4561,In_1347,In_437);
nor U4562 (N_4562,In_1041,In_256);
or U4563 (N_4563,In_2312,In_2415);
nor U4564 (N_4564,In_735,In_51);
nand U4565 (N_4565,In_1097,In_2028);
nand U4566 (N_4566,In_1254,In_24);
nor U4567 (N_4567,In_588,In_1206);
nand U4568 (N_4568,In_1443,In_543);
or U4569 (N_4569,In_1765,In_1753);
or U4570 (N_4570,In_2276,In_913);
or U4571 (N_4571,In_2495,In_1214);
nand U4572 (N_4572,In_141,In_1154);
or U4573 (N_4573,In_2447,In_2022);
or U4574 (N_4574,In_108,In_928);
nand U4575 (N_4575,In_1209,In_2300);
nor U4576 (N_4576,In_2352,In_1472);
nand U4577 (N_4577,In_1682,In_339);
nand U4578 (N_4578,In_195,In_955);
nor U4579 (N_4579,In_2071,In_450);
or U4580 (N_4580,In_860,In_645);
and U4581 (N_4581,In_2097,In_421);
or U4582 (N_4582,In_1194,In_723);
xnor U4583 (N_4583,In_702,In_735);
and U4584 (N_4584,In_1825,In_2085);
nand U4585 (N_4585,In_1561,In_2472);
xor U4586 (N_4586,In_881,In_1810);
nor U4587 (N_4587,In_345,In_137);
nand U4588 (N_4588,In_1996,In_1649);
nand U4589 (N_4589,In_23,In_1547);
or U4590 (N_4590,In_668,In_1077);
nor U4591 (N_4591,In_467,In_280);
nor U4592 (N_4592,In_884,In_190);
and U4593 (N_4593,In_1710,In_2116);
nor U4594 (N_4594,In_1938,In_1329);
xor U4595 (N_4595,In_620,In_327);
and U4596 (N_4596,In_806,In_1927);
nand U4597 (N_4597,In_2399,In_1604);
nand U4598 (N_4598,In_715,In_810);
nor U4599 (N_4599,In_1549,In_1910);
nor U4600 (N_4600,In_644,In_153);
and U4601 (N_4601,In_1942,In_1048);
or U4602 (N_4602,In_1363,In_2498);
nand U4603 (N_4603,In_1825,In_1556);
xnor U4604 (N_4604,In_416,In_1454);
nand U4605 (N_4605,In_208,In_153);
and U4606 (N_4606,In_1982,In_305);
xor U4607 (N_4607,In_1656,In_1267);
and U4608 (N_4608,In_101,In_10);
nor U4609 (N_4609,In_485,In_1435);
xor U4610 (N_4610,In_1913,In_600);
and U4611 (N_4611,In_388,In_360);
or U4612 (N_4612,In_1497,In_51);
nand U4613 (N_4613,In_2401,In_1974);
xnor U4614 (N_4614,In_1590,In_82);
and U4615 (N_4615,In_95,In_1924);
xnor U4616 (N_4616,In_1578,In_1143);
nand U4617 (N_4617,In_1886,In_807);
nor U4618 (N_4618,In_1149,In_401);
or U4619 (N_4619,In_384,In_685);
or U4620 (N_4620,In_10,In_17);
and U4621 (N_4621,In_1229,In_1264);
nand U4622 (N_4622,In_89,In_190);
and U4623 (N_4623,In_461,In_922);
or U4624 (N_4624,In_1392,In_1292);
xnor U4625 (N_4625,In_1945,In_403);
and U4626 (N_4626,In_481,In_759);
and U4627 (N_4627,In_1354,In_2158);
nand U4628 (N_4628,In_1451,In_2202);
nor U4629 (N_4629,In_342,In_805);
xor U4630 (N_4630,In_450,In_1931);
or U4631 (N_4631,In_1984,In_190);
nor U4632 (N_4632,In_971,In_371);
or U4633 (N_4633,In_1844,In_2242);
nand U4634 (N_4634,In_1432,In_281);
or U4635 (N_4635,In_1379,In_2198);
nand U4636 (N_4636,In_1828,In_1444);
xnor U4637 (N_4637,In_1457,In_1795);
and U4638 (N_4638,In_422,In_432);
and U4639 (N_4639,In_808,In_190);
or U4640 (N_4640,In_1651,In_2271);
nor U4641 (N_4641,In_1191,In_784);
xor U4642 (N_4642,In_1745,In_804);
and U4643 (N_4643,In_1829,In_2477);
and U4644 (N_4644,In_1455,In_1479);
nor U4645 (N_4645,In_2178,In_1059);
or U4646 (N_4646,In_2490,In_717);
xnor U4647 (N_4647,In_1816,In_1203);
xor U4648 (N_4648,In_768,In_1330);
or U4649 (N_4649,In_200,In_1086);
nor U4650 (N_4650,In_245,In_919);
xnor U4651 (N_4651,In_67,In_1407);
xor U4652 (N_4652,In_19,In_1217);
nand U4653 (N_4653,In_570,In_366);
xnor U4654 (N_4654,In_368,In_1633);
nor U4655 (N_4655,In_38,In_565);
nand U4656 (N_4656,In_45,In_1248);
or U4657 (N_4657,In_1613,In_428);
xnor U4658 (N_4658,In_1037,In_1702);
nand U4659 (N_4659,In_881,In_188);
and U4660 (N_4660,In_1769,In_1205);
or U4661 (N_4661,In_15,In_228);
nor U4662 (N_4662,In_1884,In_393);
or U4663 (N_4663,In_1055,In_1292);
xor U4664 (N_4664,In_1059,In_911);
nand U4665 (N_4665,In_1658,In_1457);
and U4666 (N_4666,In_810,In_1665);
or U4667 (N_4667,In_666,In_1);
and U4668 (N_4668,In_1216,In_1847);
xor U4669 (N_4669,In_341,In_1904);
or U4670 (N_4670,In_731,In_674);
nand U4671 (N_4671,In_517,In_646);
nor U4672 (N_4672,In_1496,In_1565);
xnor U4673 (N_4673,In_350,In_386);
nand U4674 (N_4674,In_2038,In_1301);
xor U4675 (N_4675,In_702,In_1403);
and U4676 (N_4676,In_442,In_1361);
nand U4677 (N_4677,In_2115,In_210);
xor U4678 (N_4678,In_2079,In_572);
or U4679 (N_4679,In_2002,In_1697);
or U4680 (N_4680,In_2488,In_1231);
xnor U4681 (N_4681,In_949,In_1746);
nand U4682 (N_4682,In_375,In_1763);
nand U4683 (N_4683,In_1760,In_677);
nand U4684 (N_4684,In_2322,In_632);
nor U4685 (N_4685,In_2234,In_2094);
nor U4686 (N_4686,In_1192,In_1726);
nand U4687 (N_4687,In_813,In_1145);
xor U4688 (N_4688,In_9,In_363);
nor U4689 (N_4689,In_1077,In_1926);
xor U4690 (N_4690,In_1302,In_605);
nand U4691 (N_4691,In_2196,In_131);
nor U4692 (N_4692,In_183,In_1821);
and U4693 (N_4693,In_2498,In_614);
nor U4694 (N_4694,In_156,In_1728);
or U4695 (N_4695,In_1392,In_2208);
nand U4696 (N_4696,In_742,In_1880);
xor U4697 (N_4697,In_477,In_451);
nor U4698 (N_4698,In_1885,In_1458);
and U4699 (N_4699,In_1972,In_2113);
or U4700 (N_4700,In_792,In_2211);
xor U4701 (N_4701,In_1008,In_55);
or U4702 (N_4702,In_1876,In_1385);
or U4703 (N_4703,In_205,In_1985);
nand U4704 (N_4704,In_337,In_1351);
xor U4705 (N_4705,In_1215,In_2129);
xor U4706 (N_4706,In_1537,In_1672);
xor U4707 (N_4707,In_420,In_1381);
xnor U4708 (N_4708,In_1321,In_2365);
nand U4709 (N_4709,In_2238,In_630);
xnor U4710 (N_4710,In_1310,In_1521);
xor U4711 (N_4711,In_2119,In_416);
or U4712 (N_4712,In_1744,In_78);
xnor U4713 (N_4713,In_886,In_2145);
nand U4714 (N_4714,In_448,In_1149);
xor U4715 (N_4715,In_1830,In_428);
nand U4716 (N_4716,In_653,In_299);
or U4717 (N_4717,In_1246,In_1169);
nor U4718 (N_4718,In_1881,In_1759);
nor U4719 (N_4719,In_768,In_144);
and U4720 (N_4720,In_714,In_2075);
nand U4721 (N_4721,In_811,In_1590);
nor U4722 (N_4722,In_1645,In_2298);
nand U4723 (N_4723,In_366,In_1682);
xnor U4724 (N_4724,In_4,In_161);
and U4725 (N_4725,In_650,In_438);
or U4726 (N_4726,In_504,In_2457);
nor U4727 (N_4727,In_197,In_2294);
xnor U4728 (N_4728,In_891,In_2176);
nor U4729 (N_4729,In_501,In_1919);
nand U4730 (N_4730,In_1288,In_1715);
or U4731 (N_4731,In_1812,In_2488);
nor U4732 (N_4732,In_1189,In_775);
nand U4733 (N_4733,In_1499,In_2448);
nand U4734 (N_4734,In_530,In_2117);
or U4735 (N_4735,In_2031,In_1016);
or U4736 (N_4736,In_1004,In_502);
or U4737 (N_4737,In_958,In_1426);
nor U4738 (N_4738,In_431,In_596);
nor U4739 (N_4739,In_2317,In_1968);
and U4740 (N_4740,In_996,In_1665);
and U4741 (N_4741,In_718,In_1813);
nor U4742 (N_4742,In_162,In_2210);
or U4743 (N_4743,In_534,In_1448);
xnor U4744 (N_4744,In_1716,In_1847);
nand U4745 (N_4745,In_567,In_1125);
xor U4746 (N_4746,In_2116,In_1816);
and U4747 (N_4747,In_221,In_993);
and U4748 (N_4748,In_365,In_1527);
nand U4749 (N_4749,In_813,In_760);
xor U4750 (N_4750,In_1561,In_1903);
xnor U4751 (N_4751,In_664,In_209);
xnor U4752 (N_4752,In_1092,In_2341);
nor U4753 (N_4753,In_343,In_121);
xnor U4754 (N_4754,In_2097,In_1405);
nor U4755 (N_4755,In_1686,In_2399);
or U4756 (N_4756,In_1556,In_392);
nand U4757 (N_4757,In_531,In_1773);
and U4758 (N_4758,In_1907,In_587);
or U4759 (N_4759,In_2300,In_288);
or U4760 (N_4760,In_757,In_995);
nor U4761 (N_4761,In_1082,In_1382);
and U4762 (N_4762,In_2368,In_1924);
nor U4763 (N_4763,In_2116,In_1618);
nand U4764 (N_4764,In_1152,In_2360);
nor U4765 (N_4765,In_40,In_719);
or U4766 (N_4766,In_2472,In_129);
xnor U4767 (N_4767,In_548,In_871);
and U4768 (N_4768,In_1840,In_2091);
and U4769 (N_4769,In_866,In_1761);
and U4770 (N_4770,In_1815,In_677);
nand U4771 (N_4771,In_1257,In_578);
nand U4772 (N_4772,In_1315,In_419);
or U4773 (N_4773,In_2311,In_318);
or U4774 (N_4774,In_2341,In_1207);
nor U4775 (N_4775,In_1602,In_1259);
nand U4776 (N_4776,In_1665,In_1161);
nor U4777 (N_4777,In_287,In_1029);
or U4778 (N_4778,In_1138,In_341);
and U4779 (N_4779,In_1221,In_923);
xor U4780 (N_4780,In_1149,In_1392);
or U4781 (N_4781,In_1575,In_1799);
and U4782 (N_4782,In_1264,In_1708);
and U4783 (N_4783,In_267,In_252);
nor U4784 (N_4784,In_1653,In_719);
nor U4785 (N_4785,In_1085,In_837);
nand U4786 (N_4786,In_2165,In_2356);
nand U4787 (N_4787,In_1601,In_461);
nand U4788 (N_4788,In_584,In_588);
xor U4789 (N_4789,In_2426,In_2298);
and U4790 (N_4790,In_1007,In_2299);
or U4791 (N_4791,In_491,In_1705);
nor U4792 (N_4792,In_2180,In_1982);
nand U4793 (N_4793,In_1279,In_2474);
or U4794 (N_4794,In_380,In_2283);
and U4795 (N_4795,In_145,In_1727);
or U4796 (N_4796,In_97,In_2446);
xnor U4797 (N_4797,In_184,In_2339);
nor U4798 (N_4798,In_629,In_2161);
or U4799 (N_4799,In_2443,In_2213);
xnor U4800 (N_4800,In_1623,In_1144);
xor U4801 (N_4801,In_1369,In_450);
xnor U4802 (N_4802,In_636,In_127);
xor U4803 (N_4803,In_872,In_378);
or U4804 (N_4804,In_2206,In_1255);
xnor U4805 (N_4805,In_1590,In_1469);
or U4806 (N_4806,In_1021,In_526);
or U4807 (N_4807,In_2226,In_1546);
nand U4808 (N_4808,In_2318,In_898);
and U4809 (N_4809,In_449,In_2046);
or U4810 (N_4810,In_1508,In_2368);
or U4811 (N_4811,In_1947,In_336);
or U4812 (N_4812,In_308,In_63);
xnor U4813 (N_4813,In_2301,In_1199);
xor U4814 (N_4814,In_2236,In_2045);
xor U4815 (N_4815,In_1946,In_1202);
xor U4816 (N_4816,In_851,In_1375);
nor U4817 (N_4817,In_1056,In_1952);
nand U4818 (N_4818,In_1963,In_1126);
xnor U4819 (N_4819,In_2104,In_2438);
and U4820 (N_4820,In_1851,In_593);
nand U4821 (N_4821,In_49,In_1921);
nor U4822 (N_4822,In_2086,In_1218);
nor U4823 (N_4823,In_656,In_1942);
nor U4824 (N_4824,In_2447,In_597);
or U4825 (N_4825,In_462,In_1573);
xnor U4826 (N_4826,In_1571,In_1874);
and U4827 (N_4827,In_158,In_800);
xnor U4828 (N_4828,In_765,In_1040);
nand U4829 (N_4829,In_1815,In_47);
or U4830 (N_4830,In_1191,In_1245);
or U4831 (N_4831,In_2383,In_1311);
and U4832 (N_4832,In_2384,In_306);
or U4833 (N_4833,In_975,In_21);
or U4834 (N_4834,In_1721,In_977);
and U4835 (N_4835,In_2144,In_2044);
and U4836 (N_4836,In_51,In_2157);
xor U4837 (N_4837,In_1562,In_633);
nor U4838 (N_4838,In_2002,In_2009);
and U4839 (N_4839,In_477,In_933);
or U4840 (N_4840,In_2001,In_2045);
nand U4841 (N_4841,In_1106,In_2439);
or U4842 (N_4842,In_2021,In_2119);
nor U4843 (N_4843,In_2318,In_1400);
nand U4844 (N_4844,In_275,In_2110);
or U4845 (N_4845,In_1533,In_2458);
nor U4846 (N_4846,In_1201,In_1491);
nand U4847 (N_4847,In_859,In_486);
nand U4848 (N_4848,In_2072,In_2283);
nor U4849 (N_4849,In_2149,In_927);
nor U4850 (N_4850,In_810,In_2286);
and U4851 (N_4851,In_1938,In_1048);
and U4852 (N_4852,In_2131,In_17);
nand U4853 (N_4853,In_538,In_1063);
or U4854 (N_4854,In_1435,In_2219);
or U4855 (N_4855,In_1468,In_126);
nor U4856 (N_4856,In_2088,In_1453);
or U4857 (N_4857,In_720,In_1469);
xnor U4858 (N_4858,In_181,In_1932);
or U4859 (N_4859,In_610,In_2473);
and U4860 (N_4860,In_684,In_311);
nor U4861 (N_4861,In_1854,In_1467);
nor U4862 (N_4862,In_1377,In_2250);
or U4863 (N_4863,In_834,In_2300);
or U4864 (N_4864,In_1352,In_2038);
or U4865 (N_4865,In_1835,In_686);
or U4866 (N_4866,In_259,In_408);
or U4867 (N_4867,In_1132,In_1174);
nand U4868 (N_4868,In_2180,In_1021);
nand U4869 (N_4869,In_2326,In_586);
xor U4870 (N_4870,In_2373,In_1308);
nor U4871 (N_4871,In_1582,In_442);
nand U4872 (N_4872,In_1451,In_436);
nand U4873 (N_4873,In_2492,In_729);
and U4874 (N_4874,In_1792,In_1666);
xor U4875 (N_4875,In_228,In_1076);
nor U4876 (N_4876,In_323,In_1719);
xor U4877 (N_4877,In_1739,In_971);
xnor U4878 (N_4878,In_1837,In_2412);
nor U4879 (N_4879,In_717,In_1571);
nand U4880 (N_4880,In_1437,In_11);
nor U4881 (N_4881,In_1520,In_574);
or U4882 (N_4882,In_62,In_1990);
nand U4883 (N_4883,In_1750,In_919);
nor U4884 (N_4884,In_2107,In_571);
nor U4885 (N_4885,In_723,In_277);
xnor U4886 (N_4886,In_337,In_452);
or U4887 (N_4887,In_171,In_2249);
xor U4888 (N_4888,In_964,In_1419);
and U4889 (N_4889,In_579,In_772);
xor U4890 (N_4890,In_1843,In_2145);
xor U4891 (N_4891,In_2454,In_413);
or U4892 (N_4892,In_1368,In_825);
nand U4893 (N_4893,In_1807,In_1157);
xnor U4894 (N_4894,In_493,In_1670);
and U4895 (N_4895,In_985,In_241);
nand U4896 (N_4896,In_1538,In_2427);
nor U4897 (N_4897,In_406,In_130);
or U4898 (N_4898,In_1909,In_1313);
nand U4899 (N_4899,In_2161,In_173);
nor U4900 (N_4900,In_2061,In_466);
and U4901 (N_4901,In_1386,In_1989);
or U4902 (N_4902,In_1963,In_1400);
xor U4903 (N_4903,In_2268,In_1495);
nor U4904 (N_4904,In_1371,In_1736);
or U4905 (N_4905,In_1395,In_1769);
nand U4906 (N_4906,In_129,In_647);
nor U4907 (N_4907,In_2031,In_2072);
and U4908 (N_4908,In_513,In_2355);
nand U4909 (N_4909,In_2024,In_1795);
nand U4910 (N_4910,In_276,In_140);
nand U4911 (N_4911,In_1296,In_1536);
and U4912 (N_4912,In_1054,In_1456);
and U4913 (N_4913,In_99,In_2460);
and U4914 (N_4914,In_1800,In_1989);
and U4915 (N_4915,In_2093,In_2099);
nand U4916 (N_4916,In_1615,In_2116);
nand U4917 (N_4917,In_2293,In_420);
nor U4918 (N_4918,In_2123,In_657);
nor U4919 (N_4919,In_233,In_2191);
nand U4920 (N_4920,In_2394,In_1945);
and U4921 (N_4921,In_505,In_1156);
nor U4922 (N_4922,In_1064,In_762);
and U4923 (N_4923,In_136,In_1289);
and U4924 (N_4924,In_776,In_2262);
nand U4925 (N_4925,In_900,In_910);
nand U4926 (N_4926,In_2439,In_277);
or U4927 (N_4927,In_192,In_1757);
nand U4928 (N_4928,In_750,In_1052);
and U4929 (N_4929,In_2022,In_747);
nor U4930 (N_4930,In_1452,In_1836);
and U4931 (N_4931,In_2177,In_2095);
nor U4932 (N_4932,In_133,In_2135);
and U4933 (N_4933,In_2060,In_1092);
and U4934 (N_4934,In_387,In_1457);
nand U4935 (N_4935,In_1422,In_803);
or U4936 (N_4936,In_2220,In_605);
nand U4937 (N_4937,In_1218,In_2443);
nand U4938 (N_4938,In_1975,In_2194);
or U4939 (N_4939,In_1989,In_824);
xor U4940 (N_4940,In_1743,In_1748);
xor U4941 (N_4941,In_674,In_1026);
xor U4942 (N_4942,In_1173,In_1079);
or U4943 (N_4943,In_1381,In_190);
nor U4944 (N_4944,In_1383,In_1155);
nand U4945 (N_4945,In_65,In_2040);
nand U4946 (N_4946,In_999,In_1853);
or U4947 (N_4947,In_985,In_1489);
xnor U4948 (N_4948,In_1246,In_1963);
xor U4949 (N_4949,In_1486,In_2204);
or U4950 (N_4950,In_404,In_1662);
nor U4951 (N_4951,In_81,In_2074);
and U4952 (N_4952,In_1906,In_113);
nor U4953 (N_4953,In_2098,In_2289);
xnor U4954 (N_4954,In_1867,In_1323);
nand U4955 (N_4955,In_309,In_1529);
xor U4956 (N_4956,In_635,In_1886);
nor U4957 (N_4957,In_1964,In_2297);
nand U4958 (N_4958,In_451,In_1763);
nand U4959 (N_4959,In_2324,In_1105);
xor U4960 (N_4960,In_303,In_1734);
xnor U4961 (N_4961,In_2034,In_1427);
or U4962 (N_4962,In_2028,In_2319);
nand U4963 (N_4963,In_876,In_776);
and U4964 (N_4964,In_141,In_1566);
and U4965 (N_4965,In_990,In_1843);
xor U4966 (N_4966,In_1935,In_1388);
nand U4967 (N_4967,In_402,In_1553);
or U4968 (N_4968,In_1505,In_1422);
nand U4969 (N_4969,In_874,In_1738);
and U4970 (N_4970,In_2212,In_1735);
nand U4971 (N_4971,In_1435,In_2397);
nand U4972 (N_4972,In_802,In_1463);
nand U4973 (N_4973,In_2468,In_1329);
and U4974 (N_4974,In_845,In_1642);
and U4975 (N_4975,In_791,In_209);
nor U4976 (N_4976,In_116,In_1538);
or U4977 (N_4977,In_1674,In_1187);
and U4978 (N_4978,In_952,In_2094);
and U4979 (N_4979,In_214,In_1939);
xor U4980 (N_4980,In_1722,In_1218);
xnor U4981 (N_4981,In_1928,In_170);
nor U4982 (N_4982,In_1981,In_446);
nor U4983 (N_4983,In_1523,In_823);
nor U4984 (N_4984,In_621,In_1696);
nand U4985 (N_4985,In_493,In_1422);
nor U4986 (N_4986,In_1994,In_1614);
xor U4987 (N_4987,In_1545,In_188);
nor U4988 (N_4988,In_38,In_1821);
or U4989 (N_4989,In_2298,In_2089);
nand U4990 (N_4990,In_669,In_569);
nor U4991 (N_4991,In_2473,In_640);
nor U4992 (N_4992,In_429,In_1874);
or U4993 (N_4993,In_1429,In_450);
nand U4994 (N_4994,In_2168,In_2203);
or U4995 (N_4995,In_2274,In_2271);
nand U4996 (N_4996,In_2006,In_408);
nand U4997 (N_4997,In_1621,In_2438);
xor U4998 (N_4998,In_2352,In_689);
or U4999 (N_4999,In_2497,In_2107);
xnor U5000 (N_5000,N_3899,N_3564);
xnor U5001 (N_5001,N_1848,N_3262);
xnor U5002 (N_5002,N_3773,N_658);
nand U5003 (N_5003,N_1582,N_3378);
nand U5004 (N_5004,N_2930,N_1914);
nand U5005 (N_5005,N_4618,N_256);
or U5006 (N_5006,N_3739,N_143);
nand U5007 (N_5007,N_146,N_3430);
xnor U5008 (N_5008,N_1992,N_1382);
nor U5009 (N_5009,N_159,N_2792);
and U5010 (N_5010,N_547,N_3491);
xnor U5011 (N_5011,N_1539,N_493);
nor U5012 (N_5012,N_2785,N_4836);
or U5013 (N_5013,N_4360,N_503);
and U5014 (N_5014,N_2411,N_2441);
or U5015 (N_5015,N_4697,N_2535);
nand U5016 (N_5016,N_2439,N_2848);
or U5017 (N_5017,N_1837,N_3371);
nand U5018 (N_5018,N_29,N_1588);
nand U5019 (N_5019,N_3776,N_3627);
xor U5020 (N_5020,N_95,N_3244);
and U5021 (N_5021,N_4987,N_567);
xor U5022 (N_5022,N_2749,N_857);
and U5023 (N_5023,N_229,N_957);
and U5024 (N_5024,N_1981,N_1260);
nor U5025 (N_5025,N_2883,N_2084);
and U5026 (N_5026,N_4095,N_953);
nand U5027 (N_5027,N_2213,N_584);
and U5028 (N_5028,N_3935,N_4730);
or U5029 (N_5029,N_2038,N_4170);
and U5030 (N_5030,N_2832,N_2582);
or U5031 (N_5031,N_1909,N_3988);
nor U5032 (N_5032,N_3152,N_921);
or U5033 (N_5033,N_2207,N_4364);
and U5034 (N_5034,N_410,N_2352);
nand U5035 (N_5035,N_1092,N_1548);
and U5036 (N_5036,N_3001,N_4680);
or U5037 (N_5037,N_849,N_461);
or U5038 (N_5038,N_1891,N_2236);
nor U5039 (N_5039,N_2019,N_2590);
nor U5040 (N_5040,N_636,N_2007);
nor U5041 (N_5041,N_655,N_2363);
nand U5042 (N_5042,N_4312,N_942);
or U5043 (N_5043,N_1980,N_1551);
and U5044 (N_5044,N_994,N_3661);
and U5045 (N_5045,N_1807,N_3039);
nand U5046 (N_5046,N_376,N_4406);
and U5047 (N_5047,N_1082,N_2399);
nand U5048 (N_5048,N_3847,N_3401);
or U5049 (N_5049,N_2840,N_3216);
or U5050 (N_5050,N_2760,N_1762);
xor U5051 (N_5051,N_70,N_3275);
nor U5052 (N_5052,N_2457,N_753);
nor U5053 (N_5053,N_3377,N_3071);
or U5054 (N_5054,N_3850,N_1093);
nor U5055 (N_5055,N_506,N_16);
nor U5056 (N_5056,N_1681,N_4726);
or U5057 (N_5057,N_3867,N_880);
and U5058 (N_5058,N_3750,N_3581);
nor U5059 (N_5059,N_3408,N_3713);
nor U5060 (N_5060,N_2083,N_97);
xor U5061 (N_5061,N_1288,N_577);
and U5062 (N_5062,N_3447,N_3705);
nand U5063 (N_5063,N_228,N_3728);
and U5064 (N_5064,N_534,N_2946);
nand U5065 (N_5065,N_698,N_2464);
nor U5066 (N_5066,N_1477,N_2068);
nor U5067 (N_5067,N_2884,N_1428);
and U5068 (N_5068,N_2280,N_3568);
xnor U5069 (N_5069,N_4340,N_2981);
or U5070 (N_5070,N_3424,N_249);
xor U5071 (N_5071,N_2288,N_1400);
or U5072 (N_5072,N_1635,N_355);
xor U5073 (N_5073,N_2603,N_2526);
xor U5074 (N_5074,N_2510,N_1154);
and U5075 (N_5075,N_579,N_1562);
or U5076 (N_5076,N_3306,N_154);
nand U5077 (N_5077,N_2784,N_915);
nor U5078 (N_5078,N_1584,N_3832);
nor U5079 (N_5079,N_273,N_64);
nor U5080 (N_5080,N_543,N_158);
xor U5081 (N_5081,N_360,N_1099);
or U5082 (N_5082,N_2053,N_2716);
or U5083 (N_5083,N_2364,N_2855);
nand U5084 (N_5084,N_2931,N_1739);
or U5085 (N_5085,N_495,N_900);
nand U5086 (N_5086,N_847,N_929);
nand U5087 (N_5087,N_1102,N_601);
nor U5088 (N_5088,N_4249,N_4701);
or U5089 (N_5089,N_4642,N_3552);
xnor U5090 (N_5090,N_4556,N_4519);
xnor U5091 (N_5091,N_650,N_2091);
and U5092 (N_5092,N_4619,N_985);
or U5093 (N_5093,N_2962,N_3024);
xnor U5094 (N_5094,N_1262,N_3175);
or U5095 (N_5095,N_4757,N_3810);
nand U5096 (N_5096,N_1823,N_4808);
or U5097 (N_5097,N_4471,N_1167);
or U5098 (N_5098,N_4358,N_1341);
and U5099 (N_5099,N_3613,N_572);
nand U5100 (N_5100,N_119,N_2004);
or U5101 (N_5101,N_4121,N_2351);
and U5102 (N_5102,N_306,N_2214);
nor U5103 (N_5103,N_4806,N_4425);
and U5104 (N_5104,N_489,N_4637);
and U5105 (N_5105,N_3531,N_4275);
nand U5106 (N_5106,N_791,N_1233);
or U5107 (N_5107,N_1253,N_3629);
or U5108 (N_5108,N_3948,N_3170);
nor U5109 (N_5109,N_860,N_1537);
xnor U5110 (N_5110,N_4223,N_4778);
nand U5111 (N_5111,N_2487,N_2344);
nand U5112 (N_5112,N_751,N_4484);
nand U5113 (N_5113,N_1407,N_2852);
nor U5114 (N_5114,N_2036,N_842);
or U5115 (N_5115,N_1033,N_3906);
xor U5116 (N_5116,N_1519,N_1665);
nand U5117 (N_5117,N_4298,N_529);
xnor U5118 (N_5118,N_2908,N_3213);
nor U5119 (N_5119,N_3287,N_4220);
xor U5120 (N_5120,N_2974,N_2372);
nor U5121 (N_5121,N_3588,N_4698);
xnor U5122 (N_5122,N_2024,N_2198);
or U5123 (N_5123,N_4707,N_2401);
nor U5124 (N_5124,N_3650,N_4973);
and U5125 (N_5125,N_4874,N_394);
and U5126 (N_5126,N_3185,N_381);
xnor U5127 (N_5127,N_4168,N_3733);
nor U5128 (N_5128,N_4190,N_1388);
or U5129 (N_5129,N_2328,N_3748);
xnor U5130 (N_5130,N_3018,N_2703);
or U5131 (N_5131,N_4935,N_2326);
nor U5132 (N_5132,N_4339,N_4147);
nor U5133 (N_5133,N_2955,N_1187);
xor U5134 (N_5134,N_2641,N_3370);
nor U5135 (N_5135,N_4441,N_4611);
and U5136 (N_5136,N_1826,N_1377);
xnor U5137 (N_5137,N_1103,N_4303);
xor U5138 (N_5138,N_482,N_3188);
nand U5139 (N_5139,N_2496,N_2539);
nand U5140 (N_5140,N_426,N_205);
and U5141 (N_5141,N_233,N_4107);
nor U5142 (N_5142,N_3040,N_3577);
and U5143 (N_5143,N_33,N_983);
or U5144 (N_5144,N_3479,N_3372);
or U5145 (N_5145,N_2096,N_49);
or U5146 (N_5146,N_4467,N_3932);
xnor U5147 (N_5147,N_1277,N_1227);
xnor U5148 (N_5148,N_2062,N_2499);
and U5149 (N_5149,N_2398,N_4956);
or U5150 (N_5150,N_1581,N_21);
or U5151 (N_5151,N_121,N_469);
xnor U5152 (N_5152,N_2734,N_1575);
and U5153 (N_5153,N_2208,N_1224);
or U5154 (N_5154,N_289,N_4505);
or U5155 (N_5155,N_1613,N_581);
nor U5156 (N_5156,N_4912,N_1494);
xor U5157 (N_5157,N_1607,N_2879);
xnor U5158 (N_5158,N_3481,N_3116);
nand U5159 (N_5159,N_1905,N_1735);
nor U5160 (N_5160,N_3376,N_4126);
nor U5161 (N_5161,N_4674,N_3781);
or U5162 (N_5162,N_1803,N_1235);
nor U5163 (N_5163,N_3641,N_4338);
xor U5164 (N_5164,N_3182,N_871);
nor U5165 (N_5165,N_806,N_4954);
and U5166 (N_5166,N_855,N_1329);
nand U5167 (N_5167,N_1890,N_285);
nor U5168 (N_5168,N_1879,N_2647);
nand U5169 (N_5169,N_1660,N_1761);
and U5170 (N_5170,N_4625,N_947);
nor U5171 (N_5171,N_508,N_4672);
xnor U5172 (N_5172,N_4919,N_1675);
and U5173 (N_5173,N_2782,N_4574);
and U5174 (N_5174,N_227,N_3614);
nor U5175 (N_5175,N_2315,N_1391);
and U5176 (N_5176,N_1664,N_776);
nand U5177 (N_5177,N_3060,N_2336);
xor U5178 (N_5178,N_4034,N_4396);
and U5179 (N_5179,N_2933,N_2835);
xor U5180 (N_5180,N_3761,N_255);
xnor U5181 (N_5181,N_2559,N_3135);
xor U5182 (N_5182,N_258,N_4463);
or U5183 (N_5183,N_3426,N_3178);
or U5184 (N_5184,N_2113,N_2416);
xor U5185 (N_5185,N_1015,N_4419);
nand U5186 (N_5186,N_2893,N_896);
xor U5187 (N_5187,N_39,N_2808);
nor U5188 (N_5188,N_1107,N_4785);
xnor U5189 (N_5189,N_1789,N_3587);
or U5190 (N_5190,N_2392,N_2786);
nor U5191 (N_5191,N_905,N_60);
nand U5192 (N_5192,N_3789,N_2342);
nand U5193 (N_5193,N_4779,N_1174);
xor U5194 (N_5194,N_212,N_3454);
nor U5195 (N_5195,N_784,N_2713);
nand U5196 (N_5196,N_4663,N_859);
xor U5197 (N_5197,N_3102,N_2064);
nor U5198 (N_5198,N_976,N_3251);
xnor U5199 (N_5199,N_1579,N_3857);
and U5200 (N_5200,N_2124,N_4522);
nor U5201 (N_5201,N_1072,N_4863);
or U5202 (N_5202,N_4890,N_1819);
and U5203 (N_5203,N_3645,N_1485);
nor U5204 (N_5204,N_22,N_1609);
xnor U5205 (N_5205,N_1429,N_1044);
xor U5206 (N_5206,N_1788,N_1899);
xnor U5207 (N_5207,N_3521,N_1917);
nor U5208 (N_5208,N_3979,N_4286);
xnor U5209 (N_5209,N_4616,N_425);
or U5210 (N_5210,N_2632,N_2137);
and U5211 (N_5211,N_4201,N_1692);
or U5212 (N_5212,N_4273,N_4613);
and U5213 (N_5213,N_4938,N_742);
or U5214 (N_5214,N_2391,N_1225);
nand U5215 (N_5215,N_1744,N_1453);
or U5216 (N_5216,N_1183,N_1779);
or U5217 (N_5217,N_3276,N_1802);
and U5218 (N_5218,N_2991,N_1839);
or U5219 (N_5219,N_2339,N_1284);
and U5220 (N_5220,N_4978,N_1587);
and U5221 (N_5221,N_3502,N_626);
and U5222 (N_5222,N_1443,N_3461);
and U5223 (N_5223,N_3590,N_3089);
nand U5224 (N_5224,N_3599,N_4855);
and U5225 (N_5225,N_3319,N_755);
nor U5226 (N_5226,N_3499,N_596);
nand U5227 (N_5227,N_4124,N_3858);
and U5228 (N_5228,N_245,N_1571);
nor U5229 (N_5229,N_2039,N_897);
and U5230 (N_5230,N_2769,N_3764);
and U5231 (N_5231,N_2986,N_47);
and U5232 (N_5232,N_4239,N_803);
nor U5233 (N_5233,N_3580,N_3996);
or U5234 (N_5234,N_1658,N_2643);
nor U5235 (N_5235,N_1705,N_3140);
xor U5236 (N_5236,N_356,N_3181);
and U5237 (N_5237,N_446,N_2617);
nor U5238 (N_5238,N_1820,N_3644);
or U5239 (N_5239,N_2305,N_1643);
nor U5240 (N_5240,N_4288,N_4211);
nor U5241 (N_5241,N_261,N_3921);
and U5242 (N_5242,N_1642,N_1714);
nand U5243 (N_5243,N_3949,N_2925);
nor U5244 (N_5244,N_3266,N_4453);
xor U5245 (N_5245,N_4002,N_4622);
or U5246 (N_5246,N_169,N_2247);
and U5247 (N_5247,N_1116,N_4524);
and U5248 (N_5248,N_431,N_3673);
and U5249 (N_5249,N_4436,N_925);
nand U5250 (N_5250,N_4236,N_1129);
xnor U5251 (N_5251,N_1659,N_4770);
nor U5252 (N_5252,N_1663,N_538);
and U5253 (N_5253,N_649,N_2846);
nand U5254 (N_5254,N_1633,N_452);
and U5255 (N_5255,N_2283,N_338);
nand U5256 (N_5256,N_279,N_1368);
nand U5257 (N_5257,N_519,N_2472);
and U5258 (N_5258,N_3719,N_2999);
nor U5259 (N_5259,N_3975,N_3474);
nor U5260 (N_5260,N_3261,N_4164);
nor U5261 (N_5261,N_903,N_1046);
and U5262 (N_5262,N_3086,N_1564);
and U5263 (N_5263,N_1098,N_3692);
or U5264 (N_5264,N_3784,N_3345);
xor U5265 (N_5265,N_2122,N_1634);
and U5266 (N_5266,N_3433,N_4362);
or U5267 (N_5267,N_2164,N_1708);
nor U5268 (N_5268,N_2424,N_4825);
nor U5269 (N_5269,N_4278,N_2021);
or U5270 (N_5270,N_3007,N_789);
xnor U5271 (N_5271,N_583,N_3093);
xnor U5272 (N_5272,N_1728,N_587);
and U5273 (N_5273,N_1442,N_4035);
nand U5274 (N_5274,N_3591,N_1666);
nand U5275 (N_5275,N_3449,N_3582);
and U5276 (N_5276,N_4749,N_2141);
and U5277 (N_5277,N_1335,N_2508);
nor U5278 (N_5278,N_2229,N_4205);
xnor U5279 (N_5279,N_530,N_2005);
nor U5280 (N_5280,N_1001,N_525);
nor U5281 (N_5281,N_309,N_3745);
or U5282 (N_5282,N_250,N_2126);
and U5283 (N_5283,N_3326,N_3436);
nor U5284 (N_5284,N_3448,N_4042);
or U5285 (N_5285,N_4678,N_3090);
or U5286 (N_5286,N_4930,N_4907);
xnor U5287 (N_5287,N_4146,N_2167);
nor U5288 (N_5288,N_2919,N_702);
nand U5289 (N_5289,N_3770,N_4084);
or U5290 (N_5290,N_4646,N_2244);
nor U5291 (N_5291,N_1108,N_4866);
nand U5292 (N_5292,N_1845,N_1718);
or U5293 (N_5293,N_973,N_1282);
or U5294 (N_5294,N_4346,N_3161);
nand U5295 (N_5295,N_1482,N_1573);
or U5296 (N_5296,N_593,N_160);
xnor U5297 (N_5297,N_3277,N_4270);
nand U5298 (N_5298,N_1467,N_2204);
nor U5299 (N_5299,N_3798,N_2490);
xor U5300 (N_5300,N_2045,N_2996);
nand U5301 (N_5301,N_3626,N_2366);
xor U5302 (N_5302,N_2470,N_2248);
xor U5303 (N_5303,N_878,N_537);
or U5304 (N_5304,N_3575,N_2297);
xnor U5305 (N_5305,N_800,N_4082);
and U5306 (N_5306,N_2063,N_3368);
or U5307 (N_5307,N_1979,N_2151);
and U5308 (N_5308,N_1601,N_4569);
xor U5309 (N_5309,N_3121,N_2013);
or U5310 (N_5310,N_4652,N_100);
nand U5311 (N_5311,N_3141,N_1441);
xor U5312 (N_5312,N_4242,N_4722);
xnor U5313 (N_5313,N_1305,N_3094);
and U5314 (N_5314,N_4452,N_2829);
nand U5315 (N_5315,N_4654,N_4843);
nor U5316 (N_5316,N_2093,N_2261);
nor U5317 (N_5317,N_1012,N_1017);
or U5318 (N_5318,N_2195,N_4257);
or U5319 (N_5319,N_27,N_3680);
or U5320 (N_5320,N_1330,N_2451);
and U5321 (N_5321,N_1648,N_3523);
nand U5322 (N_5322,N_3606,N_4018);
or U5323 (N_5323,N_2767,N_2721);
nand U5324 (N_5324,N_1502,N_3555);
or U5325 (N_5325,N_295,N_3199);
and U5326 (N_5326,N_1650,N_1300);
or U5327 (N_5327,N_2147,N_2552);
or U5328 (N_5328,N_4292,N_3934);
and U5329 (N_5329,N_85,N_46);
or U5330 (N_5330,N_2961,N_4120);
nand U5331 (N_5331,N_1626,N_4050);
and U5332 (N_5332,N_1733,N_421);
nor U5333 (N_5333,N_4244,N_1593);
nor U5334 (N_5334,N_438,N_3723);
xnor U5335 (N_5335,N_3785,N_1410);
and U5336 (N_5336,N_797,N_1892);
nand U5337 (N_5337,N_1085,N_3047);
or U5338 (N_5338,N_4751,N_560);
or U5339 (N_5339,N_992,N_809);
nand U5340 (N_5340,N_1987,N_4083);
or U5341 (N_5341,N_339,N_4984);
and U5342 (N_5342,N_4832,N_1421);
nor U5343 (N_5343,N_3338,N_1431);
or U5344 (N_5344,N_4550,N_3122);
or U5345 (N_5345,N_2635,N_1876);
nand U5346 (N_5346,N_4473,N_1499);
xnor U5347 (N_5347,N_362,N_2556);
xnor U5348 (N_5348,N_4690,N_2719);
nand U5349 (N_5349,N_2048,N_2353);
xnor U5350 (N_5350,N_2221,N_3927);
nand U5351 (N_5351,N_2421,N_3232);
xnor U5352 (N_5352,N_2764,N_3752);
and U5353 (N_5353,N_4336,N_4268);
nand U5354 (N_5354,N_3970,N_677);
nor U5355 (N_5355,N_3153,N_3835);
and U5356 (N_5356,N_4066,N_1881);
xor U5357 (N_5357,N_3540,N_2870);
or U5358 (N_5358,N_1008,N_1741);
nor U5359 (N_5359,N_2702,N_59);
and U5360 (N_5360,N_1662,N_3428);
xor U5361 (N_5361,N_4658,N_4241);
nand U5362 (N_5362,N_3894,N_4943);
or U5363 (N_5363,N_1693,N_251);
or U5364 (N_5364,N_4507,N_1292);
or U5365 (N_5365,N_2254,N_2257);
and U5366 (N_5366,N_3992,N_4047);
nor U5367 (N_5367,N_475,N_4886);
nor U5368 (N_5368,N_1113,N_4536);
nand U5369 (N_5369,N_3331,N_2436);
nor U5370 (N_5370,N_3691,N_824);
and U5371 (N_5371,N_1625,N_4932);
xor U5372 (N_5372,N_3912,N_2543);
nor U5373 (N_5373,N_752,N_3330);
and U5374 (N_5374,N_1263,N_1052);
and U5375 (N_5375,N_4673,N_466);
or U5376 (N_5376,N_2751,N_203);
and U5377 (N_5377,N_3639,N_622);
nor U5378 (N_5378,N_1090,N_4297);
nand U5379 (N_5379,N_4184,N_3076);
xnor U5380 (N_5380,N_262,N_3067);
and U5381 (N_5381,N_2346,N_4160);
nand U5382 (N_5382,N_3280,N_1320);
nand U5383 (N_5383,N_1749,N_3452);
and U5384 (N_5384,N_889,N_1840);
and U5385 (N_5385,N_3074,N_1457);
and U5386 (N_5386,N_2755,N_4666);
or U5387 (N_5387,N_181,N_4192);
xnor U5388 (N_5388,N_3113,N_819);
and U5389 (N_5389,N_1967,N_3092);
and U5390 (N_5390,N_1972,N_4528);
nand U5391 (N_5391,N_2185,N_2511);
xor U5392 (N_5392,N_3109,N_4393);
and U5393 (N_5393,N_2323,N_4183);
and U5394 (N_5394,N_2652,N_683);
xnor U5395 (N_5395,N_1037,N_4173);
or U5396 (N_5396,N_2783,N_2838);
nor U5397 (N_5397,N_3061,N_3198);
xnor U5398 (N_5398,N_3444,N_3359);
xor U5399 (N_5399,N_1460,N_4057);
xnor U5400 (N_5400,N_3944,N_3603);
nand U5401 (N_5401,N_3985,N_1337);
xnor U5402 (N_5402,N_558,N_3812);
nand U5403 (N_5403,N_3226,N_123);
and U5404 (N_5404,N_1799,N_2500);
and U5405 (N_5405,N_2604,N_4596);
nand U5406 (N_5406,N_3610,N_651);
and U5407 (N_5407,N_1206,N_1661);
and U5408 (N_5408,N_868,N_3042);
nand U5409 (N_5409,N_4323,N_3088);
nand U5410 (N_5410,N_1546,N_1585);
nor U5411 (N_5411,N_2300,N_1059);
nor U5412 (N_5412,N_1996,N_1725);
and U5413 (N_5413,N_717,N_2154);
xor U5414 (N_5414,N_4308,N_3584);
xnor U5415 (N_5415,N_66,N_1264);
and U5416 (N_5416,N_3201,N_2199);
xnor U5417 (N_5417,N_2690,N_1817);
or U5418 (N_5418,N_4090,N_2377);
or U5419 (N_5419,N_3458,N_96);
or U5420 (N_5420,N_4783,N_2747);
or U5421 (N_5421,N_460,N_3139);
nand U5422 (N_5422,N_978,N_2573);
nor U5423 (N_5423,N_244,N_4144);
or U5424 (N_5424,N_4014,N_3989);
or U5425 (N_5425,N_2549,N_324);
nor U5426 (N_5426,N_366,N_736);
xor U5427 (N_5427,N_4928,N_3839);
xnor U5428 (N_5428,N_52,N_1406);
or U5429 (N_5429,N_4623,N_1976);
nand U5430 (N_5430,N_2920,N_2541);
xnor U5431 (N_5431,N_2678,N_3533);
nand U5432 (N_5432,N_681,N_4950);
nand U5433 (N_5433,N_4639,N_1403);
and U5434 (N_5434,N_3952,N_1637);
nand U5435 (N_5435,N_204,N_1653);
nand U5436 (N_5436,N_449,N_747);
or U5437 (N_5437,N_2949,N_555);
and U5438 (N_5438,N_632,N_351);
or U5439 (N_5439,N_2197,N_4994);
nor U5440 (N_5440,N_2711,N_4139);
nor U5441 (N_5441,N_2621,N_3158);
or U5442 (N_5442,N_2822,N_2970);
and U5443 (N_5443,N_9,N_663);
or U5444 (N_5444,N_3933,N_539);
xnor U5445 (N_5445,N_4335,N_4321);
nand U5446 (N_5446,N_2560,N_4359);
nand U5447 (N_5447,N_1720,N_4204);
nand U5448 (N_5448,N_3288,N_4215);
nand U5449 (N_5449,N_4077,N_4221);
or U5450 (N_5450,N_1729,N_876);
nor U5451 (N_5451,N_3248,N_3369);
or U5452 (N_5452,N_1936,N_4589);
nand U5453 (N_5453,N_2149,N_4347);
nand U5454 (N_5454,N_3615,N_2833);
and U5455 (N_5455,N_2789,N_2688);
or U5456 (N_5456,N_2433,N_3901);
nand U5457 (N_5457,N_1011,N_2);
nor U5458 (N_5458,N_4026,N_4579);
nor U5459 (N_5459,N_4755,N_457);
and U5460 (N_5460,N_479,N_252);
xnor U5461 (N_5461,N_3668,N_1970);
nand U5462 (N_5462,N_4267,N_1822);
and U5463 (N_5463,N_2224,N_1818);
and U5464 (N_5464,N_1333,N_1266);
and U5465 (N_5465,N_3395,N_3394);
or U5466 (N_5466,N_2533,N_662);
and U5467 (N_5467,N_2044,N_782);
or U5468 (N_5468,N_2956,N_176);
nand U5469 (N_5469,N_4291,N_2774);
and U5470 (N_5470,N_1062,N_2333);
and U5471 (N_5471,N_4771,N_2354);
xnor U5472 (N_5472,N_419,N_2564);
xor U5473 (N_5473,N_4934,N_1730);
and U5474 (N_5474,N_4905,N_578);
xor U5475 (N_5475,N_2799,N_3824);
and U5476 (N_5476,N_2255,N_901);
nand U5477 (N_5477,N_678,N_3656);
nand U5478 (N_5478,N_4398,N_3375);
xnor U5479 (N_5479,N_2171,N_109);
nor U5480 (N_5480,N_3163,N_1139);
nor U5481 (N_5481,N_3546,N_1684);
nand U5482 (N_5482,N_1465,N_168);
nor U5483 (N_5483,N_4085,N_4817);
and U5484 (N_5484,N_1759,N_4485);
xor U5485 (N_5485,N_2757,N_2087);
or U5486 (N_5486,N_792,N_975);
or U5487 (N_5487,N_3791,N_2885);
xor U5488 (N_5488,N_4388,N_4285);
nor U5489 (N_5489,N_4478,N_2135);
nor U5490 (N_5490,N_2601,N_1630);
xor U5491 (N_5491,N_566,N_259);
nand U5492 (N_5492,N_1157,N_805);
nor U5493 (N_5493,N_3742,N_2152);
and U5494 (N_5494,N_4007,N_3435);
nor U5495 (N_5495,N_3757,N_2612);
nor U5496 (N_5496,N_319,N_1614);
xor U5497 (N_5497,N_1021,N_2442);
or U5498 (N_5498,N_3019,N_3134);
and U5499 (N_5499,N_4094,N_2536);
or U5500 (N_5500,N_510,N_3915);
nand U5501 (N_5501,N_3786,N_4899);
and U5502 (N_5502,N_1775,N_3);
nand U5503 (N_5503,N_3482,N_1926);
nor U5504 (N_5504,N_1954,N_3616);
or U5505 (N_5505,N_1853,N_444);
nor U5506 (N_5506,N_3982,N_4967);
or U5507 (N_5507,N_4716,N_4687);
xor U5508 (N_5508,N_1409,N_3309);
or U5509 (N_5509,N_822,N_2938);
or U5510 (N_5510,N_1356,N_2588);
xor U5511 (N_5511,N_2693,N_612);
and U5512 (N_5512,N_4792,N_2355);
nand U5513 (N_5513,N_608,N_67);
and U5514 (N_5514,N_3191,N_1141);
xnor U5515 (N_5515,N_1968,N_1918);
xnor U5516 (N_5516,N_703,N_2104);
nand U5517 (N_5517,N_3462,N_4078);
nand U5518 (N_5518,N_1338,N_562);
and U5519 (N_5519,N_2928,N_697);
nor U5520 (N_5520,N_4763,N_1171);
and U5521 (N_5521,N_2273,N_3801);
nand U5522 (N_5522,N_90,N_4391);
or U5523 (N_5523,N_661,N_4586);
or U5524 (N_5524,N_4600,N_2645);
nor U5525 (N_5525,N_3402,N_2924);
xnor U5526 (N_5526,N_2085,N_1701);
and U5527 (N_5527,N_1353,N_12);
or U5528 (N_5528,N_3020,N_2679);
and U5529 (N_5529,N_4809,N_1771);
and U5530 (N_5530,N_1462,N_3016);
nor U5531 (N_5531,N_911,N_869);
nor U5532 (N_5532,N_570,N_1915);
nand U5533 (N_5533,N_2659,N_3215);
and U5534 (N_5534,N_1680,N_2405);
or U5535 (N_5535,N_175,N_2667);
or U5536 (N_5536,N_3717,N_2069);
and U5537 (N_5537,N_1523,N_2426);
nand U5538 (N_5538,N_3298,N_2922);
xnor U5539 (N_5539,N_77,N_1578);
nor U5540 (N_5540,N_45,N_418);
and U5541 (N_5541,N_1010,N_2660);
or U5542 (N_5542,N_3734,N_3831);
nor U5543 (N_5543,N_3880,N_631);
nor U5544 (N_5544,N_995,N_826);
xnor U5545 (N_5545,N_2595,N_3891);
nand U5546 (N_5546,N_3953,N_2103);
nand U5547 (N_5547,N_2456,N_1265);
or U5548 (N_5548,N_44,N_3493);
xnor U5549 (N_5549,N_321,N_946);
or U5550 (N_5550,N_1254,N_4959);
and U5551 (N_5551,N_3632,N_665);
or U5552 (N_5552,N_108,N_3302);
and U5553 (N_5553,N_1553,N_1344);
nor U5554 (N_5554,N_2950,N_2656);
nand U5555 (N_5555,N_2279,N_104);
or U5556 (N_5556,N_2724,N_4003);
and U5557 (N_5557,N_3707,N_1543);
xnor U5558 (N_5558,N_659,N_417);
or U5559 (N_5559,N_4171,N_4256);
nand U5560 (N_5560,N_4314,N_71);
xnor U5561 (N_5561,N_523,N_364);
nor U5562 (N_5562,N_1993,N_556);
nand U5563 (N_5563,N_226,N_778);
nor U5564 (N_5564,N_2150,N_987);
xor U5565 (N_5565,N_386,N_368);
and U5566 (N_5566,N_4089,N_4027);
xnor U5567 (N_5567,N_4469,N_3164);
and U5568 (N_5568,N_186,N_3939);
and U5569 (N_5569,N_1770,N_4409);
nand U5570 (N_5570,N_4629,N_4744);
or U5571 (N_5571,N_1387,N_4299);
nand U5572 (N_5572,N_2114,N_4012);
nand U5573 (N_5573,N_1624,N_1132);
xnor U5574 (N_5574,N_2010,N_1755);
nor U5575 (N_5575,N_2998,N_821);
nor U5576 (N_5576,N_2600,N_3091);
xor U5577 (N_5577,N_3688,N_1557);
nor U5578 (N_5578,N_1363,N_1311);
xnor U5579 (N_5579,N_2850,N_675);
or U5580 (N_5580,N_1466,N_4683);
xor U5581 (N_5581,N_4675,N_522);
xor U5582 (N_5582,N_4503,N_4148);
or U5583 (N_5583,N_2812,N_2616);
and U5584 (N_5584,N_1734,N_3704);
xnor U5585 (N_5585,N_269,N_2012);
nor U5586 (N_5586,N_4540,N_4696);
nor U5587 (N_5587,N_1949,N_3977);
nand U5588 (N_5588,N_4892,N_696);
and U5589 (N_5589,N_1178,N_2675);
nand U5590 (N_5590,N_3250,N_3472);
nand U5591 (N_5591,N_1615,N_470);
nor U5592 (N_5592,N_3291,N_4838);
xnor U5593 (N_5593,N_2161,N_834);
and U5594 (N_5594,N_3887,N_2052);
or U5595 (N_5595,N_308,N_4814);
xor U5596 (N_5596,N_2669,N_815);
xor U5597 (N_5597,N_2071,N_916);
and U5598 (N_5598,N_4032,N_760);
nand U5599 (N_5599,N_1763,N_833);
xnor U5600 (N_5600,N_3385,N_2348);
and U5601 (N_5601,N_73,N_617);
nor U5602 (N_5602,N_102,N_756);
and U5603 (N_5603,N_1518,N_2329);
and U5604 (N_5604,N_1813,N_580);
or U5605 (N_5605,N_498,N_2580);
xor U5606 (N_5606,N_2821,N_1036);
nor U5607 (N_5607,N_3229,N_267);
or U5608 (N_5608,N_3657,N_4315);
or U5609 (N_5609,N_1904,N_3997);
and U5610 (N_5610,N_3648,N_1706);
or U5611 (N_5611,N_6,N_2640);
and U5612 (N_5612,N_4231,N_4461);
and U5613 (N_5613,N_4705,N_2548);
and U5614 (N_5614,N_4709,N_3649);
and U5615 (N_5615,N_4252,N_3501);
nand U5616 (N_5616,N_1057,N_2697);
and U5617 (N_5617,N_3034,N_3968);
xnor U5618 (N_5618,N_4208,N_2202);
nand U5619 (N_5619,N_4914,N_4577);
nor U5620 (N_5620,N_919,N_4213);
and U5621 (N_5621,N_3706,N_3984);
or U5622 (N_5622,N_1221,N_2502);
nor U5623 (N_5623,N_2529,N_2460);
and U5624 (N_5624,N_3478,N_1472);
nand U5625 (N_5625,N_1545,N_1020);
xnor U5626 (N_5626,N_1019,N_3183);
nor U5627 (N_5627,N_2140,N_4777);
and U5628 (N_5628,N_1745,N_4897);
and U5629 (N_5629,N_960,N_1408);
nor U5630 (N_5630,N_4472,N_2963);
nor U5631 (N_5631,N_623,N_1910);
xnor U5632 (N_5632,N_629,N_462);
nand U5633 (N_5633,N_4582,N_1592);
xnor U5634 (N_5634,N_3731,N_3442);
nor U5635 (N_5635,N_4490,N_467);
and U5636 (N_5636,N_2291,N_4826);
and U5637 (N_5637,N_32,N_201);
nand U5638 (N_5638,N_129,N_453);
xor U5639 (N_5639,N_4965,N_330);
and U5640 (N_5640,N_1023,N_1097);
xor U5641 (N_5641,N_166,N_3611);
xor U5642 (N_5642,N_748,N_1686);
and U5643 (N_5643,N_3322,N_491);
xnor U5644 (N_5644,N_2361,N_342);
or U5645 (N_5645,N_2537,N_1959);
or U5646 (N_5646,N_177,N_3940);
nand U5647 (N_5647,N_624,N_3315);
xnor U5648 (N_5648,N_4948,N_3110);
nand U5649 (N_5649,N_3307,N_2598);
nand U5650 (N_5650,N_4227,N_3525);
and U5651 (N_5651,N_2425,N_1257);
nand U5652 (N_5652,N_4367,N_208);
or U5653 (N_5653,N_4196,N_3592);
nor U5654 (N_5654,N_3397,N_1886);
and U5655 (N_5655,N_3180,N_4131);
nand U5656 (N_5656,N_2759,N_1999);
nand U5657 (N_5657,N_1893,N_4022);
or U5658 (N_5658,N_795,N_3029);
xor U5659 (N_5659,N_4671,N_3744);
nor U5660 (N_5660,N_3026,N_1126);
nor U5661 (N_5661,N_2705,N_4400);
and U5662 (N_5662,N_1252,N_4);
or U5663 (N_5663,N_4086,N_2519);
or U5664 (N_5664,N_2410,N_1095);
and U5665 (N_5665,N_1986,N_2428);
xor U5666 (N_5666,N_1493,N_1261);
xor U5667 (N_5667,N_4857,N_1677);
xnor U5668 (N_5668,N_2550,N_4791);
xor U5669 (N_5669,N_1177,N_271);
nor U5670 (N_5670,N_3655,N_1142);
nand U5671 (N_5671,N_2863,N_4561);
nor U5672 (N_5672,N_1672,N_3874);
nor U5673 (N_5673,N_2644,N_4127);
nand U5674 (N_5674,N_4944,N_4682);
nor U5675 (N_5675,N_3224,N_999);
xor U5676 (N_5676,N_3317,N_2450);
xnor U5677 (N_5677,N_1942,N_670);
or U5678 (N_5678,N_4719,N_1900);
and U5679 (N_5679,N_274,N_2193);
nor U5680 (N_5680,N_2284,N_2018);
nor U5681 (N_5681,N_4782,N_2454);
and U5682 (N_5682,N_404,N_1812);
or U5683 (N_5683,N_501,N_557);
and U5684 (N_5684,N_1689,N_4877);
nor U5685 (N_5685,N_4688,N_3299);
nor U5686 (N_5686,N_192,N_4405);
xnor U5687 (N_5687,N_811,N_4964);
xor U5688 (N_5688,N_4432,N_619);
xnor U5689 (N_5689,N_2877,N_3720);
nor U5690 (N_5690,N_3818,N_4445);
nand U5691 (N_5691,N_3936,N_3886);
and U5692 (N_5692,N_3822,N_4499);
and U5693 (N_5693,N_3925,N_4839);
and U5694 (N_5694,N_4456,N_4376);
or U5695 (N_5695,N_2658,N_3281);
nor U5696 (N_5696,N_373,N_3443);
xor U5697 (N_5697,N_349,N_2237);
and U5698 (N_5698,N_2347,N_473);
xor U5699 (N_5699,N_1199,N_2929);
xnor U5700 (N_5700,N_344,N_1245);
and U5701 (N_5701,N_11,N_3922);
nand U5702 (N_5702,N_2331,N_4302);
nand U5703 (N_5703,N_3270,N_4643);
xor U5704 (N_5704,N_1773,N_3412);
xor U5705 (N_5705,N_2754,N_4210);
nor U5706 (N_5706,N_952,N_3593);
or U5707 (N_5707,N_841,N_4565);
or U5708 (N_5708,N_2256,N_744);
nor U5709 (N_5709,N_1882,N_3220);
xnor U5710 (N_5710,N_1832,N_3516);
xor U5711 (N_5711,N_1323,N_118);
and U5712 (N_5712,N_1181,N_3926);
nor U5713 (N_5713,N_1032,N_866);
or U5714 (N_5714,N_2725,N_3498);
xor U5715 (N_5715,N_4860,N_699);
or U5716 (N_5716,N_282,N_4353);
nor U5717 (N_5717,N_4988,N_829);
nand U5718 (N_5718,N_4901,N_656);
and U5719 (N_5719,N_316,N_4097);
or U5720 (N_5720,N_2982,N_2089);
nand U5721 (N_5721,N_2271,N_357);
nor U5722 (N_5722,N_1489,N_1373);
nor U5723 (N_5723,N_4816,N_3131);
or U5724 (N_5724,N_2837,N_2127);
nor U5725 (N_5725,N_56,N_3604);
nor U5726 (N_5726,N_2748,N_3779);
xor U5727 (N_5727,N_477,N_48);
and U5728 (N_5728,N_3621,N_3529);
xor U5729 (N_5729,N_3179,N_904);
xnor U5730 (N_5730,N_3631,N_1451);
or U5731 (N_5731,N_2967,N_3082);
nor U5732 (N_5732,N_4356,N_3123);
nor U5733 (N_5733,N_630,N_1956);
nor U5734 (N_5734,N_1379,N_2220);
xnor U5735 (N_5735,N_1039,N_4721);
or U5736 (N_5736,N_1314,N_2239);
xor U5737 (N_5737,N_260,N_1374);
or U5738 (N_5738,N_2264,N_239);
and U5739 (N_5739,N_363,N_2058);
xnor U5740 (N_5740,N_367,N_2455);
nand U5741 (N_5741,N_2910,N_4296);
nand U5742 (N_5742,N_1836,N_427);
or U5743 (N_5743,N_4605,N_1595);
or U5744 (N_5744,N_1707,N_1160);
nor U5745 (N_5745,N_3025,N_2359);
nor U5746 (N_5746,N_1043,N_3233);
xnor U5747 (N_5747,N_153,N_4927);
or U5748 (N_5748,N_4437,N_283);
nor U5749 (N_5749,N_2142,N_4888);
or U5750 (N_5750,N_2097,N_891);
and U5751 (N_5751,N_74,N_4523);
or U5752 (N_5752,N_3379,N_2939);
and U5753 (N_5753,N_2209,N_2059);
xnor U5754 (N_5754,N_3166,N_1173);
or U5755 (N_5755,N_3380,N_1751);
nand U5756 (N_5756,N_2820,N_3227);
nor U5757 (N_5757,N_2976,N_2159);
or U5758 (N_5758,N_3396,N_1933);
nand U5759 (N_5759,N_155,N_4000);
nor U5760 (N_5760,N_4497,N_2174);
or U5761 (N_5761,N_3441,N_1727);
xnor U5762 (N_5762,N_1948,N_3490);
or U5763 (N_5763,N_4650,N_4081);
nor U5764 (N_5764,N_3962,N_2779);
or U5765 (N_5765,N_1217,N_257);
xor U5766 (N_5766,N_2423,N_2277);
and U5767 (N_5767,N_711,N_14);
nand U5768 (N_5768,N_965,N_4966);
nand U5769 (N_5769,N_2403,N_2872);
xnor U5770 (N_5770,N_407,N_434);
xor U5771 (N_5771,N_2873,N_2116);
nand U5772 (N_5772,N_4198,N_41);
and U5773 (N_5773,N_4151,N_1047);
and U5774 (N_5774,N_2917,N_4767);
nand U5775 (N_5775,N_2153,N_4667);
nand U5776 (N_5776,N_2406,N_4554);
and U5777 (N_5777,N_4822,N_3990);
nand U5778 (N_5778,N_2793,N_1475);
or U5779 (N_5779,N_3011,N_4365);
or U5780 (N_5780,N_4945,N_967);
nor U5781 (N_5781,N_1656,N_1874);
xnor U5782 (N_5782,N_4982,N_4617);
nor U5783 (N_5783,N_810,N_3554);
nand U5784 (N_5784,N_3146,N_72);
xor U5785 (N_5785,N_1715,N_899);
or U5786 (N_5786,N_600,N_1651);
or U5787 (N_5787,N_1975,N_3943);
and U5788 (N_5788,N_1509,N_492);
or U5789 (N_5789,N_648,N_1737);
or U5790 (N_5790,N_2434,N_4063);
and U5791 (N_5791,N_3618,N_4074);
nand U5792 (N_5792,N_4819,N_582);
nand U5793 (N_5793,N_1709,N_1829);
and U5794 (N_5794,N_3138,N_2886);
nor U5795 (N_5795,N_1760,N_4341);
or U5796 (N_5796,N_3312,N_405);
xnor U5797 (N_5797,N_3562,N_3646);
or U5798 (N_5798,N_2497,N_3169);
xor U5799 (N_5799,N_87,N_2483);
and U5800 (N_5800,N_2437,N_4849);
nor U5801 (N_5801,N_1858,N_1831);
nand U5802 (N_5802,N_3059,N_4804);
xnor U5803 (N_5803,N_2567,N_1084);
and U5804 (N_5804,N_2301,N_4232);
and U5805 (N_5805,N_1130,N_1241);
or U5806 (N_5806,N_2270,N_1732);
and U5807 (N_5807,N_3362,N_1497);
xnor U5808 (N_5808,N_2586,N_2014);
or U5809 (N_5809,N_2492,N_4059);
xor U5810 (N_5810,N_1947,N_2138);
nand U5811 (N_5811,N_1852,N_172);
nor U5812 (N_5812,N_1385,N_4853);
xor U5813 (N_5813,N_4941,N_2088);
nand U5814 (N_5814,N_3573,N_1731);
nor U5815 (N_5815,N_1149,N_3366);
nor U5816 (N_5816,N_2592,N_4812);
or U5817 (N_5817,N_4803,N_962);
or U5818 (N_5818,N_4450,N_4762);
or U5819 (N_5819,N_4800,N_463);
nor U5820 (N_5820,N_3545,N_4372);
nand U5821 (N_5821,N_1086,N_1963);
or U5822 (N_5822,N_101,N_709);
or U5823 (N_5823,N_286,N_3854);
nor U5824 (N_5824,N_4883,N_3100);
xor U5825 (N_5825,N_4209,N_1246);
nor U5826 (N_5826,N_3464,N_814);
or U5827 (N_5827,N_3861,N_2480);
or U5828 (N_5828,N_1285,N_390);
nor U5829 (N_5829,N_2054,N_388);
nand U5830 (N_5830,N_2412,N_2638);
nor U5831 (N_5831,N_4330,N_1654);
xor U5832 (N_5832,N_3409,N_2685);
or U5833 (N_5833,N_3844,N_2302);
and U5834 (N_5834,N_2095,N_3350);
nor U5835 (N_5835,N_3314,N_145);
and U5836 (N_5836,N_1617,N_2106);
and U5837 (N_5837,N_2234,N_1106);
nor U5838 (N_5838,N_2101,N_2290);
or U5839 (N_5839,N_3900,N_2634);
and U5840 (N_5840,N_1782,N_568);
or U5841 (N_5841,N_4194,N_403);
or U5842 (N_5842,N_2394,N_3205);
xor U5843 (N_5843,N_1810,N_2384);
xor U5844 (N_5844,N_920,N_3222);
nor U5845 (N_5845,N_3022,N_36);
or U5846 (N_5846,N_2311,N_2365);
nor U5847 (N_5847,N_2180,N_1331);
nor U5848 (N_5848,N_3783,N_1158);
and U5849 (N_5849,N_327,N_595);
nand U5850 (N_5850,N_3868,N_217);
nor U5851 (N_5851,N_4475,N_1550);
nor U5852 (N_5852,N_333,N_3347);
nand U5853 (N_5853,N_125,N_2923);
and U5854 (N_5854,N_1877,N_3775);
and U5855 (N_5855,N_1561,N_4802);
nor U5856 (N_5856,N_2896,N_4756);
nor U5857 (N_5857,N_2327,N_3830);
nand U5858 (N_5858,N_4724,N_3361);
or U5859 (N_5859,N_3301,N_1446);
nor U5860 (N_5860,N_1505,N_3009);
nor U5861 (N_5861,N_4043,N_4679);
nand U5862 (N_5862,N_30,N_116);
and U5863 (N_5863,N_4111,N_3814);
nor U5864 (N_5864,N_1104,N_2110);
nand U5865 (N_5865,N_4833,N_4092);
or U5866 (N_5866,N_2370,N_1004);
nand U5867 (N_5867,N_2163,N_680);
or U5868 (N_5868,N_1412,N_913);
or U5869 (N_5869,N_4939,N_4830);
nor U5870 (N_5870,N_645,N_2723);
or U5871 (N_5871,N_3388,N_2531);
and U5872 (N_5872,N_862,N_1906);
nand U5873 (N_5873,N_2299,N_4344);
and U5874 (N_5874,N_1053,N_1411);
nand U5875 (N_5875,N_2217,N_684);
and U5876 (N_5876,N_3421,N_2210);
and U5877 (N_5877,N_1835,N_3732);
xnor U5878 (N_5878,N_1163,N_2466);
nor U5879 (N_5879,N_4921,N_977);
xnor U5880 (N_5880,N_4636,N_1982);
xor U5881 (N_5881,N_532,N_1185);
xnor U5882 (N_5882,N_954,N_2727);
or U5883 (N_5883,N_472,N_2578);
and U5884 (N_5884,N_3756,N_2325);
and U5885 (N_5885,N_682,N_858);
or U5886 (N_5886,N_302,N_4435);
nor U5887 (N_5887,N_2722,N_1850);
nor U5888 (N_5888,N_4717,N_1416);
xor U5889 (N_5889,N_705,N_2429);
and U5890 (N_5890,N_2322,N_2332);
xor U5891 (N_5891,N_4850,N_2750);
nand U5892 (N_5892,N_3033,N_4193);
xor U5893 (N_5893,N_1247,N_2123);
nor U5894 (N_5894,N_361,N_3792);
xnor U5895 (N_5895,N_3043,N_990);
xor U5896 (N_5896,N_1212,N_4106);
nor U5897 (N_5897,N_2086,N_3260);
or U5898 (N_5898,N_4029,N_1153);
xor U5899 (N_5899,N_2320,N_2788);
xnor U5900 (N_5900,N_1568,N_4976);
xor U5901 (N_5901,N_2081,N_1131);
and U5902 (N_5902,N_1903,N_524);
nor U5903 (N_5903,N_432,N_1349);
nor U5904 (N_5904,N_3702,N_3833);
or U5905 (N_5905,N_1924,N_1977);
xor U5906 (N_5906,N_2687,N_4790);
nor U5907 (N_5907,N_3896,N_2358);
nand U5908 (N_5908,N_1598,N_4774);
nand U5909 (N_5909,N_2968,N_2570);
nor U5910 (N_5910,N_2546,N_3703);
and U5911 (N_5911,N_3928,N_563);
or U5912 (N_5912,N_801,N_3108);
nor U5913 (N_5913,N_3609,N_2488);
and U5914 (N_5914,N_490,N_3068);
xnor U5915 (N_5915,N_2853,N_3107);
nor U5916 (N_5916,N_906,N_136);
or U5917 (N_5917,N_2684,N_1944);
xnor U5918 (N_5918,N_1989,N_3660);
and U5919 (N_5919,N_786,N_4243);
nor U5920 (N_5920,N_1583,N_2420);
xnor U5921 (N_5921,N_2814,N_1594);
xor U5922 (N_5922,N_3675,N_4985);
and U5923 (N_5923,N_1514,N_2031);
and U5924 (N_5924,N_3827,N_2744);
nor U5925 (N_5925,N_1280,N_1767);
and U5926 (N_5926,N_3787,N_485);
nand U5927 (N_5927,N_1362,N_2269);
and U5928 (N_5928,N_396,N_4451);
nor U5929 (N_5929,N_2115,N_933);
nor U5930 (N_5930,N_3400,N_2804);
xor U5931 (N_5931,N_4794,N_3754);
xnor U5932 (N_5932,N_2983,N_2033);
and U5933 (N_5933,N_2518,N_2268);
nor U5934 (N_5934,N_329,N_1951);
nand U5935 (N_5935,N_3382,N_320);
xor U5936 (N_5936,N_4143,N_465);
nand U5937 (N_5937,N_2532,N_2413);
and U5938 (N_5938,N_178,N_708);
xor U5939 (N_5939,N_4882,N_4240);
nand U5940 (N_5940,N_4560,N_3054);
nor U5941 (N_5941,N_3677,N_266);
nand U5942 (N_5942,N_4474,N_3200);
nor U5943 (N_5943,N_1640,N_3151);
xor U5944 (N_5944,N_569,N_2609);
and U5945 (N_5945,N_480,N_3729);
and U5946 (N_5946,N_3678,N_1586);
nor U5947 (N_5947,N_2047,N_416);
and U5948 (N_5948,N_781,N_1971);
or U5949 (N_5949,N_3543,N_2565);
and U5950 (N_5950,N_2554,N_7);
and U5951 (N_5951,N_1478,N_3457);
or U5952 (N_5952,N_2887,N_2430);
nand U5953 (N_5953,N_4181,N_3696);
nand U5954 (N_5954,N_718,N_278);
and U5955 (N_5955,N_4591,N_4571);
xor U5956 (N_5956,N_1962,N_1503);
xor U5957 (N_5957,N_4510,N_3308);
or U5958 (N_5958,N_512,N_1242);
nor U5959 (N_5959,N_3885,N_3144);
and U5960 (N_5960,N_4797,N_3849);
or U5961 (N_5961,N_3095,N_4179);
nand U5962 (N_5962,N_1602,N_2915);
nand U5963 (N_5963,N_2628,N_4222);
or U5964 (N_5964,N_2651,N_2371);
nand U5965 (N_5965,N_4319,N_843);
or U5966 (N_5966,N_4604,N_741);
xor U5967 (N_5967,N_4266,N_1075);
xor U5968 (N_5968,N_2065,N_3902);
or U5969 (N_5969,N_4433,N_1234);
xnor U5970 (N_5970,N_4895,N_2238);
or U5971 (N_5971,N_1118,N_2316);
or U5972 (N_5972,N_552,N_3878);
nand U5973 (N_5973,N_1830,N_179);
nand U5974 (N_5974,N_2899,N_4006);
nor U5975 (N_5975,N_1682,N_3578);
or U5976 (N_5976,N_3081,N_3404);
xnor U5977 (N_5977,N_3537,N_4033);
xnor U5978 (N_5978,N_2073,N_2479);
nand U5979 (N_5979,N_2078,N_4504);
nor U5980 (N_5980,N_3320,N_1367);
or U5981 (N_5981,N_2797,N_1710);
xnor U5982 (N_5982,N_4929,N_326);
xor U5983 (N_5983,N_3268,N_1480);
xor U5984 (N_5984,N_1286,N_4546);
or U5985 (N_5985,N_4884,N_3530);
nor U5986 (N_5986,N_3053,N_1110);
nand U5987 (N_5987,N_2109,N_4431);
nand U5988 (N_5988,N_15,N_1051);
nand U5989 (N_5989,N_4410,N_3557);
nand U5990 (N_5990,N_3296,N_62);
nor U5991 (N_5991,N_4995,N_707);
and U5992 (N_5992,N_1372,N_1880);
nand U5993 (N_5993,N_437,N_674);
and U5994 (N_5994,N_701,N_1952);
nand U5995 (N_5995,N_2825,N_2646);
or U5996 (N_5996,N_3202,N_76);
nor U5997 (N_5997,N_1612,N_4689);
nand U5998 (N_5998,N_1359,N_3242);
and U5999 (N_5999,N_313,N_917);
xnor U6000 (N_6000,N_3194,N_391);
nor U6001 (N_6001,N_3777,N_4021);
and U6002 (N_6002,N_1512,N_3566);
nor U6003 (N_6003,N_185,N_4037);
xor U6004 (N_6004,N_4466,N_788);
or U6005 (N_6005,N_2121,N_372);
nand U6006 (N_6006,N_1860,N_4394);
nand U6007 (N_6007,N_106,N_1237);
or U6008 (N_6008,N_315,N_853);
or U6009 (N_6009,N_3710,N_1259);
xor U6010 (N_6010,N_4087,N_1137);
nor U6011 (N_6011,N_1769,N_884);
nor U6012 (N_6012,N_2098,N_4494);
or U6013 (N_6013,N_2944,N_2249);
or U6014 (N_6014,N_1746,N_216);
and U6015 (N_6015,N_606,N_3741);
nor U6016 (N_6016,N_3055,N_4119);
xor U6017 (N_6017,N_615,N_719);
nor U6018 (N_6018,N_759,N_2182);
nand U6019 (N_6019,N_2025,N_4655);
nand U6020 (N_6020,N_3586,N_2927);
or U6021 (N_6021,N_4130,N_4185);
or U6022 (N_6022,N_2892,N_970);
nand U6023 (N_6023,N_2664,N_3841);
nor U6024 (N_6024,N_167,N_1427);
nand U6025 (N_6025,N_1394,N_408);
xor U6026 (N_6026,N_1766,N_1793);
and U6027 (N_6027,N_1081,N_4906);
and U6028 (N_6028,N_4327,N_688);
xnor U6029 (N_6029,N_1101,N_1795);
and U6030 (N_6030,N_3075,N_1554);
or U6031 (N_6031,N_3736,N_4624);
nor U6032 (N_6032,N_3105,N_844);
and U6033 (N_6033,N_2794,N_2622);
nand U6034 (N_6034,N_1078,N_4251);
xor U6035 (N_6035,N_1029,N_3860);
or U6036 (N_6036,N_2181,N_1805);
nor U6037 (N_6037,N_2287,N_447);
or U6038 (N_6038,N_4858,N_423);
nor U6039 (N_6039,N_1366,N_4703);
nand U6040 (N_6040,N_1496,N_3475);
nand U6041 (N_6041,N_218,N_3489);
xnor U6042 (N_6042,N_1226,N_4161);
and U6043 (N_6043,N_4295,N_1041);
nand U6044 (N_6044,N_2626,N_3204);
xor U6045 (N_6045,N_1649,N_2051);
xor U6046 (N_6046,N_2452,N_949);
xor U6047 (N_6047,N_2285,N_2443);
nand U6048 (N_6048,N_1821,N_4427);
xnor U6049 (N_6049,N_3851,N_4887);
or U6050 (N_6050,N_2773,N_1483);
nor U6051 (N_6051,N_3955,N_909);
and U6052 (N_6052,N_4136,N_825);
nand U6053 (N_6053,N_69,N_3799);
and U6054 (N_6054,N_616,N_4535);
nor U6055 (N_6055,N_3355,N_881);
or U6056 (N_6056,N_1000,N_4305);
nand U6057 (N_6057,N_1469,N_1145);
or U6058 (N_6058,N_3959,N_1190);
or U6059 (N_6059,N_4827,N_2619);
xor U6060 (N_6060,N_4317,N_3349);
nand U6061 (N_6061,N_3693,N_318);
xor U6062 (N_6062,N_2921,N_2194);
xor U6063 (N_6063,N_932,N_183);
xor U6064 (N_6064,N_2446,N_2303);
xor U6065 (N_6065,N_2187,N_2259);
or U6066 (N_6066,N_4926,N_2189);
nand U6067 (N_6067,N_2596,N_3002);
or U6068 (N_6068,N_2400,N_2233);
nor U6069 (N_6069,N_1308,N_3348);
and U6070 (N_6070,N_195,N_1953);
or U6071 (N_6071,N_2615,N_2916);
and U6072 (N_6072,N_91,N_2906);
nand U6073 (N_6073,N_4429,N_1898);
nand U6074 (N_6074,N_2666,N_3802);
xor U6075 (N_6075,N_574,N_1031);
nand U6076 (N_6076,N_4810,N_1056);
nand U6077 (N_6077,N_764,N_3589);
nor U6078 (N_6078,N_2739,N_2002);
and U6079 (N_6079,N_1833,N_2655);
or U6080 (N_6080,N_3807,N_4660);
nor U6081 (N_6081,N_2542,N_3013);
nor U6082 (N_6082,N_918,N_1393);
or U6083 (N_6083,N_4038,N_604);
and U6084 (N_6084,N_1974,N_1847);
nand U6085 (N_6085,N_1238,N_2388);
and U6086 (N_6086,N_3875,N_1940);
xor U6087 (N_6087,N_2262,N_398);
xnor U6088 (N_6088,N_1350,N_3569);
nand U6089 (N_6089,N_1878,N_4152);
nor U6090 (N_6090,N_585,N_1447);
nor U6091 (N_6091,N_852,N_37);
nor U6092 (N_6092,N_773,N_1283);
and U6093 (N_6093,N_1608,N_4720);
or U6094 (N_6094,N_2293,N_439);
nor U6095 (N_6095,N_528,N_1291);
and U6096 (N_6096,N_4951,N_554);
nor U6097 (N_6097,N_3186,N_3049);
xnor U6098 (N_6098,N_2240,N_2493);
or U6099 (N_6099,N_3681,N_542);
nand U6100 (N_6100,N_1487,N_1490);
xor U6101 (N_6101,N_3271,N_2390);
nor U6102 (N_6102,N_854,N_3192);
xor U6103 (N_6103,N_82,N_4390);
nor U6104 (N_6104,N_1863,N_1360);
and U6105 (N_6105,N_499,N_3684);
and U6106 (N_6106,N_2540,N_669);
nor U6107 (N_6107,N_2683,N_2060);
nand U6108 (N_6108,N_2844,N_110);
nor U6109 (N_6109,N_4313,N_3815);
nor U6110 (N_6110,N_4909,N_2624);
xor U6111 (N_6111,N_2419,N_745);
nor U6112 (N_6112,N_4733,N_79);
and U6113 (N_6113,N_4448,N_937);
xor U6114 (N_6114,N_2330,N_211);
nand U6115 (N_6115,N_1842,N_1670);
or U6116 (N_6116,N_4845,N_3148);
xor U6117 (N_6117,N_2708,N_1866);
nand U6118 (N_6118,N_4608,N_4781);
xor U6119 (N_6119,N_2545,N_1629);
nand U6120 (N_6120,N_4403,N_2505);
nor U6121 (N_6121,N_738,N_382);
xnor U6122 (N_6122,N_4073,N_4805);
xnor U6123 (N_6123,N_4118,N_2781);
nor U6124 (N_6124,N_1434,N_4468);
nand U6125 (N_6125,N_2791,N_3104);
or U6126 (N_6126,N_4583,N_4740);
nand U6127 (N_6127,N_2686,N_2513);
or U6128 (N_6128,N_3195,N_981);
and U6129 (N_6129,N_731,N_3782);
or U6130 (N_6130,N_4495,N_3788);
or U6131 (N_6131,N_4754,N_3155);
nor U6132 (N_6132,N_4199,N_2294);
xor U6133 (N_6133,N_2128,N_2874);
xnor U6134 (N_6134,N_1555,N_2842);
nand U6135 (N_6135,N_20,N_2817);
nand U6136 (N_6136,N_2473,N_2942);
and U6137 (N_6137,N_685,N_2292);
xor U6138 (N_6138,N_2932,N_164);
and U6139 (N_6139,N_1211,N_496);
nand U6140 (N_6140,N_42,N_325);
xnor U6141 (N_6141,N_3560,N_3399);
nor U6142 (N_6142,N_3041,N_2000);
or U6143 (N_6143,N_4041,N_1096);
nor U6144 (N_6144,N_247,N_4274);
or U6145 (N_6145,N_3506,N_1792);
or U6146 (N_6146,N_2823,N_4521);
nand U6147 (N_6147,N_322,N_3438);
xor U6148 (N_6148,N_758,N_3931);
xor U6149 (N_6149,N_2649,N_2099);
xor U6150 (N_6150,N_3813,N_307);
nor U6151 (N_6151,N_4389,N_4692);
or U6152 (N_6152,N_4732,N_291);
nand U6153 (N_6153,N_1925,N_3207);
or U6154 (N_6154,N_2030,N_4873);
nor U6155 (N_6155,N_785,N_331);
and U6156 (N_6156,N_2509,N_4894);
nor U6157 (N_6157,N_1354,N_2859);
nor U6158 (N_6158,N_4366,N_4971);
nor U6159 (N_6159,N_3130,N_1794);
and U6160 (N_6160,N_3243,N_4920);
or U6161 (N_6161,N_3328,N_2937);
and U6162 (N_6162,N_531,N_3285);
nand U6163 (N_6163,N_265,N_4182);
xor U6164 (N_6164,N_1997,N_4272);
or U6165 (N_6165,N_1440,N_137);
or U6166 (N_6166,N_941,N_1576);
or U6167 (N_6167,N_695,N_2780);
and U6168 (N_6168,N_1574,N_1641);
nor U6169 (N_6169,N_4289,N_3037);
xor U6170 (N_6170,N_2514,N_1533);
and U6171 (N_6171,N_3340,N_2745);
nor U6172 (N_6172,N_4933,N_1510);
nand U6173 (N_6173,N_2211,N_4345);
nand U6174 (N_6174,N_4122,N_2286);
and U6175 (N_6175,N_1146,N_4706);
nor U6176 (N_6176,N_2011,N_1690);
xnor U6177 (N_6177,N_4506,N_2296);
nand U6178 (N_6178,N_3842,N_724);
or U6179 (N_6179,N_2691,N_350);
or U6180 (N_6180,N_371,N_3103);
xor U6181 (N_6181,N_2402,N_4138);
xor U6182 (N_6182,N_75,N_1674);
xor U6183 (N_6183,N_2761,N_4374);
nor U6184 (N_6184,N_4045,N_1589);
nand U6185 (N_6185,N_3221,N_2528);
and U6186 (N_6186,N_2313,N_4020);
nor U6187 (N_6187,N_963,N_1340);
nor U6188 (N_6188,N_4910,N_3162);
nor U6189 (N_6189,N_127,N_230);
or U6190 (N_6190,N_1120,N_1486);
nor U6191 (N_6191,N_1558,N_1937);
or U6192 (N_6192,N_2639,N_1932);
or U6193 (N_6193,N_2740,N_3267);
nand U6194 (N_6194,N_142,N_2599);
nor U6195 (N_6195,N_3663,N_1541);
and U6196 (N_6196,N_2334,N_2650);
nor U6197 (N_6197,N_3583,N_1599);
or U6198 (N_6198,N_2964,N_4656);
nor U6199 (N_6199,N_3120,N_2965);
xnor U6200 (N_6200,N_3467,N_839);
xor U6201 (N_6201,N_4219,N_117);
xnor U6202 (N_6202,N_2935,N_4156);
and U6203 (N_6203,N_1864,N_2913);
and U6204 (N_6204,N_2633,N_1088);
nor U6205 (N_6205,N_1889,N_3697);
and U6206 (N_6206,N_149,N_2737);
and U6207 (N_6207,N_4891,N_1208);
or U6208 (N_6208,N_548,N_1426);
and U6209 (N_6209,N_4135,N_2317);
xor U6210 (N_6210,N_873,N_4114);
xnor U6211 (N_6211,N_3283,N_2112);
nand U6212 (N_6212,N_3666,N_594);
and U6213 (N_6213,N_415,N_4363);
nand U6214 (N_6214,N_3341,N_3427);
and U6215 (N_6215,N_2816,N_4108);
nand U6216 (N_6216,N_817,N_4936);
nor U6217 (N_6217,N_934,N_2040);
or U6218 (N_6218,N_4316,N_1445);
and U6219 (N_6219,N_883,N_140);
nor U6220 (N_6220,N_605,N_3456);
nor U6221 (N_6221,N_3329,N_4752);
nor U6222 (N_6222,N_2266,N_4595);
nand U6223 (N_6223,N_3714,N_4290);
nor U6224 (N_6224,N_725,N_1328);
nor U6225 (N_6225,N_1375,N_3469);
nor U6226 (N_6226,N_476,N_3126);
xor U6227 (N_6227,N_3219,N_588);
or U6228 (N_6228,N_4580,N_3503);
nor U6229 (N_6229,N_3415,N_1606);
nand U6230 (N_6230,N_3553,N_128);
nand U6231 (N_6231,N_3625,N_3420);
or U6232 (N_6232,N_3494,N_392);
and U6233 (N_6233,N_2847,N_3156);
xnor U6234 (N_6234,N_277,N_2807);
nor U6235 (N_6235,N_2155,N_1600);
or U6236 (N_6236,N_3923,N_4067);
nand U6237 (N_6237,N_1563,N_3237);
and U6238 (N_6238,N_3513,N_666);
or U6239 (N_6239,N_4913,N_943);
nor U6240 (N_6240,N_4870,N_3670);
and U6241 (N_6241,N_3690,N_2858);
or U6242 (N_6242,N_4915,N_84);
nor U6243 (N_6243,N_3811,N_1310);
xor U6244 (N_6244,N_2524,N_1380);
nor U6245 (N_6245,N_4975,N_4842);
and U6246 (N_6246,N_2758,N_1289);
nand U6247 (N_6247,N_715,N_4530);
and U6248 (N_6248,N_779,N_3548);
xnor U6249 (N_6249,N_2985,N_3999);
nor U6250 (N_6250,N_1454,N_1644);
or U6251 (N_6251,N_2843,N_2875);
xor U6252 (N_6252,N_1439,N_743);
xor U6253 (N_6253,N_888,N_1297);
and U6254 (N_6254,N_4538,N_3008);
nor U6255 (N_6255,N_1702,N_515);
nor U6256 (N_6256,N_4626,N_2343);
xnor U6257 (N_6257,N_1908,N_2977);
xnor U6258 (N_6258,N_686,N_4568);
and U6259 (N_6259,N_3913,N_2868);
and U6260 (N_6260,N_4727,N_1067);
or U6261 (N_6261,N_2125,N_2803);
or U6262 (N_6262,N_2698,N_3304);
nor U6263 (N_6263,N_4786,N_1616);
nand U6264 (N_6264,N_4900,N_242);
nand U6265 (N_6265,N_1318,N_4864);
and U6266 (N_6266,N_1223,N_3476);
nor U6267 (N_6267,N_2557,N_236);
xor U6268 (N_6268,N_246,N_2482);
nand U6269 (N_6269,N_1919,N_4355);
nor U6270 (N_6270,N_1797,N_4375);
nand U6271 (N_6271,N_3871,N_3147);
and U6272 (N_6272,N_4772,N_3774);
or U6273 (N_6273,N_4065,N_988);
and U6274 (N_6274,N_3658,N_3898);
xor U6275 (N_6275,N_2696,N_4331);
nand U6276 (N_6276,N_2763,N_2074);
and U6277 (N_6277,N_982,N_2337);
xor U6278 (N_6278,N_359,N_474);
nor U6279 (N_6279,N_2631,N_3524);
and U6280 (N_6280,N_4324,N_1006);
or U6281 (N_6281,N_1418,N_4969);
xnor U6282 (N_6282,N_1198,N_507);
nand U6283 (N_6283,N_4686,N_4711);
and U6284 (N_6284,N_4699,N_1444);
nand U6285 (N_6285,N_516,N_2465);
nor U6286 (N_6286,N_3507,N_3892);
nor U6287 (N_6287,N_4493,N_3236);
xnor U6288 (N_6288,N_3893,N_2132);
nor U6289 (N_6289,N_4881,N_383);
and U6290 (N_6290,N_3111,N_4230);
nor U6291 (N_6291,N_3574,N_43);
xor U6292 (N_6292,N_3679,N_2813);
nor U6293 (N_6293,N_1521,N_314);
nor U6294 (N_6294,N_3414,N_2694);
xnor U6295 (N_6295,N_2117,N_4957);
nor U6296 (N_6296,N_1182,N_2022);
xor U6297 (N_6297,N_2735,N_3012);
or U6298 (N_6298,N_667,N_3571);
or U6299 (N_6299,N_2260,N_3235);
or U6300 (N_6300,N_607,N_4349);
xor U6301 (N_6301,N_3730,N_706);
xnor U6302 (N_6302,N_2538,N_4259);
and U6303 (N_6303,N_750,N_1694);
nand U6304 (N_6304,N_4922,N_1244);
nand U6305 (N_6305,N_1003,N_1687);
xor U6306 (N_6306,N_3410,N_545);
or U6307 (N_6307,N_2941,N_2815);
xor U6308 (N_6308,N_5,N_428);
nand U6309 (N_6309,N_2225,N_1220);
nand U6310 (N_6310,N_3051,N_4277);
xnor U6311 (N_6311,N_1776,N_646);
nand U6312 (N_6312,N_1425,N_28);
nor U6313 (N_6313,N_3969,N_1894);
or U6314 (N_6314,N_2170,N_1887);
nor U6315 (N_6315,N_1610,N_4896);
or U6316 (N_6316,N_1432,N_3313);
or U6317 (N_6317,N_3173,N_4852);
nor U6318 (N_6318,N_2278,N_4516);
and U6319 (N_6319,N_4539,N_3769);
and U6320 (N_6320,N_2795,N_337);
nand U6321 (N_6321,N_3517,N_3003);
and U6322 (N_6322,N_2023,N_2953);
nand U6323 (N_6323,N_3995,N_3740);
nor U6324 (N_6324,N_2094,N_550);
and U6325 (N_6325,N_2712,N_1248);
nand U6326 (N_6326,N_3597,N_4512);
nand U6327 (N_6327,N_1801,N_939);
xor U6328 (N_6328,N_2057,N_2139);
and U6329 (N_6329,N_3746,N_2258);
nor U6330 (N_6330,N_78,N_1990);
xor U6331 (N_6331,N_1392,N_2042);
nor U6332 (N_6332,N_2381,N_2515);
nor U6333 (N_6333,N_3834,N_2046);
nand U6334 (N_6334,N_4735,N_3115);
and U6335 (N_6335,N_1195,N_2061);
nor U6336 (N_6336,N_3136,N_3079);
and U6337 (N_6337,N_221,N_1239);
nand U6338 (N_6338,N_38,N_2608);
nand U6339 (N_6339,N_2796,N_4502);
nand U6340 (N_6340,N_1984,N_1202);
and U6341 (N_6341,N_61,N_3947);
or U6342 (N_6342,N_130,N_3978);
xor U6343 (N_6343,N_1365,N_3440);
nand U6344 (N_6344,N_4684,N_1897);
or U6345 (N_6345,N_2275,N_2307);
or U6346 (N_6346,N_3505,N_1218);
and U6347 (N_6347,N_1295,N_922);
nor U6348 (N_6348,N_4924,N_2801);
xor U6349 (N_6349,N_436,N_288);
and U6350 (N_6350,N_3335,N_3231);
or U6351 (N_6351,N_790,N_1632);
xnor U6352 (N_6352,N_210,N_936);
and U6353 (N_6353,N_126,N_2625);
and U6354 (N_6354,N_4854,N_694);
and U6355 (N_6355,N_1276,N_4076);
nor U6356 (N_6356,N_3439,N_4195);
nor U6357 (N_6357,N_1995,N_2775);
nand U6358 (N_6358,N_3845,N_1450);
or U6359 (N_6359,N_51,N_370);
or U6360 (N_6360,N_1184,N_4415);
and U6361 (N_6361,N_4486,N_26);
and U6362 (N_6362,N_1312,N_393);
or U6363 (N_6363,N_4379,N_2373);
xnor U6364 (N_6364,N_328,N_3066);
nor U6365 (N_6365,N_4465,N_1115);
nand U6366 (N_6366,N_2629,N_3453);
nor U6367 (N_6367,N_4309,N_1313);
xor U6368 (N_6368,N_4300,N_3087);
xnor U6369 (N_6369,N_808,N_248);
nand U6370 (N_6370,N_910,N_4633);
nor U6371 (N_6371,N_894,N_4492);
xnor U6372 (N_6372,N_2904,N_3759);
nand U6373 (N_6373,N_1696,N_2215);
or U6374 (N_6374,N_2111,N_93);
nand U6375 (N_6375,N_1549,N_802);
nand U6376 (N_6376,N_4430,N_424);
or U6377 (N_6377,N_1269,N_2491);
nand U6378 (N_6378,N_882,N_2971);
and U6379 (N_6379,N_1532,N_4955);
and U6380 (N_6380,N_2980,N_3228);
and U6381 (N_6381,N_2186,N_401);
and U6382 (N_6382,N_628,N_3819);
and U6383 (N_6383,N_2250,N_264);
and U6384 (N_6384,N_1,N_1143);
nand U6385 (N_6385,N_966,N_767);
nand U6386 (N_6386,N_551,N_2092);
nand U6387 (N_6387,N_1916,N_4694);
nor U6388 (N_6388,N_4477,N_1870);
xnor U6389 (N_6389,N_1713,N_4378);
xor U6390 (N_6390,N_3983,N_2477);
or U6391 (N_6391,N_968,N_2427);
nand U6392 (N_6392,N_4387,N_1268);
or U6393 (N_6393,N_2369,N_2253);
nor U6394 (N_6394,N_2975,N_3667);
xor U6395 (N_6395,N_1207,N_2729);
nand U6396 (N_6396,N_735,N_1214);
nor U6397 (N_6397,N_4416,N_1007);
nand U6398 (N_6398,N_3976,N_3069);
nor U6399 (N_6399,N_1645,N_25);
and U6400 (N_6400,N_4402,N_4049);
or U6401 (N_6401,N_2681,N_3294);
and U6402 (N_6402,N_2902,N_4237);
nor U6403 (N_6403,N_1048,N_400);
nor U6404 (N_6404,N_4011,N_2530);
or U6405 (N_6405,N_420,N_4594);
or U6406 (N_6406,N_1231,N_4903);
and U6407 (N_6407,N_4835,N_746);
or U6408 (N_6408,N_4056,N_2321);
or U6409 (N_6409,N_55,N_1657);
xnor U6410 (N_6410,N_3608,N_1811);
or U6411 (N_6411,N_3998,N_4867);
nor U6412 (N_6412,N_1203,N_4069);
nor U6413 (N_6413,N_4520,N_3118);
xor U6414 (N_6414,N_1695,N_3132);
nor U6415 (N_6415,N_726,N_4129);
nand U6416 (N_6416,N_4310,N_4031);
and U6417 (N_6417,N_1929,N_2387);
or U6418 (N_6418,N_1824,N_4109);
nand U6419 (N_6419,N_4408,N_478);
or U6420 (N_6420,N_1913,N_4665);
nor U6421 (N_6421,N_2133,N_1250);
xor U6422 (N_6422,N_2736,N_4200);
xor U6423 (N_6423,N_893,N_3425);
and U6424 (N_6424,N_4368,N_2265);
or U6425 (N_6425,N_3856,N_335);
nor U6426 (N_6426,N_993,N_3333);
nand U6427 (N_6427,N_3295,N_4861);
xnor U6428 (N_6428,N_225,N_4028);
nand U6429 (N_6429,N_1530,N_3908);
and U6430 (N_6430,N_2699,N_2184);
nand U6431 (N_6431,N_4224,N_4294);
xnor U6432 (N_6432,N_3119,N_4228);
or U6433 (N_6433,N_4166,N_3522);
or U6434 (N_6434,N_1704,N_4592);
nor U6435 (N_6435,N_4265,N_3431);
xnor U6436 (N_6436,N_3598,N_4742);
nand U6437 (N_6437,N_2841,N_4820);
xor U6438 (N_6438,N_4008,N_2576);
and U6439 (N_6439,N_590,N_1196);
nand U6440 (N_6440,N_1204,N_298);
and U6441 (N_6441,N_182,N_2743);
xor U6442 (N_6442,N_1960,N_1798);
or U6443 (N_6443,N_1136,N_1309);
and U6444 (N_6444,N_2717,N_1205);
xor U6445 (N_6445,N_4635,N_3674);
xnor U6446 (N_6446,N_1147,N_358);
and U6447 (N_6447,N_4868,N_3620);
nand U6448 (N_6448,N_2157,N_4333);
nor U6449 (N_6449,N_2654,N_4865);
nand U6450 (N_6450,N_875,N_1415);
and U6451 (N_6451,N_4603,N_2338);
and U6452 (N_6452,N_4534,N_353);
or U6453 (N_6453,N_1188,N_1089);
and U6454 (N_6454,N_4384,N_2898);
xor U6455 (N_6455,N_2969,N_3036);
nand U6456 (N_6456,N_1540,N_4620);
nand U6457 (N_6457,N_3353,N_3904);
nand U6458 (N_6458,N_2341,N_2368);
nor U6459 (N_6459,N_1369,N_1024);
nand U6460 (N_6460,N_1159,N_1570);
nand U6461 (N_6461,N_1389,N_263);
and U6462 (N_6462,N_2589,N_1827);
nand U6463 (N_6463,N_134,N_3336);
xor U6464 (N_6464,N_4385,N_3255);
or U6465 (N_6465,N_4382,N_4664);
or U6466 (N_6466,N_2880,N_2520);
nor U6467 (N_6467,N_1526,N_820);
or U6468 (N_6468,N_3895,N_3334);
nand U6469 (N_6469,N_4602,N_2597);
and U6470 (N_6470,N_1869,N_3032);
nand U6471 (N_6471,N_1895,N_1172);
xnor U6472 (N_6472,N_3470,N_3986);
or U6473 (N_6473,N_3403,N_1872);
or U6474 (N_6474,N_4736,N_1319);
nand U6475 (N_6475,N_1459,N_3567);
or U6476 (N_6476,N_3184,N_2584);
or U6477 (N_6477,N_4961,N_4869);
and U6478 (N_6478,N_923,N_80);
or U6479 (N_6479,N_997,N_4761);
or U6480 (N_6480,N_618,N_3480);
and U6481 (N_6481,N_2742,N_1941);
xnor U6482 (N_6482,N_53,N_2447);
xor U6483 (N_6483,N_1778,N_4404);
and U6484 (N_6484,N_4807,N_4172);
or U6485 (N_6485,N_575,N_4737);
nand U6486 (N_6486,N_89,N_4233);
xnor U6487 (N_6487,N_380,N_3843);
nor U6488 (N_6488,N_2444,N_290);
nor U6489 (N_6489,N_4700,N_535);
nand U6490 (N_6490,N_1240,N_1117);
nand U6491 (N_6491,N_3445,N_4789);
and U6492 (N_6492,N_1621,N_3628);
xor U6493 (N_6493,N_3010,N_938);
nand U6494 (N_6494,N_1683,N_3488);
and U6495 (N_6495,N_4627,N_4548);
nor U6496 (N_6496,N_240,N_1371);
or U6497 (N_6497,N_3882,N_1272);
nand U6498 (N_6498,N_1524,N_1513);
or U6499 (N_6499,N_1787,N_4563);
xor U6500 (N_6500,N_1324,N_4149);
and U6501 (N_6501,N_4515,N_402);
and U6502 (N_6502,N_68,N_1169);
xnor U6503 (N_6503,N_1390,N_1396);
or U6504 (N_6504,N_597,N_1747);
and U6505 (N_6505,N_3623,N_4091);
and U6506 (N_6506,N_3367,N_4325);
nand U6507 (N_6507,N_4036,N_2866);
or U6508 (N_6508,N_3796,N_4634);
xor U6509 (N_6509,N_2730,N_193);
nor U6510 (N_6510,N_4612,N_4280);
xnor U6511 (N_6511,N_4061,N_1270);
and U6512 (N_6512,N_3743,N_1128);
and U6513 (N_6513,N_2216,N_3044);
and U6514 (N_6514,N_4581,N_3712);
nand U6515 (N_6515,N_1068,N_827);
xor U6516 (N_6516,N_4071,N_3715);
or U6517 (N_6517,N_4216,N_3683);
nor U6518 (N_6518,N_3709,N_3514);
and U6519 (N_6519,N_4947,N_851);
nand U6520 (N_6520,N_1074,N_2914);
nand U6521 (N_6521,N_3532,N_3535);
nor U6522 (N_6522,N_1841,N_4271);
and U6523 (N_6523,N_1875,N_3559);
nor U6524 (N_6524,N_2034,N_4040);
nor U6525 (N_6525,N_961,N_1676);
xnor U6526 (N_6526,N_115,N_3617);
and U6527 (N_6527,N_4052,N_2623);
xor U6528 (N_6528,N_1780,N_971);
nand U6529 (N_6529,N_2134,N_3484);
nor U6530 (N_6530,N_1422,N_1473);
nor U6531 (N_6531,N_4167,N_1920);
nand U6532 (N_6532,N_984,N_625);
xor U6533 (N_6533,N_592,N_3945);
xor U6534 (N_6534,N_2026,N_2252);
xnor U6535 (N_6535,N_3038,N_4447);
and U6536 (N_6536,N_1267,N_887);
nand U6537 (N_6537,N_838,N_1152);
nand U6538 (N_6538,N_2732,N_3124);
or U6539 (N_6539,N_4177,N_3364);
and U6540 (N_6540,N_296,N_931);
nor U6541 (N_6541,N_4621,N_3762);
xnor U6542 (N_6542,N_4631,N_3468);
or U6543 (N_6543,N_4017,N_2934);
or U6544 (N_6544,N_4176,N_3471);
or U6545 (N_6545,N_1342,N_757);
xnor U6546 (N_6546,N_4653,N_4080);
nor U6547 (N_6547,N_2075,N_4823);
nand U6548 (N_6548,N_196,N_3343);
nor U6549 (N_6549,N_940,N_3485);
nand U6550 (N_6550,N_3422,N_1844);
xnor U6551 (N_6551,N_2762,N_2864);
or U6552 (N_6552,N_864,N_1100);
nor U6553 (N_6553,N_3321,N_879);
nor U6554 (N_6554,N_2954,N_3881);
or U6555 (N_6555,N_4713,N_693);
nand U6556 (N_6556,N_2379,N_2620);
and U6557 (N_6557,N_762,N_856);
nor U6558 (N_6558,N_3778,N_4992);
and U6559 (N_6559,N_4668,N_293);
nor U6560 (N_6560,N_2871,N_4908);
xnor U6561 (N_6561,N_241,N_1133);
nand U6562 (N_6562,N_1162,N_1961);
or U6563 (N_6563,N_374,N_945);
nand U6564 (N_6564,N_1679,N_3633);
nand U6565 (N_6565,N_1397,N_4154);
xnor U6566 (N_6566,N_133,N_3866);
nand U6567 (N_6567,N_4328,N_3918);
nor U6568 (N_6568,N_2636,N_2776);
nor U6569 (N_6569,N_1273,N_4386);
and U6570 (N_6570,N_4326,N_1527);
nor U6571 (N_6571,N_2478,N_2306);
or U6572 (N_6572,N_1063,N_4116);
or U6573 (N_6573,N_1186,N_234);
and U6574 (N_6574,N_2453,N_536);
nand U6575 (N_6575,N_2521,N_1030);
or U6576 (N_6576,N_1127,N_4306);
xor U6577 (N_6577,N_2701,N_4517);
xor U6578 (N_6578,N_1871,N_2035);
nand U6579 (N_6579,N_1209,N_2489);
nor U6580 (N_6580,N_749,N_4725);
xor U6581 (N_6581,N_2839,N_3596);
nand U6582 (N_6582,N_1405,N_3099);
nand U6583 (N_6583,N_2367,N_3030);
nand U6584 (N_6584,N_31,N_1851);
nor U6585 (N_6585,N_2459,N_4979);
and U6586 (N_6586,N_761,N_2706);
or U6587 (N_6587,N_3510,N_865);
or U6588 (N_6588,N_1035,N_3699);
nor U6589 (N_6589,N_766,N_2027);
nand U6590 (N_6590,N_1619,N_4322);
nand U6591 (N_6591,N_238,N_375);
and U6592 (N_6592,N_1316,N_2484);
or U6593 (N_6593,N_4551,N_777);
or U6594 (N_6594,N_3065,N_1786);
nor U6595 (N_6595,N_4981,N_1347);
and U6596 (N_6596,N_614,N_2766);
nor U6597 (N_6597,N_1306,N_4053);
xnor U6598 (N_6598,N_4801,N_2657);
xnor U6599 (N_6599,N_207,N_955);
or U6600 (N_6600,N_4753,N_3972);
and U6601 (N_6601,N_4878,N_3924);
xor U6602 (N_6602,N_4424,N_3058);
nor U6603 (N_6603,N_3492,N_451);
xor U6604 (N_6604,N_4369,N_836);
or U6605 (N_6605,N_4715,N_4587);
xnor U6606 (N_6606,N_1175,N_1191);
nor U6607 (N_6607,N_638,N_19);
nor U6608 (N_6608,N_2130,N_4970);
nor U6609 (N_6609,N_2865,N_4407);
and U6610 (N_6610,N_771,N_3635);
xor U6611 (N_6611,N_1757,N_2231);
nand U6612 (N_6612,N_3859,N_4986);
xor U6613 (N_6613,N_958,N_2752);
or U6614 (N_6614,N_163,N_2066);
nor U6615 (N_6615,N_1378,N_4585);
xnor U6616 (N_6616,N_4741,N_1279);
nor U6617 (N_6617,N_1258,N_1436);
and U6618 (N_6618,N_2568,N_1491);
and U6619 (N_6619,N_276,N_996);
nor U6620 (N_6620,N_1790,N_4573);
nand U6621 (N_6621,N_1943,N_1215);
xor U6622 (N_6622,N_1456,N_1865);
and U6623 (N_6623,N_1448,N_2618);
nor U6624 (N_6624,N_2516,N_2952);
xnor U6625 (N_6625,N_35,N_2765);
or U6626 (N_6626,N_3413,N_3558);
and U6627 (N_6627,N_122,N_4132);
xor U6628 (N_6628,N_4980,N_4207);
nor U6629 (N_6629,N_2834,N_2415);
or U6630 (N_6630,N_2911,N_1590);
nand U6631 (N_6631,N_2562,N_3735);
xor U6632 (N_6632,N_3640,N_151);
xnor U6633 (N_6633,N_4392,N_4544);
and U6634 (N_6634,N_3150,N_3323);
nand U6635 (N_6635,N_4844,N_3434);
and U6636 (N_6636,N_1784,N_3286);
nand U6637 (N_6637,N_3920,N_3225);
nand U6638 (N_6638,N_2912,N_3716);
or U6639 (N_6639,N_2718,N_4103);
or U6640 (N_6640,N_1148,N_4811);
nor U6641 (N_6641,N_1957,N_484);
nand U6642 (N_6642,N_2445,N_635);
or U6643 (N_6643,N_1535,N_4283);
or U6644 (N_6644,N_3217,N_4599);
or U6645 (N_6645,N_4880,N_1591);
xor U6646 (N_6646,N_2230,N_1781);
and U6647 (N_6647,N_2395,N_3914);
nand U6648 (N_6648,N_3600,N_3919);
or U6649 (N_6649,N_720,N_3938);
nor U6650 (N_6650,N_323,N_4743);
nor U6651 (N_6651,N_2506,N_1176);
nor U6652 (N_6652,N_4991,N_4983);
and U6653 (N_6653,N_94,N_4229);
nand U6654 (N_6654,N_3653,N_3112);
and U6655 (N_6655,N_152,N_2674);
or U6656 (N_6656,N_2148,N_3930);
or U6657 (N_6657,N_2386,N_3877);
xor U6658 (N_6658,N_3463,N_2945);
xnor U6659 (N_6659,N_1381,N_640);
or U6660 (N_6660,N_3751,N_220);
xnor U6661 (N_6661,N_4413,N_4601);
nor U6662 (N_6662,N_2080,N_4511);
or U6663 (N_6663,N_3758,N_3143);
nor U6664 (N_6664,N_959,N_235);
and U6665 (N_6665,N_1712,N_2695);
nor U6666 (N_6666,N_1210,N_518);
or U6667 (N_6667,N_1105,N_3450);
xor U6668 (N_6668,N_4630,N_4159);
nand U6669 (N_6669,N_4902,N_4526);
xnor U6670 (N_6670,N_4088,N_3987);
nor U6671 (N_6671,N_317,N_1399);
xnor U6672 (N_6672,N_1069,N_3686);
and U6673 (N_6673,N_1639,N_399);
and U6674 (N_6674,N_4543,N_1506);
and U6675 (N_6675,N_639,N_2475);
and U6676 (N_6676,N_310,N_1094);
or U6677 (N_6677,N_2563,N_4470);
xnor U6678 (N_6678,N_150,N_4174);
and U6679 (N_6679,N_4282,N_1716);
xor U6680 (N_6680,N_830,N_4158);
or U6681 (N_6681,N_3840,N_4659);
nor U6682 (N_6682,N_2581,N_3176);
nand U6683 (N_6683,N_4311,N_928);
and U6684 (N_6684,N_2029,N_4918);
nor U6685 (N_6685,N_3508,N_1470);
or U6686 (N_6686,N_369,N_4641);
nand U6687 (N_6687,N_412,N_1901);
nor U6688 (N_6688,N_1076,N_214);
nor U6689 (N_6689,N_4509,N_3942);
nor U6690 (N_6690,N_497,N_332);
nand U6691 (N_6691,N_1222,N_2417);
nand U6692 (N_6692,N_445,N_3993);
or U6693 (N_6693,N_4871,N_4480);
or U6694 (N_6694,N_2720,N_1255);
nor U6695 (N_6695,N_2070,N_732);
nand U6696 (N_6696,N_284,N_3245);
and U6697 (N_6697,N_1022,N_1343);
and U6698 (N_6698,N_3310,N_1070);
and U6699 (N_6699,N_1161,N_2947);
nor U6700 (N_6700,N_4112,N_3218);
xnor U6701 (N_6701,N_2611,N_3950);
nor U6702 (N_6702,N_198,N_4383);
xnor U6703 (N_6703,N_2806,N_4075);
or U6704 (N_6704,N_2746,N_1867);
xor U6705 (N_6705,N_232,N_1958);
nor U6706 (N_6706,N_4142,N_4718);
and U6707 (N_6707,N_189,N_2577);
xor U6708 (N_6708,N_4799,N_1711);
nor U6709 (N_6709,N_690,N_1723);
nand U6710 (N_6710,N_2146,N_3230);
nand U6711 (N_6711,N_2246,N_4304);
xnor U6712 (N_6712,N_603,N_2677);
and U6713 (N_6713,N_729,N_2183);
nor U6714 (N_6714,N_1547,N_2050);
and U6715 (N_6715,N_4916,N_2309);
nand U6716 (N_6716,N_3495,N_3612);
nand U6717 (N_6717,N_4060,N_3070);
and U6718 (N_6718,N_4062,N_4649);
and U6719 (N_6719,N_4044,N_1627);
and U6720 (N_6720,N_3097,N_354);
nand U6721 (N_6721,N_3838,N_3045);
or U6722 (N_6722,N_4009,N_4098);
nand U6723 (N_6723,N_2993,N_3258);
nand U6724 (N_6724,N_652,N_1468);
and U6725 (N_6725,N_1921,N_2017);
nor U6726 (N_6726,N_4829,N_3911);
nand U6727 (N_6727,N_2276,N_1896);
xor U6728 (N_6728,N_832,N_914);
nor U6729 (N_6729,N_1668,N_1888);
xnor U6730 (N_6730,N_989,N_1073);
or U6731 (N_6731,N_3269,N_2350);
nor U6732 (N_6732,N_4593,N_1965);
and U6733 (N_6733,N_4269,N_1423);
xnor U6734 (N_6734,N_1724,N_2362);
xor U6735 (N_6735,N_3223,N_3389);
nor U6736 (N_6736,N_4417,N_2055);
nor U6737 (N_6737,N_4137,N_3406);
nor U6738 (N_6738,N_526,N_1144);
and U6739 (N_6739,N_1461,N_223);
nor U6740 (N_6740,N_2909,N_2777);
nor U6741 (N_6741,N_156,N_3795);
or U6742 (N_6742,N_3332,N_2173);
xor U6743 (N_6743,N_4607,N_1376);
or U6744 (N_6744,N_3253,N_2627);
or U6745 (N_6745,N_1352,N_2037);
nand U6746 (N_6746,N_4411,N_3836);
or U6747 (N_6747,N_3460,N_448);
or U6748 (N_6748,N_2710,N_1449);
or U6749 (N_6749,N_1463,N_2494);
nor U6750 (N_6750,N_2960,N_1520);
and U6751 (N_6751,N_2435,N_828);
nand U6752 (N_6752,N_1474,N_1565);
and U6753 (N_6753,N_2558,N_4567);
xnor U6754 (N_6754,N_1401,N_1438);
nand U6755 (N_6755,N_2861,N_131);
or U6756 (N_6756,N_787,N_4189);
and U6757 (N_6757,N_1814,N_2120);
and U6758 (N_6758,N_4645,N_3157);
and U6759 (N_6759,N_877,N_2102);
nand U6760 (N_6760,N_4889,N_3352);
and U6761 (N_6761,N_1064,N_197);
or U6762 (N_6762,N_3477,N_3487);
nor U6763 (N_6763,N_3423,N_4449);
and U6764 (N_6764,N_2360,N_1861);
or U6765 (N_6765,N_4153,N_1542);
nand U6766 (N_6766,N_4093,N_1685);
xnor U6767 (N_6767,N_511,N_312);
nand U6768 (N_6768,N_124,N_3290);
nand U6769 (N_6769,N_799,N_1859);
nor U6770 (N_6770,N_2375,N_3941);
nand U6771 (N_6771,N_728,N_2862);
and U6772 (N_6772,N_4004,N_1671);
or U6773 (N_6773,N_3419,N_4925);
and U6774 (N_6774,N_2145,N_3542);
nand U6775 (N_6775,N_98,N_161);
and U6776 (N_6776,N_3325,N_2918);
nor U6777 (N_6777,N_3536,N_1414);
and U6778 (N_6778,N_872,N_1134);
xor U6779 (N_6779,N_1304,N_4165);
nand U6780 (N_6780,N_2988,N_2191);
nor U6781 (N_6781,N_2594,N_763);
nand U6782 (N_6782,N_3417,N_2049);
nor U6783 (N_6783,N_2860,N_4489);
nand U6784 (N_6784,N_3473,N_347);
and U6785 (N_6785,N_1930,N_3991);
and U6786 (N_6786,N_3465,N_3096);
nor U6787 (N_6787,N_3643,N_4640);
xnor U6788 (N_6788,N_2994,N_4030);
xnor U6789 (N_6789,N_3429,N_3722);
or U6790 (N_6790,N_598,N_2503);
or U6791 (N_6791,N_2547,N_2798);
xor U6792 (N_6792,N_3651,N_2587);
nor U6793 (N_6793,N_3652,N_4245);
nor U6794 (N_6794,N_4760,N_4293);
xnor U6795 (N_6795,N_2787,N_2077);
and U6796 (N_6796,N_174,N_611);
nand U6797 (N_6797,N_1935,N_1058);
xnor U6798 (N_6798,N_346,N_1857);
nor U6799 (N_6799,N_4454,N_2802);
nand U6800 (N_6800,N_4960,N_2606);
xor U6801 (N_6801,N_1631,N_2715);
nand U6802 (N_6802,N_4876,N_1066);
nand U6803 (N_6803,N_2178,N_1299);
nand U6804 (N_6804,N_4738,N_3279);
and U6805 (N_6805,N_2144,N_4426);
and U6806 (N_6806,N_3077,N_700);
nand U6807 (N_6807,N_280,N_1156);
or U6808 (N_6808,N_2585,N_187);
nand U6809 (N_6809,N_3056,N_2824);
and U6810 (N_6810,N_1077,N_4847);
and U6811 (N_6811,N_1326,N_4828);
and U6812 (N_6812,N_4039,N_3888);
nor U6813 (N_6813,N_886,N_722);
or U6814 (N_6814,N_3966,N_1927);
and U6815 (N_6815,N_237,N_3638);
nand U6816 (N_6816,N_4917,N_3432);
xnor U6817 (N_6817,N_487,N_774);
and U6818 (N_6818,N_3853,N_2888);
or U6819 (N_6819,N_3212,N_3520);
or U6820 (N_6820,N_4284,N_4834);
xor U6821 (N_6821,N_505,N_1071);
xnor U6822 (N_6822,N_1087,N_2940);
nor U6823 (N_6823,N_2382,N_3264);
nand U6824 (N_6824,N_3828,N_2943);
nor U6825 (N_6825,N_3576,N_4848);
xor U6826 (N_6826,N_1969,N_3240);
or U6827 (N_6827,N_2709,N_4157);
or U6828 (N_6828,N_845,N_99);
and U6829 (N_6829,N_2298,N_908);
or U6830 (N_6830,N_4101,N_3117);
and U6831 (N_6831,N_2201,N_1302);
and U6832 (N_6832,N_714,N_2704);
nor U6833 (N_6833,N_3342,N_657);
nor U6834 (N_6834,N_4879,N_2895);
nor U6835 (N_6835,N_2571,N_4998);
nor U6836 (N_6836,N_4279,N_3249);
and U6837 (N_6837,N_268,N_1114);
nor U6838 (N_6838,N_4261,N_3550);
nand U6839 (N_6839,N_540,N_1150);
nand U6840 (N_6840,N_3189,N_2357);
nand U6841 (N_6841,N_3193,N_4525);
xnor U6842 (N_6842,N_4661,N_794);
and U6843 (N_6843,N_3672,N_4422);
nor U6844 (N_6844,N_4488,N_2222);
or U6845 (N_6845,N_3365,N_1846);
nor U6846 (N_6846,N_1955,N_3411);
and U6847 (N_6847,N_2267,N_768);
and U6848 (N_6848,N_3563,N_2020);
nor U6849 (N_6849,N_3738,N_3771);
xor U6850 (N_6850,N_4019,N_3167);
or U6851 (N_6851,N_184,N_2335);
and U6852 (N_6852,N_2486,N_504);
or U6853 (N_6853,N_3821,N_2422);
and U6854 (N_6854,N_3023,N_3316);
and U6855 (N_6855,N_2067,N_3549);
nand U6856 (N_6856,N_1170,N_1700);
and U6857 (N_6857,N_4695,N_1346);
or U6858 (N_6858,N_430,N_4255);
nand U6859 (N_6859,N_3052,N_3826);
nand U6860 (N_6860,N_2389,N_4361);
xnor U6861 (N_6861,N_1849,N_1165);
and U6862 (N_6862,N_4990,N_213);
nor U6863 (N_6863,N_2409,N_206);
or U6864 (N_6864,N_2856,N_1985);
nand U6865 (N_6865,N_3870,N_2028);
and U6866 (N_6866,N_739,N_3374);
and U6867 (N_6867,N_4898,N_1054);
nand U6868 (N_6868,N_527,N_2845);
nand U6869 (N_6869,N_3137,N_4746);
xnor U6870 (N_6870,N_34,N_1109);
xor U6871 (N_6871,N_4418,N_3910);
xnor U6872 (N_6872,N_83,N_4557);
nor U6873 (N_6873,N_3154,N_2770);
nand U6874 (N_6874,N_2016,N_4937);
or U6875 (N_6875,N_1855,N_3272);
nand U6876 (N_6876,N_3062,N_571);
nand U6877 (N_6877,N_336,N_2356);
nand U6878 (N_6878,N_4481,N_2738);
nand U6879 (N_6879,N_4128,N_1854);
and U6880 (N_6880,N_2642,N_2200);
xor U6881 (N_6881,N_4058,N_2219);
xor U6882 (N_6882,N_3050,N_861);
nand U6883 (N_6883,N_1717,N_1452);
nand U6884 (N_6884,N_147,N_2196);
nor U6885 (N_6885,N_2469,N_2676);
and U6886 (N_6886,N_3360,N_3145);
and U6887 (N_6887,N_3390,N_3273);
nor U6888 (N_6888,N_3960,N_4234);
or U6889 (N_6889,N_194,N_4079);
or U6890 (N_6890,N_1603,N_3685);
nor U6891 (N_6891,N_3005,N_3017);
xnor U6892 (N_6892,N_2143,N_3416);
nor U6893 (N_6893,N_2972,N_173);
and U6894 (N_6894,N_200,N_3659);
xor U6895 (N_6895,N_1458,N_4096);
xor U6896 (N_6896,N_4180,N_4769);
xnor U6897 (N_6897,N_4999,N_816);
nor U6898 (N_6898,N_3006,N_1495);
and U6899 (N_6899,N_2553,N_2973);
or U6900 (N_6900,N_1994,N_1481);
or U6901 (N_6901,N_3035,N_969);
nor U6902 (N_6902,N_775,N_1538);
nand U6903 (N_6903,N_2397,N_672);
xor U6904 (N_6904,N_2903,N_1902);
nor U6905 (N_6905,N_2118,N_2041);
or U6906 (N_6906,N_772,N_1278);
and U6907 (N_6907,N_1275,N_1384);
nand U6908 (N_6908,N_1618,N_1567);
xor U6909 (N_6909,N_3354,N_4178);
nor U6910 (N_6910,N_3133,N_3876);
or U6911 (N_6911,N_1435,N_1395);
xnor U6912 (N_6912,N_2212,N_3561);
and U6913 (N_6913,N_2951,N_3031);
nand U6914 (N_6914,N_3823,N_1112);
or U6915 (N_6915,N_3418,N_796);
and U6916 (N_6916,N_3809,N_1293);
nand U6917 (N_6917,N_3790,N_647);
nor U6918 (N_6918,N_4440,N_1236);
and U6919 (N_6919,N_502,N_1018);
nand U6920 (N_6920,N_4421,N_4527);
or U6921 (N_6921,N_1358,N_2205);
nand U6922 (N_6922,N_2090,N_4584);
and U6923 (N_6923,N_951,N_1168);
nand U6924 (N_6924,N_898,N_4714);
nor U6925 (N_6925,N_3455,N_3292);
nor U6926 (N_6926,N_4428,N_4963);
or U6927 (N_6927,N_4647,N_4953);
nand U6928 (N_6928,N_2175,N_1271);
xnor U6929 (N_6929,N_1230,N_3889);
xor U6930 (N_6930,N_1479,N_4748);
nor U6931 (N_6931,N_4731,N_1370);
and U6932 (N_6932,N_54,N_3556);
xnor U6933 (N_6933,N_3504,N_1402);
nor U6934 (N_6934,N_1484,N_4377);
xor U6935 (N_6935,N_4113,N_4145);
nand U6936 (N_6936,N_1528,N_4100);
or U6937 (N_6937,N_3073,N_2431);
nand U6938 (N_6938,N_1045,N_837);
and U6939 (N_6939,N_1697,N_2811);
or U6940 (N_6940,N_3565,N_4226);
nor U6941 (N_6941,N_4739,N_1522);
nand U6942 (N_6942,N_435,N_3800);
nor U6943 (N_6943,N_2218,N_1005);
nand U6944 (N_6944,N_2637,N_2481);
nor U6945 (N_6945,N_4253,N_3647);
or U6946 (N_6946,N_1764,N_3539);
nor U6947 (N_6947,N_1055,N_2566);
nand U6948 (N_6948,N_3805,N_1348);
or U6949 (N_6949,N_1525,N_2984);
or U6950 (N_6950,N_4476,N_1357);
and U6951 (N_6951,N_4187,N_3165);
xor U6952 (N_6952,N_4262,N_1287);
or U6953 (N_6953,N_4455,N_2176);
nand U6954 (N_6954,N_1796,N_2136);
or U6955 (N_6955,N_1200,N_2318);
nand U6956 (N_6956,N_65,N_4529);
or U6957 (N_6957,N_520,N_885);
or U6958 (N_6958,N_4676,N_292);
or U6959 (N_6959,N_2992,N_1016);
xnor U6960 (N_6960,N_1939,N_2282);
and U6961 (N_6961,N_1652,N_3381);
xnor U6962 (N_6962,N_1828,N_2561);
and U6963 (N_6963,N_406,N_2006);
or U6964 (N_6964,N_793,N_1531);
or U6965 (N_6965,N_4482,N_459);
or U6966 (N_6966,N_2314,N_4370);
nand U6967 (N_6967,N_1398,N_1945);
or U6968 (N_6968,N_287,N_1455);
nor U6969 (N_6969,N_3724,N_2630);
nand U6970 (N_6970,N_4238,N_4712);
xnor U6971 (N_6971,N_4606,N_1303);
xor U6972 (N_6972,N_691,N_4260);
xor U6973 (N_6973,N_4669,N_2857);
xnor U6974 (N_6974,N_4533,N_4846);
xnor U6975 (N_6975,N_2572,N_1166);
or U6976 (N_6976,N_1868,N_1748);
xor U6977 (N_6977,N_2179,N_3172);
xor U6978 (N_6978,N_2177,N_468);
nand U6979 (N_6979,N_3254,N_972);
xor U6980 (N_6980,N_3305,N_3004);
nand U6981 (N_6981,N_4704,N_1364);
or U6982 (N_6982,N_3767,N_3190);
and U6983 (N_6983,N_818,N_272);
xnor U6984 (N_6984,N_4875,N_4657);
nand U6985 (N_6985,N_2575,N_3951);
nand U6986 (N_6986,N_3946,N_4343);
and U6987 (N_6987,N_4342,N_1197);
nand U6988 (N_6988,N_716,N_3682);
nand U6989 (N_6989,N_3114,N_1301);
nor U6990 (N_6990,N_1504,N_456);
and U6991 (N_6991,N_1566,N_180);
xnor U6992 (N_6992,N_1042,N_1228);
and U6993 (N_6993,N_804,N_2653);
or U6994 (N_6994,N_454,N_4276);
and U6995 (N_6995,N_1498,N_769);
or U6996 (N_6996,N_10,N_2753);
nor U6997 (N_6997,N_673,N_144);
nand U6998 (N_6998,N_3373,N_1061);
xor U6999 (N_6999,N_4597,N_2979);
xor U7000 (N_7000,N_2957,N_305);
nand U7001 (N_7001,N_2771,N_2251);
xor U7002 (N_7002,N_2995,N_1752);
or U7003 (N_7003,N_4247,N_4552);
and U7004 (N_7004,N_3538,N_1934);
xor U7005 (N_7005,N_2591,N_441);
or U7006 (N_7006,N_1420,N_1500);
xor U7007 (N_7007,N_1722,N_3398);
xnor U7008 (N_7008,N_3252,N_2661);
nand U7009 (N_7009,N_148,N_1699);
and U7010 (N_7010,N_4977,N_4968);
xor U7011 (N_7011,N_231,N_927);
xor U7012 (N_7012,N_471,N_111);
nor U7013 (N_7013,N_1111,N_4150);
nand U7014 (N_7014,N_4479,N_4254);
or U7015 (N_7015,N_1507,N_1437);
and U7016 (N_7016,N_2830,N_2393);
nor U7017 (N_7017,N_1193,N_1180);
and U7018 (N_7018,N_4776,N_4553);
nand U7019 (N_7019,N_1912,N_4250);
xor U7020 (N_7020,N_4856,N_2188);
and U7021 (N_7021,N_107,N_924);
or U7022 (N_7022,N_1983,N_4542);
nand U7023 (N_7023,N_4972,N_1907);
or U7024 (N_7024,N_4016,N_1911);
nand U7025 (N_7025,N_301,N_3701);
nand U7026 (N_7026,N_4301,N_3846);
and U7027 (N_7027,N_2227,N_486);
or U7028 (N_7028,N_3907,N_1413);
nand U7029 (N_7029,N_2440,N_1321);
nand U7030 (N_7030,N_1430,N_3174);
nor U7031 (N_7031,N_4541,N_4572);
and U7032 (N_7032,N_4588,N_835);
nor U7033 (N_7033,N_1355,N_2407);
or U7034 (N_7034,N_63,N_3384);
nor U7035 (N_7035,N_783,N_3654);
and U7036 (N_7036,N_3980,N_3825);
nand U7037 (N_7037,N_3247,N_2003);
nor U7038 (N_7038,N_3619,N_2158);
nand U7039 (N_7039,N_3958,N_2579);
xor U7040 (N_7040,N_3187,N_165);
xnor U7041 (N_7041,N_483,N_4708);
and U7042 (N_7042,N_3848,N_2768);
xor U7043 (N_7043,N_1027,N_3057);
nand U7044 (N_7044,N_4155,N_4747);
or U7045 (N_7045,N_2449,N_4212);
or U7046 (N_7046,N_2987,N_1726);
xor U7047 (N_7047,N_3937,N_3864);
and U7048 (N_7048,N_352,N_3624);
and U7049 (N_7049,N_3551,N_3630);
and U7050 (N_7050,N_2223,N_4055);
nor U7051 (N_7051,N_4952,N_4414);
or U7052 (N_7052,N_4775,N_0);
and U7053 (N_7053,N_17,N_1688);
nor U7054 (N_7054,N_2989,N_4186);
or U7055 (N_7055,N_1179,N_2310);
or U7056 (N_7056,N_1534,N_3356);
nand U7057 (N_7057,N_1838,N_377);
xnor U7058 (N_7058,N_3957,N_892);
nor U7059 (N_7059,N_4023,N_3358);
xnor U7060 (N_7060,N_3974,N_2274);
nor U7061 (N_7061,N_723,N_2897);
xnor U7062 (N_7062,N_2108,N_4263);
or U7063 (N_7063,N_1758,N_4048);
nand U7064 (N_7064,N_3177,N_1559);
and U7065 (N_7065,N_1339,N_4628);
nand U7066 (N_7066,N_2907,N_1060);
nand U7067 (N_7067,N_3257,N_3747);
xor U7068 (N_7068,N_3339,N_1201);
nand U7069 (N_7069,N_2408,N_3903);
xnor U7070 (N_7070,N_4859,N_3284);
xor U7071 (N_7071,N_2160,N_1804);
or U7072 (N_7072,N_1025,N_1471);
or U7073 (N_7073,N_3862,N_365);
xnor U7074 (N_7074,N_4514,N_2485);
nor U7075 (N_7075,N_4051,N_2162);
nand U7076 (N_7076,N_2778,N_721);
nor U7077 (N_7077,N_2894,N_3196);
xor U7078 (N_7078,N_3393,N_3083);
nor U7079 (N_7079,N_4046,N_1419);
xnor U7080 (N_7080,N_1256,N_3605);
and U7081 (N_7081,N_2728,N_4068);
nand U7082 (N_7082,N_3282,N_2272);
nand U7083 (N_7083,N_2810,N_3797);
xor U7084 (N_7084,N_2882,N_850);
xor U7085 (N_7085,N_840,N_4638);
and U7086 (N_7086,N_2504,N_3534);
and U7087 (N_7087,N_3883,N_2165);
nand U7088 (N_7088,N_4483,N_2527);
xor U7089 (N_7089,N_1834,N_2156);
and U7090 (N_7090,N_1698,N_135);
nand U7091 (N_7091,N_1383,N_3015);
and U7092 (N_7092,N_4001,N_2076);
nand U7093 (N_7093,N_3241,N_3721);
or U7094 (N_7094,N_3246,N_2881);
and U7095 (N_7095,N_4728,N_4632);
nor U7096 (N_7096,N_1560,N_2079);
nand U7097 (N_7097,N_494,N_2376);
and U7098 (N_7098,N_4175,N_1703);
nor U7099 (N_7099,N_1140,N_4348);
and U7100 (N_7100,N_4443,N_1511);
nand U7101 (N_7101,N_4923,N_668);
nor U7102 (N_7102,N_3028,N_621);
xor U7103 (N_7103,N_541,N_641);
or U7104 (N_7104,N_2613,N_3634);
and U7105 (N_7105,N_3967,N_3063);
xor U7106 (N_7106,N_3601,N_2190);
or U7107 (N_7107,N_4380,N_3526);
or U7108 (N_7108,N_3511,N_4307);
xnor U7109 (N_7109,N_712,N_2380);
nand U7110 (N_7110,N_676,N_1125);
and U7111 (N_7111,N_3405,N_171);
and U7112 (N_7112,N_3916,N_4070);
or U7113 (N_7113,N_4798,N_3274);
nand U7114 (N_7114,N_2790,N_2082);
xor U7115 (N_7115,N_2129,N_215);
or U7116 (N_7116,N_4513,N_1433);
xnor U7117 (N_7117,N_488,N_4203);
or U7118 (N_7118,N_422,N_141);
xnor U7119 (N_7119,N_4258,N_4013);
and U7120 (N_7120,N_4133,N_3206);
or U7121 (N_7121,N_1243,N_2772);
nand U7122 (N_7122,N_4759,N_4590);
and U7123 (N_7123,N_613,N_4357);
nor U7124 (N_7124,N_1620,N_3128);
xor U7125 (N_7125,N_3259,N_926);
xor U7126 (N_7126,N_3159,N_1884);
and U7127 (N_7127,N_4102,N_4434);
xor U7128 (N_7128,N_734,N_1809);
or U7129 (N_7129,N_4491,N_3665);
and U7130 (N_7130,N_2831,N_1806);
nand U7131 (N_7131,N_4134,N_948);
xnor U7132 (N_7132,N_4831,N_120);
nor U7133 (N_7133,N_573,N_3865);
nand U7134 (N_7134,N_2959,N_1552);
xor U7135 (N_7135,N_733,N_3209);
xor U7136 (N_7136,N_3879,N_3234);
or U7137 (N_7137,N_4371,N_3964);
nand U7138 (N_7138,N_2119,N_689);
nand U7139 (N_7139,N_4750,N_2009);
nand U7140 (N_7140,N_384,N_4559);
xor U7141 (N_7141,N_3971,N_679);
nor U7142 (N_7142,N_561,N_653);
and U7143 (N_7143,N_1742,N_1928);
nor U7144 (N_7144,N_450,N_1785);
and U7145 (N_7145,N_1978,N_4764);
nand U7146 (N_7146,N_4464,N_553);
or U7147 (N_7147,N_1332,N_1885);
xnor U7148 (N_7148,N_3098,N_2507);
xnor U7149 (N_7149,N_1815,N_2522);
nand U7150 (N_7150,N_3897,N_902);
xor U7151 (N_7151,N_4997,N_1151);
xnor U7152 (N_7152,N_1873,N_660);
xnor U7153 (N_7153,N_2809,N_4815);
nand U7154 (N_7154,N_549,N_4796);
or U7155 (N_7155,N_3698,N_1189);
and U7156 (N_7156,N_1843,N_1611);
xor U7157 (N_7157,N_4460,N_1774);
and U7158 (N_7158,N_740,N_4446);
nor U7159 (N_7159,N_1298,N_138);
and U7160 (N_7160,N_3676,N_4498);
and U7161 (N_7161,N_4399,N_3337);
xnor U7162 (N_7162,N_3642,N_88);
nand U7163 (N_7163,N_2281,N_4225);
nand U7164 (N_7164,N_191,N_3483);
and U7165 (N_7165,N_2733,N_1973);
nand U7166 (N_7166,N_4758,N_3872);
nor U7167 (N_7167,N_2432,N_4218);
nand U7168 (N_7168,N_2396,N_1294);
nor U7169 (N_7169,N_3718,N_2463);
xnor U7170 (N_7170,N_944,N_3459);
nand U7171 (N_7171,N_2295,N_2534);
and U7172 (N_7172,N_4287,N_4681);
and U7173 (N_7173,N_4141,N_1580);
nand U7174 (N_7174,N_4015,N_2242);
xnor U7175 (N_7175,N_2671,N_2072);
xnor U7176 (N_7176,N_3664,N_2672);
and U7177 (N_7177,N_3327,N_1772);
or U7178 (N_7178,N_3689,N_727);
nor U7179 (N_7179,N_3753,N_3671);
or U7180 (N_7180,N_637,N_4549);
or U7181 (N_7181,N_2474,N_863);
xor U7182 (N_7182,N_1119,N_3500);
nor U7183 (N_7183,N_2168,N_1135);
nand U7184 (N_7184,N_3965,N_3737);
xor U7185 (N_7185,N_4537,N_224);
or U7186 (N_7186,N_4501,N_4459);
nand U7187 (N_7187,N_1213,N_3981);
xnor U7188 (N_7188,N_253,N_2889);
nand U7189 (N_7189,N_3572,N_4214);
and U7190 (N_7190,N_1922,N_2905);
nand U7191 (N_7191,N_3407,N_2876);
xor U7192 (N_7192,N_848,N_4662);
xor U7193 (N_7193,N_1750,N_481);
and U7194 (N_7194,N_4862,N_458);
and U7195 (N_7195,N_2707,N_3806);
or U7196 (N_7196,N_633,N_4872);
xnor U7197 (N_7197,N_1317,N_297);
and U7198 (N_7198,N_4217,N_429);
nand U7199 (N_7199,N_1825,N_4412);
or U7200 (N_7200,N_3837,N_3127);
xnor U7201 (N_7201,N_4381,N_2476);
and U7202 (N_7202,N_385,N_3203);
and U7203 (N_7203,N_2680,N_4840);
and U7204 (N_7204,N_3863,N_1623);
xor U7205 (N_7205,N_4989,N_1219);
nand U7206 (N_7206,N_4206,N_2662);
nor U7207 (N_7207,N_2826,N_1229);
nand U7208 (N_7208,N_2819,N_1753);
and U7209 (N_7209,N_4904,N_3263);
xor U7210 (N_7210,N_3636,N_4765);
or U7211 (N_7211,N_713,N_2990);
or U7212 (N_7212,N_2665,N_1281);
and U7213 (N_7213,N_2245,N_2015);
and U7214 (N_7214,N_4824,N_533);
or U7215 (N_7215,N_3708,N_4558);
and U7216 (N_7216,N_4729,N_3772);
or U7217 (N_7217,N_3961,N_2670);
nor U7218 (N_7218,N_3027,N_4320);
nand U7219 (N_7219,N_311,N_4246);
nor U7220 (N_7220,N_907,N_4117);
nand U7221 (N_7221,N_4115,N_2448);
xor U7222 (N_7222,N_1080,N_627);
or U7223 (N_7223,N_1492,N_2345);
or U7224 (N_7224,N_3084,N_334);
and U7225 (N_7225,N_3311,N_4691);
or U7226 (N_7226,N_2404,N_3021);
xnor U7227 (N_7227,N_1296,N_343);
xnor U7228 (N_7228,N_190,N_964);
nor U7229 (N_7229,N_546,N_4576);
nand U7230 (N_7230,N_4188,N_1536);
or U7231 (N_7231,N_867,N_586);
and U7232 (N_7232,N_3519,N_1667);
and U7233 (N_7233,N_3760,N_86);
nand U7234 (N_7234,N_2692,N_4248);
nor U7235 (N_7235,N_1404,N_2827);
nor U7236 (N_7236,N_991,N_4837);
and U7237 (N_7237,N_2340,N_1754);
nor U7238 (N_7238,N_4191,N_692);
and U7239 (N_7239,N_3080,N_2458);
nand U7240 (N_7240,N_219,N_1155);
and U7241 (N_7241,N_780,N_4264);
nand U7242 (N_7242,N_3763,N_3211);
nor U7243 (N_7243,N_3637,N_1556);
nor U7244 (N_7244,N_3518,N_2867);
xor U7245 (N_7245,N_3160,N_4163);
or U7246 (N_7246,N_4996,N_4458);
or U7247 (N_7247,N_1646,N_2849);
or U7248 (N_7248,N_807,N_4962);
xnor U7249 (N_7249,N_3829,N_1572);
nand U7250 (N_7250,N_4354,N_4564);
nand U7251 (N_7251,N_1290,N_2936);
nand U7252 (N_7252,N_4337,N_2607);
or U7253 (N_7253,N_874,N_3437);
xor U7254 (N_7254,N_4745,N_4202);
nand U7255 (N_7255,N_4974,N_1192);
nand U7256 (N_7256,N_3544,N_3386);
xor U7257 (N_7257,N_3766,N_642);
nand U7258 (N_7258,N_4677,N_1083);
and U7259 (N_7259,N_2206,N_1274);
xnor U7260 (N_7260,N_303,N_3064);
and U7261 (N_7261,N_1991,N_3794);
or U7262 (N_7262,N_2966,N_3727);
xor U7263 (N_7263,N_2512,N_3527);
and U7264 (N_7264,N_2700,N_1123);
nor U7265 (N_7265,N_389,N_1361);
and U7266 (N_7266,N_1386,N_1028);
and U7267 (N_7267,N_2756,N_4064);
or U7268 (N_7268,N_4841,N_4420);
nor U7269 (N_7269,N_1946,N_2203);
nor U7270 (N_7270,N_378,N_2836);
xor U7271 (N_7271,N_671,N_1808);
xor U7272 (N_7272,N_1322,N_2166);
nor U7273 (N_7273,N_1345,N_209);
nor U7274 (N_7274,N_4784,N_2800);
nor U7275 (N_7275,N_2312,N_4010);
nor U7276 (N_7276,N_1038,N_4462);
and U7277 (N_7277,N_591,N_4885);
xor U7278 (N_7278,N_139,N_3695);
nor U7279 (N_7279,N_1738,N_4788);
and U7280 (N_7280,N_294,N_92);
xor U7281 (N_7281,N_2385,N_3803);
or U7282 (N_7282,N_2378,N_1315);
nand U7283 (N_7283,N_1049,N_3318);
nand U7284 (N_7284,N_1544,N_348);
nand U7285 (N_7285,N_4795,N_341);
nor U7286 (N_7286,N_4110,N_3214);
xnor U7287 (N_7287,N_3884,N_397);
nand U7288 (N_7288,N_1577,N_998);
nor U7289 (N_7289,N_1740,N_3755);
nand U7290 (N_7290,N_4197,N_3595);
or U7291 (N_7291,N_4766,N_1334);
nor U7292 (N_7292,N_2731,N_576);
or U7293 (N_7293,N_4710,N_2569);
nor U7294 (N_7294,N_3669,N_4072);
nor U7295 (N_7295,N_4350,N_4685);
nor U7296 (N_7296,N_870,N_2263);
or U7297 (N_7297,N_2890,N_664);
nor U7298 (N_7298,N_3749,N_2523);
xnor U7299 (N_7299,N_4787,N_1783);
xnor U7300 (N_7300,N_4318,N_2438);
or U7301 (N_7301,N_3297,N_4439);
and U7302 (N_7302,N_4024,N_3046);
xnor U7303 (N_7303,N_1194,N_4423);
nor U7304 (N_7304,N_3929,N_1816);
and U7305 (N_7305,N_2228,N_4352);
and U7306 (N_7306,N_2673,N_24);
and U7307 (N_7307,N_1862,N_1121);
nor U7308 (N_7308,N_4818,N_57);
and U7309 (N_7309,N_1476,N_105);
nor U7310 (N_7310,N_23,N_1597);
and U7311 (N_7311,N_4578,N_559);
xor U7312 (N_7312,N_379,N_589);
nor U7313 (N_7313,N_3909,N_1026);
and U7314 (N_7314,N_3963,N_500);
or U7315 (N_7315,N_387,N_4518);
xor U7316 (N_7316,N_4123,N_2131);
nand U7317 (N_7317,N_3793,N_1122);
and U7318 (N_7318,N_1938,N_3662);
nor U7319 (N_7319,N_3579,N_2741);
or U7320 (N_7320,N_132,N_1756);
xnor U7321 (N_7321,N_1034,N_1417);
nor U7322 (N_7322,N_1988,N_4457);
or U7323 (N_7323,N_3570,N_2169);
xor U7324 (N_7324,N_895,N_345);
and U7325 (N_7325,N_1777,N_4169);
xor U7326 (N_7326,N_2495,N_514);
nand U7327 (N_7327,N_3780,N_986);
or U7328 (N_7328,N_4614,N_4105);
xnor U7329 (N_7329,N_2555,N_4949);
and U7330 (N_7330,N_1009,N_1002);
nor U7331 (N_7331,N_3512,N_112);
xor U7332 (N_7332,N_2900,N_2319);
and U7333 (N_7333,N_2226,N_2614);
or U7334 (N_7334,N_4562,N_1628);
or U7335 (N_7335,N_4496,N_2304);
xnor U7336 (N_7336,N_4054,N_4555);
and U7337 (N_7337,N_3954,N_1721);
or U7338 (N_7338,N_956,N_890);
nand U7339 (N_7339,N_2498,N_3129);
nor U7340 (N_7340,N_1501,N_521);
or U7341 (N_7341,N_1327,N_4768);
nand U7342 (N_7342,N_2008,N_950);
nor U7343 (N_7343,N_4702,N_2593);
and U7344 (N_7344,N_3804,N_1464);
nand U7345 (N_7345,N_2308,N_4401);
nor U7346 (N_7346,N_3585,N_2978);
or U7347 (N_7347,N_3357,N_2551);
xnor U7348 (N_7348,N_564,N_3300);
or U7349 (N_7349,N_3486,N_2243);
and U7350 (N_7350,N_443,N_4125);
or U7351 (N_7351,N_1065,N_1050);
xor U7352 (N_7352,N_3149,N_1636);
nand U7353 (N_7353,N_544,N_2418);
or U7354 (N_7354,N_644,N_114);
xor U7355 (N_7355,N_4693,N_413);
xor U7356 (N_7356,N_3541,N_710);
nand U7357 (N_7357,N_3344,N_4099);
nor U7358 (N_7358,N_3303,N_2958);
xor U7359 (N_7359,N_464,N_4566);
nand U7360 (N_7360,N_3622,N_3392);
nand U7361 (N_7361,N_704,N_1691);
nor U7362 (N_7362,N_2462,N_2948);
nor U7363 (N_7363,N_4395,N_798);
nand U7364 (N_7364,N_4575,N_4532);
and U7365 (N_7365,N_3072,N_1336);
nor U7366 (N_7366,N_2891,N_395);
xnor U7367 (N_7367,N_3383,N_4531);
nand U7368 (N_7368,N_3496,N_199);
nand U7369 (N_7369,N_1743,N_4570);
or U7370 (N_7370,N_3208,N_1249);
and U7371 (N_7371,N_1515,N_4444);
nor U7372 (N_7372,N_1488,N_730);
xnor U7373 (N_7373,N_3168,N_3547);
nor U7374 (N_7374,N_340,N_4500);
and U7375 (N_7375,N_3239,N_304);
nor U7376 (N_7376,N_4851,N_4946);
xor U7377 (N_7377,N_3324,N_3446);
xor U7378 (N_7378,N_4373,N_1719);
or U7379 (N_7379,N_4025,N_609);
nor U7380 (N_7380,N_737,N_3210);
nor U7381 (N_7381,N_3278,N_4648);
or U7382 (N_7382,N_3293,N_13);
xnor U7383 (N_7383,N_4508,N_3142);
nand U7384 (N_7384,N_4931,N_414);
nand U7385 (N_7385,N_2851,N_1079);
nor U7386 (N_7386,N_3014,N_4940);
nor U7387 (N_7387,N_411,N_4487);
or U7388 (N_7388,N_3594,N_2032);
or U7389 (N_7389,N_2805,N_4547);
and U7390 (N_7390,N_243,N_254);
nor U7391 (N_7391,N_1040,N_3466);
nand U7392 (N_7392,N_1768,N_188);
and U7393 (N_7393,N_4670,N_770);
nand U7394 (N_7394,N_1569,N_2232);
nor U7395 (N_7395,N_2349,N_3817);
or U7396 (N_7396,N_157,N_1950);
or U7397 (N_7397,N_3101,N_1966);
and U7398 (N_7398,N_620,N_2235);
nand U7399 (N_7399,N_4942,N_765);
nand U7400 (N_7400,N_2289,N_1091);
nor U7401 (N_7401,N_4793,N_2583);
or U7402 (N_7402,N_3816,N_974);
nor U7403 (N_7403,N_40,N_4334);
nand U7404 (N_7404,N_1931,N_4397);
nand U7405 (N_7405,N_2107,N_3387);
xnor U7406 (N_7406,N_2818,N_2668);
nand U7407 (N_7407,N_509,N_409);
nand U7408 (N_7408,N_2501,N_643);
and U7409 (N_7409,N_1529,N_270);
nor U7410 (N_7410,N_3289,N_2901);
or U7411 (N_7411,N_2854,N_1678);
xnor U7412 (N_7412,N_2574,N_2324);
or U7413 (N_7413,N_3869,N_8);
xnor U7414 (N_7414,N_3085,N_1647);
nand U7415 (N_7415,N_602,N_3048);
or U7416 (N_7416,N_300,N_275);
or U7417 (N_7417,N_823,N_4651);
or U7418 (N_7418,N_3363,N_3509);
and U7419 (N_7419,N_1307,N_1638);
and U7420 (N_7420,N_4140,N_3852);
nand U7421 (N_7421,N_1013,N_81);
nand U7422 (N_7422,N_1216,N_3820);
and U7423 (N_7423,N_442,N_1596);
nand U7424 (N_7424,N_1883,N_1138);
and U7425 (N_7425,N_3873,N_2726);
or U7426 (N_7426,N_935,N_3726);
xnor U7427 (N_7427,N_654,N_2689);
nand U7428 (N_7428,N_4610,N_687);
nand U7429 (N_7429,N_4545,N_1964);
or U7430 (N_7430,N_3855,N_1765);
nand U7431 (N_7431,N_2878,N_3528);
nand U7432 (N_7432,N_4958,N_1014);
xor U7433 (N_7433,N_3765,N_3238);
xor U7434 (N_7434,N_2610,N_912);
xor U7435 (N_7435,N_170,N_2100);
and U7436 (N_7436,N_4332,N_4911);
nor U7437 (N_7437,N_2663,N_4644);
nor U7438 (N_7438,N_281,N_3351);
or U7439 (N_7439,N_2001,N_3973);
or U7440 (N_7440,N_1516,N_3171);
nand U7441 (N_7441,N_2172,N_1351);
nand U7442 (N_7442,N_3000,N_4609);
nand U7443 (N_7443,N_4734,N_3994);
xnor U7444 (N_7444,N_3917,N_2468);
nor U7445 (N_7445,N_565,N_299);
xor U7446 (N_7446,N_455,N_3700);
nand U7447 (N_7447,N_2414,N_3890);
and U7448 (N_7448,N_1517,N_2043);
xor U7449 (N_7449,N_50,N_1232);
xor U7450 (N_7450,N_3725,N_1622);
and U7451 (N_7451,N_610,N_4329);
and U7452 (N_7452,N_2056,N_4893);
xor U7453 (N_7453,N_1164,N_1856);
nor U7454 (N_7454,N_2525,N_3602);
nor U7455 (N_7455,N_1508,N_202);
xnor U7456 (N_7456,N_4813,N_2869);
nor U7457 (N_7457,N_3391,N_831);
nand U7458 (N_7458,N_517,N_634);
or U7459 (N_7459,N_4281,N_3346);
nand U7460 (N_7460,N_754,N_4442);
and U7461 (N_7461,N_18,N_4615);
and U7462 (N_7462,N_3497,N_599);
xnor U7463 (N_7463,N_2682,N_2241);
xor U7464 (N_7464,N_3256,N_846);
nand U7465 (N_7465,N_2605,N_4780);
nor U7466 (N_7466,N_1800,N_2192);
nand U7467 (N_7467,N_3687,N_3905);
xnor U7468 (N_7468,N_4993,N_2648);
nor U7469 (N_7469,N_1673,N_3711);
xor U7470 (N_7470,N_2517,N_1791);
nand U7471 (N_7471,N_433,N_3197);
nand U7472 (N_7472,N_2467,N_4598);
or U7473 (N_7473,N_1923,N_440);
xnor U7474 (N_7474,N_4723,N_4235);
or U7475 (N_7475,N_2602,N_2383);
or U7476 (N_7476,N_4773,N_2544);
nand U7477 (N_7477,N_1424,N_979);
or U7478 (N_7478,N_2828,N_222);
nor U7479 (N_7479,N_4438,N_3125);
and U7480 (N_7480,N_4005,N_2926);
nor U7481 (N_7481,N_1655,N_3515);
nor U7482 (N_7482,N_813,N_3956);
nand U7483 (N_7483,N_3265,N_2374);
nor U7484 (N_7484,N_3808,N_4104);
xnor U7485 (N_7485,N_930,N_4821);
and U7486 (N_7486,N_1669,N_1604);
nor U7487 (N_7487,N_3607,N_162);
nand U7488 (N_7488,N_2471,N_980);
nor U7489 (N_7489,N_1736,N_103);
nand U7490 (N_7490,N_4351,N_113);
nor U7491 (N_7491,N_4162,N_1605);
or U7492 (N_7492,N_3451,N_2105);
nand U7493 (N_7493,N_2461,N_1325);
nand U7494 (N_7494,N_1251,N_3768);
nor U7495 (N_7495,N_3078,N_2714);
xor U7496 (N_7496,N_812,N_58);
nand U7497 (N_7497,N_1124,N_3106);
xor U7498 (N_7498,N_513,N_3694);
nor U7499 (N_7499,N_1998,N_2997);
and U7500 (N_7500,N_1944,N_4663);
nor U7501 (N_7501,N_806,N_4752);
nor U7502 (N_7502,N_3879,N_3788);
nor U7503 (N_7503,N_4653,N_2386);
or U7504 (N_7504,N_3257,N_4981);
or U7505 (N_7505,N_1912,N_4690);
xnor U7506 (N_7506,N_1280,N_3614);
nand U7507 (N_7507,N_3260,N_3282);
nor U7508 (N_7508,N_4793,N_2866);
xor U7509 (N_7509,N_4618,N_55);
nor U7510 (N_7510,N_3989,N_1681);
nor U7511 (N_7511,N_3219,N_653);
and U7512 (N_7512,N_3200,N_117);
nand U7513 (N_7513,N_2418,N_4897);
nor U7514 (N_7514,N_1483,N_4821);
xnor U7515 (N_7515,N_2553,N_978);
or U7516 (N_7516,N_1522,N_3791);
and U7517 (N_7517,N_2508,N_3394);
and U7518 (N_7518,N_4754,N_1877);
nand U7519 (N_7519,N_1366,N_2230);
nor U7520 (N_7520,N_3993,N_2485);
or U7521 (N_7521,N_2932,N_2445);
or U7522 (N_7522,N_833,N_3839);
xnor U7523 (N_7523,N_2610,N_4532);
nor U7524 (N_7524,N_12,N_1062);
xnor U7525 (N_7525,N_1079,N_1890);
and U7526 (N_7526,N_1441,N_3773);
or U7527 (N_7527,N_1158,N_3295);
nand U7528 (N_7528,N_1287,N_3950);
xnor U7529 (N_7529,N_114,N_3384);
and U7530 (N_7530,N_3086,N_3994);
or U7531 (N_7531,N_204,N_4856);
and U7532 (N_7532,N_1401,N_4307);
or U7533 (N_7533,N_3125,N_592);
xor U7534 (N_7534,N_1254,N_2689);
or U7535 (N_7535,N_3062,N_607);
xnor U7536 (N_7536,N_941,N_3073);
or U7537 (N_7537,N_779,N_946);
nand U7538 (N_7538,N_1189,N_727);
nor U7539 (N_7539,N_4828,N_4367);
nand U7540 (N_7540,N_4762,N_3869);
and U7541 (N_7541,N_2211,N_4295);
and U7542 (N_7542,N_1261,N_2584);
and U7543 (N_7543,N_1353,N_786);
xnor U7544 (N_7544,N_4034,N_1641);
or U7545 (N_7545,N_2358,N_1839);
nand U7546 (N_7546,N_158,N_2490);
and U7547 (N_7547,N_1313,N_1519);
nor U7548 (N_7548,N_4527,N_1117);
nand U7549 (N_7549,N_2883,N_2800);
or U7550 (N_7550,N_3330,N_3478);
nand U7551 (N_7551,N_809,N_1754);
nor U7552 (N_7552,N_2691,N_3825);
or U7553 (N_7553,N_2545,N_1600);
xnor U7554 (N_7554,N_4262,N_310);
xnor U7555 (N_7555,N_674,N_2842);
or U7556 (N_7556,N_2628,N_3287);
nand U7557 (N_7557,N_933,N_4263);
nor U7558 (N_7558,N_4930,N_4786);
and U7559 (N_7559,N_3131,N_3567);
xnor U7560 (N_7560,N_3483,N_3245);
and U7561 (N_7561,N_1624,N_1086);
and U7562 (N_7562,N_3128,N_2337);
nand U7563 (N_7563,N_3116,N_3484);
nor U7564 (N_7564,N_2203,N_2350);
nand U7565 (N_7565,N_1092,N_777);
nand U7566 (N_7566,N_2893,N_1311);
nor U7567 (N_7567,N_673,N_1122);
or U7568 (N_7568,N_3023,N_883);
xor U7569 (N_7569,N_1471,N_1644);
nor U7570 (N_7570,N_1770,N_594);
and U7571 (N_7571,N_3738,N_4144);
or U7572 (N_7572,N_1022,N_4209);
nor U7573 (N_7573,N_392,N_2760);
or U7574 (N_7574,N_4786,N_4421);
or U7575 (N_7575,N_3844,N_1714);
or U7576 (N_7576,N_886,N_4362);
nand U7577 (N_7577,N_2928,N_480);
nor U7578 (N_7578,N_3851,N_70);
nand U7579 (N_7579,N_127,N_2241);
xnor U7580 (N_7580,N_234,N_3635);
or U7581 (N_7581,N_2059,N_2822);
nand U7582 (N_7582,N_2328,N_2329);
or U7583 (N_7583,N_1848,N_1666);
or U7584 (N_7584,N_1024,N_2694);
xor U7585 (N_7585,N_924,N_286);
or U7586 (N_7586,N_487,N_4540);
xnor U7587 (N_7587,N_548,N_3001);
nand U7588 (N_7588,N_341,N_3685);
xnor U7589 (N_7589,N_4738,N_4097);
and U7590 (N_7590,N_2099,N_3582);
xor U7591 (N_7591,N_243,N_3605);
nand U7592 (N_7592,N_3832,N_3403);
or U7593 (N_7593,N_735,N_1730);
xnor U7594 (N_7594,N_4884,N_3515);
xnor U7595 (N_7595,N_89,N_3729);
xnor U7596 (N_7596,N_3606,N_2402);
nand U7597 (N_7597,N_1405,N_443);
nand U7598 (N_7598,N_2165,N_2);
xnor U7599 (N_7599,N_1651,N_4845);
or U7600 (N_7600,N_2247,N_4682);
xnor U7601 (N_7601,N_2053,N_1982);
nor U7602 (N_7602,N_2449,N_1205);
xor U7603 (N_7603,N_4334,N_1608);
nor U7604 (N_7604,N_2886,N_2668);
nor U7605 (N_7605,N_4618,N_151);
nor U7606 (N_7606,N_3340,N_4190);
nand U7607 (N_7607,N_896,N_440);
nor U7608 (N_7608,N_4856,N_2751);
or U7609 (N_7609,N_4957,N_2410);
and U7610 (N_7610,N_322,N_1438);
or U7611 (N_7611,N_3135,N_992);
and U7612 (N_7612,N_4309,N_1515);
nor U7613 (N_7613,N_3566,N_1558);
xor U7614 (N_7614,N_4969,N_1120);
nand U7615 (N_7615,N_2120,N_3978);
or U7616 (N_7616,N_680,N_80);
xor U7617 (N_7617,N_1622,N_2637);
nand U7618 (N_7618,N_77,N_310);
nor U7619 (N_7619,N_76,N_3644);
and U7620 (N_7620,N_4707,N_3981);
and U7621 (N_7621,N_1174,N_4692);
nand U7622 (N_7622,N_1519,N_4991);
or U7623 (N_7623,N_1278,N_1106);
and U7624 (N_7624,N_669,N_3358);
and U7625 (N_7625,N_2336,N_3392);
or U7626 (N_7626,N_252,N_3304);
nand U7627 (N_7627,N_2972,N_1580);
or U7628 (N_7628,N_2055,N_4415);
or U7629 (N_7629,N_2765,N_909);
xor U7630 (N_7630,N_70,N_1977);
nor U7631 (N_7631,N_1659,N_3457);
or U7632 (N_7632,N_2121,N_4184);
nor U7633 (N_7633,N_4704,N_559);
nor U7634 (N_7634,N_1808,N_2857);
nor U7635 (N_7635,N_2776,N_1459);
or U7636 (N_7636,N_3523,N_4076);
nand U7637 (N_7637,N_3464,N_1473);
or U7638 (N_7638,N_1851,N_884);
and U7639 (N_7639,N_2204,N_2921);
nand U7640 (N_7640,N_3211,N_1142);
xnor U7641 (N_7641,N_3397,N_1875);
nor U7642 (N_7642,N_3896,N_4604);
nand U7643 (N_7643,N_2520,N_1374);
and U7644 (N_7644,N_2594,N_3119);
and U7645 (N_7645,N_118,N_4666);
nand U7646 (N_7646,N_1686,N_302);
nand U7647 (N_7647,N_4202,N_4538);
xor U7648 (N_7648,N_528,N_3706);
nand U7649 (N_7649,N_1013,N_295);
or U7650 (N_7650,N_987,N_3680);
nand U7651 (N_7651,N_4024,N_423);
or U7652 (N_7652,N_3525,N_202);
or U7653 (N_7653,N_4391,N_4668);
nor U7654 (N_7654,N_4214,N_3447);
nor U7655 (N_7655,N_702,N_1336);
or U7656 (N_7656,N_1078,N_1699);
nor U7657 (N_7657,N_1834,N_3811);
nor U7658 (N_7658,N_1391,N_2103);
xor U7659 (N_7659,N_4106,N_4083);
or U7660 (N_7660,N_81,N_313);
or U7661 (N_7661,N_4348,N_2716);
xor U7662 (N_7662,N_2075,N_3942);
nand U7663 (N_7663,N_3062,N_4548);
nor U7664 (N_7664,N_3686,N_100);
and U7665 (N_7665,N_2423,N_2421);
or U7666 (N_7666,N_1827,N_1973);
xor U7667 (N_7667,N_1477,N_4890);
nor U7668 (N_7668,N_885,N_1853);
xor U7669 (N_7669,N_2070,N_2002);
or U7670 (N_7670,N_4818,N_4402);
and U7671 (N_7671,N_1201,N_4706);
nand U7672 (N_7672,N_923,N_1882);
xor U7673 (N_7673,N_329,N_1989);
nor U7674 (N_7674,N_2549,N_4491);
nor U7675 (N_7675,N_1415,N_4974);
or U7676 (N_7676,N_2327,N_4253);
nand U7677 (N_7677,N_1266,N_1699);
nand U7678 (N_7678,N_2739,N_3940);
or U7679 (N_7679,N_4126,N_4643);
xor U7680 (N_7680,N_4362,N_4026);
nand U7681 (N_7681,N_3556,N_3863);
nand U7682 (N_7682,N_4437,N_2712);
and U7683 (N_7683,N_1774,N_2626);
xor U7684 (N_7684,N_3479,N_4224);
nand U7685 (N_7685,N_476,N_4975);
xor U7686 (N_7686,N_4292,N_2985);
and U7687 (N_7687,N_4550,N_1727);
nand U7688 (N_7688,N_2518,N_4381);
or U7689 (N_7689,N_3819,N_3656);
nor U7690 (N_7690,N_851,N_4047);
nand U7691 (N_7691,N_4583,N_226);
and U7692 (N_7692,N_465,N_1908);
or U7693 (N_7693,N_2379,N_3939);
nor U7694 (N_7694,N_383,N_1106);
or U7695 (N_7695,N_454,N_4068);
nor U7696 (N_7696,N_3212,N_608);
or U7697 (N_7697,N_4553,N_2458);
nor U7698 (N_7698,N_939,N_2538);
xor U7699 (N_7699,N_1119,N_679);
or U7700 (N_7700,N_1550,N_39);
nor U7701 (N_7701,N_2184,N_3369);
nor U7702 (N_7702,N_488,N_820);
nor U7703 (N_7703,N_2245,N_3841);
or U7704 (N_7704,N_2996,N_3553);
and U7705 (N_7705,N_1038,N_686);
or U7706 (N_7706,N_572,N_1647);
and U7707 (N_7707,N_2048,N_4593);
and U7708 (N_7708,N_599,N_4939);
xor U7709 (N_7709,N_565,N_2505);
xor U7710 (N_7710,N_4917,N_380);
xor U7711 (N_7711,N_3570,N_1992);
nand U7712 (N_7712,N_1647,N_4044);
and U7713 (N_7713,N_1390,N_4586);
or U7714 (N_7714,N_696,N_4645);
nand U7715 (N_7715,N_4454,N_4530);
nand U7716 (N_7716,N_838,N_1328);
and U7717 (N_7717,N_2708,N_4446);
or U7718 (N_7718,N_535,N_1954);
nand U7719 (N_7719,N_2384,N_3390);
and U7720 (N_7720,N_3184,N_2481);
xor U7721 (N_7721,N_3263,N_1785);
or U7722 (N_7722,N_4317,N_4060);
and U7723 (N_7723,N_2919,N_1515);
nor U7724 (N_7724,N_3289,N_3570);
xnor U7725 (N_7725,N_3664,N_4237);
or U7726 (N_7726,N_541,N_4973);
xnor U7727 (N_7727,N_1157,N_5);
or U7728 (N_7728,N_3185,N_79);
nor U7729 (N_7729,N_1678,N_4680);
and U7730 (N_7730,N_303,N_1729);
or U7731 (N_7731,N_1287,N_2588);
nand U7732 (N_7732,N_992,N_3726);
xor U7733 (N_7733,N_325,N_4937);
nor U7734 (N_7734,N_3621,N_4306);
xnor U7735 (N_7735,N_1400,N_148);
nor U7736 (N_7736,N_841,N_1189);
and U7737 (N_7737,N_4524,N_2920);
nor U7738 (N_7738,N_2553,N_4507);
and U7739 (N_7739,N_4449,N_1820);
nand U7740 (N_7740,N_3414,N_3908);
nor U7741 (N_7741,N_3254,N_3655);
nor U7742 (N_7742,N_1649,N_1260);
nand U7743 (N_7743,N_2077,N_2490);
xnor U7744 (N_7744,N_1701,N_3296);
and U7745 (N_7745,N_658,N_1645);
nor U7746 (N_7746,N_1526,N_3787);
or U7747 (N_7747,N_1159,N_506);
nor U7748 (N_7748,N_1720,N_1196);
or U7749 (N_7749,N_2613,N_3983);
or U7750 (N_7750,N_2929,N_2014);
nor U7751 (N_7751,N_4353,N_1905);
and U7752 (N_7752,N_2916,N_4763);
and U7753 (N_7753,N_2623,N_901);
or U7754 (N_7754,N_2929,N_4394);
and U7755 (N_7755,N_797,N_293);
xnor U7756 (N_7756,N_4574,N_2957);
nand U7757 (N_7757,N_2960,N_1987);
or U7758 (N_7758,N_2514,N_4887);
xnor U7759 (N_7759,N_1882,N_3381);
and U7760 (N_7760,N_4728,N_4062);
and U7761 (N_7761,N_1615,N_4412);
or U7762 (N_7762,N_3878,N_2802);
and U7763 (N_7763,N_54,N_2479);
nand U7764 (N_7764,N_4710,N_2194);
or U7765 (N_7765,N_3247,N_3406);
or U7766 (N_7766,N_3048,N_260);
nand U7767 (N_7767,N_1840,N_3309);
xor U7768 (N_7768,N_4841,N_1576);
nor U7769 (N_7769,N_4729,N_3721);
xnor U7770 (N_7770,N_391,N_1310);
or U7771 (N_7771,N_1457,N_2013);
nand U7772 (N_7772,N_692,N_1075);
xor U7773 (N_7773,N_4365,N_889);
or U7774 (N_7774,N_3830,N_1381);
or U7775 (N_7775,N_2107,N_2467);
and U7776 (N_7776,N_4940,N_526);
xor U7777 (N_7777,N_3461,N_4183);
and U7778 (N_7778,N_2198,N_1018);
nand U7779 (N_7779,N_634,N_804);
or U7780 (N_7780,N_2988,N_2947);
or U7781 (N_7781,N_1421,N_1957);
and U7782 (N_7782,N_3375,N_517);
nand U7783 (N_7783,N_203,N_4939);
xnor U7784 (N_7784,N_943,N_1265);
or U7785 (N_7785,N_2615,N_543);
or U7786 (N_7786,N_4727,N_250);
nor U7787 (N_7787,N_3223,N_1144);
and U7788 (N_7788,N_2427,N_3998);
nand U7789 (N_7789,N_106,N_1855);
nor U7790 (N_7790,N_2302,N_2803);
and U7791 (N_7791,N_4766,N_4910);
and U7792 (N_7792,N_3313,N_3837);
xor U7793 (N_7793,N_3931,N_3920);
or U7794 (N_7794,N_3836,N_4027);
and U7795 (N_7795,N_2596,N_2683);
xnor U7796 (N_7796,N_3625,N_662);
nand U7797 (N_7797,N_2462,N_2426);
or U7798 (N_7798,N_2134,N_941);
xor U7799 (N_7799,N_4293,N_4450);
nand U7800 (N_7800,N_642,N_1581);
and U7801 (N_7801,N_110,N_2371);
and U7802 (N_7802,N_214,N_3592);
xor U7803 (N_7803,N_4514,N_2412);
or U7804 (N_7804,N_2830,N_3889);
or U7805 (N_7805,N_3073,N_2442);
xnor U7806 (N_7806,N_1054,N_2639);
nor U7807 (N_7807,N_3495,N_990);
or U7808 (N_7808,N_3835,N_1132);
and U7809 (N_7809,N_1957,N_4394);
and U7810 (N_7810,N_55,N_1080);
and U7811 (N_7811,N_4190,N_3034);
or U7812 (N_7812,N_4758,N_3839);
nand U7813 (N_7813,N_4198,N_509);
or U7814 (N_7814,N_3516,N_1634);
or U7815 (N_7815,N_2123,N_2457);
and U7816 (N_7816,N_793,N_577);
nor U7817 (N_7817,N_2328,N_4286);
and U7818 (N_7818,N_2477,N_4772);
or U7819 (N_7819,N_390,N_569);
and U7820 (N_7820,N_3205,N_4771);
nor U7821 (N_7821,N_3096,N_1170);
nor U7822 (N_7822,N_1058,N_902);
xor U7823 (N_7823,N_1632,N_1714);
xnor U7824 (N_7824,N_4522,N_3482);
and U7825 (N_7825,N_258,N_4395);
and U7826 (N_7826,N_4351,N_586);
or U7827 (N_7827,N_4901,N_4101);
nand U7828 (N_7828,N_3501,N_2363);
and U7829 (N_7829,N_652,N_4877);
and U7830 (N_7830,N_1708,N_2681);
or U7831 (N_7831,N_1976,N_395);
xnor U7832 (N_7832,N_3220,N_4255);
nor U7833 (N_7833,N_3640,N_2701);
nand U7834 (N_7834,N_3164,N_2509);
nand U7835 (N_7835,N_1265,N_1469);
nor U7836 (N_7836,N_4018,N_1965);
and U7837 (N_7837,N_2178,N_1386);
nor U7838 (N_7838,N_515,N_121);
or U7839 (N_7839,N_2638,N_4911);
xnor U7840 (N_7840,N_326,N_3658);
or U7841 (N_7841,N_3212,N_648);
xnor U7842 (N_7842,N_2223,N_4611);
or U7843 (N_7843,N_374,N_4309);
and U7844 (N_7844,N_4005,N_4042);
nand U7845 (N_7845,N_165,N_3261);
nand U7846 (N_7846,N_2992,N_1855);
or U7847 (N_7847,N_835,N_732);
nand U7848 (N_7848,N_1308,N_3094);
or U7849 (N_7849,N_3642,N_2834);
nor U7850 (N_7850,N_858,N_1976);
and U7851 (N_7851,N_2448,N_1195);
xor U7852 (N_7852,N_3452,N_2802);
xnor U7853 (N_7853,N_4639,N_258);
nor U7854 (N_7854,N_2173,N_956);
or U7855 (N_7855,N_4970,N_4217);
nand U7856 (N_7856,N_870,N_650);
nor U7857 (N_7857,N_1465,N_3340);
nor U7858 (N_7858,N_2689,N_3745);
and U7859 (N_7859,N_4716,N_2293);
or U7860 (N_7860,N_1942,N_2587);
or U7861 (N_7861,N_3912,N_2715);
and U7862 (N_7862,N_455,N_404);
xnor U7863 (N_7863,N_2175,N_256);
nor U7864 (N_7864,N_398,N_4208);
and U7865 (N_7865,N_3756,N_1131);
or U7866 (N_7866,N_4244,N_743);
nor U7867 (N_7867,N_2071,N_398);
nor U7868 (N_7868,N_3120,N_1307);
nor U7869 (N_7869,N_527,N_1982);
nor U7870 (N_7870,N_4560,N_1227);
or U7871 (N_7871,N_3564,N_2910);
or U7872 (N_7872,N_198,N_3353);
nand U7873 (N_7873,N_762,N_0);
and U7874 (N_7874,N_2039,N_1061);
nand U7875 (N_7875,N_258,N_2383);
or U7876 (N_7876,N_4472,N_2262);
xnor U7877 (N_7877,N_4268,N_1480);
nor U7878 (N_7878,N_1254,N_3287);
nor U7879 (N_7879,N_2376,N_1963);
nand U7880 (N_7880,N_1164,N_2481);
or U7881 (N_7881,N_2103,N_457);
or U7882 (N_7882,N_4801,N_4160);
or U7883 (N_7883,N_2528,N_1720);
nor U7884 (N_7884,N_3621,N_1648);
and U7885 (N_7885,N_2926,N_2883);
xnor U7886 (N_7886,N_4098,N_4703);
nand U7887 (N_7887,N_4125,N_1755);
or U7888 (N_7888,N_3896,N_1691);
nor U7889 (N_7889,N_4296,N_3266);
or U7890 (N_7890,N_4342,N_3744);
and U7891 (N_7891,N_3534,N_3162);
and U7892 (N_7892,N_1712,N_1590);
nand U7893 (N_7893,N_4746,N_2891);
and U7894 (N_7894,N_4099,N_4936);
xor U7895 (N_7895,N_3331,N_811);
or U7896 (N_7896,N_4816,N_318);
nand U7897 (N_7897,N_4699,N_4819);
and U7898 (N_7898,N_2113,N_577);
nand U7899 (N_7899,N_1771,N_4566);
and U7900 (N_7900,N_3732,N_615);
and U7901 (N_7901,N_3843,N_2348);
or U7902 (N_7902,N_4026,N_1646);
xnor U7903 (N_7903,N_4101,N_56);
or U7904 (N_7904,N_587,N_4704);
nor U7905 (N_7905,N_4740,N_3276);
xor U7906 (N_7906,N_805,N_3319);
nand U7907 (N_7907,N_395,N_4046);
xnor U7908 (N_7908,N_2742,N_2186);
or U7909 (N_7909,N_4137,N_2085);
and U7910 (N_7910,N_1823,N_934);
and U7911 (N_7911,N_4336,N_3690);
xor U7912 (N_7912,N_122,N_3086);
or U7913 (N_7913,N_1122,N_2633);
and U7914 (N_7914,N_4350,N_4195);
nand U7915 (N_7915,N_2410,N_907);
xnor U7916 (N_7916,N_3983,N_1925);
nand U7917 (N_7917,N_3495,N_3046);
nor U7918 (N_7918,N_2993,N_3094);
or U7919 (N_7919,N_1763,N_540);
nand U7920 (N_7920,N_4952,N_929);
and U7921 (N_7921,N_2654,N_3196);
xor U7922 (N_7922,N_1697,N_2548);
xnor U7923 (N_7923,N_1177,N_3025);
nand U7924 (N_7924,N_3672,N_4160);
xor U7925 (N_7925,N_3186,N_1984);
nand U7926 (N_7926,N_3196,N_794);
and U7927 (N_7927,N_1368,N_1533);
nand U7928 (N_7928,N_201,N_1803);
xnor U7929 (N_7929,N_2350,N_2528);
or U7930 (N_7930,N_3303,N_2353);
or U7931 (N_7931,N_3711,N_1703);
xor U7932 (N_7932,N_3704,N_3785);
and U7933 (N_7933,N_3213,N_3583);
nor U7934 (N_7934,N_4679,N_2577);
xor U7935 (N_7935,N_3724,N_1525);
and U7936 (N_7936,N_17,N_258);
nand U7937 (N_7937,N_2405,N_3027);
nand U7938 (N_7938,N_2603,N_1552);
or U7939 (N_7939,N_2089,N_1346);
nand U7940 (N_7940,N_2636,N_4655);
xor U7941 (N_7941,N_390,N_61);
nor U7942 (N_7942,N_2966,N_4707);
and U7943 (N_7943,N_3970,N_2232);
nand U7944 (N_7944,N_4215,N_4046);
nor U7945 (N_7945,N_2745,N_4809);
or U7946 (N_7946,N_1679,N_978);
or U7947 (N_7947,N_2279,N_4358);
nand U7948 (N_7948,N_789,N_549);
nand U7949 (N_7949,N_3349,N_1232);
nor U7950 (N_7950,N_2650,N_1435);
nor U7951 (N_7951,N_1598,N_4285);
or U7952 (N_7952,N_2174,N_1290);
nor U7953 (N_7953,N_4733,N_3989);
and U7954 (N_7954,N_448,N_1853);
or U7955 (N_7955,N_2422,N_732);
or U7956 (N_7956,N_848,N_2187);
nor U7957 (N_7957,N_3230,N_297);
or U7958 (N_7958,N_2999,N_735);
nand U7959 (N_7959,N_1865,N_3205);
xnor U7960 (N_7960,N_343,N_27);
xor U7961 (N_7961,N_3331,N_4411);
nor U7962 (N_7962,N_326,N_3031);
nor U7963 (N_7963,N_583,N_1862);
nand U7964 (N_7964,N_8,N_2160);
and U7965 (N_7965,N_3236,N_3989);
xor U7966 (N_7966,N_3980,N_1340);
nand U7967 (N_7967,N_889,N_435);
or U7968 (N_7968,N_87,N_1803);
nor U7969 (N_7969,N_1248,N_551);
and U7970 (N_7970,N_3383,N_2749);
or U7971 (N_7971,N_4569,N_3774);
nand U7972 (N_7972,N_1746,N_83);
and U7973 (N_7973,N_3472,N_1242);
xor U7974 (N_7974,N_4372,N_1790);
nor U7975 (N_7975,N_255,N_56);
or U7976 (N_7976,N_3696,N_4768);
or U7977 (N_7977,N_3944,N_3891);
xor U7978 (N_7978,N_2510,N_2844);
and U7979 (N_7979,N_4121,N_3664);
xor U7980 (N_7980,N_378,N_2903);
nor U7981 (N_7981,N_4263,N_22);
and U7982 (N_7982,N_3579,N_263);
xor U7983 (N_7983,N_2305,N_2331);
nor U7984 (N_7984,N_1765,N_1109);
nor U7985 (N_7985,N_2337,N_588);
or U7986 (N_7986,N_438,N_2345);
and U7987 (N_7987,N_973,N_3257);
or U7988 (N_7988,N_4733,N_3582);
nor U7989 (N_7989,N_3020,N_2633);
nand U7990 (N_7990,N_2388,N_1591);
or U7991 (N_7991,N_4111,N_3170);
xor U7992 (N_7992,N_477,N_3544);
nor U7993 (N_7993,N_1258,N_3855);
and U7994 (N_7994,N_3354,N_4061);
xor U7995 (N_7995,N_2861,N_2629);
nand U7996 (N_7996,N_1288,N_1090);
xnor U7997 (N_7997,N_4952,N_3246);
or U7998 (N_7998,N_1679,N_665);
or U7999 (N_7999,N_1806,N_4353);
and U8000 (N_8000,N_218,N_1214);
or U8001 (N_8001,N_4139,N_2062);
and U8002 (N_8002,N_1179,N_855);
xnor U8003 (N_8003,N_2189,N_1725);
nand U8004 (N_8004,N_2684,N_3174);
nand U8005 (N_8005,N_4485,N_3017);
xor U8006 (N_8006,N_2811,N_2910);
xor U8007 (N_8007,N_704,N_1696);
nor U8008 (N_8008,N_2073,N_4613);
xnor U8009 (N_8009,N_3870,N_42);
xnor U8010 (N_8010,N_1626,N_4994);
xor U8011 (N_8011,N_2137,N_4669);
and U8012 (N_8012,N_1441,N_1018);
nand U8013 (N_8013,N_4494,N_56);
or U8014 (N_8014,N_2200,N_2056);
nand U8015 (N_8015,N_2265,N_3334);
nor U8016 (N_8016,N_66,N_2993);
nand U8017 (N_8017,N_2299,N_3597);
xnor U8018 (N_8018,N_1539,N_4886);
nand U8019 (N_8019,N_1219,N_1525);
nor U8020 (N_8020,N_25,N_3463);
nand U8021 (N_8021,N_2381,N_42);
or U8022 (N_8022,N_245,N_4200);
xnor U8023 (N_8023,N_931,N_2927);
and U8024 (N_8024,N_3009,N_3052);
nand U8025 (N_8025,N_866,N_4760);
nor U8026 (N_8026,N_3431,N_264);
nor U8027 (N_8027,N_213,N_743);
xor U8028 (N_8028,N_2480,N_2976);
and U8029 (N_8029,N_4676,N_3326);
or U8030 (N_8030,N_3337,N_1885);
and U8031 (N_8031,N_3743,N_2900);
nand U8032 (N_8032,N_1148,N_4180);
nand U8033 (N_8033,N_2204,N_4545);
nand U8034 (N_8034,N_4318,N_3347);
nand U8035 (N_8035,N_2867,N_4079);
nand U8036 (N_8036,N_709,N_1917);
and U8037 (N_8037,N_1374,N_2836);
xnor U8038 (N_8038,N_1335,N_3795);
and U8039 (N_8039,N_1567,N_685);
nand U8040 (N_8040,N_4421,N_640);
nor U8041 (N_8041,N_1382,N_4144);
nand U8042 (N_8042,N_2761,N_715);
nor U8043 (N_8043,N_4766,N_1108);
nor U8044 (N_8044,N_2716,N_3766);
or U8045 (N_8045,N_3589,N_3508);
nor U8046 (N_8046,N_1297,N_4817);
xor U8047 (N_8047,N_872,N_3490);
nor U8048 (N_8048,N_2495,N_652);
nor U8049 (N_8049,N_3264,N_2113);
or U8050 (N_8050,N_2662,N_3550);
nor U8051 (N_8051,N_2018,N_1236);
nand U8052 (N_8052,N_436,N_4808);
nor U8053 (N_8053,N_394,N_1825);
or U8054 (N_8054,N_2069,N_1643);
nand U8055 (N_8055,N_4108,N_3804);
or U8056 (N_8056,N_4607,N_749);
nand U8057 (N_8057,N_330,N_1254);
nand U8058 (N_8058,N_98,N_577);
xor U8059 (N_8059,N_66,N_4170);
and U8060 (N_8060,N_826,N_3382);
nand U8061 (N_8061,N_486,N_4653);
nor U8062 (N_8062,N_362,N_4893);
and U8063 (N_8063,N_3134,N_1037);
or U8064 (N_8064,N_3326,N_1795);
nand U8065 (N_8065,N_2973,N_4775);
and U8066 (N_8066,N_2957,N_3642);
or U8067 (N_8067,N_4074,N_3703);
and U8068 (N_8068,N_2006,N_2986);
or U8069 (N_8069,N_1252,N_631);
nor U8070 (N_8070,N_2240,N_2211);
and U8071 (N_8071,N_2178,N_1819);
nor U8072 (N_8072,N_4237,N_1490);
or U8073 (N_8073,N_2718,N_1135);
and U8074 (N_8074,N_2401,N_1180);
and U8075 (N_8075,N_1465,N_3372);
nand U8076 (N_8076,N_4633,N_1102);
nand U8077 (N_8077,N_527,N_1976);
nand U8078 (N_8078,N_3689,N_3551);
xor U8079 (N_8079,N_2784,N_126);
and U8080 (N_8080,N_2660,N_3292);
nand U8081 (N_8081,N_4410,N_220);
xor U8082 (N_8082,N_71,N_3829);
and U8083 (N_8083,N_658,N_3741);
xor U8084 (N_8084,N_2202,N_1799);
xnor U8085 (N_8085,N_4918,N_4878);
or U8086 (N_8086,N_3741,N_3829);
or U8087 (N_8087,N_3819,N_3349);
nor U8088 (N_8088,N_3227,N_1339);
nor U8089 (N_8089,N_3369,N_970);
or U8090 (N_8090,N_3028,N_1678);
or U8091 (N_8091,N_3906,N_975);
and U8092 (N_8092,N_4954,N_4112);
xor U8093 (N_8093,N_3953,N_1801);
nor U8094 (N_8094,N_2766,N_4323);
nor U8095 (N_8095,N_2180,N_1138);
xnor U8096 (N_8096,N_3053,N_1313);
nand U8097 (N_8097,N_3869,N_3068);
nor U8098 (N_8098,N_4147,N_34);
xor U8099 (N_8099,N_2261,N_1507);
nor U8100 (N_8100,N_3603,N_861);
xor U8101 (N_8101,N_4394,N_4177);
nor U8102 (N_8102,N_2090,N_2639);
nor U8103 (N_8103,N_2954,N_154);
nand U8104 (N_8104,N_4816,N_2901);
nand U8105 (N_8105,N_1957,N_3623);
or U8106 (N_8106,N_4755,N_3705);
and U8107 (N_8107,N_4709,N_4882);
nand U8108 (N_8108,N_2041,N_3108);
xor U8109 (N_8109,N_3439,N_2407);
xnor U8110 (N_8110,N_732,N_1736);
and U8111 (N_8111,N_2220,N_3742);
nand U8112 (N_8112,N_2103,N_1714);
nor U8113 (N_8113,N_2937,N_3077);
or U8114 (N_8114,N_4657,N_500);
nand U8115 (N_8115,N_1130,N_450);
nor U8116 (N_8116,N_1453,N_3498);
xor U8117 (N_8117,N_3310,N_4112);
or U8118 (N_8118,N_4896,N_1678);
nand U8119 (N_8119,N_3524,N_2783);
or U8120 (N_8120,N_4533,N_2713);
nor U8121 (N_8121,N_4006,N_2614);
nor U8122 (N_8122,N_539,N_2433);
nor U8123 (N_8123,N_2554,N_2109);
nand U8124 (N_8124,N_1791,N_2659);
and U8125 (N_8125,N_4204,N_791);
nand U8126 (N_8126,N_3056,N_4182);
nand U8127 (N_8127,N_2015,N_4807);
or U8128 (N_8128,N_2060,N_1240);
xnor U8129 (N_8129,N_2626,N_3273);
nor U8130 (N_8130,N_752,N_3320);
nand U8131 (N_8131,N_4264,N_3460);
nand U8132 (N_8132,N_2733,N_1809);
nand U8133 (N_8133,N_116,N_1745);
or U8134 (N_8134,N_1260,N_4678);
nor U8135 (N_8135,N_2746,N_599);
and U8136 (N_8136,N_4730,N_3944);
nor U8137 (N_8137,N_2865,N_1466);
or U8138 (N_8138,N_3454,N_1134);
xor U8139 (N_8139,N_4216,N_3716);
nand U8140 (N_8140,N_1213,N_3619);
and U8141 (N_8141,N_3080,N_4560);
nor U8142 (N_8142,N_1871,N_1372);
nand U8143 (N_8143,N_3543,N_4329);
nor U8144 (N_8144,N_1809,N_4321);
nor U8145 (N_8145,N_4901,N_2813);
and U8146 (N_8146,N_1513,N_2419);
or U8147 (N_8147,N_799,N_1750);
and U8148 (N_8148,N_417,N_1223);
and U8149 (N_8149,N_996,N_693);
and U8150 (N_8150,N_907,N_4803);
nand U8151 (N_8151,N_3639,N_2175);
nor U8152 (N_8152,N_4559,N_2298);
xor U8153 (N_8153,N_4223,N_2197);
nor U8154 (N_8154,N_641,N_932);
and U8155 (N_8155,N_1424,N_4931);
or U8156 (N_8156,N_2731,N_4198);
xnor U8157 (N_8157,N_3685,N_3324);
and U8158 (N_8158,N_3876,N_3520);
nand U8159 (N_8159,N_3982,N_35);
and U8160 (N_8160,N_124,N_3337);
xor U8161 (N_8161,N_3736,N_3115);
nor U8162 (N_8162,N_2366,N_1502);
xor U8163 (N_8163,N_1268,N_1154);
xor U8164 (N_8164,N_4780,N_44);
nor U8165 (N_8165,N_1331,N_4107);
nor U8166 (N_8166,N_1717,N_2809);
and U8167 (N_8167,N_959,N_3118);
or U8168 (N_8168,N_2535,N_2718);
nand U8169 (N_8169,N_2761,N_3981);
and U8170 (N_8170,N_3387,N_1588);
or U8171 (N_8171,N_4340,N_2695);
nand U8172 (N_8172,N_4349,N_2380);
and U8173 (N_8173,N_4454,N_4199);
and U8174 (N_8174,N_782,N_2522);
nand U8175 (N_8175,N_2003,N_4206);
xnor U8176 (N_8176,N_3286,N_4915);
or U8177 (N_8177,N_1530,N_1593);
nand U8178 (N_8178,N_3845,N_1165);
nand U8179 (N_8179,N_2462,N_4828);
xnor U8180 (N_8180,N_3161,N_4605);
xnor U8181 (N_8181,N_3275,N_4802);
and U8182 (N_8182,N_1387,N_1663);
and U8183 (N_8183,N_2089,N_184);
nor U8184 (N_8184,N_3582,N_731);
nand U8185 (N_8185,N_2424,N_2099);
nand U8186 (N_8186,N_4052,N_4622);
and U8187 (N_8187,N_2937,N_2466);
nand U8188 (N_8188,N_4305,N_3674);
and U8189 (N_8189,N_3688,N_4423);
xor U8190 (N_8190,N_313,N_4306);
or U8191 (N_8191,N_2290,N_1236);
and U8192 (N_8192,N_3370,N_2590);
or U8193 (N_8193,N_2599,N_4981);
nor U8194 (N_8194,N_2309,N_3891);
nand U8195 (N_8195,N_3987,N_1780);
and U8196 (N_8196,N_2456,N_2735);
xor U8197 (N_8197,N_707,N_999);
or U8198 (N_8198,N_3586,N_2638);
nor U8199 (N_8199,N_1836,N_400);
and U8200 (N_8200,N_3394,N_1662);
or U8201 (N_8201,N_3893,N_1867);
xnor U8202 (N_8202,N_3260,N_4723);
or U8203 (N_8203,N_3839,N_2422);
xor U8204 (N_8204,N_3609,N_4161);
and U8205 (N_8205,N_4276,N_4186);
and U8206 (N_8206,N_4108,N_31);
or U8207 (N_8207,N_3676,N_1056);
and U8208 (N_8208,N_857,N_2994);
xor U8209 (N_8209,N_3762,N_3085);
or U8210 (N_8210,N_1774,N_4505);
nor U8211 (N_8211,N_2754,N_3203);
nor U8212 (N_8212,N_2765,N_3161);
and U8213 (N_8213,N_348,N_122);
or U8214 (N_8214,N_2049,N_2591);
nor U8215 (N_8215,N_3404,N_3325);
xnor U8216 (N_8216,N_3761,N_1364);
xor U8217 (N_8217,N_918,N_7);
xor U8218 (N_8218,N_1317,N_1681);
nand U8219 (N_8219,N_3536,N_2773);
xnor U8220 (N_8220,N_2961,N_1444);
xnor U8221 (N_8221,N_2444,N_1849);
xnor U8222 (N_8222,N_167,N_2231);
nand U8223 (N_8223,N_3544,N_2549);
xnor U8224 (N_8224,N_754,N_3532);
nand U8225 (N_8225,N_382,N_1641);
and U8226 (N_8226,N_3530,N_1922);
xnor U8227 (N_8227,N_4997,N_3302);
or U8228 (N_8228,N_2199,N_1684);
nand U8229 (N_8229,N_3370,N_2025);
xor U8230 (N_8230,N_3139,N_1763);
or U8231 (N_8231,N_3949,N_2104);
and U8232 (N_8232,N_3950,N_3171);
or U8233 (N_8233,N_475,N_4108);
and U8234 (N_8234,N_2468,N_3329);
xor U8235 (N_8235,N_2293,N_2675);
and U8236 (N_8236,N_4199,N_4326);
and U8237 (N_8237,N_4819,N_108);
and U8238 (N_8238,N_1478,N_2618);
nor U8239 (N_8239,N_663,N_3686);
nor U8240 (N_8240,N_177,N_95);
or U8241 (N_8241,N_1662,N_1587);
nor U8242 (N_8242,N_170,N_4262);
xnor U8243 (N_8243,N_4718,N_1211);
nand U8244 (N_8244,N_4122,N_4629);
nand U8245 (N_8245,N_2756,N_612);
xor U8246 (N_8246,N_714,N_2908);
nor U8247 (N_8247,N_3316,N_899);
or U8248 (N_8248,N_997,N_4703);
nand U8249 (N_8249,N_4010,N_2995);
xor U8250 (N_8250,N_1425,N_125);
nand U8251 (N_8251,N_1205,N_1639);
and U8252 (N_8252,N_4878,N_3355);
nand U8253 (N_8253,N_1094,N_715);
xnor U8254 (N_8254,N_10,N_698);
nand U8255 (N_8255,N_3379,N_3989);
or U8256 (N_8256,N_3850,N_3421);
xor U8257 (N_8257,N_3295,N_4694);
nor U8258 (N_8258,N_102,N_1504);
xor U8259 (N_8259,N_4804,N_4518);
nor U8260 (N_8260,N_4577,N_2434);
and U8261 (N_8261,N_4205,N_2843);
nor U8262 (N_8262,N_3864,N_2197);
and U8263 (N_8263,N_4122,N_3122);
or U8264 (N_8264,N_1708,N_1228);
and U8265 (N_8265,N_2843,N_4928);
and U8266 (N_8266,N_1220,N_4389);
nor U8267 (N_8267,N_489,N_361);
xnor U8268 (N_8268,N_2383,N_3843);
nand U8269 (N_8269,N_265,N_4460);
or U8270 (N_8270,N_134,N_1519);
and U8271 (N_8271,N_3377,N_4863);
nor U8272 (N_8272,N_4976,N_1922);
xnor U8273 (N_8273,N_4253,N_3130);
nand U8274 (N_8274,N_875,N_606);
xnor U8275 (N_8275,N_4719,N_2604);
nor U8276 (N_8276,N_1730,N_2265);
or U8277 (N_8277,N_875,N_1391);
or U8278 (N_8278,N_793,N_4557);
nand U8279 (N_8279,N_1021,N_2434);
or U8280 (N_8280,N_4763,N_2683);
xor U8281 (N_8281,N_3685,N_1537);
xnor U8282 (N_8282,N_472,N_1694);
nor U8283 (N_8283,N_1461,N_953);
or U8284 (N_8284,N_4282,N_1780);
nor U8285 (N_8285,N_2912,N_3417);
xor U8286 (N_8286,N_3619,N_2929);
and U8287 (N_8287,N_2164,N_3353);
xnor U8288 (N_8288,N_2979,N_4970);
nand U8289 (N_8289,N_1170,N_616);
xnor U8290 (N_8290,N_3490,N_239);
nor U8291 (N_8291,N_2341,N_2677);
nand U8292 (N_8292,N_3943,N_2110);
xor U8293 (N_8293,N_1126,N_4818);
and U8294 (N_8294,N_2311,N_182);
and U8295 (N_8295,N_518,N_289);
nor U8296 (N_8296,N_235,N_3446);
xnor U8297 (N_8297,N_3089,N_3772);
nor U8298 (N_8298,N_1482,N_3055);
xor U8299 (N_8299,N_2167,N_3463);
nor U8300 (N_8300,N_10,N_2600);
and U8301 (N_8301,N_3736,N_1427);
and U8302 (N_8302,N_1216,N_3322);
nand U8303 (N_8303,N_496,N_2316);
xor U8304 (N_8304,N_207,N_560);
nor U8305 (N_8305,N_362,N_1359);
and U8306 (N_8306,N_214,N_2793);
or U8307 (N_8307,N_4735,N_1292);
nor U8308 (N_8308,N_3542,N_2445);
xor U8309 (N_8309,N_1644,N_185);
nor U8310 (N_8310,N_3096,N_3581);
and U8311 (N_8311,N_100,N_3221);
nor U8312 (N_8312,N_4889,N_186);
or U8313 (N_8313,N_116,N_3060);
nand U8314 (N_8314,N_3811,N_4028);
nand U8315 (N_8315,N_1040,N_2515);
nand U8316 (N_8316,N_19,N_3393);
xor U8317 (N_8317,N_4253,N_1138);
xor U8318 (N_8318,N_3781,N_1226);
nand U8319 (N_8319,N_2309,N_443);
nor U8320 (N_8320,N_2331,N_1240);
or U8321 (N_8321,N_2258,N_1721);
or U8322 (N_8322,N_4447,N_2725);
and U8323 (N_8323,N_3405,N_1501);
or U8324 (N_8324,N_1327,N_282);
nor U8325 (N_8325,N_4586,N_4317);
nand U8326 (N_8326,N_1780,N_3736);
and U8327 (N_8327,N_4838,N_3436);
nand U8328 (N_8328,N_2825,N_2266);
or U8329 (N_8329,N_1495,N_3064);
and U8330 (N_8330,N_3157,N_4855);
or U8331 (N_8331,N_103,N_1613);
nor U8332 (N_8332,N_1425,N_4400);
and U8333 (N_8333,N_3132,N_4043);
or U8334 (N_8334,N_1682,N_2224);
xor U8335 (N_8335,N_1172,N_3174);
nand U8336 (N_8336,N_1054,N_4063);
nor U8337 (N_8337,N_4362,N_788);
nand U8338 (N_8338,N_4168,N_3578);
or U8339 (N_8339,N_1923,N_4199);
or U8340 (N_8340,N_761,N_2284);
nor U8341 (N_8341,N_801,N_2717);
xnor U8342 (N_8342,N_1992,N_2864);
nand U8343 (N_8343,N_2643,N_4298);
xnor U8344 (N_8344,N_3524,N_2719);
nor U8345 (N_8345,N_4645,N_2464);
xnor U8346 (N_8346,N_585,N_4896);
or U8347 (N_8347,N_2431,N_3201);
and U8348 (N_8348,N_842,N_1780);
and U8349 (N_8349,N_1463,N_492);
nor U8350 (N_8350,N_4592,N_4216);
nor U8351 (N_8351,N_2910,N_2779);
nand U8352 (N_8352,N_3724,N_872);
and U8353 (N_8353,N_2323,N_1347);
nand U8354 (N_8354,N_1925,N_689);
or U8355 (N_8355,N_1230,N_1015);
or U8356 (N_8356,N_2738,N_2714);
or U8357 (N_8357,N_3466,N_2180);
nand U8358 (N_8358,N_573,N_4571);
xor U8359 (N_8359,N_2810,N_4935);
nor U8360 (N_8360,N_3064,N_3050);
nor U8361 (N_8361,N_26,N_2623);
nor U8362 (N_8362,N_512,N_1620);
and U8363 (N_8363,N_1152,N_4189);
xor U8364 (N_8364,N_2333,N_3264);
nor U8365 (N_8365,N_2506,N_3307);
nor U8366 (N_8366,N_3319,N_959);
xor U8367 (N_8367,N_4349,N_4105);
nand U8368 (N_8368,N_3775,N_493);
xnor U8369 (N_8369,N_4501,N_2428);
xnor U8370 (N_8370,N_2057,N_4040);
and U8371 (N_8371,N_2929,N_2354);
or U8372 (N_8372,N_1067,N_2727);
nor U8373 (N_8373,N_812,N_4315);
and U8374 (N_8374,N_1160,N_2325);
nand U8375 (N_8375,N_664,N_454);
and U8376 (N_8376,N_3783,N_646);
nand U8377 (N_8377,N_3547,N_2766);
or U8378 (N_8378,N_2433,N_3280);
nor U8379 (N_8379,N_2006,N_4767);
and U8380 (N_8380,N_3020,N_2297);
or U8381 (N_8381,N_382,N_1170);
or U8382 (N_8382,N_1689,N_1317);
or U8383 (N_8383,N_4212,N_3741);
nor U8384 (N_8384,N_4765,N_1684);
and U8385 (N_8385,N_4155,N_2114);
and U8386 (N_8386,N_3386,N_591);
xnor U8387 (N_8387,N_1245,N_1617);
and U8388 (N_8388,N_4140,N_3938);
nor U8389 (N_8389,N_4195,N_201);
xor U8390 (N_8390,N_2257,N_248);
nand U8391 (N_8391,N_2448,N_1183);
nand U8392 (N_8392,N_3225,N_2810);
xor U8393 (N_8393,N_2127,N_645);
and U8394 (N_8394,N_2891,N_3332);
nor U8395 (N_8395,N_3184,N_2891);
and U8396 (N_8396,N_3119,N_3927);
xnor U8397 (N_8397,N_2164,N_3649);
xnor U8398 (N_8398,N_2634,N_820);
xnor U8399 (N_8399,N_3969,N_3454);
nand U8400 (N_8400,N_255,N_4077);
or U8401 (N_8401,N_469,N_4329);
and U8402 (N_8402,N_3202,N_4436);
xor U8403 (N_8403,N_4111,N_929);
xnor U8404 (N_8404,N_2556,N_2517);
and U8405 (N_8405,N_2927,N_1652);
nand U8406 (N_8406,N_204,N_4239);
nor U8407 (N_8407,N_1306,N_500);
nor U8408 (N_8408,N_4352,N_2633);
nor U8409 (N_8409,N_3826,N_3254);
and U8410 (N_8410,N_574,N_177);
or U8411 (N_8411,N_1756,N_1471);
and U8412 (N_8412,N_2375,N_2528);
xor U8413 (N_8413,N_3475,N_2924);
nor U8414 (N_8414,N_4242,N_2550);
or U8415 (N_8415,N_4862,N_4562);
nand U8416 (N_8416,N_2770,N_2940);
nand U8417 (N_8417,N_4259,N_3275);
and U8418 (N_8418,N_615,N_4536);
or U8419 (N_8419,N_3176,N_78);
nand U8420 (N_8420,N_2041,N_4085);
nand U8421 (N_8421,N_2497,N_1909);
nand U8422 (N_8422,N_260,N_87);
and U8423 (N_8423,N_4664,N_3355);
xor U8424 (N_8424,N_254,N_2561);
or U8425 (N_8425,N_2704,N_2105);
xnor U8426 (N_8426,N_1319,N_1685);
and U8427 (N_8427,N_4667,N_4549);
and U8428 (N_8428,N_1896,N_2073);
nand U8429 (N_8429,N_1554,N_293);
nor U8430 (N_8430,N_3668,N_2172);
nand U8431 (N_8431,N_1893,N_4341);
xor U8432 (N_8432,N_2267,N_887);
nand U8433 (N_8433,N_3378,N_4991);
xnor U8434 (N_8434,N_3654,N_517);
and U8435 (N_8435,N_1469,N_3294);
nor U8436 (N_8436,N_2941,N_3889);
xnor U8437 (N_8437,N_1332,N_1911);
nand U8438 (N_8438,N_4463,N_3842);
nor U8439 (N_8439,N_2059,N_2351);
or U8440 (N_8440,N_474,N_4526);
or U8441 (N_8441,N_883,N_1300);
or U8442 (N_8442,N_1869,N_1321);
nand U8443 (N_8443,N_115,N_1459);
nor U8444 (N_8444,N_1825,N_1037);
nor U8445 (N_8445,N_3706,N_1993);
or U8446 (N_8446,N_1947,N_2885);
nor U8447 (N_8447,N_3896,N_3764);
or U8448 (N_8448,N_2192,N_631);
nor U8449 (N_8449,N_1915,N_1389);
xor U8450 (N_8450,N_3337,N_513);
or U8451 (N_8451,N_1962,N_1682);
nand U8452 (N_8452,N_1091,N_2790);
xor U8453 (N_8453,N_2099,N_1358);
nor U8454 (N_8454,N_4472,N_1396);
and U8455 (N_8455,N_4363,N_4351);
nand U8456 (N_8456,N_1730,N_625);
or U8457 (N_8457,N_3253,N_2887);
nand U8458 (N_8458,N_2486,N_4346);
nand U8459 (N_8459,N_1503,N_3765);
xor U8460 (N_8460,N_3943,N_1321);
nand U8461 (N_8461,N_943,N_1425);
and U8462 (N_8462,N_505,N_3081);
nor U8463 (N_8463,N_3793,N_2559);
xor U8464 (N_8464,N_3362,N_275);
nand U8465 (N_8465,N_3995,N_191);
xor U8466 (N_8466,N_1535,N_2168);
or U8467 (N_8467,N_3293,N_323);
and U8468 (N_8468,N_4815,N_612);
and U8469 (N_8469,N_3797,N_2162);
nand U8470 (N_8470,N_2988,N_1429);
nand U8471 (N_8471,N_922,N_4512);
and U8472 (N_8472,N_3898,N_197);
and U8473 (N_8473,N_2164,N_4299);
nor U8474 (N_8474,N_3561,N_3532);
or U8475 (N_8475,N_2987,N_1558);
nand U8476 (N_8476,N_3372,N_1871);
nand U8477 (N_8477,N_1695,N_4748);
nand U8478 (N_8478,N_4419,N_3828);
and U8479 (N_8479,N_4894,N_3236);
or U8480 (N_8480,N_4718,N_1781);
nand U8481 (N_8481,N_150,N_122);
and U8482 (N_8482,N_2867,N_3793);
nand U8483 (N_8483,N_2891,N_624);
or U8484 (N_8484,N_2981,N_4754);
nand U8485 (N_8485,N_2039,N_4883);
nand U8486 (N_8486,N_3964,N_3556);
and U8487 (N_8487,N_2730,N_3101);
nand U8488 (N_8488,N_3536,N_2557);
and U8489 (N_8489,N_335,N_2156);
and U8490 (N_8490,N_4877,N_2243);
nand U8491 (N_8491,N_1124,N_3962);
and U8492 (N_8492,N_2035,N_3978);
nor U8493 (N_8493,N_1992,N_197);
nor U8494 (N_8494,N_226,N_1028);
xnor U8495 (N_8495,N_2813,N_4308);
xor U8496 (N_8496,N_2044,N_3439);
or U8497 (N_8497,N_2168,N_514);
nand U8498 (N_8498,N_3196,N_2312);
or U8499 (N_8499,N_3288,N_694);
nand U8500 (N_8500,N_1914,N_3957);
xor U8501 (N_8501,N_1948,N_936);
and U8502 (N_8502,N_4738,N_2690);
and U8503 (N_8503,N_1617,N_3880);
and U8504 (N_8504,N_1565,N_1953);
nor U8505 (N_8505,N_2466,N_3431);
or U8506 (N_8506,N_3369,N_340);
or U8507 (N_8507,N_3983,N_452);
or U8508 (N_8508,N_4663,N_3041);
xnor U8509 (N_8509,N_1832,N_3537);
nor U8510 (N_8510,N_705,N_4926);
nand U8511 (N_8511,N_792,N_595);
xor U8512 (N_8512,N_886,N_3005);
nand U8513 (N_8513,N_3292,N_3694);
nor U8514 (N_8514,N_4276,N_3283);
or U8515 (N_8515,N_332,N_1527);
or U8516 (N_8516,N_3885,N_528);
nand U8517 (N_8517,N_4564,N_3780);
nand U8518 (N_8518,N_2111,N_3699);
nand U8519 (N_8519,N_275,N_3325);
or U8520 (N_8520,N_1744,N_3247);
nor U8521 (N_8521,N_4464,N_4715);
xor U8522 (N_8522,N_3692,N_3083);
xnor U8523 (N_8523,N_2976,N_2816);
nand U8524 (N_8524,N_2393,N_3622);
xor U8525 (N_8525,N_4812,N_4232);
xnor U8526 (N_8526,N_4132,N_3237);
or U8527 (N_8527,N_4217,N_1449);
nor U8528 (N_8528,N_2021,N_145);
and U8529 (N_8529,N_2499,N_3116);
nand U8530 (N_8530,N_4833,N_1233);
xnor U8531 (N_8531,N_2114,N_2666);
and U8532 (N_8532,N_1598,N_1768);
or U8533 (N_8533,N_350,N_4641);
nand U8534 (N_8534,N_660,N_3594);
xor U8535 (N_8535,N_3207,N_638);
nor U8536 (N_8536,N_1321,N_2522);
xor U8537 (N_8537,N_328,N_3376);
nor U8538 (N_8538,N_418,N_603);
nand U8539 (N_8539,N_1397,N_3002);
nor U8540 (N_8540,N_2007,N_1736);
and U8541 (N_8541,N_483,N_683);
xor U8542 (N_8542,N_1174,N_4819);
or U8543 (N_8543,N_4317,N_1110);
nor U8544 (N_8544,N_1174,N_4568);
xor U8545 (N_8545,N_4703,N_592);
nand U8546 (N_8546,N_3082,N_2279);
and U8547 (N_8547,N_2842,N_91);
and U8548 (N_8548,N_4019,N_1642);
or U8549 (N_8549,N_2213,N_3163);
or U8550 (N_8550,N_902,N_2061);
xnor U8551 (N_8551,N_437,N_3061);
nand U8552 (N_8552,N_4272,N_4938);
or U8553 (N_8553,N_1815,N_3205);
and U8554 (N_8554,N_4942,N_1053);
nor U8555 (N_8555,N_3493,N_3487);
and U8556 (N_8556,N_1504,N_3927);
and U8557 (N_8557,N_127,N_1273);
and U8558 (N_8558,N_1289,N_3632);
nor U8559 (N_8559,N_4188,N_982);
nor U8560 (N_8560,N_807,N_3925);
or U8561 (N_8561,N_4931,N_2646);
nand U8562 (N_8562,N_4268,N_479);
and U8563 (N_8563,N_526,N_1289);
nor U8564 (N_8564,N_3336,N_2113);
and U8565 (N_8565,N_4046,N_2579);
xnor U8566 (N_8566,N_2038,N_4847);
and U8567 (N_8567,N_4118,N_3713);
and U8568 (N_8568,N_3571,N_2901);
or U8569 (N_8569,N_1805,N_3846);
nor U8570 (N_8570,N_292,N_1814);
nor U8571 (N_8571,N_3122,N_3229);
nor U8572 (N_8572,N_2945,N_3629);
and U8573 (N_8573,N_1592,N_2246);
xnor U8574 (N_8574,N_4294,N_942);
or U8575 (N_8575,N_2332,N_4920);
or U8576 (N_8576,N_2854,N_2538);
or U8577 (N_8577,N_1256,N_4722);
xor U8578 (N_8578,N_1446,N_2603);
or U8579 (N_8579,N_2577,N_3783);
nor U8580 (N_8580,N_4993,N_1974);
nor U8581 (N_8581,N_534,N_1941);
or U8582 (N_8582,N_4857,N_252);
or U8583 (N_8583,N_978,N_3077);
nor U8584 (N_8584,N_1014,N_1630);
or U8585 (N_8585,N_2459,N_4470);
and U8586 (N_8586,N_4022,N_3984);
nand U8587 (N_8587,N_4423,N_3227);
and U8588 (N_8588,N_4800,N_1184);
xor U8589 (N_8589,N_3222,N_4727);
and U8590 (N_8590,N_591,N_2156);
nand U8591 (N_8591,N_2977,N_837);
xnor U8592 (N_8592,N_2639,N_2454);
xor U8593 (N_8593,N_481,N_3391);
or U8594 (N_8594,N_1105,N_1900);
and U8595 (N_8595,N_1241,N_3158);
xor U8596 (N_8596,N_843,N_4065);
xnor U8597 (N_8597,N_3631,N_3934);
nand U8598 (N_8598,N_3091,N_4130);
nor U8599 (N_8599,N_563,N_2096);
or U8600 (N_8600,N_2554,N_4503);
xor U8601 (N_8601,N_3207,N_1452);
xor U8602 (N_8602,N_83,N_1094);
nor U8603 (N_8603,N_3856,N_1060);
xnor U8604 (N_8604,N_1057,N_3042);
nand U8605 (N_8605,N_1004,N_1739);
xnor U8606 (N_8606,N_4138,N_2397);
xor U8607 (N_8607,N_4941,N_3799);
nor U8608 (N_8608,N_2456,N_1850);
and U8609 (N_8609,N_4936,N_400);
nand U8610 (N_8610,N_2967,N_3407);
xor U8611 (N_8611,N_4568,N_2997);
xor U8612 (N_8612,N_2455,N_617);
xnor U8613 (N_8613,N_4651,N_665);
nor U8614 (N_8614,N_1530,N_2489);
or U8615 (N_8615,N_1794,N_1846);
nand U8616 (N_8616,N_4120,N_3509);
nor U8617 (N_8617,N_1447,N_2933);
nand U8618 (N_8618,N_2967,N_3975);
nand U8619 (N_8619,N_2380,N_3775);
xor U8620 (N_8620,N_1774,N_3257);
nand U8621 (N_8621,N_3305,N_1968);
and U8622 (N_8622,N_4334,N_4516);
and U8623 (N_8623,N_2198,N_3980);
or U8624 (N_8624,N_2340,N_701);
and U8625 (N_8625,N_3026,N_1213);
or U8626 (N_8626,N_1433,N_1264);
xnor U8627 (N_8627,N_533,N_3102);
or U8628 (N_8628,N_3632,N_2379);
nand U8629 (N_8629,N_3888,N_4881);
nand U8630 (N_8630,N_3519,N_2754);
nand U8631 (N_8631,N_391,N_1019);
xnor U8632 (N_8632,N_1144,N_2976);
nand U8633 (N_8633,N_1516,N_4064);
and U8634 (N_8634,N_1874,N_1747);
nor U8635 (N_8635,N_59,N_302);
nand U8636 (N_8636,N_2859,N_221);
nor U8637 (N_8637,N_1765,N_57);
nor U8638 (N_8638,N_2535,N_345);
and U8639 (N_8639,N_2946,N_365);
and U8640 (N_8640,N_2015,N_2975);
nor U8641 (N_8641,N_4259,N_4096);
and U8642 (N_8642,N_3527,N_3692);
nor U8643 (N_8643,N_299,N_583);
or U8644 (N_8644,N_2207,N_3267);
nor U8645 (N_8645,N_3006,N_2424);
and U8646 (N_8646,N_957,N_912);
or U8647 (N_8647,N_2433,N_2723);
nor U8648 (N_8648,N_224,N_3566);
nand U8649 (N_8649,N_315,N_762);
and U8650 (N_8650,N_837,N_3834);
xor U8651 (N_8651,N_924,N_4669);
and U8652 (N_8652,N_2755,N_4782);
xor U8653 (N_8653,N_980,N_1916);
and U8654 (N_8654,N_776,N_2191);
or U8655 (N_8655,N_1491,N_235);
nand U8656 (N_8656,N_1890,N_2331);
or U8657 (N_8657,N_1088,N_1278);
or U8658 (N_8658,N_3124,N_1028);
nand U8659 (N_8659,N_4208,N_322);
nand U8660 (N_8660,N_114,N_3841);
nor U8661 (N_8661,N_1155,N_2942);
or U8662 (N_8662,N_601,N_3096);
nand U8663 (N_8663,N_4804,N_3743);
xor U8664 (N_8664,N_4627,N_584);
or U8665 (N_8665,N_725,N_4662);
xnor U8666 (N_8666,N_3933,N_4401);
xnor U8667 (N_8667,N_2492,N_3839);
nand U8668 (N_8668,N_4007,N_1566);
and U8669 (N_8669,N_4875,N_3246);
nand U8670 (N_8670,N_3669,N_4998);
or U8671 (N_8671,N_4708,N_3546);
or U8672 (N_8672,N_1776,N_2407);
nor U8673 (N_8673,N_2605,N_2801);
or U8674 (N_8674,N_965,N_3605);
nor U8675 (N_8675,N_2404,N_944);
xor U8676 (N_8676,N_1683,N_98);
nand U8677 (N_8677,N_3451,N_2750);
nand U8678 (N_8678,N_2523,N_606);
and U8679 (N_8679,N_480,N_4674);
or U8680 (N_8680,N_23,N_4207);
nor U8681 (N_8681,N_878,N_4802);
nand U8682 (N_8682,N_3225,N_1636);
nor U8683 (N_8683,N_2344,N_542);
xnor U8684 (N_8684,N_1351,N_4355);
xor U8685 (N_8685,N_753,N_3271);
nand U8686 (N_8686,N_1288,N_729);
nor U8687 (N_8687,N_2586,N_3754);
nand U8688 (N_8688,N_4395,N_3929);
xnor U8689 (N_8689,N_3007,N_4816);
nand U8690 (N_8690,N_3226,N_933);
and U8691 (N_8691,N_4840,N_4079);
nor U8692 (N_8692,N_4602,N_1026);
nor U8693 (N_8693,N_3137,N_734);
or U8694 (N_8694,N_1256,N_3678);
nor U8695 (N_8695,N_911,N_3801);
or U8696 (N_8696,N_3093,N_2729);
or U8697 (N_8697,N_3355,N_758);
nand U8698 (N_8698,N_2417,N_4976);
nand U8699 (N_8699,N_4925,N_2079);
xor U8700 (N_8700,N_2506,N_4674);
and U8701 (N_8701,N_4321,N_2541);
nand U8702 (N_8702,N_4680,N_616);
xnor U8703 (N_8703,N_24,N_1001);
xnor U8704 (N_8704,N_446,N_3355);
nand U8705 (N_8705,N_696,N_4185);
nand U8706 (N_8706,N_2957,N_74);
xnor U8707 (N_8707,N_1718,N_199);
or U8708 (N_8708,N_130,N_3353);
nand U8709 (N_8709,N_3056,N_3258);
nand U8710 (N_8710,N_3101,N_4961);
xnor U8711 (N_8711,N_2047,N_2191);
and U8712 (N_8712,N_3793,N_2964);
or U8713 (N_8713,N_2859,N_4658);
and U8714 (N_8714,N_253,N_936);
and U8715 (N_8715,N_3458,N_3765);
xor U8716 (N_8716,N_1543,N_1298);
or U8717 (N_8717,N_1916,N_7);
and U8718 (N_8718,N_2025,N_3054);
or U8719 (N_8719,N_3608,N_3390);
nor U8720 (N_8720,N_4802,N_1578);
or U8721 (N_8721,N_301,N_503);
and U8722 (N_8722,N_4587,N_3886);
xor U8723 (N_8723,N_3130,N_1538);
xnor U8724 (N_8724,N_2537,N_2352);
nand U8725 (N_8725,N_4964,N_1717);
nor U8726 (N_8726,N_1987,N_1830);
xor U8727 (N_8727,N_4136,N_3387);
xnor U8728 (N_8728,N_2935,N_2127);
nand U8729 (N_8729,N_984,N_4620);
nand U8730 (N_8730,N_4828,N_1642);
nand U8731 (N_8731,N_3297,N_2595);
and U8732 (N_8732,N_4141,N_319);
nand U8733 (N_8733,N_941,N_1533);
xnor U8734 (N_8734,N_1561,N_2233);
or U8735 (N_8735,N_3630,N_2119);
and U8736 (N_8736,N_588,N_85);
or U8737 (N_8737,N_243,N_1028);
xor U8738 (N_8738,N_4194,N_1870);
nor U8739 (N_8739,N_59,N_782);
nand U8740 (N_8740,N_2122,N_3251);
xor U8741 (N_8741,N_1186,N_2127);
xnor U8742 (N_8742,N_1846,N_1602);
and U8743 (N_8743,N_1544,N_1014);
nand U8744 (N_8744,N_2697,N_4676);
or U8745 (N_8745,N_4870,N_4748);
xnor U8746 (N_8746,N_3052,N_3864);
or U8747 (N_8747,N_3400,N_1827);
or U8748 (N_8748,N_3324,N_609);
and U8749 (N_8749,N_4430,N_4983);
nand U8750 (N_8750,N_2765,N_1699);
or U8751 (N_8751,N_4044,N_1526);
and U8752 (N_8752,N_1803,N_2658);
nor U8753 (N_8753,N_4031,N_3166);
nand U8754 (N_8754,N_253,N_2377);
xnor U8755 (N_8755,N_3302,N_1613);
and U8756 (N_8756,N_3805,N_1612);
and U8757 (N_8757,N_1917,N_867);
nor U8758 (N_8758,N_1424,N_1071);
nand U8759 (N_8759,N_646,N_4963);
xnor U8760 (N_8760,N_4669,N_156);
nor U8761 (N_8761,N_2651,N_4771);
nor U8762 (N_8762,N_4912,N_1431);
xnor U8763 (N_8763,N_2867,N_1033);
or U8764 (N_8764,N_1820,N_4035);
xnor U8765 (N_8765,N_4090,N_2289);
xnor U8766 (N_8766,N_2822,N_1801);
or U8767 (N_8767,N_1893,N_4988);
nor U8768 (N_8768,N_4623,N_242);
or U8769 (N_8769,N_2071,N_1);
nand U8770 (N_8770,N_855,N_1369);
or U8771 (N_8771,N_4515,N_3904);
nor U8772 (N_8772,N_3424,N_4128);
xor U8773 (N_8773,N_1758,N_2599);
nor U8774 (N_8774,N_1563,N_3991);
nor U8775 (N_8775,N_4749,N_2580);
nor U8776 (N_8776,N_3762,N_3050);
and U8777 (N_8777,N_3585,N_3265);
or U8778 (N_8778,N_1377,N_1598);
xor U8779 (N_8779,N_3947,N_3073);
or U8780 (N_8780,N_1850,N_3622);
xnor U8781 (N_8781,N_4669,N_1352);
and U8782 (N_8782,N_4076,N_683);
nand U8783 (N_8783,N_4122,N_1773);
nand U8784 (N_8784,N_4920,N_2473);
nor U8785 (N_8785,N_2990,N_666);
and U8786 (N_8786,N_2171,N_4134);
and U8787 (N_8787,N_4736,N_4163);
xor U8788 (N_8788,N_4180,N_98);
xnor U8789 (N_8789,N_424,N_503);
nand U8790 (N_8790,N_1751,N_1112);
xnor U8791 (N_8791,N_504,N_588);
or U8792 (N_8792,N_281,N_1016);
nand U8793 (N_8793,N_3927,N_3726);
or U8794 (N_8794,N_388,N_1665);
xnor U8795 (N_8795,N_1963,N_871);
nand U8796 (N_8796,N_1068,N_1512);
or U8797 (N_8797,N_424,N_1610);
xor U8798 (N_8798,N_2967,N_3898);
nor U8799 (N_8799,N_125,N_3119);
nand U8800 (N_8800,N_4625,N_3923);
and U8801 (N_8801,N_2443,N_2276);
nor U8802 (N_8802,N_1672,N_1528);
xor U8803 (N_8803,N_4021,N_4636);
xnor U8804 (N_8804,N_2302,N_3119);
and U8805 (N_8805,N_3878,N_2548);
nand U8806 (N_8806,N_1980,N_4962);
xor U8807 (N_8807,N_4379,N_2644);
nor U8808 (N_8808,N_4558,N_2996);
or U8809 (N_8809,N_3291,N_1145);
and U8810 (N_8810,N_1483,N_4126);
nand U8811 (N_8811,N_1705,N_1870);
or U8812 (N_8812,N_2347,N_43);
xor U8813 (N_8813,N_4546,N_4017);
and U8814 (N_8814,N_294,N_2064);
nor U8815 (N_8815,N_879,N_3408);
xnor U8816 (N_8816,N_4349,N_1081);
nor U8817 (N_8817,N_720,N_3639);
or U8818 (N_8818,N_310,N_593);
or U8819 (N_8819,N_834,N_843);
nor U8820 (N_8820,N_4815,N_1797);
xor U8821 (N_8821,N_4508,N_4940);
or U8822 (N_8822,N_1635,N_3980);
nand U8823 (N_8823,N_1113,N_2755);
nand U8824 (N_8824,N_4968,N_2799);
xnor U8825 (N_8825,N_4059,N_1385);
nor U8826 (N_8826,N_3012,N_2108);
xnor U8827 (N_8827,N_1113,N_3563);
or U8828 (N_8828,N_3788,N_4791);
nand U8829 (N_8829,N_1115,N_1045);
nand U8830 (N_8830,N_464,N_1761);
nor U8831 (N_8831,N_1131,N_259);
nand U8832 (N_8832,N_436,N_211);
and U8833 (N_8833,N_675,N_1778);
nor U8834 (N_8834,N_4418,N_1229);
nor U8835 (N_8835,N_3113,N_237);
nand U8836 (N_8836,N_1421,N_1834);
nor U8837 (N_8837,N_59,N_4271);
nor U8838 (N_8838,N_1688,N_878);
nand U8839 (N_8839,N_2857,N_3425);
nor U8840 (N_8840,N_977,N_4986);
and U8841 (N_8841,N_4966,N_328);
nand U8842 (N_8842,N_4901,N_2442);
and U8843 (N_8843,N_693,N_207);
nor U8844 (N_8844,N_3050,N_1428);
nand U8845 (N_8845,N_2500,N_2255);
xor U8846 (N_8846,N_234,N_1043);
xnor U8847 (N_8847,N_3170,N_699);
nor U8848 (N_8848,N_3778,N_1283);
or U8849 (N_8849,N_4225,N_4616);
nand U8850 (N_8850,N_4148,N_435);
xor U8851 (N_8851,N_3974,N_2683);
nor U8852 (N_8852,N_346,N_4181);
or U8853 (N_8853,N_598,N_324);
nor U8854 (N_8854,N_1462,N_61);
and U8855 (N_8855,N_1658,N_2767);
and U8856 (N_8856,N_2160,N_1281);
and U8857 (N_8857,N_3157,N_4266);
or U8858 (N_8858,N_4702,N_3292);
and U8859 (N_8859,N_615,N_1497);
and U8860 (N_8860,N_3112,N_4543);
and U8861 (N_8861,N_2883,N_4900);
nand U8862 (N_8862,N_1590,N_4699);
or U8863 (N_8863,N_3389,N_2324);
and U8864 (N_8864,N_4263,N_429);
nand U8865 (N_8865,N_2425,N_1412);
xor U8866 (N_8866,N_4646,N_4495);
nor U8867 (N_8867,N_3671,N_1404);
or U8868 (N_8868,N_4948,N_4940);
nor U8869 (N_8869,N_4410,N_4983);
xor U8870 (N_8870,N_2329,N_3394);
or U8871 (N_8871,N_5,N_3883);
xnor U8872 (N_8872,N_838,N_4802);
xor U8873 (N_8873,N_4776,N_2393);
nand U8874 (N_8874,N_3614,N_4065);
nor U8875 (N_8875,N_1995,N_742);
xnor U8876 (N_8876,N_2249,N_464);
xor U8877 (N_8877,N_952,N_2531);
and U8878 (N_8878,N_35,N_4139);
xor U8879 (N_8879,N_877,N_459);
and U8880 (N_8880,N_4162,N_2953);
nor U8881 (N_8881,N_627,N_142);
or U8882 (N_8882,N_4971,N_1006);
nor U8883 (N_8883,N_1546,N_3495);
and U8884 (N_8884,N_341,N_4516);
nor U8885 (N_8885,N_4598,N_230);
xor U8886 (N_8886,N_4411,N_4380);
nand U8887 (N_8887,N_1810,N_570);
or U8888 (N_8888,N_3241,N_320);
nor U8889 (N_8889,N_990,N_2528);
xnor U8890 (N_8890,N_4427,N_2410);
and U8891 (N_8891,N_2978,N_3861);
and U8892 (N_8892,N_2934,N_788);
nor U8893 (N_8893,N_455,N_1386);
or U8894 (N_8894,N_4773,N_1576);
nor U8895 (N_8895,N_3153,N_2322);
and U8896 (N_8896,N_1282,N_104);
xnor U8897 (N_8897,N_4008,N_3024);
nor U8898 (N_8898,N_4033,N_3275);
nand U8899 (N_8899,N_1004,N_3173);
nor U8900 (N_8900,N_2446,N_4966);
nand U8901 (N_8901,N_1763,N_52);
nand U8902 (N_8902,N_3873,N_825);
nand U8903 (N_8903,N_2623,N_1122);
and U8904 (N_8904,N_1051,N_349);
nand U8905 (N_8905,N_3969,N_4015);
nor U8906 (N_8906,N_2136,N_1364);
nor U8907 (N_8907,N_1936,N_2531);
nand U8908 (N_8908,N_3784,N_3619);
and U8909 (N_8909,N_1739,N_1460);
xor U8910 (N_8910,N_3676,N_3900);
nor U8911 (N_8911,N_849,N_4834);
or U8912 (N_8912,N_2745,N_1839);
nor U8913 (N_8913,N_2350,N_2599);
xnor U8914 (N_8914,N_912,N_4251);
and U8915 (N_8915,N_1260,N_1181);
nor U8916 (N_8916,N_4376,N_1539);
nand U8917 (N_8917,N_1419,N_3545);
or U8918 (N_8918,N_4149,N_123);
and U8919 (N_8919,N_4169,N_3010);
nor U8920 (N_8920,N_1936,N_1705);
or U8921 (N_8921,N_1365,N_3129);
xnor U8922 (N_8922,N_1417,N_2569);
nand U8923 (N_8923,N_2466,N_3608);
xnor U8924 (N_8924,N_3535,N_807);
or U8925 (N_8925,N_4159,N_4657);
and U8926 (N_8926,N_4256,N_2982);
or U8927 (N_8927,N_1837,N_1954);
xnor U8928 (N_8928,N_810,N_3271);
xor U8929 (N_8929,N_2461,N_126);
xnor U8930 (N_8930,N_986,N_2263);
xnor U8931 (N_8931,N_4975,N_200);
xor U8932 (N_8932,N_225,N_3398);
xnor U8933 (N_8933,N_2692,N_3998);
xnor U8934 (N_8934,N_4054,N_1136);
nand U8935 (N_8935,N_1577,N_2825);
and U8936 (N_8936,N_1239,N_2602);
or U8937 (N_8937,N_2260,N_2203);
or U8938 (N_8938,N_1058,N_3220);
nand U8939 (N_8939,N_3486,N_4220);
xor U8940 (N_8940,N_3805,N_3736);
or U8941 (N_8941,N_3914,N_4487);
nand U8942 (N_8942,N_3828,N_4436);
nand U8943 (N_8943,N_3374,N_4091);
or U8944 (N_8944,N_3727,N_1905);
or U8945 (N_8945,N_2870,N_3582);
xor U8946 (N_8946,N_3075,N_1593);
xnor U8947 (N_8947,N_4974,N_3074);
and U8948 (N_8948,N_666,N_3060);
and U8949 (N_8949,N_554,N_198);
nand U8950 (N_8950,N_448,N_3511);
nand U8951 (N_8951,N_272,N_1956);
xor U8952 (N_8952,N_3826,N_3891);
nand U8953 (N_8953,N_2456,N_1661);
and U8954 (N_8954,N_325,N_3409);
nand U8955 (N_8955,N_4462,N_4064);
and U8956 (N_8956,N_1720,N_373);
xnor U8957 (N_8957,N_4192,N_1486);
and U8958 (N_8958,N_1579,N_1298);
and U8959 (N_8959,N_4885,N_2888);
and U8960 (N_8960,N_4093,N_4811);
or U8961 (N_8961,N_4570,N_3972);
or U8962 (N_8962,N_2344,N_791);
and U8963 (N_8963,N_4102,N_3654);
nor U8964 (N_8964,N_1433,N_3418);
nand U8965 (N_8965,N_3753,N_2244);
xor U8966 (N_8966,N_772,N_4775);
and U8967 (N_8967,N_920,N_707);
nand U8968 (N_8968,N_1261,N_136);
nor U8969 (N_8969,N_2646,N_2199);
nor U8970 (N_8970,N_4703,N_4126);
and U8971 (N_8971,N_1745,N_2037);
and U8972 (N_8972,N_3758,N_625);
xnor U8973 (N_8973,N_3701,N_3531);
and U8974 (N_8974,N_1296,N_2876);
nand U8975 (N_8975,N_2564,N_1006);
xnor U8976 (N_8976,N_1974,N_122);
xor U8977 (N_8977,N_1441,N_3556);
nor U8978 (N_8978,N_4288,N_4521);
and U8979 (N_8979,N_3145,N_4);
nand U8980 (N_8980,N_2605,N_4314);
or U8981 (N_8981,N_1051,N_1691);
or U8982 (N_8982,N_1484,N_4774);
xnor U8983 (N_8983,N_4090,N_1614);
xnor U8984 (N_8984,N_3618,N_122);
and U8985 (N_8985,N_38,N_3247);
nand U8986 (N_8986,N_2331,N_2801);
and U8987 (N_8987,N_4616,N_4018);
or U8988 (N_8988,N_4451,N_1426);
xor U8989 (N_8989,N_849,N_873);
nand U8990 (N_8990,N_1154,N_576);
nor U8991 (N_8991,N_3117,N_1237);
nor U8992 (N_8992,N_873,N_2090);
or U8993 (N_8993,N_2449,N_1681);
nand U8994 (N_8994,N_1136,N_3635);
and U8995 (N_8995,N_2552,N_3909);
xor U8996 (N_8996,N_1407,N_2589);
or U8997 (N_8997,N_3765,N_924);
or U8998 (N_8998,N_4550,N_215);
or U8999 (N_8999,N_10,N_1277);
xor U9000 (N_9000,N_235,N_391);
or U9001 (N_9001,N_2822,N_2387);
or U9002 (N_9002,N_2141,N_2372);
xnor U9003 (N_9003,N_1600,N_1070);
xnor U9004 (N_9004,N_1636,N_3295);
nor U9005 (N_9005,N_3452,N_4072);
and U9006 (N_9006,N_3468,N_209);
and U9007 (N_9007,N_1467,N_4603);
nand U9008 (N_9008,N_1543,N_3031);
or U9009 (N_9009,N_773,N_397);
and U9010 (N_9010,N_3801,N_4033);
nand U9011 (N_9011,N_1447,N_2889);
and U9012 (N_9012,N_2960,N_4011);
nor U9013 (N_9013,N_4718,N_2472);
xor U9014 (N_9014,N_862,N_353);
nand U9015 (N_9015,N_4556,N_3623);
xor U9016 (N_9016,N_2620,N_825);
nand U9017 (N_9017,N_83,N_2291);
and U9018 (N_9018,N_3954,N_4518);
and U9019 (N_9019,N_3016,N_2931);
or U9020 (N_9020,N_139,N_612);
xnor U9021 (N_9021,N_3259,N_1830);
xnor U9022 (N_9022,N_2898,N_4008);
nor U9023 (N_9023,N_170,N_596);
nor U9024 (N_9024,N_2809,N_1638);
xor U9025 (N_9025,N_216,N_234);
nor U9026 (N_9026,N_3163,N_3958);
and U9027 (N_9027,N_1132,N_235);
nor U9028 (N_9028,N_4763,N_3868);
nand U9029 (N_9029,N_390,N_1277);
xnor U9030 (N_9030,N_222,N_2937);
xor U9031 (N_9031,N_308,N_4901);
nand U9032 (N_9032,N_2381,N_3025);
nor U9033 (N_9033,N_4694,N_3304);
and U9034 (N_9034,N_4602,N_2136);
or U9035 (N_9035,N_4258,N_3721);
and U9036 (N_9036,N_4211,N_4555);
nor U9037 (N_9037,N_1954,N_3503);
nand U9038 (N_9038,N_1694,N_3480);
nand U9039 (N_9039,N_2036,N_359);
xnor U9040 (N_9040,N_912,N_3670);
or U9041 (N_9041,N_138,N_2711);
or U9042 (N_9042,N_3441,N_63);
nor U9043 (N_9043,N_1817,N_1252);
nor U9044 (N_9044,N_4543,N_3311);
nand U9045 (N_9045,N_738,N_114);
nor U9046 (N_9046,N_233,N_845);
nand U9047 (N_9047,N_217,N_733);
nand U9048 (N_9048,N_2462,N_3315);
xnor U9049 (N_9049,N_4604,N_2540);
and U9050 (N_9050,N_4440,N_3874);
xor U9051 (N_9051,N_2202,N_2901);
nand U9052 (N_9052,N_4566,N_1756);
xor U9053 (N_9053,N_4098,N_2518);
xor U9054 (N_9054,N_3318,N_1713);
xor U9055 (N_9055,N_2853,N_2835);
or U9056 (N_9056,N_4856,N_4524);
nor U9057 (N_9057,N_2579,N_3884);
or U9058 (N_9058,N_3449,N_440);
or U9059 (N_9059,N_2732,N_1402);
nor U9060 (N_9060,N_1266,N_4209);
nand U9061 (N_9061,N_4250,N_4612);
nand U9062 (N_9062,N_494,N_4885);
nand U9063 (N_9063,N_26,N_3515);
or U9064 (N_9064,N_1380,N_701);
xor U9065 (N_9065,N_59,N_839);
nor U9066 (N_9066,N_3239,N_91);
or U9067 (N_9067,N_3441,N_627);
nor U9068 (N_9068,N_4629,N_4295);
nand U9069 (N_9069,N_3437,N_3582);
nand U9070 (N_9070,N_4938,N_4157);
xor U9071 (N_9071,N_2328,N_3927);
xnor U9072 (N_9072,N_400,N_4253);
or U9073 (N_9073,N_368,N_964);
nand U9074 (N_9074,N_4205,N_2376);
nand U9075 (N_9075,N_2083,N_3936);
nor U9076 (N_9076,N_547,N_221);
and U9077 (N_9077,N_687,N_4555);
or U9078 (N_9078,N_135,N_1063);
and U9079 (N_9079,N_1858,N_4546);
nor U9080 (N_9080,N_3020,N_2769);
xnor U9081 (N_9081,N_1708,N_2010);
or U9082 (N_9082,N_4046,N_288);
nor U9083 (N_9083,N_4570,N_682);
or U9084 (N_9084,N_3610,N_2239);
xor U9085 (N_9085,N_3722,N_1390);
nand U9086 (N_9086,N_2950,N_2035);
and U9087 (N_9087,N_4902,N_3453);
xor U9088 (N_9088,N_4559,N_3461);
and U9089 (N_9089,N_4701,N_1994);
nand U9090 (N_9090,N_4714,N_4211);
or U9091 (N_9091,N_1986,N_4444);
xnor U9092 (N_9092,N_2384,N_2925);
or U9093 (N_9093,N_1012,N_4094);
or U9094 (N_9094,N_3218,N_637);
or U9095 (N_9095,N_3029,N_4393);
and U9096 (N_9096,N_157,N_3475);
nand U9097 (N_9097,N_1431,N_4686);
and U9098 (N_9098,N_302,N_2404);
and U9099 (N_9099,N_3247,N_2090);
and U9100 (N_9100,N_4187,N_3376);
and U9101 (N_9101,N_123,N_4163);
xor U9102 (N_9102,N_4387,N_2109);
or U9103 (N_9103,N_3288,N_4067);
and U9104 (N_9104,N_4861,N_2637);
and U9105 (N_9105,N_4467,N_4574);
and U9106 (N_9106,N_2768,N_3494);
and U9107 (N_9107,N_4421,N_2121);
nand U9108 (N_9108,N_4776,N_1417);
xnor U9109 (N_9109,N_1501,N_58);
nor U9110 (N_9110,N_1832,N_4056);
nor U9111 (N_9111,N_1205,N_4425);
nand U9112 (N_9112,N_1216,N_4048);
and U9113 (N_9113,N_4263,N_3952);
nor U9114 (N_9114,N_1587,N_4678);
xnor U9115 (N_9115,N_3725,N_3636);
and U9116 (N_9116,N_4812,N_946);
nand U9117 (N_9117,N_887,N_1235);
or U9118 (N_9118,N_3275,N_3396);
or U9119 (N_9119,N_4367,N_3097);
nand U9120 (N_9120,N_1430,N_97);
nor U9121 (N_9121,N_4939,N_2264);
nand U9122 (N_9122,N_4002,N_2267);
or U9123 (N_9123,N_89,N_224);
or U9124 (N_9124,N_1445,N_3250);
xnor U9125 (N_9125,N_4932,N_349);
or U9126 (N_9126,N_463,N_1375);
xor U9127 (N_9127,N_3926,N_4491);
or U9128 (N_9128,N_4710,N_3601);
xor U9129 (N_9129,N_150,N_4763);
xor U9130 (N_9130,N_1657,N_225);
xnor U9131 (N_9131,N_408,N_1334);
and U9132 (N_9132,N_591,N_4440);
or U9133 (N_9133,N_4427,N_2278);
nor U9134 (N_9134,N_1602,N_1042);
xor U9135 (N_9135,N_440,N_2803);
nand U9136 (N_9136,N_18,N_3300);
nand U9137 (N_9137,N_3904,N_3731);
and U9138 (N_9138,N_155,N_2667);
or U9139 (N_9139,N_3357,N_1390);
and U9140 (N_9140,N_280,N_65);
and U9141 (N_9141,N_2936,N_381);
nor U9142 (N_9142,N_2783,N_2527);
nand U9143 (N_9143,N_2055,N_1641);
and U9144 (N_9144,N_1343,N_4603);
or U9145 (N_9145,N_1235,N_274);
nor U9146 (N_9146,N_3094,N_3226);
nand U9147 (N_9147,N_3282,N_625);
and U9148 (N_9148,N_4387,N_1938);
xnor U9149 (N_9149,N_2058,N_2138);
and U9150 (N_9150,N_1448,N_4368);
nor U9151 (N_9151,N_4776,N_1065);
or U9152 (N_9152,N_3358,N_2045);
or U9153 (N_9153,N_4293,N_4868);
and U9154 (N_9154,N_3494,N_3639);
and U9155 (N_9155,N_3139,N_3677);
nor U9156 (N_9156,N_1306,N_801);
nand U9157 (N_9157,N_1189,N_3986);
xor U9158 (N_9158,N_2559,N_3794);
and U9159 (N_9159,N_4096,N_361);
and U9160 (N_9160,N_2065,N_1884);
and U9161 (N_9161,N_230,N_4080);
nor U9162 (N_9162,N_2009,N_2250);
or U9163 (N_9163,N_1180,N_21);
nand U9164 (N_9164,N_838,N_2270);
nand U9165 (N_9165,N_3566,N_1976);
nand U9166 (N_9166,N_37,N_4356);
nand U9167 (N_9167,N_4456,N_1818);
nor U9168 (N_9168,N_2796,N_4347);
nor U9169 (N_9169,N_337,N_4635);
xnor U9170 (N_9170,N_1233,N_4926);
or U9171 (N_9171,N_4124,N_4765);
or U9172 (N_9172,N_3258,N_1892);
nor U9173 (N_9173,N_1079,N_1996);
xor U9174 (N_9174,N_2274,N_4711);
or U9175 (N_9175,N_347,N_1694);
xnor U9176 (N_9176,N_4556,N_3193);
nor U9177 (N_9177,N_733,N_4770);
xnor U9178 (N_9178,N_1676,N_4400);
nand U9179 (N_9179,N_3331,N_583);
nor U9180 (N_9180,N_409,N_2398);
or U9181 (N_9181,N_3258,N_1441);
xor U9182 (N_9182,N_2929,N_115);
and U9183 (N_9183,N_919,N_516);
xnor U9184 (N_9184,N_4920,N_2231);
nor U9185 (N_9185,N_319,N_1311);
and U9186 (N_9186,N_85,N_788);
and U9187 (N_9187,N_4370,N_4235);
and U9188 (N_9188,N_3756,N_4642);
xnor U9189 (N_9189,N_915,N_4593);
and U9190 (N_9190,N_3584,N_610);
xnor U9191 (N_9191,N_2785,N_913);
and U9192 (N_9192,N_4792,N_1939);
nand U9193 (N_9193,N_2709,N_668);
nand U9194 (N_9194,N_2052,N_169);
xnor U9195 (N_9195,N_3308,N_4791);
and U9196 (N_9196,N_921,N_135);
nor U9197 (N_9197,N_1226,N_331);
nand U9198 (N_9198,N_3648,N_4116);
or U9199 (N_9199,N_2545,N_2962);
nand U9200 (N_9200,N_1556,N_2982);
xnor U9201 (N_9201,N_2638,N_4219);
nor U9202 (N_9202,N_3944,N_1618);
and U9203 (N_9203,N_3425,N_3646);
nor U9204 (N_9204,N_2512,N_3939);
or U9205 (N_9205,N_1818,N_4195);
or U9206 (N_9206,N_1186,N_4896);
xnor U9207 (N_9207,N_982,N_4002);
nor U9208 (N_9208,N_906,N_903);
nor U9209 (N_9209,N_4751,N_2209);
nor U9210 (N_9210,N_2575,N_524);
nand U9211 (N_9211,N_4649,N_534);
or U9212 (N_9212,N_3049,N_3327);
nand U9213 (N_9213,N_756,N_2145);
xnor U9214 (N_9214,N_106,N_2366);
nor U9215 (N_9215,N_4021,N_2080);
nand U9216 (N_9216,N_2419,N_3944);
xnor U9217 (N_9217,N_628,N_2917);
and U9218 (N_9218,N_528,N_1552);
nand U9219 (N_9219,N_3811,N_3628);
xor U9220 (N_9220,N_2178,N_2546);
nor U9221 (N_9221,N_3659,N_2027);
nor U9222 (N_9222,N_1988,N_772);
xnor U9223 (N_9223,N_3371,N_2075);
and U9224 (N_9224,N_1978,N_1816);
xnor U9225 (N_9225,N_259,N_1704);
or U9226 (N_9226,N_449,N_2258);
nand U9227 (N_9227,N_1315,N_4571);
nand U9228 (N_9228,N_1339,N_4530);
nor U9229 (N_9229,N_2929,N_3017);
nand U9230 (N_9230,N_3146,N_2593);
or U9231 (N_9231,N_2444,N_2060);
or U9232 (N_9232,N_2756,N_1098);
and U9233 (N_9233,N_1293,N_2503);
nor U9234 (N_9234,N_3751,N_4771);
or U9235 (N_9235,N_621,N_1039);
xnor U9236 (N_9236,N_3164,N_11);
nand U9237 (N_9237,N_3117,N_476);
xnor U9238 (N_9238,N_417,N_1597);
nor U9239 (N_9239,N_4741,N_1502);
and U9240 (N_9240,N_2400,N_2280);
nor U9241 (N_9241,N_65,N_1971);
xor U9242 (N_9242,N_1070,N_334);
and U9243 (N_9243,N_1110,N_4981);
nor U9244 (N_9244,N_578,N_1097);
nor U9245 (N_9245,N_772,N_2746);
nand U9246 (N_9246,N_2905,N_895);
nor U9247 (N_9247,N_750,N_4058);
and U9248 (N_9248,N_4949,N_4150);
xor U9249 (N_9249,N_4597,N_832);
nor U9250 (N_9250,N_3176,N_4832);
nor U9251 (N_9251,N_2418,N_3357);
or U9252 (N_9252,N_2354,N_389);
or U9253 (N_9253,N_864,N_2057);
nor U9254 (N_9254,N_3919,N_1786);
xnor U9255 (N_9255,N_105,N_1112);
xor U9256 (N_9256,N_4459,N_1907);
and U9257 (N_9257,N_2153,N_3460);
xor U9258 (N_9258,N_1540,N_2404);
and U9259 (N_9259,N_4341,N_1911);
and U9260 (N_9260,N_1073,N_1492);
nand U9261 (N_9261,N_4899,N_1792);
or U9262 (N_9262,N_4671,N_2956);
nor U9263 (N_9263,N_4087,N_4661);
xor U9264 (N_9264,N_3401,N_3025);
nand U9265 (N_9265,N_515,N_2140);
or U9266 (N_9266,N_682,N_150);
or U9267 (N_9267,N_1994,N_979);
nor U9268 (N_9268,N_1621,N_2771);
or U9269 (N_9269,N_3601,N_4445);
and U9270 (N_9270,N_2990,N_3029);
or U9271 (N_9271,N_1468,N_4985);
nor U9272 (N_9272,N_1797,N_4498);
or U9273 (N_9273,N_3952,N_4192);
xnor U9274 (N_9274,N_3524,N_443);
nor U9275 (N_9275,N_2963,N_2221);
or U9276 (N_9276,N_3479,N_189);
and U9277 (N_9277,N_4237,N_4993);
nand U9278 (N_9278,N_3677,N_981);
or U9279 (N_9279,N_2357,N_3870);
nand U9280 (N_9280,N_889,N_2009);
and U9281 (N_9281,N_4565,N_2440);
or U9282 (N_9282,N_272,N_1835);
or U9283 (N_9283,N_513,N_173);
nor U9284 (N_9284,N_4593,N_3315);
and U9285 (N_9285,N_2816,N_3357);
nor U9286 (N_9286,N_481,N_4705);
or U9287 (N_9287,N_245,N_3523);
nor U9288 (N_9288,N_3556,N_366);
nand U9289 (N_9289,N_2002,N_4200);
or U9290 (N_9290,N_1760,N_4742);
xnor U9291 (N_9291,N_1080,N_3633);
nand U9292 (N_9292,N_2482,N_1841);
and U9293 (N_9293,N_4598,N_4309);
nand U9294 (N_9294,N_1024,N_1569);
xnor U9295 (N_9295,N_3919,N_2290);
or U9296 (N_9296,N_682,N_2915);
nor U9297 (N_9297,N_4687,N_1286);
nor U9298 (N_9298,N_1188,N_3904);
and U9299 (N_9299,N_1069,N_2615);
nand U9300 (N_9300,N_3956,N_3492);
nor U9301 (N_9301,N_1203,N_175);
and U9302 (N_9302,N_2952,N_3086);
and U9303 (N_9303,N_4328,N_2587);
and U9304 (N_9304,N_2875,N_1072);
nand U9305 (N_9305,N_4665,N_4210);
nand U9306 (N_9306,N_1955,N_2112);
xnor U9307 (N_9307,N_1544,N_2462);
nand U9308 (N_9308,N_114,N_532);
nand U9309 (N_9309,N_4601,N_791);
nor U9310 (N_9310,N_4731,N_249);
nor U9311 (N_9311,N_1271,N_269);
nor U9312 (N_9312,N_1919,N_3836);
nor U9313 (N_9313,N_1236,N_3217);
nand U9314 (N_9314,N_1988,N_2582);
and U9315 (N_9315,N_1602,N_1704);
xnor U9316 (N_9316,N_57,N_762);
and U9317 (N_9317,N_3019,N_2761);
nand U9318 (N_9318,N_4,N_3812);
and U9319 (N_9319,N_2696,N_383);
or U9320 (N_9320,N_1185,N_4899);
and U9321 (N_9321,N_2672,N_1499);
nor U9322 (N_9322,N_799,N_3516);
or U9323 (N_9323,N_1616,N_506);
and U9324 (N_9324,N_2116,N_1584);
and U9325 (N_9325,N_1402,N_433);
or U9326 (N_9326,N_2546,N_4821);
or U9327 (N_9327,N_1076,N_2736);
or U9328 (N_9328,N_3570,N_3967);
or U9329 (N_9329,N_851,N_2610);
and U9330 (N_9330,N_4706,N_3835);
nor U9331 (N_9331,N_772,N_2871);
or U9332 (N_9332,N_4800,N_1804);
and U9333 (N_9333,N_566,N_515);
nor U9334 (N_9334,N_120,N_2840);
or U9335 (N_9335,N_3908,N_393);
and U9336 (N_9336,N_854,N_1517);
nor U9337 (N_9337,N_545,N_801);
nor U9338 (N_9338,N_3858,N_1702);
xnor U9339 (N_9339,N_3690,N_2499);
nand U9340 (N_9340,N_2715,N_4479);
nand U9341 (N_9341,N_1548,N_3842);
or U9342 (N_9342,N_1595,N_3204);
or U9343 (N_9343,N_2521,N_2364);
nor U9344 (N_9344,N_2605,N_3777);
or U9345 (N_9345,N_2629,N_4313);
and U9346 (N_9346,N_2272,N_921);
and U9347 (N_9347,N_200,N_2107);
and U9348 (N_9348,N_2459,N_2245);
and U9349 (N_9349,N_2094,N_2062);
or U9350 (N_9350,N_3814,N_4498);
nand U9351 (N_9351,N_60,N_1143);
and U9352 (N_9352,N_3586,N_1750);
xor U9353 (N_9353,N_4444,N_2961);
and U9354 (N_9354,N_4102,N_3027);
nor U9355 (N_9355,N_3767,N_3952);
nand U9356 (N_9356,N_170,N_3529);
nor U9357 (N_9357,N_4563,N_4054);
nor U9358 (N_9358,N_1014,N_4996);
nor U9359 (N_9359,N_3004,N_3588);
nand U9360 (N_9360,N_2841,N_2244);
or U9361 (N_9361,N_4002,N_1847);
nor U9362 (N_9362,N_4673,N_3423);
nand U9363 (N_9363,N_2225,N_1786);
or U9364 (N_9364,N_1254,N_4427);
or U9365 (N_9365,N_3835,N_3834);
nor U9366 (N_9366,N_3672,N_3077);
nor U9367 (N_9367,N_979,N_3255);
nor U9368 (N_9368,N_4755,N_4992);
xnor U9369 (N_9369,N_4889,N_4560);
xnor U9370 (N_9370,N_1091,N_3657);
xnor U9371 (N_9371,N_1203,N_36);
or U9372 (N_9372,N_4213,N_546);
and U9373 (N_9373,N_3494,N_3273);
and U9374 (N_9374,N_2467,N_4022);
nor U9375 (N_9375,N_1183,N_851);
or U9376 (N_9376,N_4487,N_3290);
nor U9377 (N_9377,N_307,N_1958);
nand U9378 (N_9378,N_481,N_3600);
and U9379 (N_9379,N_3594,N_4362);
or U9380 (N_9380,N_946,N_2079);
nand U9381 (N_9381,N_2228,N_3532);
or U9382 (N_9382,N_193,N_3671);
and U9383 (N_9383,N_672,N_1844);
xnor U9384 (N_9384,N_4465,N_1565);
nor U9385 (N_9385,N_3131,N_4234);
nand U9386 (N_9386,N_214,N_3197);
xor U9387 (N_9387,N_974,N_4588);
nor U9388 (N_9388,N_4474,N_2038);
nand U9389 (N_9389,N_2635,N_2507);
or U9390 (N_9390,N_3298,N_410);
xnor U9391 (N_9391,N_650,N_210);
xor U9392 (N_9392,N_4390,N_1158);
nand U9393 (N_9393,N_679,N_4686);
nor U9394 (N_9394,N_2783,N_2704);
and U9395 (N_9395,N_2810,N_1812);
nand U9396 (N_9396,N_3120,N_1457);
xor U9397 (N_9397,N_898,N_256);
and U9398 (N_9398,N_3922,N_1787);
xnor U9399 (N_9399,N_957,N_3363);
xnor U9400 (N_9400,N_3094,N_4713);
nor U9401 (N_9401,N_307,N_4401);
nor U9402 (N_9402,N_3885,N_1003);
nor U9403 (N_9403,N_2804,N_4616);
nor U9404 (N_9404,N_4628,N_4947);
nor U9405 (N_9405,N_995,N_2185);
nand U9406 (N_9406,N_1767,N_1009);
and U9407 (N_9407,N_3986,N_4309);
and U9408 (N_9408,N_447,N_2203);
and U9409 (N_9409,N_293,N_3237);
nand U9410 (N_9410,N_4394,N_3565);
nand U9411 (N_9411,N_4448,N_819);
xor U9412 (N_9412,N_3866,N_1833);
and U9413 (N_9413,N_4758,N_886);
or U9414 (N_9414,N_2107,N_223);
and U9415 (N_9415,N_2229,N_334);
and U9416 (N_9416,N_3386,N_761);
and U9417 (N_9417,N_4783,N_2919);
or U9418 (N_9418,N_2707,N_1857);
or U9419 (N_9419,N_2586,N_2108);
or U9420 (N_9420,N_2400,N_4301);
nand U9421 (N_9421,N_2372,N_3502);
nand U9422 (N_9422,N_333,N_4907);
xor U9423 (N_9423,N_2360,N_4585);
xnor U9424 (N_9424,N_3815,N_3534);
xnor U9425 (N_9425,N_3601,N_491);
or U9426 (N_9426,N_4587,N_2986);
nand U9427 (N_9427,N_280,N_1064);
nor U9428 (N_9428,N_4515,N_2292);
xnor U9429 (N_9429,N_1882,N_881);
xnor U9430 (N_9430,N_2589,N_1006);
and U9431 (N_9431,N_3891,N_106);
xnor U9432 (N_9432,N_1610,N_3423);
or U9433 (N_9433,N_3594,N_2293);
or U9434 (N_9434,N_942,N_553);
nor U9435 (N_9435,N_1915,N_4089);
xnor U9436 (N_9436,N_153,N_472);
nor U9437 (N_9437,N_2803,N_4600);
nand U9438 (N_9438,N_1282,N_3676);
nor U9439 (N_9439,N_77,N_269);
xor U9440 (N_9440,N_491,N_1212);
or U9441 (N_9441,N_3363,N_1297);
or U9442 (N_9442,N_2301,N_1766);
nor U9443 (N_9443,N_1582,N_567);
nand U9444 (N_9444,N_4808,N_3739);
nor U9445 (N_9445,N_36,N_2591);
or U9446 (N_9446,N_4925,N_1017);
nand U9447 (N_9447,N_1555,N_3211);
xnor U9448 (N_9448,N_3581,N_4322);
xor U9449 (N_9449,N_4580,N_4051);
nand U9450 (N_9450,N_2706,N_2689);
or U9451 (N_9451,N_2720,N_3165);
or U9452 (N_9452,N_386,N_4677);
xnor U9453 (N_9453,N_2350,N_1843);
or U9454 (N_9454,N_3268,N_3697);
or U9455 (N_9455,N_336,N_4504);
and U9456 (N_9456,N_3838,N_250);
xnor U9457 (N_9457,N_487,N_3095);
and U9458 (N_9458,N_1266,N_3405);
and U9459 (N_9459,N_2383,N_3720);
nand U9460 (N_9460,N_1840,N_4362);
nand U9461 (N_9461,N_2939,N_4332);
or U9462 (N_9462,N_2996,N_2506);
nor U9463 (N_9463,N_2223,N_1352);
nor U9464 (N_9464,N_769,N_3569);
nor U9465 (N_9465,N_844,N_4071);
nand U9466 (N_9466,N_3252,N_906);
and U9467 (N_9467,N_2681,N_3117);
and U9468 (N_9468,N_3816,N_167);
nand U9469 (N_9469,N_922,N_3150);
xor U9470 (N_9470,N_256,N_4477);
nand U9471 (N_9471,N_3995,N_732);
xnor U9472 (N_9472,N_2352,N_3850);
nor U9473 (N_9473,N_153,N_4667);
nor U9474 (N_9474,N_1764,N_3026);
or U9475 (N_9475,N_262,N_1294);
or U9476 (N_9476,N_981,N_3432);
xor U9477 (N_9477,N_1809,N_1438);
and U9478 (N_9478,N_2026,N_22);
nand U9479 (N_9479,N_2123,N_1070);
xnor U9480 (N_9480,N_2799,N_1821);
nand U9481 (N_9481,N_2497,N_4853);
nor U9482 (N_9482,N_2725,N_1534);
or U9483 (N_9483,N_2412,N_252);
nor U9484 (N_9484,N_752,N_4112);
nand U9485 (N_9485,N_2543,N_4808);
nand U9486 (N_9486,N_4963,N_4841);
or U9487 (N_9487,N_3337,N_4404);
nand U9488 (N_9488,N_1186,N_520);
nor U9489 (N_9489,N_1615,N_3454);
and U9490 (N_9490,N_1458,N_4467);
nor U9491 (N_9491,N_1678,N_3296);
nand U9492 (N_9492,N_2739,N_3043);
or U9493 (N_9493,N_3542,N_4490);
and U9494 (N_9494,N_3415,N_3543);
and U9495 (N_9495,N_254,N_1237);
and U9496 (N_9496,N_2137,N_652);
or U9497 (N_9497,N_3856,N_4960);
xnor U9498 (N_9498,N_3313,N_2793);
and U9499 (N_9499,N_3414,N_3804);
and U9500 (N_9500,N_3344,N_479);
nor U9501 (N_9501,N_2095,N_3242);
nor U9502 (N_9502,N_2259,N_2681);
and U9503 (N_9503,N_3454,N_376);
nand U9504 (N_9504,N_1635,N_2889);
or U9505 (N_9505,N_311,N_2818);
nor U9506 (N_9506,N_2778,N_4897);
and U9507 (N_9507,N_3860,N_630);
xnor U9508 (N_9508,N_2019,N_4576);
nor U9509 (N_9509,N_3487,N_315);
nand U9510 (N_9510,N_4364,N_2996);
xnor U9511 (N_9511,N_2109,N_2133);
and U9512 (N_9512,N_3044,N_4621);
or U9513 (N_9513,N_351,N_993);
or U9514 (N_9514,N_2478,N_1963);
or U9515 (N_9515,N_3871,N_1401);
nor U9516 (N_9516,N_4784,N_720);
nor U9517 (N_9517,N_2530,N_3679);
xor U9518 (N_9518,N_3330,N_4918);
nand U9519 (N_9519,N_1026,N_2923);
nand U9520 (N_9520,N_1253,N_377);
nand U9521 (N_9521,N_4162,N_917);
nand U9522 (N_9522,N_2005,N_2079);
and U9523 (N_9523,N_4349,N_3203);
nand U9524 (N_9524,N_4674,N_2291);
xor U9525 (N_9525,N_1219,N_3017);
nand U9526 (N_9526,N_1558,N_1648);
nor U9527 (N_9527,N_4600,N_4984);
nand U9528 (N_9528,N_4599,N_3590);
xor U9529 (N_9529,N_2594,N_3521);
and U9530 (N_9530,N_4589,N_4075);
nor U9531 (N_9531,N_342,N_2345);
or U9532 (N_9532,N_3969,N_3942);
nor U9533 (N_9533,N_3161,N_2531);
nand U9534 (N_9534,N_975,N_591);
nor U9535 (N_9535,N_4938,N_4676);
nand U9536 (N_9536,N_2103,N_439);
xor U9537 (N_9537,N_1378,N_862);
or U9538 (N_9538,N_4134,N_4270);
and U9539 (N_9539,N_3382,N_3106);
or U9540 (N_9540,N_34,N_2285);
nand U9541 (N_9541,N_4565,N_409);
nand U9542 (N_9542,N_3977,N_1493);
nand U9543 (N_9543,N_516,N_61);
or U9544 (N_9544,N_1991,N_3908);
nand U9545 (N_9545,N_2203,N_2102);
nor U9546 (N_9546,N_4887,N_4306);
nand U9547 (N_9547,N_3987,N_3592);
and U9548 (N_9548,N_4695,N_4563);
and U9549 (N_9549,N_473,N_3450);
nor U9550 (N_9550,N_4447,N_106);
nand U9551 (N_9551,N_262,N_576);
nor U9552 (N_9552,N_2385,N_2906);
nand U9553 (N_9553,N_17,N_472);
xnor U9554 (N_9554,N_4459,N_3926);
xnor U9555 (N_9555,N_4918,N_4516);
xnor U9556 (N_9556,N_4622,N_3510);
xor U9557 (N_9557,N_4685,N_4055);
xnor U9558 (N_9558,N_1631,N_2561);
nor U9559 (N_9559,N_4468,N_3982);
and U9560 (N_9560,N_4541,N_2802);
nor U9561 (N_9561,N_638,N_475);
xnor U9562 (N_9562,N_131,N_2188);
and U9563 (N_9563,N_4391,N_3225);
or U9564 (N_9564,N_3375,N_4623);
xor U9565 (N_9565,N_1744,N_339);
xor U9566 (N_9566,N_1248,N_4802);
or U9567 (N_9567,N_3632,N_3147);
nand U9568 (N_9568,N_4786,N_3250);
xnor U9569 (N_9569,N_4604,N_384);
or U9570 (N_9570,N_421,N_3233);
and U9571 (N_9571,N_1846,N_1822);
and U9572 (N_9572,N_4910,N_1592);
or U9573 (N_9573,N_3046,N_2752);
nor U9574 (N_9574,N_4923,N_3368);
nand U9575 (N_9575,N_1520,N_2711);
nor U9576 (N_9576,N_2075,N_1996);
and U9577 (N_9577,N_2879,N_887);
xnor U9578 (N_9578,N_4752,N_4541);
and U9579 (N_9579,N_3339,N_3976);
xnor U9580 (N_9580,N_1342,N_2544);
and U9581 (N_9581,N_3403,N_2467);
or U9582 (N_9582,N_37,N_1899);
nor U9583 (N_9583,N_1733,N_3992);
or U9584 (N_9584,N_4598,N_1796);
and U9585 (N_9585,N_3312,N_3633);
or U9586 (N_9586,N_3264,N_368);
xnor U9587 (N_9587,N_1595,N_1426);
and U9588 (N_9588,N_4889,N_872);
nand U9589 (N_9589,N_4966,N_1998);
and U9590 (N_9590,N_2258,N_2244);
nor U9591 (N_9591,N_1431,N_2688);
nor U9592 (N_9592,N_1871,N_1237);
nor U9593 (N_9593,N_2548,N_2411);
nand U9594 (N_9594,N_31,N_3006);
and U9595 (N_9595,N_312,N_3055);
nor U9596 (N_9596,N_4433,N_1124);
nor U9597 (N_9597,N_694,N_2520);
nand U9598 (N_9598,N_4005,N_1721);
and U9599 (N_9599,N_2698,N_166);
or U9600 (N_9600,N_1540,N_848);
or U9601 (N_9601,N_3115,N_4767);
xor U9602 (N_9602,N_4428,N_4228);
nor U9603 (N_9603,N_202,N_1567);
nand U9604 (N_9604,N_4466,N_3883);
nand U9605 (N_9605,N_2730,N_1355);
nand U9606 (N_9606,N_2637,N_977);
nand U9607 (N_9607,N_3036,N_3428);
and U9608 (N_9608,N_561,N_3211);
and U9609 (N_9609,N_1197,N_4561);
or U9610 (N_9610,N_2147,N_2055);
and U9611 (N_9611,N_2662,N_4644);
xnor U9612 (N_9612,N_2042,N_2610);
and U9613 (N_9613,N_734,N_1089);
or U9614 (N_9614,N_358,N_3829);
nor U9615 (N_9615,N_3944,N_1084);
and U9616 (N_9616,N_2113,N_4006);
xnor U9617 (N_9617,N_1810,N_4284);
xnor U9618 (N_9618,N_4003,N_2861);
xnor U9619 (N_9619,N_4102,N_3147);
and U9620 (N_9620,N_2755,N_4537);
nand U9621 (N_9621,N_237,N_2127);
nor U9622 (N_9622,N_270,N_2865);
nor U9623 (N_9623,N_1912,N_1078);
nand U9624 (N_9624,N_3645,N_1552);
or U9625 (N_9625,N_1560,N_1352);
or U9626 (N_9626,N_4603,N_2022);
xnor U9627 (N_9627,N_3900,N_4701);
xnor U9628 (N_9628,N_1054,N_3793);
or U9629 (N_9629,N_2125,N_702);
or U9630 (N_9630,N_4608,N_3356);
or U9631 (N_9631,N_3458,N_3127);
and U9632 (N_9632,N_4968,N_4425);
or U9633 (N_9633,N_3094,N_3624);
and U9634 (N_9634,N_2271,N_1961);
xor U9635 (N_9635,N_2144,N_3207);
or U9636 (N_9636,N_2548,N_2489);
and U9637 (N_9637,N_4709,N_69);
or U9638 (N_9638,N_4308,N_1491);
and U9639 (N_9639,N_825,N_4429);
or U9640 (N_9640,N_1280,N_2049);
nor U9641 (N_9641,N_1309,N_4740);
or U9642 (N_9642,N_2488,N_4742);
nand U9643 (N_9643,N_3495,N_4237);
xnor U9644 (N_9644,N_3157,N_1011);
xor U9645 (N_9645,N_1776,N_1023);
xnor U9646 (N_9646,N_4829,N_114);
and U9647 (N_9647,N_3068,N_2370);
or U9648 (N_9648,N_1310,N_3279);
nor U9649 (N_9649,N_4639,N_4689);
xor U9650 (N_9650,N_4669,N_2673);
nand U9651 (N_9651,N_2347,N_929);
or U9652 (N_9652,N_788,N_2383);
or U9653 (N_9653,N_1150,N_2353);
nor U9654 (N_9654,N_389,N_2563);
and U9655 (N_9655,N_2121,N_4127);
and U9656 (N_9656,N_1253,N_2554);
and U9657 (N_9657,N_1693,N_158);
nor U9658 (N_9658,N_4599,N_542);
nand U9659 (N_9659,N_4645,N_3008);
or U9660 (N_9660,N_2489,N_1508);
or U9661 (N_9661,N_1642,N_3198);
nand U9662 (N_9662,N_2320,N_2989);
and U9663 (N_9663,N_3002,N_4574);
or U9664 (N_9664,N_3964,N_2897);
or U9665 (N_9665,N_2614,N_2105);
nand U9666 (N_9666,N_2181,N_507);
and U9667 (N_9667,N_3873,N_471);
and U9668 (N_9668,N_2787,N_4729);
xnor U9669 (N_9669,N_4523,N_3286);
nor U9670 (N_9670,N_4199,N_2030);
or U9671 (N_9671,N_4715,N_4488);
nand U9672 (N_9672,N_1879,N_275);
and U9673 (N_9673,N_2635,N_93);
or U9674 (N_9674,N_370,N_1333);
nor U9675 (N_9675,N_4278,N_2446);
nand U9676 (N_9676,N_4553,N_2085);
and U9677 (N_9677,N_1867,N_991);
nand U9678 (N_9678,N_1174,N_4019);
and U9679 (N_9679,N_4236,N_4445);
and U9680 (N_9680,N_1058,N_648);
or U9681 (N_9681,N_4646,N_3564);
or U9682 (N_9682,N_251,N_331);
or U9683 (N_9683,N_3873,N_2213);
and U9684 (N_9684,N_3632,N_2089);
xor U9685 (N_9685,N_2984,N_4792);
xor U9686 (N_9686,N_7,N_1583);
and U9687 (N_9687,N_3889,N_582);
xnor U9688 (N_9688,N_399,N_1380);
nor U9689 (N_9689,N_3021,N_593);
nor U9690 (N_9690,N_1987,N_178);
nand U9691 (N_9691,N_1078,N_119);
nor U9692 (N_9692,N_2689,N_518);
nand U9693 (N_9693,N_621,N_1400);
xnor U9694 (N_9694,N_2570,N_430);
nand U9695 (N_9695,N_2355,N_3704);
xor U9696 (N_9696,N_2222,N_394);
or U9697 (N_9697,N_143,N_4732);
nor U9698 (N_9698,N_911,N_2316);
and U9699 (N_9699,N_2966,N_1644);
and U9700 (N_9700,N_1260,N_1248);
nand U9701 (N_9701,N_3110,N_4193);
or U9702 (N_9702,N_2619,N_2920);
nand U9703 (N_9703,N_886,N_3168);
nand U9704 (N_9704,N_2161,N_4216);
xnor U9705 (N_9705,N_3117,N_4418);
nand U9706 (N_9706,N_3296,N_4378);
nor U9707 (N_9707,N_2949,N_4063);
xor U9708 (N_9708,N_1276,N_1846);
and U9709 (N_9709,N_4024,N_1386);
nand U9710 (N_9710,N_3905,N_1891);
nand U9711 (N_9711,N_4733,N_3789);
and U9712 (N_9712,N_194,N_3657);
xnor U9713 (N_9713,N_910,N_4793);
nand U9714 (N_9714,N_2160,N_3939);
nor U9715 (N_9715,N_3935,N_4680);
nand U9716 (N_9716,N_1238,N_2954);
or U9717 (N_9717,N_2182,N_4733);
and U9718 (N_9718,N_3737,N_745);
and U9719 (N_9719,N_1641,N_3850);
or U9720 (N_9720,N_4818,N_4837);
nor U9721 (N_9721,N_2832,N_2439);
and U9722 (N_9722,N_2569,N_3529);
xor U9723 (N_9723,N_3652,N_3359);
and U9724 (N_9724,N_4344,N_1261);
nor U9725 (N_9725,N_1148,N_4602);
xor U9726 (N_9726,N_2726,N_499);
xor U9727 (N_9727,N_3763,N_280);
nand U9728 (N_9728,N_2658,N_1106);
nor U9729 (N_9729,N_1779,N_4502);
and U9730 (N_9730,N_1739,N_41);
nor U9731 (N_9731,N_1504,N_143);
nand U9732 (N_9732,N_1774,N_2010);
xor U9733 (N_9733,N_484,N_4042);
xnor U9734 (N_9734,N_1712,N_1200);
xnor U9735 (N_9735,N_4490,N_4230);
xnor U9736 (N_9736,N_306,N_3446);
xnor U9737 (N_9737,N_2213,N_229);
nand U9738 (N_9738,N_4276,N_4755);
nor U9739 (N_9739,N_2986,N_4033);
nor U9740 (N_9740,N_1996,N_4361);
nand U9741 (N_9741,N_3659,N_636);
nor U9742 (N_9742,N_1227,N_2534);
nor U9743 (N_9743,N_4708,N_807);
or U9744 (N_9744,N_1335,N_2487);
nand U9745 (N_9745,N_1057,N_4645);
nor U9746 (N_9746,N_2045,N_3201);
nor U9747 (N_9747,N_4975,N_2534);
nand U9748 (N_9748,N_2209,N_3777);
nor U9749 (N_9749,N_4987,N_3562);
nand U9750 (N_9750,N_3765,N_1021);
xor U9751 (N_9751,N_4223,N_803);
nor U9752 (N_9752,N_421,N_4918);
or U9753 (N_9753,N_1004,N_4299);
or U9754 (N_9754,N_3156,N_562);
and U9755 (N_9755,N_821,N_4862);
and U9756 (N_9756,N_4265,N_370);
nor U9757 (N_9757,N_2787,N_1751);
xor U9758 (N_9758,N_4649,N_2143);
and U9759 (N_9759,N_2131,N_4573);
nand U9760 (N_9760,N_314,N_1571);
nor U9761 (N_9761,N_4918,N_1700);
nor U9762 (N_9762,N_4148,N_3086);
or U9763 (N_9763,N_614,N_3787);
nor U9764 (N_9764,N_944,N_4053);
xnor U9765 (N_9765,N_413,N_913);
nand U9766 (N_9766,N_2033,N_395);
or U9767 (N_9767,N_4993,N_3576);
nand U9768 (N_9768,N_3713,N_4793);
nand U9769 (N_9769,N_2616,N_3750);
or U9770 (N_9770,N_1395,N_692);
nor U9771 (N_9771,N_2253,N_2499);
xor U9772 (N_9772,N_2479,N_3692);
or U9773 (N_9773,N_4196,N_676);
nor U9774 (N_9774,N_4803,N_846);
and U9775 (N_9775,N_4124,N_1034);
nand U9776 (N_9776,N_1006,N_68);
nand U9777 (N_9777,N_413,N_3955);
nand U9778 (N_9778,N_2453,N_373);
xor U9779 (N_9779,N_1007,N_4353);
and U9780 (N_9780,N_2364,N_436);
xnor U9781 (N_9781,N_4517,N_2573);
and U9782 (N_9782,N_4096,N_3775);
and U9783 (N_9783,N_3631,N_643);
nor U9784 (N_9784,N_956,N_1042);
xnor U9785 (N_9785,N_4011,N_1357);
nor U9786 (N_9786,N_2138,N_341);
nand U9787 (N_9787,N_61,N_3122);
and U9788 (N_9788,N_2951,N_4788);
nor U9789 (N_9789,N_819,N_311);
or U9790 (N_9790,N_1853,N_4263);
nor U9791 (N_9791,N_5,N_2770);
or U9792 (N_9792,N_3131,N_1539);
nand U9793 (N_9793,N_485,N_1799);
or U9794 (N_9794,N_4939,N_1513);
and U9795 (N_9795,N_1115,N_4434);
and U9796 (N_9796,N_2197,N_725);
nor U9797 (N_9797,N_3370,N_2996);
or U9798 (N_9798,N_1564,N_512);
nand U9799 (N_9799,N_4577,N_2185);
nand U9800 (N_9800,N_603,N_2358);
nor U9801 (N_9801,N_1270,N_3553);
nand U9802 (N_9802,N_623,N_3809);
xnor U9803 (N_9803,N_3191,N_4758);
nor U9804 (N_9804,N_729,N_79);
xor U9805 (N_9805,N_4017,N_2587);
xor U9806 (N_9806,N_3831,N_4875);
xnor U9807 (N_9807,N_1427,N_493);
nor U9808 (N_9808,N_4272,N_4204);
nand U9809 (N_9809,N_3826,N_2863);
nand U9810 (N_9810,N_3608,N_1614);
and U9811 (N_9811,N_3974,N_2757);
nand U9812 (N_9812,N_4415,N_3103);
and U9813 (N_9813,N_4768,N_4);
nor U9814 (N_9814,N_4924,N_3458);
or U9815 (N_9815,N_1843,N_1446);
or U9816 (N_9816,N_3785,N_3689);
nor U9817 (N_9817,N_4701,N_1533);
xnor U9818 (N_9818,N_3042,N_4685);
and U9819 (N_9819,N_2498,N_2614);
nand U9820 (N_9820,N_2344,N_973);
or U9821 (N_9821,N_3853,N_2473);
nand U9822 (N_9822,N_1753,N_4617);
xnor U9823 (N_9823,N_3624,N_3256);
nand U9824 (N_9824,N_4344,N_3546);
or U9825 (N_9825,N_3116,N_3858);
and U9826 (N_9826,N_2227,N_4018);
nand U9827 (N_9827,N_216,N_2785);
or U9828 (N_9828,N_4889,N_762);
and U9829 (N_9829,N_1360,N_3302);
nand U9830 (N_9830,N_2795,N_3342);
nand U9831 (N_9831,N_547,N_1978);
or U9832 (N_9832,N_4998,N_3361);
or U9833 (N_9833,N_3211,N_4295);
nor U9834 (N_9834,N_3745,N_470);
nor U9835 (N_9835,N_107,N_1137);
nand U9836 (N_9836,N_69,N_2980);
or U9837 (N_9837,N_647,N_4931);
or U9838 (N_9838,N_3421,N_1671);
xor U9839 (N_9839,N_2785,N_345);
nor U9840 (N_9840,N_1649,N_4948);
nor U9841 (N_9841,N_496,N_2928);
or U9842 (N_9842,N_4779,N_4909);
nor U9843 (N_9843,N_176,N_3740);
or U9844 (N_9844,N_3928,N_189);
nand U9845 (N_9845,N_1174,N_3807);
xnor U9846 (N_9846,N_1564,N_2818);
and U9847 (N_9847,N_3423,N_3500);
nor U9848 (N_9848,N_4637,N_4067);
and U9849 (N_9849,N_2561,N_4648);
and U9850 (N_9850,N_4577,N_2586);
or U9851 (N_9851,N_3404,N_2932);
or U9852 (N_9852,N_4611,N_1089);
xor U9853 (N_9853,N_1899,N_1342);
nor U9854 (N_9854,N_3150,N_545);
nor U9855 (N_9855,N_3461,N_476);
or U9856 (N_9856,N_246,N_1418);
nand U9857 (N_9857,N_2773,N_282);
or U9858 (N_9858,N_855,N_2698);
and U9859 (N_9859,N_2478,N_4293);
and U9860 (N_9860,N_3965,N_1970);
xnor U9861 (N_9861,N_150,N_859);
nor U9862 (N_9862,N_541,N_3398);
or U9863 (N_9863,N_1052,N_4325);
nor U9864 (N_9864,N_1942,N_1404);
nor U9865 (N_9865,N_4500,N_3732);
nand U9866 (N_9866,N_3447,N_4334);
nor U9867 (N_9867,N_2845,N_1784);
xor U9868 (N_9868,N_2853,N_2452);
or U9869 (N_9869,N_599,N_3647);
nor U9870 (N_9870,N_2376,N_218);
or U9871 (N_9871,N_2771,N_2497);
or U9872 (N_9872,N_56,N_3044);
and U9873 (N_9873,N_339,N_1933);
nor U9874 (N_9874,N_3786,N_1593);
or U9875 (N_9875,N_63,N_1319);
xor U9876 (N_9876,N_3290,N_2005);
and U9877 (N_9877,N_1144,N_4606);
nand U9878 (N_9878,N_3889,N_3074);
xnor U9879 (N_9879,N_4869,N_2538);
nand U9880 (N_9880,N_1946,N_4318);
nor U9881 (N_9881,N_3316,N_2682);
and U9882 (N_9882,N_2712,N_4560);
and U9883 (N_9883,N_3782,N_1407);
nor U9884 (N_9884,N_3462,N_3846);
xnor U9885 (N_9885,N_1425,N_4574);
nor U9886 (N_9886,N_4169,N_2039);
nand U9887 (N_9887,N_4313,N_4285);
nor U9888 (N_9888,N_2819,N_568);
nand U9889 (N_9889,N_3019,N_906);
and U9890 (N_9890,N_1260,N_3416);
nand U9891 (N_9891,N_4747,N_4202);
nand U9892 (N_9892,N_1668,N_2269);
nand U9893 (N_9893,N_725,N_1417);
xnor U9894 (N_9894,N_2690,N_2581);
and U9895 (N_9895,N_3402,N_4119);
or U9896 (N_9896,N_1409,N_231);
xnor U9897 (N_9897,N_4259,N_4101);
and U9898 (N_9898,N_3417,N_4184);
nand U9899 (N_9899,N_4413,N_1686);
nand U9900 (N_9900,N_536,N_90);
or U9901 (N_9901,N_512,N_3952);
and U9902 (N_9902,N_3449,N_2416);
nor U9903 (N_9903,N_4874,N_2422);
xnor U9904 (N_9904,N_37,N_4237);
or U9905 (N_9905,N_4789,N_1918);
and U9906 (N_9906,N_4050,N_3555);
nor U9907 (N_9907,N_3590,N_4325);
xnor U9908 (N_9908,N_3320,N_4437);
nor U9909 (N_9909,N_2532,N_4866);
xnor U9910 (N_9910,N_3581,N_361);
xnor U9911 (N_9911,N_2020,N_2366);
or U9912 (N_9912,N_576,N_4254);
xnor U9913 (N_9913,N_3865,N_952);
xor U9914 (N_9914,N_710,N_764);
xor U9915 (N_9915,N_4897,N_2817);
nor U9916 (N_9916,N_1744,N_3050);
or U9917 (N_9917,N_3295,N_2574);
or U9918 (N_9918,N_4661,N_2335);
nand U9919 (N_9919,N_3872,N_3381);
or U9920 (N_9920,N_2903,N_3502);
nand U9921 (N_9921,N_958,N_701);
nor U9922 (N_9922,N_3717,N_3199);
and U9923 (N_9923,N_59,N_959);
nor U9924 (N_9924,N_1520,N_4420);
and U9925 (N_9925,N_2427,N_738);
xor U9926 (N_9926,N_4539,N_4385);
or U9927 (N_9927,N_4006,N_241);
nand U9928 (N_9928,N_669,N_2221);
or U9929 (N_9929,N_90,N_753);
xor U9930 (N_9930,N_4474,N_3452);
nor U9931 (N_9931,N_4820,N_2279);
nor U9932 (N_9932,N_1238,N_3680);
and U9933 (N_9933,N_753,N_3938);
and U9934 (N_9934,N_4961,N_1286);
nand U9935 (N_9935,N_3297,N_1749);
and U9936 (N_9936,N_3851,N_3762);
nor U9937 (N_9937,N_1003,N_3803);
xnor U9938 (N_9938,N_4406,N_4292);
nand U9939 (N_9939,N_2564,N_4776);
nor U9940 (N_9940,N_3285,N_3032);
or U9941 (N_9941,N_3925,N_4483);
or U9942 (N_9942,N_343,N_2700);
nand U9943 (N_9943,N_116,N_976);
and U9944 (N_9944,N_245,N_1829);
or U9945 (N_9945,N_4922,N_3976);
nor U9946 (N_9946,N_2931,N_3978);
nand U9947 (N_9947,N_1898,N_2459);
and U9948 (N_9948,N_3451,N_4856);
or U9949 (N_9949,N_2376,N_878);
nor U9950 (N_9950,N_1021,N_3871);
and U9951 (N_9951,N_3994,N_2417);
and U9952 (N_9952,N_3695,N_386);
nor U9953 (N_9953,N_4233,N_4777);
nand U9954 (N_9954,N_527,N_4665);
xor U9955 (N_9955,N_556,N_2443);
nand U9956 (N_9956,N_1152,N_126);
and U9957 (N_9957,N_2080,N_1524);
and U9958 (N_9958,N_844,N_4031);
and U9959 (N_9959,N_1636,N_3416);
nand U9960 (N_9960,N_2897,N_4451);
nand U9961 (N_9961,N_39,N_1160);
or U9962 (N_9962,N_3024,N_10);
or U9963 (N_9963,N_2034,N_1035);
nor U9964 (N_9964,N_2037,N_2225);
nor U9965 (N_9965,N_3913,N_2474);
nor U9966 (N_9966,N_3859,N_2753);
nor U9967 (N_9967,N_253,N_2337);
nor U9968 (N_9968,N_2214,N_4738);
and U9969 (N_9969,N_483,N_2834);
nand U9970 (N_9970,N_590,N_4936);
and U9971 (N_9971,N_3683,N_1398);
and U9972 (N_9972,N_706,N_2038);
or U9973 (N_9973,N_2810,N_429);
or U9974 (N_9974,N_2115,N_4755);
xnor U9975 (N_9975,N_1776,N_1658);
nand U9976 (N_9976,N_2207,N_292);
nor U9977 (N_9977,N_4721,N_361);
nand U9978 (N_9978,N_1582,N_2147);
xnor U9979 (N_9979,N_3908,N_1950);
nand U9980 (N_9980,N_3726,N_3393);
xnor U9981 (N_9981,N_2703,N_2131);
nor U9982 (N_9982,N_1226,N_3667);
xor U9983 (N_9983,N_3661,N_694);
xnor U9984 (N_9984,N_988,N_781);
xnor U9985 (N_9985,N_4230,N_838);
and U9986 (N_9986,N_2690,N_2572);
or U9987 (N_9987,N_3390,N_3763);
xnor U9988 (N_9988,N_345,N_1269);
nor U9989 (N_9989,N_1518,N_4521);
xor U9990 (N_9990,N_2479,N_3892);
nor U9991 (N_9991,N_586,N_946);
xnor U9992 (N_9992,N_861,N_3532);
nor U9993 (N_9993,N_1481,N_3744);
and U9994 (N_9994,N_1980,N_641);
nand U9995 (N_9995,N_1652,N_583);
and U9996 (N_9996,N_2143,N_3329);
nor U9997 (N_9997,N_2198,N_1670);
and U9998 (N_9998,N_1007,N_2007);
and U9999 (N_9999,N_1695,N_3057);
and U10000 (N_10000,N_5743,N_7856);
xnor U10001 (N_10001,N_6416,N_5716);
or U10002 (N_10002,N_8555,N_6451);
nor U10003 (N_10003,N_5019,N_7538);
nand U10004 (N_10004,N_9529,N_6097);
nand U10005 (N_10005,N_7158,N_6759);
nor U10006 (N_10006,N_9724,N_6757);
nor U10007 (N_10007,N_8739,N_9502);
nor U10008 (N_10008,N_7597,N_8842);
or U10009 (N_10009,N_6488,N_8805);
nand U10010 (N_10010,N_7672,N_8799);
and U10011 (N_10011,N_9609,N_8085);
xor U10012 (N_10012,N_5401,N_8229);
and U10013 (N_10013,N_6153,N_5062);
or U10014 (N_10014,N_9001,N_8408);
nand U10015 (N_10015,N_6010,N_9931);
nor U10016 (N_10016,N_9339,N_9872);
xor U10017 (N_10017,N_9287,N_5273);
xor U10018 (N_10018,N_6234,N_5519);
nand U10019 (N_10019,N_8852,N_6732);
and U10020 (N_10020,N_7199,N_7507);
and U10021 (N_10021,N_7652,N_6252);
and U10022 (N_10022,N_8250,N_9186);
nand U10023 (N_10023,N_8437,N_6976);
and U10024 (N_10024,N_6029,N_9436);
nor U10025 (N_10025,N_7426,N_6989);
or U10026 (N_10026,N_9024,N_9478);
nand U10027 (N_10027,N_6077,N_9362);
and U10028 (N_10028,N_5683,N_8557);
or U10029 (N_10029,N_8966,N_7907);
nor U10030 (N_10030,N_8271,N_9707);
and U10031 (N_10031,N_8477,N_5003);
nor U10032 (N_10032,N_7220,N_5837);
and U10033 (N_10033,N_8279,N_5241);
xor U10034 (N_10034,N_5321,N_5014);
nor U10035 (N_10035,N_8157,N_8330);
and U10036 (N_10036,N_7843,N_5574);
nor U10037 (N_10037,N_6668,N_8158);
nor U10038 (N_10038,N_5841,N_8562);
xnor U10039 (N_10039,N_5736,N_5784);
xnor U10040 (N_10040,N_6959,N_8201);
and U10041 (N_10041,N_9515,N_5714);
nand U10042 (N_10042,N_9503,N_6808);
xnor U10043 (N_10043,N_9979,N_5575);
nand U10044 (N_10044,N_9813,N_8683);
nand U10045 (N_10045,N_8320,N_6677);
and U10046 (N_10046,N_9603,N_8627);
nor U10047 (N_10047,N_9135,N_5506);
and U10048 (N_10048,N_5825,N_9884);
nand U10049 (N_10049,N_9610,N_9927);
and U10050 (N_10050,N_6586,N_5843);
nor U10051 (N_10051,N_9901,N_8749);
and U10052 (N_10052,N_6862,N_8273);
xor U10053 (N_10053,N_9162,N_7600);
nand U10054 (N_10054,N_5269,N_5620);
nor U10055 (N_10055,N_5525,N_9010);
nor U10056 (N_10056,N_8360,N_9561);
xnor U10057 (N_10057,N_6223,N_5383);
or U10058 (N_10058,N_9732,N_8440);
xor U10059 (N_10059,N_9743,N_8137);
nor U10060 (N_10060,N_7295,N_7928);
or U10061 (N_10061,N_6710,N_5036);
nand U10062 (N_10062,N_7228,N_8570);
and U10063 (N_10063,N_7513,N_5486);
nor U10064 (N_10064,N_7211,N_5319);
or U10065 (N_10065,N_7953,N_8632);
nand U10066 (N_10066,N_8057,N_8877);
nor U10067 (N_10067,N_9881,N_8608);
nor U10068 (N_10068,N_8192,N_8658);
nor U10069 (N_10069,N_5938,N_9595);
nor U10070 (N_10070,N_5758,N_7410);
nor U10071 (N_10071,N_8011,N_5667);
nand U10072 (N_10072,N_7607,N_5788);
or U10073 (N_10073,N_9134,N_5262);
nand U10074 (N_10074,N_6267,N_7742);
nor U10075 (N_10075,N_8630,N_5524);
and U10076 (N_10076,N_9768,N_8552);
or U10077 (N_10077,N_7684,N_7188);
nand U10078 (N_10078,N_8342,N_8663);
and U10079 (N_10079,N_6339,N_9267);
and U10080 (N_10080,N_7187,N_9656);
xor U10081 (N_10081,N_8776,N_8017);
or U10082 (N_10082,N_9705,N_8582);
xnor U10083 (N_10083,N_8080,N_8371);
nand U10084 (N_10084,N_9363,N_7519);
nor U10085 (N_10085,N_8896,N_9305);
xor U10086 (N_10086,N_7479,N_8003);
nand U10087 (N_10087,N_8078,N_6548);
or U10088 (N_10088,N_9941,N_5129);
nor U10089 (N_10089,N_8864,N_9326);
or U10090 (N_10090,N_8621,N_9952);
nor U10091 (N_10091,N_8432,N_6094);
nand U10092 (N_10092,N_7157,N_6038);
or U10093 (N_10093,N_7891,N_8024);
nor U10094 (N_10094,N_5451,N_7074);
nor U10095 (N_10095,N_6408,N_8275);
nor U10096 (N_10096,N_7235,N_5426);
and U10097 (N_10097,N_6600,N_5655);
nor U10098 (N_10098,N_8379,N_6888);
nor U10099 (N_10099,N_7952,N_6560);
or U10100 (N_10100,N_7807,N_6944);
or U10101 (N_10101,N_8083,N_6167);
nor U10102 (N_10102,N_8669,N_6333);
or U10103 (N_10103,N_7583,N_9421);
nor U10104 (N_10104,N_8269,N_8216);
nand U10105 (N_10105,N_8678,N_6680);
nand U10106 (N_10106,N_9713,N_9906);
nand U10107 (N_10107,N_5406,N_9585);
xnor U10108 (N_10108,N_8975,N_6442);
nand U10109 (N_10109,N_6265,N_8890);
nand U10110 (N_10110,N_5284,N_7564);
xnor U10111 (N_10111,N_5674,N_7967);
xnor U10112 (N_10112,N_6447,N_7333);
nand U10113 (N_10113,N_5007,N_7109);
nand U10114 (N_10114,N_9160,N_8266);
nand U10115 (N_10115,N_5992,N_9356);
xor U10116 (N_10116,N_8846,N_6222);
or U10117 (N_10117,N_9727,N_5404);
and U10118 (N_10118,N_7556,N_7795);
nor U10119 (N_10119,N_8052,N_9679);
or U10120 (N_10120,N_8478,N_7865);
nor U10121 (N_10121,N_5460,N_6357);
and U10122 (N_10122,N_9350,N_8455);
and U10123 (N_10123,N_6389,N_6512);
nand U10124 (N_10124,N_5698,N_9064);
xnor U10125 (N_10125,N_9265,N_7570);
nor U10126 (N_10126,N_5991,N_6742);
nor U10127 (N_10127,N_7822,N_9127);
nand U10128 (N_10128,N_9216,N_7572);
xor U10129 (N_10129,N_8285,N_6707);
and U10130 (N_10130,N_5447,N_8396);
and U10131 (N_10131,N_8809,N_8036);
nand U10132 (N_10132,N_8573,N_8998);
nand U10133 (N_10133,N_5098,N_8891);
and U10134 (N_10134,N_8999,N_9439);
or U10135 (N_10135,N_7540,N_5921);
or U10136 (N_10136,N_5564,N_7981);
xnor U10137 (N_10137,N_8122,N_8687);
nand U10138 (N_10138,N_8077,N_7728);
and U10139 (N_10139,N_7683,N_5597);
and U10140 (N_10140,N_7450,N_8177);
xnor U10141 (N_10141,N_8832,N_5151);
nor U10142 (N_10142,N_7924,N_7960);
nand U10143 (N_10143,N_6427,N_8466);
nor U10144 (N_10144,N_8480,N_8924);
or U10145 (N_10145,N_9678,N_8248);
nand U10146 (N_10146,N_7948,N_7330);
or U10147 (N_10147,N_7222,N_8067);
nor U10148 (N_10148,N_8114,N_8556);
and U10149 (N_10149,N_9379,N_8005);
xnor U10150 (N_10150,N_7251,N_9654);
xnor U10151 (N_10151,N_9956,N_7743);
and U10152 (N_10152,N_7255,N_8539);
xor U10153 (N_10153,N_6289,N_6392);
nand U10154 (N_10154,N_6486,N_9596);
xor U10155 (N_10155,N_5144,N_9555);
or U10156 (N_10156,N_5027,N_6510);
or U10157 (N_10157,N_7497,N_6343);
xnor U10158 (N_10158,N_9735,N_9976);
nand U10159 (N_10159,N_7879,N_5982);
nand U10160 (N_10160,N_5797,N_6918);
xor U10161 (N_10161,N_8131,N_7777);
or U10162 (N_10162,N_8037,N_8741);
and U10163 (N_10163,N_5711,N_5158);
xnor U10164 (N_10164,N_6605,N_8033);
or U10165 (N_10165,N_5817,N_8151);
nor U10166 (N_10166,N_8811,N_6365);
nor U10167 (N_10167,N_8344,N_9057);
nand U10168 (N_10168,N_7037,N_7551);
and U10169 (N_10169,N_8824,N_9950);
nand U10170 (N_10170,N_5851,N_7150);
or U10171 (N_10171,N_9761,N_9964);
nand U10172 (N_10172,N_8215,N_6549);
nor U10173 (N_10173,N_7403,N_8786);
nor U10174 (N_10174,N_9161,N_9327);
and U10175 (N_10175,N_7580,N_6579);
or U10176 (N_10176,N_5412,N_7798);
or U10177 (N_10177,N_7653,N_7820);
xor U10178 (N_10178,N_5068,N_6156);
or U10179 (N_10179,N_5505,N_8372);
xor U10180 (N_10180,N_5816,N_5111);
or U10181 (N_10181,N_9554,N_5940);
xor U10182 (N_10182,N_9907,N_7099);
nand U10183 (N_10183,N_9445,N_8921);
and U10184 (N_10184,N_8245,N_8093);
and U10185 (N_10185,N_6975,N_5916);
nor U10186 (N_10186,N_7462,N_7136);
and U10187 (N_10187,N_7951,N_7622);
or U10188 (N_10188,N_7306,N_8606);
or U10189 (N_10189,N_9206,N_6305);
or U10190 (N_10190,N_9259,N_9660);
nor U10191 (N_10191,N_6601,N_7522);
and U10192 (N_10192,N_8381,N_9062);
xor U10193 (N_10193,N_6613,N_6202);
and U10194 (N_10194,N_5004,N_9429);
or U10195 (N_10195,N_6482,N_9709);
nor U10196 (N_10196,N_8544,N_5353);
nor U10197 (N_10197,N_5117,N_7260);
xor U10198 (N_10198,N_6310,N_8542);
nand U10199 (N_10199,N_7353,N_9132);
xnor U10200 (N_10200,N_6940,N_7495);
or U10201 (N_10201,N_7598,N_7892);
and U10202 (N_10202,N_8563,N_6228);
xor U10203 (N_10203,N_6409,N_8291);
nand U10204 (N_10204,N_7297,N_8667);
xor U10205 (N_10205,N_5956,N_5185);
or U10206 (N_10206,N_6373,N_8348);
nand U10207 (N_10207,N_5116,N_7047);
xor U10208 (N_10208,N_6868,N_6595);
or U10209 (N_10209,N_6316,N_9408);
nor U10210 (N_10210,N_8431,N_7024);
nand U10211 (N_10211,N_5021,N_5266);
xor U10212 (N_10212,N_9310,N_7261);
or U10213 (N_10213,N_5918,N_5427);
nor U10214 (N_10214,N_6509,N_7417);
nor U10215 (N_10215,N_7853,N_7175);
nor U10216 (N_10216,N_7249,N_6514);
xnor U10217 (N_10217,N_7609,N_7758);
xnor U10218 (N_10218,N_5961,N_9980);
nand U10219 (N_10219,N_8347,N_6826);
and U10220 (N_10220,N_6647,N_6928);
nand U10221 (N_10221,N_8735,N_9215);
xor U10222 (N_10222,N_7613,N_9525);
or U10223 (N_10223,N_5678,N_9171);
nor U10224 (N_10224,N_8888,N_5696);
nor U10225 (N_10225,N_5310,N_9639);
nor U10226 (N_10226,N_5794,N_8117);
nor U10227 (N_10227,N_9164,N_8536);
nand U10228 (N_10228,N_7573,N_9295);
and U10229 (N_10229,N_7046,N_5218);
nor U10230 (N_10230,N_9203,N_7760);
nor U10231 (N_10231,N_9812,N_8341);
and U10232 (N_10232,N_8338,N_5490);
and U10233 (N_10233,N_6602,N_6456);
or U10234 (N_10234,N_6270,N_8754);
nor U10235 (N_10235,N_8618,N_8287);
nor U10236 (N_10236,N_5294,N_8700);
nor U10237 (N_10237,N_8583,N_6513);
and U10238 (N_10238,N_5933,N_7091);
nand U10239 (N_10239,N_6492,N_5687);
nor U10240 (N_10240,N_6268,N_5081);
nand U10241 (N_10241,N_6627,N_5782);
nand U10242 (N_10242,N_9366,N_9225);
xnor U10243 (N_10243,N_5779,N_6000);
and U10244 (N_10244,N_6069,N_6847);
xor U10245 (N_10245,N_6977,N_5077);
and U10246 (N_10246,N_7170,N_6922);
nand U10247 (N_10247,N_7088,N_8997);
nand U10248 (N_10248,N_9069,N_5413);
and U10249 (N_10249,N_6239,N_7991);
and U10250 (N_10250,N_5217,N_7398);
nand U10251 (N_10251,N_8985,N_5768);
nor U10252 (N_10252,N_7481,N_8064);
or U10253 (N_10253,N_7869,N_9170);
or U10254 (N_10254,N_7491,N_9005);
and U10255 (N_10255,N_7102,N_5285);
nor U10256 (N_10256,N_7367,N_8744);
nor U10257 (N_10257,N_6532,N_7282);
nand U10258 (N_10258,N_9462,N_8870);
or U10259 (N_10259,N_9371,N_6042);
nor U10260 (N_10260,N_9888,N_5156);
xnor U10261 (N_10261,N_7453,N_6886);
or U10262 (N_10262,N_8300,N_5610);
xnor U10263 (N_10263,N_5234,N_5160);
and U10264 (N_10264,N_5393,N_5330);
nand U10265 (N_10265,N_9521,N_8402);
and U10266 (N_10266,N_6429,N_8427);
nand U10267 (N_10267,N_8407,N_7802);
nor U10268 (N_10268,N_9229,N_6621);
or U10269 (N_10269,N_7900,N_6494);
xor U10270 (N_10270,N_9859,N_8254);
or U10271 (N_10271,N_9627,N_6506);
xnor U10272 (N_10272,N_8205,N_9681);
nand U10273 (N_10273,N_5465,N_7849);
xnor U10274 (N_10274,N_9833,N_7120);
nand U10275 (N_10275,N_8170,N_7499);
or U10276 (N_10276,N_6338,N_6947);
or U10277 (N_10277,N_9061,N_5015);
nor U10278 (N_10278,N_7016,N_5638);
and U10279 (N_10279,N_5442,N_6011);
nand U10280 (N_10280,N_9940,N_9255);
nor U10281 (N_10281,N_8740,N_8762);
nor U10282 (N_10282,N_9882,N_8858);
nor U10283 (N_10283,N_9054,N_7221);
and U10284 (N_10284,N_6235,N_6195);
nand U10285 (N_10285,N_5939,N_5508);
and U10286 (N_10286,N_7544,N_6511);
nand U10287 (N_10287,N_6583,N_8369);
and U10288 (N_10288,N_9332,N_6297);
nand U10289 (N_10289,N_9574,N_8127);
or U10290 (N_10290,N_8299,N_5229);
nand U10291 (N_10291,N_6303,N_7180);
nor U10292 (N_10292,N_7717,N_7234);
or U10293 (N_10293,N_8825,N_5879);
xnor U10294 (N_10294,N_5001,N_8867);
and U10295 (N_10295,N_8394,N_8847);
and U10296 (N_10296,N_6775,N_9273);
and U10297 (N_10297,N_7986,N_7394);
xor U10298 (N_10298,N_6271,N_9110);
or U10299 (N_10299,N_8804,N_5188);
or U10300 (N_10300,N_6971,N_9370);
nand U10301 (N_10301,N_5187,N_5346);
nand U10302 (N_10302,N_5484,N_6051);
xnor U10303 (N_10303,N_5733,N_9607);
and U10304 (N_10304,N_6585,N_8990);
xor U10305 (N_10305,N_7794,N_6708);
nand U10306 (N_10306,N_9424,N_8186);
and U10307 (N_10307,N_7686,N_9214);
nor U10308 (N_10308,N_7612,N_7941);
xnor U10309 (N_10309,N_6645,N_5553);
and U10310 (N_10310,N_6903,N_6430);
nand U10311 (N_10311,N_9891,N_5863);
xnor U10312 (N_10312,N_7662,N_6873);
or U10313 (N_10313,N_7217,N_9645);
and U10314 (N_10314,N_5417,N_5142);
nand U10315 (N_10315,N_5350,N_6230);
nand U10316 (N_10316,N_7329,N_6712);
xor U10317 (N_10317,N_7336,N_5225);
nand U10318 (N_10318,N_6170,N_5685);
or U10319 (N_10319,N_8717,N_9348);
xor U10320 (N_10320,N_7732,N_9114);
or U10321 (N_10321,N_8937,N_8983);
or U10322 (N_10322,N_5260,N_6899);
and U10323 (N_10323,N_8500,N_5541);
xor U10324 (N_10324,N_7937,N_8419);
xor U10325 (N_10325,N_8472,N_9205);
nand U10326 (N_10326,N_7006,N_5361);
nand U10327 (N_10327,N_6005,N_5497);
nand U10328 (N_10328,N_5201,N_6821);
nand U10329 (N_10329,N_6150,N_5325);
or U10330 (N_10330,N_8110,N_7880);
xnor U10331 (N_10331,N_8522,N_6876);
xor U10332 (N_10332,N_6299,N_9672);
or U10333 (N_10333,N_9826,N_5379);
nand U10334 (N_10334,N_6412,N_6795);
nor U10335 (N_10335,N_9663,N_9772);
nor U10336 (N_10336,N_6288,N_8682);
or U10337 (N_10337,N_5334,N_6452);
or U10338 (N_10338,N_6386,N_6898);
nor U10339 (N_10339,N_9376,N_9815);
and U10340 (N_10340,N_8958,N_6641);
nand U10341 (N_10341,N_6981,N_7793);
nor U10342 (N_10342,N_6371,N_9464);
nor U10343 (N_10343,N_7940,N_9676);
xor U10344 (N_10344,N_9232,N_5594);
or U10345 (N_10345,N_8212,N_7123);
nor U10346 (N_10346,N_9451,N_9150);
nand U10347 (N_10347,N_7774,N_7355);
or U10348 (N_10348,N_9290,N_6973);
nand U10349 (N_10349,N_6652,N_5555);
or U10350 (N_10350,N_8227,N_7989);
xnor U10351 (N_10351,N_5540,N_6151);
nand U10352 (N_10352,N_5086,N_5787);
or U10353 (N_10353,N_9105,N_8495);
and U10354 (N_10354,N_6220,N_8617);
xor U10355 (N_10355,N_6881,N_7232);
and U10356 (N_10356,N_8412,N_9612);
and U10357 (N_10357,N_5141,N_5504);
or U10358 (N_10358,N_8593,N_7862);
xor U10359 (N_10359,N_8884,N_8878);
nor U10360 (N_10360,N_5898,N_7208);
nand U10361 (N_10361,N_6073,N_9702);
and U10362 (N_10362,N_6395,N_8054);
and U10363 (N_10363,N_8920,N_5263);
and U10364 (N_10364,N_9988,N_9674);
nand U10365 (N_10365,N_9469,N_6672);
nor U10366 (N_10366,N_6980,N_8359);
nor U10367 (N_10367,N_7008,N_7974);
or U10368 (N_10368,N_9869,N_9716);
and U10369 (N_10369,N_7466,N_5029);
or U10370 (N_10370,N_8088,N_5643);
or U10371 (N_10371,N_7325,N_8420);
nand U10372 (N_10372,N_9775,N_5513);
xnor U10373 (N_10373,N_9092,N_9159);
xor U10374 (N_10374,N_7811,N_5205);
nor U10375 (N_10375,N_8189,N_8084);
nor U10376 (N_10376,N_6747,N_7204);
nor U10377 (N_10377,N_9182,N_7542);
nor U10378 (N_10378,N_6032,N_8406);
and U10379 (N_10379,N_8453,N_7801);
xor U10380 (N_10380,N_6105,N_7553);
nor U10381 (N_10381,N_8863,N_8032);
and U10382 (N_10382,N_7831,N_8709);
xnor U10383 (N_10383,N_8268,N_6469);
nand U10384 (N_10384,N_5291,N_6164);
or U10385 (N_10385,N_5152,N_5060);
and U10386 (N_10386,N_5536,N_7638);
and U10387 (N_10387,N_8307,N_6114);
and U10388 (N_10388,N_5411,N_5778);
or U10389 (N_10389,N_6694,N_5629);
xor U10390 (N_10390,N_7098,N_8520);
nor U10391 (N_10391,N_7292,N_5588);
xnor U10392 (N_10392,N_6612,N_5599);
and U10393 (N_10393,N_7778,N_7510);
nor U10394 (N_10394,N_7428,N_7000);
nor U10395 (N_10395,N_9359,N_6183);
and U10396 (N_10396,N_9741,N_7281);
nand U10397 (N_10397,N_9151,N_5755);
nand U10398 (N_10398,N_7841,N_9999);
xnor U10399 (N_10399,N_6537,N_9187);
nor U10400 (N_10400,N_9841,N_9994);
xnor U10401 (N_10401,N_7197,N_6807);
xnor U10402 (N_10402,N_7119,N_7272);
nor U10403 (N_10403,N_9051,N_9116);
xnor U10404 (N_10404,N_7241,N_9889);
and U10405 (N_10405,N_5010,N_5011);
and U10406 (N_10406,N_6120,N_8029);
nand U10407 (N_10407,N_5181,N_9819);
and U10408 (N_10408,N_5364,N_5979);
nor U10409 (N_10409,N_5226,N_9723);
nor U10410 (N_10410,N_5198,N_5178);
or U10411 (N_10411,N_7177,N_8767);
or U10412 (N_10412,N_5107,N_7547);
and U10413 (N_10413,N_5924,N_6019);
nor U10414 (N_10414,N_8071,N_5750);
nand U10415 (N_10415,N_8930,N_7144);
nand U10416 (N_10416,N_5022,N_6967);
nand U10417 (N_10417,N_5623,N_8725);
and U10418 (N_10418,N_7876,N_9306);
and U10419 (N_10419,N_8885,N_7302);
nand U10420 (N_10420,N_5164,N_6589);
and U10421 (N_10421,N_5071,N_6180);
nand U10422 (N_10422,N_6609,N_6477);
nor U10423 (N_10423,N_5416,N_7451);
xnor U10424 (N_10424,N_7032,N_6246);
nand U10425 (N_10425,N_9349,N_7238);
and U10426 (N_10426,N_9280,N_8236);
or U10427 (N_10427,N_6705,N_9825);
xor U10428 (N_10428,N_6330,N_5231);
and U10429 (N_10429,N_8604,N_6553);
xor U10430 (N_10430,N_5532,N_9294);
and U10431 (N_10431,N_9410,N_5965);
and U10432 (N_10432,N_9246,N_7995);
xor U10433 (N_10433,N_6340,N_6249);
xor U10434 (N_10434,N_8730,N_8311);
and U10435 (N_10435,N_8546,N_6772);
nand U10436 (N_10436,N_5437,N_7723);
or U10437 (N_10437,N_6162,N_5814);
and U10438 (N_10438,N_8686,N_7964);
xnor U10439 (N_10439,N_8043,N_5405);
or U10440 (N_10440,N_8816,N_8304);
and U10441 (N_10441,N_7909,N_9773);
nor U10442 (N_10442,N_9390,N_5340);
nand U10443 (N_10443,N_9354,N_5089);
or U10444 (N_10444,N_6804,N_9067);
and U10445 (N_10445,N_6467,N_8684);
nor U10446 (N_10446,N_7141,N_8136);
nand U10447 (N_10447,N_7184,N_6474);
xnor U10448 (N_10448,N_6367,N_7867);
and U10449 (N_10449,N_8174,N_7489);
nand U10450 (N_10450,N_7602,N_9947);
xor U10451 (N_10451,N_9423,N_7796);
or U10452 (N_10452,N_6139,N_5335);
or U10453 (N_10453,N_8302,N_7779);
nand U10454 (N_10454,N_6161,N_9873);
or U10455 (N_10455,N_5562,N_8833);
and U10456 (N_10456,N_8397,N_6013);
nand U10457 (N_10457,N_5966,N_5084);
and U10458 (N_10458,N_9890,N_6885);
or U10459 (N_10459,N_6949,N_7029);
or U10460 (N_10460,N_7111,N_6352);
nor U10461 (N_10461,N_8538,N_7198);
nand U10462 (N_10462,N_8792,N_9718);
nand U10463 (N_10463,N_5927,N_7165);
nor U10464 (N_10464,N_5095,N_7461);
xnor U10465 (N_10465,N_9567,N_5292);
nand U10466 (N_10466,N_5547,N_7915);
nor U10467 (N_10467,N_9626,N_5728);
xnor U10468 (N_10468,N_7244,N_6072);
and U10469 (N_10469,N_5018,N_7236);
xor U10470 (N_10470,N_5873,N_8906);
xnor U10471 (N_10471,N_6950,N_5516);
nor U10472 (N_10472,N_8654,N_7945);
nor U10473 (N_10473,N_8610,N_5835);
nor U10474 (N_10474,N_7344,N_6279);
nand U10475 (N_10475,N_9406,N_7145);
and U10476 (N_10476,N_7289,N_5131);
and U10477 (N_10477,N_7508,N_6901);
or U10478 (N_10478,N_6358,N_9018);
xor U10479 (N_10479,N_8973,N_7746);
xor U10480 (N_10480,N_5351,N_5459);
xnor U10481 (N_10481,N_6264,N_5359);
nor U10482 (N_10482,N_6656,N_7854);
nand U10483 (N_10483,N_9427,N_5043);
nand U10484 (N_10484,N_7017,N_5313);
nand U10485 (N_10485,N_9396,N_6536);
xor U10486 (N_10486,N_7106,N_9892);
or U10487 (N_10487,N_7923,N_5434);
or U10488 (N_10488,N_8154,N_6729);
or U10489 (N_10489,N_5414,N_6178);
and U10490 (N_10490,N_9395,N_7290);
xor U10491 (N_10491,N_9028,N_6021);
xor U10492 (N_10492,N_8991,N_9447);
xnor U10493 (N_10493,N_6762,N_5368);
and U10494 (N_10494,N_5661,N_9081);
xnor U10495 (N_10495,N_7692,N_9830);
or U10496 (N_10496,N_9391,N_5469);
and U10497 (N_10497,N_9719,N_6052);
and U10498 (N_10498,N_7690,N_9043);
xnor U10499 (N_10499,N_6250,N_7322);
nor U10500 (N_10500,N_9856,N_5509);
and U10501 (N_10501,N_9703,N_9085);
nand U10502 (N_10502,N_8944,N_6860);
nor U10503 (N_10503,N_5170,N_6321);
or U10504 (N_10504,N_7166,N_8492);
or U10505 (N_10505,N_5482,N_8993);
or U10506 (N_10506,N_8979,N_7472);
and U10507 (N_10507,N_8642,N_8637);
nor U10508 (N_10508,N_5637,N_6640);
and U10509 (N_10509,N_7335,N_7339);
nor U10510 (N_10510,N_5867,N_6720);
and U10511 (N_10511,N_9806,N_8599);
and U10512 (N_10512,N_6314,N_7870);
and U10513 (N_10513,N_8162,N_6691);
or U10514 (N_10514,N_9250,N_5189);
xor U10515 (N_10515,N_9710,N_5862);
nand U10516 (N_10516,N_7716,N_8872);
or U10517 (N_10517,N_8156,N_7360);
or U10518 (N_10518,N_9090,N_7294);
and U10519 (N_10519,N_7040,N_7087);
and U10520 (N_10520,N_5688,N_7825);
nand U10521 (N_10521,N_8545,N_7308);
and U10522 (N_10522,N_8075,N_8173);
nor U10523 (N_10523,N_6820,N_8855);
xnor U10524 (N_10524,N_9628,N_5311);
xor U10525 (N_10525,N_7803,N_8515);
nand U10526 (N_10526,N_6085,N_9572);
nor U10527 (N_10527,N_7035,N_6238);
nor U10528 (N_10528,N_6123,N_7471);
xnor U10529 (N_10529,N_6964,N_7839);
or U10530 (N_10530,N_7557,N_6112);
nand U10531 (N_10531,N_5571,N_6438);
nor U10532 (N_10532,N_7832,N_6923);
nand U10533 (N_10533,N_8380,N_6206);
and U10534 (N_10534,N_9934,N_7163);
or U10535 (N_10535,N_5283,N_8796);
nor U10536 (N_10536,N_9341,N_6133);
or U10537 (N_10537,N_5208,N_6622);
nand U10538 (N_10538,N_9311,N_9983);
nand U10539 (N_10539,N_6154,N_8827);
nor U10540 (N_10540,N_9477,N_8178);
and U10541 (N_10541,N_6909,N_6660);
or U10542 (N_10542,N_9823,N_7435);
nand U10543 (N_10543,N_7068,N_7515);
nand U10544 (N_10544,N_7164,N_6683);
xnor U10545 (N_10545,N_6911,N_7757);
or U10546 (N_10546,N_9333,N_6990);
or U10547 (N_10547,N_8274,N_5120);
and U10548 (N_10548,N_6778,N_8566);
or U10549 (N_10549,N_6382,N_9898);
and U10550 (N_10550,N_8228,N_6972);
or U10551 (N_10551,N_8176,N_9293);
and U10552 (N_10552,N_5920,N_9103);
and U10553 (N_10553,N_5093,N_6015);
and U10554 (N_10554,N_9321,N_6527);
nor U10555 (N_10555,N_5658,N_8022);
nor U10556 (N_10556,N_6730,N_7056);
nand U10557 (N_10557,N_6931,N_6484);
nand U10558 (N_10558,N_8184,N_9699);
xor U10559 (N_10559,N_6725,N_5054);
and U10560 (N_10560,N_8124,N_6070);
or U10561 (N_10561,N_8977,N_9531);
xor U10562 (N_10562,N_9641,N_5202);
and U10563 (N_10563,N_9975,N_9494);
or U10564 (N_10564,N_5183,N_8561);
nor U10565 (N_10565,N_5849,N_9543);
or U10566 (N_10566,N_8710,N_9909);
nor U10567 (N_10567,N_5650,N_7376);
and U10568 (N_10568,N_5922,N_5384);
nor U10569 (N_10569,N_8759,N_5094);
xor U10570 (N_10570,N_9811,N_6925);
and U10571 (N_10571,N_5605,N_5478);
nor U10572 (N_10572,N_9244,N_9506);
xor U10573 (N_10573,N_7590,N_7110);
or U10574 (N_10574,N_5549,N_7483);
and U10575 (N_10575,N_7064,N_9692);
xnor U10576 (N_10576,N_9108,N_5378);
and U10577 (N_10577,N_5125,N_5489);
xor U10578 (N_10578,N_5430,N_9600);
xor U10579 (N_10579,N_9804,N_9698);
xor U10580 (N_10580,N_5828,N_5893);
nand U10581 (N_10581,N_9433,N_6719);
nor U10582 (N_10582,N_8336,N_9517);
xor U10583 (N_10583,N_6397,N_7620);
nand U10584 (N_10584,N_7767,N_6059);
or U10585 (N_10585,N_6750,N_7762);
or U10586 (N_10586,N_6086,N_7368);
xnor U10587 (N_10587,N_6581,N_7399);
xor U10588 (N_10588,N_8375,N_6004);
and U10589 (N_10589,N_7894,N_6460);
xor U10590 (N_10590,N_7725,N_5507);
nor U10591 (N_10591,N_6377,N_9711);
nor U10592 (N_10592,N_7284,N_6364);
or U10593 (N_10593,N_9495,N_8012);
and U10594 (N_10594,N_5352,N_6446);
xnor U10595 (N_10595,N_8652,N_8272);
and U10596 (N_10596,N_6251,N_5477);
nand U10597 (N_10597,N_9669,N_5753);
nor U10598 (N_10598,N_5989,N_8760);
or U10599 (N_10599,N_9516,N_9673);
and U10600 (N_10600,N_6044,N_8028);
nand U10601 (N_10601,N_8756,N_8413);
nor U10602 (N_10602,N_6906,N_5031);
nor U10603 (N_10603,N_6221,N_6748);
or U10604 (N_10604,N_7392,N_7206);
xor U10605 (N_10605,N_9850,N_5288);
or U10606 (N_10606,N_8309,N_6796);
xor U10607 (N_10607,N_6932,N_9185);
nand U10608 (N_10608,N_5423,N_5847);
xor U10609 (N_10609,N_9158,N_8059);
or U10610 (N_10610,N_5075,N_5207);
or U10611 (N_10611,N_6121,N_9799);
and U10612 (N_10612,N_8788,N_7840);
and U10613 (N_10613,N_5398,N_9649);
nor U10614 (N_10614,N_8263,N_6929);
and U10615 (N_10615,N_6328,N_8861);
and U10616 (N_10616,N_6100,N_8010);
xnor U10617 (N_10617,N_9328,N_8871);
xnor U10618 (N_10618,N_6275,N_7625);
nand U10619 (N_10619,N_9721,N_7500);
nor U10620 (N_10620,N_5567,N_7946);
xor U10621 (N_10621,N_8535,N_8956);
or U10622 (N_10622,N_8649,N_9760);
and U10623 (N_10623,N_5037,N_8079);
nand U10624 (N_10624,N_8253,N_9720);
nor U10625 (N_10625,N_9714,N_7022);
and U10626 (N_10626,N_9694,N_5586);
and U10627 (N_10627,N_9284,N_7711);
and U10628 (N_10628,N_5885,N_6788);
or U10629 (N_10629,N_9917,N_9510);
and U10630 (N_10630,N_5689,N_6383);
and U10631 (N_10631,N_5391,N_6942);
xnor U10632 (N_10632,N_9345,N_9569);
or U10633 (N_10633,N_8941,N_5595);
nor U10634 (N_10634,N_6493,N_8260);
nand U10635 (N_10635,N_7484,N_7162);
nor U10636 (N_10636,N_6002,N_8175);
nand U10637 (N_10637,N_8167,N_8957);
and U10638 (N_10638,N_7469,N_9896);
or U10639 (N_10639,N_5474,N_6814);
nand U10640 (N_10640,N_6580,N_8246);
nor U10641 (N_10641,N_8945,N_6381);
xnor U10642 (N_10642,N_7280,N_5118);
and U10643 (N_10643,N_5407,N_9014);
xor U10644 (N_10644,N_8065,N_8249);
xnor U10645 (N_10645,N_7671,N_8913);
xnor U10646 (N_10646,N_7097,N_7262);
nor U10647 (N_10647,N_6472,N_5140);
nand U10648 (N_10648,N_7784,N_9682);
nor U10649 (N_10649,N_7722,N_9473);
xnor U10650 (N_10650,N_5487,N_5772);
xnor U10651 (N_10651,N_6090,N_7247);
or U10652 (N_10652,N_7709,N_7385);
or U10653 (N_10653,N_5115,N_8994);
or U10654 (N_10654,N_6630,N_7738);
xor U10655 (N_10655,N_7407,N_8257);
xnor U10656 (N_10656,N_6274,N_5360);
nand U10657 (N_10657,N_9374,N_9653);
xor U10658 (N_10658,N_9832,N_5278);
or U10659 (N_10659,N_8335,N_5357);
nor U10660 (N_10660,N_6877,N_9706);
and U10661 (N_10661,N_9211,N_6777);
and U10662 (N_10662,N_9008,N_8423);
and U10663 (N_10663,N_5826,N_5827);
and U10664 (N_10664,N_5771,N_6674);
xnor U10665 (N_10665,N_8537,N_6017);
or U10666 (N_10666,N_7473,N_5631);
xor U10667 (N_10667,N_9996,N_6434);
xor U10668 (N_10668,N_9748,N_6829);
nor U10669 (N_10669,N_7025,N_6917);
or U10670 (N_10670,N_6780,N_8363);
or U10671 (N_10671,N_6812,N_5972);
nor U10672 (N_10672,N_5559,N_8531);
or U10673 (N_10673,N_5237,N_9693);
or U10674 (N_10674,N_8231,N_8699);
nand U10675 (N_10675,N_9109,N_5366);
nor U10676 (N_10676,N_5815,N_8401);
xor U10677 (N_10677,N_6626,N_8690);
xnor U10678 (N_10678,N_6620,N_7051);
nand U10679 (N_10679,N_5764,N_7081);
nor U10680 (N_10680,N_9136,N_7543);
nand U10681 (N_10681,N_6496,N_9807);
xor U10682 (N_10682,N_5734,N_7458);
and U10683 (N_10683,N_7182,N_7026);
and U10684 (N_10684,N_6521,N_8448);
and U10685 (N_10685,N_9128,N_5880);
xor U10686 (N_10686,N_5840,N_5641);
nor U10687 (N_10687,N_7388,N_6457);
nand U10688 (N_10688,N_8283,N_7303);
xnor U10689 (N_10689,N_5067,N_8575);
nor U10690 (N_10690,N_5980,N_5791);
and U10691 (N_10691,N_8770,N_8826);
and U10692 (N_10692,N_9876,N_5762);
xor U10693 (N_10693,N_7786,N_5611);
or U10694 (N_10694,N_6026,N_6827);
or U10695 (N_10695,N_6131,N_8479);
or U10696 (N_10696,N_5727,N_7943);
nand U10697 (N_10697,N_7107,N_7581);
and U10698 (N_10698,N_7124,N_6722);
or U10699 (N_10699,N_9455,N_7352);
and U10700 (N_10700,N_8806,N_9838);
or U10701 (N_10701,N_7408,N_9000);
or U10702 (N_10702,N_5389,N_8595);
and U10703 (N_10703,N_7586,N_5370);
and U10704 (N_10704,N_8499,N_9144);
xor U10705 (N_10705,N_7808,N_6767);
nor U10706 (N_10706,N_5006,N_8326);
nand U10707 (N_10707,N_5860,N_9659);
and U10708 (N_10708,N_6740,N_7372);
or U10709 (N_10709,N_7833,N_8035);
xnor U10710 (N_10710,N_5109,N_9526);
xnor U10711 (N_10711,N_6577,N_5162);
nor U10712 (N_10712,N_9686,N_9604);
or U10713 (N_10713,N_5177,N_5561);
nor U10714 (N_10714,N_6398,N_8679);
or U10715 (N_10715,N_5254,N_7756);
xor U10716 (N_10716,N_5929,N_7185);
or U10717 (N_10717,N_5646,N_5228);
and U10718 (N_10718,N_9095,N_9454);
and U10719 (N_10719,N_8881,N_8485);
xor U10720 (N_10720,N_5382,N_7440);
xnor U10721 (N_10721,N_6046,N_9071);
xnor U10722 (N_10722,N_5420,N_8925);
nand U10723 (N_10723,N_9755,N_9750);
xor U10724 (N_10724,N_8633,N_6113);
nor U10725 (N_10725,N_9809,N_8066);
xnor U10726 (N_10726,N_6968,N_7886);
nand U10727 (N_10727,N_6341,N_7980);
and U10728 (N_10728,N_5617,N_7918);
or U10729 (N_10729,N_9082,N_5299);
and U10730 (N_10730,N_9446,N_6089);
xnor U10731 (N_10731,N_8600,N_7210);
xnor U10732 (N_10732,N_7882,N_5954);
nand U10733 (N_10733,N_6960,N_9323);
nor U10734 (N_10734,N_7094,N_6181);
nand U10735 (N_10735,N_9708,N_8619);
or U10736 (N_10736,N_6802,N_7701);
nand U10737 (N_10737,N_8421,N_7475);
nand U10738 (N_10738,N_5510,N_6501);
nand U10739 (N_10739,N_8962,N_5809);
nor U10740 (N_10740,N_6902,N_9858);
and U10741 (N_10741,N_8434,N_7871);
nor U10742 (N_10742,N_6558,N_5763);
nor U10743 (N_10743,N_7151,N_8724);
or U10744 (N_10744,N_7276,N_6394);
and U10745 (N_10745,N_6449,N_7651);
and U10746 (N_10746,N_5433,N_9304);
or U10747 (N_10747,N_6978,N_9904);
xnor U10748 (N_10748,N_7978,N_7283);
and U10749 (N_10749,N_8109,N_5362);
nor U10750 (N_10750,N_8384,N_5642);
nor U10751 (N_10751,N_8830,N_7036);
or U10752 (N_10752,N_7212,N_8643);
nor U10753 (N_10753,N_6410,N_7114);
or U10754 (N_10754,N_9793,N_9801);
nor U10755 (N_10755,N_5348,N_6024);
and U10756 (N_10756,N_7585,N_7769);
xnor U10757 (N_10757,N_9033,N_7524);
and U10758 (N_10758,N_5239,N_5876);
and U10759 (N_10759,N_7341,N_5881);
and U10760 (N_10760,N_8651,N_5537);
nand U10761 (N_10761,N_7468,N_6143);
nor U10762 (N_10762,N_9301,N_5977);
or U10763 (N_10763,N_8668,N_5221);
or U10764 (N_10764,N_7396,N_5634);
nand U10765 (N_10765,N_7639,N_8940);
nand U10766 (N_10766,N_5316,N_8696);
or U10767 (N_10767,N_6716,N_8390);
and U10768 (N_10768,N_7614,N_8954);
nor U10769 (N_10769,N_8992,N_5886);
and U10770 (N_10770,N_5846,N_5978);
nand U10771 (N_10771,N_8547,N_8130);
or U10772 (N_10772,N_5830,N_7791);
nor U10773 (N_10773,N_9180,N_5122);
nand U10774 (N_10774,N_8422,N_8284);
and U10775 (N_10775,N_5590,N_6604);
nor U10776 (N_10776,N_8625,N_6618);
or U10777 (N_10777,N_6666,N_7171);
or U10778 (N_10778,N_7447,N_9951);
and U10779 (N_10779,N_7670,N_8337);
nand U10780 (N_10780,N_7868,N_9605);
and U10781 (N_10781,N_9897,N_8521);
nand U10782 (N_10782,N_5545,N_5580);
and U10783 (N_10783,N_5964,N_7237);
or U10784 (N_10784,N_7009,N_6129);
xnor U10785 (N_10785,N_6280,N_5041);
nor U10786 (N_10786,N_5626,N_7193);
nor U10787 (N_10787,N_6118,N_7628);
nor U10788 (N_10788,N_5960,N_9428);
or U10789 (N_10789,N_9153,N_5328);
nor U10790 (N_10790,N_8780,N_9101);
nor U10791 (N_10791,N_9399,N_5377);
or U10792 (N_10792,N_9191,N_5431);
nand U10793 (N_10793,N_9549,N_6502);
nand U10794 (N_10794,N_6065,N_6603);
or U10795 (N_10795,N_9272,N_6561);
and U10796 (N_10796,N_7361,N_9300);
nand U10797 (N_10797,N_8771,N_9420);
nor U10798 (N_10798,N_5079,N_7582);
xor U10799 (N_10799,N_7323,N_6662);
or U10800 (N_10800,N_7270,N_9118);
and U10801 (N_10801,N_5531,N_6594);
or U10802 (N_10802,N_9021,N_8111);
or U10803 (N_10803,N_6322,N_5955);
and U10804 (N_10804,N_8578,N_7874);
xor U10805 (N_10805,N_7837,N_6701);
nand U10806 (N_10806,N_7365,N_7359);
xnor U10807 (N_10807,N_9683,N_5251);
nand U10808 (N_10808,N_5676,N_5725);
nand U10809 (N_10809,N_5705,N_8040);
nand U10810 (N_10810,N_6992,N_5833);
or U10811 (N_10811,N_6215,N_9668);
and U10812 (N_10812,N_7438,N_6282);
nand U10813 (N_10813,N_7888,N_9509);
nand U10814 (N_10814,N_7754,N_9622);
xor U10815 (N_10815,N_9107,N_8584);
nand U10816 (N_10816,N_6646,N_9080);
xor U10817 (N_10817,N_5498,N_9177);
xor U10818 (N_10818,N_7286,N_6489);
nand U10819 (N_10819,N_5056,N_6490);
nor U10820 (N_10820,N_5495,N_9369);
xnor U10821 (N_10821,N_6713,N_9857);
nand U10822 (N_10822,N_5926,N_9816);
nand U10823 (N_10823,N_9523,N_9296);
xnor U10824 (N_10824,N_5473,N_5822);
or U10825 (N_10825,N_7358,N_8484);
and U10826 (N_10826,N_6999,N_8353);
nand U10827 (N_10827,N_6669,N_8923);
xnor U10828 (N_10828,N_7587,N_8355);
or U10829 (N_10829,N_5930,N_9288);
or U10830 (N_10830,N_7863,N_9093);
or U10831 (N_10831,N_6919,N_9285);
xnor U10832 (N_10832,N_8609,N_8482);
and U10833 (N_10833,N_6840,N_9237);
nand U10834 (N_10834,N_9416,N_9277);
and U10835 (N_10835,N_5657,N_6704);
nor U10836 (N_10836,N_9539,N_7082);
nand U10837 (N_10837,N_6035,N_9945);
nor U10838 (N_10838,N_6770,N_7730);
nand U10839 (N_10839,N_8091,N_6284);
and U10840 (N_10840,N_7054,N_6728);
and U10841 (N_10841,N_6961,N_8405);
or U10842 (N_10842,N_7264,N_6296);
or U10843 (N_10843,N_6768,N_7389);
xor U10844 (N_10844,N_9330,N_5773);
or U10845 (N_10845,N_6634,N_7851);
or U10846 (N_10846,N_6657,N_5408);
and U10847 (N_10847,N_6459,N_6945);
and U10848 (N_10848,N_9995,N_6499);
nand U10849 (N_10849,N_8144,N_6593);
and U10850 (N_10850,N_9695,N_8807);
or U10851 (N_10851,N_6592,N_7809);
or U10852 (N_10852,N_5745,N_7893);
or U10853 (N_10853,N_7657,N_7216);
or U10854 (N_10854,N_5538,N_9157);
xnor U10855 (N_10855,N_6053,N_6791);
xor U10856 (N_10856,N_5697,N_5191);
xnor U10857 (N_10857,N_5558,N_7565);
nand U10858 (N_10858,N_9233,N_6141);
nor U10859 (N_10859,N_9015,N_5517);
or U10860 (N_10860,N_7311,N_8290);
nand U10861 (N_10861,N_7736,N_6880);
nor U10862 (N_10862,N_7050,N_6998);
and U10863 (N_10863,N_5645,N_8876);
nor U10864 (N_10864,N_9998,N_5857);
or U10865 (N_10865,N_7030,N_5543);
xor U10866 (N_10866,N_6095,N_7420);
or U10867 (N_10867,N_5059,N_8383);
or U10868 (N_10868,N_5195,N_9106);
xor U10869 (N_10869,N_5952,N_7340);
nand U10870 (N_10870,N_7337,N_5604);
or U10871 (N_10871,N_6001,N_9261);
xor U10872 (N_10872,N_9091,N_8164);
and U10873 (N_10873,N_9864,N_9959);
nand U10874 (N_10874,N_9032,N_6743);
xnor U10875 (N_10875,N_5962,N_5692);
nor U10876 (N_10876,N_7086,N_7305);
nor U10877 (N_10877,N_6294,N_8911);
xor U10878 (N_10878,N_5320,N_8854);
nand U10879 (N_10879,N_8317,N_6838);
nand U10880 (N_10880,N_5168,N_9452);
or U10881 (N_10881,N_7299,N_5103);
nor U10882 (N_10882,N_7812,N_7621);
nor U10883 (N_10883,N_8938,N_7608);
nand U10884 (N_10884,N_9230,N_5592);
and U10885 (N_10885,N_6405,N_6190);
nor U10886 (N_10886,N_8331,N_7773);
and U10887 (N_10887,N_8146,N_8340);
or U10888 (N_10888,N_8234,N_6455);
and U10889 (N_10889,N_9785,N_6043);
nor U10890 (N_10890,N_6068,N_8688);
nand U10891 (N_10891,N_9124,N_7258);
and U10892 (N_10892,N_8015,N_9778);
and U10893 (N_10893,N_8752,N_6943);
xnor U10894 (N_10894,N_5813,N_7089);
and U10895 (N_10895,N_7380,N_8213);
nor U10896 (N_10896,N_9562,N_9963);
nor U10897 (N_10897,N_8674,N_9734);
nand U10898 (N_10898,N_9925,N_9336);
nand U10899 (N_10899,N_6889,N_7984);
nand U10900 (N_10900,N_5932,N_6503);
and U10901 (N_10901,N_9552,N_7449);
or U10902 (N_10902,N_8789,N_5312);
and U10903 (N_10903,N_6570,N_7317);
nand U10904 (N_10904,N_6517,N_8656);
xor U10905 (N_10905,N_5332,N_7816);
xor U10906 (N_10906,N_7147,N_9430);
and U10907 (N_10907,N_6610,N_8819);
nand U10908 (N_10908,N_6281,N_8296);
and U10909 (N_10909,N_6098,N_6148);
or U10910 (N_10910,N_6136,N_7805);
nand U10911 (N_10911,N_8882,N_8660);
nor U10912 (N_10912,N_9023,N_7482);
xnor U10913 (N_10913,N_5998,N_8447);
and U10914 (N_10914,N_8820,N_5730);
and U10915 (N_10915,N_8090,N_8490);
nand U10916 (N_10916,N_8142,N_7155);
and U10917 (N_10917,N_5456,N_7910);
or U10918 (N_10918,N_5695,N_5712);
nor U10919 (N_10919,N_5726,N_8182);
nor U10920 (N_10920,N_5786,N_6211);
nand U10921 (N_10921,N_6466,N_7326);
or U10922 (N_10922,N_8732,N_7548);
nand U10923 (N_10923,N_7632,N_8141);
nand U10924 (N_10924,N_9965,N_5868);
and U10925 (N_10925,N_7539,N_6957);
nand U10926 (N_10926,N_6030,N_6475);
or U10927 (N_10927,N_9894,N_6080);
or U10928 (N_10928,N_7998,N_7954);
xor U10929 (N_10929,N_7667,N_9803);
or U10930 (N_10930,N_7965,N_8598);
nand U10931 (N_10931,N_6805,N_5600);
xnor U10932 (N_10932,N_8697,N_5210);
or U10933 (N_10933,N_9666,N_7427);
nand U10934 (N_10934,N_6415,N_7346);
nand U10935 (N_10935,N_7059,N_8076);
or U10936 (N_10936,N_6566,N_8506);
xor U10937 (N_10937,N_5483,N_7887);
nand U10938 (N_10938,N_6016,N_9744);
and U10939 (N_10939,N_5875,N_9331);
nand U10940 (N_10940,N_6257,N_5526);
xnor U10941 (N_10941,N_5005,N_6984);
and U10942 (N_10942,N_9989,N_8831);
nor U10943 (N_10943,N_8960,N_9968);
nand U10944 (N_10944,N_9579,N_9601);
xor U10945 (N_10945,N_8241,N_8702);
and U10946 (N_10946,N_8160,N_5963);
nor U10947 (N_10947,N_6733,N_9367);
or U10948 (N_10948,N_5854,N_8791);
or U10949 (N_10949,N_9358,N_6819);
or U10950 (N_10950,N_8240,N_6498);
nand U10951 (N_10951,N_9044,N_9139);
nand U10952 (N_10952,N_7525,N_8969);
xor U10953 (N_10953,N_8238,N_5974);
xnor U10954 (N_10954,N_6843,N_7963);
and U10955 (N_10955,N_6958,N_6327);
nor U10956 (N_10956,N_7366,N_7203);
or U10957 (N_10957,N_9235,N_6644);
and U10958 (N_10958,N_7027,N_6751);
nand U10959 (N_10959,N_5719,N_7231);
or U10960 (N_10960,N_9195,N_8840);
nand U10961 (N_10961,N_7496,N_5785);
nor U10962 (N_10962,N_8392,N_6543);
nor U10963 (N_10963,N_7605,N_9475);
nor U10964 (N_10964,N_7085,N_7645);
or U10965 (N_10965,N_9535,N_5464);
or U10966 (N_10966,N_9871,N_9365);
and U10967 (N_10967,N_9593,N_9733);
nand U10968 (N_10968,N_8465,N_9966);
nor U10969 (N_10969,N_5902,N_8790);
or U10970 (N_10970,N_5842,N_8147);
xor U10971 (N_10971,N_5307,N_7021);
and U10972 (N_10972,N_8483,N_9460);
and U10973 (N_10973,N_6237,N_8721);
nor U10974 (N_10974,N_9742,N_9836);
and U10975 (N_10975,N_8350,N_9582);
nand U10976 (N_10976,N_6867,N_8297);
nor U10977 (N_10977,N_8163,N_7413);
nand U10978 (N_10978,N_9575,N_9498);
nand U10979 (N_10979,N_8488,N_6247);
or U10980 (N_10980,N_9392,N_6817);
xnor U10981 (N_10981,N_8471,N_5219);
nor U10982 (N_10982,N_6854,N_8589);
and U10983 (N_10983,N_7457,N_8454);
nor U10984 (N_10984,N_8782,N_5102);
nor U10985 (N_10985,N_6057,N_7414);
and U10986 (N_10986,N_6615,N_9147);
or U10987 (N_10987,N_8753,N_7935);
and U10988 (N_10988,N_8596,N_5552);
or U10989 (N_10989,N_7121,N_6803);
nor U10990 (N_10990,N_9784,N_9558);
nor U10991 (N_10991,N_6844,N_6738);
nand U10992 (N_10992,N_9753,N_5400);
or U10993 (N_10993,N_8443,N_5166);
xor U10994 (N_10994,N_5128,N_5884);
xor U10995 (N_10995,N_8153,N_5020);
nand U10996 (N_10996,N_6308,N_5942);
xor U10997 (N_10997,N_5356,N_9141);
xor U10998 (N_10998,N_6547,N_9113);
and U10999 (N_10999,N_6291,N_6792);
nor U11000 (N_11000,N_7494,N_6941);
nand U11001 (N_11001,N_7705,N_5349);
xnor U11002 (N_11002,N_9227,N_9397);
nor U11003 (N_11003,N_6700,N_9338);
or U11004 (N_11004,N_5723,N_6419);
nand U11005 (N_11005,N_9929,N_6648);
nor U11006 (N_11006,N_5635,N_5184);
or U11007 (N_11007,N_5891,N_5983);
nand U11008 (N_11008,N_7256,N_7445);
nand U11009 (N_11009,N_8769,N_5652);
nor U11010 (N_11010,N_6879,N_6841);
nor U11011 (N_11011,N_5375,N_9468);
xnor U11012 (N_11012,N_8414,N_8532);
and U11013 (N_11013,N_7504,N_6315);
and U11014 (N_11014,N_7993,N_7242);
xnor U11015 (N_11015,N_8497,N_5100);
nand U11016 (N_11016,N_9334,N_6784);
nand U11017 (N_11017,N_5371,N_8376);
xor U11018 (N_11018,N_6101,N_8750);
nor U11019 (N_11019,N_7635,N_5302);
nand U11020 (N_11020,N_7269,N_8452);
nand U11021 (N_11021,N_5169,N_8030);
nand U11022 (N_11022,N_5441,N_8571);
xnor U11023 (N_11023,N_6815,N_7243);
or U11024 (N_11024,N_6411,N_9992);
xor U11025 (N_11025,N_6444,N_5934);
and U11026 (N_11026,N_8374,N_6096);
or U11027 (N_11027,N_9619,N_7579);
and U11028 (N_11028,N_7080,N_9789);
and U11029 (N_11029,N_5243,N_8543);
nor U11030 (N_11030,N_6706,N_7561);
nand U11031 (N_11031,N_7530,N_7615);
xor U11032 (N_11032,N_8459,N_7594);
nand U11033 (N_11033,N_8661,N_9817);
and U11034 (N_11034,N_8281,N_5909);
or U11035 (N_11035,N_7486,N_5214);
xor U11036 (N_11036,N_7343,N_9176);
and U11037 (N_11037,N_6334,N_8441);
xnor U11038 (N_11038,N_6736,N_6749);
nand U11039 (N_11039,N_7492,N_8701);
or U11040 (N_11040,N_5281,N_6693);
and U11041 (N_11041,N_8007,N_6699);
xnor U11042 (N_11042,N_8103,N_9667);
and U11043 (N_11043,N_7629,N_7487);
or U11044 (N_11044,N_6951,N_8239);
or U11045 (N_11045,N_7753,N_7503);
nor U11046 (N_11046,N_7881,N_7702);
or U11047 (N_11047,N_7850,N_8622);
nand U11048 (N_11048,N_6723,N_5810);
nor U11049 (N_11049,N_8021,N_7552);
or U11050 (N_11050,N_8680,N_9501);
xnor U11051 (N_11051,N_7933,N_9745);
nor U11052 (N_11052,N_6003,N_9401);
or U11053 (N_11053,N_9986,N_9343);
xor U11054 (N_11054,N_9096,N_9449);
nand U11055 (N_11055,N_9347,N_5450);
and U11056 (N_11056,N_8425,N_7493);
or U11057 (N_11057,N_9885,N_9129);
or U11058 (N_11058,N_5808,N_8446);
and U11059 (N_11059,N_5297,N_8777);
nor U11060 (N_11060,N_9765,N_5176);
and U11061 (N_11061,N_8148,N_8046);
and U11062 (N_11062,N_5618,N_9839);
nor U11063 (N_11063,N_9505,N_6326);
nand U11064 (N_11064,N_8915,N_9780);
or U11065 (N_11065,N_7633,N_6061);
nand U11066 (N_11066,N_9922,N_6200);
xor U11067 (N_11067,N_5134,N_5175);
nor U11068 (N_11068,N_8594,N_7463);
xnor U11069 (N_11069,N_6418,N_7285);
or U11070 (N_11070,N_5193,N_9541);
nand U11071 (N_11071,N_7455,N_7838);
or U11072 (N_11072,N_8288,N_6259);
or U11073 (N_11073,N_6062,N_6295);
xor U11074 (N_11074,N_8898,N_6538);
nor U11075 (N_11075,N_9463,N_8797);
xor U11076 (N_11076,N_5831,N_9834);
and U11077 (N_11077,N_8051,N_9623);
xnor U11078 (N_11078,N_8041,N_6505);
xnor U11079 (N_11079,N_7105,N_8428);
xnor U11080 (N_11080,N_9398,N_7922);
xnor U11081 (N_11081,N_6018,N_7700);
or U11082 (N_11082,N_7362,N_5528);
and U11083 (N_11083,N_6629,N_9342);
and U11084 (N_11084,N_5563,N_5523);
and U11085 (N_11085,N_8386,N_9030);
xor U11086 (N_11086,N_5088,N_5770);
nor U11087 (N_11087,N_7518,N_5061);
xor U11088 (N_11088,N_8473,N_7431);
and U11089 (N_11089,N_9352,N_6924);
or U11090 (N_11090,N_7693,N_7654);
nor U11091 (N_11091,N_8572,N_5877);
nand U11092 (N_11092,N_7669,N_7319);
and U11093 (N_11093,N_9993,N_5072);
or U11094 (N_11094,N_8294,N_8841);
or U11095 (N_11095,N_5394,N_9847);
nand U11096 (N_11096,N_5323,N_9647);
or U11097 (N_11097,N_6856,N_9751);
xor U11098 (N_11098,N_6556,N_8125);
nor U11099 (N_11099,N_7044,N_7739);
and U11100 (N_11100,N_9181,N_5780);
nand U11101 (N_11101,N_9912,N_8629);
nor U11102 (N_11102,N_5665,N_5702);
nand U11103 (N_11103,N_6524,N_6822);
nand U11104 (N_11104,N_8303,N_7514);
nand U11105 (N_11105,N_6935,N_6776);
nor U11106 (N_11106,N_9730,N_6137);
or U11107 (N_11107,N_7688,N_7416);
nor U11108 (N_11108,N_8403,N_7464);
xor U11109 (N_11109,N_9643,N_6863);
xor U11110 (N_11110,N_5171,N_6354);
xor U11111 (N_11111,N_5163,N_5123);
xnor U11112 (N_11112,N_9236,N_6476);
and U11113 (N_11113,N_6058,N_9930);
nor U11114 (N_11114,N_5581,N_7033);
xnor U11115 (N_11115,N_6420,N_9684);
nand U11116 (N_11116,N_5988,N_5130);
nor U11117 (N_11117,N_9489,N_5295);
or U11118 (N_11118,N_7505,N_9957);
nor U11119 (N_11119,N_5025,N_7298);
xor U11120 (N_11120,N_5403,N_7277);
xor U11121 (N_11121,N_5796,N_6692);
nor U11122 (N_11122,N_6350,N_6651);
nand U11123 (N_11123,N_8073,N_9843);
xor U11124 (N_11124,N_7485,N_9212);
xor U11125 (N_11125,N_8946,N_9219);
xor U11126 (N_11126,N_7095,N_8430);
nand U11127 (N_11127,N_5138,N_8244);
xnor U11128 (N_11128,N_9353,N_8972);
xor U11129 (N_11129,N_7977,N_8276);
nand U11130 (N_11130,N_5613,N_9414);
xor U11131 (N_11131,N_6140,N_5182);
xnor U11132 (N_11132,N_8838,N_7122);
nand U11133 (N_11133,N_9419,N_9842);
or U11134 (N_11134,N_9411,N_6465);
nor U11135 (N_11135,N_8519,N_6714);
nand U11136 (N_11136,N_6497,N_9783);
or U11137 (N_11137,N_9769,N_9491);
xor U11138 (N_11138,N_9774,N_5987);
nor U11139 (N_11139,N_8955,N_6424);
and U11140 (N_11140,N_8196,N_9412);
nor U11141 (N_11141,N_8282,N_5869);
nor U11142 (N_11142,N_9849,N_6763);
and U11143 (N_11143,N_5024,N_8436);
nand U11144 (N_11144,N_7768,N_9875);
nor U11145 (N_11145,N_8647,N_5197);
nand U11146 (N_11146,N_9481,N_7536);
nor U11147 (N_11147,N_8469,N_5633);
nand U11148 (N_11148,N_5584,N_8758);
nand U11149 (N_11149,N_6277,N_6952);
and U11150 (N_11150,N_9242,N_6428);
or U11151 (N_11151,N_7152,N_8460);
or U11152 (N_11152,N_9779,N_7558);
xor U11153 (N_11153,N_5579,N_7061);
or U11154 (N_11154,N_5622,N_6956);
or U11155 (N_11155,N_8491,N_7409);
xor U11156 (N_11156,N_8763,N_5834);
nor U11157 (N_11157,N_8061,N_5132);
and U11158 (N_11158,N_8783,N_5502);
xor U11159 (N_11159,N_5850,N_6611);
and U11160 (N_11160,N_9402,N_6551);
nor U11161 (N_11161,N_5415,N_6103);
or U11162 (N_11162,N_6892,N_9545);
nor U11163 (N_11163,N_7190,N_7118);
nor U11164 (N_11164,N_8264,N_9072);
nand U11165 (N_11165,N_9650,N_7253);
xor U11166 (N_11166,N_8518,N_9313);
or U11167 (N_11167,N_7312,N_8233);
and U11168 (N_11168,N_5440,N_7906);
nand U11169 (N_11169,N_9387,N_6519);
or U11170 (N_11170,N_6625,N_7406);
or U11171 (N_11171,N_5428,N_7640);
or U11172 (N_11172,N_6242,N_6818);
and U11173 (N_11173,N_8121,N_9074);
nor U11174 (N_11174,N_7528,N_7411);
nand U11175 (N_11175,N_8931,N_9796);
and U11176 (N_11176,N_9100,N_7546);
and U11177 (N_11177,N_5315,N_6125);
xnor U11178 (N_11178,N_6782,N_9564);
nor U11179 (N_11179,N_7067,N_7631);
nor U11180 (N_11180,N_9969,N_7861);
nor U11181 (N_11181,N_6040,N_9289);
xnor U11182 (N_11182,N_8974,N_5949);
nor U11183 (N_11183,N_5864,N_5593);
nor U11184 (N_11184,N_7836,N_9059);
nor U11185 (N_11185,N_5647,N_9644);
xor U11186 (N_11186,N_8850,N_9981);
and U11187 (N_11187,N_5783,N_6020);
xor U11188 (N_11188,N_9479,N_9611);
nand U11189 (N_11189,N_6913,N_9758);
nand U11190 (N_11190,N_7624,N_5690);
or U11191 (N_11191,N_7351,N_8225);
and U11192 (N_11192,N_5475,N_8237);
nor U11193 (N_11193,N_8968,N_6399);
xnor U11194 (N_11194,N_7092,N_8366);
nand U11195 (N_11195,N_8462,N_9228);
nor U11196 (N_11196,N_7859,N_9852);
nor U11197 (N_11197,N_6276,N_9448);
and U11198 (N_11198,N_9094,N_5805);
nor U11199 (N_11199,N_6676,N_8720);
nor U11200 (N_11200,N_7215,N_7828);
or U11201 (N_11201,N_7619,N_5048);
xnor U11202 (N_11202,N_9004,N_9193);
xor U11203 (N_11203,N_5557,N_7476);
xor U11204 (N_11204,N_5503,N_8388);
nor U11205 (N_11205,N_8256,N_6546);
xnor U11206 (N_11206,N_8638,N_6773);
or U11207 (N_11207,N_6983,N_5731);
and U11208 (N_11208,N_5073,N_5640);
or U11209 (N_11209,N_7927,N_5738);
and U11210 (N_11210,N_7897,N_9291);
and U11211 (N_11211,N_8726,N_8879);
nor U11212 (N_11212,N_6300,N_8856);
xnor U11213 (N_11213,N_5331,N_8567);
nand U11214 (N_11214,N_8074,N_7246);
and U11215 (N_11215,N_7789,N_9618);
xor U11216 (N_11216,N_9202,N_6318);
and U11217 (N_11217,N_7959,N_8224);
nor U11218 (N_11218,N_5765,N_6813);
xor U11219 (N_11219,N_5682,N_5732);
nand U11220 (N_11220,N_6916,N_5931);
or U11221 (N_11221,N_6724,N_7610);
or U11222 (N_11222,N_9577,N_8255);
or U11223 (N_11223,N_9747,N_6781);
nor U11224 (N_11224,N_5249,N_7167);
and U11225 (N_11225,N_7161,N_5028);
nand U11226 (N_11226,N_9899,N_8489);
xnor U11227 (N_11227,N_8967,N_6355);
xnor U11228 (N_11228,N_9086,N_8361);
nand U11229 (N_11229,N_9252,N_7254);
xor U11230 (N_11230,N_7827,N_6426);
nand U11231 (N_11231,N_7153,N_7834);
nor U11232 (N_11232,N_5925,N_9821);
and U11233 (N_11233,N_5369,N_7745);
nor U11234 (N_11234,N_8597,N_9022);
nor U11235 (N_11235,N_6799,N_5257);
xnor U11236 (N_11236,N_6370,N_6667);
nor U11237 (N_11237,N_6520,N_5560);
xnor U11238 (N_11238,N_7117,N_9079);
xnor U11239 (N_11239,N_5453,N_5057);
xnor U11240 (N_11240,N_7800,N_5390);
nand U11241 (N_11241,N_5108,N_5589);
nor U11242 (N_11242,N_7437,N_6507);
or U11243 (N_11243,N_7031,N_5230);
and U11244 (N_11244,N_6450,N_7310);
xor U11245 (N_11245,N_8810,N_7973);
and U11246 (N_11246,N_9098,N_6111);
or U11247 (N_11247,N_9997,N_8650);
xnor U11248 (N_11248,N_9844,N_5253);
and U11249 (N_11249,N_6632,N_8734);
or U11250 (N_11250,N_6554,N_7858);
or U11251 (N_11251,N_6869,N_5344);
nor U11252 (N_11252,N_9500,N_9337);
nand U11253 (N_11253,N_8665,N_5901);
and U11254 (N_11254,N_7884,N_5585);
and U11255 (N_11255,N_7990,N_6033);
or U11256 (N_11256,N_7304,N_5945);
nor U11257 (N_11257,N_5135,N_5746);
nor U11258 (N_11258,N_6933,N_9982);
nand U11259 (N_11259,N_8905,N_6734);
nor U11260 (N_11260,N_7129,N_8435);
and U11261 (N_11261,N_8458,N_9470);
and U11262 (N_11262,N_9790,N_6797);
nor U11263 (N_11263,N_5713,N_8526);
nor U11264 (N_11264,N_9933,N_6204);
nand U11265 (N_11265,N_5539,N_8470);
xor U11266 (N_11266,N_7535,N_7309);
xnor U11267 (N_11267,N_9344,N_7921);
or U11268 (N_11268,N_5751,N_5454);
and U11269 (N_11269,N_8180,N_5296);
or U11270 (N_11270,N_6171,N_6329);
xor U11271 (N_11271,N_8862,N_6179);
xor U11272 (N_11272,N_7441,N_5521);
nand U11273 (N_11273,N_8143,N_9440);
or U11274 (N_11274,N_6481,N_9687);
xor U11275 (N_11275,N_7646,N_8042);
xnor U11276 (N_11276,N_7425,N_7521);
nor U11277 (N_11277,N_6464,N_5708);
xnor U11278 (N_11278,N_5052,N_9608);
nor U11279 (N_11279,N_8221,N_6988);
and U11280 (N_11280,N_8947,N_8100);
xor U11281 (N_11281,N_9167,N_8576);
or U11282 (N_11282,N_9736,N_6263);
and U11283 (N_11283,N_7815,N_5105);
nand U11284 (N_11284,N_5757,N_8553);
xor U11285 (N_11285,N_8315,N_8026);
nor U11286 (N_11286,N_6236,N_7007);
nand U11287 (N_11287,N_9514,N_9767);
and U11288 (N_11288,N_6544,N_7710);
and U11289 (N_11289,N_5907,N_6485);
or U11290 (N_11290,N_5421,N_5457);
or U11291 (N_11291,N_5248,N_9657);
and U11292 (N_11292,N_5154,N_8070);
nor U11293 (N_11293,N_8505,N_8768);
nor U11294 (N_11294,N_6064,N_9407);
xor U11295 (N_11295,N_9559,N_6912);
nand U11296 (N_11296,N_7149,N_5614);
nand U11297 (N_11297,N_6874,N_8191);
nand U11298 (N_11298,N_8952,N_8716);
and U11299 (N_11299,N_9916,N_7666);
nand U11300 (N_11300,N_8265,N_8866);
or U11301 (N_11301,N_8541,N_5468);
xnor U11302 (N_11302,N_7189,N_7656);
xor U11303 (N_11303,N_6540,N_8895);
and U11304 (N_11304,N_6286,N_8900);
or U11305 (N_11305,N_5848,N_6198);
nor U11306 (N_11306,N_6027,N_9065);
nand U11307 (N_11307,N_8934,N_9025);
xor U11308 (N_11308,N_5114,N_5038);
and U11309 (N_11309,N_6786,N_8209);
nor U11310 (N_11310,N_5943,N_9757);
and U11311 (N_11311,N_8092,N_5542);
and U11312 (N_11312,N_8018,N_8308);
nand U11313 (N_11313,N_7218,N_6159);
xor U11314 (N_11314,N_6440,N_9697);
nand U11315 (N_11315,N_8685,N_7687);
nor U11316 (N_11316,N_8293,N_7781);
nor U11317 (N_11317,N_6022,N_8982);
and U11318 (N_11318,N_8014,N_5681);
or U11319 (N_11319,N_7133,N_9883);
xor U11320 (N_11320,N_6127,N_6939);
xnor U11321 (N_11321,N_8252,N_8068);
or U11322 (N_11322,N_7172,N_8996);
and U11323 (N_11323,N_9027,N_8586);
or U11324 (N_11324,N_9029,N_5717);
and U11325 (N_11325,N_6765,N_5709);
and U11326 (N_11326,N_8463,N_5718);
and U11327 (N_11327,N_6317,N_5327);
xor U11328 (N_11328,N_7999,N_9263);
and U11329 (N_11329,N_8635,N_8063);
nor U11330 (N_11330,N_7641,N_6292);
nand U11331 (N_11331,N_9013,N_5146);
or U11332 (N_11332,N_9052,N_6332);
and U11333 (N_11333,N_7315,N_8493);
nor U11334 (N_11334,N_6655,N_9788);
nand U11335 (N_11335,N_6266,N_5800);
nor U11336 (N_11336,N_7348,N_7517);
nor U11337 (N_11337,N_9863,N_5432);
nor U11338 (N_11338,N_8605,N_5264);
nand U11339 (N_11339,N_6682,N_5091);
nor U11340 (N_11340,N_8322,N_5121);
nand U11341 (N_11341,N_6208,N_8902);
or U11342 (N_11342,N_6650,N_9490);
nor U11343 (N_11343,N_6182,N_5823);
nand U11344 (N_11344,N_8135,N_6596);
and U11345 (N_11345,N_5653,N_6393);
nor U11346 (N_11346,N_8501,N_9198);
or U11347 (N_11347,N_7156,N_9009);
and U11348 (N_11348,N_6895,N_6937);
nor U11349 (N_11349,N_6529,N_7676);
nand U11350 (N_11350,N_9642,N_6851);
nor U11351 (N_11351,N_5085,N_7932);
nor U11352 (N_11352,N_5271,N_9329);
xor U11353 (N_11353,N_6639,N_9527);
and U11354 (N_11354,N_9874,N_8169);
xnor U11355 (N_11355,N_8438,N_9140);
nand U11356 (N_11356,N_7501,N_9437);
nor U11357 (N_11357,N_7313,N_8464);
and U11358 (N_11358,N_5016,N_7327);
nor U11359 (N_11359,N_5606,N_7069);
nor U11360 (N_11360,N_9637,N_7112);
nand U11361 (N_11361,N_6783,N_7627);
nand U11362 (N_11362,N_5272,N_7397);
xnor U11363 (N_11363,N_6590,N_7576);
nand U11364 (N_11364,N_6849,N_6233);
nand U11365 (N_11365,N_7516,N_6954);
xor U11366 (N_11366,N_6240,N_5452);
and U11367 (N_11367,N_9264,N_7930);
nor U11368 (N_11368,N_9319,N_7474);
and U11369 (N_11369,N_9066,N_8551);
xor U11370 (N_11370,N_7983,N_8880);
nand U11371 (N_11371,N_6828,N_6891);
or U11372 (N_11372,N_8704,N_7048);
and U11373 (N_11373,N_8926,N_8207);
or U11374 (N_11374,N_5889,N_6698);
nand U11375 (N_11375,N_7987,N_7096);
and U11376 (N_11376,N_6523,N_5861);
or U11377 (N_11377,N_6014,N_5050);
nor U11378 (N_11378,N_6953,N_8305);
or U11379 (N_11379,N_9537,N_5616);
and U11380 (N_11380,N_8140,N_5720);
or U11381 (N_11381,N_5212,N_7020);
nand U11382 (N_11382,N_8310,N_7975);
nor U11383 (N_11383,N_6304,N_7259);
nand U11384 (N_11384,N_5703,N_8738);
or U11385 (N_11385,N_8319,N_5865);
or U11386 (N_11386,N_6760,N_6661);
nor U11387 (N_11387,N_5858,N_8772);
nand U11388 (N_11388,N_9378,N_7911);
xor U11389 (N_11389,N_7764,N_8295);
and U11390 (N_11390,N_8662,N_7316);
nand U11391 (N_11391,N_8082,N_5040);
and U11392 (N_11392,N_7334,N_7134);
nand U11393 (N_11393,N_7045,N_9199);
nand U11394 (N_11394,N_9661,N_8653);
nor U11395 (N_11395,N_8056,N_7195);
or U11396 (N_11396,N_6755,N_5333);
nor U11397 (N_11397,N_5993,N_7783);
xnor U11398 (N_11398,N_5148,N_6007);
nor U11399 (N_11399,N_9792,N_5820);
and U11400 (N_11400,N_5113,N_8139);
and U11401 (N_11401,N_9974,N_6166);
nand U11402 (N_11402,N_9621,N_6219);
nand U11403 (N_11403,N_5968,N_7659);
nand U11404 (N_11404,N_6896,N_5973);
xnor U11405 (N_11405,N_6110,N_9224);
or U11406 (N_11406,N_9312,N_9731);
xor U11407 (N_11407,N_9512,N_9274);
or U11408 (N_11408,N_9987,N_5887);
and U11409 (N_11409,N_8844,N_9482);
or U11410 (N_11410,N_9620,N_7685);
nand U11411 (N_11411,N_5000,N_8301);
nand U11412 (N_11412,N_5275,N_8914);
and U11413 (N_11413,N_5078,N_6572);
nand U11414 (N_11414,N_7379,N_9598);
or U11415 (N_11415,N_9880,N_9409);
nand U11416 (N_11416,N_9893,N_6146);
nand U11417 (N_11417,N_6825,N_6462);
nor U11418 (N_11418,N_9048,N_8659);
xor U11419 (N_11419,N_6454,N_8671);
nand U11420 (N_11420,N_9131,N_9828);
or U11421 (N_11421,N_9260,N_7864);
nor U11422 (N_11422,N_7140,N_9335);
nor U11423 (N_11423,N_5179,N_7005);
nand U11424 (N_11424,N_6126,N_6764);
and U11425 (N_11425,N_6480,N_9496);
and U11426 (N_11426,N_5790,N_9578);
or U11427 (N_11427,N_7958,N_5802);
or U11428 (N_11428,N_5990,N_7201);
and U11429 (N_11429,N_8400,N_6037);
and U11430 (N_11430,N_6771,N_9099);
nand U11431 (N_11431,N_8038,N_9047);
or U11432 (N_11432,N_7611,N_7988);
or U11433 (N_11433,N_9638,N_7356);
xor U11434 (N_11434,N_6067,N_5306);
and U11435 (N_11435,N_8467,N_9776);
nor U11436 (N_11436,N_7018,N_6307);
or U11437 (N_11437,N_6028,N_6996);
xor U11438 (N_11438,N_5044,N_7593);
nand U11439 (N_11439,N_8445,N_6174);
nand U11440 (N_11440,N_5871,N_5583);
xor U11441 (N_11441,N_9532,N_5832);
and U11442 (N_11442,N_5446,N_8152);
and U11443 (N_11443,N_9786,N_7391);
nand U11444 (N_11444,N_9268,N_7433);
xor U11445 (N_11445,N_8869,N_8904);
nand U11446 (N_11446,N_9805,N_5039);
or U11447 (N_11447,N_5259,N_5894);
nand U11448 (N_11448,N_9218,N_6787);
nand U11449 (N_11449,N_8778,N_8280);
nor U11450 (N_11450,N_5511,N_5675);
xor U11451 (N_11451,N_7209,N_5354);
nand U11452 (N_11452,N_5912,N_5941);
xor U11453 (N_11453,N_6995,N_8907);
and U11454 (N_11454,N_8150,N_9375);
nor U11455 (N_11455,N_7950,N_7374);
xnor U11456 (N_11456,N_7568,N_9715);
xor U11457 (N_11457,N_6135,N_5204);
or U11458 (N_11458,N_6060,N_7257);
or U11459 (N_11459,N_7079,N_8179);
nand U11460 (N_11460,N_8009,N_8524);
and U11461 (N_11461,N_5985,N_9070);
and U11462 (N_11462,N_8020,N_5844);
and U11463 (N_11463,N_5092,N_5648);
and U11464 (N_11464,N_8187,N_6184);
and U11465 (N_11465,N_9245,N_6104);
nor U11466 (N_11466,N_9318,N_7125);
nor U11467 (N_11467,N_6689,N_7814);
xnor U11468 (N_11468,N_6201,N_5455);
and U11469 (N_11469,N_6479,N_9886);
xor U11470 (N_11470,N_7714,N_5298);
nand U11471 (N_11471,N_6076,N_8235);
nand U11472 (N_11472,N_7956,N_8115);
or U11473 (N_11473,N_6088,N_9019);
or U11474 (N_11474,N_5387,N_6574);
or U11475 (N_11475,N_7456,N_7630);
nand U11476 (N_11476,N_8675,N_7502);
and U11477 (N_11477,N_8286,N_6388);
xnor U11478 (N_11478,N_5781,N_9275);
nand U11479 (N_11479,N_7039,N_9102);
or U11480 (N_11480,N_8612,N_7636);
and U11481 (N_11481,N_7898,N_5326);
xnor U11482 (N_11482,N_6664,N_7373);
and U11483 (N_11483,N_7955,N_5215);
and U11484 (N_11484,N_8845,N_6845);
xnor U11485 (N_11485,N_9936,N_8705);
or U11486 (N_11486,N_9039,N_6187);
nor U11487 (N_11487,N_5222,N_6108);
or U11488 (N_11488,N_6910,N_7541);
xnor U11489 (N_11489,N_9746,N_9097);
xor U11490 (N_11490,N_6116,N_8607);
or U11491 (N_11491,N_6168,N_8577);
or U11492 (N_11492,N_5601,N_6273);
and U11493 (N_11493,N_9346,N_6816);
or U11494 (N_11494,N_9403,N_7028);
and U11495 (N_11495,N_5911,N_8746);
xor U11496 (N_11496,N_9361,N_5897);
and U11497 (N_11497,N_5300,N_9587);
and U11498 (N_11498,N_9528,N_6963);
xnor U11499 (N_11499,N_7245,N_6172);
nor U11500 (N_11500,N_8950,N_6934);
or U11501 (N_11501,N_5436,N_5855);
and U11502 (N_11502,N_8533,N_9115);
xnor U11503 (N_11503,N_9201,N_6134);
xnor U11504 (N_11504,N_6287,N_5481);
and U11505 (N_11505,N_9156,N_8172);
xor U11506 (N_11506,N_9016,N_9213);
nand U11507 (N_11507,N_9851,N_6193);
nand U11508 (N_11508,N_9309,N_8289);
and U11509 (N_11509,N_7419,N_9076);
nor U11510 (N_11510,N_7584,N_7829);
or U11511 (N_11511,N_5975,N_6670);
or U11512 (N_11512,N_7655,N_8243);
and U11513 (N_11513,N_6746,N_7775);
xor U11514 (N_11514,N_9297,N_7506);
xor U11515 (N_11515,N_6448,N_6752);
xor U11516 (N_11516,N_6850,N_9688);
nand U11517 (N_11517,N_7680,N_8314);
nand U11518 (N_11518,N_9740,N_5721);
or U11519 (N_11519,N_8218,N_6852);
xnor U11520 (N_11520,N_6753,N_5374);
xnor U11521 (N_11521,N_8615,N_9315);
or U11522 (N_11522,N_5157,N_6515);
nor U11523 (N_11523,N_8468,N_9939);
nand U11524 (N_11524,N_6717,N_7712);
nor U11525 (N_11525,N_9492,N_7429);
or U11526 (N_11526,N_6525,N_6735);
xnor U11527 (N_11527,N_8277,N_5282);
and U11528 (N_11528,N_9142,N_9955);
xor U11529 (N_11529,N_8585,N_7696);
nand U11530 (N_11530,N_9207,N_5220);
nor U11531 (N_11531,N_9566,N_9011);
nand U11532 (N_11532,N_6337,N_7142);
and U11533 (N_11533,N_6396,N_9652);
xnor U11534 (N_11534,N_6290,N_8086);
and U11535 (N_11535,N_6099,N_6695);
or U11536 (N_11536,N_5301,N_6986);
xnor U11537 (N_11537,N_7219,N_8978);
nor U11538 (N_11538,N_6443,N_6837);
xnor U11539 (N_11539,N_7192,N_5318);
or U11540 (N_11540,N_8094,N_5903);
nand U11541 (N_11541,N_5649,N_9606);
or U11542 (N_11542,N_7574,N_6157);
or U11543 (N_11543,N_7681,N_5915);
and U11544 (N_11544,N_8614,N_5664);
xor U11545 (N_11545,N_5396,N_6599);
nand U11546 (N_11546,N_8382,N_5632);
or U11547 (N_11547,N_5967,N_7526);
nand U11548 (N_11548,N_6390,N_8298);
and U11549 (N_11549,N_8183,N_9738);
or U11550 (N_11550,N_6638,N_7691);
and U11551 (N_11551,N_8195,N_5971);
and U11552 (N_11552,N_8089,N_9474);
nor U11553 (N_11553,N_8409,N_7015);
xor U11554 (N_11554,N_7644,N_8917);
xor U11555 (N_11555,N_5654,N_9443);
xnor U11556 (N_11556,N_5811,N_8365);
or U11557 (N_11557,N_9307,N_5669);
xor U11558 (N_11558,N_9133,N_7148);
nor U11559 (N_11559,N_8411,N_8728);
xnor U11560 (N_11560,N_5896,N_9944);
and U11561 (N_11561,N_9553,N_5147);
and U11562 (N_11562,N_7143,N_6260);
nand U11563 (N_11563,N_5002,N_7925);
and U11564 (N_11564,N_6908,N_6688);
nor U11565 (N_11565,N_9155,N_6591);
nor U11566 (N_11566,N_7592,N_5691);
nor U11567 (N_11567,N_7844,N_9680);
nor U11568 (N_11568,N_9651,N_8751);
and U11569 (N_11569,N_7766,N_8574);
nor U11570 (N_11570,N_8935,N_5917);
nand U11571 (N_11571,N_5947,N_9557);
xor U11572 (N_11572,N_7797,N_5190);
or U11573 (N_11573,N_7307,N_8641);
nand U11574 (N_11574,N_6423,N_8802);
nand U11575 (N_11575,N_8356,N_6619);
nor U11576 (N_11576,N_8204,N_6766);
or U11577 (N_11577,N_6066,N_8208);
xor U11578 (N_11578,N_7126,N_7038);
nand U11579 (N_11579,N_7649,N_6152);
nor U11580 (N_11580,N_5544,N_5969);
nand U11581 (N_11581,N_5238,N_9787);
nor U11582 (N_11582,N_9241,N_8736);
and U11583 (N_11583,N_7737,N_6681);
or U11584 (N_11584,N_5386,N_5919);
xnor U11585 (N_11585,N_6569,N_5522);
xnor U11586 (N_11586,N_9991,N_8313);
xnor U11587 (N_11587,N_6353,N_7452);
or U11588 (N_11588,N_8516,N_8081);
xnor U11589 (N_11589,N_5270,N_9283);
xnor U11590 (N_11590,N_9629,N_9020);
nor U11591 (N_11591,N_9453,N_6160);
xnor U11592 (N_11592,N_6213,N_8549);
xnor U11593 (N_11593,N_6607,N_9413);
nor U11594 (N_11594,N_7626,N_9194);
xor U11595 (N_11595,N_9149,N_5256);
nand U11596 (N_11596,N_8587,N_7763);
or U11597 (N_11597,N_5615,N_7444);
xor U11598 (N_11598,N_9217,N_8112);
nand U11599 (N_11599,N_6346,N_6272);
or U11600 (N_11600,N_7043,N_6232);
or U11601 (N_11601,N_6711,N_7055);
xnor U11602 (N_11602,N_5795,N_9210);
or U11603 (N_11603,N_9533,N_5293);
nand U11604 (N_11604,N_9722,N_6555);
and U11605 (N_11605,N_7750,N_8166);
nand U11606 (N_11606,N_6721,N_7830);
nand U11607 (N_11607,N_5355,N_5265);
xor U11608 (N_11608,N_9385,N_7531);
xor U11609 (N_11609,N_7477,N_5970);
or U11610 (N_11610,N_8901,N_6407);
nor U11611 (N_11611,N_5338,N_7601);
or U11612 (N_11612,N_6417,N_7616);
and U11613 (N_11613,N_6362,N_8961);
nand U11614 (N_11614,N_7470,N_8258);
nor U11615 (N_11615,N_7357,N_6907);
and U11616 (N_11616,N_5905,N_8118);
nor U11617 (N_11617,N_5358,N_8677);
and U11618 (N_11618,N_9499,N_9442);
and U11619 (N_11619,N_6191,N_5030);
and U11620 (N_11620,N_6904,N_6853);
and U11621 (N_11621,N_9143,N_9243);
or U11622 (N_11622,N_6936,N_5602);
nor U11623 (N_11623,N_8620,N_7665);
and U11624 (N_11624,N_8418,N_9855);
nor U11625 (N_11625,N_9700,N_9249);
or U11626 (N_11626,N_5063,N_7012);
or U11627 (N_11627,N_5119,N_9373);
xnor U11628 (N_11628,N_9822,N_9690);
nand U11629 (N_11629,N_6071,N_5621);
nand U11630 (N_11630,N_9797,N_9902);
nand U11631 (N_11631,N_5596,N_5628);
nor U11632 (N_11632,N_7178,N_7271);
nand U11633 (N_11633,N_9913,N_8779);
nor U11634 (N_11634,N_8145,N_9878);
nand U11635 (N_11635,N_8785,N_6606);
xnor U11636 (N_11636,N_8722,N_9146);
nor U11637 (N_11637,N_6987,N_6079);
or U11638 (N_11638,N_7066,N_5097);
nor U11639 (N_11639,N_6031,N_5494);
nand U11640 (N_11640,N_7623,N_6737);
nand U11641 (N_11641,N_5395,N_8874);
or U11642 (N_11642,N_6421,N_8694);
or U11643 (N_11643,N_7338,N_6571);
or U11644 (N_11644,N_8226,N_7826);
xnor U11645 (N_11645,N_9905,N_9701);
or U11646 (N_11646,N_6439,N_6074);
nand U11647 (N_11647,N_5180,N_6834);
xnor U11648 (N_11648,N_9121,N_9571);
nor U11649 (N_11649,N_8932,N_9749);
nand U11650 (N_11650,N_6177,N_8171);
nor U11651 (N_11651,N_9189,N_8787);
xnor U11652 (N_11652,N_7214,N_7713);
xor U11653 (N_11653,N_6756,N_5448);
nand U11654 (N_11654,N_5381,N_5910);
or U11655 (N_11655,N_6550,N_6830);
xor U11656 (N_11656,N_6199,N_8883);
and U11657 (N_11657,N_5167,N_9258);
or U11658 (N_11658,N_7384,N_5761);
and U11659 (N_11659,N_5749,N_5324);
or U11660 (N_11660,N_8072,N_8708);
nand U11661 (N_11661,N_5066,N_6905);
or U11662 (N_11662,N_5240,N_7729);
or U11663 (N_11663,N_6385,N_9308);
xnor U11664 (N_11664,N_8648,N_9324);
xor U11665 (N_11665,N_8149,N_8050);
or U11666 (N_11666,N_8367,N_6378);
nand U11667 (N_11667,N_5277,N_5747);
and U11668 (N_11668,N_9056,N_9031);
xor U11669 (N_11669,N_6970,N_6533);
and U11670 (N_11670,N_9756,N_8096);
and U11671 (N_11671,N_6445,N_5422);
and U11672 (N_11672,N_7617,N_6349);
nand U11673 (N_11673,N_8527,N_8329);
or U11674 (N_11674,N_8312,N_6483);
nand U11675 (N_11675,N_9949,N_9594);
and U11676 (N_11676,N_7041,N_7436);
or U11677 (N_11677,N_8004,N_6718);
nand U11678 (N_11678,N_7369,N_5995);
xor U11679 (N_11679,N_6653,N_5026);
nor U11680 (N_11680,N_8817,N_6401);
nor U11681 (N_11681,N_9286,N_7076);
nand U11682 (N_11682,N_7400,N_8534);
xor U11683 (N_11683,N_6487,N_7883);
nor U11684 (N_11684,N_9860,N_8712);
and U11685 (N_11685,N_8410,N_6573);
xnor U11686 (N_11686,N_7698,N_6036);
nor U11687 (N_11687,N_6582,N_6578);
xor U11688 (N_11688,N_8835,N_5279);
nor U11689 (N_11689,N_5906,N_7770);
nand U11690 (N_11690,N_7168,N_8378);
nand U11691 (N_11691,N_8377,N_9591);
nor U11692 (N_11692,N_8251,N_5047);
or U11693 (N_11693,N_6709,N_6793);
xor U11694 (N_11694,N_8230,N_7878);
xor U11695 (N_11695,N_9685,N_7154);
and U11696 (N_11696,N_5812,N_6703);
or U11697 (N_11697,N_7480,N_8138);
or U11698 (N_11698,N_8803,N_5627);
and U11699 (N_11699,N_5556,N_5304);
nor U11700 (N_11700,N_7070,N_5314);
or U11701 (N_11701,N_7658,N_5568);
and U11702 (N_11702,N_5984,N_9943);
and U11703 (N_11703,N_5899,N_9762);
and U11704 (N_11704,N_9325,N_9034);
or U11705 (N_11705,N_7146,N_5493);
xnor U11706 (N_11706,N_9111,N_9810);
xnor U11707 (N_11707,N_7603,N_8565);
or U11708 (N_11708,N_9266,N_6158);
xnor U11709 (N_11709,N_8002,N_7512);
and U11710 (N_11710,N_5347,N_9818);
nand U11711 (N_11711,N_6050,N_6785);
xnor U11712 (N_11712,N_9368,N_6119);
nand U11713 (N_11713,N_6535,N_7248);
nand U11714 (N_11714,N_5467,N_9068);
and U11715 (N_11715,N_8087,N_8964);
or U11716 (N_11716,N_8099,N_7527);
nand U11717 (N_11717,N_6739,N_6324);
or U11718 (N_11718,N_9895,N_9357);
or U11719 (N_11719,N_9935,N_9417);
nor U11720 (N_11720,N_7207,N_9820);
nand U11721 (N_11721,N_5603,N_9511);
and U11722 (N_11722,N_5890,N_6894);
nor U11723 (N_11723,N_5948,N_7866);
or U11724 (N_11724,N_9602,N_6810);
xor U11725 (N_11725,N_9485,N_5133);
xor U11726 (N_11726,N_8034,N_8892);
and U11727 (N_11727,N_8645,N_7668);
nand U11728 (N_11728,N_7695,N_6848);
xor U11729 (N_11729,N_6900,N_7128);
and U11730 (N_11730,N_5376,N_7780);
or U11731 (N_11731,N_8116,N_9962);
nor U11732 (N_11732,N_5017,N_5582);
nor U11733 (N_11733,N_6083,N_8217);
and U11734 (N_11734,N_7917,N_7233);
xnor U11735 (N_11735,N_8989,N_9431);
xnor U11736 (N_11736,N_7223,N_8590);
nor U11737 (N_11737,N_5058,N_8108);
nand U11738 (N_11738,N_7819,N_5410);
nand U11739 (N_11739,N_9977,N_8132);
and U11740 (N_11740,N_9704,N_5591);
and U11741 (N_11741,N_5082,N_6262);
xor U11742 (N_11742,N_7901,N_6678);
or U11743 (N_11743,N_5194,N_8731);
nand U11744 (N_11744,N_8242,N_5656);
or U11745 (N_11745,N_9739,N_8995);
nor U11746 (N_11746,N_7448,N_5209);
nor U11747 (N_11747,N_8101,N_7718);
xor U11748 (N_11748,N_8948,N_6835);
nand U11749 (N_11749,N_6744,N_7412);
xor U11750 (N_11750,N_9675,N_7979);
or U11751 (N_11751,N_8631,N_9717);
or U11752 (N_11752,N_8851,N_5462);
nand U11753 (N_11753,N_8481,N_7939);
nand U11754 (N_11754,N_5853,N_9712);
nand U11755 (N_11755,N_5744,N_5461);
or U11756 (N_11756,N_6864,N_9802);
and U11757 (N_11757,N_7589,N_7533);
nor U11758 (N_11758,N_8194,N_7889);
or U11759 (N_11759,N_5165,N_5463);
or U11760 (N_11760,N_8193,N_6425);
and U11761 (N_11761,N_6255,N_8354);
xor U11762 (N_11762,N_5227,N_8062);
nor U11763 (N_11763,N_6254,N_6938);
nand U11764 (N_11764,N_7523,N_6565);
xor U11765 (N_11765,N_9854,N_9918);
and U11766 (N_11766,N_6790,N_5578);
xnor U11767 (N_11767,N_5535,N_5838);
nand U11768 (N_11768,N_9480,N_5774);
nor U11769 (N_11769,N_8426,N_7230);
or U11770 (N_11770,N_7459,N_8159);
and U11771 (N_11771,N_9251,N_7699);
or U11772 (N_11772,N_6092,N_5821);
and U11773 (N_11773,N_8664,N_6870);
nand U11774 (N_11774,N_5518,N_7873);
nand U11775 (N_11775,N_8976,N_6997);
nand U11776 (N_11776,N_6557,N_8352);
or U11777 (N_11777,N_6897,N_6531);
xor U11778 (N_11778,N_5776,N_8695);
nand U11779 (N_11779,N_5485,N_7377);
or U11780 (N_11780,N_5443,N_7733);
and U11781 (N_11781,N_7749,N_6214);
xor U11782 (N_11782,N_9870,N_7731);
xor U11783 (N_11783,N_6687,N_7771);
nor U11784 (N_11784,N_8601,N_5937);
nand U11785 (N_11785,N_8626,N_7173);
or U11786 (N_11786,N_9221,N_5818);
or U11787 (N_11787,N_9384,N_9519);
nor U11788 (N_11788,N_7415,N_5663);
or U11789 (N_11789,N_9386,N_6278);
or U11790 (N_11790,N_9117,N_5224);
nor U11791 (N_11791,N_6859,N_8834);
or U11792 (N_11792,N_9484,N_7395);
xnor U11793 (N_11793,N_9292,N_5112);
or U11794 (N_11794,N_6614,N_9467);
xnor U11795 (N_11795,N_7439,N_6025);
or U11796 (N_11796,N_9634,N_9493);
nor U11797 (N_11797,N_5892,N_5409);
xor U11798 (N_11798,N_8929,N_5363);
nor U11799 (N_11799,N_6754,N_8591);
xor U11800 (N_11800,N_9791,N_6617);
or U11801 (N_11801,N_5789,N_7139);
xor U11802 (N_11802,N_9377,N_6453);
nand U11803 (N_11803,N_6147,N_9978);
nor U11804 (N_11804,N_8126,N_7588);
xnor U11805 (N_11805,N_7371,N_5137);
nand U11806 (N_11806,N_7010,N_7752);
nor U11807 (N_11807,N_6227,N_7650);
nand U11808 (N_11808,N_6458,N_5342);
or U11809 (N_11809,N_6836,N_8155);
and U11810 (N_11810,N_9320,N_9405);
and U11811 (N_11811,N_9827,N_9172);
nand U11812 (N_11812,N_9752,N_9497);
and U11813 (N_11813,N_5677,N_5106);
or U11814 (N_11814,N_9130,N_6861);
xor U11815 (N_11815,N_5139,N_8053);
xnor U11816 (N_11816,N_9837,N_7637);
nand U11817 (N_11817,N_8188,N_7363);
or U11818 (N_11818,N_8165,N_9278);
xnor U11819 (N_11819,N_9985,N_9921);
xnor U11820 (N_11820,N_6075,N_9050);
nor U11821 (N_11821,N_6969,N_8821);
or U11822 (N_11822,N_8393,N_6690);
xnor U11823 (N_11823,N_6175,N_9126);
or U11824 (N_11824,N_9914,N_8399);
and U11825 (N_11825,N_7788,N_8476);
xnor U11826 (N_11826,N_5671,N_8903);
xnor U11827 (N_11827,N_7559,N_8550);
xor U11828 (N_11828,N_7772,N_9536);
and U11829 (N_11829,N_9534,N_6210);
and U11830 (N_11830,N_8623,N_7135);
xnor U11831 (N_11831,N_7132,N_5775);
nand U11832 (N_11832,N_9389,N_8965);
nand U11833 (N_11833,N_6528,N_9520);
nand U11834 (N_11834,N_5707,N_5624);
nor U11835 (N_11835,N_6130,N_5530);
nand U11836 (N_11836,N_9188,N_6312);
xor U11837 (N_11837,N_8514,N_6047);
and U11838 (N_11838,N_9599,N_5076);
nor U11839 (N_11839,N_6045,N_7823);
nor U11840 (N_11840,N_7179,N_9946);
nand U11841 (N_11841,N_5276,N_6658);
and U11842 (N_11842,N_5032,N_5769);
nor U11843 (N_11843,N_5799,N_5439);
or U11844 (N_11844,N_7968,N_5399);
nand U11845 (N_11845,N_7404,N_6063);
nand U11846 (N_11846,N_9351,N_6865);
nor U11847 (N_11847,N_8343,N_5329);
and U11848 (N_11848,N_9197,N_8703);
or U11849 (N_11849,N_9060,N_7961);
nor U11850 (N_11850,N_9282,N_7332);
nand U11851 (N_11851,N_6633,N_9655);
xor U11852 (N_11852,N_5946,N_9222);
nor U11853 (N_11853,N_9513,N_9570);
nor U11854 (N_11854,N_7446,N_8214);
or U11855 (N_11855,N_7674,N_8389);
nor U11856 (N_11856,N_5914,N_5159);
and U11857 (N_11857,N_5174,N_5373);
and U11858 (N_11858,N_5882,N_7755);
nor U11859 (N_11859,N_8742,N_9163);
or U11860 (N_11860,N_5694,N_7549);
or U11861 (N_11861,N_7821,N_7130);
nand U11862 (N_11862,N_6048,N_5402);
nor U11863 (N_11863,N_5951,N_5065);
xor U11864 (N_11864,N_7200,N_7004);
or U11865 (N_11865,N_9372,N_6348);
or U11866 (N_11866,N_7679,N_7560);
or U11867 (N_11867,N_8616,N_5928);
and U11868 (N_11868,N_5756,N_8815);
xnor U11869 (N_11869,N_9006,N_5127);
or U11870 (N_11870,N_8391,N_9435);
nand U11871 (N_11871,N_5150,N_9040);
and U11872 (N_11872,N_5792,N_5501);
and U11873 (N_11873,N_6132,N_8044);
nor U11874 (N_11874,N_8267,N_5529);
xnor U11875 (N_11875,N_7159,N_5425);
xor U11876 (N_11876,N_5913,N_8681);
nor U11877 (N_11877,N_5737,N_8069);
nand U11878 (N_11878,N_7364,N_8581);
nand U11879 (N_11879,N_9846,N_9248);
and U11880 (N_11880,N_9299,N_6823);
nor U11881 (N_11881,N_8922,N_9972);
or U11882 (N_11882,N_7537,N_9544);
or U11883 (N_11883,N_6189,N_9763);
nor U11884 (N_11884,N_6205,N_7751);
and U11885 (N_11885,N_8339,N_8120);
nor U11886 (N_11886,N_6731,N_6800);
nor U11887 (N_11887,N_9119,N_5741);
nor U11888 (N_11888,N_7824,N_8715);
nor U11889 (N_11889,N_9648,N_6256);
nand U11890 (N_11890,N_5836,N_6298);
and U11891 (N_11891,N_9450,N_9441);
or U11892 (N_11892,N_7787,N_9691);
nor U11893 (N_11893,N_7454,N_7137);
and U11894 (N_11894,N_7634,N_8232);
and U11895 (N_11895,N_6361,N_9862);
and U11896 (N_11896,N_5252,N_7296);
nand U11897 (N_11897,N_8794,N_8775);
and U11898 (N_11898,N_6715,N_7848);
or U11899 (N_11899,N_5289,N_6824);
xor U11900 (N_11900,N_6806,N_7799);
and U11901 (N_11901,N_6855,N_9002);
nor U11902 (N_11902,N_7176,N_8456);
or U11903 (N_11903,N_8474,N_8933);
and U11904 (N_11904,N_9466,N_5587);
nor U11905 (N_11905,N_6539,N_5250);
and U11906 (N_11906,N_6372,N_6363);
and U11907 (N_11907,N_9540,N_9617);
nor U11908 (N_11908,N_6974,N_7817);
nand U11909 (N_11909,N_8512,N_9340);
xor U11910 (N_11910,N_5680,N_9137);
nor U11911 (N_11911,N_5878,N_9677);
or U11912 (N_11912,N_7181,N_8358);
or U11913 (N_11913,N_5904,N_5950);
nor U11914 (N_11914,N_8580,N_6643);
and U11915 (N_11915,N_8899,N_6403);
xor U11916 (N_11916,N_9737,N_9049);
and U11917 (N_11917,N_7899,N_7460);
or U11918 (N_11918,N_6575,N_5679);
nand U11919 (N_11919,N_6518,N_9472);
nor U11920 (N_11920,N_9636,N_7606);
xor U11921 (N_11921,N_6176,N_5267);
nor U11922 (N_11922,N_8748,N_5803);
nand U11923 (N_11923,N_7890,N_6196);
xnor U11924 (N_11924,N_7034,N_8097);
and U11925 (N_11925,N_6857,N_5438);
and U11926 (N_11926,N_5804,N_8047);
xnor U11927 (N_11927,N_6761,N_6741);
nand U11928 (N_11928,N_6635,N_8502);
and U11929 (N_11929,N_7913,N_5754);
xor U11930 (N_11930,N_5211,N_8324);
nor U11931 (N_11931,N_8588,N_6686);
xnor U11932 (N_11932,N_6608,N_5104);
nand U11933 (N_11933,N_5630,N_9958);
xnor U11934 (N_11934,N_7903,N_7936);
and U11935 (N_11935,N_9017,N_7806);
or U11936 (N_11936,N_8970,N_6122);
nand U11937 (N_11937,N_8853,N_9635);
xnor U11938 (N_11938,N_8503,N_8743);
or U11939 (N_11939,N_5724,N_5491);
nand U11940 (N_11940,N_6758,N_6093);
or U11941 (N_11941,N_6930,N_6508);
or U11942 (N_11942,N_5023,N_6197);
or U11943 (N_11943,N_9835,N_7857);
nand U11944 (N_11944,N_8719,N_7566);
and U11945 (N_11945,N_9588,N_5287);
nor U11946 (N_11946,N_9432,N_8927);
xor U11947 (N_11947,N_7213,N_5074);
xor U11948 (N_11948,N_7563,N_6039);
and U11949 (N_11949,N_7274,N_5499);
or U11950 (N_11950,N_7023,N_5573);
xor U11951 (N_11951,N_7402,N_9262);
nand U11952 (N_11952,N_5668,N_8800);
nand U11953 (N_11953,N_8332,N_7520);
and U11954 (N_11954,N_8808,N_7545);
nand U11955 (N_11955,N_8494,N_7301);
xor U11956 (N_11956,N_7378,N_8657);
xor U11957 (N_11957,N_6207,N_6368);
xnor U11958 (N_11958,N_5527,N_9954);
xor U11959 (N_11959,N_7942,N_8613);
nor U11960 (N_11960,N_6078,N_7229);
or U11961 (N_11961,N_6530,N_7314);
xnor U11962 (N_11962,N_7678,N_5859);
xor U11963 (N_11963,N_7421,N_8019);
and U11964 (N_11964,N_6927,N_6696);
or U11965 (N_11965,N_5852,N_9581);
and U11966 (N_11966,N_5445,N_9269);
nand U11967 (N_11967,N_5693,N_8168);
nor U11968 (N_11968,N_5533,N_9058);
and U11969 (N_11969,N_5161,N_9078);
nor U11970 (N_11970,N_9853,N_8765);
or U11971 (N_11971,N_6225,N_6320);
and U11972 (N_11972,N_7062,N_8439);
and U11973 (N_11973,N_7011,N_9239);
nor U11974 (N_11974,N_6832,N_8639);
xnor U11975 (N_11975,N_5101,N_7908);
nor U11976 (N_11976,N_9829,N_5472);
nor U11977 (N_11977,N_8223,N_6229);
nand U11978 (N_11978,N_6253,N_5449);
or U11979 (N_11979,N_7321,N_5806);
xor U11980 (N_11980,N_8640,N_5997);
xnor U11981 (N_11981,N_9169,N_6186);
nor U11982 (N_11982,N_8259,N_7643);
and U11983 (N_11983,N_6359,N_9487);
xor U11984 (N_11984,N_7721,N_7949);
and U11985 (N_11985,N_6979,N_5480);
and U11986 (N_11986,N_7994,N_8868);
or U11987 (N_11987,N_8417,N_9729);
xor U11988 (N_11988,N_8603,N_6588);
nand U11989 (N_11989,N_8323,N_5639);
or U11990 (N_11990,N_8346,N_7724);
nor U11991 (N_11991,N_9471,N_6124);
or U11992 (N_11992,N_5793,N_6584);
nand U11993 (N_11993,N_9848,N_8008);
nand U11994 (N_11994,N_7375,N_9538);
and U11995 (N_11995,N_9394,N_7618);
xnor U11996 (N_11996,N_7970,N_8875);
and U11997 (N_11997,N_6379,N_8102);
nand U11998 (N_11998,N_5908,N_8357);
or U11999 (N_11999,N_6471,N_8559);
xnor U12000 (N_12000,N_8813,N_5339);
and U12001 (N_12001,N_8318,N_8106);
or U12002 (N_12002,N_8691,N_8814);
or U12003 (N_12003,N_9173,N_5444);
xnor U12004 (N_12004,N_8055,N_8672);
nand U12005 (N_12005,N_7846,N_7902);
or U12006 (N_12006,N_6926,N_9404);
or U12007 (N_12007,N_6376,N_5636);
nand U12008 (N_12008,N_6144,N_9865);
nor U12009 (N_12009,N_5008,N_8943);
xor U12010 (N_12010,N_8857,N_6313);
nand U12011 (N_12011,N_6360,N_6366);
nor U12012 (N_12012,N_9037,N_6008);
nor U12013 (N_12013,N_9725,N_7578);
and U12014 (N_12014,N_6406,N_7912);
nand U12015 (N_12015,N_9208,N_6241);
xnor U12016 (N_12016,N_9900,N_6356);
nor U12017 (N_12017,N_6552,N_7934);
or U12018 (N_12018,N_8498,N_6587);
xor U12019 (N_12019,N_7490,N_9302);
nor U12020 (N_12020,N_9926,N_5612);
or U12021 (N_12021,N_9204,N_7063);
nand U12022 (N_12022,N_6347,N_7962);
xnor U12023 (N_12023,N_9589,N_8134);
or U12024 (N_12024,N_6915,N_9613);
nand U12025 (N_12025,N_7761,N_8886);
nor U12026 (N_12026,N_9179,N_9270);
nor U12027 (N_12027,N_7734,N_8262);
or U12028 (N_12028,N_8416,N_5684);
xnor U12029 (N_12029,N_5735,N_5233);
xnor U12030 (N_12030,N_8558,N_9728);
nor U12031 (N_12031,N_7741,N_6598);
or U12032 (N_12032,N_6301,N_5186);
or U12033 (N_12033,N_5424,N_5223);
nand U12034 (N_12034,N_8049,N_7191);
nand U12035 (N_12035,N_6801,N_7938);
xnor U12036 (N_12036,N_9971,N_5087);
nand U12037 (N_12037,N_8105,N_8554);
xor U12038 (N_12038,N_9580,N_8306);
nor U12039 (N_12039,N_5839,N_5471);
nor U12040 (N_12040,N_6649,N_8646);
nand U12041 (N_12041,N_9089,N_9908);
nand U12042 (N_12042,N_9696,N_5936);
or U12043 (N_12043,N_7071,N_8666);
or U12044 (N_12044,N_8496,N_5308);
or U12045 (N_12045,N_8027,N_5290);
xnor U12046 (N_12046,N_5090,N_5673);
and U12047 (N_12047,N_6217,N_9794);
nor U12048 (N_12048,N_8757,N_7996);
or U12049 (N_12049,N_7562,N_6871);
or U12050 (N_12050,N_6375,N_6500);
and U12051 (N_12051,N_6055,N_5701);
or U12052 (N_12052,N_7847,N_7478);
nand U12053 (N_12053,N_6866,N_5083);
xnor U12054 (N_12054,N_7084,N_8706);
and U12055 (N_12055,N_5706,N_8568);
xnor U12056 (N_12056,N_6345,N_6285);
nand U12057 (N_12057,N_7383,N_5888);
nor U12058 (N_12058,N_5286,N_9861);
and U12059 (N_12059,N_7842,N_9220);
or U12060 (N_12060,N_6659,N_8673);
or U12061 (N_12061,N_7707,N_6012);
or U12062 (N_12062,N_6809,N_9120);
and U12063 (N_12063,N_6991,N_9154);
or U12064 (N_12064,N_9671,N_9530);
xnor U12065 (N_12065,N_8128,N_5268);
xor U12066 (N_12066,N_8865,N_5598);
xor U12067 (N_12067,N_9592,N_8444);
xor U12068 (N_12068,N_5686,N_6194);
or U12069 (N_12069,N_6212,N_6261);
xnor U12070 (N_12070,N_9355,N_6920);
nand U12071 (N_12071,N_5345,N_7053);
or U12072 (N_12072,N_8107,N_8523);
and U12073 (N_12073,N_7855,N_7291);
and U12074 (N_12074,N_6673,N_7776);
or U12075 (N_12075,N_5874,N_7785);
xnor U12076 (N_12076,N_8836,N_9630);
xor U12077 (N_12077,N_8939,N_7328);
nor U12078 (N_12078,N_6858,N_5322);
xnor U12079 (N_12079,N_7422,N_8316);
nand U12080 (N_12080,N_6811,N_9542);
xor U12081 (N_12081,N_5801,N_7919);
or U12082 (N_12082,N_9257,N_9910);
or U12083 (N_12083,N_7073,N_9845);
or U12084 (N_12084,N_7108,N_8963);
nor U12085 (N_12085,N_9364,N_9633);
or U12086 (N_12086,N_5609,N_5704);
nand U12087 (N_12087,N_9771,N_5380);
nand U12088 (N_12088,N_8971,N_8887);
xor U12089 (N_12089,N_5659,N_6789);
xor U12090 (N_12090,N_6542,N_7266);
nor U12091 (N_12091,N_7424,N_7599);
nor U12092 (N_12092,N_8203,N_8823);
and U12093 (N_12093,N_9063,N_8098);
xnor U12094 (N_12094,N_7382,N_8161);
and U12095 (N_12095,N_5143,N_6041);
xor U12096 (N_12096,N_9183,N_5883);
nor U12097 (N_12097,N_9271,N_5124);
and U12098 (N_12098,N_9759,N_6087);
or U12099 (N_12099,N_9632,N_9038);
and U12100 (N_12100,N_9547,N_5385);
nand U12101 (N_12101,N_9055,N_7735);
xnor U12102 (N_12102,N_7224,N_5550);
or U12103 (N_12103,N_8200,N_8859);
or U12104 (N_12104,N_6344,N_8270);
and U12105 (N_12105,N_9168,N_5798);
nor U12106 (N_12106,N_9766,N_9026);
nand U12107 (N_12107,N_8060,N_9184);
xor U12108 (N_12108,N_5819,N_7196);
xnor U12109 (N_12109,N_7985,N_9814);
nand U12110 (N_12110,N_7268,N_6091);
xor U12111 (N_12111,N_5046,N_7875);
xnor U12112 (N_12112,N_9456,N_5739);
xnor U12113 (N_12113,N_6243,N_8185);
nor U12114 (N_12114,N_6679,N_5577);
xnor U12115 (N_12115,N_6504,N_9764);
and U12116 (N_12116,N_8292,N_8781);
or U12117 (N_12117,N_7001,N_7972);
nand U12118 (N_12118,N_5554,N_6914);
xor U12119 (N_12119,N_9381,N_8001);
or U12120 (N_12120,N_9459,N_7320);
and U12121 (N_12121,N_9990,N_6675);
or U12122 (N_12122,N_7957,N_8119);
or U12123 (N_12123,N_5145,N_8897);
and U12124 (N_12124,N_9868,N_7818);
nor U12125 (N_12125,N_8199,N_7904);
nor U12126 (N_12126,N_9400,N_7205);
or U12127 (N_12127,N_9138,N_8475);
and U12128 (N_12128,N_6559,N_7577);
or U12129 (N_12129,N_9415,N_8321);
and U12130 (N_12130,N_9625,N_9504);
and U12131 (N_12131,N_8611,N_9075);
and U12132 (N_12132,N_7782,N_6882);
and U12133 (N_12133,N_6102,N_8936);
and U12134 (N_12134,N_7442,N_7104);
nor U12135 (N_12135,N_9112,N_8424);
and U12136 (N_12136,N_9077,N_7342);
xor U12137 (N_12137,N_9486,N_5722);
and U12138 (N_12138,N_9317,N_9088);
or U12139 (N_12139,N_8784,N_6209);
nand U12140 (N_12140,N_5429,N_8689);
nor U12141 (N_12141,N_7090,N_5999);
nand U12142 (N_12142,N_8839,N_7202);
nand U12143 (N_12143,N_8206,N_7703);
or U12144 (N_12144,N_6082,N_9915);
nand U12145 (N_12145,N_8793,N_6948);
xnor U12146 (N_12146,N_8016,N_7273);
nor U12147 (N_12147,N_9073,N_8013);
xnor U12148 (N_12148,N_8894,N_6568);
xnor U12149 (N_12149,N_8755,N_7885);
nor U12150 (N_12150,N_8928,N_5126);
nor U12151 (N_12151,N_8670,N_6023);
or U12152 (N_12152,N_6224,N_5569);
xor U12153 (N_12153,N_7430,N_9932);
nand U12154 (N_12154,N_8345,N_6149);
nand U12155 (N_12155,N_6842,N_9664);
nand U12156 (N_12156,N_6564,N_9924);
and U12157 (N_12157,N_8349,N_6258);
xor U12158 (N_12158,N_5715,N_5670);
and U12159 (N_12159,N_8822,N_6616);
and U12160 (N_12160,N_6306,N_8486);
nor U12161 (N_12161,N_7275,N_6697);
xor U12162 (N_12162,N_6374,N_7065);
xnor U12163 (N_12163,N_6883,N_9192);
xnor U12164 (N_12164,N_9425,N_5317);
nand U12165 (N_12165,N_7101,N_9967);
nor U12166 (N_12166,N_7872,N_8328);
nor U12167 (N_12167,N_8764,N_6631);
or U12168 (N_12168,N_8548,N_7804);
xnor U12169 (N_12169,N_7719,N_6384);
nand U12170 (N_12170,N_7381,N_7926);
or U12171 (N_12171,N_5466,N_7052);
or U12172 (N_12172,N_9798,N_9795);
or U12173 (N_12173,N_7810,N_5546);
nor U12174 (N_12174,N_7529,N_5367);
nor U12175 (N_12175,N_8737,N_7370);
xor U12176 (N_12176,N_9046,N_5512);
xor U12177 (N_12177,N_5051,N_6994);
nor U12178 (N_12178,N_6516,N_6831);
nor U12179 (N_12179,N_7288,N_6875);
nand U12180 (N_12180,N_7660,N_9631);
or U12181 (N_12181,N_6311,N_7115);
or U12182 (N_12182,N_6269,N_5514);
nand U12183 (N_12183,N_7550,N_5110);
xor U12184 (N_12184,N_6563,N_8893);
nand U12185 (N_12185,N_6955,N_6115);
and U12186 (N_12186,N_6163,N_6637);
nor U12187 (N_12187,N_7689,N_5255);
nand U12188 (N_12188,N_8795,N_7896);
nor U12189 (N_12189,N_5136,N_6145);
xor U12190 (N_12190,N_8981,N_7100);
and U12191 (N_12191,N_6006,N_8711);
and U12192 (N_12192,N_7252,N_7511);
and U12193 (N_12193,N_6562,N_5829);
nand U12194 (N_12194,N_7354,N_5055);
or U12195 (N_12195,N_8517,N_7534);
nor U12196 (N_12196,N_8602,N_7401);
nand U12197 (N_12197,N_9824,N_6665);
and U12198 (N_12198,N_8723,N_7418);
xor U12199 (N_12199,N_5274,N_5996);
xor U12200 (N_12200,N_5305,N_6726);
nor U12201 (N_12201,N_7443,N_9770);
and U12202 (N_12202,N_8848,N_7225);
and U12203 (N_12203,N_9726,N_6893);
nor U12204 (N_12204,N_6117,N_5548);
and U12205 (N_12205,N_9303,N_5699);
and U12206 (N_12206,N_8509,N_7014);
and U12207 (N_12207,N_5235,N_9461);
nor U12208 (N_12208,N_5012,N_5625);
xnor U12209 (N_12209,N_9041,N_9253);
nand U12210 (N_12210,N_6084,N_9083);
or U12211 (N_12211,N_6283,N_9276);
nor U12212 (N_12212,N_9012,N_7792);
nor U12213 (N_12213,N_6106,N_5419);
xor U12214 (N_12214,N_5651,N_9556);
or U12215 (N_12215,N_5343,N_8457);
and U12216 (N_12216,N_5192,N_7265);
nor U12217 (N_12217,N_7759,N_7532);
and U12218 (N_12218,N_9614,N_7554);
nand U12219 (N_12219,N_9573,N_8370);
or U12220 (N_12220,N_9973,N_5035);
nand U12221 (N_12221,N_6293,N_7748);
nand U12222 (N_12222,N_5247,N_5748);
xor U12223 (N_12223,N_5246,N_6463);
nor U12224 (N_12224,N_9190,N_5053);
and U12225 (N_12225,N_6231,N_5155);
xor U12226 (N_12226,N_9003,N_7186);
nand U12227 (N_12227,N_8713,N_8202);
nor U12228 (N_12228,N_5172,N_7387);
xor U12229 (N_12229,N_9053,N_8181);
nand U12230 (N_12230,N_7727,N_7765);
and U12231 (N_12231,N_8451,N_8761);
and U12232 (N_12232,N_5740,N_6628);
nor U12233 (N_12233,N_5672,N_9781);
or U12234 (N_12234,N_8325,N_7160);
or U12235 (N_12235,N_9438,N_7113);
nand U12236 (N_12236,N_6522,N_8916);
nand U12237 (N_12237,N_8729,N_8525);
and U12238 (N_12238,N_8222,N_8048);
nand U12239 (N_12239,N_9279,N_7976);
and U12240 (N_12240,N_6872,N_9256);
nand U12241 (N_12241,N_7744,N_7567);
nor U12242 (N_12242,N_6336,N_6128);
xnor U12243 (N_12243,N_6567,N_5303);
nand U12244 (N_12244,N_8634,N_6081);
and U12245 (N_12245,N_9616,N_6049);
or U12246 (N_12246,N_9565,N_5242);
or U12247 (N_12247,N_9360,N_6323);
or U12248 (N_12248,N_8909,N_9382);
and U12249 (N_12249,N_9928,N_9388);
nand U12250 (N_12250,N_9045,N_5365);
or U12251 (N_12251,N_9434,N_6495);
and U12252 (N_12252,N_7072,N_8540);
and U12253 (N_12253,N_8644,N_6887);
xor U12254 (N_12254,N_9938,N_6188);
xnor U12255 (N_12255,N_6685,N_5576);
xnor U12256 (N_12256,N_5944,N_5515);
nand U12257 (N_12257,N_9923,N_8529);
or U12258 (N_12258,N_7596,N_7240);
and U12259 (N_12259,N_9383,N_6138);
and U12260 (N_12260,N_5470,N_9879);
nand U12261 (N_12261,N_6526,N_9584);
nand U12262 (N_12262,N_9624,N_8133);
nor U12263 (N_12263,N_7131,N_5824);
nor U12264 (N_12264,N_9782,N_6165);
nor U12265 (N_12265,N_9658,N_8798);
or U12266 (N_12266,N_7013,N_7279);
and U12267 (N_12267,N_8398,N_6946);
nor U12268 (N_12268,N_9840,N_7060);
xor U12269 (N_12269,N_6491,N_8510);
or U12270 (N_12270,N_6331,N_6624);
or U12271 (N_12271,N_8949,N_8095);
or U12272 (N_12272,N_6727,N_9911);
nand U12273 (N_12273,N_6884,N_6056);
nor U12274 (N_12274,N_8219,N_5199);
nand U12275 (N_12275,N_5153,N_5856);
nand U12276 (N_12276,N_9689,N_6192);
or U12277 (N_12277,N_9122,N_7318);
nand U12278 (N_12278,N_9123,N_5099);
xnor U12279 (N_12279,N_7467,N_7664);
xnor U12280 (N_12280,N_6654,N_8261);
and U12281 (N_12281,N_5245,N_7982);
xor U12282 (N_12282,N_8197,N_6244);
nand U12283 (N_12283,N_9551,N_9524);
nand U12284 (N_12284,N_6702,N_7083);
or U12285 (N_12285,N_9640,N_8843);
nor U12286 (N_12286,N_7726,N_8528);
nand U12287 (N_12287,N_6433,N_6319);
xnor U12288 (N_12288,N_5203,N_8023);
xor U12289 (N_12289,N_5923,N_5845);
xor U12290 (N_12290,N_8837,N_8113);
nor U12291 (N_12291,N_9937,N_8980);
and U12292 (N_12292,N_9576,N_7347);
nor U12293 (N_12293,N_7966,N_6203);
nand U12294 (N_12294,N_7331,N_5033);
nor U12295 (N_12295,N_8698,N_7498);
and U12296 (N_12296,N_8129,N_7647);
nand U12297 (N_12297,N_6921,N_9560);
or U12298 (N_12298,N_8873,N_5565);
or U12299 (N_12299,N_8624,N_6745);
and U12300 (N_12300,N_5372,N_7931);
and U12301 (N_12301,N_5034,N_7677);
nand U12302 (N_12302,N_5244,N_9488);
or U12303 (N_12303,N_9148,N_6985);
nor U12304 (N_12304,N_5479,N_9984);
nor U12305 (N_12305,N_8449,N_8507);
xnor U12306 (N_12306,N_9178,N_9507);
xor U12307 (N_12307,N_5435,N_6436);
nor U12308 (N_12308,N_7324,N_8045);
or U12309 (N_12309,N_8334,N_7250);
xor U12310 (N_12310,N_5196,N_5096);
nor U12311 (N_12311,N_8000,N_8918);
nand U12312 (N_12312,N_5009,N_7393);
nand U12313 (N_12313,N_9254,N_5566);
xor U12314 (N_12314,N_5729,N_7604);
and U12315 (N_12315,N_9200,N_8987);
and U12316 (N_12316,N_7992,N_6185);
or U12317 (N_12317,N_7947,N_6878);
and U12318 (N_12318,N_9970,N_9007);
or U12319 (N_12319,N_6400,N_7058);
and U12320 (N_12320,N_9174,N_5994);
nand U12321 (N_12321,N_9226,N_5064);
xnor U12322 (N_12322,N_5213,N_9960);
xnor U12323 (N_12323,N_5149,N_8442);
nor U12324 (N_12324,N_5570,N_5777);
nand U12325 (N_12325,N_8579,N_5492);
nor U12326 (N_12326,N_8676,N_9087);
and U12327 (N_12327,N_7642,N_5752);
xnor U12328 (N_12328,N_8385,N_9145);
or U12329 (N_12329,N_6302,N_8747);
nor U12330 (N_12330,N_7682,N_8327);
or U12331 (N_12331,N_7569,N_5069);
nor U12332 (N_12332,N_6794,N_8025);
xor U12333 (N_12333,N_9035,N_6798);
or U12334 (N_12334,N_7971,N_8508);
and U12335 (N_12335,N_8211,N_5895);
nand U12336 (N_12336,N_6216,N_8368);
nor U12337 (N_12337,N_9887,N_5013);
or U12338 (N_12338,N_5520,N_9476);
or U12339 (N_12339,N_8560,N_9238);
or U12340 (N_12340,N_5759,N_5200);
nand U12341 (N_12341,N_6441,N_7127);
and U12342 (N_12342,N_9234,N_6034);
nor U12343 (N_12343,N_7042,N_8912);
nor U12344 (N_12344,N_9240,N_8247);
or U12345 (N_12345,N_9457,N_5173);
and U12346 (N_12346,N_9953,N_6461);
and U12347 (N_12347,N_9961,N_8942);
or U12348 (N_12348,N_7944,N_8849);
xnor U12349 (N_12349,N_9165,N_8333);
or U12350 (N_12350,N_5710,N_9223);
nand U12351 (N_12351,N_7675,N_7790);
nor U12352 (N_12352,N_7488,N_5500);
nand U12353 (N_12353,N_6684,N_8210);
nand U12354 (N_12354,N_8774,N_7239);
nor U12355 (N_12355,N_5953,N_9458);
and U12356 (N_12356,N_6335,N_6404);
xnor U12357 (N_12357,N_6846,N_9322);
nor U12358 (N_12358,N_7019,N_9444);
nor U12359 (N_12359,N_8395,N_7183);
or U12360 (N_12360,N_6663,N_6435);
xnor U12361 (N_12361,N_9597,N_8569);
nor U12362 (N_12362,N_8636,N_9483);
and U12363 (N_12363,N_7078,N_5049);
xor U12364 (N_12364,N_9754,N_7278);
nor U12365 (N_12365,N_6325,N_8733);
nor U12366 (N_12366,N_5388,N_9586);
or U12367 (N_12367,N_7386,N_7914);
xor U12368 (N_12368,N_8745,N_8415);
nand U12369 (N_12369,N_7432,N_7706);
nor U12370 (N_12370,N_8564,N_5760);
or U12371 (N_12371,N_6623,N_9665);
nor U12372 (N_12372,N_5341,N_7174);
nand U12373 (N_12373,N_6009,N_6142);
nand U12374 (N_12374,N_7845,N_7405);
nand U12375 (N_12375,N_8278,N_7423);
or U12376 (N_12376,N_9196,N_7835);
or U12377 (N_12377,N_9175,N_6391);
xnor U12378 (N_12378,N_9563,N_5080);
nor U12379 (N_12379,N_7997,N_9646);
or U12380 (N_12380,N_8198,N_8919);
or U12381 (N_12381,N_7747,N_7905);
and U12382 (N_12382,N_8429,N_8801);
xnor U12383 (N_12383,N_7103,N_6576);
nand U12384 (N_12384,N_5042,N_5551);
and U12385 (N_12385,N_7194,N_8984);
nand U12386 (N_12386,N_5392,N_7077);
nor U12387 (N_12387,N_9316,N_7002);
nand U12388 (N_12388,N_8104,N_8959);
xnor U12389 (N_12389,N_9583,N_7287);
xnor U12390 (N_12390,N_5958,N_9831);
and U12391 (N_12391,N_6054,N_8387);
and U12392 (N_12392,N_9166,N_7465);
xor U12393 (N_12393,N_7116,N_6226);
and U12394 (N_12394,N_7300,N_8006);
xor U12395 (N_12395,N_6155,N_5935);
xor U12396 (N_12396,N_8910,N_5045);
xnor U12397 (N_12397,N_9042,N_5534);
and U12398 (N_12398,N_9590,N_7708);
or U12399 (N_12399,N_7673,N_8951);
or U12400 (N_12400,N_6473,N_6541);
xor U12401 (N_12401,N_6671,N_9125);
and U12402 (N_12402,N_5488,N_7715);
xnor U12403 (N_12403,N_5261,N_8692);
nand U12404 (N_12404,N_8693,N_9670);
nor U12405 (N_12405,N_6833,N_8812);
and U12406 (N_12406,N_7263,N_9422);
xor U12407 (N_12407,N_8362,N_5957);
and U12408 (N_12408,N_8718,N_9418);
nand U12409 (N_12409,N_5619,N_6109);
or U12410 (N_12410,N_5976,N_8986);
and U12411 (N_12411,N_8889,N_7555);
nand U12412 (N_12412,N_5607,N_7895);
or U12413 (N_12413,N_6636,N_7350);
nor U12414 (N_12414,N_5476,N_5807);
xnor U12415 (N_12415,N_5981,N_9314);
nand U12416 (N_12416,N_8433,N_7648);
and U12417 (N_12417,N_6965,N_8592);
or U12418 (N_12418,N_6431,N_5496);
or U12419 (N_12419,N_5666,N_7969);
or U12420 (N_12420,N_7093,N_8220);
or U12421 (N_12421,N_9104,N_6351);
nor U12422 (N_12422,N_6890,N_6218);
xor U12423 (N_12423,N_6380,N_6779);
or U12424 (N_12424,N_9518,N_7877);
xnor U12425 (N_12425,N_7575,N_7390);
nor U12426 (N_12426,N_6422,N_6642);
xor U12427 (N_12427,N_8450,N_6413);
nand U12428 (N_12428,N_5742,N_8530);
nand U12429 (N_12429,N_5070,N_8351);
nor U12430 (N_12430,N_8364,N_9942);
xor U12431 (N_12431,N_7267,N_7694);
and U12432 (N_12432,N_6534,N_9298);
and U12433 (N_12433,N_5700,N_6169);
and U12434 (N_12434,N_9393,N_8829);
nor U12435 (N_12435,N_9522,N_5870);
nand U12436 (N_12436,N_7226,N_9919);
and U12437 (N_12437,N_7057,N_7929);
and U12438 (N_12438,N_5660,N_9800);
nor U12439 (N_12439,N_6387,N_6309);
or U12440 (N_12440,N_9152,N_6597);
xor U12441 (N_12441,N_7075,N_6402);
nand U12442 (N_12442,N_8031,N_7916);
nor U12443 (N_12443,N_8190,N_6774);
and U12444 (N_12444,N_9209,N_9615);
xnor U12445 (N_12445,N_7720,N_7571);
and U12446 (N_12446,N_6173,N_5236);
nor U12447 (N_12447,N_9808,N_5458);
nand U12448 (N_12448,N_9546,N_9084);
or U12449 (N_12449,N_6342,N_7349);
nor U12450 (N_12450,N_5872,N_5280);
xnor U12451 (N_12451,N_5766,N_6839);
nor U12452 (N_12452,N_5644,N_7434);
nand U12453 (N_12453,N_6966,N_5767);
and U12454 (N_12454,N_9877,N_8953);
nor U12455 (N_12455,N_6248,N_5959);
nor U12456 (N_12456,N_7227,N_5216);
or U12457 (N_12457,N_7003,N_6468);
nor U12458 (N_12458,N_8707,N_7169);
nand U12459 (N_12459,N_9920,N_7663);
nor U12460 (N_12460,N_9903,N_6470);
xor U12461 (N_12461,N_9281,N_5337);
or U12462 (N_12462,N_9465,N_9777);
and U12463 (N_12463,N_5397,N_8655);
or U12464 (N_12464,N_7920,N_9550);
nor U12465 (N_12465,N_8988,N_6982);
and U12466 (N_12466,N_6437,N_9231);
nor U12467 (N_12467,N_8908,N_7049);
nand U12468 (N_12468,N_7591,N_5900);
nand U12469 (N_12469,N_8714,N_8373);
nand U12470 (N_12470,N_8628,N_9426);
or U12471 (N_12471,N_8504,N_6993);
and U12472 (N_12472,N_8766,N_8123);
nor U12473 (N_12473,N_6432,N_5309);
and U12474 (N_12474,N_8727,N_7661);
or U12475 (N_12475,N_7697,N_8773);
or U12476 (N_12476,N_9548,N_6545);
nand U12477 (N_12477,N_7852,N_5258);
or U12478 (N_12478,N_7293,N_7138);
xor U12479 (N_12479,N_7860,N_9568);
nor U12480 (N_12480,N_5572,N_6245);
or U12481 (N_12481,N_7813,N_8513);
nand U12482 (N_12482,N_5232,N_8487);
or U12483 (N_12483,N_5662,N_6107);
nand U12484 (N_12484,N_6414,N_6369);
and U12485 (N_12485,N_9036,N_6769);
xnor U12486 (N_12486,N_5986,N_8404);
and U12487 (N_12487,N_8511,N_5608);
and U12488 (N_12488,N_5418,N_8860);
nand U12489 (N_12489,N_8818,N_9662);
nand U12490 (N_12490,N_8058,N_8828);
xnor U12491 (N_12491,N_9948,N_9380);
nor U12492 (N_12492,N_9867,N_9247);
and U12493 (N_12493,N_5866,N_8461);
and U12494 (N_12494,N_9866,N_6962);
nand U12495 (N_12495,N_7509,N_6478);
nand U12496 (N_12496,N_5206,N_8039);
and U12497 (N_12497,N_7345,N_7704);
xnor U12498 (N_12498,N_5336,N_7740);
and U12499 (N_12499,N_9508,N_7595);
or U12500 (N_12500,N_5834,N_5913);
nand U12501 (N_12501,N_9466,N_9323);
and U12502 (N_12502,N_9257,N_9994);
and U12503 (N_12503,N_9646,N_8642);
nor U12504 (N_12504,N_7007,N_7143);
or U12505 (N_12505,N_5075,N_9642);
or U12506 (N_12506,N_6113,N_6377);
xor U12507 (N_12507,N_8951,N_8323);
nor U12508 (N_12508,N_9354,N_8271);
nor U12509 (N_12509,N_9928,N_9549);
and U12510 (N_12510,N_7548,N_5889);
nor U12511 (N_12511,N_9640,N_6275);
nor U12512 (N_12512,N_9719,N_5165);
and U12513 (N_12513,N_5329,N_8517);
nor U12514 (N_12514,N_6330,N_8831);
nor U12515 (N_12515,N_5066,N_9640);
nand U12516 (N_12516,N_8706,N_6069);
xnor U12517 (N_12517,N_8115,N_6737);
nor U12518 (N_12518,N_5498,N_6462);
or U12519 (N_12519,N_6210,N_7787);
nor U12520 (N_12520,N_6114,N_5792);
and U12521 (N_12521,N_8582,N_7660);
xor U12522 (N_12522,N_7456,N_8288);
nand U12523 (N_12523,N_9642,N_8159);
and U12524 (N_12524,N_9123,N_7900);
xnor U12525 (N_12525,N_7659,N_5095);
or U12526 (N_12526,N_6097,N_5830);
nand U12527 (N_12527,N_9634,N_7673);
xor U12528 (N_12528,N_5965,N_6253);
nand U12529 (N_12529,N_5327,N_6922);
xnor U12530 (N_12530,N_7295,N_9578);
nand U12531 (N_12531,N_6629,N_7147);
xor U12532 (N_12532,N_8423,N_7013);
xnor U12533 (N_12533,N_7641,N_9690);
and U12534 (N_12534,N_9717,N_5361);
and U12535 (N_12535,N_6733,N_7026);
nand U12536 (N_12536,N_7705,N_7910);
xor U12537 (N_12537,N_8574,N_9546);
or U12538 (N_12538,N_5452,N_7751);
xnor U12539 (N_12539,N_5884,N_6851);
nand U12540 (N_12540,N_8185,N_5154);
or U12541 (N_12541,N_8371,N_9365);
nand U12542 (N_12542,N_9447,N_5571);
and U12543 (N_12543,N_9690,N_9477);
and U12544 (N_12544,N_9721,N_5418);
nand U12545 (N_12545,N_9441,N_8922);
or U12546 (N_12546,N_9039,N_6193);
and U12547 (N_12547,N_8415,N_8289);
and U12548 (N_12548,N_7144,N_8487);
or U12549 (N_12549,N_8898,N_7726);
and U12550 (N_12550,N_9494,N_8677);
and U12551 (N_12551,N_6993,N_6579);
nand U12552 (N_12552,N_9117,N_5530);
or U12553 (N_12553,N_9666,N_9072);
xnor U12554 (N_12554,N_8125,N_9605);
nor U12555 (N_12555,N_6865,N_5167);
xor U12556 (N_12556,N_8986,N_7653);
or U12557 (N_12557,N_6851,N_9261);
and U12558 (N_12558,N_5366,N_8430);
or U12559 (N_12559,N_6564,N_8647);
nand U12560 (N_12560,N_9774,N_7260);
or U12561 (N_12561,N_5750,N_8083);
nor U12562 (N_12562,N_6670,N_7293);
xnor U12563 (N_12563,N_5592,N_7764);
and U12564 (N_12564,N_8683,N_9891);
and U12565 (N_12565,N_5902,N_6005);
and U12566 (N_12566,N_7771,N_6485);
or U12567 (N_12567,N_8490,N_5066);
nand U12568 (N_12568,N_6463,N_5395);
nor U12569 (N_12569,N_8919,N_9996);
nand U12570 (N_12570,N_7641,N_8761);
and U12571 (N_12571,N_9506,N_6253);
nand U12572 (N_12572,N_8581,N_8985);
or U12573 (N_12573,N_8044,N_5562);
xor U12574 (N_12574,N_6766,N_9281);
nand U12575 (N_12575,N_8231,N_7021);
nand U12576 (N_12576,N_8492,N_8147);
xor U12577 (N_12577,N_9386,N_9673);
nand U12578 (N_12578,N_7727,N_6046);
nand U12579 (N_12579,N_8469,N_6575);
nand U12580 (N_12580,N_9070,N_7883);
nand U12581 (N_12581,N_9384,N_5613);
nand U12582 (N_12582,N_7011,N_6087);
xor U12583 (N_12583,N_6241,N_9995);
nor U12584 (N_12584,N_5158,N_9203);
xnor U12585 (N_12585,N_9647,N_5402);
xnor U12586 (N_12586,N_6287,N_9423);
or U12587 (N_12587,N_5403,N_9046);
or U12588 (N_12588,N_5905,N_5445);
nand U12589 (N_12589,N_7224,N_9641);
or U12590 (N_12590,N_8363,N_5502);
nand U12591 (N_12591,N_8446,N_6270);
xor U12592 (N_12592,N_8924,N_9533);
and U12593 (N_12593,N_8264,N_6048);
nor U12594 (N_12594,N_9436,N_7614);
nor U12595 (N_12595,N_8046,N_6040);
or U12596 (N_12596,N_8813,N_6590);
nand U12597 (N_12597,N_7979,N_7189);
and U12598 (N_12598,N_8699,N_5282);
or U12599 (N_12599,N_6923,N_5130);
or U12600 (N_12600,N_8940,N_6204);
xor U12601 (N_12601,N_5010,N_5525);
or U12602 (N_12602,N_5829,N_9960);
nand U12603 (N_12603,N_7937,N_5131);
xor U12604 (N_12604,N_5287,N_7903);
and U12605 (N_12605,N_8768,N_9193);
nor U12606 (N_12606,N_7823,N_5825);
nand U12607 (N_12607,N_9456,N_7274);
or U12608 (N_12608,N_7168,N_6501);
nand U12609 (N_12609,N_5373,N_9484);
nor U12610 (N_12610,N_8695,N_7101);
and U12611 (N_12611,N_7449,N_7892);
nor U12612 (N_12612,N_7062,N_9326);
xor U12613 (N_12613,N_5315,N_9825);
nor U12614 (N_12614,N_7377,N_9520);
or U12615 (N_12615,N_5356,N_9795);
or U12616 (N_12616,N_6973,N_9954);
nand U12617 (N_12617,N_5666,N_9099);
nand U12618 (N_12618,N_6056,N_6171);
nand U12619 (N_12619,N_8417,N_6698);
or U12620 (N_12620,N_5878,N_8475);
nor U12621 (N_12621,N_9788,N_9334);
or U12622 (N_12622,N_7564,N_9670);
and U12623 (N_12623,N_7758,N_6975);
nand U12624 (N_12624,N_8886,N_7391);
nand U12625 (N_12625,N_7638,N_8654);
and U12626 (N_12626,N_9557,N_7225);
nor U12627 (N_12627,N_8953,N_8807);
or U12628 (N_12628,N_5365,N_5401);
or U12629 (N_12629,N_7943,N_6516);
xnor U12630 (N_12630,N_6945,N_5320);
or U12631 (N_12631,N_9740,N_9734);
nor U12632 (N_12632,N_6554,N_7081);
xor U12633 (N_12633,N_7368,N_9606);
nand U12634 (N_12634,N_8940,N_8730);
xor U12635 (N_12635,N_7260,N_5585);
xnor U12636 (N_12636,N_7017,N_8241);
xnor U12637 (N_12637,N_6682,N_5288);
or U12638 (N_12638,N_5814,N_7149);
xnor U12639 (N_12639,N_7045,N_8586);
or U12640 (N_12640,N_8961,N_7751);
xnor U12641 (N_12641,N_9968,N_7788);
and U12642 (N_12642,N_7405,N_8654);
nor U12643 (N_12643,N_7078,N_5937);
xor U12644 (N_12644,N_6719,N_5980);
xnor U12645 (N_12645,N_6413,N_5174);
nand U12646 (N_12646,N_6338,N_9049);
nor U12647 (N_12647,N_9186,N_8595);
xnor U12648 (N_12648,N_7045,N_7634);
nor U12649 (N_12649,N_7559,N_8668);
xnor U12650 (N_12650,N_8100,N_9231);
nor U12651 (N_12651,N_9584,N_8501);
xor U12652 (N_12652,N_5353,N_5681);
or U12653 (N_12653,N_5786,N_5863);
xor U12654 (N_12654,N_5953,N_6697);
nand U12655 (N_12655,N_9354,N_7486);
or U12656 (N_12656,N_8502,N_7789);
and U12657 (N_12657,N_6775,N_5124);
xor U12658 (N_12658,N_6058,N_8659);
or U12659 (N_12659,N_7898,N_6037);
nor U12660 (N_12660,N_7053,N_7155);
or U12661 (N_12661,N_6163,N_6281);
and U12662 (N_12662,N_7966,N_9186);
and U12663 (N_12663,N_5468,N_5864);
xnor U12664 (N_12664,N_6714,N_7271);
nor U12665 (N_12665,N_9466,N_8848);
xnor U12666 (N_12666,N_9255,N_8430);
and U12667 (N_12667,N_7009,N_9817);
nand U12668 (N_12668,N_6136,N_8189);
nand U12669 (N_12669,N_7245,N_8343);
nor U12670 (N_12670,N_8978,N_5082);
nor U12671 (N_12671,N_6615,N_5208);
and U12672 (N_12672,N_5094,N_9695);
xor U12673 (N_12673,N_8021,N_9816);
nand U12674 (N_12674,N_9699,N_6944);
and U12675 (N_12675,N_5077,N_7249);
nand U12676 (N_12676,N_9153,N_6452);
nand U12677 (N_12677,N_7926,N_8511);
nand U12678 (N_12678,N_8338,N_6661);
nand U12679 (N_12679,N_7477,N_6958);
xnor U12680 (N_12680,N_5982,N_6828);
nor U12681 (N_12681,N_6116,N_5524);
or U12682 (N_12682,N_7580,N_5259);
nor U12683 (N_12683,N_8978,N_6280);
xnor U12684 (N_12684,N_7940,N_6191);
nand U12685 (N_12685,N_5586,N_8069);
xor U12686 (N_12686,N_8341,N_7267);
nand U12687 (N_12687,N_9004,N_7246);
or U12688 (N_12688,N_8539,N_9844);
or U12689 (N_12689,N_8796,N_5333);
nand U12690 (N_12690,N_8810,N_6555);
nor U12691 (N_12691,N_9490,N_9048);
and U12692 (N_12692,N_8559,N_6134);
nor U12693 (N_12693,N_6404,N_5670);
or U12694 (N_12694,N_6995,N_7257);
or U12695 (N_12695,N_6456,N_8223);
or U12696 (N_12696,N_5567,N_8540);
xor U12697 (N_12697,N_6692,N_9967);
nor U12698 (N_12698,N_6483,N_7907);
or U12699 (N_12699,N_7524,N_9425);
nand U12700 (N_12700,N_6213,N_8289);
nand U12701 (N_12701,N_5981,N_7631);
nand U12702 (N_12702,N_8752,N_5612);
and U12703 (N_12703,N_9196,N_9470);
nand U12704 (N_12704,N_5798,N_5322);
or U12705 (N_12705,N_6258,N_5006);
xor U12706 (N_12706,N_7132,N_6670);
nor U12707 (N_12707,N_8587,N_5356);
nor U12708 (N_12708,N_5925,N_6692);
or U12709 (N_12709,N_5163,N_6826);
nand U12710 (N_12710,N_5551,N_9942);
and U12711 (N_12711,N_9629,N_8998);
or U12712 (N_12712,N_7375,N_5060);
nand U12713 (N_12713,N_7585,N_5064);
and U12714 (N_12714,N_5969,N_7776);
xor U12715 (N_12715,N_6219,N_7993);
xnor U12716 (N_12716,N_6041,N_7345);
or U12717 (N_12717,N_9780,N_9203);
and U12718 (N_12718,N_9046,N_9198);
xor U12719 (N_12719,N_8491,N_6025);
and U12720 (N_12720,N_7956,N_9536);
nand U12721 (N_12721,N_9723,N_9002);
nand U12722 (N_12722,N_6705,N_6337);
and U12723 (N_12723,N_7986,N_9151);
nor U12724 (N_12724,N_8320,N_7652);
nor U12725 (N_12725,N_9636,N_6283);
nand U12726 (N_12726,N_8833,N_8646);
and U12727 (N_12727,N_9901,N_5851);
nand U12728 (N_12728,N_7079,N_9957);
xor U12729 (N_12729,N_9343,N_9015);
xnor U12730 (N_12730,N_8151,N_9794);
nor U12731 (N_12731,N_9662,N_5857);
or U12732 (N_12732,N_5998,N_7868);
or U12733 (N_12733,N_5681,N_8770);
xnor U12734 (N_12734,N_6537,N_5711);
nand U12735 (N_12735,N_9387,N_6841);
xnor U12736 (N_12736,N_5547,N_9269);
nand U12737 (N_12737,N_8236,N_8221);
or U12738 (N_12738,N_7815,N_5887);
and U12739 (N_12739,N_7178,N_7785);
or U12740 (N_12740,N_7845,N_9735);
or U12741 (N_12741,N_6837,N_6845);
nor U12742 (N_12742,N_5376,N_9361);
nand U12743 (N_12743,N_8859,N_8761);
xnor U12744 (N_12744,N_8372,N_6317);
or U12745 (N_12745,N_8460,N_7885);
or U12746 (N_12746,N_8959,N_6637);
and U12747 (N_12747,N_5956,N_5202);
and U12748 (N_12748,N_7534,N_6104);
nand U12749 (N_12749,N_6854,N_7188);
nor U12750 (N_12750,N_9365,N_9182);
and U12751 (N_12751,N_6620,N_7064);
nor U12752 (N_12752,N_9941,N_5361);
xnor U12753 (N_12753,N_9472,N_6168);
xnor U12754 (N_12754,N_6227,N_6194);
or U12755 (N_12755,N_6957,N_6505);
or U12756 (N_12756,N_8994,N_8654);
or U12757 (N_12757,N_9418,N_8419);
xnor U12758 (N_12758,N_5203,N_8045);
or U12759 (N_12759,N_6732,N_7887);
and U12760 (N_12760,N_8119,N_7250);
and U12761 (N_12761,N_5515,N_6843);
or U12762 (N_12762,N_5546,N_7968);
nand U12763 (N_12763,N_9706,N_5888);
or U12764 (N_12764,N_9178,N_6298);
xor U12765 (N_12765,N_7353,N_7149);
and U12766 (N_12766,N_5095,N_8323);
or U12767 (N_12767,N_9062,N_6750);
and U12768 (N_12768,N_6976,N_6302);
nor U12769 (N_12769,N_9473,N_7291);
and U12770 (N_12770,N_8485,N_8792);
nor U12771 (N_12771,N_9859,N_5108);
nor U12772 (N_12772,N_5710,N_8466);
or U12773 (N_12773,N_6320,N_8280);
nor U12774 (N_12774,N_9873,N_7742);
xnor U12775 (N_12775,N_5430,N_5195);
and U12776 (N_12776,N_6801,N_5500);
and U12777 (N_12777,N_7253,N_9371);
nor U12778 (N_12778,N_8336,N_5088);
or U12779 (N_12779,N_5821,N_8155);
nand U12780 (N_12780,N_9287,N_7225);
or U12781 (N_12781,N_7240,N_6015);
nand U12782 (N_12782,N_9386,N_7066);
nor U12783 (N_12783,N_7297,N_5096);
nand U12784 (N_12784,N_6991,N_8785);
or U12785 (N_12785,N_8691,N_8689);
nand U12786 (N_12786,N_7138,N_7830);
xnor U12787 (N_12787,N_6012,N_5469);
or U12788 (N_12788,N_8974,N_7037);
xor U12789 (N_12789,N_9955,N_5481);
and U12790 (N_12790,N_9803,N_9732);
nor U12791 (N_12791,N_5800,N_8695);
xnor U12792 (N_12792,N_7443,N_8998);
xnor U12793 (N_12793,N_8479,N_6508);
and U12794 (N_12794,N_9666,N_5211);
xnor U12795 (N_12795,N_9217,N_5642);
and U12796 (N_12796,N_8212,N_5092);
and U12797 (N_12797,N_8398,N_9575);
and U12798 (N_12798,N_8006,N_8149);
nor U12799 (N_12799,N_6605,N_9764);
nor U12800 (N_12800,N_6666,N_9650);
or U12801 (N_12801,N_9968,N_9878);
nor U12802 (N_12802,N_6519,N_6268);
xnor U12803 (N_12803,N_8911,N_7788);
xnor U12804 (N_12804,N_6777,N_5878);
xor U12805 (N_12805,N_5892,N_6366);
and U12806 (N_12806,N_9921,N_9892);
or U12807 (N_12807,N_5766,N_6497);
nor U12808 (N_12808,N_8408,N_7318);
nor U12809 (N_12809,N_6762,N_7998);
nor U12810 (N_12810,N_6435,N_6925);
nor U12811 (N_12811,N_9004,N_6733);
nand U12812 (N_12812,N_8379,N_8575);
and U12813 (N_12813,N_8195,N_8931);
xor U12814 (N_12814,N_5122,N_8320);
nor U12815 (N_12815,N_9187,N_9248);
xnor U12816 (N_12816,N_6768,N_6123);
nor U12817 (N_12817,N_5082,N_7222);
and U12818 (N_12818,N_6377,N_9625);
and U12819 (N_12819,N_5624,N_8862);
and U12820 (N_12820,N_7504,N_8655);
and U12821 (N_12821,N_5613,N_5770);
nor U12822 (N_12822,N_7538,N_9586);
and U12823 (N_12823,N_7572,N_7462);
nand U12824 (N_12824,N_9861,N_8781);
and U12825 (N_12825,N_5874,N_8794);
xnor U12826 (N_12826,N_9260,N_9697);
nor U12827 (N_12827,N_7725,N_8263);
and U12828 (N_12828,N_9018,N_7037);
or U12829 (N_12829,N_5923,N_7897);
or U12830 (N_12830,N_5744,N_5212);
nor U12831 (N_12831,N_8359,N_9406);
or U12832 (N_12832,N_7512,N_5441);
and U12833 (N_12833,N_6127,N_7275);
or U12834 (N_12834,N_5032,N_6956);
nor U12835 (N_12835,N_8467,N_8903);
and U12836 (N_12836,N_8684,N_7968);
xor U12837 (N_12837,N_7743,N_8858);
nand U12838 (N_12838,N_6336,N_6922);
xor U12839 (N_12839,N_8187,N_5401);
and U12840 (N_12840,N_6047,N_8597);
and U12841 (N_12841,N_7086,N_7586);
nand U12842 (N_12842,N_6977,N_7913);
xor U12843 (N_12843,N_5407,N_7682);
and U12844 (N_12844,N_5996,N_6045);
nor U12845 (N_12845,N_5317,N_7170);
and U12846 (N_12846,N_7336,N_6830);
nand U12847 (N_12847,N_9396,N_6169);
nand U12848 (N_12848,N_6517,N_9352);
nor U12849 (N_12849,N_8555,N_7564);
nor U12850 (N_12850,N_6826,N_9407);
nor U12851 (N_12851,N_5141,N_5530);
and U12852 (N_12852,N_5847,N_9306);
and U12853 (N_12853,N_7218,N_6000);
nor U12854 (N_12854,N_5356,N_7058);
or U12855 (N_12855,N_5793,N_8364);
nand U12856 (N_12856,N_8828,N_6239);
nand U12857 (N_12857,N_7149,N_8010);
or U12858 (N_12858,N_7285,N_8924);
or U12859 (N_12859,N_6081,N_9329);
or U12860 (N_12860,N_8808,N_9620);
and U12861 (N_12861,N_5600,N_9423);
nand U12862 (N_12862,N_8139,N_6429);
or U12863 (N_12863,N_7583,N_6101);
xor U12864 (N_12864,N_6154,N_9158);
nor U12865 (N_12865,N_7040,N_8378);
or U12866 (N_12866,N_8108,N_5830);
or U12867 (N_12867,N_6107,N_9140);
nor U12868 (N_12868,N_6064,N_9823);
or U12869 (N_12869,N_8649,N_8023);
xor U12870 (N_12870,N_5060,N_7853);
nor U12871 (N_12871,N_9074,N_9827);
or U12872 (N_12872,N_9865,N_7277);
nand U12873 (N_12873,N_9725,N_9450);
nor U12874 (N_12874,N_8422,N_9277);
nor U12875 (N_12875,N_8927,N_5566);
nand U12876 (N_12876,N_5688,N_5422);
or U12877 (N_12877,N_9977,N_7531);
nor U12878 (N_12878,N_7828,N_7273);
xnor U12879 (N_12879,N_5217,N_5947);
or U12880 (N_12880,N_8598,N_8934);
or U12881 (N_12881,N_8509,N_6879);
xor U12882 (N_12882,N_8589,N_5850);
and U12883 (N_12883,N_5931,N_8503);
and U12884 (N_12884,N_6432,N_5799);
xnor U12885 (N_12885,N_9672,N_9679);
and U12886 (N_12886,N_7196,N_6657);
xor U12887 (N_12887,N_8496,N_9025);
nor U12888 (N_12888,N_6833,N_7471);
xnor U12889 (N_12889,N_9485,N_9175);
and U12890 (N_12890,N_5107,N_6478);
nor U12891 (N_12891,N_5267,N_8651);
nor U12892 (N_12892,N_5354,N_7449);
and U12893 (N_12893,N_7723,N_7460);
nor U12894 (N_12894,N_9850,N_9340);
nand U12895 (N_12895,N_9846,N_7124);
xor U12896 (N_12896,N_8423,N_6002);
xor U12897 (N_12897,N_5296,N_8864);
nor U12898 (N_12898,N_6157,N_8037);
nand U12899 (N_12899,N_9434,N_6442);
or U12900 (N_12900,N_7893,N_8836);
and U12901 (N_12901,N_6395,N_7642);
or U12902 (N_12902,N_9395,N_6342);
xnor U12903 (N_12903,N_5513,N_5685);
xor U12904 (N_12904,N_7569,N_6794);
nand U12905 (N_12905,N_7877,N_5886);
nor U12906 (N_12906,N_5090,N_5415);
or U12907 (N_12907,N_6198,N_9146);
nor U12908 (N_12908,N_9165,N_8527);
and U12909 (N_12909,N_7444,N_6690);
and U12910 (N_12910,N_9083,N_6380);
nor U12911 (N_12911,N_8611,N_6634);
nand U12912 (N_12912,N_5052,N_8136);
nand U12913 (N_12913,N_7942,N_7524);
xnor U12914 (N_12914,N_7254,N_8392);
and U12915 (N_12915,N_7301,N_7068);
and U12916 (N_12916,N_8616,N_7659);
xor U12917 (N_12917,N_7176,N_5586);
xnor U12918 (N_12918,N_6475,N_6394);
nor U12919 (N_12919,N_7445,N_6615);
and U12920 (N_12920,N_9468,N_8575);
and U12921 (N_12921,N_6272,N_5048);
xor U12922 (N_12922,N_9471,N_5871);
xor U12923 (N_12923,N_9975,N_7500);
nand U12924 (N_12924,N_8495,N_9299);
xnor U12925 (N_12925,N_9417,N_9092);
xor U12926 (N_12926,N_5241,N_5959);
nand U12927 (N_12927,N_8577,N_8959);
or U12928 (N_12928,N_8154,N_9968);
nor U12929 (N_12929,N_8455,N_8154);
xor U12930 (N_12930,N_9822,N_5219);
nor U12931 (N_12931,N_8954,N_7016);
or U12932 (N_12932,N_9737,N_7710);
and U12933 (N_12933,N_6882,N_8271);
nand U12934 (N_12934,N_5473,N_7882);
or U12935 (N_12935,N_5466,N_7969);
and U12936 (N_12936,N_5060,N_9905);
or U12937 (N_12937,N_5960,N_7264);
or U12938 (N_12938,N_7897,N_8231);
and U12939 (N_12939,N_8952,N_6066);
xor U12940 (N_12940,N_6538,N_6688);
xor U12941 (N_12941,N_9246,N_9888);
xor U12942 (N_12942,N_8775,N_7159);
and U12943 (N_12943,N_5480,N_6091);
xor U12944 (N_12944,N_6590,N_6035);
and U12945 (N_12945,N_5137,N_7109);
or U12946 (N_12946,N_8416,N_6011);
xor U12947 (N_12947,N_9387,N_6280);
nand U12948 (N_12948,N_5650,N_9707);
nor U12949 (N_12949,N_5009,N_9397);
and U12950 (N_12950,N_5974,N_9154);
or U12951 (N_12951,N_5596,N_5807);
nor U12952 (N_12952,N_6357,N_7176);
and U12953 (N_12953,N_6022,N_6116);
and U12954 (N_12954,N_5951,N_9259);
and U12955 (N_12955,N_6793,N_9810);
and U12956 (N_12956,N_9198,N_5941);
and U12957 (N_12957,N_8533,N_6084);
xnor U12958 (N_12958,N_8719,N_9816);
nor U12959 (N_12959,N_7457,N_8886);
xor U12960 (N_12960,N_7575,N_7340);
and U12961 (N_12961,N_5596,N_7519);
xnor U12962 (N_12962,N_5110,N_8774);
xor U12963 (N_12963,N_6380,N_7143);
and U12964 (N_12964,N_5431,N_6269);
nand U12965 (N_12965,N_7266,N_8417);
xor U12966 (N_12966,N_6723,N_7228);
nand U12967 (N_12967,N_5020,N_5398);
and U12968 (N_12968,N_9976,N_9900);
and U12969 (N_12969,N_5903,N_7543);
or U12970 (N_12970,N_6501,N_6039);
xor U12971 (N_12971,N_7209,N_8456);
or U12972 (N_12972,N_8019,N_6661);
nor U12973 (N_12973,N_7596,N_9388);
and U12974 (N_12974,N_8503,N_5030);
and U12975 (N_12975,N_5548,N_6489);
xnor U12976 (N_12976,N_7792,N_5523);
or U12977 (N_12977,N_8982,N_6355);
and U12978 (N_12978,N_9381,N_9423);
nand U12979 (N_12979,N_7493,N_5908);
or U12980 (N_12980,N_7364,N_5171);
or U12981 (N_12981,N_7950,N_5111);
or U12982 (N_12982,N_9530,N_5967);
xnor U12983 (N_12983,N_8969,N_6886);
or U12984 (N_12984,N_5251,N_9669);
and U12985 (N_12985,N_7641,N_8246);
nor U12986 (N_12986,N_6532,N_9818);
nand U12987 (N_12987,N_6090,N_6350);
and U12988 (N_12988,N_5855,N_9824);
nand U12989 (N_12989,N_8334,N_9306);
or U12990 (N_12990,N_8449,N_5276);
xor U12991 (N_12991,N_7763,N_7797);
xor U12992 (N_12992,N_6444,N_8818);
nor U12993 (N_12993,N_6732,N_5992);
or U12994 (N_12994,N_8090,N_9539);
xor U12995 (N_12995,N_9602,N_5420);
xor U12996 (N_12996,N_6762,N_7921);
and U12997 (N_12997,N_8813,N_7146);
xnor U12998 (N_12998,N_6586,N_5708);
xnor U12999 (N_12999,N_8006,N_7692);
or U13000 (N_13000,N_5392,N_8947);
or U13001 (N_13001,N_8744,N_8760);
and U13002 (N_13002,N_5911,N_8398);
xnor U13003 (N_13003,N_9674,N_8863);
nand U13004 (N_13004,N_6535,N_8354);
and U13005 (N_13005,N_8408,N_9350);
xnor U13006 (N_13006,N_7689,N_7184);
nor U13007 (N_13007,N_6736,N_8111);
nor U13008 (N_13008,N_9556,N_5498);
nand U13009 (N_13009,N_6665,N_7863);
nor U13010 (N_13010,N_7344,N_9236);
or U13011 (N_13011,N_5533,N_9818);
nor U13012 (N_13012,N_8093,N_8243);
and U13013 (N_13013,N_8132,N_8327);
xnor U13014 (N_13014,N_9991,N_5238);
nor U13015 (N_13015,N_8900,N_7835);
nand U13016 (N_13016,N_9912,N_7218);
and U13017 (N_13017,N_5362,N_5246);
and U13018 (N_13018,N_7917,N_9095);
nand U13019 (N_13019,N_7003,N_8604);
or U13020 (N_13020,N_5173,N_5334);
xnor U13021 (N_13021,N_8918,N_9938);
xor U13022 (N_13022,N_6408,N_5957);
or U13023 (N_13023,N_5848,N_9862);
xnor U13024 (N_13024,N_9999,N_9314);
xnor U13025 (N_13025,N_8486,N_8131);
and U13026 (N_13026,N_9828,N_8534);
nor U13027 (N_13027,N_6570,N_5845);
or U13028 (N_13028,N_8611,N_5251);
or U13029 (N_13029,N_9050,N_6257);
nor U13030 (N_13030,N_9043,N_8249);
nand U13031 (N_13031,N_9999,N_8638);
and U13032 (N_13032,N_9691,N_6358);
or U13033 (N_13033,N_6927,N_8243);
nand U13034 (N_13034,N_8046,N_7281);
and U13035 (N_13035,N_6502,N_7991);
or U13036 (N_13036,N_9565,N_8553);
nor U13037 (N_13037,N_7354,N_6996);
xnor U13038 (N_13038,N_8026,N_5496);
xor U13039 (N_13039,N_8430,N_8190);
xnor U13040 (N_13040,N_5412,N_9025);
nand U13041 (N_13041,N_6482,N_9515);
nand U13042 (N_13042,N_7962,N_9504);
nand U13043 (N_13043,N_9388,N_7521);
xnor U13044 (N_13044,N_5395,N_9793);
and U13045 (N_13045,N_6811,N_5554);
and U13046 (N_13046,N_8584,N_9290);
nor U13047 (N_13047,N_7148,N_5113);
and U13048 (N_13048,N_5569,N_6339);
nor U13049 (N_13049,N_5883,N_5003);
xor U13050 (N_13050,N_5233,N_7773);
or U13051 (N_13051,N_7292,N_8277);
nand U13052 (N_13052,N_9839,N_9478);
and U13053 (N_13053,N_7552,N_7644);
or U13054 (N_13054,N_5925,N_5284);
nand U13055 (N_13055,N_5751,N_6315);
and U13056 (N_13056,N_7123,N_8957);
nand U13057 (N_13057,N_9985,N_6358);
and U13058 (N_13058,N_8499,N_6799);
and U13059 (N_13059,N_9562,N_9344);
or U13060 (N_13060,N_9118,N_9547);
nor U13061 (N_13061,N_6938,N_6884);
or U13062 (N_13062,N_6501,N_9898);
or U13063 (N_13063,N_5249,N_9913);
xor U13064 (N_13064,N_9084,N_9364);
xor U13065 (N_13065,N_7752,N_7992);
and U13066 (N_13066,N_7449,N_9446);
or U13067 (N_13067,N_8936,N_5172);
nand U13068 (N_13068,N_8271,N_8857);
nand U13069 (N_13069,N_7794,N_8067);
nor U13070 (N_13070,N_6901,N_7777);
nor U13071 (N_13071,N_9558,N_9497);
and U13072 (N_13072,N_7173,N_8285);
xor U13073 (N_13073,N_5051,N_5073);
nand U13074 (N_13074,N_7325,N_7087);
nand U13075 (N_13075,N_7911,N_9311);
and U13076 (N_13076,N_9713,N_8961);
or U13077 (N_13077,N_7514,N_6584);
or U13078 (N_13078,N_7843,N_9805);
or U13079 (N_13079,N_7830,N_5503);
or U13080 (N_13080,N_7525,N_8001);
and U13081 (N_13081,N_6319,N_5204);
and U13082 (N_13082,N_9501,N_9911);
nand U13083 (N_13083,N_7343,N_6643);
and U13084 (N_13084,N_8903,N_5659);
or U13085 (N_13085,N_9078,N_9411);
nand U13086 (N_13086,N_9089,N_5980);
nand U13087 (N_13087,N_5750,N_8168);
and U13088 (N_13088,N_6248,N_5847);
xor U13089 (N_13089,N_9382,N_5208);
nor U13090 (N_13090,N_5052,N_7251);
nor U13091 (N_13091,N_6981,N_5397);
nor U13092 (N_13092,N_8663,N_9521);
nor U13093 (N_13093,N_5446,N_9033);
nor U13094 (N_13094,N_6077,N_6927);
or U13095 (N_13095,N_9878,N_5817);
or U13096 (N_13096,N_6447,N_5612);
xor U13097 (N_13097,N_5124,N_8903);
xnor U13098 (N_13098,N_7022,N_5107);
nand U13099 (N_13099,N_5557,N_7973);
and U13100 (N_13100,N_8856,N_5313);
nor U13101 (N_13101,N_7980,N_9800);
nor U13102 (N_13102,N_6221,N_6746);
xor U13103 (N_13103,N_6365,N_7850);
and U13104 (N_13104,N_8450,N_8372);
xor U13105 (N_13105,N_7576,N_8275);
nor U13106 (N_13106,N_8339,N_5056);
and U13107 (N_13107,N_5228,N_8087);
nor U13108 (N_13108,N_6617,N_9693);
nand U13109 (N_13109,N_5072,N_5955);
or U13110 (N_13110,N_6208,N_5467);
nor U13111 (N_13111,N_5407,N_7349);
nor U13112 (N_13112,N_6876,N_6117);
and U13113 (N_13113,N_7311,N_6691);
and U13114 (N_13114,N_7911,N_6550);
xor U13115 (N_13115,N_9501,N_8690);
nand U13116 (N_13116,N_8978,N_8464);
or U13117 (N_13117,N_7456,N_7427);
nor U13118 (N_13118,N_5874,N_7202);
and U13119 (N_13119,N_8551,N_5780);
nor U13120 (N_13120,N_5720,N_5806);
nand U13121 (N_13121,N_5556,N_8392);
or U13122 (N_13122,N_5160,N_8400);
xor U13123 (N_13123,N_9631,N_5677);
xor U13124 (N_13124,N_7152,N_8613);
and U13125 (N_13125,N_7622,N_8757);
and U13126 (N_13126,N_7636,N_8912);
or U13127 (N_13127,N_7042,N_9252);
xor U13128 (N_13128,N_5370,N_5941);
xnor U13129 (N_13129,N_8823,N_7710);
nand U13130 (N_13130,N_8045,N_9240);
nand U13131 (N_13131,N_6003,N_5429);
and U13132 (N_13132,N_9171,N_5838);
xor U13133 (N_13133,N_6834,N_5609);
xor U13134 (N_13134,N_9831,N_5571);
and U13135 (N_13135,N_9372,N_8615);
and U13136 (N_13136,N_9911,N_9226);
xnor U13137 (N_13137,N_9718,N_8300);
nor U13138 (N_13138,N_6720,N_9091);
xnor U13139 (N_13139,N_6505,N_7700);
or U13140 (N_13140,N_5672,N_9944);
nor U13141 (N_13141,N_7056,N_9375);
nor U13142 (N_13142,N_5634,N_5602);
or U13143 (N_13143,N_8646,N_9311);
nor U13144 (N_13144,N_7022,N_5048);
nor U13145 (N_13145,N_6431,N_6688);
and U13146 (N_13146,N_8510,N_9330);
xor U13147 (N_13147,N_5888,N_7272);
nor U13148 (N_13148,N_6670,N_9292);
or U13149 (N_13149,N_9036,N_7226);
and U13150 (N_13150,N_6991,N_8226);
nand U13151 (N_13151,N_9531,N_6792);
and U13152 (N_13152,N_9128,N_9901);
xor U13153 (N_13153,N_6964,N_7151);
nor U13154 (N_13154,N_5031,N_6846);
xor U13155 (N_13155,N_8079,N_8835);
or U13156 (N_13156,N_6724,N_7584);
nand U13157 (N_13157,N_6336,N_9287);
and U13158 (N_13158,N_9565,N_7482);
nor U13159 (N_13159,N_8535,N_9470);
xnor U13160 (N_13160,N_7409,N_7667);
nand U13161 (N_13161,N_7805,N_6829);
and U13162 (N_13162,N_6215,N_6130);
or U13163 (N_13163,N_6351,N_8418);
or U13164 (N_13164,N_7249,N_8321);
or U13165 (N_13165,N_7092,N_6754);
nor U13166 (N_13166,N_7051,N_9212);
nor U13167 (N_13167,N_5523,N_5151);
nor U13168 (N_13168,N_5031,N_8496);
or U13169 (N_13169,N_6989,N_9401);
or U13170 (N_13170,N_7936,N_5077);
xor U13171 (N_13171,N_8469,N_7032);
nor U13172 (N_13172,N_6112,N_5042);
nor U13173 (N_13173,N_8391,N_9165);
and U13174 (N_13174,N_5191,N_9323);
nand U13175 (N_13175,N_6112,N_8977);
or U13176 (N_13176,N_9275,N_5955);
nand U13177 (N_13177,N_7047,N_9525);
nand U13178 (N_13178,N_5869,N_9576);
and U13179 (N_13179,N_7994,N_6225);
or U13180 (N_13180,N_8428,N_5464);
and U13181 (N_13181,N_6359,N_5946);
nor U13182 (N_13182,N_9379,N_9388);
or U13183 (N_13183,N_9774,N_6840);
nor U13184 (N_13184,N_6952,N_9014);
or U13185 (N_13185,N_5518,N_5427);
xor U13186 (N_13186,N_6028,N_9768);
xor U13187 (N_13187,N_6737,N_7475);
nand U13188 (N_13188,N_9111,N_6244);
nor U13189 (N_13189,N_9446,N_6802);
and U13190 (N_13190,N_8137,N_5503);
or U13191 (N_13191,N_9982,N_6181);
and U13192 (N_13192,N_5360,N_6745);
nand U13193 (N_13193,N_5945,N_7586);
xor U13194 (N_13194,N_9994,N_6786);
or U13195 (N_13195,N_6772,N_5562);
and U13196 (N_13196,N_9147,N_8484);
nor U13197 (N_13197,N_6757,N_6729);
or U13198 (N_13198,N_7745,N_6533);
nor U13199 (N_13199,N_6263,N_7676);
nand U13200 (N_13200,N_5430,N_5021);
nor U13201 (N_13201,N_5443,N_5313);
and U13202 (N_13202,N_8042,N_8975);
nand U13203 (N_13203,N_7237,N_6971);
and U13204 (N_13204,N_5356,N_5050);
and U13205 (N_13205,N_5677,N_9460);
and U13206 (N_13206,N_7360,N_5136);
or U13207 (N_13207,N_5180,N_5518);
or U13208 (N_13208,N_9036,N_8320);
or U13209 (N_13209,N_8152,N_7020);
xor U13210 (N_13210,N_6159,N_9542);
or U13211 (N_13211,N_7390,N_5233);
nand U13212 (N_13212,N_6028,N_5123);
or U13213 (N_13213,N_5875,N_6356);
xor U13214 (N_13214,N_7817,N_7540);
xnor U13215 (N_13215,N_5225,N_7120);
xor U13216 (N_13216,N_5283,N_8387);
and U13217 (N_13217,N_8319,N_9523);
or U13218 (N_13218,N_7228,N_5106);
nor U13219 (N_13219,N_5159,N_8226);
and U13220 (N_13220,N_6426,N_7124);
or U13221 (N_13221,N_5901,N_7541);
and U13222 (N_13222,N_5381,N_6105);
nand U13223 (N_13223,N_8868,N_6042);
or U13224 (N_13224,N_6113,N_5820);
xnor U13225 (N_13225,N_6317,N_6860);
or U13226 (N_13226,N_7432,N_8269);
and U13227 (N_13227,N_5039,N_9521);
nand U13228 (N_13228,N_8043,N_6805);
and U13229 (N_13229,N_6391,N_9702);
or U13230 (N_13230,N_9345,N_6447);
nand U13231 (N_13231,N_5038,N_6220);
xor U13232 (N_13232,N_8298,N_8446);
nand U13233 (N_13233,N_8143,N_8532);
or U13234 (N_13234,N_6291,N_7223);
nor U13235 (N_13235,N_6257,N_5191);
and U13236 (N_13236,N_7460,N_7797);
nand U13237 (N_13237,N_8279,N_5938);
nor U13238 (N_13238,N_6441,N_6298);
nand U13239 (N_13239,N_7622,N_6139);
and U13240 (N_13240,N_5259,N_8719);
and U13241 (N_13241,N_7708,N_9906);
or U13242 (N_13242,N_9280,N_7554);
xor U13243 (N_13243,N_7570,N_7577);
nand U13244 (N_13244,N_8888,N_6428);
nand U13245 (N_13245,N_9634,N_7616);
nand U13246 (N_13246,N_9932,N_6527);
or U13247 (N_13247,N_9244,N_6154);
and U13248 (N_13248,N_6411,N_9933);
nor U13249 (N_13249,N_7327,N_8816);
and U13250 (N_13250,N_9948,N_8740);
xnor U13251 (N_13251,N_9925,N_6089);
or U13252 (N_13252,N_5866,N_7263);
nor U13253 (N_13253,N_5809,N_7957);
xor U13254 (N_13254,N_7787,N_9108);
nor U13255 (N_13255,N_9588,N_7568);
nor U13256 (N_13256,N_8064,N_7266);
and U13257 (N_13257,N_6015,N_7331);
nor U13258 (N_13258,N_8673,N_8936);
and U13259 (N_13259,N_8676,N_6169);
and U13260 (N_13260,N_9854,N_6530);
and U13261 (N_13261,N_9899,N_9912);
and U13262 (N_13262,N_5156,N_8263);
xnor U13263 (N_13263,N_7811,N_8979);
xnor U13264 (N_13264,N_5359,N_7551);
nor U13265 (N_13265,N_6578,N_9685);
xnor U13266 (N_13266,N_9698,N_6325);
or U13267 (N_13267,N_6631,N_5997);
or U13268 (N_13268,N_8193,N_6744);
nand U13269 (N_13269,N_8559,N_8436);
or U13270 (N_13270,N_9782,N_8606);
and U13271 (N_13271,N_9017,N_6735);
nand U13272 (N_13272,N_5540,N_6070);
nor U13273 (N_13273,N_5445,N_7361);
nor U13274 (N_13274,N_5612,N_7591);
xor U13275 (N_13275,N_5197,N_9414);
xor U13276 (N_13276,N_7325,N_5184);
or U13277 (N_13277,N_6563,N_7525);
or U13278 (N_13278,N_8015,N_8197);
xnor U13279 (N_13279,N_6464,N_6961);
xor U13280 (N_13280,N_8859,N_7874);
and U13281 (N_13281,N_5293,N_9671);
and U13282 (N_13282,N_9036,N_7219);
and U13283 (N_13283,N_9899,N_8263);
nand U13284 (N_13284,N_8382,N_6232);
xor U13285 (N_13285,N_9521,N_7944);
nand U13286 (N_13286,N_7878,N_8738);
nor U13287 (N_13287,N_6220,N_7286);
xor U13288 (N_13288,N_9644,N_8114);
nand U13289 (N_13289,N_6150,N_9121);
nor U13290 (N_13290,N_8643,N_9779);
and U13291 (N_13291,N_5000,N_6087);
xor U13292 (N_13292,N_8723,N_5404);
nor U13293 (N_13293,N_7895,N_6277);
nor U13294 (N_13294,N_6913,N_8534);
and U13295 (N_13295,N_8053,N_9111);
or U13296 (N_13296,N_6132,N_8614);
and U13297 (N_13297,N_8082,N_9865);
nor U13298 (N_13298,N_8922,N_9290);
or U13299 (N_13299,N_7420,N_7601);
nand U13300 (N_13300,N_5576,N_5615);
or U13301 (N_13301,N_7500,N_9672);
nand U13302 (N_13302,N_8587,N_5231);
nor U13303 (N_13303,N_5942,N_7520);
nand U13304 (N_13304,N_6576,N_7172);
xnor U13305 (N_13305,N_5428,N_6382);
xor U13306 (N_13306,N_9578,N_7407);
or U13307 (N_13307,N_6149,N_8845);
or U13308 (N_13308,N_8744,N_9689);
nand U13309 (N_13309,N_5701,N_5906);
or U13310 (N_13310,N_5601,N_7349);
and U13311 (N_13311,N_8756,N_7947);
nand U13312 (N_13312,N_9110,N_8831);
xnor U13313 (N_13313,N_6746,N_5884);
and U13314 (N_13314,N_5059,N_8503);
xnor U13315 (N_13315,N_6682,N_5041);
xnor U13316 (N_13316,N_6144,N_5589);
xnor U13317 (N_13317,N_8416,N_6376);
or U13318 (N_13318,N_6440,N_6387);
nor U13319 (N_13319,N_9226,N_5845);
nor U13320 (N_13320,N_5674,N_7972);
nor U13321 (N_13321,N_6068,N_5665);
and U13322 (N_13322,N_7828,N_7376);
xor U13323 (N_13323,N_5661,N_5718);
xor U13324 (N_13324,N_7903,N_7630);
xnor U13325 (N_13325,N_8076,N_6947);
and U13326 (N_13326,N_7478,N_5934);
xnor U13327 (N_13327,N_6165,N_8111);
or U13328 (N_13328,N_7483,N_8536);
and U13329 (N_13329,N_6659,N_7979);
nand U13330 (N_13330,N_8489,N_6671);
and U13331 (N_13331,N_6396,N_5116);
xor U13332 (N_13332,N_6087,N_9486);
nor U13333 (N_13333,N_6398,N_7250);
nand U13334 (N_13334,N_5745,N_5195);
and U13335 (N_13335,N_6949,N_6386);
nor U13336 (N_13336,N_9317,N_5150);
or U13337 (N_13337,N_6763,N_5117);
nand U13338 (N_13338,N_8778,N_7102);
xor U13339 (N_13339,N_8918,N_6289);
and U13340 (N_13340,N_8914,N_5509);
nor U13341 (N_13341,N_7983,N_8521);
xor U13342 (N_13342,N_9782,N_5764);
nand U13343 (N_13343,N_9174,N_6924);
nand U13344 (N_13344,N_9480,N_7416);
nand U13345 (N_13345,N_6066,N_7338);
nor U13346 (N_13346,N_5905,N_8805);
or U13347 (N_13347,N_6791,N_9222);
or U13348 (N_13348,N_6404,N_6301);
or U13349 (N_13349,N_7470,N_6369);
xor U13350 (N_13350,N_6517,N_6779);
or U13351 (N_13351,N_8682,N_5219);
and U13352 (N_13352,N_8056,N_8314);
nor U13353 (N_13353,N_5301,N_8347);
and U13354 (N_13354,N_6721,N_6452);
nand U13355 (N_13355,N_6087,N_9324);
nor U13356 (N_13356,N_5988,N_7869);
and U13357 (N_13357,N_7104,N_8031);
or U13358 (N_13358,N_5409,N_8498);
xor U13359 (N_13359,N_7385,N_7180);
nor U13360 (N_13360,N_8622,N_8815);
nand U13361 (N_13361,N_8277,N_9770);
xor U13362 (N_13362,N_8565,N_7880);
or U13363 (N_13363,N_7739,N_9897);
nor U13364 (N_13364,N_8966,N_7742);
nand U13365 (N_13365,N_7891,N_6834);
nand U13366 (N_13366,N_8380,N_7848);
nand U13367 (N_13367,N_8816,N_9400);
and U13368 (N_13368,N_5577,N_6926);
and U13369 (N_13369,N_8878,N_6609);
and U13370 (N_13370,N_5217,N_8935);
xnor U13371 (N_13371,N_6891,N_6897);
and U13372 (N_13372,N_9519,N_5829);
xor U13373 (N_13373,N_6768,N_7136);
nor U13374 (N_13374,N_9890,N_6265);
xor U13375 (N_13375,N_6225,N_7120);
or U13376 (N_13376,N_7734,N_7789);
nand U13377 (N_13377,N_9469,N_7878);
and U13378 (N_13378,N_7540,N_9102);
or U13379 (N_13379,N_8276,N_5866);
xor U13380 (N_13380,N_5404,N_9194);
nor U13381 (N_13381,N_9734,N_9376);
xor U13382 (N_13382,N_8521,N_9290);
nor U13383 (N_13383,N_7907,N_5280);
nor U13384 (N_13384,N_6624,N_7943);
nand U13385 (N_13385,N_7912,N_9244);
nand U13386 (N_13386,N_8088,N_5642);
nor U13387 (N_13387,N_5145,N_7245);
xor U13388 (N_13388,N_5940,N_5122);
or U13389 (N_13389,N_7089,N_8028);
xor U13390 (N_13390,N_6812,N_6469);
or U13391 (N_13391,N_6552,N_7150);
nor U13392 (N_13392,N_6184,N_6031);
nor U13393 (N_13393,N_5144,N_7209);
xnor U13394 (N_13394,N_5939,N_7692);
xor U13395 (N_13395,N_9427,N_8239);
or U13396 (N_13396,N_7754,N_9909);
nand U13397 (N_13397,N_9702,N_5879);
and U13398 (N_13398,N_8171,N_8511);
nor U13399 (N_13399,N_7285,N_6758);
and U13400 (N_13400,N_9161,N_5750);
xnor U13401 (N_13401,N_7731,N_9577);
or U13402 (N_13402,N_6395,N_9739);
nor U13403 (N_13403,N_7815,N_5873);
or U13404 (N_13404,N_9395,N_7832);
nand U13405 (N_13405,N_6869,N_7678);
or U13406 (N_13406,N_6580,N_8648);
or U13407 (N_13407,N_5598,N_8288);
and U13408 (N_13408,N_9878,N_8302);
xor U13409 (N_13409,N_8957,N_5200);
xor U13410 (N_13410,N_7110,N_8037);
nand U13411 (N_13411,N_5956,N_6185);
or U13412 (N_13412,N_5340,N_8762);
nand U13413 (N_13413,N_5807,N_8846);
nor U13414 (N_13414,N_8388,N_7632);
or U13415 (N_13415,N_7996,N_5661);
or U13416 (N_13416,N_5825,N_9021);
or U13417 (N_13417,N_6128,N_6960);
and U13418 (N_13418,N_9182,N_9360);
nor U13419 (N_13419,N_7629,N_8319);
nand U13420 (N_13420,N_6493,N_5066);
nand U13421 (N_13421,N_8593,N_6172);
nand U13422 (N_13422,N_8394,N_8879);
and U13423 (N_13423,N_6214,N_6488);
nand U13424 (N_13424,N_6709,N_9524);
and U13425 (N_13425,N_9556,N_6782);
nand U13426 (N_13426,N_7324,N_8835);
nand U13427 (N_13427,N_8808,N_9109);
nor U13428 (N_13428,N_6475,N_6964);
xnor U13429 (N_13429,N_5231,N_6218);
or U13430 (N_13430,N_5437,N_9955);
and U13431 (N_13431,N_5302,N_6853);
xor U13432 (N_13432,N_6309,N_8342);
and U13433 (N_13433,N_8688,N_7470);
xnor U13434 (N_13434,N_5225,N_5691);
nor U13435 (N_13435,N_7671,N_8205);
xor U13436 (N_13436,N_8275,N_5986);
nor U13437 (N_13437,N_8307,N_6154);
or U13438 (N_13438,N_8587,N_5706);
nand U13439 (N_13439,N_5493,N_8686);
nand U13440 (N_13440,N_9150,N_7669);
nand U13441 (N_13441,N_5097,N_8994);
nand U13442 (N_13442,N_7468,N_8698);
xor U13443 (N_13443,N_7072,N_7174);
nand U13444 (N_13444,N_5639,N_6552);
xor U13445 (N_13445,N_6846,N_5927);
nor U13446 (N_13446,N_9900,N_7056);
xor U13447 (N_13447,N_5478,N_7725);
or U13448 (N_13448,N_9305,N_6299);
nand U13449 (N_13449,N_6142,N_6963);
nand U13450 (N_13450,N_5041,N_5031);
and U13451 (N_13451,N_8577,N_7837);
and U13452 (N_13452,N_8929,N_5296);
xnor U13453 (N_13453,N_7526,N_6908);
nor U13454 (N_13454,N_6122,N_6980);
xor U13455 (N_13455,N_6380,N_8064);
and U13456 (N_13456,N_8408,N_9219);
nand U13457 (N_13457,N_9734,N_8343);
or U13458 (N_13458,N_9062,N_9042);
or U13459 (N_13459,N_7394,N_8354);
or U13460 (N_13460,N_6846,N_9265);
xor U13461 (N_13461,N_5706,N_7088);
nand U13462 (N_13462,N_6511,N_8067);
nor U13463 (N_13463,N_7244,N_6732);
nand U13464 (N_13464,N_9737,N_6123);
xnor U13465 (N_13465,N_7454,N_5265);
or U13466 (N_13466,N_8855,N_6630);
nand U13467 (N_13467,N_7006,N_9562);
or U13468 (N_13468,N_7007,N_7384);
xnor U13469 (N_13469,N_7492,N_7895);
or U13470 (N_13470,N_9518,N_5858);
nand U13471 (N_13471,N_7720,N_6934);
nand U13472 (N_13472,N_9771,N_6652);
nor U13473 (N_13473,N_7085,N_9437);
or U13474 (N_13474,N_9499,N_6879);
nor U13475 (N_13475,N_9311,N_5729);
nor U13476 (N_13476,N_7898,N_6790);
or U13477 (N_13477,N_9009,N_6535);
xnor U13478 (N_13478,N_5070,N_8409);
nand U13479 (N_13479,N_8653,N_6788);
nor U13480 (N_13480,N_9468,N_5655);
and U13481 (N_13481,N_8603,N_9871);
nor U13482 (N_13482,N_5639,N_6202);
nor U13483 (N_13483,N_9701,N_5634);
nand U13484 (N_13484,N_7865,N_8348);
and U13485 (N_13485,N_6330,N_8559);
nand U13486 (N_13486,N_7660,N_5874);
and U13487 (N_13487,N_9675,N_5453);
and U13488 (N_13488,N_5879,N_8619);
nor U13489 (N_13489,N_7635,N_5821);
or U13490 (N_13490,N_8536,N_7752);
nand U13491 (N_13491,N_8087,N_6377);
nand U13492 (N_13492,N_7559,N_8500);
nand U13493 (N_13493,N_5747,N_7954);
nor U13494 (N_13494,N_5222,N_5072);
or U13495 (N_13495,N_7941,N_7444);
nand U13496 (N_13496,N_6034,N_9213);
nand U13497 (N_13497,N_9996,N_7978);
and U13498 (N_13498,N_6708,N_7664);
nor U13499 (N_13499,N_9617,N_8453);
xor U13500 (N_13500,N_7459,N_5836);
or U13501 (N_13501,N_5448,N_9993);
or U13502 (N_13502,N_6725,N_7555);
nor U13503 (N_13503,N_5869,N_7414);
and U13504 (N_13504,N_9022,N_7754);
nor U13505 (N_13505,N_8467,N_7386);
nor U13506 (N_13506,N_9227,N_9845);
nand U13507 (N_13507,N_7721,N_9909);
or U13508 (N_13508,N_8466,N_7679);
or U13509 (N_13509,N_6080,N_5816);
or U13510 (N_13510,N_6289,N_8424);
or U13511 (N_13511,N_6194,N_5014);
or U13512 (N_13512,N_5827,N_8083);
and U13513 (N_13513,N_7036,N_5959);
nor U13514 (N_13514,N_7233,N_7176);
or U13515 (N_13515,N_9169,N_8509);
xor U13516 (N_13516,N_6267,N_9880);
nor U13517 (N_13517,N_5763,N_9074);
nand U13518 (N_13518,N_8613,N_5361);
xor U13519 (N_13519,N_5495,N_7034);
or U13520 (N_13520,N_7123,N_8214);
and U13521 (N_13521,N_9923,N_5122);
xnor U13522 (N_13522,N_8775,N_7319);
nor U13523 (N_13523,N_8433,N_7722);
or U13524 (N_13524,N_9430,N_5378);
xor U13525 (N_13525,N_5672,N_9209);
xnor U13526 (N_13526,N_5044,N_8582);
and U13527 (N_13527,N_7495,N_5433);
or U13528 (N_13528,N_5618,N_9303);
nand U13529 (N_13529,N_6127,N_6982);
nand U13530 (N_13530,N_8788,N_6773);
and U13531 (N_13531,N_5835,N_6375);
xor U13532 (N_13532,N_7080,N_9764);
or U13533 (N_13533,N_6208,N_6507);
nand U13534 (N_13534,N_7380,N_8553);
xnor U13535 (N_13535,N_7074,N_6519);
nor U13536 (N_13536,N_6409,N_6704);
or U13537 (N_13537,N_7320,N_8367);
and U13538 (N_13538,N_5771,N_5802);
xor U13539 (N_13539,N_5002,N_8119);
xnor U13540 (N_13540,N_7312,N_8993);
xor U13541 (N_13541,N_7470,N_9738);
nand U13542 (N_13542,N_9546,N_5916);
nand U13543 (N_13543,N_9165,N_5357);
nor U13544 (N_13544,N_5633,N_9691);
and U13545 (N_13545,N_7733,N_6455);
and U13546 (N_13546,N_7503,N_9950);
nand U13547 (N_13547,N_7624,N_7212);
and U13548 (N_13548,N_9868,N_6702);
or U13549 (N_13549,N_9391,N_5155);
or U13550 (N_13550,N_9263,N_9764);
and U13551 (N_13551,N_6940,N_9339);
nand U13552 (N_13552,N_5593,N_5463);
xnor U13553 (N_13553,N_5894,N_9929);
or U13554 (N_13554,N_5547,N_5695);
xor U13555 (N_13555,N_6598,N_7844);
or U13556 (N_13556,N_6450,N_9848);
xor U13557 (N_13557,N_6392,N_6252);
xor U13558 (N_13558,N_5962,N_7343);
and U13559 (N_13559,N_9515,N_6187);
nand U13560 (N_13560,N_6784,N_8810);
or U13561 (N_13561,N_7645,N_9261);
or U13562 (N_13562,N_6160,N_9442);
and U13563 (N_13563,N_8352,N_7002);
nand U13564 (N_13564,N_7108,N_9399);
or U13565 (N_13565,N_6231,N_5247);
xor U13566 (N_13566,N_5347,N_5597);
xor U13567 (N_13567,N_5308,N_7469);
or U13568 (N_13568,N_6296,N_5259);
and U13569 (N_13569,N_7765,N_8032);
nor U13570 (N_13570,N_8662,N_9629);
and U13571 (N_13571,N_6187,N_8488);
and U13572 (N_13572,N_9765,N_7994);
and U13573 (N_13573,N_5988,N_7129);
xnor U13574 (N_13574,N_5023,N_8683);
or U13575 (N_13575,N_7702,N_9723);
xor U13576 (N_13576,N_6099,N_7367);
or U13577 (N_13577,N_6666,N_8251);
nor U13578 (N_13578,N_5548,N_6490);
xnor U13579 (N_13579,N_8925,N_5588);
and U13580 (N_13580,N_9418,N_8530);
xnor U13581 (N_13581,N_6996,N_9633);
or U13582 (N_13582,N_7609,N_8848);
and U13583 (N_13583,N_6807,N_8396);
nand U13584 (N_13584,N_9588,N_7327);
or U13585 (N_13585,N_5591,N_8713);
or U13586 (N_13586,N_9732,N_6513);
nand U13587 (N_13587,N_9458,N_6766);
and U13588 (N_13588,N_6699,N_9252);
or U13589 (N_13589,N_8271,N_6915);
nand U13590 (N_13590,N_7094,N_8487);
or U13591 (N_13591,N_6036,N_8706);
or U13592 (N_13592,N_6102,N_9192);
xor U13593 (N_13593,N_6518,N_6023);
or U13594 (N_13594,N_9217,N_6268);
or U13595 (N_13595,N_5519,N_5085);
xnor U13596 (N_13596,N_7409,N_6321);
xnor U13597 (N_13597,N_7899,N_9699);
and U13598 (N_13598,N_9218,N_7816);
and U13599 (N_13599,N_8778,N_7507);
and U13600 (N_13600,N_8215,N_9455);
nor U13601 (N_13601,N_8032,N_7959);
nor U13602 (N_13602,N_6869,N_7670);
nand U13603 (N_13603,N_6895,N_5311);
xor U13604 (N_13604,N_9836,N_6387);
nor U13605 (N_13605,N_6565,N_8054);
or U13606 (N_13606,N_6095,N_7187);
xnor U13607 (N_13607,N_9664,N_7305);
nor U13608 (N_13608,N_6914,N_6867);
xnor U13609 (N_13609,N_8063,N_8195);
xor U13610 (N_13610,N_8105,N_9320);
xor U13611 (N_13611,N_5641,N_8302);
and U13612 (N_13612,N_8955,N_7459);
nor U13613 (N_13613,N_5403,N_9374);
nand U13614 (N_13614,N_5648,N_8002);
nor U13615 (N_13615,N_9268,N_5376);
or U13616 (N_13616,N_8034,N_8928);
nor U13617 (N_13617,N_8333,N_9893);
or U13618 (N_13618,N_8777,N_9936);
nor U13619 (N_13619,N_7947,N_7374);
or U13620 (N_13620,N_7201,N_5685);
and U13621 (N_13621,N_6209,N_9745);
nor U13622 (N_13622,N_6922,N_9728);
and U13623 (N_13623,N_5775,N_5067);
xor U13624 (N_13624,N_8159,N_6308);
xor U13625 (N_13625,N_5853,N_7979);
nand U13626 (N_13626,N_5938,N_9556);
nor U13627 (N_13627,N_9375,N_6832);
xor U13628 (N_13628,N_9444,N_7745);
nand U13629 (N_13629,N_8057,N_9096);
nor U13630 (N_13630,N_8933,N_8435);
nor U13631 (N_13631,N_6667,N_9917);
nand U13632 (N_13632,N_9623,N_9394);
xor U13633 (N_13633,N_8497,N_7702);
or U13634 (N_13634,N_8236,N_9528);
nand U13635 (N_13635,N_9161,N_6160);
nand U13636 (N_13636,N_8208,N_7477);
xor U13637 (N_13637,N_8823,N_7246);
xor U13638 (N_13638,N_5611,N_9668);
nor U13639 (N_13639,N_5199,N_6489);
nand U13640 (N_13640,N_8253,N_7519);
nand U13641 (N_13641,N_6359,N_8717);
or U13642 (N_13642,N_5536,N_5071);
or U13643 (N_13643,N_5526,N_6939);
nor U13644 (N_13644,N_9945,N_8116);
and U13645 (N_13645,N_9322,N_8146);
xor U13646 (N_13646,N_8193,N_5766);
and U13647 (N_13647,N_8339,N_8077);
nand U13648 (N_13648,N_9833,N_7877);
nand U13649 (N_13649,N_9432,N_8911);
or U13650 (N_13650,N_7453,N_7165);
or U13651 (N_13651,N_7032,N_5515);
nor U13652 (N_13652,N_5642,N_9948);
xnor U13653 (N_13653,N_6998,N_6647);
and U13654 (N_13654,N_7768,N_7319);
xnor U13655 (N_13655,N_5531,N_9554);
and U13656 (N_13656,N_9377,N_9513);
and U13657 (N_13657,N_8789,N_7891);
nor U13658 (N_13658,N_6745,N_5376);
nand U13659 (N_13659,N_9334,N_7463);
xnor U13660 (N_13660,N_7358,N_6860);
xnor U13661 (N_13661,N_7825,N_8557);
nand U13662 (N_13662,N_8852,N_6314);
and U13663 (N_13663,N_5155,N_8550);
and U13664 (N_13664,N_5091,N_7580);
and U13665 (N_13665,N_7707,N_7331);
and U13666 (N_13666,N_5421,N_7840);
nand U13667 (N_13667,N_5144,N_6380);
and U13668 (N_13668,N_6546,N_6234);
nand U13669 (N_13669,N_5163,N_5795);
and U13670 (N_13670,N_9501,N_5077);
nor U13671 (N_13671,N_7060,N_8311);
or U13672 (N_13672,N_6445,N_9841);
nand U13673 (N_13673,N_9788,N_9900);
and U13674 (N_13674,N_5798,N_8926);
nor U13675 (N_13675,N_6815,N_5001);
and U13676 (N_13676,N_6074,N_6318);
nor U13677 (N_13677,N_9609,N_8321);
nand U13678 (N_13678,N_5383,N_9458);
or U13679 (N_13679,N_5358,N_7947);
nor U13680 (N_13680,N_8590,N_6684);
xor U13681 (N_13681,N_8789,N_6080);
and U13682 (N_13682,N_9164,N_8300);
or U13683 (N_13683,N_6447,N_5311);
nor U13684 (N_13684,N_6008,N_6793);
and U13685 (N_13685,N_6517,N_8364);
nand U13686 (N_13686,N_7173,N_7374);
nor U13687 (N_13687,N_6360,N_5579);
xnor U13688 (N_13688,N_6268,N_5123);
xor U13689 (N_13689,N_6639,N_7231);
or U13690 (N_13690,N_6707,N_6272);
xnor U13691 (N_13691,N_7576,N_6360);
or U13692 (N_13692,N_7611,N_8760);
xor U13693 (N_13693,N_9494,N_9623);
nor U13694 (N_13694,N_6085,N_6937);
nor U13695 (N_13695,N_7786,N_6519);
nor U13696 (N_13696,N_6589,N_6883);
xnor U13697 (N_13697,N_8630,N_5262);
nor U13698 (N_13698,N_5073,N_6247);
and U13699 (N_13699,N_5559,N_8474);
xor U13700 (N_13700,N_7880,N_5328);
or U13701 (N_13701,N_9110,N_7534);
nor U13702 (N_13702,N_9067,N_7001);
xor U13703 (N_13703,N_5501,N_5720);
nand U13704 (N_13704,N_6237,N_9829);
or U13705 (N_13705,N_5002,N_7028);
nor U13706 (N_13706,N_8639,N_6026);
nor U13707 (N_13707,N_7382,N_8440);
and U13708 (N_13708,N_7160,N_6111);
xor U13709 (N_13709,N_9116,N_6310);
xor U13710 (N_13710,N_9820,N_5376);
and U13711 (N_13711,N_8170,N_9494);
or U13712 (N_13712,N_7972,N_6865);
xnor U13713 (N_13713,N_7628,N_8084);
xor U13714 (N_13714,N_9692,N_5043);
xor U13715 (N_13715,N_5481,N_6610);
or U13716 (N_13716,N_7329,N_8364);
or U13717 (N_13717,N_5418,N_6477);
and U13718 (N_13718,N_7361,N_7964);
or U13719 (N_13719,N_6951,N_6755);
and U13720 (N_13720,N_7597,N_7507);
or U13721 (N_13721,N_8292,N_7764);
or U13722 (N_13722,N_6170,N_5069);
nor U13723 (N_13723,N_8603,N_5140);
or U13724 (N_13724,N_9485,N_6720);
xor U13725 (N_13725,N_6660,N_6967);
xnor U13726 (N_13726,N_9708,N_9286);
nor U13727 (N_13727,N_7993,N_5616);
and U13728 (N_13728,N_5664,N_9355);
nand U13729 (N_13729,N_9878,N_5120);
nor U13730 (N_13730,N_9137,N_8241);
nor U13731 (N_13731,N_7028,N_7687);
nand U13732 (N_13732,N_5123,N_7407);
nor U13733 (N_13733,N_9061,N_6192);
and U13734 (N_13734,N_5133,N_7519);
or U13735 (N_13735,N_8354,N_9996);
xor U13736 (N_13736,N_5039,N_9378);
xor U13737 (N_13737,N_8476,N_7344);
xor U13738 (N_13738,N_6409,N_9990);
xor U13739 (N_13739,N_5666,N_7341);
or U13740 (N_13740,N_7679,N_6845);
xnor U13741 (N_13741,N_9646,N_6782);
and U13742 (N_13742,N_5419,N_8323);
or U13743 (N_13743,N_5355,N_9280);
and U13744 (N_13744,N_9138,N_5457);
nor U13745 (N_13745,N_7420,N_8604);
and U13746 (N_13746,N_6792,N_5831);
or U13747 (N_13747,N_9457,N_9884);
or U13748 (N_13748,N_5947,N_7069);
nand U13749 (N_13749,N_7027,N_9350);
xor U13750 (N_13750,N_9755,N_5061);
nand U13751 (N_13751,N_6189,N_5121);
nor U13752 (N_13752,N_5877,N_7375);
xor U13753 (N_13753,N_5273,N_7954);
or U13754 (N_13754,N_8270,N_5307);
or U13755 (N_13755,N_6622,N_8134);
nor U13756 (N_13756,N_7153,N_8437);
nor U13757 (N_13757,N_5213,N_5822);
nand U13758 (N_13758,N_7401,N_7776);
nor U13759 (N_13759,N_6601,N_6918);
xor U13760 (N_13760,N_5284,N_8955);
nor U13761 (N_13761,N_9025,N_9382);
nand U13762 (N_13762,N_9335,N_5016);
xor U13763 (N_13763,N_9553,N_6418);
nor U13764 (N_13764,N_8068,N_7015);
and U13765 (N_13765,N_9121,N_9477);
or U13766 (N_13766,N_6538,N_6328);
and U13767 (N_13767,N_7153,N_5955);
xnor U13768 (N_13768,N_6194,N_9644);
nand U13769 (N_13769,N_9576,N_7658);
or U13770 (N_13770,N_9951,N_9093);
or U13771 (N_13771,N_5295,N_6049);
nor U13772 (N_13772,N_9063,N_7000);
nor U13773 (N_13773,N_8684,N_9437);
xnor U13774 (N_13774,N_7198,N_7991);
or U13775 (N_13775,N_9150,N_7533);
xnor U13776 (N_13776,N_5102,N_5931);
nand U13777 (N_13777,N_7682,N_9219);
and U13778 (N_13778,N_6693,N_6936);
nand U13779 (N_13779,N_8629,N_7234);
nand U13780 (N_13780,N_9574,N_8450);
or U13781 (N_13781,N_5256,N_7241);
xnor U13782 (N_13782,N_5026,N_6666);
and U13783 (N_13783,N_8293,N_9514);
xnor U13784 (N_13784,N_5338,N_5554);
nor U13785 (N_13785,N_5173,N_5568);
nor U13786 (N_13786,N_5845,N_6590);
nand U13787 (N_13787,N_5844,N_9610);
nor U13788 (N_13788,N_6706,N_7433);
nor U13789 (N_13789,N_6605,N_6317);
nand U13790 (N_13790,N_6449,N_5305);
nand U13791 (N_13791,N_6746,N_9987);
nand U13792 (N_13792,N_6381,N_9047);
or U13793 (N_13793,N_8780,N_7667);
and U13794 (N_13794,N_6020,N_9946);
nor U13795 (N_13795,N_6030,N_7528);
or U13796 (N_13796,N_9553,N_5037);
nor U13797 (N_13797,N_9814,N_8840);
nor U13798 (N_13798,N_7034,N_8805);
nand U13799 (N_13799,N_9105,N_5378);
and U13800 (N_13800,N_7838,N_6500);
and U13801 (N_13801,N_8901,N_6868);
nor U13802 (N_13802,N_6289,N_5072);
or U13803 (N_13803,N_9449,N_5740);
nand U13804 (N_13804,N_5751,N_8544);
or U13805 (N_13805,N_6469,N_7929);
or U13806 (N_13806,N_9743,N_9084);
and U13807 (N_13807,N_9115,N_7790);
nor U13808 (N_13808,N_6502,N_8560);
nand U13809 (N_13809,N_6802,N_9801);
and U13810 (N_13810,N_5602,N_9916);
nand U13811 (N_13811,N_8412,N_9142);
or U13812 (N_13812,N_7566,N_9719);
and U13813 (N_13813,N_9228,N_7447);
nor U13814 (N_13814,N_6775,N_8537);
and U13815 (N_13815,N_9992,N_6432);
nor U13816 (N_13816,N_8311,N_8110);
or U13817 (N_13817,N_6226,N_8892);
xnor U13818 (N_13818,N_9297,N_6471);
nor U13819 (N_13819,N_5228,N_6751);
nor U13820 (N_13820,N_6279,N_9375);
nor U13821 (N_13821,N_9676,N_9239);
nand U13822 (N_13822,N_6827,N_9496);
nor U13823 (N_13823,N_8823,N_9414);
xnor U13824 (N_13824,N_5996,N_8882);
or U13825 (N_13825,N_6793,N_6822);
and U13826 (N_13826,N_6934,N_7923);
or U13827 (N_13827,N_6033,N_6164);
nor U13828 (N_13828,N_8348,N_8786);
nor U13829 (N_13829,N_6243,N_8146);
or U13830 (N_13830,N_5103,N_6314);
nand U13831 (N_13831,N_9952,N_7192);
nand U13832 (N_13832,N_5031,N_7243);
or U13833 (N_13833,N_6271,N_8246);
or U13834 (N_13834,N_6802,N_6526);
or U13835 (N_13835,N_5035,N_8939);
or U13836 (N_13836,N_7862,N_8081);
nor U13837 (N_13837,N_8633,N_9948);
nor U13838 (N_13838,N_5191,N_7383);
xor U13839 (N_13839,N_5393,N_5609);
nand U13840 (N_13840,N_8405,N_5457);
nor U13841 (N_13841,N_8031,N_7480);
nor U13842 (N_13842,N_8244,N_9793);
and U13843 (N_13843,N_9855,N_6329);
nand U13844 (N_13844,N_7027,N_8421);
xnor U13845 (N_13845,N_5253,N_6239);
or U13846 (N_13846,N_8894,N_7223);
nand U13847 (N_13847,N_7012,N_9263);
or U13848 (N_13848,N_5653,N_7202);
xor U13849 (N_13849,N_8203,N_5823);
and U13850 (N_13850,N_6888,N_7859);
or U13851 (N_13851,N_6076,N_5745);
nor U13852 (N_13852,N_8882,N_9086);
nor U13853 (N_13853,N_5139,N_9414);
and U13854 (N_13854,N_9314,N_8898);
nand U13855 (N_13855,N_7867,N_5081);
and U13856 (N_13856,N_9160,N_5253);
or U13857 (N_13857,N_6029,N_9033);
nand U13858 (N_13858,N_9492,N_6018);
xor U13859 (N_13859,N_6765,N_6040);
xnor U13860 (N_13860,N_7886,N_6885);
xor U13861 (N_13861,N_7736,N_5614);
and U13862 (N_13862,N_5158,N_7683);
xnor U13863 (N_13863,N_9467,N_5838);
nand U13864 (N_13864,N_7571,N_5667);
and U13865 (N_13865,N_6670,N_7771);
or U13866 (N_13866,N_9976,N_6206);
nor U13867 (N_13867,N_7247,N_5953);
and U13868 (N_13868,N_8010,N_7310);
and U13869 (N_13869,N_8873,N_6662);
or U13870 (N_13870,N_6659,N_7830);
nor U13871 (N_13871,N_9288,N_5691);
xnor U13872 (N_13872,N_8868,N_8967);
or U13873 (N_13873,N_7483,N_7089);
xor U13874 (N_13874,N_5548,N_5382);
or U13875 (N_13875,N_9387,N_9350);
xor U13876 (N_13876,N_8223,N_6653);
and U13877 (N_13877,N_9496,N_9212);
and U13878 (N_13878,N_7211,N_7951);
or U13879 (N_13879,N_5017,N_8430);
nor U13880 (N_13880,N_5741,N_7150);
and U13881 (N_13881,N_7881,N_6124);
and U13882 (N_13882,N_8447,N_7238);
xnor U13883 (N_13883,N_6048,N_6292);
xnor U13884 (N_13884,N_8990,N_6744);
or U13885 (N_13885,N_5272,N_7617);
nand U13886 (N_13886,N_7356,N_5283);
nor U13887 (N_13887,N_8471,N_6941);
nor U13888 (N_13888,N_6175,N_9942);
and U13889 (N_13889,N_9916,N_9152);
or U13890 (N_13890,N_5732,N_6503);
and U13891 (N_13891,N_7051,N_9305);
nor U13892 (N_13892,N_8355,N_7717);
and U13893 (N_13893,N_7189,N_5129);
xnor U13894 (N_13894,N_7770,N_8792);
xnor U13895 (N_13895,N_8994,N_7251);
or U13896 (N_13896,N_9596,N_7880);
nand U13897 (N_13897,N_5350,N_9972);
nor U13898 (N_13898,N_7879,N_5431);
and U13899 (N_13899,N_8813,N_7843);
xnor U13900 (N_13900,N_8385,N_5384);
xnor U13901 (N_13901,N_9044,N_6811);
nor U13902 (N_13902,N_7775,N_9519);
and U13903 (N_13903,N_9138,N_9956);
and U13904 (N_13904,N_5451,N_6093);
nand U13905 (N_13905,N_6905,N_7703);
xnor U13906 (N_13906,N_8800,N_6996);
or U13907 (N_13907,N_6365,N_6032);
nand U13908 (N_13908,N_7314,N_6921);
xnor U13909 (N_13909,N_8048,N_8339);
nor U13910 (N_13910,N_7985,N_6164);
or U13911 (N_13911,N_5327,N_5891);
or U13912 (N_13912,N_9906,N_9536);
nor U13913 (N_13913,N_5313,N_6469);
and U13914 (N_13914,N_8796,N_5433);
xnor U13915 (N_13915,N_9539,N_7228);
nor U13916 (N_13916,N_6699,N_8034);
and U13917 (N_13917,N_7772,N_6752);
or U13918 (N_13918,N_6152,N_6058);
nor U13919 (N_13919,N_7140,N_9069);
and U13920 (N_13920,N_6815,N_8384);
or U13921 (N_13921,N_8972,N_5230);
or U13922 (N_13922,N_6534,N_7939);
and U13923 (N_13923,N_8324,N_6286);
nor U13924 (N_13924,N_8219,N_8569);
xnor U13925 (N_13925,N_5003,N_5706);
nand U13926 (N_13926,N_6330,N_8202);
and U13927 (N_13927,N_6143,N_5458);
nor U13928 (N_13928,N_6312,N_8041);
xnor U13929 (N_13929,N_9568,N_5384);
nand U13930 (N_13930,N_6822,N_6259);
and U13931 (N_13931,N_8733,N_6038);
nor U13932 (N_13932,N_5153,N_5352);
and U13933 (N_13933,N_8210,N_7985);
nor U13934 (N_13934,N_7181,N_9177);
and U13935 (N_13935,N_5066,N_9725);
and U13936 (N_13936,N_9107,N_6444);
nand U13937 (N_13937,N_5647,N_5688);
nor U13938 (N_13938,N_9452,N_5225);
xor U13939 (N_13939,N_8625,N_9546);
nor U13940 (N_13940,N_6522,N_9535);
nor U13941 (N_13941,N_9546,N_7534);
nand U13942 (N_13942,N_9167,N_5535);
nor U13943 (N_13943,N_7837,N_5957);
nor U13944 (N_13944,N_9179,N_9866);
and U13945 (N_13945,N_7615,N_7115);
and U13946 (N_13946,N_5985,N_6216);
or U13947 (N_13947,N_5871,N_5730);
nand U13948 (N_13948,N_9800,N_5719);
xnor U13949 (N_13949,N_6800,N_5627);
xnor U13950 (N_13950,N_8078,N_6989);
and U13951 (N_13951,N_5533,N_7503);
nor U13952 (N_13952,N_5458,N_9533);
or U13953 (N_13953,N_6980,N_8835);
or U13954 (N_13954,N_6391,N_9337);
and U13955 (N_13955,N_8465,N_5486);
nand U13956 (N_13956,N_5962,N_9272);
and U13957 (N_13957,N_5606,N_6679);
nand U13958 (N_13958,N_8566,N_9971);
and U13959 (N_13959,N_7507,N_8706);
and U13960 (N_13960,N_8348,N_9243);
nand U13961 (N_13961,N_5229,N_5362);
or U13962 (N_13962,N_8082,N_9091);
and U13963 (N_13963,N_9068,N_7743);
xnor U13964 (N_13964,N_9284,N_8880);
nand U13965 (N_13965,N_6575,N_6100);
or U13966 (N_13966,N_9867,N_9837);
xor U13967 (N_13967,N_8412,N_9552);
nand U13968 (N_13968,N_6469,N_9088);
or U13969 (N_13969,N_8177,N_5949);
xnor U13970 (N_13970,N_9230,N_5310);
xor U13971 (N_13971,N_9511,N_5232);
nand U13972 (N_13972,N_7455,N_5471);
or U13973 (N_13973,N_8615,N_7155);
nand U13974 (N_13974,N_5100,N_5553);
nor U13975 (N_13975,N_7514,N_6689);
nor U13976 (N_13976,N_7805,N_9341);
and U13977 (N_13977,N_8913,N_9399);
xnor U13978 (N_13978,N_6883,N_9638);
and U13979 (N_13979,N_7374,N_6728);
or U13980 (N_13980,N_5369,N_5003);
nand U13981 (N_13981,N_8928,N_6227);
xnor U13982 (N_13982,N_8244,N_9938);
and U13983 (N_13983,N_9259,N_6916);
or U13984 (N_13984,N_6824,N_5628);
xnor U13985 (N_13985,N_5510,N_9584);
or U13986 (N_13986,N_9351,N_6737);
nor U13987 (N_13987,N_9533,N_6344);
xnor U13988 (N_13988,N_9517,N_9031);
or U13989 (N_13989,N_6788,N_8402);
or U13990 (N_13990,N_5450,N_9028);
nor U13991 (N_13991,N_6075,N_5817);
nor U13992 (N_13992,N_7740,N_8283);
and U13993 (N_13993,N_5199,N_5106);
and U13994 (N_13994,N_5600,N_6942);
or U13995 (N_13995,N_7101,N_8898);
nor U13996 (N_13996,N_5327,N_6159);
nor U13997 (N_13997,N_7885,N_8538);
xnor U13998 (N_13998,N_7650,N_5410);
nand U13999 (N_13999,N_8351,N_7075);
nor U14000 (N_14000,N_5052,N_5586);
xnor U14001 (N_14001,N_8178,N_7761);
nand U14002 (N_14002,N_6937,N_7885);
xor U14003 (N_14003,N_8533,N_8346);
or U14004 (N_14004,N_9266,N_9636);
and U14005 (N_14005,N_5941,N_8794);
and U14006 (N_14006,N_6272,N_8204);
or U14007 (N_14007,N_8084,N_5952);
nor U14008 (N_14008,N_6706,N_8316);
or U14009 (N_14009,N_6805,N_7174);
or U14010 (N_14010,N_7007,N_7068);
and U14011 (N_14011,N_6681,N_8275);
nor U14012 (N_14012,N_5048,N_5024);
nand U14013 (N_14013,N_9186,N_5391);
or U14014 (N_14014,N_8755,N_7291);
nor U14015 (N_14015,N_9028,N_8295);
and U14016 (N_14016,N_9501,N_9392);
xor U14017 (N_14017,N_7230,N_7888);
and U14018 (N_14018,N_7154,N_9284);
or U14019 (N_14019,N_5130,N_9520);
nand U14020 (N_14020,N_9245,N_6966);
and U14021 (N_14021,N_8106,N_6874);
nand U14022 (N_14022,N_6954,N_5102);
xnor U14023 (N_14023,N_7412,N_7460);
and U14024 (N_14024,N_8336,N_9155);
xnor U14025 (N_14025,N_7930,N_6923);
xnor U14026 (N_14026,N_6221,N_7763);
nand U14027 (N_14027,N_7471,N_6610);
nor U14028 (N_14028,N_9311,N_5382);
and U14029 (N_14029,N_8458,N_5996);
and U14030 (N_14030,N_6492,N_6623);
xnor U14031 (N_14031,N_9165,N_6129);
and U14032 (N_14032,N_8948,N_9582);
and U14033 (N_14033,N_6581,N_5114);
or U14034 (N_14034,N_8476,N_6077);
nand U14035 (N_14035,N_6190,N_5685);
nor U14036 (N_14036,N_9707,N_9095);
and U14037 (N_14037,N_9196,N_9947);
xor U14038 (N_14038,N_5037,N_5565);
and U14039 (N_14039,N_8886,N_9726);
nor U14040 (N_14040,N_9823,N_8912);
nand U14041 (N_14041,N_6005,N_9257);
nand U14042 (N_14042,N_7006,N_7026);
or U14043 (N_14043,N_8188,N_6810);
and U14044 (N_14044,N_5438,N_7597);
nor U14045 (N_14045,N_9599,N_9670);
or U14046 (N_14046,N_5120,N_5988);
xnor U14047 (N_14047,N_9061,N_8704);
nand U14048 (N_14048,N_6851,N_9777);
nor U14049 (N_14049,N_8204,N_7865);
and U14050 (N_14050,N_6707,N_8168);
xnor U14051 (N_14051,N_5069,N_9307);
nor U14052 (N_14052,N_7995,N_7867);
and U14053 (N_14053,N_5680,N_7210);
or U14054 (N_14054,N_9708,N_8926);
nor U14055 (N_14055,N_6939,N_7523);
nand U14056 (N_14056,N_6546,N_5489);
and U14057 (N_14057,N_6531,N_5694);
and U14058 (N_14058,N_6774,N_9534);
xnor U14059 (N_14059,N_5586,N_9282);
and U14060 (N_14060,N_8552,N_6199);
xor U14061 (N_14061,N_7864,N_7725);
or U14062 (N_14062,N_6605,N_7489);
nand U14063 (N_14063,N_7966,N_9762);
nand U14064 (N_14064,N_9662,N_9778);
and U14065 (N_14065,N_5957,N_8068);
nor U14066 (N_14066,N_7296,N_8941);
nor U14067 (N_14067,N_7523,N_6093);
nand U14068 (N_14068,N_5448,N_5585);
and U14069 (N_14069,N_5827,N_6407);
nand U14070 (N_14070,N_8574,N_5116);
or U14071 (N_14071,N_7064,N_5916);
or U14072 (N_14072,N_9728,N_6363);
nand U14073 (N_14073,N_8371,N_6947);
and U14074 (N_14074,N_6446,N_5947);
nor U14075 (N_14075,N_7597,N_7757);
xor U14076 (N_14076,N_5245,N_8436);
or U14077 (N_14077,N_7679,N_6678);
or U14078 (N_14078,N_9451,N_9956);
or U14079 (N_14079,N_8500,N_5583);
or U14080 (N_14080,N_7049,N_9595);
or U14081 (N_14081,N_5337,N_8010);
or U14082 (N_14082,N_5402,N_8295);
xor U14083 (N_14083,N_7419,N_5839);
and U14084 (N_14084,N_5802,N_6375);
and U14085 (N_14085,N_6473,N_7749);
nand U14086 (N_14086,N_5210,N_8333);
xor U14087 (N_14087,N_6844,N_9948);
xor U14088 (N_14088,N_5970,N_9799);
and U14089 (N_14089,N_7269,N_9479);
nor U14090 (N_14090,N_9751,N_8792);
or U14091 (N_14091,N_8817,N_5119);
xnor U14092 (N_14092,N_6153,N_5818);
and U14093 (N_14093,N_8506,N_5563);
nand U14094 (N_14094,N_6951,N_5540);
nor U14095 (N_14095,N_8275,N_6838);
nand U14096 (N_14096,N_8242,N_6075);
xnor U14097 (N_14097,N_6988,N_7261);
nor U14098 (N_14098,N_8120,N_8779);
nor U14099 (N_14099,N_5690,N_8790);
nor U14100 (N_14100,N_7283,N_5545);
nor U14101 (N_14101,N_7967,N_5133);
xor U14102 (N_14102,N_7099,N_7353);
and U14103 (N_14103,N_7466,N_8786);
and U14104 (N_14104,N_5370,N_8048);
or U14105 (N_14105,N_8262,N_6041);
xor U14106 (N_14106,N_5792,N_6863);
or U14107 (N_14107,N_7681,N_5671);
or U14108 (N_14108,N_7342,N_7005);
and U14109 (N_14109,N_8854,N_8578);
or U14110 (N_14110,N_6079,N_9518);
nand U14111 (N_14111,N_5996,N_5028);
and U14112 (N_14112,N_6594,N_7871);
nor U14113 (N_14113,N_5019,N_6490);
nand U14114 (N_14114,N_7269,N_8744);
nand U14115 (N_14115,N_5734,N_6731);
or U14116 (N_14116,N_8027,N_8756);
or U14117 (N_14117,N_7487,N_5484);
nand U14118 (N_14118,N_8242,N_7525);
or U14119 (N_14119,N_5140,N_6491);
xor U14120 (N_14120,N_5035,N_7430);
and U14121 (N_14121,N_9069,N_9081);
and U14122 (N_14122,N_8197,N_5517);
and U14123 (N_14123,N_6107,N_6933);
nand U14124 (N_14124,N_9913,N_8249);
xor U14125 (N_14125,N_5199,N_5213);
or U14126 (N_14126,N_9559,N_8282);
or U14127 (N_14127,N_5270,N_5778);
nor U14128 (N_14128,N_6537,N_6267);
nand U14129 (N_14129,N_5197,N_7628);
xnor U14130 (N_14130,N_8021,N_8900);
nand U14131 (N_14131,N_5152,N_5858);
nor U14132 (N_14132,N_8819,N_6097);
or U14133 (N_14133,N_5811,N_7067);
nand U14134 (N_14134,N_7274,N_8797);
and U14135 (N_14135,N_6994,N_9260);
nor U14136 (N_14136,N_5471,N_5043);
xor U14137 (N_14137,N_8075,N_5374);
or U14138 (N_14138,N_7992,N_9849);
nor U14139 (N_14139,N_6338,N_9577);
and U14140 (N_14140,N_6008,N_8255);
xor U14141 (N_14141,N_9795,N_6215);
nor U14142 (N_14142,N_9111,N_5770);
and U14143 (N_14143,N_9191,N_8604);
and U14144 (N_14144,N_6229,N_5720);
or U14145 (N_14145,N_8217,N_7749);
nand U14146 (N_14146,N_6494,N_8389);
xnor U14147 (N_14147,N_9915,N_9794);
or U14148 (N_14148,N_6816,N_9146);
or U14149 (N_14149,N_7863,N_9803);
nand U14150 (N_14150,N_8303,N_8081);
xor U14151 (N_14151,N_5471,N_5831);
and U14152 (N_14152,N_9854,N_9076);
or U14153 (N_14153,N_5927,N_5656);
and U14154 (N_14154,N_7516,N_9385);
and U14155 (N_14155,N_6473,N_9698);
and U14156 (N_14156,N_8909,N_8555);
and U14157 (N_14157,N_6164,N_5619);
nand U14158 (N_14158,N_7455,N_7096);
nor U14159 (N_14159,N_9849,N_5080);
nand U14160 (N_14160,N_8457,N_5310);
xor U14161 (N_14161,N_9051,N_7468);
xnor U14162 (N_14162,N_6034,N_8288);
xor U14163 (N_14163,N_9579,N_7465);
nand U14164 (N_14164,N_6313,N_9049);
xor U14165 (N_14165,N_8579,N_7657);
and U14166 (N_14166,N_7435,N_8836);
nor U14167 (N_14167,N_6971,N_7810);
nand U14168 (N_14168,N_8834,N_6010);
nand U14169 (N_14169,N_5954,N_8017);
nand U14170 (N_14170,N_6229,N_9321);
or U14171 (N_14171,N_5889,N_8988);
nor U14172 (N_14172,N_7462,N_9060);
or U14173 (N_14173,N_7599,N_8076);
or U14174 (N_14174,N_5840,N_6741);
nor U14175 (N_14175,N_6707,N_7323);
nand U14176 (N_14176,N_5170,N_5436);
or U14177 (N_14177,N_5909,N_7191);
nor U14178 (N_14178,N_5545,N_5190);
and U14179 (N_14179,N_8192,N_7893);
xor U14180 (N_14180,N_8564,N_6850);
nand U14181 (N_14181,N_5203,N_9680);
or U14182 (N_14182,N_5038,N_5932);
nand U14183 (N_14183,N_5660,N_7097);
or U14184 (N_14184,N_7902,N_6231);
and U14185 (N_14185,N_9924,N_8042);
and U14186 (N_14186,N_6931,N_5973);
and U14187 (N_14187,N_5400,N_7202);
and U14188 (N_14188,N_7177,N_5001);
nand U14189 (N_14189,N_7504,N_6788);
nor U14190 (N_14190,N_6186,N_9969);
xnor U14191 (N_14191,N_6764,N_7161);
xnor U14192 (N_14192,N_5066,N_5838);
nor U14193 (N_14193,N_5522,N_5630);
and U14194 (N_14194,N_8567,N_8286);
xor U14195 (N_14195,N_8229,N_5603);
xor U14196 (N_14196,N_5563,N_7710);
xnor U14197 (N_14197,N_9598,N_8903);
nor U14198 (N_14198,N_7231,N_6792);
and U14199 (N_14199,N_8419,N_9305);
and U14200 (N_14200,N_8983,N_9541);
xor U14201 (N_14201,N_5832,N_6467);
and U14202 (N_14202,N_6192,N_8554);
nor U14203 (N_14203,N_9878,N_5719);
or U14204 (N_14204,N_7640,N_8092);
nand U14205 (N_14205,N_8035,N_7232);
nand U14206 (N_14206,N_8313,N_7947);
nand U14207 (N_14207,N_8538,N_7271);
and U14208 (N_14208,N_9589,N_9890);
and U14209 (N_14209,N_9067,N_7411);
nand U14210 (N_14210,N_5302,N_5872);
or U14211 (N_14211,N_8978,N_9918);
xor U14212 (N_14212,N_6832,N_6584);
nor U14213 (N_14213,N_6216,N_7234);
xor U14214 (N_14214,N_6187,N_6159);
and U14215 (N_14215,N_9194,N_5225);
nor U14216 (N_14216,N_5411,N_6549);
nor U14217 (N_14217,N_7471,N_6037);
nand U14218 (N_14218,N_9929,N_6607);
and U14219 (N_14219,N_9641,N_6520);
nor U14220 (N_14220,N_8071,N_8128);
and U14221 (N_14221,N_7675,N_8624);
nor U14222 (N_14222,N_8688,N_6514);
nor U14223 (N_14223,N_5757,N_7623);
and U14224 (N_14224,N_8542,N_8830);
or U14225 (N_14225,N_7004,N_9635);
nor U14226 (N_14226,N_7040,N_6358);
or U14227 (N_14227,N_7922,N_5778);
or U14228 (N_14228,N_9293,N_5338);
nor U14229 (N_14229,N_8025,N_7751);
nor U14230 (N_14230,N_8744,N_6936);
nor U14231 (N_14231,N_6986,N_8366);
nand U14232 (N_14232,N_8065,N_7564);
and U14233 (N_14233,N_9979,N_7192);
nand U14234 (N_14234,N_5817,N_9608);
nand U14235 (N_14235,N_6596,N_9657);
nor U14236 (N_14236,N_7317,N_9256);
nor U14237 (N_14237,N_8374,N_7993);
or U14238 (N_14238,N_6527,N_8703);
or U14239 (N_14239,N_7009,N_8648);
nand U14240 (N_14240,N_9209,N_7001);
and U14241 (N_14241,N_5357,N_5093);
nor U14242 (N_14242,N_5457,N_6374);
and U14243 (N_14243,N_9138,N_6074);
nand U14244 (N_14244,N_8094,N_7848);
xor U14245 (N_14245,N_8188,N_7297);
xor U14246 (N_14246,N_6020,N_5461);
nand U14247 (N_14247,N_9566,N_7319);
nor U14248 (N_14248,N_7779,N_7303);
and U14249 (N_14249,N_7770,N_5211);
nor U14250 (N_14250,N_5481,N_6930);
and U14251 (N_14251,N_9728,N_6204);
xor U14252 (N_14252,N_5299,N_7567);
nor U14253 (N_14253,N_9394,N_5296);
and U14254 (N_14254,N_9269,N_6312);
nor U14255 (N_14255,N_5237,N_8849);
and U14256 (N_14256,N_9102,N_9641);
xnor U14257 (N_14257,N_6139,N_5336);
nand U14258 (N_14258,N_8566,N_9695);
or U14259 (N_14259,N_6287,N_6427);
or U14260 (N_14260,N_5644,N_8045);
xor U14261 (N_14261,N_6651,N_8907);
or U14262 (N_14262,N_7474,N_9606);
xnor U14263 (N_14263,N_7628,N_5547);
or U14264 (N_14264,N_8936,N_9708);
nor U14265 (N_14265,N_5468,N_5326);
nor U14266 (N_14266,N_7490,N_9497);
and U14267 (N_14267,N_7918,N_6220);
or U14268 (N_14268,N_5216,N_7977);
xor U14269 (N_14269,N_9213,N_9537);
and U14270 (N_14270,N_5069,N_8819);
xor U14271 (N_14271,N_8879,N_9258);
xor U14272 (N_14272,N_7901,N_7075);
nor U14273 (N_14273,N_7733,N_7465);
or U14274 (N_14274,N_6467,N_7210);
nor U14275 (N_14275,N_8167,N_9836);
xor U14276 (N_14276,N_8842,N_6435);
and U14277 (N_14277,N_6239,N_6038);
or U14278 (N_14278,N_7867,N_7993);
nor U14279 (N_14279,N_5782,N_9901);
nand U14280 (N_14280,N_6551,N_5688);
nor U14281 (N_14281,N_7959,N_9998);
xor U14282 (N_14282,N_9685,N_8710);
and U14283 (N_14283,N_8690,N_8657);
nor U14284 (N_14284,N_6157,N_5771);
or U14285 (N_14285,N_8658,N_6995);
nand U14286 (N_14286,N_8542,N_7171);
nor U14287 (N_14287,N_7358,N_7574);
and U14288 (N_14288,N_5077,N_7067);
and U14289 (N_14289,N_5607,N_5020);
nor U14290 (N_14290,N_7562,N_9067);
or U14291 (N_14291,N_9488,N_8170);
or U14292 (N_14292,N_6861,N_9961);
and U14293 (N_14293,N_8134,N_6619);
xnor U14294 (N_14294,N_9456,N_7303);
and U14295 (N_14295,N_8942,N_8556);
nand U14296 (N_14296,N_6088,N_9893);
and U14297 (N_14297,N_6671,N_6431);
nand U14298 (N_14298,N_5380,N_5868);
or U14299 (N_14299,N_8067,N_5050);
nand U14300 (N_14300,N_6753,N_7109);
and U14301 (N_14301,N_6546,N_9972);
nor U14302 (N_14302,N_7182,N_5062);
nand U14303 (N_14303,N_6013,N_8800);
nand U14304 (N_14304,N_6742,N_9679);
xor U14305 (N_14305,N_7185,N_9011);
nand U14306 (N_14306,N_8065,N_9732);
and U14307 (N_14307,N_6776,N_8796);
and U14308 (N_14308,N_8532,N_5453);
and U14309 (N_14309,N_5622,N_5487);
xor U14310 (N_14310,N_6245,N_8844);
nand U14311 (N_14311,N_8830,N_6995);
or U14312 (N_14312,N_7695,N_9937);
nand U14313 (N_14313,N_9916,N_8057);
xnor U14314 (N_14314,N_9811,N_9633);
xnor U14315 (N_14315,N_5438,N_6647);
nor U14316 (N_14316,N_6518,N_9052);
nor U14317 (N_14317,N_9610,N_9907);
xor U14318 (N_14318,N_9457,N_5146);
nor U14319 (N_14319,N_5661,N_5813);
xnor U14320 (N_14320,N_9356,N_5269);
or U14321 (N_14321,N_6542,N_9823);
and U14322 (N_14322,N_5137,N_5706);
or U14323 (N_14323,N_9604,N_5345);
or U14324 (N_14324,N_9373,N_9197);
nand U14325 (N_14325,N_9206,N_9237);
nor U14326 (N_14326,N_7966,N_9670);
nor U14327 (N_14327,N_8388,N_7464);
nor U14328 (N_14328,N_5679,N_8420);
and U14329 (N_14329,N_7291,N_5920);
nor U14330 (N_14330,N_7765,N_8316);
nand U14331 (N_14331,N_7099,N_9981);
nand U14332 (N_14332,N_6320,N_6001);
or U14333 (N_14333,N_9252,N_7821);
nand U14334 (N_14334,N_9069,N_9650);
nand U14335 (N_14335,N_7564,N_7221);
nor U14336 (N_14336,N_6556,N_5740);
or U14337 (N_14337,N_5633,N_9779);
or U14338 (N_14338,N_5149,N_7649);
or U14339 (N_14339,N_5883,N_8952);
and U14340 (N_14340,N_5759,N_9222);
nor U14341 (N_14341,N_7563,N_9655);
or U14342 (N_14342,N_7756,N_6268);
nor U14343 (N_14343,N_6184,N_6255);
xor U14344 (N_14344,N_5824,N_5697);
and U14345 (N_14345,N_8127,N_8134);
nand U14346 (N_14346,N_6921,N_7877);
and U14347 (N_14347,N_5760,N_7497);
and U14348 (N_14348,N_5558,N_6893);
nand U14349 (N_14349,N_5430,N_7425);
and U14350 (N_14350,N_9359,N_5746);
nor U14351 (N_14351,N_8118,N_6169);
or U14352 (N_14352,N_8546,N_5057);
xor U14353 (N_14353,N_6795,N_8693);
nor U14354 (N_14354,N_7278,N_8248);
nor U14355 (N_14355,N_6660,N_6716);
or U14356 (N_14356,N_5869,N_9961);
nand U14357 (N_14357,N_7452,N_7992);
xor U14358 (N_14358,N_5716,N_9817);
xnor U14359 (N_14359,N_7023,N_8805);
nor U14360 (N_14360,N_8814,N_6528);
nor U14361 (N_14361,N_6799,N_9024);
nor U14362 (N_14362,N_8153,N_6473);
or U14363 (N_14363,N_7322,N_9725);
and U14364 (N_14364,N_8003,N_7789);
and U14365 (N_14365,N_6256,N_6942);
nand U14366 (N_14366,N_7041,N_9154);
nand U14367 (N_14367,N_8465,N_8749);
xor U14368 (N_14368,N_5380,N_8163);
nand U14369 (N_14369,N_7536,N_5016);
or U14370 (N_14370,N_9698,N_8290);
nand U14371 (N_14371,N_7768,N_6960);
nand U14372 (N_14372,N_5460,N_9010);
xnor U14373 (N_14373,N_9478,N_8449);
or U14374 (N_14374,N_5199,N_9980);
and U14375 (N_14375,N_8033,N_6496);
nor U14376 (N_14376,N_9203,N_6782);
nand U14377 (N_14377,N_9673,N_8638);
xor U14378 (N_14378,N_7841,N_8611);
xnor U14379 (N_14379,N_9456,N_5821);
or U14380 (N_14380,N_5083,N_5048);
or U14381 (N_14381,N_6181,N_9831);
xnor U14382 (N_14382,N_7198,N_8475);
nand U14383 (N_14383,N_9481,N_9048);
nand U14384 (N_14384,N_9030,N_5168);
nand U14385 (N_14385,N_6333,N_7647);
xor U14386 (N_14386,N_9882,N_7983);
and U14387 (N_14387,N_7416,N_5901);
xnor U14388 (N_14388,N_9865,N_6730);
xnor U14389 (N_14389,N_9958,N_8612);
xnor U14390 (N_14390,N_8051,N_7325);
nand U14391 (N_14391,N_6062,N_9278);
xor U14392 (N_14392,N_9913,N_7644);
nor U14393 (N_14393,N_5483,N_5014);
xor U14394 (N_14394,N_6340,N_9026);
or U14395 (N_14395,N_8048,N_7773);
and U14396 (N_14396,N_5359,N_5890);
nand U14397 (N_14397,N_8952,N_9735);
or U14398 (N_14398,N_7782,N_5609);
or U14399 (N_14399,N_8416,N_7309);
nand U14400 (N_14400,N_6255,N_5787);
nand U14401 (N_14401,N_7644,N_8745);
and U14402 (N_14402,N_7879,N_5497);
nand U14403 (N_14403,N_6330,N_6798);
xor U14404 (N_14404,N_7378,N_6030);
nand U14405 (N_14405,N_5041,N_7610);
and U14406 (N_14406,N_9706,N_9222);
or U14407 (N_14407,N_6754,N_5301);
nor U14408 (N_14408,N_7101,N_5183);
nor U14409 (N_14409,N_9882,N_9090);
or U14410 (N_14410,N_8540,N_9928);
or U14411 (N_14411,N_8967,N_9709);
nand U14412 (N_14412,N_7442,N_9467);
and U14413 (N_14413,N_5215,N_7902);
nand U14414 (N_14414,N_6651,N_7509);
nand U14415 (N_14415,N_9325,N_5721);
xor U14416 (N_14416,N_7086,N_5804);
or U14417 (N_14417,N_8917,N_9198);
nand U14418 (N_14418,N_5187,N_6646);
nand U14419 (N_14419,N_9236,N_6367);
nand U14420 (N_14420,N_6919,N_5206);
nor U14421 (N_14421,N_8154,N_7022);
or U14422 (N_14422,N_7452,N_8907);
or U14423 (N_14423,N_9687,N_8408);
and U14424 (N_14424,N_9852,N_9672);
nor U14425 (N_14425,N_8043,N_7202);
nor U14426 (N_14426,N_6190,N_6251);
or U14427 (N_14427,N_6196,N_7715);
xor U14428 (N_14428,N_5390,N_5558);
nand U14429 (N_14429,N_8938,N_9896);
nand U14430 (N_14430,N_5460,N_7299);
nand U14431 (N_14431,N_7495,N_7870);
and U14432 (N_14432,N_9892,N_7352);
or U14433 (N_14433,N_9338,N_5096);
and U14434 (N_14434,N_9239,N_9098);
and U14435 (N_14435,N_9925,N_6465);
nor U14436 (N_14436,N_5549,N_8778);
or U14437 (N_14437,N_6240,N_7234);
nor U14438 (N_14438,N_5069,N_5312);
or U14439 (N_14439,N_9415,N_8088);
nor U14440 (N_14440,N_5579,N_7543);
xor U14441 (N_14441,N_6607,N_5624);
nor U14442 (N_14442,N_5941,N_6528);
nand U14443 (N_14443,N_8294,N_9815);
or U14444 (N_14444,N_5309,N_7727);
xnor U14445 (N_14445,N_8432,N_9062);
or U14446 (N_14446,N_6914,N_5981);
nor U14447 (N_14447,N_8861,N_9514);
nand U14448 (N_14448,N_8040,N_9718);
nor U14449 (N_14449,N_8999,N_8496);
or U14450 (N_14450,N_9947,N_9814);
nand U14451 (N_14451,N_9850,N_8205);
and U14452 (N_14452,N_7650,N_7383);
nand U14453 (N_14453,N_8986,N_9000);
xor U14454 (N_14454,N_9362,N_7636);
and U14455 (N_14455,N_6937,N_8363);
and U14456 (N_14456,N_5256,N_8498);
xor U14457 (N_14457,N_5352,N_5900);
and U14458 (N_14458,N_5582,N_5727);
and U14459 (N_14459,N_5196,N_8834);
nand U14460 (N_14460,N_8868,N_7386);
xor U14461 (N_14461,N_8877,N_7402);
xnor U14462 (N_14462,N_6967,N_9587);
or U14463 (N_14463,N_7691,N_5183);
and U14464 (N_14464,N_7563,N_8173);
nand U14465 (N_14465,N_5526,N_8396);
or U14466 (N_14466,N_8304,N_9853);
xor U14467 (N_14467,N_5662,N_5522);
nand U14468 (N_14468,N_7129,N_9658);
and U14469 (N_14469,N_9377,N_9490);
or U14470 (N_14470,N_9296,N_6230);
nor U14471 (N_14471,N_8880,N_7347);
xnor U14472 (N_14472,N_9375,N_9747);
xnor U14473 (N_14473,N_8060,N_7233);
and U14474 (N_14474,N_7666,N_6408);
or U14475 (N_14475,N_7382,N_8923);
nand U14476 (N_14476,N_6832,N_8308);
and U14477 (N_14477,N_9483,N_9104);
nand U14478 (N_14478,N_5428,N_8174);
xor U14479 (N_14479,N_7081,N_6947);
and U14480 (N_14480,N_9579,N_9718);
and U14481 (N_14481,N_6356,N_9164);
and U14482 (N_14482,N_9658,N_9971);
nand U14483 (N_14483,N_8404,N_8270);
nand U14484 (N_14484,N_6557,N_8829);
and U14485 (N_14485,N_7062,N_9669);
and U14486 (N_14486,N_9660,N_9561);
xor U14487 (N_14487,N_6145,N_6498);
nand U14488 (N_14488,N_5369,N_7506);
nor U14489 (N_14489,N_5019,N_6766);
nand U14490 (N_14490,N_8943,N_8986);
and U14491 (N_14491,N_7538,N_6909);
nand U14492 (N_14492,N_8654,N_8022);
and U14493 (N_14493,N_5783,N_7741);
xnor U14494 (N_14494,N_8459,N_7953);
nor U14495 (N_14495,N_9180,N_8242);
nand U14496 (N_14496,N_7475,N_7818);
or U14497 (N_14497,N_5621,N_6031);
nand U14498 (N_14498,N_7949,N_7989);
xnor U14499 (N_14499,N_7550,N_9334);
and U14500 (N_14500,N_8269,N_5713);
nor U14501 (N_14501,N_6739,N_9165);
or U14502 (N_14502,N_8646,N_6388);
or U14503 (N_14503,N_5599,N_9651);
nor U14504 (N_14504,N_8499,N_5073);
nor U14505 (N_14505,N_9253,N_6081);
and U14506 (N_14506,N_5216,N_6040);
or U14507 (N_14507,N_8960,N_7974);
and U14508 (N_14508,N_8044,N_5988);
or U14509 (N_14509,N_7930,N_8780);
xnor U14510 (N_14510,N_7605,N_8373);
and U14511 (N_14511,N_5753,N_5917);
or U14512 (N_14512,N_5767,N_7271);
and U14513 (N_14513,N_5947,N_8546);
nor U14514 (N_14514,N_5485,N_5121);
or U14515 (N_14515,N_5953,N_9162);
nand U14516 (N_14516,N_6311,N_8048);
nor U14517 (N_14517,N_8545,N_9500);
nand U14518 (N_14518,N_8125,N_5485);
or U14519 (N_14519,N_5092,N_6980);
nand U14520 (N_14520,N_5493,N_5492);
or U14521 (N_14521,N_6382,N_9756);
nand U14522 (N_14522,N_5398,N_8082);
nand U14523 (N_14523,N_5081,N_7900);
xnor U14524 (N_14524,N_5767,N_7096);
nor U14525 (N_14525,N_9311,N_9701);
nor U14526 (N_14526,N_6662,N_8030);
nor U14527 (N_14527,N_6874,N_7576);
nand U14528 (N_14528,N_9478,N_8328);
nor U14529 (N_14529,N_6757,N_5875);
nor U14530 (N_14530,N_8231,N_8544);
nor U14531 (N_14531,N_5262,N_6710);
nand U14532 (N_14532,N_6845,N_9649);
or U14533 (N_14533,N_7502,N_6812);
xor U14534 (N_14534,N_5357,N_6774);
xnor U14535 (N_14535,N_9265,N_8660);
xor U14536 (N_14536,N_6484,N_8045);
and U14537 (N_14537,N_5592,N_9010);
xor U14538 (N_14538,N_7404,N_6491);
nor U14539 (N_14539,N_9403,N_5677);
nand U14540 (N_14540,N_9103,N_5848);
nand U14541 (N_14541,N_9929,N_6816);
or U14542 (N_14542,N_6768,N_8755);
or U14543 (N_14543,N_7323,N_7825);
xor U14544 (N_14544,N_7661,N_6781);
xor U14545 (N_14545,N_6367,N_5818);
nor U14546 (N_14546,N_9273,N_8652);
and U14547 (N_14547,N_5651,N_6055);
nand U14548 (N_14548,N_5978,N_6957);
xor U14549 (N_14549,N_8560,N_5439);
and U14550 (N_14550,N_7652,N_6417);
nor U14551 (N_14551,N_5202,N_7206);
nor U14552 (N_14552,N_7189,N_7238);
nor U14553 (N_14553,N_6375,N_5997);
and U14554 (N_14554,N_5939,N_7118);
nand U14555 (N_14555,N_8037,N_5319);
and U14556 (N_14556,N_8805,N_9542);
nand U14557 (N_14557,N_6152,N_6979);
and U14558 (N_14558,N_5618,N_8876);
nor U14559 (N_14559,N_6418,N_7404);
xnor U14560 (N_14560,N_7847,N_5584);
xnor U14561 (N_14561,N_7506,N_7720);
or U14562 (N_14562,N_5740,N_8452);
and U14563 (N_14563,N_8346,N_6300);
or U14564 (N_14564,N_8235,N_5631);
and U14565 (N_14565,N_7594,N_5874);
nand U14566 (N_14566,N_5626,N_5308);
nand U14567 (N_14567,N_7192,N_6565);
xnor U14568 (N_14568,N_8863,N_5532);
or U14569 (N_14569,N_5900,N_9373);
and U14570 (N_14570,N_6521,N_8540);
xor U14571 (N_14571,N_7184,N_6853);
xnor U14572 (N_14572,N_8929,N_9545);
nand U14573 (N_14573,N_5191,N_9366);
nand U14574 (N_14574,N_8978,N_9515);
nor U14575 (N_14575,N_8611,N_5559);
nor U14576 (N_14576,N_8700,N_9706);
or U14577 (N_14577,N_8987,N_9571);
xor U14578 (N_14578,N_7531,N_9286);
nand U14579 (N_14579,N_8198,N_6275);
nand U14580 (N_14580,N_9477,N_7869);
or U14581 (N_14581,N_7196,N_8530);
or U14582 (N_14582,N_9287,N_8186);
xor U14583 (N_14583,N_5313,N_8114);
nor U14584 (N_14584,N_8098,N_6262);
nand U14585 (N_14585,N_5659,N_5217);
nor U14586 (N_14586,N_8559,N_5811);
xor U14587 (N_14587,N_8937,N_9150);
nor U14588 (N_14588,N_8090,N_9186);
or U14589 (N_14589,N_9205,N_7980);
and U14590 (N_14590,N_5670,N_8230);
nand U14591 (N_14591,N_9355,N_6864);
xor U14592 (N_14592,N_9844,N_6099);
or U14593 (N_14593,N_5102,N_7301);
nor U14594 (N_14594,N_7443,N_9530);
and U14595 (N_14595,N_5258,N_9512);
or U14596 (N_14596,N_8729,N_7002);
nand U14597 (N_14597,N_5831,N_6848);
or U14598 (N_14598,N_7232,N_5443);
xnor U14599 (N_14599,N_8171,N_8605);
xnor U14600 (N_14600,N_6285,N_9370);
nand U14601 (N_14601,N_5473,N_9910);
and U14602 (N_14602,N_8180,N_7133);
and U14603 (N_14603,N_8036,N_5828);
or U14604 (N_14604,N_6259,N_6345);
nand U14605 (N_14605,N_8619,N_7780);
and U14606 (N_14606,N_9041,N_7785);
or U14607 (N_14607,N_8167,N_8328);
and U14608 (N_14608,N_5189,N_7327);
nor U14609 (N_14609,N_8210,N_7188);
nand U14610 (N_14610,N_8265,N_8303);
nand U14611 (N_14611,N_6745,N_9905);
nor U14612 (N_14612,N_7650,N_5143);
or U14613 (N_14613,N_7317,N_9602);
or U14614 (N_14614,N_5805,N_9454);
nor U14615 (N_14615,N_7804,N_9462);
or U14616 (N_14616,N_9380,N_8021);
and U14617 (N_14617,N_6464,N_5197);
xnor U14618 (N_14618,N_9444,N_7163);
xor U14619 (N_14619,N_5951,N_9264);
or U14620 (N_14620,N_5956,N_6659);
xor U14621 (N_14621,N_6362,N_7352);
xnor U14622 (N_14622,N_9952,N_5231);
nand U14623 (N_14623,N_8591,N_8309);
nand U14624 (N_14624,N_9593,N_7872);
nand U14625 (N_14625,N_6502,N_9307);
nor U14626 (N_14626,N_9838,N_8664);
nand U14627 (N_14627,N_5660,N_7443);
nor U14628 (N_14628,N_5392,N_7874);
nor U14629 (N_14629,N_6976,N_9518);
and U14630 (N_14630,N_6580,N_6000);
xnor U14631 (N_14631,N_6526,N_7307);
nand U14632 (N_14632,N_7867,N_6128);
or U14633 (N_14633,N_6196,N_7245);
xnor U14634 (N_14634,N_7844,N_6566);
xnor U14635 (N_14635,N_5224,N_6527);
xnor U14636 (N_14636,N_8361,N_6704);
nor U14637 (N_14637,N_9291,N_6052);
nand U14638 (N_14638,N_9174,N_6595);
nor U14639 (N_14639,N_9674,N_7326);
nor U14640 (N_14640,N_6648,N_6652);
and U14641 (N_14641,N_8585,N_5364);
nor U14642 (N_14642,N_6769,N_6295);
or U14643 (N_14643,N_8569,N_7855);
nor U14644 (N_14644,N_6525,N_9509);
nor U14645 (N_14645,N_9357,N_8002);
and U14646 (N_14646,N_5839,N_7266);
or U14647 (N_14647,N_8579,N_5725);
nand U14648 (N_14648,N_9846,N_8332);
and U14649 (N_14649,N_8189,N_9732);
xor U14650 (N_14650,N_5424,N_7153);
nand U14651 (N_14651,N_7622,N_7352);
nand U14652 (N_14652,N_7307,N_7368);
and U14653 (N_14653,N_7784,N_9233);
xnor U14654 (N_14654,N_9486,N_5236);
or U14655 (N_14655,N_6169,N_8968);
nor U14656 (N_14656,N_7657,N_7029);
or U14657 (N_14657,N_7125,N_8288);
or U14658 (N_14658,N_6318,N_5796);
nor U14659 (N_14659,N_8753,N_5911);
or U14660 (N_14660,N_6197,N_8628);
nand U14661 (N_14661,N_5455,N_6971);
and U14662 (N_14662,N_8688,N_6760);
xnor U14663 (N_14663,N_9879,N_8451);
and U14664 (N_14664,N_6583,N_7333);
or U14665 (N_14665,N_7886,N_7170);
nor U14666 (N_14666,N_9942,N_7234);
nand U14667 (N_14667,N_6238,N_8746);
or U14668 (N_14668,N_9585,N_5345);
nand U14669 (N_14669,N_8441,N_5810);
and U14670 (N_14670,N_7259,N_9247);
nand U14671 (N_14671,N_9430,N_6613);
or U14672 (N_14672,N_6221,N_6130);
or U14673 (N_14673,N_9221,N_8185);
or U14674 (N_14674,N_9445,N_6994);
nor U14675 (N_14675,N_5337,N_5499);
nor U14676 (N_14676,N_5812,N_7610);
nor U14677 (N_14677,N_5234,N_5654);
xnor U14678 (N_14678,N_5775,N_9586);
xor U14679 (N_14679,N_7547,N_5041);
or U14680 (N_14680,N_8230,N_6270);
nor U14681 (N_14681,N_8499,N_5889);
nor U14682 (N_14682,N_8171,N_6926);
nor U14683 (N_14683,N_9608,N_5501);
nand U14684 (N_14684,N_5555,N_5263);
nand U14685 (N_14685,N_8803,N_5414);
xor U14686 (N_14686,N_5554,N_7921);
and U14687 (N_14687,N_9032,N_9465);
nand U14688 (N_14688,N_6049,N_9705);
and U14689 (N_14689,N_6183,N_6774);
xor U14690 (N_14690,N_6830,N_9524);
and U14691 (N_14691,N_7661,N_7354);
and U14692 (N_14692,N_9865,N_6754);
and U14693 (N_14693,N_9764,N_5567);
xor U14694 (N_14694,N_6332,N_7094);
or U14695 (N_14695,N_5479,N_9073);
or U14696 (N_14696,N_7519,N_7670);
nand U14697 (N_14697,N_8107,N_7654);
or U14698 (N_14698,N_5888,N_7488);
nor U14699 (N_14699,N_8781,N_5949);
xor U14700 (N_14700,N_8342,N_5114);
and U14701 (N_14701,N_6707,N_9500);
and U14702 (N_14702,N_5283,N_5421);
or U14703 (N_14703,N_7484,N_9674);
nor U14704 (N_14704,N_6427,N_8187);
nor U14705 (N_14705,N_5250,N_9526);
and U14706 (N_14706,N_8764,N_7504);
nor U14707 (N_14707,N_7616,N_9970);
xnor U14708 (N_14708,N_7806,N_5095);
xnor U14709 (N_14709,N_8716,N_7787);
or U14710 (N_14710,N_6103,N_8234);
or U14711 (N_14711,N_6665,N_8914);
nand U14712 (N_14712,N_6053,N_7978);
nand U14713 (N_14713,N_9210,N_9344);
or U14714 (N_14714,N_5545,N_7562);
nor U14715 (N_14715,N_5083,N_5246);
or U14716 (N_14716,N_5970,N_8354);
nand U14717 (N_14717,N_5422,N_9638);
or U14718 (N_14718,N_8577,N_5035);
xnor U14719 (N_14719,N_7372,N_9871);
and U14720 (N_14720,N_8405,N_7918);
xor U14721 (N_14721,N_5741,N_8840);
nor U14722 (N_14722,N_7868,N_9468);
or U14723 (N_14723,N_8535,N_8465);
xor U14724 (N_14724,N_9908,N_5750);
xnor U14725 (N_14725,N_8216,N_9384);
xor U14726 (N_14726,N_8962,N_9371);
nand U14727 (N_14727,N_6801,N_9279);
xor U14728 (N_14728,N_5402,N_9785);
nand U14729 (N_14729,N_9223,N_9807);
or U14730 (N_14730,N_9517,N_7977);
xnor U14731 (N_14731,N_9991,N_5383);
nor U14732 (N_14732,N_6894,N_9586);
and U14733 (N_14733,N_8008,N_8631);
or U14734 (N_14734,N_8898,N_5610);
nand U14735 (N_14735,N_6446,N_9881);
and U14736 (N_14736,N_5247,N_7921);
nand U14737 (N_14737,N_8158,N_6737);
nor U14738 (N_14738,N_8690,N_5739);
or U14739 (N_14739,N_5701,N_6485);
nor U14740 (N_14740,N_6592,N_9393);
nor U14741 (N_14741,N_8621,N_5864);
and U14742 (N_14742,N_7751,N_5154);
nand U14743 (N_14743,N_5958,N_5586);
nor U14744 (N_14744,N_6592,N_7948);
or U14745 (N_14745,N_7120,N_7002);
xor U14746 (N_14746,N_8538,N_7484);
nor U14747 (N_14747,N_8583,N_9713);
nand U14748 (N_14748,N_9988,N_9551);
xnor U14749 (N_14749,N_7793,N_7145);
nand U14750 (N_14750,N_6384,N_8556);
nor U14751 (N_14751,N_5413,N_8376);
and U14752 (N_14752,N_9724,N_9005);
xor U14753 (N_14753,N_8618,N_9816);
or U14754 (N_14754,N_8328,N_8762);
nor U14755 (N_14755,N_7762,N_5187);
nor U14756 (N_14756,N_5591,N_6686);
nand U14757 (N_14757,N_7095,N_8801);
or U14758 (N_14758,N_5912,N_5248);
nor U14759 (N_14759,N_5838,N_6673);
nand U14760 (N_14760,N_7729,N_6030);
and U14761 (N_14761,N_7907,N_6847);
and U14762 (N_14762,N_5690,N_9028);
xnor U14763 (N_14763,N_9962,N_9648);
or U14764 (N_14764,N_7813,N_8540);
nor U14765 (N_14765,N_6114,N_9616);
xnor U14766 (N_14766,N_5728,N_7777);
nand U14767 (N_14767,N_7990,N_9415);
and U14768 (N_14768,N_5742,N_6501);
or U14769 (N_14769,N_5768,N_5879);
or U14770 (N_14770,N_8536,N_7761);
xnor U14771 (N_14771,N_9190,N_7839);
nand U14772 (N_14772,N_8632,N_8104);
and U14773 (N_14773,N_6151,N_7580);
nor U14774 (N_14774,N_7701,N_6332);
nand U14775 (N_14775,N_7989,N_9035);
nand U14776 (N_14776,N_6471,N_9068);
nand U14777 (N_14777,N_6774,N_7849);
nand U14778 (N_14778,N_6872,N_8121);
nor U14779 (N_14779,N_9411,N_6315);
nor U14780 (N_14780,N_7105,N_5213);
xnor U14781 (N_14781,N_5397,N_5746);
or U14782 (N_14782,N_6163,N_9425);
nor U14783 (N_14783,N_9555,N_6151);
nand U14784 (N_14784,N_8810,N_9755);
nand U14785 (N_14785,N_7615,N_9321);
or U14786 (N_14786,N_9066,N_7498);
nand U14787 (N_14787,N_5210,N_7410);
nor U14788 (N_14788,N_6504,N_9612);
and U14789 (N_14789,N_6396,N_8693);
or U14790 (N_14790,N_8596,N_8771);
nand U14791 (N_14791,N_6403,N_7581);
and U14792 (N_14792,N_8672,N_5839);
nor U14793 (N_14793,N_5261,N_9934);
nand U14794 (N_14794,N_5813,N_8746);
nand U14795 (N_14795,N_5446,N_6003);
and U14796 (N_14796,N_7123,N_7496);
nand U14797 (N_14797,N_6917,N_7182);
nor U14798 (N_14798,N_7166,N_7877);
nor U14799 (N_14799,N_5240,N_9716);
or U14800 (N_14800,N_8175,N_8092);
or U14801 (N_14801,N_8860,N_6345);
nand U14802 (N_14802,N_7929,N_7818);
xnor U14803 (N_14803,N_8519,N_7781);
nor U14804 (N_14804,N_5477,N_9441);
xor U14805 (N_14805,N_7618,N_5823);
nor U14806 (N_14806,N_5185,N_8221);
xor U14807 (N_14807,N_5033,N_8747);
nand U14808 (N_14808,N_9870,N_5516);
xnor U14809 (N_14809,N_6251,N_9999);
or U14810 (N_14810,N_9947,N_7084);
and U14811 (N_14811,N_8252,N_5145);
nand U14812 (N_14812,N_5952,N_7623);
nand U14813 (N_14813,N_8771,N_7780);
xor U14814 (N_14814,N_6961,N_9451);
xor U14815 (N_14815,N_7550,N_7976);
nor U14816 (N_14816,N_5758,N_8010);
xor U14817 (N_14817,N_5311,N_7217);
xnor U14818 (N_14818,N_6597,N_6362);
nand U14819 (N_14819,N_9740,N_7056);
nand U14820 (N_14820,N_6109,N_8064);
and U14821 (N_14821,N_7992,N_7354);
nand U14822 (N_14822,N_7810,N_7840);
and U14823 (N_14823,N_8054,N_5786);
xor U14824 (N_14824,N_7229,N_6684);
or U14825 (N_14825,N_9241,N_9104);
nor U14826 (N_14826,N_9594,N_9783);
and U14827 (N_14827,N_9873,N_9034);
nor U14828 (N_14828,N_6141,N_5501);
and U14829 (N_14829,N_5559,N_5364);
nand U14830 (N_14830,N_9067,N_7369);
xnor U14831 (N_14831,N_7955,N_5315);
and U14832 (N_14832,N_8956,N_9506);
and U14833 (N_14833,N_7648,N_7470);
nor U14834 (N_14834,N_5447,N_8996);
nor U14835 (N_14835,N_6578,N_9460);
xnor U14836 (N_14836,N_6344,N_6949);
nor U14837 (N_14837,N_8778,N_7258);
or U14838 (N_14838,N_8807,N_6543);
nor U14839 (N_14839,N_8308,N_7937);
xor U14840 (N_14840,N_6216,N_6939);
and U14841 (N_14841,N_6751,N_8060);
and U14842 (N_14842,N_6494,N_5896);
or U14843 (N_14843,N_6372,N_6203);
and U14844 (N_14844,N_7983,N_7711);
or U14845 (N_14845,N_7297,N_5289);
nand U14846 (N_14846,N_7209,N_7330);
or U14847 (N_14847,N_8559,N_9226);
nor U14848 (N_14848,N_6405,N_9069);
nor U14849 (N_14849,N_5999,N_9291);
and U14850 (N_14850,N_9153,N_8742);
and U14851 (N_14851,N_7606,N_6830);
and U14852 (N_14852,N_5335,N_9354);
or U14853 (N_14853,N_5749,N_8316);
and U14854 (N_14854,N_5569,N_8813);
nand U14855 (N_14855,N_8842,N_6586);
xor U14856 (N_14856,N_7534,N_5991);
nand U14857 (N_14857,N_6412,N_5682);
xnor U14858 (N_14858,N_9775,N_5377);
nor U14859 (N_14859,N_9767,N_6869);
nand U14860 (N_14860,N_6596,N_9289);
or U14861 (N_14861,N_5939,N_9927);
and U14862 (N_14862,N_6334,N_8151);
or U14863 (N_14863,N_5592,N_9290);
or U14864 (N_14864,N_5942,N_8990);
and U14865 (N_14865,N_8206,N_9997);
nor U14866 (N_14866,N_9389,N_5075);
nand U14867 (N_14867,N_9592,N_9686);
nor U14868 (N_14868,N_6312,N_6945);
and U14869 (N_14869,N_9939,N_9132);
nand U14870 (N_14870,N_7548,N_8352);
and U14871 (N_14871,N_6339,N_9049);
xnor U14872 (N_14872,N_8627,N_9674);
or U14873 (N_14873,N_9407,N_8012);
or U14874 (N_14874,N_6418,N_7806);
nand U14875 (N_14875,N_5912,N_5688);
nand U14876 (N_14876,N_7000,N_7237);
xnor U14877 (N_14877,N_9461,N_6773);
or U14878 (N_14878,N_5949,N_7980);
xnor U14879 (N_14879,N_6874,N_9951);
nor U14880 (N_14880,N_5572,N_5709);
xor U14881 (N_14881,N_6863,N_7609);
xor U14882 (N_14882,N_9319,N_7762);
nor U14883 (N_14883,N_8451,N_8211);
and U14884 (N_14884,N_5745,N_6306);
and U14885 (N_14885,N_5587,N_7374);
xor U14886 (N_14886,N_5321,N_9155);
nand U14887 (N_14887,N_6458,N_9425);
and U14888 (N_14888,N_6784,N_7434);
xor U14889 (N_14889,N_8999,N_9204);
and U14890 (N_14890,N_6166,N_6667);
nor U14891 (N_14891,N_5318,N_6303);
and U14892 (N_14892,N_5521,N_9053);
nand U14893 (N_14893,N_9185,N_6814);
xor U14894 (N_14894,N_5511,N_5990);
nand U14895 (N_14895,N_8538,N_8994);
or U14896 (N_14896,N_8458,N_7847);
nand U14897 (N_14897,N_5604,N_8935);
nor U14898 (N_14898,N_5610,N_7182);
nand U14899 (N_14899,N_8483,N_6306);
nor U14900 (N_14900,N_6081,N_8089);
xor U14901 (N_14901,N_9816,N_9114);
nand U14902 (N_14902,N_8831,N_7566);
and U14903 (N_14903,N_7376,N_6365);
nor U14904 (N_14904,N_7800,N_5598);
xnor U14905 (N_14905,N_8131,N_6546);
xnor U14906 (N_14906,N_7563,N_7338);
nand U14907 (N_14907,N_6651,N_7489);
nand U14908 (N_14908,N_6806,N_6153);
nor U14909 (N_14909,N_6546,N_8051);
and U14910 (N_14910,N_6467,N_7700);
nand U14911 (N_14911,N_8283,N_7690);
nor U14912 (N_14912,N_5898,N_7999);
nand U14913 (N_14913,N_8887,N_5784);
nor U14914 (N_14914,N_5913,N_6791);
nand U14915 (N_14915,N_9263,N_9109);
xnor U14916 (N_14916,N_5682,N_7362);
xnor U14917 (N_14917,N_6172,N_9850);
nor U14918 (N_14918,N_8494,N_6389);
nor U14919 (N_14919,N_5029,N_8940);
or U14920 (N_14920,N_7098,N_5805);
or U14921 (N_14921,N_7874,N_7055);
and U14922 (N_14922,N_9188,N_7689);
xnor U14923 (N_14923,N_8165,N_9080);
and U14924 (N_14924,N_5282,N_7178);
nand U14925 (N_14925,N_8498,N_9368);
or U14926 (N_14926,N_5295,N_7397);
xnor U14927 (N_14927,N_5598,N_5233);
and U14928 (N_14928,N_7787,N_9624);
nor U14929 (N_14929,N_9887,N_6682);
xnor U14930 (N_14930,N_7661,N_9200);
and U14931 (N_14931,N_5742,N_7463);
or U14932 (N_14932,N_8075,N_9267);
nand U14933 (N_14933,N_7179,N_7035);
and U14934 (N_14934,N_8497,N_5114);
or U14935 (N_14935,N_5473,N_8453);
or U14936 (N_14936,N_5027,N_7504);
xnor U14937 (N_14937,N_8120,N_7376);
nor U14938 (N_14938,N_5334,N_5356);
nand U14939 (N_14939,N_6220,N_6729);
nand U14940 (N_14940,N_7523,N_6739);
nor U14941 (N_14941,N_8552,N_5639);
nand U14942 (N_14942,N_8804,N_8844);
nand U14943 (N_14943,N_6627,N_8902);
nand U14944 (N_14944,N_6102,N_7251);
and U14945 (N_14945,N_8456,N_6878);
nor U14946 (N_14946,N_9364,N_5889);
nand U14947 (N_14947,N_7225,N_5758);
and U14948 (N_14948,N_7944,N_7160);
or U14949 (N_14949,N_6315,N_7073);
nor U14950 (N_14950,N_6418,N_6032);
nor U14951 (N_14951,N_6531,N_9857);
and U14952 (N_14952,N_8418,N_9933);
nor U14953 (N_14953,N_7726,N_9577);
nor U14954 (N_14954,N_8044,N_6663);
nor U14955 (N_14955,N_7920,N_9222);
xor U14956 (N_14956,N_6629,N_7647);
nor U14957 (N_14957,N_9245,N_9178);
nand U14958 (N_14958,N_9036,N_6211);
or U14959 (N_14959,N_5413,N_9649);
nor U14960 (N_14960,N_8270,N_5373);
nor U14961 (N_14961,N_5068,N_7245);
nand U14962 (N_14962,N_7903,N_7938);
or U14963 (N_14963,N_7932,N_5813);
or U14964 (N_14964,N_9383,N_8526);
xor U14965 (N_14965,N_8850,N_9045);
xor U14966 (N_14966,N_6648,N_6456);
nand U14967 (N_14967,N_7994,N_7081);
nor U14968 (N_14968,N_5507,N_6356);
xor U14969 (N_14969,N_7449,N_7404);
nand U14970 (N_14970,N_6907,N_5989);
or U14971 (N_14971,N_8037,N_8042);
nor U14972 (N_14972,N_7128,N_8588);
nand U14973 (N_14973,N_7383,N_9613);
xnor U14974 (N_14974,N_9954,N_8949);
nand U14975 (N_14975,N_7929,N_8650);
or U14976 (N_14976,N_9974,N_8640);
or U14977 (N_14977,N_9765,N_7303);
nor U14978 (N_14978,N_6208,N_9218);
nand U14979 (N_14979,N_5870,N_5805);
xnor U14980 (N_14980,N_5956,N_8904);
or U14981 (N_14981,N_9063,N_5828);
or U14982 (N_14982,N_7219,N_6628);
xnor U14983 (N_14983,N_8361,N_9837);
and U14984 (N_14984,N_7320,N_8742);
and U14985 (N_14985,N_5864,N_9833);
nor U14986 (N_14986,N_9942,N_5754);
nor U14987 (N_14987,N_5473,N_5627);
or U14988 (N_14988,N_7420,N_6272);
nor U14989 (N_14989,N_8635,N_9006);
xor U14990 (N_14990,N_8389,N_7982);
and U14991 (N_14991,N_7688,N_8836);
and U14992 (N_14992,N_7606,N_7391);
and U14993 (N_14993,N_9477,N_5504);
nor U14994 (N_14994,N_7236,N_6221);
nand U14995 (N_14995,N_8038,N_8478);
and U14996 (N_14996,N_9377,N_8830);
nand U14997 (N_14997,N_6811,N_7256);
or U14998 (N_14998,N_9601,N_5125);
xor U14999 (N_14999,N_8793,N_5490);
nand U15000 (N_15000,N_10035,N_11910);
or U15001 (N_15001,N_14653,N_12899);
xnor U15002 (N_15002,N_10520,N_12012);
and U15003 (N_15003,N_11587,N_13469);
and U15004 (N_15004,N_10358,N_13029);
xor U15005 (N_15005,N_13838,N_14755);
nor U15006 (N_15006,N_11275,N_11245);
nor U15007 (N_15007,N_10327,N_12351);
xor U15008 (N_15008,N_11929,N_14379);
nor U15009 (N_15009,N_10749,N_13586);
nand U15010 (N_15010,N_11339,N_11725);
or U15011 (N_15011,N_12652,N_11482);
or U15012 (N_15012,N_14642,N_13863);
and U15013 (N_15013,N_13743,N_10343);
or U15014 (N_15014,N_11206,N_13898);
and U15015 (N_15015,N_10100,N_14896);
xor U15016 (N_15016,N_12013,N_13950);
or U15017 (N_15017,N_13584,N_12076);
xnor U15018 (N_15018,N_10257,N_11370);
nand U15019 (N_15019,N_11078,N_12122);
and U15020 (N_15020,N_12363,N_14699);
nand U15021 (N_15021,N_10978,N_14992);
and U15022 (N_15022,N_12781,N_14544);
xor U15023 (N_15023,N_10124,N_14621);
xor U15024 (N_15024,N_11267,N_11333);
xnor U15025 (N_15025,N_13250,N_11118);
xor U15026 (N_15026,N_12699,N_11302);
xnor U15027 (N_15027,N_12901,N_14469);
or U15028 (N_15028,N_14672,N_12043);
or U15029 (N_15029,N_11262,N_10466);
and U15030 (N_15030,N_11697,N_13120);
and U15031 (N_15031,N_10965,N_10345);
or U15032 (N_15032,N_13585,N_13240);
and U15033 (N_15033,N_10059,N_12026);
nor U15034 (N_15034,N_12609,N_10033);
nand U15035 (N_15035,N_13078,N_10092);
or U15036 (N_15036,N_12033,N_13079);
nand U15037 (N_15037,N_13775,N_13464);
xnor U15038 (N_15038,N_10564,N_14768);
nor U15039 (N_15039,N_14499,N_13038);
and U15040 (N_15040,N_12660,N_12923);
or U15041 (N_15041,N_11885,N_12961);
nor U15042 (N_15042,N_13714,N_11678);
nor U15043 (N_15043,N_11556,N_14888);
and U15044 (N_15044,N_13566,N_11427);
and U15045 (N_15045,N_11379,N_14721);
or U15046 (N_15046,N_13961,N_10933);
nand U15047 (N_15047,N_14317,N_13049);
nor U15048 (N_15048,N_12889,N_10648);
nand U15049 (N_15049,N_13657,N_13210);
xnor U15050 (N_15050,N_12665,N_13242);
xor U15051 (N_15051,N_11840,N_12563);
and U15052 (N_15052,N_10006,N_13612);
or U15053 (N_15053,N_10819,N_10783);
and U15054 (N_15054,N_14675,N_13902);
and U15055 (N_15055,N_10444,N_11684);
nand U15056 (N_15056,N_11581,N_14904);
nand U15057 (N_15057,N_13670,N_12502);
and U15058 (N_15058,N_12397,N_11366);
nand U15059 (N_15059,N_10793,N_13747);
xnor U15060 (N_15060,N_11374,N_12814);
or U15061 (N_15061,N_12433,N_11500);
and U15062 (N_15062,N_14879,N_14179);
nand U15063 (N_15063,N_14032,N_10646);
and U15064 (N_15064,N_11726,N_13324);
xnor U15065 (N_15065,N_11720,N_13036);
xnor U15066 (N_15066,N_12119,N_10116);
or U15067 (N_15067,N_12361,N_12559);
or U15068 (N_15068,N_14163,N_14223);
nor U15069 (N_15069,N_13191,N_10080);
or U15070 (N_15070,N_14853,N_13713);
nand U15071 (N_15071,N_10065,N_14463);
xnor U15072 (N_15072,N_11942,N_10890);
and U15073 (N_15073,N_13248,N_13587);
nor U15074 (N_15074,N_14685,N_11598);
or U15075 (N_15075,N_11316,N_12913);
xor U15076 (N_15076,N_11130,N_11026);
xor U15077 (N_15077,N_14292,N_11924);
nor U15078 (N_15078,N_11681,N_11735);
and U15079 (N_15079,N_14016,N_11306);
or U15080 (N_15080,N_10150,N_13255);
nand U15081 (N_15081,N_12545,N_12516);
nand U15082 (N_15082,N_12843,N_13589);
nor U15083 (N_15083,N_11852,N_13223);
nor U15084 (N_15084,N_13619,N_13938);
nand U15085 (N_15085,N_14967,N_11994);
xnor U15086 (N_15086,N_14489,N_14341);
and U15087 (N_15087,N_10631,N_12943);
xnor U15088 (N_15088,N_11979,N_14459);
or U15089 (N_15089,N_14765,N_11626);
nor U15090 (N_15090,N_12170,N_12975);
and U15091 (N_15091,N_10392,N_12746);
nand U15092 (N_15092,N_10692,N_10587);
xnor U15093 (N_15093,N_10740,N_10734);
nand U15094 (N_15094,N_14156,N_13075);
nor U15095 (N_15095,N_11619,N_10312);
or U15096 (N_15096,N_14322,N_12616);
nand U15097 (N_15097,N_14940,N_14411);
and U15098 (N_15098,N_12256,N_10229);
xor U15099 (N_15099,N_12275,N_13606);
nor U15100 (N_15100,N_13887,N_14662);
xnor U15101 (N_15101,N_10976,N_14885);
xor U15102 (N_15102,N_11935,N_10627);
xnor U15103 (N_15103,N_11080,N_14218);
or U15104 (N_15104,N_13245,N_13087);
and U15105 (N_15105,N_12242,N_13328);
or U15106 (N_15106,N_13807,N_14628);
nand U15107 (N_15107,N_14878,N_14908);
xor U15108 (N_15108,N_14789,N_10338);
nand U15109 (N_15109,N_14188,N_13795);
xor U15110 (N_15110,N_10313,N_10908);
nor U15111 (N_15111,N_13802,N_14894);
xnor U15112 (N_15112,N_14217,N_11066);
and U15113 (N_15113,N_14356,N_11165);
or U15114 (N_15114,N_11522,N_10613);
xnor U15115 (N_15115,N_11722,N_11595);
nand U15116 (N_15116,N_10935,N_10544);
nor U15117 (N_15117,N_14187,N_13820);
nor U15118 (N_15118,N_12022,N_12530);
or U15119 (N_15119,N_13572,N_13972);
or U15120 (N_15120,N_12954,N_13192);
and U15121 (N_15121,N_13900,N_13234);
nor U15122 (N_15122,N_11006,N_11955);
nand U15123 (N_15123,N_11831,N_14503);
nand U15124 (N_15124,N_14998,N_14727);
and U15125 (N_15125,N_14668,N_11624);
or U15126 (N_15126,N_13721,N_11393);
nor U15127 (N_15127,N_10770,N_10836);
and U15128 (N_15128,N_12542,N_10738);
and U15129 (N_15129,N_14603,N_14763);
and U15130 (N_15130,N_10282,N_10295);
and U15131 (N_15131,N_13065,N_14947);
nand U15132 (N_15132,N_11644,N_11279);
and U15133 (N_15133,N_12598,N_12115);
xor U15134 (N_15134,N_10974,N_13487);
and U15135 (N_15135,N_14679,N_12876);
xnor U15136 (N_15136,N_11934,N_13733);
xnor U15137 (N_15137,N_10478,N_11304);
nor U15138 (N_15138,N_11421,N_14135);
nand U15139 (N_15139,N_11780,N_12558);
nor U15140 (N_15140,N_10326,N_11752);
xnor U15141 (N_15141,N_12164,N_11639);
xor U15142 (N_15142,N_12072,N_11822);
nor U15143 (N_15143,N_12168,N_11751);
xor U15144 (N_15144,N_10781,N_13856);
nor U15145 (N_15145,N_10460,N_13549);
xnor U15146 (N_15146,N_14029,N_12509);
or U15147 (N_15147,N_13564,N_11582);
xnor U15148 (N_15148,N_12780,N_10996);
nor U15149 (N_15149,N_14663,N_12527);
nand U15150 (N_15150,N_11982,N_10024);
nand U15151 (N_15151,N_12725,N_14019);
xnor U15152 (N_15152,N_10171,N_11219);
and U15153 (N_15153,N_12903,N_13405);
nand U15154 (N_15154,N_12310,N_11159);
xor U15155 (N_15155,N_14722,N_13921);
nor U15156 (N_15156,N_11826,N_10046);
xor U15157 (N_15157,N_12649,N_14664);
nor U15158 (N_15158,N_14932,N_12970);
xnor U15159 (N_15159,N_10379,N_11378);
nor U15160 (N_15160,N_10652,N_10166);
or U15161 (N_15161,N_13720,N_11569);
nor U15162 (N_15162,N_14866,N_13004);
nand U15163 (N_15163,N_11693,N_12192);
and U15164 (N_15164,N_13243,N_12474);
nor U15165 (N_15165,N_14512,N_14733);
xnor U15166 (N_15166,N_10412,N_11170);
or U15167 (N_15167,N_12133,N_13423);
xnor U15168 (N_15168,N_11001,N_11322);
nand U15169 (N_15169,N_12618,N_10626);
or U15170 (N_15170,N_13574,N_14625);
nor U15171 (N_15171,N_13647,N_13035);
nor U15172 (N_15172,N_11814,N_10195);
xnor U15173 (N_15173,N_13579,N_12511);
or U15174 (N_15174,N_10797,N_12146);
and U15175 (N_15175,N_12657,N_10363);
and U15176 (N_15176,N_13292,N_13077);
nor U15177 (N_15177,N_13497,N_10403);
or U15178 (N_15178,N_10804,N_13744);
or U15179 (N_15179,N_10001,N_14980);
nand U15180 (N_15180,N_11583,N_14263);
nor U15181 (N_15181,N_11612,N_11793);
nand U15182 (N_15182,N_13148,N_10243);
or U15183 (N_15183,N_12944,N_13851);
nand U15184 (N_15184,N_10141,N_11059);
and U15185 (N_15185,N_13433,N_12856);
and U15186 (N_15186,N_13417,N_10639);
xor U15187 (N_15187,N_13013,N_10490);
and U15188 (N_15188,N_13793,N_10433);
nor U15189 (N_15189,N_14073,N_14922);
or U15190 (N_15190,N_11796,N_14192);
and U15191 (N_15191,N_13053,N_13341);
nor U15192 (N_15192,N_12764,N_10228);
xor U15193 (N_15193,N_13421,N_11155);
nor U15194 (N_15194,N_10027,N_10757);
xnor U15195 (N_15195,N_11860,N_12708);
and U15196 (N_15196,N_13395,N_13490);
nand U15197 (N_15197,N_12960,N_14429);
xor U15198 (N_15198,N_13129,N_13225);
nor U15199 (N_15199,N_11889,N_10203);
xor U15200 (N_15200,N_11097,N_12514);
nand U15201 (N_15201,N_14375,N_11489);
nor U15202 (N_15202,N_10108,N_14149);
and U15203 (N_15203,N_11090,N_12243);
or U15204 (N_15204,N_13704,N_14775);
and U15205 (N_15205,N_11638,N_10842);
nor U15206 (N_15206,N_10088,N_14288);
nor U15207 (N_15207,N_13609,N_12315);
xnor U15208 (N_15208,N_11975,N_11252);
and U15209 (N_15209,N_14123,N_11133);
and U15210 (N_15210,N_10484,N_14307);
xnor U15211 (N_15211,N_14510,N_13684);
nand U15212 (N_15212,N_12297,N_10849);
nand U15213 (N_15213,N_14027,N_12157);
nand U15214 (N_15214,N_12495,N_10920);
xor U15215 (N_15215,N_13529,N_12633);
or U15216 (N_15216,N_11347,N_12829);
and U15217 (N_15217,N_12393,N_10630);
or U15218 (N_15218,N_12600,N_10402);
nand U15219 (N_15219,N_11677,N_11178);
nor U15220 (N_15220,N_14600,N_13452);
nor U15221 (N_15221,N_10875,N_13352);
nor U15222 (N_15222,N_13147,N_13880);
xnor U15223 (N_15223,N_14801,N_10720);
xnor U15224 (N_15224,N_14630,N_10763);
and U15225 (N_15225,N_10794,N_12679);
or U15226 (N_15226,N_14207,N_14482);
and U15227 (N_15227,N_12670,N_13888);
nor U15228 (N_15228,N_14654,N_14020);
xor U15229 (N_15229,N_10410,N_13396);
nand U15230 (N_15230,N_12084,N_10064);
and U15231 (N_15231,N_12064,N_10208);
xnor U15232 (N_15232,N_13336,N_10120);
nand U15233 (N_15233,N_14779,N_13629);
nand U15234 (N_15234,N_14046,N_14959);
nor U15235 (N_15235,N_11862,N_12668);
or U15236 (N_15236,N_10084,N_11151);
nor U15237 (N_15237,N_11498,N_14846);
xnor U15238 (N_15238,N_13310,N_14077);
or U15239 (N_15239,N_11691,N_14747);
and U15240 (N_15240,N_11487,N_14911);
xor U15241 (N_15241,N_10661,N_14443);
or U15242 (N_15242,N_12544,N_10917);
or U15243 (N_15243,N_12127,N_12196);
or U15244 (N_15244,N_11832,N_14355);
xor U15245 (N_15245,N_14816,N_12244);
nand U15246 (N_15246,N_13694,N_14232);
xor U15247 (N_15247,N_13555,N_12367);
xor U15248 (N_15248,N_10384,N_10651);
nand U15249 (N_15249,N_13932,N_14152);
nor U15250 (N_15250,N_13548,N_12571);
xor U15251 (N_15251,N_11880,N_14487);
and U15252 (N_15252,N_14971,N_11939);
nor U15253 (N_15253,N_13127,N_13788);
and U15254 (N_15254,N_11108,N_10562);
xor U15255 (N_15255,N_13528,N_13655);
nor U15256 (N_15256,N_11235,N_11485);
nand U15257 (N_15257,N_11396,N_10638);
xor U15258 (N_15258,N_13088,N_12295);
nor U15259 (N_15259,N_14395,N_10514);
nor U15260 (N_15260,N_10971,N_11398);
or U15261 (N_15261,N_14277,N_10669);
nor U15262 (N_15262,N_10168,N_10553);
xor U15263 (N_15263,N_12352,N_10095);
or U15264 (N_15264,N_11403,N_11968);
nand U15265 (N_15265,N_11911,N_12933);
nand U15266 (N_15266,N_12240,N_14891);
nand U15267 (N_15267,N_10915,N_12160);
nand U15268 (N_15268,N_14072,N_13832);
and U15269 (N_15269,N_11286,N_12309);
xor U15270 (N_15270,N_14478,N_12650);
nand U15271 (N_15271,N_14890,N_13617);
nand U15272 (N_15272,N_14227,N_11740);
xor U15273 (N_15273,N_12925,N_11315);
xnor U15274 (N_15274,N_12967,N_11011);
nand U15275 (N_15275,N_14514,N_11341);
nand U15276 (N_15276,N_10710,N_10011);
nor U15277 (N_15277,N_10409,N_14414);
nor U15278 (N_15278,N_13169,N_12015);
nor U15279 (N_15279,N_13446,N_11513);
nor U15280 (N_15280,N_12184,N_11652);
nor U15281 (N_15281,N_10887,N_11297);
and U15282 (N_15282,N_13136,N_10582);
nand U15283 (N_15283,N_11953,N_10950);
nand U15284 (N_15284,N_11258,N_13749);
and U15285 (N_15285,N_12258,N_14354);
nor U15286 (N_15286,N_10707,N_12999);
or U15287 (N_15287,N_14731,N_13676);
or U15288 (N_15288,N_11292,N_12890);
nor U15289 (N_15289,N_13030,N_12178);
and U15290 (N_15290,N_12197,N_13910);
xnor U15291 (N_15291,N_11041,N_12448);
and U15292 (N_15292,N_13906,N_14391);
and U15293 (N_15293,N_14465,N_12507);
xnor U15294 (N_15294,N_11147,N_10489);
xnor U15295 (N_15295,N_13484,N_10016);
nand U15296 (N_15296,N_11864,N_12892);
nand U15297 (N_15297,N_10142,N_14559);
or U15298 (N_15298,N_12117,N_12150);
or U15299 (N_15299,N_14047,N_14678);
xnor U15300 (N_15300,N_10317,N_11457);
or U15301 (N_15301,N_11153,N_12199);
or U15302 (N_15302,N_14126,N_13442);
xor U15303 (N_15303,N_14538,N_12344);
nor U15304 (N_15304,N_12910,N_11137);
and U15305 (N_15305,N_13154,N_10350);
and U15306 (N_15306,N_10383,N_12902);
xnor U15307 (N_15307,N_12019,N_13343);
nor U15308 (N_15308,N_12938,N_11891);
or U15309 (N_15309,N_11372,N_10139);
and U15310 (N_15310,N_12947,N_11318);
nand U15311 (N_15311,N_10276,N_14105);
or U15312 (N_15312,N_10333,N_12748);
nor U15313 (N_15313,N_14726,N_13739);
nand U15314 (N_15314,N_12800,N_11463);
xnor U15315 (N_15315,N_13847,N_13259);
nand U15316 (N_15316,N_14370,N_14208);
nor U15317 (N_15317,N_11280,N_12723);
nand U15318 (N_15318,N_14210,N_14169);
or U15319 (N_15319,N_10795,N_14404);
nand U15320 (N_15320,N_13841,N_11818);
nor U15321 (N_15321,N_12267,N_11761);
and U15322 (N_15322,N_12908,N_12341);
or U15323 (N_15323,N_11283,N_11524);
nand U15324 (N_15324,N_13717,N_10604);
nand U15325 (N_15325,N_11656,N_14068);
xnor U15326 (N_15326,N_11486,N_14457);
xnor U15327 (N_15327,N_13023,N_14636);
and U15328 (N_15328,N_13355,N_14461);
xor U15329 (N_15329,N_12586,N_12532);
nand U15330 (N_15330,N_14573,N_12758);
or U15331 (N_15331,N_10921,N_12928);
and U15332 (N_15332,N_14724,N_11892);
nor U15333 (N_15333,N_10833,N_11674);
nor U15334 (N_15334,N_13089,N_11266);
xor U15335 (N_15335,N_11932,N_12840);
nor U15336 (N_15336,N_11950,N_13440);
or U15337 (N_15337,N_11958,N_11127);
nor U15338 (N_15338,N_12667,N_11695);
nor U15339 (N_15339,N_10019,N_13545);
and U15340 (N_15340,N_11749,N_11085);
nor U15341 (N_15341,N_12365,N_13418);
or U15342 (N_15342,N_11949,N_13507);
nand U15343 (N_15343,N_11961,N_10411);
nor U15344 (N_15344,N_12986,N_11301);
nand U15345 (N_15345,N_13881,N_10187);
or U15346 (N_15346,N_10873,N_14641);
nand U15347 (N_15347,N_11107,N_14661);
nand U15348 (N_15348,N_12741,N_10464);
nand U15349 (N_15349,N_12317,N_11801);
or U15350 (N_15350,N_11661,N_12203);
xnor U15351 (N_15351,N_13295,N_11764);
or U15352 (N_15352,N_14591,N_11923);
nor U15353 (N_15353,N_12305,N_10518);
nor U15354 (N_15354,N_13687,N_10854);
and U15355 (N_15355,N_13400,N_14114);
nor U15356 (N_15356,N_14336,N_10815);
or U15357 (N_15357,N_11050,N_12038);
nand U15358 (N_15358,N_14083,N_14570);
or U15359 (N_15359,N_11918,N_13297);
or U15360 (N_15360,N_14780,N_11914);
and U15361 (N_15361,N_11597,N_13133);
or U15362 (N_15362,N_10808,N_10280);
nor U15363 (N_15363,N_10928,N_11040);
or U15364 (N_15364,N_14874,N_13215);
nor U15365 (N_15365,N_11857,N_11493);
nand U15366 (N_15366,N_11744,N_10633);
nand U15367 (N_15367,N_12370,N_13422);
nor U15368 (N_15368,N_10185,N_12381);
or U15369 (N_15369,N_10247,N_12328);
nand U15370 (N_15370,N_13812,N_10759);
nand U15371 (N_15371,N_13673,N_11909);
and U15372 (N_15372,N_10913,N_10113);
nor U15373 (N_15373,N_12624,N_10086);
nand U15374 (N_15374,N_12035,N_11998);
xnor U15375 (N_15375,N_10264,N_14914);
nor U15376 (N_15376,N_14310,N_13196);
and U15377 (N_15377,N_11613,N_14583);
or U15378 (N_15378,N_11590,N_12217);
and U15379 (N_15379,N_11988,N_13517);
xor U15380 (N_15380,N_11441,N_14753);
or U15381 (N_15381,N_10292,N_11972);
nand U15382 (N_15382,N_13068,N_10048);
nor U15383 (N_15383,N_13115,N_12483);
and U15384 (N_15384,N_14593,N_13000);
or U15385 (N_15385,N_14071,N_11380);
nand U15386 (N_15386,N_11736,N_13045);
xor U15387 (N_15387,N_14001,N_13185);
nor U15388 (N_15388,N_12603,N_14587);
and U15389 (N_15389,N_11284,N_13176);
nand U15390 (N_15390,N_13924,N_13311);
xnor U15391 (N_15391,N_14554,N_13244);
or U15392 (N_15392,N_11896,N_11064);
or U15393 (N_15393,N_14855,N_10746);
or U15394 (N_15394,N_14546,N_10625);
and U15395 (N_15395,N_10956,N_13506);
and U15396 (N_15396,N_10285,N_10737);
or U15397 (N_15397,N_12612,N_11999);
nor U15398 (N_15398,N_11675,N_11476);
or U15399 (N_15399,N_10507,N_13450);
nor U15400 (N_15400,N_13971,N_10936);
xor U15401 (N_15401,N_13489,N_13104);
or U15402 (N_15402,N_13016,N_12429);
nor U15403 (N_15403,N_10161,N_14342);
or U15404 (N_15404,N_12587,N_14939);
nand U15405 (N_15405,N_11765,N_12059);
xor U15406 (N_15406,N_12697,N_10910);
and U15407 (N_15407,N_12086,N_10330);
nand U15408 (N_15408,N_13407,N_10752);
xor U15409 (N_15409,N_14245,N_11629);
nand U15410 (N_15410,N_10762,N_11508);
or U15411 (N_15411,N_12354,N_14820);
nor U15412 (N_15412,N_11960,N_10445);
nand U15413 (N_15413,N_12732,N_13680);
or U15414 (N_15414,N_14669,N_14455);
and U15415 (N_15415,N_10602,N_10703);
and U15416 (N_15416,N_11802,N_12226);
nor U15417 (N_15417,N_12120,N_10642);
xor U15418 (N_15418,N_10101,N_14657);
and U15419 (N_15419,N_10422,N_10127);
xor U15420 (N_15420,N_14344,N_10975);
nor U15421 (N_15421,N_11854,N_14225);
xor U15422 (N_15422,N_12109,N_10533);
nand U15423 (N_15423,N_13685,N_12394);
nor U15424 (N_15424,N_13597,N_14204);
nor U15425 (N_15425,N_12093,N_11231);
nor U15426 (N_15426,N_11803,N_10431);
or U15427 (N_15427,N_11188,N_10586);
xor U15428 (N_15428,N_10784,N_10199);
nor U15429 (N_15429,N_10463,N_14873);
or U15430 (N_15430,N_12081,N_10342);
xnor U15431 (N_15431,N_13897,N_11732);
xnor U15432 (N_15432,N_11196,N_12137);
or U15433 (N_15433,N_13062,N_14979);
and U15434 (N_15434,N_14623,N_11076);
and U15435 (N_15435,N_13019,N_13956);
or U15436 (N_15436,N_13552,N_10684);
or U15437 (N_15437,N_12687,N_12833);
nor U15438 (N_15438,N_11827,N_13042);
or U15439 (N_15439,N_10066,N_14451);
and U15440 (N_15440,N_12460,N_10365);
xor U15441 (N_15441,N_11992,N_11230);
xnor U15442 (N_15442,N_14248,N_12294);
xor U15443 (N_15443,N_11824,N_11883);
xor U15444 (N_15444,N_11409,N_13153);
or U15445 (N_15445,N_10308,N_10140);
or U15446 (N_15446,N_13630,N_13535);
nand U15447 (N_15447,N_13372,N_14427);
xnor U15448 (N_15448,N_13190,N_14962);
nand U15449 (N_15449,N_14371,N_14303);
nor U15450 (N_15450,N_14045,N_10013);
or U15451 (N_15451,N_10690,N_13928);
or U15452 (N_15452,N_12490,N_14024);
nand U15453 (N_15453,N_14334,N_14863);
xnor U15454 (N_15454,N_12391,N_14677);
and U15455 (N_15455,N_14405,N_13622);
xor U15456 (N_15456,N_11669,N_13702);
nor U15457 (N_15457,N_12279,N_13282);
nor U15458 (N_15458,N_10114,N_14576);
xor U15459 (N_15459,N_14580,N_10443);
or U15460 (N_15460,N_14422,N_11468);
nor U15461 (N_15461,N_11634,N_11614);
or U15462 (N_15462,N_11637,N_12060);
or U15463 (N_15463,N_12976,N_14617);
nand U15464 (N_15464,N_12054,N_11326);
xnor U15465 (N_15465,N_12034,N_11220);
nand U15466 (N_15466,N_14644,N_12782);
or U15467 (N_15467,N_14133,N_11828);
and U15468 (N_15468,N_12247,N_13025);
nand U15469 (N_15469,N_12557,N_10827);
nand U15470 (N_15470,N_11298,N_14445);
nand U15471 (N_15471,N_13010,N_11753);
or U15472 (N_15472,N_13594,N_12037);
nand U15473 (N_15473,N_11271,N_10503);
nand U15474 (N_15474,N_11375,N_14782);
xnor U15475 (N_15475,N_10271,N_10611);
or U15476 (N_15476,N_11841,N_12783);
or U15477 (N_15477,N_13868,N_10432);
nor U15478 (N_15478,N_10045,N_11213);
and U15479 (N_15479,N_13050,N_12734);
and U15480 (N_15480,N_10126,N_12271);
nand U15481 (N_15481,N_14869,N_12148);
and U15482 (N_15482,N_13985,N_13844);
nand U15483 (N_15483,N_10964,N_11715);
and U15484 (N_15484,N_11943,N_10122);
or U15485 (N_15485,N_13709,N_12266);
and U15486 (N_15486,N_13699,N_10820);
xnor U15487 (N_15487,N_13911,N_10717);
nand U15488 (N_15488,N_11983,N_12424);
or U15489 (N_15489,N_11743,N_12193);
xor U15490 (N_15490,N_10335,N_10942);
and U15491 (N_15491,N_13759,N_13893);
nor U15492 (N_15492,N_11676,N_12291);
xor U15493 (N_15493,N_12531,N_13117);
nor U15494 (N_15494,N_13438,N_10550);
nor U15495 (N_15495,N_10987,N_13351);
or U15496 (N_15496,N_12916,N_14881);
nand U15497 (N_15497,N_11173,N_10796);
nand U15498 (N_15498,N_14774,N_13536);
or U15499 (N_15499,N_10198,N_10089);
or U15500 (N_15500,N_12255,N_10014);
xnor U15501 (N_15501,N_11451,N_13247);
nor U15502 (N_15502,N_12039,N_14825);
xor U15503 (N_15503,N_13819,N_11115);
nand U15504 (N_15504,N_10773,N_14452);
or U15505 (N_15505,N_12503,N_11847);
nor U15506 (N_15506,N_10760,N_12103);
or U15507 (N_15507,N_13451,N_14471);
nand U15508 (N_15508,N_13278,N_14950);
or U15509 (N_15509,N_14448,N_10647);
xnor U15510 (N_15510,N_12324,N_10315);
and U15511 (N_15511,N_10961,N_13140);
nand U15512 (N_15512,N_12068,N_11881);
nand U15513 (N_15513,N_12658,N_10191);
nand U15514 (N_15514,N_14244,N_14498);
nand U15515 (N_15515,N_11989,N_11533);
xor U15516 (N_15516,N_11705,N_14707);
nor U15517 (N_15517,N_10217,N_12036);
nand U15518 (N_15518,N_10702,N_14148);
nand U15519 (N_15519,N_12191,N_12770);
xor U15520 (N_15520,N_14106,N_12823);
xnor U15521 (N_15521,N_10552,N_10778);
xnor U15522 (N_15522,N_12619,N_10307);
nand U15523 (N_15523,N_13272,N_14477);
nor U15524 (N_15524,N_11855,N_10202);
nor U15525 (N_15525,N_11816,N_10968);
or U15526 (N_15526,N_13514,N_13799);
xor U15527 (N_15527,N_14970,N_12853);
nor U15528 (N_15528,N_14807,N_12578);
xnor U15529 (N_15529,N_10509,N_11215);
xor U15530 (N_15530,N_13095,N_13951);
xnor U15531 (N_15531,N_14502,N_12525);
or U15532 (N_15532,N_14095,N_12614);
and U15533 (N_15533,N_11716,N_14285);
and U15534 (N_15534,N_10026,N_11861);
and U15535 (N_15535,N_10578,N_14257);
and U15536 (N_15536,N_11323,N_10709);
nand U15537 (N_15537,N_10272,N_10779);
or U15538 (N_15538,N_12232,N_12946);
nand U15539 (N_15539,N_12470,N_11324);
or U15540 (N_15540,N_13556,N_11194);
xnor U15541 (N_15541,N_10818,N_14655);
xor U15542 (N_15542,N_13992,N_11377);
nor U15543 (N_15543,N_13659,N_14075);
nor U15544 (N_15544,N_11022,N_11264);
nand U15545 (N_15545,N_11340,N_11986);
nand U15546 (N_15546,N_13842,N_11707);
nand U15547 (N_15547,N_11210,N_14633);
xor U15548 (N_15548,N_10325,N_12069);
nor U15549 (N_15549,N_13508,N_14042);
nor U15550 (N_15550,N_11865,N_10672);
nand U15551 (N_15551,N_11466,N_14886);
nor U15552 (N_15552,N_14629,N_12506);
nor U15553 (N_15553,N_10306,N_11241);
and U15554 (N_15554,N_13866,N_10377);
nor U15555 (N_15555,N_10385,N_10667);
or U15556 (N_15556,N_13108,N_14013);
and U15557 (N_15557,N_14826,N_14361);
xor U15558 (N_15558,N_11905,N_11680);
or U15559 (N_15559,N_10269,N_10851);
xnor U15560 (N_15560,N_12410,N_11850);
xnor U15561 (N_15561,N_12898,N_12759);
and U15562 (N_15562,N_11520,N_10858);
or U15563 (N_15563,N_11250,N_14534);
nand U15564 (N_15564,N_13503,N_13873);
nand U15565 (N_15565,N_13895,N_12994);
and U15566 (N_15566,N_14040,N_13430);
nand U15567 (N_15567,N_14719,N_11700);
nand U15568 (N_15568,N_11083,N_13063);
nand U15569 (N_15569,N_12216,N_12466);
xor U15570 (N_15570,N_14057,N_10025);
and U15571 (N_15571,N_10905,N_14390);
or U15572 (N_15572,N_12834,N_13304);
nand U15573 (N_15573,N_14279,N_13265);
or U15574 (N_15574,N_11048,N_13009);
or U15575 (N_15575,N_12597,N_13066);
xnor U15576 (N_15576,N_13679,N_10575);
xor U15577 (N_15577,N_11430,N_12447);
and U15578 (N_15578,N_10641,N_13738);
and U15579 (N_15579,N_10153,N_12893);
xor U15580 (N_15580,N_14986,N_10018);
nand U15581 (N_15581,N_13313,N_10215);
and U15582 (N_15582,N_11407,N_13661);
xnor U15583 (N_15583,N_11390,N_10303);
nand U15584 (N_15584,N_10294,N_14278);
and U15585 (N_15585,N_13220,N_13974);
or U15586 (N_15586,N_12175,N_11564);
and U15587 (N_15587,N_12135,N_10049);
nand U15588 (N_15588,N_13591,N_13779);
or U15589 (N_15589,N_14194,N_14144);
nand U15590 (N_15590,N_14735,N_12302);
nand U15591 (N_15591,N_14978,N_12980);
or U15592 (N_15592,N_12413,N_11207);
nand U15593 (N_15593,N_13157,N_11654);
and U15594 (N_15594,N_13273,N_14828);
xnor U15595 (N_15595,N_14612,N_12897);
nor U15596 (N_15596,N_14030,N_11906);
nor U15597 (N_15597,N_11072,N_11470);
or U15598 (N_15598,N_11104,N_11603);
xnor U15599 (N_15599,N_11788,N_11530);
xnor U15600 (N_15600,N_14938,N_13792);
and U15601 (N_15601,N_10525,N_14900);
or U15602 (N_15602,N_14955,N_12071);
and U15603 (N_15603,N_12812,N_10321);
nor U15604 (N_15604,N_14738,N_13816);
and U15605 (N_15605,N_13886,N_11555);
xnor U15606 (N_15606,N_12128,N_14741);
or U15607 (N_15607,N_14615,N_11887);
xor U15608 (N_15608,N_10146,N_10495);
or U15609 (N_15609,N_13482,N_11208);
nor U15610 (N_15610,N_12768,N_10696);
or U15611 (N_15611,N_10284,N_12924);
nor U15612 (N_15612,N_10390,N_10590);
or U15613 (N_15613,N_13712,N_12499);
nand U15614 (N_15614,N_14078,N_14053);
nor U15615 (N_15615,N_10429,N_12231);
or U15616 (N_15616,N_12468,N_14080);
nand U15617 (N_15617,N_13745,N_12162);
nand U15618 (N_15618,N_14118,N_13693);
or U15619 (N_15619,N_13151,N_11016);
nor U15620 (N_15620,N_13773,N_11360);
nand U15621 (N_15621,N_11825,N_13286);
xnor U15622 (N_15622,N_13058,N_13354);
nor U15623 (N_15623,N_11094,N_14748);
nor U15624 (N_15624,N_12779,N_10724);
nor U15625 (N_15625,N_10994,N_10052);
or U15626 (N_15626,N_13138,N_13100);
and U15627 (N_15627,N_10008,N_14839);
nand U15628 (N_15628,N_11413,N_14810);
or U15629 (N_15629,N_11823,N_11941);
xnor U15630 (N_15630,N_10871,N_10539);
nor U15631 (N_15631,N_13654,N_11521);
nor U15632 (N_15632,N_11658,N_10555);
xor U15633 (N_15633,N_13750,N_14222);
or U15634 (N_15634,N_13258,N_13275);
or U15635 (N_15635,N_12224,N_10666);
nor U15636 (N_15636,N_12337,N_12885);
xor U15637 (N_15637,N_12227,N_14400);
nor U15638 (N_15638,N_12742,N_12607);
nand U15639 (N_15639,N_13486,N_11647);
or U15640 (N_15640,N_14960,N_13020);
and U15641 (N_15641,N_13189,N_12561);
nand U15642 (N_15642,N_14343,N_11868);
nand U15643 (N_15643,N_14973,N_14505);
xor U15644 (N_15644,N_13329,N_11757);
xor U15645 (N_15645,N_14293,N_12286);
or U15646 (N_15646,N_13323,N_10426);
or U15647 (N_15647,N_13696,N_14433);
or U15648 (N_15648,N_14928,N_11337);
or U15649 (N_15649,N_11174,N_11770);
or U15650 (N_15650,N_14331,N_11931);
or U15651 (N_15651,N_11578,N_14140);
nor U15652 (N_15652,N_13783,N_10549);
nor U15653 (N_15653,N_14237,N_12273);
nor U15654 (N_15654,N_13160,N_12387);
xor U15655 (N_15655,N_11733,N_12042);
or U15656 (N_15656,N_10991,N_13753);
and U15657 (N_15657,N_14790,N_13305);
xnor U15658 (N_15658,N_10554,N_10959);
nor U15659 (N_15659,N_14151,N_10861);
xor U15660 (N_15660,N_12265,N_14530);
nand U15661 (N_15661,N_10143,N_10111);
nand U15662 (N_15662,N_14848,N_11186);
nor U15663 (N_15663,N_11778,N_11534);
nor U15664 (N_15664,N_12661,N_14092);
or U15665 (N_15665,N_12818,N_11003);
and U15666 (N_15666,N_12684,N_14142);
or U15667 (N_15667,N_14170,N_13970);
xor U15668 (N_15668,N_11842,N_11969);
nor U15669 (N_15669,N_11124,N_10838);
nor U15670 (N_15670,N_13607,N_13159);
xnor U15671 (N_15671,N_10816,N_12321);
and U15672 (N_15672,N_11452,N_14906);
nor U15673 (N_15673,N_13209,N_10896);
nand U15674 (N_15674,N_12570,N_14200);
nand U15675 (N_15675,N_11499,N_13983);
xor U15676 (N_15676,N_11335,N_10891);
and U15677 (N_15677,N_11060,N_10471);
or U15678 (N_15678,N_10664,N_10912);
nand U15679 (N_15679,N_14814,N_14112);
and U15680 (N_15680,N_12056,N_10580);
and U15681 (N_15681,N_14524,N_11401);
xor U15682 (N_15682,N_14632,N_14725);
nor U15683 (N_15683,N_12142,N_14284);
xor U15684 (N_15684,N_12366,N_10121);
or U15685 (N_15685,N_12605,N_14520);
or U15686 (N_15686,N_14266,N_12827);
or U15687 (N_15687,N_11357,N_14746);
or U15688 (N_15688,N_11946,N_11954);
and U15689 (N_15689,N_13144,N_13943);
nand U15690 (N_15690,N_10662,N_11947);
xor U15691 (N_15691,N_14176,N_11020);
or U15692 (N_15692,N_14660,N_12235);
or U15693 (N_15693,N_10218,N_10522);
or U15694 (N_15694,N_10864,N_10356);
xor U15695 (N_15695,N_14501,N_14067);
xnor U15696 (N_15696,N_12956,N_12739);
or U15697 (N_15697,N_11376,N_12234);
and U15698 (N_15698,N_11143,N_11872);
or U15699 (N_15699,N_10175,N_10360);
and U15700 (N_15700,N_10758,N_14832);
and U15701 (N_15701,N_12692,N_11904);
xor U15702 (N_15702,N_10683,N_11070);
nor U15703 (N_15703,N_12891,N_11718);
and U15704 (N_15704,N_10105,N_11185);
nand U15705 (N_15705,N_11248,N_12214);
xor U15706 (N_15706,N_11201,N_11024);
xor U15707 (N_15707,N_11609,N_13123);
nand U15708 (N_15708,N_10448,N_12883);
and U15709 (N_15709,N_14516,N_14037);
nand U15710 (N_15710,N_10085,N_13408);
nor U15711 (N_15711,N_10386,N_11240);
nand U15712 (N_15712,N_14249,N_12909);
xor U15713 (N_15713,N_10398,N_10591);
xnor U15714 (N_15714,N_12220,N_11167);
nor U15715 (N_15715,N_11767,N_13746);
or U15716 (N_15716,N_14771,N_12481);
or U15717 (N_15717,N_12263,N_14330);
and U15718 (N_15718,N_12085,N_10435);
xor U15719 (N_15719,N_11300,N_12958);
nand U15720 (N_15720,N_14480,N_13580);
and U15721 (N_15721,N_10748,N_13067);
nand U15722 (N_15722,N_13414,N_14945);
nor U15723 (N_15723,N_14550,N_13741);
or U15724 (N_15724,N_12438,N_12459);
nand U15725 (N_15725,N_12795,N_12123);
xnor U15726 (N_15726,N_12631,N_12663);
nor U15727 (N_15727,N_13491,N_14766);
or U15728 (N_15728,N_10878,N_11336);
xnor U15729 (N_15729,N_13183,N_10010);
nand U15730 (N_15730,N_13086,N_14665);
and U15731 (N_15731,N_14260,N_12575);
xor U15732 (N_15732,N_14085,N_10922);
nor U15733 (N_15733,N_11991,N_13797);
and U15734 (N_15734,N_11502,N_12140);
nor U15735 (N_15735,N_11148,N_11251);
nor U15736 (N_15736,N_10856,N_14298);
or U15737 (N_15737,N_11205,N_12412);
nor U15738 (N_15738,N_11144,N_10107);
nand U15739 (N_15739,N_10826,N_10062);
nand U15740 (N_15740,N_10919,N_14350);
nor U15741 (N_15741,N_13803,N_12152);
and U15742 (N_15742,N_12816,N_14511);
nand U15743 (N_15743,N_11044,N_11731);
nand U15744 (N_15744,N_13142,N_11685);
and U15745 (N_15745,N_13271,N_12865);
and U15746 (N_15746,N_12482,N_10351);
nor U15747 (N_15747,N_10513,N_13736);
nor U15748 (N_15748,N_13377,N_13052);
and U15749 (N_15749,N_11694,N_11038);
nand U15750 (N_15750,N_12048,N_10494);
nand U15751 (N_15751,N_11308,N_14683);
nor U15752 (N_15752,N_14539,N_10268);
and U15753 (N_15753,N_14394,N_11189);
nor U15754 (N_15754,N_11666,N_10131);
nand U15755 (N_15755,N_13485,N_12832);
and U15756 (N_15756,N_11507,N_11035);
xor U15757 (N_15757,N_10954,N_11249);
nand U15758 (N_15758,N_11665,N_11544);
nand U15759 (N_15759,N_14374,N_14026);
or U15760 (N_15760,N_10699,N_13064);
or U15761 (N_15761,N_12331,N_14506);
xor U15762 (N_15762,N_14235,N_13602);
xor U15763 (N_15763,N_11877,N_13785);
and U15764 (N_15764,N_11162,N_13582);
nand U15765 (N_15765,N_13945,N_13061);
nand U15766 (N_15766,N_12982,N_13706);
and U15767 (N_15767,N_12733,N_13397);
xnor U15768 (N_15768,N_13260,N_11243);
nand U15769 (N_15769,N_12002,N_13768);
nand U15770 (N_15770,N_12786,N_10865);
nor U15771 (N_15771,N_14365,N_14584);
or U15772 (N_15772,N_12659,N_10259);
nor U15773 (N_15773,N_11787,N_14723);
nand U15774 (N_15774,N_12896,N_10806);
nand U15775 (N_15775,N_12338,N_13903);
xor U15776 (N_15776,N_11807,N_13686);
and U15777 (N_15777,N_13390,N_10031);
xor U15778 (N_15778,N_13501,N_14515);
nand U15779 (N_15779,N_13977,N_12269);
nand U15780 (N_15780,N_13611,N_12504);
nor U15781 (N_15781,N_13321,N_11096);
nand U15782 (N_15782,N_14836,N_12336);
or U15783 (N_15783,N_13625,N_10493);
and U15784 (N_15784,N_13006,N_13082);
xnor U15785 (N_15785,N_11512,N_12236);
xnor U15786 (N_15786,N_10148,N_10246);
nand U15787 (N_15787,N_11423,N_12003);
nand U15788 (N_15788,N_13703,N_11591);
nor U15789 (N_15789,N_12368,N_12950);
nand U15790 (N_15790,N_11599,N_14213);
nand U15791 (N_15791,N_12067,N_12807);
and U15792 (N_15792,N_11135,N_13861);
and U15793 (N_15793,N_11829,N_10624);
or U15794 (N_15794,N_13794,N_13998);
and U15795 (N_15795,N_13776,N_10480);
xor U15796 (N_15796,N_10070,N_12259);
xor U15797 (N_15797,N_10742,N_12991);
nor U15798 (N_15798,N_14813,N_11728);
and U15799 (N_15799,N_13604,N_10104);
and U15800 (N_15800,N_11849,N_10328);
and U15801 (N_15801,N_12000,N_12147);
and U15802 (N_15802,N_11089,N_11138);
nor U15803 (N_15803,N_14543,N_13568);
and U15804 (N_15804,N_12566,N_14897);
and U15805 (N_15805,N_11776,N_14488);
and U15806 (N_15806,N_10862,N_14410);
nor U15807 (N_15807,N_10524,N_10370);
nand U15808 (N_15808,N_13986,N_11539);
or U15809 (N_15809,N_12398,N_13007);
and U15810 (N_15810,N_12884,N_14005);
and U15811 (N_15811,N_12751,N_11576);
nand U15812 (N_15812,N_13386,N_12154);
xnor U15813 (N_15813,N_11381,N_13815);
nor U15814 (N_15814,N_11321,N_13018);
nand U15815 (N_15815,N_10204,N_10629);
nand U15816 (N_15816,N_11704,N_12456);
and U15817 (N_15817,N_13907,N_14792);
xor U15818 (N_15818,N_12858,N_11573);
xnor U15819 (N_15819,N_12046,N_11808);
or U15820 (N_15820,N_12850,N_13758);
nor U15821 (N_15821,N_11702,N_10894);
and U15822 (N_15822,N_11171,N_13091);
or U15823 (N_15823,N_11256,N_13818);
and U15824 (N_15824,N_14996,N_14737);
and U15825 (N_15825,N_13202,N_12492);
and U15826 (N_15826,N_14286,N_14018);
or U15827 (N_15827,N_13558,N_11054);
nand U15828 (N_15828,N_10387,N_13224);
xor U15829 (N_15829,N_11981,N_14061);
or U15830 (N_15830,N_12964,N_12078);
xnor U15831 (N_15831,N_12882,N_10788);
and U15832 (N_15832,N_13211,N_14376);
and U15833 (N_15833,N_12919,N_14901);
and U15834 (N_15834,N_10157,N_14745);
and U15835 (N_15835,N_13667,N_14104);
xor U15836 (N_15836,N_13551,N_12820);
xor U15837 (N_15837,N_13922,N_11547);
and U15838 (N_15838,N_12489,N_10821);
and U15839 (N_15839,N_11759,N_14802);
nand U15840 (N_15840,N_11371,N_12787);
or U15841 (N_15841,N_13969,N_14173);
and U15842 (N_15842,N_14238,N_11996);
or U15843 (N_15843,N_14366,N_14066);
nand U15844 (N_15844,N_10711,N_12857);
xnor U15845 (N_15845,N_10017,N_12396);
or U15846 (N_15846,N_14346,N_11029);
nor U15847 (N_15847,N_11608,N_14486);
nand U15848 (N_15848,N_13074,N_12841);
nand U15849 (N_15849,N_12907,N_12446);
nand U15850 (N_15850,N_10137,N_11146);
and U15851 (N_15851,N_14659,N_12044);
xnor U15852 (N_15852,N_11331,N_11884);
and U15853 (N_15853,N_10152,N_12329);
nor U15854 (N_15854,N_10042,N_14734);
nor U15855 (N_15855,N_14177,N_12132);
nor U15856 (N_15856,N_12601,N_14406);
nand U15857 (N_15857,N_12737,N_10231);
or U15858 (N_15858,N_14555,N_13033);
and U15859 (N_15859,N_11848,N_13362);
and U15860 (N_15860,N_13577,N_10687);
or U15861 (N_15861,N_12299,N_11699);
and U15862 (N_15862,N_10076,N_10252);
or U15863 (N_15863,N_14440,N_11785);
nand U15864 (N_15864,N_13635,N_13695);
and U15865 (N_15865,N_10782,N_10075);
and U15866 (N_15866,N_10361,N_12798);
xor U15867 (N_15867,N_12075,N_14714);
and U15868 (N_15868,N_13266,N_10261);
nor U15869 (N_15869,N_10021,N_11226);
xor U15870 (N_15870,N_10984,N_11584);
or U15871 (N_15871,N_13641,N_14605);
nor U15872 (N_15872,N_11668,N_11930);
and U15873 (N_15873,N_12828,N_14942);
xor U15874 (N_15874,N_14476,N_11529);
and U15875 (N_15875,N_10481,N_14689);
xnor U15876 (N_15876,N_13356,N_10069);
xor U15877 (N_15877,N_14953,N_13737);
nand U15878 (N_15878,N_10305,N_10888);
nand U15879 (N_15879,N_10012,N_11327);
and U15880 (N_15880,N_14215,N_11464);
xor U15881 (N_15881,N_10465,N_11806);
nor U15882 (N_15882,N_13173,N_12988);
nand U15883 (N_15883,N_12983,N_14313);
nand U15884 (N_15884,N_10441,N_10487);
nor U15885 (N_15885,N_14301,N_11447);
or U15886 (N_15886,N_14132,N_10044);
or U15887 (N_15887,N_13523,N_10178);
nand U15888 (N_15888,N_13110,N_12996);
and U15889 (N_15889,N_11913,N_10551);
nor U15890 (N_15890,N_11293,N_14048);
or U15891 (N_15891,N_14561,N_10623);
nor U15892 (N_15892,N_11181,N_14262);
or U15893 (N_15893,N_13836,N_10837);
xnor U15894 (N_15894,N_14711,N_14527);
or U15895 (N_15895,N_12620,N_11944);
nand U15896 (N_15896,N_11565,N_11713);
xor U15897 (N_15897,N_13389,N_10598);
xnor U15898 (N_15898,N_13821,N_10442);
or U15899 (N_15899,N_11993,N_12400);
nor U15900 (N_15900,N_13811,N_12683);
or U15901 (N_15901,N_11545,N_13885);
or U15902 (N_15902,N_14401,N_13284);
nand U15903 (N_15903,N_13829,N_14983);
or U15904 (N_15904,N_12070,N_12007);
and U15905 (N_15905,N_10932,N_14111);
xnor U15906 (N_15906,N_11837,N_14348);
or U15907 (N_15907,N_12535,N_13521);
xor U15908 (N_15908,N_13479,N_13102);
nand U15909 (N_15909,N_11460,N_13480);
nand U15910 (N_15910,N_10947,N_14347);
or U15911 (N_15911,N_13718,N_14328);
nor U15912 (N_15912,N_13462,N_14599);
or U15913 (N_15913,N_11782,N_14357);
and U15914 (N_15914,N_10428,N_14158);
or U15915 (N_15915,N_13437,N_12785);
or U15916 (N_15916,N_13345,N_14425);
nor U15917 (N_15917,N_10072,N_11494);
or U15918 (N_15918,N_14658,N_14315);
nand U15919 (N_15919,N_12202,N_10258);
nand U15920 (N_15920,N_11005,N_14023);
nor U15921 (N_15921,N_13652,N_14776);
or U15922 (N_15922,N_10323,N_13388);
nand U15923 (N_15923,N_13504,N_14178);
and U15924 (N_15924,N_11492,N_13626);
and U15925 (N_15925,N_13270,N_12540);
nand U15926 (N_15926,N_13393,N_14526);
nand U15927 (N_15927,N_12198,N_12395);
xnor U15928 (N_15928,N_14470,N_10607);
nor U15929 (N_15929,N_14861,N_14058);
and U15930 (N_15930,N_10475,N_13378);
nor U15931 (N_15931,N_10595,N_10291);
and U15932 (N_15932,N_13349,N_13860);
or U15933 (N_15933,N_13541,N_14508);
or U15934 (N_15934,N_14239,N_13964);
and U15935 (N_15935,N_10566,N_10205);
and U15936 (N_15936,N_11263,N_10620);
and U15937 (N_15937,N_12374,N_10698);
xnor U15938 (N_15938,N_12420,N_10277);
or U15939 (N_15939,N_13730,N_14521);
and U15940 (N_15940,N_14608,N_10572);
and U15941 (N_15941,N_14718,N_10298);
and U15942 (N_15942,N_12444,N_13874);
nand U15943 (N_15943,N_12577,N_12125);
or U15944 (N_15944,N_11897,N_10456);
nor U15945 (N_15945,N_13166,N_14070);
or U15946 (N_15946,N_10400,N_14359);
or U15947 (N_15947,N_14884,N_13360);
nor U15948 (N_15948,N_13199,N_11907);
nand U15949 (N_15949,N_14119,N_13634);
nand U15950 (N_15950,N_10340,N_10156);
nand U15951 (N_15951,N_12704,N_10537);
nand U15952 (N_15952,N_13613,N_10354);
and U15953 (N_15953,N_11364,N_14185);
nor U15954 (N_15954,N_14229,N_12104);
and U15955 (N_15955,N_13995,N_11879);
or U15956 (N_15956,N_12941,N_13015);
xor U15957 (N_15957,N_13522,N_14949);
xor U15958 (N_15958,N_10420,N_11714);
or U15959 (N_15959,N_12775,N_11027);
nor U15960 (N_15960,N_12548,N_14464);
nand U15961 (N_15961,N_12819,N_13913);
xnor U15962 (N_15962,N_10678,N_12161);
or U15963 (N_15963,N_14398,N_12904);
and U15964 (N_15964,N_10723,N_12174);
nor U15965 (N_15965,N_12682,N_11687);
xnor U15966 (N_15966,N_14147,N_10941);
or U15967 (N_15967,N_11724,N_14234);
and U15968 (N_15968,N_10579,N_13748);
nor U15969 (N_15969,N_14130,N_10502);
nor U15970 (N_15970,N_12077,N_13217);
xnor U15971 (N_15971,N_12940,N_12435);
xor U15972 (N_15972,N_11846,N_10830);
or U15973 (N_15973,N_12881,N_12917);
nor U15974 (N_15974,N_13139,N_12599);
xnor U15975 (N_15975,N_10735,N_10569);
xor U15976 (N_15976,N_12092,N_14622);
nand U15977 (N_15977,N_13167,N_11739);
and U15978 (N_15978,N_14624,N_11062);
and U15979 (N_15979,N_14137,N_12952);
and U15980 (N_15980,N_10727,N_11551);
nand U15981 (N_15981,N_13398,N_10877);
or U15982 (N_15982,N_12409,N_13994);
nor U15983 (N_15983,N_11025,N_11633);
nand U15984 (N_15984,N_11798,N_12626);
nor U15985 (N_15985,N_11086,N_10957);
or U15986 (N_15986,N_14918,N_10395);
xor U15987 (N_15987,N_14291,N_13027);
xnor U15988 (N_15988,N_13161,N_14212);
xnor U15989 (N_15989,N_11190,N_10169);
nor U15990 (N_15990,N_13560,N_10123);
or U15991 (N_15991,N_10382,N_13565);
or U15992 (N_15992,N_14099,N_13288);
and U15993 (N_15993,N_10043,N_11400);
and U15994 (N_15994,N_12763,N_14003);
nand U15995 (N_15995,N_11277,N_14916);
or U15996 (N_15996,N_10792,N_13353);
nand U15997 (N_15997,N_12730,N_13188);
or U15998 (N_15998,N_10074,N_11719);
or U15999 (N_15999,N_10951,N_14821);
nor U16000 (N_16000,N_12686,N_10504);
or U16001 (N_16001,N_12488,N_12750);
xor U16002 (N_16002,N_11352,N_12445);
or U16003 (N_16003,N_11577,N_12702);
and U16004 (N_16004,N_14692,N_11388);
or U16005 (N_16005,N_14713,N_12475);
or U16006 (N_16006,N_12736,N_14671);
nand U16007 (N_16007,N_13512,N_11527);
nand U16008 (N_16008,N_11833,N_14872);
and U16009 (N_16009,N_11018,N_12210);
or U16010 (N_16010,N_14141,N_13307);
nand U16011 (N_16011,N_10177,N_14392);
nand U16012 (N_16012,N_11655,N_14153);
xnor U16013 (N_16013,N_12130,N_10918);
and U16014 (N_16014,N_13325,N_10654);
nand U16015 (N_16015,N_11766,N_10596);
nand U16016 (N_16016,N_13592,N_11734);
or U16017 (N_16017,N_14822,N_11566);
or U16018 (N_16018,N_11588,N_13890);
or U16019 (N_16019,N_12993,N_13467);
or U16020 (N_16020,N_13990,N_11199);
nand U16021 (N_16021,N_13302,N_13333);
xnor U16022 (N_16022,N_14154,N_13385);
nand U16023 (N_16023,N_12851,N_10674);
nand U16024 (N_16024,N_11260,N_13834);
and U16025 (N_16025,N_13691,N_13342);
nand U16026 (N_16026,N_11032,N_11789);
nand U16027 (N_16027,N_12772,N_12306);
nand U16028 (N_16028,N_12844,N_14703);
nand U16029 (N_16029,N_14253,N_10739);
xnor U16030 (N_16030,N_11792,N_10560);
and U16031 (N_16031,N_10728,N_11087);
nand U16032 (N_16032,N_14449,N_11160);
or U16033 (N_16033,N_10375,N_12110);
and U16034 (N_16034,N_14812,N_10176);
nor U16035 (N_16035,N_13177,N_12707);
and U16036 (N_16036,N_12796,N_12848);
xnor U16037 (N_16037,N_13090,N_12094);
xnor U16038 (N_16038,N_13172,N_10235);
nor U16039 (N_16039,N_14558,N_13774);
and U16040 (N_16040,N_14698,N_14708);
xnor U16041 (N_16041,N_14199,N_10834);
nand U16042 (N_16042,N_12549,N_10245);
nor U16043 (N_16043,N_12998,N_11291);
xor U16044 (N_16044,N_14627,N_13081);
nor U16045 (N_16045,N_10421,N_10995);
nand U16046 (N_16046,N_13835,N_10632);
xor U16047 (N_16047,N_11406,N_10884);
and U16048 (N_16048,N_12773,N_12051);
nand U16049 (N_16049,N_11937,N_12671);
and U16050 (N_16050,N_13632,N_11325);
nand U16051 (N_16051,N_10874,N_13870);
nor U16052 (N_16052,N_12278,N_13201);
nand U16053 (N_16053,N_14712,N_14739);
and U16054 (N_16054,N_11478,N_13174);
or U16055 (N_16055,N_14214,N_11859);
nor U16056 (N_16056,N_13946,N_10545);
nor U16057 (N_16057,N_11479,N_14389);
or U16058 (N_16058,N_12582,N_10650);
nor U16059 (N_16059,N_14740,N_10103);
nor U16060 (N_16060,N_12017,N_13493);
nor U16061 (N_16061,N_12621,N_13527);
nand U16062 (N_16062,N_11519,N_13171);
or U16063 (N_16063,N_13952,N_12568);
nor U16064 (N_16064,N_13181,N_11330);
nand U16065 (N_16065,N_14335,N_12300);
nor U16066 (N_16066,N_13936,N_11903);
or U16067 (N_16067,N_11428,N_10557);
and U16068 (N_16068,N_14143,N_13727);
or U16069 (N_16069,N_12806,N_10160);
nor U16070 (N_16070,N_10172,N_12871);
nor U16071 (N_16071,N_14730,N_10015);
or U16072 (N_16072,N_14377,N_12421);
nor U16073 (N_16073,N_12134,N_12280);
nor U16074 (N_16074,N_14845,N_14198);
xnor U16075 (N_16075,N_14485,N_10531);
nor U16076 (N_16076,N_12769,N_11511);
and U16077 (N_16077,N_12487,N_11886);
nand U16078 (N_16078,N_12188,N_14162);
nor U16079 (N_16079,N_12089,N_14681);
or U16080 (N_16080,N_11559,N_13472);
nor U16081 (N_16081,N_14064,N_12246);
or U16082 (N_16082,N_14598,N_12866);
or U16083 (N_16083,N_13496,N_11109);
xor U16084 (N_16084,N_14552,N_10584);
nor U16085 (N_16085,N_13516,N_12284);
xnor U16086 (N_16086,N_11437,N_10612);
nand U16087 (N_16087,N_14093,N_12644);
nand U16088 (N_16088,N_13978,N_11622);
nor U16089 (N_16089,N_13474,N_12464);
xor U16090 (N_16090,N_14705,N_11121);
xnor U16091 (N_16091,N_11074,N_12647);
xnor U16092 (N_16092,N_13459,N_14157);
nand U16093 (N_16093,N_13967,N_12441);
or U16094 (N_16094,N_13427,N_12756);
nor U16095 (N_16095,N_11572,N_14261);
nor U16096 (N_16096,N_10353,N_13228);
xnor U16097 (N_16097,N_13658,N_13182);
xor U16098 (N_16098,N_11557,N_11505);
nor U16099 (N_16099,N_11593,N_13428);
xnor U16100 (N_16100,N_11495,N_10180);
nor U16101 (N_16101,N_14509,N_10597);
nor U16102 (N_16102,N_12845,N_12431);
nor U16103 (N_16103,N_12155,N_10225);
nand U16104 (N_16104,N_14224,N_13751);
nor U16105 (N_16105,N_14582,N_12632);
xor U16106 (N_16106,N_10073,N_13618);
or U16107 (N_16107,N_14937,N_12143);
nor U16108 (N_16108,N_12555,N_13760);
xor U16109 (N_16109,N_13005,N_11184);
and U16110 (N_16110,N_12428,N_13158);
nor U16111 (N_16111,N_14800,N_14882);
or U16112 (N_16112,N_13303,N_13331);
xor U16113 (N_16113,N_11425,N_12016);
nand U16114 (N_16114,N_14923,N_10610);
nor U16115 (N_16115,N_14251,N_11100);
xnor U16116 (N_16116,N_12526,N_10182);
and U16117 (N_16117,N_14014,N_13530);
and U16118 (N_16118,N_13599,N_13949);
xor U16119 (N_16119,N_13755,N_11077);
or U16120 (N_16120,N_13884,N_11870);
nand U16121 (N_16121,N_11052,N_10346);
or U16122 (N_16122,N_13947,N_14450);
nor U16123 (N_16123,N_14091,N_12285);
and U16124 (N_16124,N_13678,N_13419);
or U16125 (N_16125,N_13195,N_11532);
or U16126 (N_16126,N_13546,N_11164);
and U16127 (N_16127,N_14172,N_13358);
or U16128 (N_16128,N_13476,N_12467);
nor U16129 (N_16129,N_14351,N_12382);
and U16130 (N_16130,N_10986,N_12915);
nor U16131 (N_16131,N_11332,N_11819);
xor U16132 (N_16132,N_13804,N_14952);
nor U16133 (N_16133,N_14065,N_14021);
xnor U16134 (N_16134,N_10068,N_13784);
nor U16135 (N_16135,N_11216,N_14586);
nor U16136 (N_16136,N_14397,N_10606);
xnor U16137 (N_16137,N_12211,N_10022);
and U16138 (N_16138,N_11014,N_12418);
xor U16139 (N_16139,N_14383,N_10499);
and U16140 (N_16140,N_10841,N_12453);
nand U16141 (N_16141,N_12345,N_10538);
nor U16142 (N_16142,N_12113,N_10125);
nand U16143 (N_16143,N_14929,N_12451);
or U16144 (N_16144,N_13926,N_11422);
and U16145 (N_16145,N_10731,N_11061);
or U16146 (N_16146,N_11514,N_12765);
or U16147 (N_16147,N_12159,N_14393);
nor U16148 (N_16148,N_10581,N_11355);
xor U16149 (N_16149,N_12018,N_13253);
or U16150 (N_16150,N_13620,N_13403);
and U16151 (N_16151,N_14378,N_10329);
nand U16152 (N_16152,N_13916,N_12972);
or U16153 (N_16153,N_13537,N_11711);
nor U16154 (N_16154,N_13383,N_10616);
nor U16155 (N_16155,N_10903,N_12674);
xnor U16156 (N_16156,N_10847,N_12588);
or U16157 (N_16157,N_13498,N_11596);
xor U16158 (N_16158,N_12373,N_13263);
nor U16159 (N_16159,N_12515,N_12762);
and U16160 (N_16160,N_14146,N_13155);
nand U16161 (N_16161,N_12030,N_14647);
xnor U16162 (N_16162,N_14006,N_12606);
or U16163 (N_16163,N_11193,N_12486);
and U16164 (N_16164,N_12053,N_14327);
nand U16165 (N_16165,N_14693,N_13059);
nand U16166 (N_16166,N_12927,N_12401);
nor U16167 (N_16167,N_10892,N_12701);
xnor U16168 (N_16168,N_10673,N_12745);
and U16169 (N_16169,N_14420,N_13690);
nand U16170 (N_16170,N_13764,N_14761);
nand U16171 (N_16171,N_12556,N_11561);
nor U16172 (N_16172,N_10439,N_11454);
or U16173 (N_16173,N_13092,N_13865);
nor U16174 (N_16174,N_12932,N_14273);
and U16175 (N_16175,N_13772,N_11282);
or U16176 (N_16176,N_12529,N_11786);
or U16177 (N_16177,N_10615,N_13105);
and U16178 (N_16178,N_13028,N_11140);
nor U16179 (N_16179,N_10814,N_10479);
xor U16180 (N_16180,N_13848,N_12987);
nor U16181 (N_16181,N_10953,N_10857);
xnor U16182 (N_16182,N_13854,N_12245);
nor U16183 (N_16183,N_11900,N_14715);
nor U16184 (N_16184,N_10985,N_10697);
nor U16185 (N_16185,N_12562,N_14369);
xor U16186 (N_16186,N_10424,N_12951);
or U16187 (N_16187,N_11709,N_10902);
and U16188 (N_16188,N_10938,N_14667);
and U16189 (N_16189,N_12861,N_14231);
xnor U16190 (N_16190,N_11775,N_12718);
nand U16191 (N_16191,N_10600,N_13084);
nand U16192 (N_16192,N_10592,N_13441);
nand U16193 (N_16193,N_13357,N_11592);
or U16194 (N_16194,N_10241,N_13534);
nand U16195 (N_16195,N_12112,N_13763);
or U16196 (N_16196,N_10036,N_10047);
and U16197 (N_16197,N_10914,N_14493);
xor U16198 (N_16198,N_14468,N_13665);
nor U16199 (N_16199,N_13674,N_10844);
xnor U16200 (N_16200,N_10714,N_12645);
or U16201 (N_16201,N_11434,N_13338);
nor U16202 (N_16202,N_11353,N_14935);
xnor U16203 (N_16203,N_10474,N_11290);
xnor U16204 (N_16204,N_11176,N_12842);
and U16205 (N_16205,N_12189,N_14166);
or U16206 (N_16206,N_10163,N_14793);
or U16207 (N_16207,N_14631,N_13346);
or U16208 (N_16208,N_11594,N_13770);
and U16209 (N_16209,N_13833,N_10061);
nand U16210 (N_16210,N_13162,N_13603);
or U16211 (N_16211,N_12835,N_11329);
nor U16212 (N_16212,N_11469,N_12425);
and U16213 (N_16213,N_10923,N_12984);
or U16214 (N_16214,N_11311,N_10764);
or U16215 (N_16215,N_11132,N_11139);
nor U16216 (N_16216,N_12740,N_14255);
nand U16217 (N_16217,N_14028,N_14254);
and U16218 (N_16218,N_11838,N_14205);
and U16219 (N_16219,N_10355,N_14860);
or U16220 (N_16220,N_14460,N_13101);
nand U16221 (N_16221,N_13348,N_10336);
nand U16222 (N_16222,N_12942,N_11057);
and U16223 (N_16223,N_10263,N_10689);
and U16224 (N_16224,N_12793,N_14545);
nor U16225 (N_16225,N_13235,N_14859);
nand U16226 (N_16226,N_13252,N_14551);
or U16227 (N_16227,N_10497,N_14830);
xor U16228 (N_16228,N_13344,N_13689);
xnor U16229 (N_16229,N_11689,N_14134);
or U16230 (N_16230,N_12058,N_12895);
or U16231 (N_16231,N_11804,N_14887);
nand U16232 (N_16232,N_14536,N_13475);
or U16233 (N_16233,N_11007,N_12314);
and U16234 (N_16234,N_14175,N_11628);
nor U16235 (N_16235,N_14069,N_10407);
nor U16236 (N_16236,N_10972,N_12239);
nor U16237 (N_16237,N_13017,N_14340);
xor U16238 (N_16238,N_14358,N_12789);
and U16239 (N_16239,N_10437,N_13488);
and U16240 (N_16240,N_14557,N_11586);
or U16241 (N_16241,N_10159,N_12355);
nor U16242 (N_16242,N_12872,N_10149);
and U16243 (N_16243,N_12494,N_11049);
or U16244 (N_16244,N_11809,N_10963);
and U16245 (N_16245,N_10081,N_12990);
nand U16246 (N_16246,N_12213,N_12384);
nand U16247 (N_16247,N_14649,N_11625);
xnor U16248 (N_16248,N_13707,N_10415);
xor U16249 (N_16249,N_13662,N_14290);
nand U16250 (N_16250,N_10288,N_10009);
or U16251 (N_16251,N_14931,N_11537);
and U16252 (N_16252,N_14271,N_14994);
xor U16253 (N_16253,N_14306,N_14613);
and U16254 (N_16254,N_12979,N_11169);
xnor U16255 (N_16255,N_12032,N_14430);
nand U16256 (N_16256,N_13456,N_10643);
and U16257 (N_16257,N_14441,N_13249);
xnor U16258 (N_16258,N_14316,N_10546);
nor U16259 (N_16259,N_11546,N_10535);
and U16260 (N_16260,N_13571,N_10381);
or U16261 (N_16261,N_14041,N_11717);
nor U16262 (N_16262,N_13511,N_10452);
and U16263 (N_16263,N_14352,N_10835);
nor U16264 (N_16264,N_14297,N_10083);
and U16265 (N_16265,N_11420,N_11046);
or U16266 (N_16266,N_10034,N_10469);
or U16267 (N_16267,N_12874,N_10174);
and U16268 (N_16268,N_10970,N_12594);
nor U16269 (N_16269,N_12696,N_13119);
or U16270 (N_16270,N_13226,N_13069);
nor U16271 (N_16271,N_14870,N_13553);
nand U16272 (N_16272,N_14933,N_12592);
nand U16273 (N_16273,N_14436,N_14767);
xor U16274 (N_16274,N_10196,N_14190);
or U16275 (N_16275,N_10547,N_14743);
and U16276 (N_16276,N_11209,N_12417);
nand U16277 (N_16277,N_12797,N_11015);
nor U16278 (N_16278,N_14183,N_13118);
xnor U16279 (N_16279,N_13777,N_11976);
and U16280 (N_16280,N_13781,N_10997);
xor U16281 (N_16281,N_11754,N_12929);
nand U16282 (N_16282,N_14744,N_12478);
and U16283 (N_16283,N_14674,N_12864);
and U16284 (N_16284,N_13590,N_14090);
xor U16285 (N_16285,N_11227,N_12680);
xnor U16286 (N_16286,N_10254,N_13614);
and U16287 (N_16287,N_11198,N_13991);
nand U16288 (N_16288,N_12179,N_11429);
nor U16289 (N_16289,N_11800,N_14907);
nor U16290 (N_16290,N_12860,N_14697);
or U16291 (N_16291,N_10067,N_12139);
and U16292 (N_16292,N_10040,N_14528);
or U16293 (N_16293,N_10374,N_10603);
xor U16294 (N_16294,N_11150,N_14597);
nand U16295 (N_16295,N_13672,N_10393);
nand U16296 (N_16296,N_10165,N_13175);
nand U16297 (N_16297,N_10655,N_11660);
and U16298 (N_16298,N_10516,N_10399);
xor U16299 (N_16299,N_12407,N_10214);
nor U16300 (N_16300,N_14880,N_14589);
and U16301 (N_16301,N_13026,N_14975);
nor U16302 (N_16302,N_14862,N_14865);
xor U16303 (N_16303,N_13369,N_13808);
nor U16304 (N_16304,N_10568,N_11925);
and U16305 (N_16305,N_12318,N_12830);
nand U16306 (N_16306,N_11281,N_12821);
nand U16307 (N_16307,N_13705,N_10800);
xnor U16308 (N_16308,N_13557,N_11154);
nor U16309 (N_16309,N_10824,N_12595);
nor U16310 (N_16310,N_13901,N_11750);
nand U16311 (N_16311,N_13131,N_11563);
or U16312 (N_16312,N_10799,N_10158);
or U16313 (N_16313,N_11009,N_10028);
or U16314 (N_16314,N_12590,N_11523);
nand U16315 (N_16315,N_11246,N_10286);
and U16316 (N_16316,N_10496,N_12172);
xnor U16317 (N_16317,N_12356,N_13363);
and U16318 (N_16318,N_14088,N_10003);
xnor U16319 (N_16319,N_12653,N_11997);
xor U16320 (N_16320,N_12817,N_14274);
or U16321 (N_16321,N_13631,N_13518);
nand U16322 (N_16322,N_12706,N_10519);
xor U16323 (N_16323,N_10946,N_11621);
nand U16324 (N_16324,N_12274,N_13925);
xor U16325 (N_16325,N_11202,N_14927);
nor U16326 (N_16326,N_14265,N_14854);
xnor U16327 (N_16327,N_13515,N_14372);
xnor U16328 (N_16328,N_13623,N_14637);
or U16329 (N_16329,N_13968,N_11334);
nand U16330 (N_16330,N_12439,N_11387);
nor U16331 (N_16331,N_14164,N_12905);
nand U16332 (N_16332,N_14439,N_13099);
xor U16333 (N_16333,N_10934,N_12332);
or U16334 (N_16334,N_13276,N_11783);
xor U16335 (N_16335,N_11157,N_14760);
or U16336 (N_16336,N_11365,N_13261);
xnor U16337 (N_16337,N_10979,N_13608);
nor U16338 (N_16338,N_12200,N_10477);
or U16339 (N_16339,N_13012,N_11698);
xor U16340 (N_16340,N_14421,N_10425);
and U16341 (N_16341,N_13085,N_12749);
nand U16342 (N_16342,N_12547,N_13197);
nor U16343 (N_16343,N_10803,N_11088);
and U16344 (N_16344,N_14305,N_12145);
nand U16345 (N_16345,N_11481,N_10810);
or U16346 (N_16346,N_14595,N_13767);
nand U16347 (N_16347,N_12700,N_11446);
xnor U16348 (N_16348,N_14423,N_12802);
nor U16349 (N_16349,N_13315,N_14367);
nand U16350 (N_16350,N_11328,N_14742);
xnor U16351 (N_16351,N_14196,N_10944);
and U16352 (N_16352,N_12442,N_12877);
xor U16353 (N_16353,N_12727,N_11471);
nor U16354 (N_16354,N_10344,N_13022);
nand U16355 (N_16355,N_14124,N_12219);
or U16356 (N_16356,N_12449,N_11294);
nand U16357 (N_16357,N_10162,N_11093);
nor U16358 (N_16358,N_14876,N_12799);
xnor U16359 (N_16359,N_12153,N_12826);
nor U16360 (N_16360,N_14611,N_12006);
or U16361 (N_16361,N_10670,N_11562);
nor U16362 (N_16362,N_10515,N_13359);
and U16363 (N_16363,N_12181,N_13128);
nor U16364 (N_16364,N_13207,N_13905);
xor U16365 (N_16365,N_14993,N_13111);
nor U16366 (N_16366,N_13236,N_11103);
nor U16367 (N_16367,N_12339,N_10691);
xnor U16368 (N_16368,N_13578,N_11344);
or U16369 (N_16369,N_13891,N_12576);
xnor U16370 (N_16370,N_12238,N_10438);
nand U16371 (N_16371,N_10829,N_12257);
or U16372 (N_16372,N_13238,N_13698);
or U16373 (N_16373,N_11771,N_12287);
nand U16374 (N_16374,N_13610,N_13757);
or U16375 (N_16375,N_10279,N_12497);
and U16376 (N_16376,N_13850,N_13559);
nor U16377 (N_16377,N_11784,N_14094);
and U16378 (N_16378,N_10485,N_12681);
xor U16379 (N_16379,N_14987,N_11610);
xor U16380 (N_16380,N_11632,N_10609);
nand U16381 (N_16381,N_10766,N_10679);
xnor U16382 (N_16382,N_12703,N_13810);
nand U16383 (N_16383,N_12888,N_14673);
or U16384 (N_16384,N_14602,N_11111);
nor U16385 (N_16385,N_12638,N_12926);
or U16386 (N_16386,N_13149,N_10256);
nand U16387 (N_16387,N_14182,N_12550);
or U16388 (N_16388,N_13231,N_13646);
nor U16389 (N_16389,N_10893,N_13230);
nand U16390 (N_16390,N_12025,N_12215);
and U16391 (N_16391,N_10283,N_11503);
xor U16392 (N_16392,N_13595,N_10508);
and U16393 (N_16393,N_10188,N_12546);
and U16394 (N_16394,N_10754,N_13180);
or U16395 (N_16395,N_12591,N_12206);
nand U16396 (N_16396,N_14915,N_12849);
nand U16397 (N_16397,N_10223,N_12379);
xnor U16398 (N_16398,N_12694,N_12501);
nand U16399 (N_16399,N_12362,N_12608);
or U16400 (N_16400,N_11664,N_13570);
nor U16401 (N_16401,N_13668,N_13554);
nand U16402 (N_16402,N_13444,N_10109);
or U16403 (N_16403,N_10775,N_13845);
and U16404 (N_16404,N_12496,N_13719);
nand U16405 (N_16405,N_11475,N_12552);
nor U16406 (N_16406,N_11021,N_12322);
or U16407 (N_16407,N_14553,N_12754);
or U16408 (N_16408,N_14110,N_12434);
nand U16409 (N_16409,N_11987,N_11163);
or U16410 (N_16410,N_10132,N_12129);
nor U16411 (N_16411,N_12939,N_12900);
and U16412 (N_16412,N_11738,N_14787);
nand U16413 (N_16413,N_11156,N_13040);
or U16414 (N_16414,N_10686,N_11456);
nor U16415 (N_16415,N_12610,N_13274);
nand U16416 (N_16416,N_11878,N_12308);
and U16417 (N_16417,N_10467,N_10904);
xnor U16418 (N_16418,N_13716,N_11367);
and U16419 (N_16419,N_10753,N_14010);
and U16420 (N_16420,N_12333,N_12301);
nor U16421 (N_16421,N_12183,N_14577);
nand U16422 (N_16422,N_13379,N_12063);
nand U16423 (N_16423,N_13852,N_10020);
and U16424 (N_16424,N_10977,N_10588);
nor U16425 (N_16425,N_10266,N_14483);
and U16426 (N_16426,N_11081,N_14857);
or U16427 (N_16427,N_12101,N_11113);
and U16428 (N_16428,N_10680,N_10369);
or U16429 (N_16429,N_10380,N_10106);
and U16430 (N_16430,N_14382,N_10721);
and U16431 (N_16431,N_10743,N_13550);
xor U16432 (N_16432,N_14240,N_11542);
xor U16433 (N_16433,N_12004,N_13984);
xor U16434 (N_16434,N_10542,N_11570);
xnor U16435 (N_16435,N_10726,N_12953);
nor U16436 (N_16436,N_10364,N_13682);
or U16437 (N_16437,N_11580,N_10491);
nand U16438 (N_16438,N_11416,N_10565);
xor U16439 (N_16439,N_14844,N_14181);
xor U16440 (N_16440,N_11729,N_13509);
or U16441 (N_16441,N_14399,N_12688);
or U16442 (N_16442,N_10505,N_10897);
and U16443 (N_16443,N_14656,N_11497);
nand U16444 (N_16444,N_14808,N_14381);
nand U16445 (N_16445,N_11843,N_10868);
or U16446 (N_16446,N_14495,N_13367);
nand U16447 (N_16447,N_13843,N_11708);
nand U16448 (N_16448,N_13561,N_10151);
or U16449 (N_16449,N_10450,N_14684);
or U16450 (N_16450,N_14560,N_14604);
nand U16451 (N_16451,N_12237,N_10880);
or U16452 (N_16452,N_14494,N_14736);
nor U16453 (N_16453,N_12436,N_10732);
and U16454 (N_16454,N_14283,N_13908);
and U16455 (N_16455,N_10099,N_10924);
or U16456 (N_16456,N_12312,N_13281);
nor U16457 (N_16457,N_14601,N_10309);
and U16458 (N_16458,N_13300,N_10736);
nand U16459 (N_16459,N_10998,N_10197);
or U16460 (N_16460,N_12995,N_12767);
and U16461 (N_16461,N_10454,N_14384);
xor U16462 (N_16462,N_10712,N_12124);
nand U16463 (N_16463,N_14803,N_12082);
or U16464 (N_16464,N_11126,N_12248);
and U16465 (N_16465,N_10388,N_10787);
and U16466 (N_16466,N_14120,N_14108);
nand U16467 (N_16467,N_10147,N_13332);
nor U16468 (N_16468,N_11010,N_10540);
xor U16469 (N_16469,N_11936,N_11223);
or U16470 (N_16470,N_14666,N_13470);
nand U16471 (N_16471,N_12985,N_13347);
nor U16472 (N_16472,N_10423,N_13780);
and U16473 (N_16473,N_14363,N_13831);
xnor U16474 (N_16474,N_12560,N_14786);
xnor U16475 (N_16475,N_11696,N_14523);
nor U16476 (N_16476,N_12513,N_13729);
nor U16477 (N_16477,N_12992,N_13361);
nor U16478 (N_16478,N_13538,N_12057);
nor U16479 (N_16479,N_13114,N_10281);
and U16480 (N_16480,N_12375,N_14000);
and U16481 (N_16481,N_13241,N_13814);
and U16482 (N_16482,N_13483,N_10451);
and U16483 (N_16483,N_12973,N_14211);
and U16484 (N_16484,N_13857,N_13203);
nor U16485 (N_16485,N_13233,N_14716);
or U16486 (N_16486,N_10293,N_10265);
xnor U16487 (N_16487,N_12187,N_10534);
or U16488 (N_16488,N_11774,N_10192);
and U16489 (N_16489,N_11305,N_13449);
xor U16490 (N_16490,N_10331,N_13198);
and U16491 (N_16491,N_12629,N_13871);
and U16492 (N_16492,N_10571,N_10213);
xor U16493 (N_16493,N_12690,N_10005);
and U16494 (N_16494,N_10371,N_11642);
xnor U16495 (N_16495,N_11212,N_11746);
or U16496 (N_16496,N_11526,N_14139);
or U16497 (N_16497,N_13402,N_12173);
nand U16498 (N_16498,N_13918,N_13944);
nand U16499 (N_16499,N_14115,N_10614);
or U16500 (N_16500,N_13627,N_10334);
and U16501 (N_16501,N_11543,N_13973);
nor U16502 (N_16502,N_12087,N_12228);
xor U16503 (N_16503,N_10992,N_14025);
xnor U16504 (N_16504,N_10532,N_12020);
nor U16505 (N_16505,N_14532,N_10526);
nand U16506 (N_16506,N_14186,N_13376);
nand U16507 (N_16507,N_14161,N_14033);
or U16508 (N_16508,N_14413,N_12427);
nand U16509 (N_16509,N_12151,N_11273);
nand U16510 (N_16510,N_11358,N_10405);
or U16511 (N_16511,N_11672,N_14074);
nor U16512 (N_16512,N_10789,N_11510);
nand U16513 (N_16513,N_11261,N_12498);
nor U16514 (N_16514,N_11182,N_12724);
and U16515 (N_16515,N_10665,N_13639);
xor U16516 (N_16516,N_12551,N_13892);
and U16517 (N_16517,N_11763,N_14349);
nand U16518 (N_16518,N_11449,N_10949);
nand U16519 (N_16519,N_14902,N_10744);
xnor U16520 (N_16520,N_11112,N_11033);
or U16521 (N_16521,N_13649,N_14267);
xor U16522 (N_16522,N_13896,N_12673);
and U16523 (N_16523,N_12965,N_13642);
or U16524 (N_16524,N_13809,N_13269);
xnor U16525 (N_16525,N_12116,N_12121);
xnor U16526 (N_16526,N_13039,N_13636);
or U16527 (N_16527,N_12126,N_12021);
or U16528 (N_16528,N_10635,N_12028);
xor U16529 (N_16529,N_10769,N_12536);
nand U16530 (N_16530,N_14640,N_12293);
nand U16531 (N_16531,N_14287,N_10693);
and U16532 (N_16532,N_11899,N_11483);
nand U16533 (N_16533,N_13827,N_13875);
or U16534 (N_16534,N_11187,N_14054);
xor U16535 (N_16535,N_11635,N_11926);
and U16536 (N_16536,N_11071,N_13279);
or U16537 (N_16537,N_10230,N_12669);
and U16538 (N_16538,N_11433,N_11490);
nand U16539 (N_16539,N_13935,N_12455);
xnor U16540 (N_16540,N_11630,N_12572);
nor U16541 (N_16541,N_14103,N_12491);
or U16542 (N_16542,N_11307,N_10094);
or U16543 (N_16543,N_13953,N_11888);
and U16544 (N_16544,N_12977,N_14852);
nand U16545 (N_16545,N_11541,N_12868);
nor U16546 (N_16546,N_13671,N_11224);
nand U16547 (N_16547,N_11192,N_11973);
nand U16548 (N_16548,N_13644,N_11894);
nand U16549 (N_16549,N_12422,N_13791);
and U16550 (N_16550,N_10745,N_12165);
and U16551 (N_16551,N_14634,N_10668);
and U16552 (N_16552,N_13277,N_12343);
or U16553 (N_16553,N_14541,N_13384);
or U16554 (N_16554,N_13825,N_13251);
nor U16555 (N_16555,N_13598,N_10278);
or U16556 (N_16556,N_11065,N_11813);
or U16557 (N_16557,N_12452,N_12167);
nor U16558 (N_16558,N_14454,N_10133);
or U16559 (N_16559,N_14858,N_14275);
and U16560 (N_16560,N_13999,N_10750);
nor U16561 (N_16561,N_12666,N_12330);
nand U16562 (N_16562,N_13869,N_10895);
nor U16563 (N_16563,N_10958,N_13859);
or U16564 (N_16564,N_11242,N_14339);
xor U16565 (N_16565,N_10419,N_14912);
nand U16566 (N_16566,N_12521,N_14850);
and U16567 (N_16567,N_11945,N_13616);
or U16568 (N_16568,N_10889,N_10077);
or U16569 (N_16569,N_13218,N_14921);
nand U16570 (N_16570,N_13771,N_10296);
or U16571 (N_16571,N_10023,N_14309);
nor U16572 (N_16572,N_10102,N_12935);
xor U16573 (N_16573,N_10316,N_13268);
nand U16574 (N_16574,N_10206,N_13979);
xnor U16575 (N_16575,N_11239,N_14799);
nor U16576 (N_16576,N_11558,N_10929);
nor U16577 (N_16577,N_12778,N_12836);
and U16578 (N_16578,N_11129,N_11673);
nand U16579 (N_16579,N_12074,N_13121);
xor U16580 (N_16580,N_12911,N_11615);
nand U16581 (N_16581,N_12824,N_10906);
xor U16582 (N_16582,N_14966,N_10622);
and U16583 (N_16583,N_14308,N_14345);
or U16584 (N_16584,N_11426,N_11442);
or U16585 (N_16585,N_14893,N_11548);
xor U16586 (N_16586,N_13051,N_13976);
nor U16587 (N_16587,N_10853,N_11742);
nor U16588 (N_16588,N_10112,N_14578);
and U16589 (N_16589,N_14012,N_12846);
nand U16590 (N_16590,N_11161,N_13789);
xor U16591 (N_16591,N_14758,N_12001);
xor U16592 (N_16592,N_11727,N_11309);
nor U16593 (N_16593,N_10634,N_12792);
xnor U16594 (N_16594,N_13413,N_10640);
and U16595 (N_16595,N_10349,N_14596);
nor U16596 (N_16596,N_13638,N_11439);
xor U16597 (N_16597,N_14571,N_14784);
nand U16598 (N_16598,N_13839,N_14481);
nand U16599 (N_16599,N_12981,N_11128);
xnor U16600 (N_16600,N_13322,N_13982);
nor U16601 (N_16601,N_11747,N_14556);
or U16602 (N_16602,N_13340,N_14773);
nand U16603 (N_16603,N_11560,N_10675);
or U16604 (N_16604,N_11229,N_12528);
or U16605 (N_16605,N_12554,N_14569);
or U16606 (N_16606,N_14968,N_11191);
nand U16607 (N_16607,N_13997,N_12719);
or U16608 (N_16608,N_10937,N_11002);
nand U16609 (N_16609,N_10983,N_10366);
or U16610 (N_16610,N_10056,N_11149);
xor U16611 (N_16611,N_12296,N_13146);
or U16612 (N_16612,N_13156,N_14579);
xor U16613 (N_16613,N_13853,N_14646);
nand U16614 (N_16614,N_12959,N_11399);
nor U16615 (N_16615,N_13137,N_10041);
or U16616 (N_16616,N_10128,N_10511);
nand U16617 (N_16617,N_10341,N_14819);
nand U16618 (N_16618,N_11623,N_11278);
xnor U16619 (N_16619,N_11606,N_11927);
nand U16620 (N_16620,N_13941,N_10653);
xnor U16621 (N_16621,N_13337,N_14944);
or U16622 (N_16622,N_11265,N_14129);
nor U16623 (N_16623,N_12283,N_11474);
xor U16624 (N_16624,N_12348,N_11871);
nor U16625 (N_16625,N_12111,N_13801);
or U16626 (N_16626,N_10232,N_10087);
or U16627 (N_16627,N_12957,N_13135);
nor U16628 (N_16628,N_12261,N_13531);
xor U16629 (N_16629,N_10911,N_13453);
nor U16630 (N_16630,N_11920,N_13239);
nand U16631 (N_16631,N_12879,N_10701);
or U16632 (N_16632,N_12839,N_10242);
xnor U16633 (N_16633,N_12349,N_11348);
nand U16634 (N_16634,N_11462,N_12282);
and U16635 (N_16635,N_12426,N_14491);
nand U16636 (N_16636,N_11461,N_11605);
nor U16637 (N_16637,N_11516,N_13216);
and U16638 (N_16638,N_12100,N_13732);
nand U16639 (N_16639,N_13939,N_12712);
or U16640 (N_16640,N_11928,N_11142);
xor U16641 (N_16641,N_10413,N_14783);
nand U16642 (N_16642,N_10567,N_13287);
xnor U16643 (N_16643,N_12753,N_10319);
and U16644 (N_16644,N_13416,N_13237);
xnor U16645 (N_16645,N_10663,N_14412);
and U16646 (N_16646,N_11354,N_14920);
nor U16647 (N_16647,N_14831,N_13368);
nand U16648 (N_16648,N_11670,N_10899);
and U16649 (N_16649,N_12065,N_12831);
and U16650 (N_16650,N_10682,N_12761);
nand U16651 (N_16651,N_13194,N_10577);
xnor U16652 (N_16652,N_12569,N_11518);
nor U16653 (N_16653,N_14497,N_14762);
xor U16654 (N_16654,N_11234,N_11465);
xnor U16655 (N_16655,N_10900,N_11383);
nand U16656 (N_16656,N_13254,N_12726);
xor U16657 (N_16657,N_14168,N_10765);
xor U16658 (N_16658,N_14009,N_10962);
and U16659 (N_16659,N_11553,N_13813);
and U16660 (N_16660,N_11179,N_12735);
and U16661 (N_16661,N_11232,N_10621);
nor U16662 (N_16662,N_14540,N_11604);
xnor U16663 (N_16663,N_14898,N_12357);
or U16664 (N_16664,N_13257,N_10869);
or U16665 (N_16665,N_11509,N_13769);
and U16666 (N_16666,N_12476,N_11285);
nand U16667 (N_16667,N_11295,N_11356);
nor U16668 (N_16668,N_14507,N_11359);
xnor U16669 (N_16669,N_13526,N_12260);
nor U16670 (N_16670,N_10483,N_14639);
nor U16671 (N_16671,N_10226,N_13778);
or U16672 (N_16672,N_12808,N_12720);
or U16673 (N_16673,N_11703,N_10455);
nand U16674 (N_16674,N_12049,N_14974);
nor U16675 (N_16675,N_12241,N_12867);
xor U16676 (N_16676,N_13186,N_14982);
nand U16677 (N_16677,N_12079,N_11964);
or U16678 (N_16678,N_11222,N_14910);
nand U16679 (N_16679,N_11933,N_11574);
nor U16680 (N_16680,N_13429,N_10846);
nor U16681 (N_16681,N_11921,N_14269);
nor U16682 (N_16682,N_13435,N_11890);
and U16683 (N_16683,N_11965,N_10772);
or U16684 (N_16684,N_13960,N_11875);
xnor U16685 (N_16685,N_10055,N_12744);
nor U16686 (N_16686,N_12711,N_13533);
and U16687 (N_16687,N_10848,N_10573);
or U16688 (N_16688,N_12648,N_14895);
and U16689 (N_16689,N_14428,N_12565);
xnor U16690 (N_16690,N_10649,N_11737);
and U16691 (N_16691,N_11525,N_11123);
nand U16692 (N_16692,N_12403,N_14326);
or U16693 (N_16693,N_14490,N_10948);
xor U16694 (N_16694,N_14107,N_14360);
or U16695 (N_16695,N_14442,N_14364);
xnor U16696 (N_16696,N_12774,N_11651);
xnor U16697 (N_16697,N_10785,N_13805);
nor U16698 (N_16698,N_13996,N_10091);
or U16699 (N_16699,N_10719,N_14867);
or U16700 (N_16700,N_10057,N_12581);
and U16701 (N_16701,N_12968,N_14883);
or U16702 (N_16702,N_14256,N_14416);
xor U16703 (N_16703,N_11690,N_13677);
nor U16704 (N_16704,N_13894,N_14847);
nor U16705 (N_16705,N_14079,N_13293);
and U16706 (N_16706,N_13787,N_14809);
xnor U16707 (N_16707,N_10872,N_13637);
or U16708 (N_16708,N_14650,N_14247);
xor U16709 (N_16709,N_10656,N_14043);
and U16710 (N_16710,N_11073,N_13112);
xnor U16711 (N_16711,N_13373,N_11617);
and U16712 (N_16712,N_11940,N_12930);
xnor U16713 (N_16713,N_12801,N_13963);
xnor U16714 (N_16714,N_13319,N_12863);
nand U16715 (N_16715,N_10408,N_10004);
nor U16716 (N_16716,N_12024,N_10822);
xnor U16717 (N_16717,N_12290,N_13958);
or U16718 (N_16718,N_14732,N_13562);
or U16719 (N_16719,N_11620,N_11990);
or U16720 (N_16720,N_13912,N_13966);
nor U16721 (N_16721,N_13596,N_10227);
and U16722 (N_16722,N_12962,N_14276);
nor U16723 (N_16723,N_14829,N_10144);
nand U16724 (N_16724,N_14989,N_11967);
or U16725 (N_16725,N_14954,N_13126);
or U16726 (N_16726,N_12948,N_13817);
xor U16727 (N_16727,N_10244,N_10823);
nand U16728 (N_16728,N_11043,N_13954);
and U16729 (N_16729,N_12055,N_10002);
nand U16730 (N_16730,N_14838,N_12862);
nand U16731 (N_16731,N_14517,N_14696);
nor U16732 (N_16732,N_12524,N_14128);
xnor U16733 (N_16733,N_10832,N_10054);
xor U16734 (N_16734,N_13317,N_10583);
nor U16735 (N_16735,N_13862,N_11810);
and U16736 (N_16736,N_11028,N_13681);
nor U16737 (N_16737,N_13666,N_12804);
nor U16738 (N_16738,N_10767,N_10605);
xnor U16739 (N_16739,N_13152,N_10618);
xnor U16740 (N_16740,N_14651,N_12083);
and U16741 (N_16741,N_12346,N_10468);
and U16742 (N_16742,N_11389,N_14702);
xor U16743 (N_16743,N_12141,N_12628);
nand U16744 (N_16744,N_11017,N_12493);
xor U16745 (N_16745,N_10676,N_11101);
xnor U16746 (N_16746,N_14969,N_11916);
nand U16747 (N_16747,N_12776,N_13130);
xor U16748 (N_16748,N_10251,N_14924);
nand U16749 (N_16749,N_13957,N_12574);
and U16750 (N_16750,N_14236,N_14919);
nor U16751 (N_16751,N_13170,N_14063);
nor U16752 (N_16752,N_10729,N_12182);
nand U16753 (N_16753,N_12430,N_12505);
xnor U16754 (N_16754,N_10813,N_13656);
nand U16755 (N_16755,N_13525,N_12371);
nand U16756 (N_16756,N_11549,N_12717);
and U16757 (N_16757,N_11745,N_14145);
and U16758 (N_16758,N_12790,N_10543);
nor U16759 (N_16759,N_13312,N_11455);
xnor U16760 (N_16760,N_11384,N_13917);
and U16761 (N_16761,N_10240,N_14474);
and U16762 (N_16762,N_12771,N_14806);
nand U16763 (N_16763,N_10273,N_13828);
nor U16764 (N_16764,N_11517,N_13889);
and U16765 (N_16765,N_12377,N_14701);
nor U16766 (N_16766,N_10167,N_14039);
nand U16767 (N_16767,N_10886,N_10418);
nand U16768 (N_16768,N_10414,N_12639);
nor U16769 (N_16769,N_14008,N_14125);
and U16770 (N_16770,N_14817,N_12204);
or U16771 (N_16771,N_12755,N_12463);
nor U16772 (N_16772,N_12088,N_10427);
nor U16773 (N_16773,N_14670,N_10453);
xnor U16774 (N_16774,N_11659,N_13179);
nand U16775 (N_16775,N_13494,N_11435);
nand U16776 (N_16776,N_12625,N_10138);
or U16777 (N_16777,N_12208,N_11985);
nand U16778 (N_16778,N_14362,N_10476);
nor U16779 (N_16779,N_14121,N_10644);
and U16780 (N_16780,N_10299,N_12974);
and U16781 (N_16781,N_12642,N_12847);
nand U16782 (N_16782,N_12955,N_14268);
nand U16783 (N_16783,N_12945,N_12186);
nor U16784 (N_16784,N_11412,N_10839);
xor U16785 (N_16785,N_14193,N_10190);
nor U16786 (N_16786,N_14226,N_12920);
nor U16787 (N_16787,N_11233,N_11369);
or U16788 (N_16788,N_13222,N_11158);
xor U16789 (N_16789,N_11091,N_11579);
nand U16790 (N_16790,N_10130,N_12678);
nand U16791 (N_16791,N_13477,N_13948);
or U16792 (N_16792,N_14687,N_11554);
xor U16793 (N_16793,N_14531,N_14424);
nor U16794 (N_16794,N_12385,N_13420);
or U16795 (N_16795,N_13316,N_10224);
nand U16796 (N_16796,N_10389,N_11114);
nor U16797 (N_16797,N_13878,N_14652);
and U16798 (N_16798,N_11373,N_11395);
and U16799 (N_16799,N_12009,N_12520);
xor U16800 (N_16800,N_10990,N_14562);
or U16801 (N_16801,N_12508,N_13043);
nand U16802 (N_16802,N_13927,N_12118);
and U16803 (N_16803,N_10718,N_14785);
nor U16804 (N_16804,N_13256,N_14956);
nand U16805 (N_16805,N_10671,N_14976);
nor U16806 (N_16806,N_14936,N_11276);
or U16807 (N_16807,N_14948,N_14230);
nor U16808 (N_16808,N_10097,N_13330);
or U16809 (N_16809,N_11122,N_11671);
and U16810 (N_16810,N_14228,N_11830);
xor U16811 (N_16811,N_14299,N_13448);
nor U16812 (N_16812,N_11679,N_10755);
nor U16813 (N_16813,N_11769,N_12066);
xor U16814 (N_16814,N_14620,N_11102);
nor U16815 (N_16815,N_13406,N_14197);
xor U16816 (N_16816,N_14373,N_12390);
and U16817 (N_16817,N_13692,N_11218);
xnor U16818 (N_16818,N_13143,N_11646);
nor U16819 (N_16819,N_12966,N_11540);
and U16820 (N_16820,N_10805,N_11105);
nand U16821 (N_16821,N_12651,N_14963);
nor U16822 (N_16822,N_13113,N_12825);
xnor U16823 (N_16823,N_13072,N_11361);
nor U16824 (N_16824,N_10207,N_10239);
or U16825 (N_16825,N_10320,N_10210);
and U16826 (N_16826,N_14127,N_10186);
nor U16827 (N_16827,N_12177,N_12171);
or U16828 (N_16828,N_12416,N_11536);
nor U16829 (N_16829,N_10209,N_11607);
xnor U16830 (N_16830,N_11313,N_12254);
xnor U16831 (N_16831,N_12573,N_12689);
nor U16832 (N_16832,N_11310,N_12672);
nand U16833 (N_16833,N_11092,N_11047);
nor U16834 (N_16834,N_13669,N_12303);
nor U16835 (N_16835,N_12005,N_14815);
or U16836 (N_16836,N_13246,N_12747);
and U16837 (N_16837,N_11450,N_10082);
and U16838 (N_16838,N_10733,N_12870);
nor U16839 (N_16839,N_12149,N_14610);
xnor U16840 (N_16840,N_10866,N_12949);
and U16841 (N_16841,N_14607,N_12589);
xor U16842 (N_16842,N_14964,N_10850);
xnor U16843 (N_16843,N_12102,N_10090);
nand U16844 (N_16844,N_12473,N_12537);
and U16845 (N_16845,N_13213,N_14050);
xor U16846 (N_16846,N_12715,N_12912);
and U16847 (N_16847,N_10440,N_12443);
or U16848 (N_16848,N_11368,N_13399);
and U16849 (N_16849,N_12784,N_12855);
or U16850 (N_16850,N_12743,N_13350);
or U16851 (N_16851,N_11758,N_12095);
nand U16852 (N_16852,N_11571,N_11237);
and U16853 (N_16853,N_10840,N_11445);
nand U16854 (N_16854,N_11289,N_10262);
nand U16855 (N_16855,N_12553,N_13624);
xor U16856 (N_16856,N_13955,N_14419);
nor U16857 (N_16857,N_14616,N_14565);
nor U16858 (N_16858,N_13289,N_13920);
and U16859 (N_16859,N_10855,N_13410);
and U16860 (N_16860,N_13219,N_13569);
nor U16861 (N_16861,N_12180,N_13929);
or U16862 (N_16862,N_13073,N_12646);
nor U16863 (N_16863,N_11269,N_10221);
or U16864 (N_16864,N_12480,N_13782);
xnor U16865 (N_16865,N_11453,N_13846);
and U16866 (N_16866,N_12519,N_10973);
nor U16867 (N_16867,N_14259,N_13883);
nand U16868 (N_16868,N_12997,N_11531);
or U16869 (N_16869,N_13057,N_12229);
or U16870 (N_16870,N_11686,N_14242);
nand U16871 (N_16871,N_13308,N_10930);
nand U16872 (N_16872,N_14086,N_11995);
or U16873 (N_16873,N_12326,N_13412);
nor U16874 (N_16874,N_11959,N_13280);
xnor U16875 (N_16875,N_11835,N_10348);
nor U16876 (N_16876,N_12194,N_14270);
xnor U16877 (N_16877,N_11268,N_14638);
nor U16878 (N_16878,N_13471,N_14609);
nor U16879 (N_16879,N_12880,N_13003);
or U16880 (N_16880,N_14160,N_10193);
xor U16881 (N_16881,N_13465,N_11296);
nand U16882 (N_16882,N_10876,N_10472);
nand U16883 (N_16883,N_11781,N_11362);
nand U16884 (N_16884,N_10706,N_11978);
nand U16885 (N_16885,N_11895,N_10901);
xnor U16886 (N_16886,N_11244,N_14191);
and U16887 (N_16887,N_12097,N_10510);
nor U16888 (N_16888,N_13520,N_10863);
or U16889 (N_16889,N_10777,N_12472);
and U16890 (N_16890,N_12313,N_12500);
xnor U16891 (N_16891,N_11030,N_11415);
xor U16892 (N_16892,N_14535,N_13724);
nand U16893 (N_16893,N_12656,N_10430);
nor U16894 (N_16894,N_14926,N_13688);
nand U16895 (N_16895,N_12250,N_11408);
or U16896 (N_16896,N_13502,N_14281);
nand U16897 (N_16897,N_14329,N_12304);
nand U16898 (N_16898,N_14246,N_12166);
nor U16899 (N_16899,N_12011,N_10558);
xnor U16900 (N_16900,N_10825,N_10179);
nor U16901 (N_16901,N_11211,N_10585);
and U16902 (N_16902,N_10119,N_12971);
and U16903 (N_16903,N_11272,N_14453);
nand U16904 (N_16904,N_11812,N_11338);
xor U16905 (N_16905,N_14635,N_10960);
and U16906 (N_16906,N_12523,N_10845);
and U16907 (N_16907,N_14022,N_11663);
nor U16908 (N_16908,N_11528,N_13573);
xor U16909 (N_16909,N_12342,N_13615);
and U16910 (N_16910,N_13660,N_13645);
xor U16911 (N_16911,N_14626,N_10318);
nor U16912 (N_16912,N_14011,N_14034);
nor U16913 (N_16913,N_12583,N_13455);
nor U16914 (N_16914,N_14209,N_13648);
nor U16915 (N_16915,N_11491,N_10730);
or U16916 (N_16916,N_10063,N_13326);
xnor U16917 (N_16917,N_11042,N_13937);
nor U16918 (N_16918,N_11134,N_12479);
nand U16919 (N_16919,N_13454,N_10406);
or U16920 (N_16920,N_13034,N_12593);
nor U16921 (N_16921,N_12386,N_13499);
and U16922 (N_16922,N_13510,N_12534);
nand U16923 (N_16923,N_10181,N_14272);
nor U16924 (N_16924,N_13370,N_11254);
nand U16925 (N_16925,N_11068,N_12311);
or U16926 (N_16926,N_10098,N_10201);
or U16927 (N_16927,N_11136,N_14797);
and U16928 (N_16928,N_12676,N_12729);
or U16929 (N_16929,N_13094,N_10473);
nor U16930 (N_16930,N_13701,N_14548);
and U16931 (N_16931,N_13366,N_11152);
and U16932 (N_16932,N_10512,N_12969);
xor U16933 (N_16933,N_10860,N_14338);
nand U16934 (N_16934,N_13318,N_14849);
nor U16935 (N_16935,N_13401,N_12477);
nor U16936 (N_16936,N_10521,N_13867);
or U16937 (N_16937,N_12201,N_10129);
and U16938 (N_16938,N_13593,N_14823);
or U16939 (N_16939,N_10527,N_10843);
nor U16940 (N_16940,N_11836,N_13320);
or U16941 (N_16941,N_11948,N_13055);
xnor U16942 (N_16942,N_14645,N_14682);
xnor U16943 (N_16943,N_10000,N_10337);
xor U16944 (N_16944,N_13601,N_14097);
nand U16945 (N_16945,N_12596,N_11459);
or U16946 (N_16946,N_13728,N_14418);
or U16947 (N_16947,N_10078,N_14407);
nor U16948 (N_16948,N_10780,N_10988);
xor U16949 (N_16949,N_14717,N_11008);
nor U16950 (N_16950,N_13394,N_10931);
and U16951 (N_16951,N_10155,N_14049);
nor U16952 (N_16952,N_13071,N_11131);
or U16953 (N_16953,N_12615,N_12114);
nor U16954 (N_16954,N_14017,N_10817);
xor U16955 (N_16955,N_11504,N_12040);
xnor U16956 (N_16956,N_14680,N_13283);
xor U16957 (N_16957,N_14081,N_10357);
and U16958 (N_16958,N_13466,N_12289);
nand U16959 (N_16959,N_11851,N_14435);
nand U16960 (N_16960,N_12432,N_14757);
and U16961 (N_16961,N_11779,N_12873);
and U16962 (N_16962,N_14841,N_10548);
and U16963 (N_16963,N_12404,N_14791);
xnor U16964 (N_16964,N_12512,N_12538);
nor U16965 (N_16965,N_14415,N_11394);
nand U16966 (N_16966,N_12360,N_12809);
and U16967 (N_16967,N_11195,N_14643);
xor U16968 (N_16968,N_12731,N_13989);
and U16969 (N_16969,N_14131,N_14467);
or U16970 (N_16970,N_10486,N_11351);
nand U16971 (N_16971,N_12288,N_13299);
xnor U16972 (N_16972,N_14280,N_10417);
nor U16973 (N_16973,N_12281,N_12388);
nand U16974 (N_16974,N_10060,N_11034);
nand U16975 (N_16975,N_12230,N_11480);
or U16976 (N_16976,N_11055,N_14136);
nor U16977 (N_16977,N_14402,N_13291);
and U16978 (N_16978,N_11200,N_14031);
nand U16979 (N_16979,N_13576,N_12325);
nand U16980 (N_16980,N_13208,N_14991);
or U16981 (N_16981,N_13505,N_13909);
nor U16982 (N_16982,N_14007,N_12402);
nor U16983 (N_16983,N_11204,N_14818);
or U16984 (N_16984,N_12268,N_14015);
nor U16985 (N_16985,N_11723,N_14958);
nor U16986 (N_16986,N_10237,N_10570);
xor U16987 (N_16987,N_10154,N_14250);
nand U16988 (N_16988,N_10694,N_13047);
and U16989 (N_16989,N_13663,N_14566);
nand U16990 (N_16990,N_13544,N_11768);
or U16991 (N_16991,N_12276,N_14180);
nor U16992 (N_16992,N_13824,N_12788);
nand U16993 (N_16993,N_13933,N_11012);
nand U16994 (N_16994,N_11760,N_11145);
xor U16995 (N_16995,N_10079,N_13675);
or U16996 (N_16996,N_13415,N_10449);
nor U16997 (N_16997,N_11069,N_11287);
nor U16998 (N_16998,N_14549,N_12335);
xor U16999 (N_16999,N_10234,N_13742);
or U17000 (N_17000,N_14877,N_12158);
and U17001 (N_17001,N_13731,N_14770);
nor U17002 (N_17002,N_10677,N_10882);
nor U17003 (N_17003,N_10458,N_10436);
or U17004 (N_17004,N_14431,N_13930);
or U17005 (N_17005,N_11575,N_12108);
nor U17006 (N_17006,N_11253,N_11004);
and U17007 (N_17007,N_14759,N_12922);
nor U17008 (N_17008,N_14563,N_12637);
nand U17009 (N_17009,N_13037,N_14930);
nand U17010 (N_17010,N_10233,N_11772);
or U17011 (N_17011,N_12471,N_10599);
nor U17012 (N_17012,N_11257,N_11797);
xnor U17013 (N_17013,N_12008,N_11203);
xnor U17014 (N_17014,N_14243,N_13168);
nor U17015 (N_17015,N_10883,N_13879);
nor U17016 (N_17016,N_12541,N_10194);
nand U17017 (N_17017,N_13600,N_10250);
xnor U17018 (N_17018,N_14500,N_14076);
xnor U17019 (N_17019,N_14438,N_14320);
nand U17020 (N_17020,N_12023,N_11970);
nor U17021 (N_17021,N_12383,N_12564);
nor U17022 (N_17022,N_10645,N_12262);
nand U17023 (N_17023,N_12822,N_14122);
nand U17024 (N_17024,N_10617,N_11506);
nor U17025 (N_17025,N_14525,N_10058);
or U17026 (N_17026,N_14925,N_13765);
or U17027 (N_17027,N_11084,N_10236);
xnor U17028 (N_17028,N_13060,N_12685);
nand U17029 (N_17029,N_11472,N_13387);
nand U17030 (N_17030,N_12334,N_14567);
xor U17031 (N_17031,N_13041,N_11299);
xor U17032 (N_17032,N_13640,N_11912);
and U17033 (N_17033,N_13735,N_11402);
xor U17034 (N_17034,N_12156,N_13858);
and U17035 (N_17035,N_12073,N_13876);
nor U17036 (N_17036,N_12047,N_11345);
nand U17037 (N_17037,N_13206,N_13187);
nor U17038 (N_17038,N_14202,N_12760);
or U17039 (N_17039,N_11274,N_11683);
and U17040 (N_17040,N_14387,N_10952);
nor U17041 (N_17041,N_14220,N_10885);
and U17042 (N_17042,N_14943,N_14756);
nor U17043 (N_17043,N_13141,N_14977);
and U17044 (N_17044,N_10304,N_11908);
xor U17045 (N_17045,N_12934,N_10925);
and U17046 (N_17046,N_10447,N_14834);
and U17047 (N_17047,N_13404,N_14824);
and U17048 (N_17048,N_13975,N_14426);
and U17049 (N_17049,N_13056,N_10809);
or U17050 (N_17050,N_14038,N_11259);
and U17051 (N_17051,N_14096,N_14795);
nor U17052 (N_17052,N_11386,N_11856);
and U17053 (N_17053,N_12218,N_14686);
or U17054 (N_17054,N_10529,N_10391);
xor U17055 (N_17055,N_11748,N_11391);
nor U17056 (N_17056,N_14999,N_14875);
and U17057 (N_17057,N_10255,N_14997);
and U17058 (N_17058,N_13800,N_13882);
xnor U17059 (N_17059,N_12347,N_12107);
xor U17060 (N_17060,N_14961,N_12838);
nand U17061 (N_17061,N_13334,N_13375);
nor U17062 (N_17062,N_13178,N_10852);
or U17063 (N_17063,N_13290,N_14319);
xnor U17064 (N_17064,N_11221,N_14159);
nand U17065 (N_17065,N_11643,N_11917);
or U17066 (N_17066,N_11552,N_12654);
or U17067 (N_17067,N_11177,N_10359);
and U17068 (N_17068,N_12223,N_11079);
xnor U17069 (N_17069,N_13849,N_12634);
xor U17070 (N_17070,N_13150,N_13205);
nand U17071 (N_17071,N_12272,N_14060);
nor U17072 (N_17072,N_12752,N_13540);
nand U17073 (N_17073,N_11919,N_14380);
nor U17074 (N_17074,N_14529,N_12270);
and U17075 (N_17075,N_13124,N_10302);
xnor U17076 (N_17076,N_13855,N_12662);
nor U17077 (N_17077,N_11382,N_14304);
and U17078 (N_17078,N_11873,N_12567);
nand U17079 (N_17079,N_11811,N_11342);
xor U17080 (N_17080,N_14547,N_14899);
xor U17081 (N_17081,N_11119,N_11314);
nand U17082 (N_17082,N_12205,N_14201);
xor U17083 (N_17083,N_11000,N_12757);
and U17084 (N_17084,N_13048,N_13436);
nor U17085 (N_17085,N_11067,N_14856);
and U17086 (N_17086,N_10457,N_12031);
nand U17087 (N_17087,N_10347,N_14044);
nand U17088 (N_17088,N_12978,N_13697);
and U17089 (N_17089,N_10523,N_14252);
and U17090 (N_17090,N_14764,N_14837);
xnor U17091 (N_17091,N_13722,N_11236);
nor U17092 (N_17092,N_13877,N_11036);
or U17093 (N_17093,N_13822,N_13633);
or U17094 (N_17094,N_11247,N_13547);
nand U17095 (N_17095,N_12319,N_12636);
or U17096 (N_17096,N_12411,N_14522);
xnor U17097 (N_17097,N_11641,N_12169);
nor U17098 (N_17098,N_10434,N_14504);
nor U17099 (N_17099,N_14788,N_12803);
xnor U17100 (N_17100,N_14472,N_14492);
or U17101 (N_17101,N_14417,N_14458);
nand U17102 (N_17102,N_14518,N_10705);
xor U17103 (N_17103,N_10183,N_13915);
xor U17104 (N_17104,N_10939,N_14056);
and U17105 (N_17105,N_14434,N_11501);
nand U17106 (N_17106,N_10249,N_13365);
nand U17107 (N_17107,N_13463,N_14750);
and U17108 (N_17108,N_11197,N_13940);
xnor U17109 (N_17109,N_13588,N_11901);
or U17110 (N_17110,N_13581,N_13264);
nor U17111 (N_17111,N_10289,N_10500);
nor U17112 (N_17112,N_13923,N_13381);
xnor U17113 (N_17113,N_10110,N_12584);
xor U17114 (N_17114,N_13725,N_13931);
xnor U17115 (N_17115,N_13024,N_13934);
nor U17116 (N_17116,N_13374,N_14772);
or U17117 (N_17117,N_14619,N_10713);
nor U17118 (N_17118,N_10397,N_10324);
nand U17119 (N_17119,N_14988,N_10032);
and U17120 (N_17120,N_11496,N_12691);
xor U17121 (N_17121,N_13708,N_11834);
and U17122 (N_17122,N_11858,N_12010);
nor U17123 (N_17123,N_11653,N_10628);
xor U17124 (N_17124,N_11477,N_13424);
xor U17125 (N_17125,N_14206,N_13460);
xnor U17126 (N_17126,N_11175,N_11601);
nand U17127 (N_17127,N_10459,N_10747);
xnor U17128 (N_17128,N_10260,N_11343);
or U17129 (N_17129,N_13710,N_14174);
nor U17130 (N_17130,N_13301,N_11270);
xnor U17131 (N_17131,N_13468,N_10220);
xnor U17132 (N_17132,N_12543,N_11974);
nor U17133 (N_17133,N_13628,N_10879);
and U17134 (N_17134,N_13392,N_13981);
or U17135 (N_17135,N_13031,N_10926);
or U17136 (N_17136,N_11110,N_12029);
xor U17137 (N_17137,N_13382,N_14295);
or U17138 (N_17138,N_12358,N_12195);
or U17139 (N_17139,N_13165,N_12207);
xor U17140 (N_17140,N_11172,N_10248);
nand U17141 (N_17141,N_10093,N_12380);
and U17142 (N_17142,N_14851,N_11550);
and U17143 (N_17143,N_13044,N_13740);
or U17144 (N_17144,N_14337,N_11431);
xnor U17145 (N_17145,N_11440,N_10700);
nand U17146 (N_17146,N_10658,N_11657);
nand U17147 (N_17147,N_11692,N_13335);
and U17148 (N_17148,N_12713,N_14648);
or U17149 (N_17149,N_13904,N_12485);
nand U17150 (N_17150,N_10898,N_12579);
or U17151 (N_17151,N_14695,N_14751);
and U17152 (N_17152,N_10416,N_10051);
nand U17153 (N_17153,N_11971,N_14941);
nand U17154 (N_17154,N_13434,N_11443);
xor U17155 (N_17155,N_10216,N_14835);
or U17156 (N_17156,N_14368,N_12292);
nand U17157 (N_17157,N_14318,N_12813);
nor U17158 (N_17158,N_13364,N_14052);
and U17159 (N_17159,N_14233,N_13700);
xor U17160 (N_17160,N_10927,N_14903);
nor U17161 (N_17161,N_10290,N_11631);
xnor U17162 (N_17162,N_12399,N_14117);
and U17163 (N_17163,N_12510,N_14805);
nand U17164 (N_17164,N_10940,N_10300);
xor U17165 (N_17165,N_13193,N_12225);
and U17166 (N_17166,N_11790,N_13021);
xor U17167 (N_17167,N_13327,N_13447);
nand U17168 (N_17168,N_11866,N_10993);
and U17169 (N_17169,N_13054,N_14323);
or U17170 (N_17170,N_14484,N_10219);
and U17171 (N_17171,N_13621,N_12340);
nor U17172 (N_17172,N_14564,N_14542);
nor U17173 (N_17173,N_13212,N_13076);
and U17174 (N_17174,N_13481,N_13083);
xor U17175 (N_17175,N_11053,N_13524);
xor U17176 (N_17176,N_13830,N_10212);
xnor U17177 (N_17177,N_14990,N_14905);
xor U17178 (N_17178,N_14843,N_14087);
or U17179 (N_17179,N_11701,N_10771);
or U17180 (N_17180,N_14537,N_13267);
nand U17181 (N_17181,N_13837,N_13232);
and U17182 (N_17182,N_11117,N_11820);
nor U17183 (N_17183,N_12277,N_11952);
or U17184 (N_17184,N_13563,N_12533);
and U17185 (N_17185,N_12378,N_14219);
nor U17186 (N_17186,N_13411,N_13380);
or U17187 (N_17187,N_13711,N_10812);
xnor U17188 (N_17188,N_13227,N_14594);
nand U17189 (N_17189,N_13458,N_14386);
nand U17190 (N_17190,N_11602,N_10790);
nand U17191 (N_17191,N_10118,N_10134);
nor U17192 (N_17192,N_10482,N_10270);
nor U17193 (N_17193,N_14221,N_14321);
nand U17194 (N_17194,N_13221,N_10828);
nand U17195 (N_17195,N_13109,N_14171);
and U17196 (N_17196,N_14519,N_10907);
xor U17197 (N_17197,N_11056,N_12099);
or U17198 (N_17198,N_14479,N_14432);
xor U17199 (N_17199,N_12408,N_13298);
xnor U17200 (N_17200,N_13754,N_14082);
xnor U17201 (N_17201,N_11255,N_13098);
nor U17202 (N_17202,N_10556,N_11467);
nand U17203 (N_17203,N_13959,N_12252);
and U17204 (N_17204,N_14984,N_10501);
or U17205 (N_17205,N_11228,N_10966);
nand U17206 (N_17206,N_12716,N_13650);
and U17207 (N_17207,N_13011,N_13164);
xor U17208 (N_17208,N_13204,N_12221);
xor U17209 (N_17209,N_13296,N_13798);
or U17210 (N_17210,N_14150,N_10657);
and U17211 (N_17211,N_13046,N_11166);
or U17212 (N_17212,N_10761,N_14798);
nor U17213 (N_17213,N_10376,N_14572);
nand U17214 (N_17214,N_11640,N_14704);
and U17215 (N_17215,N_14264,N_14216);
and U17216 (N_17216,N_10802,N_14496);
or U17217 (N_17217,N_13125,N_14302);
and U17218 (N_17218,N_12176,N_13184);
xor U17219 (N_17219,N_14388,N_12454);
nor U17220 (N_17220,N_12353,N_11893);
or U17221 (N_17221,N_13965,N_12722);
xnor U17222 (N_17222,N_10071,N_10310);
or U17223 (N_17223,N_12222,N_12350);
xor U17224 (N_17224,N_11882,N_10339);
xor U17225 (N_17225,N_11106,N_12045);
nor U17226 (N_17226,N_10791,N_12264);
and U17227 (N_17227,N_14475,N_13715);
and U17228 (N_17228,N_13806,N_10716);
nor U17229 (N_17229,N_14396,N_12307);
nor U17230 (N_17230,N_12837,N_14002);
and U17231 (N_17231,N_12376,N_13872);
or U17232 (N_17232,N_12630,N_11869);
xor U17233 (N_17233,N_10530,N_14985);
nor U17234 (N_17234,N_12484,N_10332);
nor U17235 (N_17235,N_12062,N_11817);
or U17236 (N_17236,N_12728,N_13371);
and U17237 (N_17237,N_13761,N_14456);
xnor U17238 (N_17238,N_12887,N_10050);
xnor U17239 (N_17239,N_10943,N_12052);
nand U17240 (N_17240,N_12014,N_14676);
xor U17241 (N_17241,N_12364,N_12253);
or U17242 (N_17242,N_11183,N_10352);
xnor U17243 (N_17243,N_12693,N_14864);
nand U17244 (N_17244,N_13726,N_14036);
xor U17245 (N_17245,N_10253,N_10362);
nand U17246 (N_17246,N_13103,N_14909);
xor U17247 (N_17247,N_10488,N_11350);
or U17248 (N_17248,N_11303,N_11414);
xnor U17249 (N_17249,N_12794,N_10619);
xnor U17250 (N_17250,N_10967,N_13786);
or U17251 (N_17251,N_12457,N_12738);
nor U17252 (N_17252,N_10287,N_12144);
xor U17253 (N_17253,N_12469,N_11662);
and U17254 (N_17254,N_13426,N_10275);
nand U17255 (N_17255,N_12852,N_12251);
nor U17256 (N_17256,N_13542,N_10751);
nand U17257 (N_17257,N_13145,N_14385);
and U17258 (N_17258,N_10999,N_13962);
and U17259 (N_17259,N_10145,N_13116);
xnor U17260 (N_17260,N_14203,N_14827);
and U17261 (N_17261,N_11404,N_11436);
nand U17262 (N_17262,N_12617,N_10267);
xor U17263 (N_17263,N_13519,N_11448);
or U17264 (N_17264,N_12623,N_13425);
nor U17265 (N_17265,N_10115,N_10636);
xor U17266 (N_17266,N_14184,N_12875);
nor U17267 (N_17267,N_14051,N_12918);
xor U17268 (N_17268,N_14804,N_12613);
or U17269 (N_17269,N_11839,N_10184);
and U17270 (N_17270,N_11484,N_10859);
and U17271 (N_17271,N_11180,N_11845);
xor U17272 (N_17272,N_14513,N_11432);
nor U17273 (N_17273,N_11418,N_14752);
and U17274 (N_17274,N_14965,N_12810);
and U17275 (N_17275,N_14729,N_11741);
nand U17276 (N_17276,N_13532,N_14353);
nor U17277 (N_17277,N_11712,N_12423);
or U17278 (N_17278,N_14314,N_11031);
nor U17279 (N_17279,N_13093,N_13583);
and U17280 (N_17280,N_14728,N_13229);
nor U17281 (N_17281,N_12465,N_11320);
nor U17282 (N_17282,N_11099,N_10136);
nand U17283 (N_17283,N_14098,N_14311);
xnor U17284 (N_17284,N_14333,N_10096);
nor U17285 (N_17285,N_12721,N_10786);
nor U17286 (N_17286,N_12914,N_12372);
and U17287 (N_17287,N_12138,N_10704);
or U17288 (N_17288,N_12931,N_12090);
xnor U17289 (N_17289,N_12298,N_14720);
nand U17290 (N_17290,N_11902,N_10982);
nand U17291 (N_17291,N_12041,N_14946);
and U17292 (N_17292,N_11844,N_12450);
or U17293 (N_17293,N_13664,N_13014);
xor U17294 (N_17294,N_14972,N_11627);
and U17295 (N_17295,N_12061,N_14995);
nand U17296 (N_17296,N_14102,N_11385);
or U17297 (N_17297,N_11867,N_12320);
xnor U17298 (N_17298,N_10688,N_14868);
xor U17299 (N_17299,N_14437,N_14957);
xor U17300 (N_17300,N_11116,N_12539);
nor U17301 (N_17301,N_13723,N_11957);
and U17302 (N_17302,N_12027,N_12080);
xor U17303 (N_17303,N_11058,N_11876);
or U17304 (N_17304,N_12811,N_11777);
nor U17305 (N_17305,N_12714,N_10053);
xnor U17306 (N_17306,N_11963,N_11417);
nand U17307 (N_17307,N_14892,N_12050);
xnor U17308 (N_17308,N_13106,N_10909);
and U17309 (N_17309,N_10368,N_14282);
nand U17310 (N_17310,N_14694,N_11438);
xor U17311 (N_17311,N_14574,N_14754);
nand U17312 (N_17312,N_14100,N_10969);
nand U17313 (N_17313,N_12655,N_10601);
nand U17314 (N_17314,N_10989,N_11915);
and U17315 (N_17315,N_12675,N_11821);
nor U17316 (N_17316,N_12640,N_10378);
xor U17317 (N_17317,N_12585,N_13391);
nor U17318 (N_17318,N_14700,N_10881);
nand U17319 (N_17319,N_10945,N_12249);
or U17320 (N_17320,N_11141,N_11791);
and U17321 (N_17321,N_13134,N_13988);
nor U17322 (N_17322,N_11805,N_13605);
nand U17323 (N_17323,N_12131,N_12709);
xnor U17324 (N_17324,N_14796,N_10774);
nand U17325 (N_17325,N_11075,N_14089);
and U17326 (N_17326,N_14296,N_11217);
nor U17327 (N_17327,N_11013,N_11312);
or U17328 (N_17328,N_10301,N_10470);
nand U17329 (N_17329,N_11346,N_10164);
xor U17330 (N_17330,N_10462,N_11616);
nand U17331 (N_17331,N_10561,N_12185);
and U17332 (N_17332,N_14690,N_14688);
or U17333 (N_17333,N_13914,N_12419);
nand U17334 (N_17334,N_12705,N_12458);
xnor U17335 (N_17335,N_10297,N_12936);
or U17336 (N_17336,N_13766,N_10528);
and U17337 (N_17337,N_10029,N_10401);
and U17338 (N_17338,N_12611,N_12766);
xnor U17339 (N_17339,N_11962,N_11238);
and U17340 (N_17340,N_11956,N_12777);
nand U17341 (N_17341,N_11585,N_13214);
and U17342 (N_17342,N_11444,N_14794);
xor U17343 (N_17343,N_11515,N_11799);
or U17344 (N_17344,N_13314,N_10695);
xor U17345 (N_17345,N_12518,N_10574);
xor U17346 (N_17346,N_12105,N_13008);
nor U17347 (N_17347,N_10373,N_11649);
nand U17348 (N_17348,N_13756,N_12091);
xnor U17349 (N_17349,N_13306,N_12209);
nor U17350 (N_17350,N_10007,N_11567);
xnor U17351 (N_17351,N_11618,N_12635);
or U17352 (N_17352,N_14614,N_12963);
nand U17353 (N_17353,N_11214,N_14462);
and U17354 (N_17354,N_13461,N_12602);
xnor U17355 (N_17355,N_10274,N_13513);
or U17356 (N_17356,N_12854,N_13762);
xor U17357 (N_17357,N_10030,N_14062);
xnor U17358 (N_17358,N_12710,N_13752);
or U17359 (N_17359,N_14588,N_11051);
or U17360 (N_17360,N_13683,N_13097);
or U17361 (N_17361,N_10170,N_10981);
or U17362 (N_17362,N_14059,N_10189);
nor U17363 (N_17363,N_10506,N_10498);
nand U17364 (N_17364,N_10536,N_13826);
and U17365 (N_17365,N_12406,N_11589);
nand U17366 (N_17366,N_14913,N_12641);
or U17367 (N_17367,N_12212,N_10980);
and U17368 (N_17368,N_11898,N_14934);
nand U17369 (N_17369,N_11794,N_14778);
and U17370 (N_17370,N_11966,N_12859);
and U17371 (N_17371,N_13445,N_14409);
xnor U17372 (N_17372,N_11063,N_12327);
and U17373 (N_17373,N_10798,N_10589);
nor U17374 (N_17374,N_11317,N_13080);
or U17375 (N_17375,N_10238,N_11650);
or U17376 (N_17376,N_11288,N_11392);
or U17377 (N_17377,N_14618,N_12389);
nand U17378 (N_17378,N_12695,N_12323);
xor U17379 (N_17379,N_14568,N_13070);
or U17380 (N_17380,N_12791,N_10222);
or U17381 (N_17381,N_12233,N_10916);
nor U17382 (N_17382,N_12604,N_11349);
or U17383 (N_17383,N_11648,N_11600);
nor U17384 (N_17384,N_13942,N_13980);
and U17385 (N_17385,N_12098,N_11410);
xnor U17386 (N_17386,N_12316,N_12627);
nor U17387 (N_17387,N_11706,N_13653);
xor U17388 (N_17388,N_12359,N_14575);
or U17389 (N_17389,N_10559,N_11120);
and U17390 (N_17390,N_13651,N_11535);
nand U17391 (N_17391,N_11853,N_10446);
xor U17392 (N_17392,N_12622,N_12989);
nand U17393 (N_17393,N_14585,N_13163);
or U17394 (N_17394,N_14606,N_12414);
or U17395 (N_17395,N_13543,N_11773);
nor U17396 (N_17396,N_13567,N_13032);
xor U17397 (N_17397,N_14811,N_11023);
or U17398 (N_17398,N_10741,N_13840);
and U17399 (N_17399,N_12677,N_10593);
or U17400 (N_17400,N_10659,N_13643);
nand U17401 (N_17401,N_13262,N_14294);
or U17402 (N_17402,N_10322,N_14155);
and U17403 (N_17403,N_13478,N_14055);
and U17404 (N_17404,N_11039,N_11363);
nor U17405 (N_17405,N_11922,N_11721);
xor U17406 (N_17406,N_10685,N_12440);
nor U17407 (N_17407,N_10576,N_14917);
or U17408 (N_17408,N_12462,N_14116);
and U17409 (N_17409,N_13309,N_12136);
xor U17410 (N_17410,N_10396,N_11419);
xnor U17411 (N_17411,N_13096,N_10367);
or U17412 (N_17412,N_13575,N_14403);
nor U17413 (N_17413,N_11473,N_10681);
and U17414 (N_17414,N_13734,N_12522);
and U17415 (N_17415,N_12921,N_11424);
nor U17416 (N_17416,N_11037,N_14581);
xnor U17417 (N_17417,N_10594,N_11098);
and U17418 (N_17418,N_10708,N_12190);
xnor U17419 (N_17419,N_11405,N_12869);
nor U17420 (N_17420,N_11795,N_12805);
xnor U17421 (N_17421,N_14871,N_10725);
xnor U17422 (N_17422,N_11611,N_11095);
or U17423 (N_17423,N_10955,N_10492);
nand U17424 (N_17424,N_14035,N_12517);
and U17425 (N_17425,N_11411,N_13107);
and U17426 (N_17426,N_10461,N_14113);
or U17427 (N_17427,N_12643,N_12894);
and U17428 (N_17428,N_13919,N_14447);
xor U17429 (N_17429,N_10807,N_10038);
xnor U17430 (N_17430,N_14749,N_14084);
nor U17431 (N_17431,N_10173,N_11636);
and U17432 (N_17432,N_14951,N_10608);
nor U17433 (N_17433,N_11645,N_11319);
xor U17434 (N_17434,N_11874,N_13132);
and U17435 (N_17435,N_12096,N_14840);
nand U17436 (N_17436,N_14258,N_14289);
or U17437 (N_17437,N_13002,N_14769);
and U17438 (N_17438,N_10404,N_12405);
xor U17439 (N_17439,N_13409,N_10637);
xnor U17440 (N_17440,N_13432,N_11125);
or U17441 (N_17441,N_13457,N_14109);
nand U17442 (N_17442,N_12461,N_13294);
and U17443 (N_17443,N_12163,N_11980);
and U17444 (N_17444,N_14473,N_10200);
and U17445 (N_17445,N_12815,N_10314);
and U17446 (N_17446,N_13431,N_13500);
or U17447 (N_17447,N_11019,N_14300);
or U17448 (N_17448,N_14706,N_13339);
nand U17449 (N_17449,N_14165,N_14889);
nor U17450 (N_17450,N_10541,N_10563);
or U17451 (N_17451,N_14312,N_11762);
nor U17452 (N_17452,N_12906,N_10394);
nor U17453 (N_17453,N_14408,N_14781);
nand U17454 (N_17454,N_10039,N_12937);
or U17455 (N_17455,N_14533,N_10135);
or U17456 (N_17456,N_10117,N_12106);
nor U17457 (N_17457,N_10372,N_11458);
nand U17458 (N_17458,N_11225,N_10811);
nand U17459 (N_17459,N_10211,N_10801);
or U17460 (N_17460,N_10776,N_14241);
and U17461 (N_17461,N_14446,N_11397);
or U17462 (N_17462,N_12580,N_14833);
nand U17463 (N_17463,N_13492,N_11977);
nor U17464 (N_17464,N_14138,N_11951);
nor U17465 (N_17465,N_13200,N_10037);
and U17466 (N_17466,N_11667,N_10517);
or U17467 (N_17467,N_14101,N_13122);
and U17468 (N_17468,N_11756,N_11688);
and U17469 (N_17469,N_14324,N_12369);
nor U17470 (N_17470,N_11045,N_14189);
nand U17471 (N_17471,N_13796,N_14444);
and U17472 (N_17472,N_13443,N_13495);
nor U17473 (N_17473,N_11682,N_11710);
nand U17474 (N_17474,N_13987,N_11568);
or U17475 (N_17475,N_10660,N_11538);
xnor U17476 (N_17476,N_10311,N_10756);
or U17477 (N_17477,N_14195,N_10768);
nor U17478 (N_17478,N_14590,N_13993);
nand U17479 (N_17479,N_12698,N_11168);
or U17480 (N_17480,N_11730,N_12878);
xnor U17481 (N_17481,N_12437,N_14709);
or U17482 (N_17482,N_11488,N_14710);
or U17483 (N_17483,N_10722,N_10867);
nand U17484 (N_17484,N_11938,N_14691);
nor U17485 (N_17485,N_11815,N_12415);
or U17486 (N_17486,N_14332,N_13790);
xor U17487 (N_17487,N_14167,N_14592);
and U17488 (N_17488,N_11755,N_14842);
nand U17489 (N_17489,N_14004,N_13823);
and U17490 (N_17490,N_13539,N_13001);
or U17491 (N_17491,N_11082,N_13473);
xor U17492 (N_17492,N_12664,N_12886);
xnor U17493 (N_17493,N_14466,N_10715);
nor U17494 (N_17494,N_10831,N_13285);
xnor U17495 (N_17495,N_14777,N_13439);
or U17496 (N_17496,N_14981,N_14325);
nor U17497 (N_17497,N_11984,N_12392);
or U17498 (N_17498,N_13899,N_13864);
nor U17499 (N_17499,N_11863,N_10870);
xnor U17500 (N_17500,N_13173,N_10240);
and U17501 (N_17501,N_14034,N_13836);
or U17502 (N_17502,N_12680,N_14826);
and U17503 (N_17503,N_11331,N_12605);
nor U17504 (N_17504,N_14406,N_14772);
nor U17505 (N_17505,N_10360,N_11022);
or U17506 (N_17506,N_10393,N_12008);
and U17507 (N_17507,N_10099,N_10495);
nand U17508 (N_17508,N_14347,N_10277);
nand U17509 (N_17509,N_11275,N_13824);
xnor U17510 (N_17510,N_14057,N_10298);
and U17511 (N_17511,N_12244,N_10267);
and U17512 (N_17512,N_13816,N_10411);
nor U17513 (N_17513,N_10607,N_13995);
or U17514 (N_17514,N_14603,N_11955);
nor U17515 (N_17515,N_11603,N_11981);
and U17516 (N_17516,N_10741,N_12798);
and U17517 (N_17517,N_10079,N_12901);
nor U17518 (N_17518,N_14376,N_10677);
nand U17519 (N_17519,N_14687,N_13231);
or U17520 (N_17520,N_10953,N_14476);
and U17521 (N_17521,N_10355,N_12112);
xnor U17522 (N_17522,N_10111,N_14490);
or U17523 (N_17523,N_10137,N_11199);
nand U17524 (N_17524,N_13565,N_13870);
or U17525 (N_17525,N_12095,N_10724);
nand U17526 (N_17526,N_13409,N_12211);
and U17527 (N_17527,N_10645,N_13960);
or U17528 (N_17528,N_13005,N_10656);
xor U17529 (N_17529,N_10004,N_13679);
nor U17530 (N_17530,N_10886,N_10812);
nor U17531 (N_17531,N_11266,N_14986);
nand U17532 (N_17532,N_14758,N_14119);
or U17533 (N_17533,N_10404,N_11651);
and U17534 (N_17534,N_13283,N_11044);
nor U17535 (N_17535,N_10245,N_12020);
nand U17536 (N_17536,N_13881,N_14086);
nand U17537 (N_17537,N_13064,N_13222);
nand U17538 (N_17538,N_14145,N_14422);
or U17539 (N_17539,N_14799,N_12894);
nor U17540 (N_17540,N_13586,N_10620);
and U17541 (N_17541,N_10690,N_11157);
xnor U17542 (N_17542,N_10361,N_13517);
nor U17543 (N_17543,N_13677,N_12126);
nor U17544 (N_17544,N_14958,N_13767);
nor U17545 (N_17545,N_13092,N_14415);
xnor U17546 (N_17546,N_11659,N_10844);
and U17547 (N_17547,N_14204,N_11737);
or U17548 (N_17548,N_11176,N_12358);
or U17549 (N_17549,N_11309,N_14655);
nand U17550 (N_17550,N_13900,N_11009);
and U17551 (N_17551,N_12167,N_11339);
nand U17552 (N_17552,N_11442,N_14016);
or U17553 (N_17553,N_14690,N_11809);
nand U17554 (N_17554,N_10959,N_10031);
nand U17555 (N_17555,N_10861,N_14892);
xor U17556 (N_17556,N_14873,N_13051);
nor U17557 (N_17557,N_13599,N_14956);
nand U17558 (N_17558,N_13365,N_12792);
or U17559 (N_17559,N_10696,N_14078);
xnor U17560 (N_17560,N_10674,N_12476);
and U17561 (N_17561,N_11057,N_11233);
and U17562 (N_17562,N_12550,N_12140);
nand U17563 (N_17563,N_14047,N_14135);
xor U17564 (N_17564,N_11153,N_12643);
xnor U17565 (N_17565,N_14254,N_14147);
xor U17566 (N_17566,N_14953,N_13883);
or U17567 (N_17567,N_14389,N_13003);
xnor U17568 (N_17568,N_10226,N_14742);
xor U17569 (N_17569,N_13080,N_12868);
nand U17570 (N_17570,N_13536,N_12601);
nor U17571 (N_17571,N_12153,N_10842);
nand U17572 (N_17572,N_14832,N_12174);
and U17573 (N_17573,N_13568,N_12253);
or U17574 (N_17574,N_13414,N_11302);
xor U17575 (N_17575,N_11374,N_10150);
and U17576 (N_17576,N_14626,N_11895);
nor U17577 (N_17577,N_10164,N_12441);
and U17578 (N_17578,N_12877,N_12619);
nand U17579 (N_17579,N_13240,N_14726);
nor U17580 (N_17580,N_12201,N_10420);
and U17581 (N_17581,N_13205,N_10259);
or U17582 (N_17582,N_14663,N_13593);
and U17583 (N_17583,N_13245,N_10263);
or U17584 (N_17584,N_12515,N_11955);
and U17585 (N_17585,N_12630,N_14632);
nor U17586 (N_17586,N_12179,N_11683);
and U17587 (N_17587,N_11100,N_10769);
xor U17588 (N_17588,N_13270,N_12742);
nand U17589 (N_17589,N_12340,N_11506);
or U17590 (N_17590,N_12289,N_13683);
or U17591 (N_17591,N_11593,N_10090);
or U17592 (N_17592,N_14581,N_13087);
or U17593 (N_17593,N_13408,N_13187);
nor U17594 (N_17594,N_13655,N_10074);
xor U17595 (N_17595,N_14179,N_14388);
or U17596 (N_17596,N_14068,N_13122);
and U17597 (N_17597,N_13681,N_14221);
and U17598 (N_17598,N_14000,N_11953);
and U17599 (N_17599,N_11160,N_11531);
or U17600 (N_17600,N_11222,N_13277);
nor U17601 (N_17601,N_13085,N_11729);
and U17602 (N_17602,N_12299,N_13906);
xnor U17603 (N_17603,N_10097,N_13164);
nand U17604 (N_17604,N_11464,N_11359);
nand U17605 (N_17605,N_14727,N_12822);
xnor U17606 (N_17606,N_13386,N_10598);
or U17607 (N_17607,N_14148,N_10407);
nand U17608 (N_17608,N_13565,N_11634);
nor U17609 (N_17609,N_14101,N_10127);
or U17610 (N_17610,N_13319,N_10109);
nor U17611 (N_17611,N_12142,N_11459);
or U17612 (N_17612,N_14286,N_13838);
nand U17613 (N_17613,N_10073,N_11165);
xnor U17614 (N_17614,N_10866,N_10724);
and U17615 (N_17615,N_14134,N_13362);
nand U17616 (N_17616,N_10944,N_13303);
nand U17617 (N_17617,N_11625,N_11030);
or U17618 (N_17618,N_12789,N_12199);
nor U17619 (N_17619,N_13182,N_13391);
or U17620 (N_17620,N_10318,N_11453);
nor U17621 (N_17621,N_13671,N_12583);
xor U17622 (N_17622,N_12396,N_13997);
nor U17623 (N_17623,N_13158,N_11402);
nor U17624 (N_17624,N_12568,N_13710);
nor U17625 (N_17625,N_10174,N_11611);
nand U17626 (N_17626,N_12282,N_14389);
nand U17627 (N_17627,N_10238,N_10524);
and U17628 (N_17628,N_11917,N_13135);
nand U17629 (N_17629,N_10664,N_14555);
xor U17630 (N_17630,N_12259,N_13939);
and U17631 (N_17631,N_11599,N_10571);
nor U17632 (N_17632,N_10968,N_10812);
nor U17633 (N_17633,N_10754,N_12230);
nand U17634 (N_17634,N_10583,N_11301);
nor U17635 (N_17635,N_14637,N_12628);
xnor U17636 (N_17636,N_10390,N_12540);
or U17637 (N_17637,N_13653,N_12666);
nand U17638 (N_17638,N_10521,N_14450);
xnor U17639 (N_17639,N_13634,N_13465);
or U17640 (N_17640,N_13128,N_12824);
nor U17641 (N_17641,N_11403,N_13542);
nor U17642 (N_17642,N_11682,N_11448);
and U17643 (N_17643,N_13503,N_11915);
nand U17644 (N_17644,N_10446,N_14290);
or U17645 (N_17645,N_11468,N_14527);
nand U17646 (N_17646,N_13564,N_14604);
or U17647 (N_17647,N_11722,N_14744);
xnor U17648 (N_17648,N_13143,N_14360);
xnor U17649 (N_17649,N_12864,N_12376);
nor U17650 (N_17650,N_10603,N_14169);
nand U17651 (N_17651,N_11546,N_11096);
nor U17652 (N_17652,N_11559,N_12285);
nor U17653 (N_17653,N_14376,N_11916);
nand U17654 (N_17654,N_12894,N_12997);
nor U17655 (N_17655,N_13418,N_14111);
xnor U17656 (N_17656,N_13742,N_14918);
xnor U17657 (N_17657,N_12267,N_11823);
and U17658 (N_17658,N_13374,N_11668);
xnor U17659 (N_17659,N_12794,N_14915);
and U17660 (N_17660,N_10859,N_12657);
or U17661 (N_17661,N_12011,N_12910);
nand U17662 (N_17662,N_14935,N_12874);
nor U17663 (N_17663,N_14254,N_12373);
and U17664 (N_17664,N_12244,N_10755);
nor U17665 (N_17665,N_11122,N_12907);
nand U17666 (N_17666,N_12962,N_11055);
nor U17667 (N_17667,N_14015,N_13629);
or U17668 (N_17668,N_10341,N_14437);
or U17669 (N_17669,N_14696,N_10541);
nand U17670 (N_17670,N_10884,N_10200);
nor U17671 (N_17671,N_11404,N_11209);
nand U17672 (N_17672,N_13625,N_10641);
and U17673 (N_17673,N_12193,N_11324);
or U17674 (N_17674,N_11470,N_13547);
xor U17675 (N_17675,N_11428,N_10084);
nor U17676 (N_17676,N_11293,N_10823);
or U17677 (N_17677,N_11436,N_11784);
nand U17678 (N_17678,N_11466,N_11235);
nor U17679 (N_17679,N_12374,N_12381);
nand U17680 (N_17680,N_14475,N_11015);
nor U17681 (N_17681,N_14078,N_10152);
and U17682 (N_17682,N_12858,N_13009);
xnor U17683 (N_17683,N_10639,N_13855);
xor U17684 (N_17684,N_13691,N_10395);
and U17685 (N_17685,N_12615,N_13910);
and U17686 (N_17686,N_11076,N_12570);
xnor U17687 (N_17687,N_12251,N_11809);
xor U17688 (N_17688,N_11607,N_11723);
xor U17689 (N_17689,N_10725,N_13826);
nor U17690 (N_17690,N_12386,N_11878);
xnor U17691 (N_17691,N_11253,N_10667);
or U17692 (N_17692,N_13247,N_11896);
and U17693 (N_17693,N_11255,N_13333);
and U17694 (N_17694,N_11060,N_13436);
or U17695 (N_17695,N_13623,N_14001);
xnor U17696 (N_17696,N_13513,N_14103);
nor U17697 (N_17697,N_14942,N_14560);
and U17698 (N_17698,N_12537,N_12665);
nand U17699 (N_17699,N_12270,N_11194);
or U17700 (N_17700,N_14880,N_14030);
and U17701 (N_17701,N_14910,N_10112);
nand U17702 (N_17702,N_13414,N_12370);
or U17703 (N_17703,N_14411,N_10945);
or U17704 (N_17704,N_10176,N_10138);
nor U17705 (N_17705,N_11483,N_12368);
nand U17706 (N_17706,N_14911,N_10719);
nand U17707 (N_17707,N_12755,N_13104);
or U17708 (N_17708,N_10475,N_10739);
xor U17709 (N_17709,N_10456,N_10265);
or U17710 (N_17710,N_10474,N_14621);
nand U17711 (N_17711,N_11418,N_13111);
nor U17712 (N_17712,N_14177,N_12367);
xnor U17713 (N_17713,N_14149,N_12278);
or U17714 (N_17714,N_11375,N_14486);
nand U17715 (N_17715,N_11345,N_14301);
and U17716 (N_17716,N_11423,N_12787);
and U17717 (N_17717,N_12863,N_12002);
or U17718 (N_17718,N_14973,N_12966);
and U17719 (N_17719,N_12626,N_13839);
nor U17720 (N_17720,N_13316,N_12253);
nand U17721 (N_17721,N_13040,N_14936);
and U17722 (N_17722,N_12618,N_14545);
nand U17723 (N_17723,N_13935,N_14050);
and U17724 (N_17724,N_10193,N_14832);
xor U17725 (N_17725,N_12946,N_11971);
and U17726 (N_17726,N_10626,N_10750);
or U17727 (N_17727,N_11106,N_14991);
nor U17728 (N_17728,N_12678,N_13049);
nand U17729 (N_17729,N_11583,N_10450);
nor U17730 (N_17730,N_14997,N_11831);
or U17731 (N_17731,N_10613,N_12413);
and U17732 (N_17732,N_12826,N_10858);
xnor U17733 (N_17733,N_11135,N_11539);
or U17734 (N_17734,N_14377,N_11231);
nor U17735 (N_17735,N_13146,N_11101);
and U17736 (N_17736,N_12998,N_11472);
nor U17737 (N_17737,N_13407,N_14752);
or U17738 (N_17738,N_12122,N_12950);
nand U17739 (N_17739,N_12759,N_11356);
or U17740 (N_17740,N_12047,N_14183);
nor U17741 (N_17741,N_12145,N_10506);
or U17742 (N_17742,N_11758,N_13038);
nand U17743 (N_17743,N_11479,N_14785);
nand U17744 (N_17744,N_13854,N_14401);
or U17745 (N_17745,N_11105,N_12072);
nand U17746 (N_17746,N_13688,N_12544);
or U17747 (N_17747,N_13658,N_13752);
nor U17748 (N_17748,N_12794,N_12636);
nand U17749 (N_17749,N_10304,N_11713);
nor U17750 (N_17750,N_14808,N_10814);
and U17751 (N_17751,N_14800,N_10138);
and U17752 (N_17752,N_10912,N_13642);
xor U17753 (N_17753,N_12212,N_10978);
and U17754 (N_17754,N_10051,N_11874);
xnor U17755 (N_17755,N_13905,N_12624);
nand U17756 (N_17756,N_12020,N_14125);
or U17757 (N_17757,N_10604,N_12248);
nand U17758 (N_17758,N_12836,N_10105);
and U17759 (N_17759,N_11417,N_11850);
nand U17760 (N_17760,N_10352,N_14364);
or U17761 (N_17761,N_10898,N_14187);
xor U17762 (N_17762,N_13952,N_11709);
nor U17763 (N_17763,N_11017,N_13432);
nor U17764 (N_17764,N_11699,N_14234);
or U17765 (N_17765,N_13878,N_10476);
nor U17766 (N_17766,N_10597,N_12159);
xnor U17767 (N_17767,N_14237,N_11809);
or U17768 (N_17768,N_13399,N_12464);
nand U17769 (N_17769,N_12835,N_12589);
and U17770 (N_17770,N_14829,N_10319);
xor U17771 (N_17771,N_12161,N_12392);
or U17772 (N_17772,N_12943,N_13344);
nand U17773 (N_17773,N_11773,N_10708);
or U17774 (N_17774,N_10933,N_14412);
nand U17775 (N_17775,N_11497,N_12593);
xnor U17776 (N_17776,N_13591,N_11527);
xor U17777 (N_17777,N_12706,N_10198);
nand U17778 (N_17778,N_13891,N_14895);
or U17779 (N_17779,N_10663,N_11842);
xor U17780 (N_17780,N_10240,N_13394);
or U17781 (N_17781,N_14794,N_12845);
nor U17782 (N_17782,N_12408,N_13423);
or U17783 (N_17783,N_11073,N_14951);
xor U17784 (N_17784,N_13912,N_11278);
nor U17785 (N_17785,N_10994,N_14381);
nand U17786 (N_17786,N_10273,N_11804);
xor U17787 (N_17787,N_13262,N_13449);
xor U17788 (N_17788,N_11835,N_10374);
and U17789 (N_17789,N_14201,N_11018);
nand U17790 (N_17790,N_13597,N_10598);
and U17791 (N_17791,N_13035,N_10935);
or U17792 (N_17792,N_11270,N_13371);
and U17793 (N_17793,N_11109,N_12239);
nor U17794 (N_17794,N_13602,N_10928);
or U17795 (N_17795,N_13333,N_14233);
and U17796 (N_17796,N_11390,N_12149);
or U17797 (N_17797,N_10710,N_14210);
xnor U17798 (N_17798,N_10058,N_12015);
xnor U17799 (N_17799,N_12254,N_10094);
or U17800 (N_17800,N_13888,N_12217);
nor U17801 (N_17801,N_12273,N_12761);
and U17802 (N_17802,N_12665,N_10978);
or U17803 (N_17803,N_11581,N_12572);
nor U17804 (N_17804,N_10285,N_14297);
nor U17805 (N_17805,N_12611,N_10759);
nand U17806 (N_17806,N_10456,N_11599);
nand U17807 (N_17807,N_11923,N_13698);
xnor U17808 (N_17808,N_11431,N_10513);
xnor U17809 (N_17809,N_10186,N_10565);
xnor U17810 (N_17810,N_12299,N_11436);
xnor U17811 (N_17811,N_12594,N_11316);
xor U17812 (N_17812,N_10885,N_10875);
or U17813 (N_17813,N_13652,N_11173);
nand U17814 (N_17814,N_13573,N_14698);
xor U17815 (N_17815,N_12572,N_10956);
and U17816 (N_17816,N_10558,N_11088);
nand U17817 (N_17817,N_12774,N_10923);
and U17818 (N_17818,N_14894,N_14387);
nor U17819 (N_17819,N_10446,N_11895);
or U17820 (N_17820,N_10613,N_13216);
or U17821 (N_17821,N_11062,N_14107);
and U17822 (N_17822,N_10871,N_10798);
nor U17823 (N_17823,N_13743,N_11189);
nand U17824 (N_17824,N_13301,N_10011);
nor U17825 (N_17825,N_12043,N_14757);
xnor U17826 (N_17826,N_12793,N_14516);
or U17827 (N_17827,N_11081,N_14119);
nand U17828 (N_17828,N_12487,N_13373);
nand U17829 (N_17829,N_12404,N_14969);
nand U17830 (N_17830,N_11108,N_13525);
xor U17831 (N_17831,N_13371,N_14483);
nor U17832 (N_17832,N_14526,N_10392);
nand U17833 (N_17833,N_10207,N_12367);
nor U17834 (N_17834,N_12416,N_14401);
nand U17835 (N_17835,N_12270,N_12806);
xnor U17836 (N_17836,N_10163,N_10550);
or U17837 (N_17837,N_10004,N_14315);
or U17838 (N_17838,N_10416,N_11653);
or U17839 (N_17839,N_11091,N_10161);
xor U17840 (N_17840,N_10103,N_10185);
nand U17841 (N_17841,N_11686,N_13703);
nand U17842 (N_17842,N_13792,N_14590);
or U17843 (N_17843,N_12461,N_10612);
and U17844 (N_17844,N_10039,N_13265);
xnor U17845 (N_17845,N_13536,N_10073);
xor U17846 (N_17846,N_10660,N_11082);
xnor U17847 (N_17847,N_10528,N_14626);
or U17848 (N_17848,N_12474,N_12096);
and U17849 (N_17849,N_11956,N_12201);
or U17850 (N_17850,N_13998,N_13025);
or U17851 (N_17851,N_11307,N_13133);
xnor U17852 (N_17852,N_13873,N_14375);
nor U17853 (N_17853,N_13581,N_11562);
and U17854 (N_17854,N_14001,N_13375);
nand U17855 (N_17855,N_14974,N_13228);
xor U17856 (N_17856,N_12811,N_11813);
nor U17857 (N_17857,N_11672,N_12783);
and U17858 (N_17858,N_13741,N_10026);
xnor U17859 (N_17859,N_13719,N_11896);
or U17860 (N_17860,N_10660,N_10851);
nor U17861 (N_17861,N_12328,N_13958);
and U17862 (N_17862,N_12512,N_14961);
or U17863 (N_17863,N_12039,N_11588);
and U17864 (N_17864,N_11908,N_10728);
nor U17865 (N_17865,N_12041,N_11078);
xor U17866 (N_17866,N_14941,N_10438);
xor U17867 (N_17867,N_10861,N_12000);
nand U17868 (N_17868,N_10478,N_12202);
xnor U17869 (N_17869,N_13458,N_10661);
or U17870 (N_17870,N_11681,N_13551);
or U17871 (N_17871,N_14567,N_10317);
nand U17872 (N_17872,N_11455,N_12031);
nor U17873 (N_17873,N_12778,N_13526);
nor U17874 (N_17874,N_10963,N_13016);
nor U17875 (N_17875,N_12667,N_13425);
and U17876 (N_17876,N_11255,N_11126);
xnor U17877 (N_17877,N_10103,N_11273);
xor U17878 (N_17878,N_13386,N_12261);
or U17879 (N_17879,N_13874,N_13574);
and U17880 (N_17880,N_13381,N_13796);
or U17881 (N_17881,N_12806,N_11121);
or U17882 (N_17882,N_10234,N_11093);
nand U17883 (N_17883,N_13011,N_14978);
xnor U17884 (N_17884,N_11050,N_10400);
or U17885 (N_17885,N_13690,N_11454);
nand U17886 (N_17886,N_14199,N_11567);
nand U17887 (N_17887,N_12327,N_14506);
nor U17888 (N_17888,N_12156,N_11874);
nor U17889 (N_17889,N_14508,N_14712);
nand U17890 (N_17890,N_12259,N_13715);
nand U17891 (N_17891,N_14686,N_12972);
or U17892 (N_17892,N_14474,N_12283);
nor U17893 (N_17893,N_13751,N_13845);
and U17894 (N_17894,N_13300,N_11142);
or U17895 (N_17895,N_14744,N_10386);
xor U17896 (N_17896,N_11975,N_10566);
and U17897 (N_17897,N_13188,N_12049);
nand U17898 (N_17898,N_11213,N_14740);
or U17899 (N_17899,N_12256,N_10749);
nor U17900 (N_17900,N_12262,N_12664);
or U17901 (N_17901,N_14125,N_14660);
nor U17902 (N_17902,N_13670,N_12758);
or U17903 (N_17903,N_12516,N_14784);
or U17904 (N_17904,N_11850,N_10204);
xnor U17905 (N_17905,N_13850,N_13125);
or U17906 (N_17906,N_13435,N_11526);
or U17907 (N_17907,N_11794,N_11607);
xor U17908 (N_17908,N_11521,N_12871);
nor U17909 (N_17909,N_12961,N_10249);
xor U17910 (N_17910,N_13369,N_11390);
and U17911 (N_17911,N_13435,N_11454);
xor U17912 (N_17912,N_14515,N_12154);
nor U17913 (N_17913,N_12936,N_10984);
nor U17914 (N_17914,N_10749,N_12546);
xor U17915 (N_17915,N_13417,N_12755);
and U17916 (N_17916,N_10788,N_14940);
nand U17917 (N_17917,N_12651,N_13725);
or U17918 (N_17918,N_12235,N_12432);
nand U17919 (N_17919,N_12103,N_10958);
and U17920 (N_17920,N_14521,N_12586);
nand U17921 (N_17921,N_12103,N_10441);
xor U17922 (N_17922,N_10700,N_14705);
nor U17923 (N_17923,N_13389,N_10342);
and U17924 (N_17924,N_11000,N_10798);
nor U17925 (N_17925,N_11189,N_14316);
nand U17926 (N_17926,N_11223,N_11918);
nand U17927 (N_17927,N_11940,N_10834);
xnor U17928 (N_17928,N_10888,N_11804);
nor U17929 (N_17929,N_11237,N_11580);
nor U17930 (N_17930,N_10592,N_14960);
and U17931 (N_17931,N_12455,N_14359);
nand U17932 (N_17932,N_13538,N_13533);
or U17933 (N_17933,N_10519,N_12631);
xnor U17934 (N_17934,N_11432,N_14754);
nand U17935 (N_17935,N_11425,N_14567);
nor U17936 (N_17936,N_10649,N_12334);
or U17937 (N_17937,N_12036,N_12787);
or U17938 (N_17938,N_11963,N_12135);
nand U17939 (N_17939,N_11223,N_13247);
nor U17940 (N_17940,N_11319,N_12997);
or U17941 (N_17941,N_12156,N_14025);
nor U17942 (N_17942,N_14936,N_12883);
nor U17943 (N_17943,N_14771,N_12428);
nor U17944 (N_17944,N_11009,N_11784);
nor U17945 (N_17945,N_10055,N_13549);
nor U17946 (N_17946,N_13650,N_10631);
and U17947 (N_17947,N_13336,N_13225);
xnor U17948 (N_17948,N_14776,N_12230);
or U17949 (N_17949,N_10464,N_13137);
or U17950 (N_17950,N_10837,N_13888);
nor U17951 (N_17951,N_11069,N_13839);
xor U17952 (N_17952,N_11227,N_10130);
nor U17953 (N_17953,N_13399,N_10469);
xor U17954 (N_17954,N_12180,N_11677);
or U17955 (N_17955,N_10059,N_10378);
xnor U17956 (N_17956,N_11478,N_13924);
and U17957 (N_17957,N_13341,N_13585);
or U17958 (N_17958,N_10859,N_10055);
nand U17959 (N_17959,N_13719,N_14030);
xnor U17960 (N_17960,N_10363,N_12855);
nor U17961 (N_17961,N_12896,N_13030);
or U17962 (N_17962,N_14497,N_14533);
nor U17963 (N_17963,N_10378,N_12662);
nor U17964 (N_17964,N_12824,N_13958);
and U17965 (N_17965,N_12651,N_11006);
or U17966 (N_17966,N_10406,N_11867);
xor U17967 (N_17967,N_14017,N_12564);
and U17968 (N_17968,N_11483,N_10363);
nor U17969 (N_17969,N_12513,N_13459);
or U17970 (N_17970,N_12796,N_13022);
nand U17971 (N_17971,N_11466,N_11552);
nor U17972 (N_17972,N_14547,N_14978);
nor U17973 (N_17973,N_13183,N_11289);
nand U17974 (N_17974,N_10211,N_11634);
or U17975 (N_17975,N_14152,N_11959);
nor U17976 (N_17976,N_10929,N_10543);
nand U17977 (N_17977,N_11325,N_14377);
or U17978 (N_17978,N_11539,N_10877);
and U17979 (N_17979,N_14848,N_10594);
nand U17980 (N_17980,N_13676,N_14682);
and U17981 (N_17981,N_12039,N_10773);
or U17982 (N_17982,N_14116,N_11760);
or U17983 (N_17983,N_14570,N_11809);
or U17984 (N_17984,N_12470,N_10590);
nor U17985 (N_17985,N_13295,N_12046);
nand U17986 (N_17986,N_13641,N_10741);
nor U17987 (N_17987,N_14603,N_13342);
nand U17988 (N_17988,N_14747,N_12779);
or U17989 (N_17989,N_10259,N_14521);
nand U17990 (N_17990,N_14815,N_10256);
or U17991 (N_17991,N_14571,N_12195);
xnor U17992 (N_17992,N_12414,N_14634);
and U17993 (N_17993,N_11872,N_13040);
and U17994 (N_17994,N_12959,N_13838);
nor U17995 (N_17995,N_12792,N_10587);
and U17996 (N_17996,N_14494,N_12160);
or U17997 (N_17997,N_14229,N_14745);
nor U17998 (N_17998,N_13933,N_13805);
or U17999 (N_17999,N_11752,N_13367);
or U18000 (N_18000,N_10068,N_13349);
nand U18001 (N_18001,N_11407,N_13802);
and U18002 (N_18002,N_14404,N_11238);
nand U18003 (N_18003,N_12228,N_11327);
xnor U18004 (N_18004,N_14071,N_10342);
and U18005 (N_18005,N_11384,N_10324);
or U18006 (N_18006,N_13203,N_13932);
or U18007 (N_18007,N_14232,N_10128);
xnor U18008 (N_18008,N_13092,N_13069);
and U18009 (N_18009,N_12296,N_14416);
nor U18010 (N_18010,N_12020,N_10045);
and U18011 (N_18011,N_14799,N_11067);
xnor U18012 (N_18012,N_13003,N_12390);
and U18013 (N_18013,N_13428,N_14834);
nand U18014 (N_18014,N_11055,N_14815);
nor U18015 (N_18015,N_10269,N_11573);
nand U18016 (N_18016,N_13611,N_12855);
nand U18017 (N_18017,N_10369,N_12738);
nand U18018 (N_18018,N_12616,N_13174);
or U18019 (N_18019,N_12813,N_14169);
and U18020 (N_18020,N_10136,N_14600);
and U18021 (N_18021,N_10218,N_10692);
or U18022 (N_18022,N_12188,N_13741);
nand U18023 (N_18023,N_10259,N_14686);
nand U18024 (N_18024,N_11012,N_10296);
xnor U18025 (N_18025,N_10555,N_10196);
xnor U18026 (N_18026,N_14344,N_11460);
xor U18027 (N_18027,N_12556,N_13571);
xor U18028 (N_18028,N_13044,N_11941);
nor U18029 (N_18029,N_13284,N_10912);
nor U18030 (N_18030,N_11493,N_10673);
nand U18031 (N_18031,N_14273,N_11508);
nor U18032 (N_18032,N_11286,N_11168);
nand U18033 (N_18033,N_11432,N_14404);
or U18034 (N_18034,N_12957,N_13240);
nor U18035 (N_18035,N_13127,N_10356);
xor U18036 (N_18036,N_10741,N_14605);
and U18037 (N_18037,N_13443,N_13007);
xnor U18038 (N_18038,N_12327,N_10728);
or U18039 (N_18039,N_12954,N_12706);
and U18040 (N_18040,N_12037,N_11721);
and U18041 (N_18041,N_11202,N_11441);
nand U18042 (N_18042,N_10018,N_11146);
and U18043 (N_18043,N_13336,N_14099);
xor U18044 (N_18044,N_14248,N_12994);
nand U18045 (N_18045,N_13786,N_14370);
or U18046 (N_18046,N_12397,N_11800);
xor U18047 (N_18047,N_11477,N_11692);
nand U18048 (N_18048,N_10419,N_12846);
nor U18049 (N_18049,N_13800,N_10903);
and U18050 (N_18050,N_14632,N_13350);
xor U18051 (N_18051,N_14931,N_12501);
nor U18052 (N_18052,N_13686,N_10332);
nor U18053 (N_18053,N_14700,N_14652);
nand U18054 (N_18054,N_13223,N_13431);
nor U18055 (N_18055,N_12775,N_10066);
xor U18056 (N_18056,N_11435,N_10882);
xor U18057 (N_18057,N_14905,N_12009);
xor U18058 (N_18058,N_14778,N_12367);
nor U18059 (N_18059,N_13726,N_13039);
nor U18060 (N_18060,N_13718,N_10897);
or U18061 (N_18061,N_12736,N_10689);
and U18062 (N_18062,N_11218,N_12260);
nand U18063 (N_18063,N_12307,N_10369);
or U18064 (N_18064,N_12947,N_10642);
xor U18065 (N_18065,N_13664,N_12522);
nor U18066 (N_18066,N_13720,N_10892);
or U18067 (N_18067,N_12206,N_12513);
nor U18068 (N_18068,N_14080,N_12033);
nor U18069 (N_18069,N_14784,N_10720);
and U18070 (N_18070,N_13556,N_12024);
xnor U18071 (N_18071,N_11608,N_10885);
nor U18072 (N_18072,N_12953,N_10081);
xnor U18073 (N_18073,N_10523,N_14850);
nor U18074 (N_18074,N_10198,N_14539);
nand U18075 (N_18075,N_11953,N_10489);
xnor U18076 (N_18076,N_11926,N_11871);
nand U18077 (N_18077,N_11565,N_10263);
or U18078 (N_18078,N_11131,N_13659);
and U18079 (N_18079,N_14633,N_12810);
and U18080 (N_18080,N_14264,N_14156);
nor U18081 (N_18081,N_14086,N_11531);
and U18082 (N_18082,N_13665,N_13025);
nand U18083 (N_18083,N_13196,N_14124);
or U18084 (N_18084,N_12648,N_12891);
nor U18085 (N_18085,N_11531,N_14532);
nor U18086 (N_18086,N_11850,N_12668);
nand U18087 (N_18087,N_12187,N_13594);
nand U18088 (N_18088,N_10965,N_10362);
nand U18089 (N_18089,N_11375,N_14321);
and U18090 (N_18090,N_12383,N_14187);
xnor U18091 (N_18091,N_12983,N_12074);
or U18092 (N_18092,N_10974,N_13033);
and U18093 (N_18093,N_14577,N_14505);
xnor U18094 (N_18094,N_10239,N_14689);
nand U18095 (N_18095,N_12177,N_14625);
or U18096 (N_18096,N_13222,N_12120);
and U18097 (N_18097,N_14083,N_10725);
xnor U18098 (N_18098,N_12259,N_13667);
or U18099 (N_18099,N_10812,N_11166);
or U18100 (N_18100,N_11446,N_10356);
nor U18101 (N_18101,N_13767,N_13750);
xor U18102 (N_18102,N_13742,N_10843);
nand U18103 (N_18103,N_12686,N_10517);
xnor U18104 (N_18104,N_14865,N_10533);
nor U18105 (N_18105,N_10251,N_13227);
nand U18106 (N_18106,N_14662,N_10566);
nor U18107 (N_18107,N_11628,N_10888);
nand U18108 (N_18108,N_10266,N_12451);
and U18109 (N_18109,N_11804,N_10089);
and U18110 (N_18110,N_14520,N_14583);
xnor U18111 (N_18111,N_12117,N_11851);
or U18112 (N_18112,N_14345,N_12210);
or U18113 (N_18113,N_13379,N_10660);
xor U18114 (N_18114,N_10388,N_14783);
and U18115 (N_18115,N_14161,N_11715);
nor U18116 (N_18116,N_12972,N_14035);
nor U18117 (N_18117,N_12314,N_12909);
xnor U18118 (N_18118,N_10689,N_12966);
nor U18119 (N_18119,N_14368,N_13308);
nand U18120 (N_18120,N_13021,N_12571);
nand U18121 (N_18121,N_14432,N_13652);
xor U18122 (N_18122,N_12225,N_14338);
nor U18123 (N_18123,N_12540,N_11730);
and U18124 (N_18124,N_11010,N_14699);
and U18125 (N_18125,N_11066,N_11984);
or U18126 (N_18126,N_13758,N_10433);
nand U18127 (N_18127,N_13874,N_10287);
nand U18128 (N_18128,N_12653,N_14458);
and U18129 (N_18129,N_11678,N_14062);
nor U18130 (N_18130,N_11427,N_13452);
xnor U18131 (N_18131,N_12645,N_11111);
and U18132 (N_18132,N_14479,N_11187);
or U18133 (N_18133,N_12208,N_13418);
and U18134 (N_18134,N_14011,N_11354);
nand U18135 (N_18135,N_10477,N_10005);
and U18136 (N_18136,N_14470,N_13774);
nor U18137 (N_18137,N_13373,N_10493);
nor U18138 (N_18138,N_13765,N_10531);
nand U18139 (N_18139,N_11361,N_11161);
nor U18140 (N_18140,N_10429,N_11579);
xor U18141 (N_18141,N_14418,N_13868);
nor U18142 (N_18142,N_14828,N_10007);
nand U18143 (N_18143,N_13444,N_13442);
or U18144 (N_18144,N_10705,N_11372);
and U18145 (N_18145,N_11871,N_14435);
xor U18146 (N_18146,N_12097,N_10999);
xor U18147 (N_18147,N_14490,N_10897);
xor U18148 (N_18148,N_14977,N_14953);
nand U18149 (N_18149,N_14237,N_13165);
or U18150 (N_18150,N_12653,N_13562);
or U18151 (N_18151,N_12332,N_10396);
nand U18152 (N_18152,N_11065,N_12574);
nand U18153 (N_18153,N_10767,N_14355);
and U18154 (N_18154,N_14596,N_12914);
nand U18155 (N_18155,N_12899,N_13126);
nand U18156 (N_18156,N_12986,N_11050);
nand U18157 (N_18157,N_12227,N_14249);
nor U18158 (N_18158,N_10963,N_13218);
and U18159 (N_18159,N_10197,N_12905);
xor U18160 (N_18160,N_13346,N_11754);
xnor U18161 (N_18161,N_11920,N_12131);
and U18162 (N_18162,N_12982,N_10453);
xnor U18163 (N_18163,N_12770,N_13274);
and U18164 (N_18164,N_10056,N_10238);
nand U18165 (N_18165,N_14871,N_10824);
nor U18166 (N_18166,N_13909,N_12922);
and U18167 (N_18167,N_10482,N_10199);
and U18168 (N_18168,N_10491,N_14895);
xnor U18169 (N_18169,N_12022,N_14214);
and U18170 (N_18170,N_10037,N_10238);
xor U18171 (N_18171,N_11566,N_12946);
and U18172 (N_18172,N_11063,N_13942);
xnor U18173 (N_18173,N_11414,N_13921);
xnor U18174 (N_18174,N_13215,N_10796);
nor U18175 (N_18175,N_10039,N_10500);
or U18176 (N_18176,N_14598,N_12946);
and U18177 (N_18177,N_13725,N_11138);
xor U18178 (N_18178,N_11848,N_14550);
or U18179 (N_18179,N_11395,N_10849);
or U18180 (N_18180,N_14749,N_13210);
nand U18181 (N_18181,N_12793,N_12569);
xor U18182 (N_18182,N_10738,N_10190);
and U18183 (N_18183,N_13592,N_10444);
nor U18184 (N_18184,N_10468,N_11462);
and U18185 (N_18185,N_11458,N_10771);
nor U18186 (N_18186,N_14030,N_12080);
or U18187 (N_18187,N_13448,N_10744);
nor U18188 (N_18188,N_12689,N_10247);
or U18189 (N_18189,N_11912,N_14580);
or U18190 (N_18190,N_10065,N_11673);
xor U18191 (N_18191,N_14297,N_10875);
nor U18192 (N_18192,N_10000,N_14952);
nor U18193 (N_18193,N_10664,N_12949);
nand U18194 (N_18194,N_10896,N_12284);
nor U18195 (N_18195,N_14117,N_10841);
nand U18196 (N_18196,N_10141,N_10899);
xnor U18197 (N_18197,N_14679,N_12547);
and U18198 (N_18198,N_13217,N_12563);
and U18199 (N_18199,N_13288,N_11625);
nor U18200 (N_18200,N_13328,N_13517);
and U18201 (N_18201,N_10517,N_14699);
and U18202 (N_18202,N_10920,N_10255);
nand U18203 (N_18203,N_13188,N_11461);
nor U18204 (N_18204,N_10319,N_12633);
nor U18205 (N_18205,N_10240,N_11939);
xor U18206 (N_18206,N_11448,N_14445);
or U18207 (N_18207,N_12904,N_12250);
nor U18208 (N_18208,N_13603,N_11150);
nor U18209 (N_18209,N_10412,N_14941);
and U18210 (N_18210,N_12846,N_11933);
xnor U18211 (N_18211,N_10916,N_14766);
and U18212 (N_18212,N_13212,N_14569);
nand U18213 (N_18213,N_14080,N_12192);
and U18214 (N_18214,N_11922,N_13485);
nor U18215 (N_18215,N_10059,N_14338);
xor U18216 (N_18216,N_10295,N_10882);
xor U18217 (N_18217,N_12188,N_14659);
or U18218 (N_18218,N_10428,N_12454);
nor U18219 (N_18219,N_11346,N_14449);
and U18220 (N_18220,N_12555,N_13170);
xnor U18221 (N_18221,N_12591,N_11782);
and U18222 (N_18222,N_13687,N_10013);
and U18223 (N_18223,N_10054,N_13305);
xor U18224 (N_18224,N_12856,N_12117);
and U18225 (N_18225,N_12760,N_12451);
xor U18226 (N_18226,N_12526,N_10297);
and U18227 (N_18227,N_11554,N_10490);
or U18228 (N_18228,N_14794,N_14611);
or U18229 (N_18229,N_11370,N_10871);
xnor U18230 (N_18230,N_12108,N_11328);
and U18231 (N_18231,N_12342,N_10699);
and U18232 (N_18232,N_14566,N_13350);
xor U18233 (N_18233,N_14067,N_10533);
or U18234 (N_18234,N_13116,N_12970);
and U18235 (N_18235,N_12404,N_12685);
or U18236 (N_18236,N_11263,N_13830);
nand U18237 (N_18237,N_13521,N_13798);
xnor U18238 (N_18238,N_12379,N_10807);
nand U18239 (N_18239,N_13800,N_11219);
xnor U18240 (N_18240,N_13037,N_12184);
nor U18241 (N_18241,N_13877,N_11800);
and U18242 (N_18242,N_12173,N_11179);
xnor U18243 (N_18243,N_11588,N_11300);
xnor U18244 (N_18244,N_13468,N_14307);
xnor U18245 (N_18245,N_13871,N_11656);
or U18246 (N_18246,N_10902,N_13355);
nand U18247 (N_18247,N_13499,N_14346);
nand U18248 (N_18248,N_10531,N_12826);
nand U18249 (N_18249,N_14233,N_13915);
or U18250 (N_18250,N_11660,N_13447);
or U18251 (N_18251,N_12382,N_10140);
xor U18252 (N_18252,N_10177,N_13612);
xnor U18253 (N_18253,N_13438,N_11596);
and U18254 (N_18254,N_12228,N_11074);
or U18255 (N_18255,N_13620,N_11212);
xor U18256 (N_18256,N_14096,N_11563);
nor U18257 (N_18257,N_14000,N_12684);
nor U18258 (N_18258,N_13182,N_12723);
xnor U18259 (N_18259,N_12597,N_10944);
nand U18260 (N_18260,N_13152,N_13910);
nor U18261 (N_18261,N_10485,N_10353);
nand U18262 (N_18262,N_14211,N_13419);
or U18263 (N_18263,N_12485,N_14757);
nor U18264 (N_18264,N_13346,N_12156);
or U18265 (N_18265,N_12016,N_14798);
xor U18266 (N_18266,N_12054,N_10230);
nor U18267 (N_18267,N_13640,N_14056);
and U18268 (N_18268,N_14041,N_10970);
and U18269 (N_18269,N_13690,N_10497);
xor U18270 (N_18270,N_13713,N_10832);
or U18271 (N_18271,N_14879,N_13501);
or U18272 (N_18272,N_14708,N_10502);
nand U18273 (N_18273,N_12675,N_12298);
nor U18274 (N_18274,N_10594,N_12868);
nor U18275 (N_18275,N_10791,N_13573);
xor U18276 (N_18276,N_11579,N_14344);
xor U18277 (N_18277,N_13450,N_13157);
xor U18278 (N_18278,N_13325,N_12904);
nand U18279 (N_18279,N_12837,N_14358);
nand U18280 (N_18280,N_11121,N_14990);
xnor U18281 (N_18281,N_12390,N_10117);
or U18282 (N_18282,N_13300,N_11587);
xnor U18283 (N_18283,N_12233,N_14598);
nand U18284 (N_18284,N_13008,N_11755);
xor U18285 (N_18285,N_14583,N_10508);
or U18286 (N_18286,N_12541,N_12259);
and U18287 (N_18287,N_11081,N_12753);
xnor U18288 (N_18288,N_14531,N_11461);
and U18289 (N_18289,N_12374,N_11084);
and U18290 (N_18290,N_13925,N_12005);
nand U18291 (N_18291,N_11642,N_13266);
xnor U18292 (N_18292,N_12681,N_10903);
nor U18293 (N_18293,N_10956,N_13606);
nor U18294 (N_18294,N_13316,N_11690);
xnor U18295 (N_18295,N_11685,N_13213);
nor U18296 (N_18296,N_14010,N_11978);
and U18297 (N_18297,N_14032,N_10113);
nor U18298 (N_18298,N_11711,N_14975);
and U18299 (N_18299,N_14351,N_13448);
and U18300 (N_18300,N_10936,N_11649);
or U18301 (N_18301,N_11303,N_12277);
or U18302 (N_18302,N_12321,N_10581);
xnor U18303 (N_18303,N_10480,N_14648);
and U18304 (N_18304,N_12885,N_12452);
and U18305 (N_18305,N_10157,N_10805);
and U18306 (N_18306,N_13521,N_13232);
or U18307 (N_18307,N_12435,N_11633);
or U18308 (N_18308,N_10617,N_11656);
nor U18309 (N_18309,N_11772,N_10301);
and U18310 (N_18310,N_10818,N_13174);
or U18311 (N_18311,N_14315,N_11166);
and U18312 (N_18312,N_10825,N_12978);
and U18313 (N_18313,N_11933,N_10497);
and U18314 (N_18314,N_10966,N_10586);
nor U18315 (N_18315,N_11483,N_10542);
xor U18316 (N_18316,N_11587,N_12800);
nand U18317 (N_18317,N_10320,N_10189);
xor U18318 (N_18318,N_11179,N_14217);
nor U18319 (N_18319,N_13951,N_12915);
nor U18320 (N_18320,N_12158,N_12054);
nor U18321 (N_18321,N_10656,N_14787);
and U18322 (N_18322,N_12784,N_11874);
or U18323 (N_18323,N_11505,N_11162);
xor U18324 (N_18324,N_14021,N_10670);
nand U18325 (N_18325,N_10159,N_13041);
nor U18326 (N_18326,N_13832,N_13561);
nand U18327 (N_18327,N_11334,N_10087);
or U18328 (N_18328,N_13790,N_14705);
nor U18329 (N_18329,N_14514,N_12923);
and U18330 (N_18330,N_14909,N_10751);
nor U18331 (N_18331,N_10033,N_13062);
nor U18332 (N_18332,N_10130,N_13179);
nand U18333 (N_18333,N_10458,N_13569);
nand U18334 (N_18334,N_12191,N_11255);
nand U18335 (N_18335,N_14222,N_11617);
nand U18336 (N_18336,N_11356,N_10616);
nor U18337 (N_18337,N_14610,N_12727);
nor U18338 (N_18338,N_12919,N_10587);
xnor U18339 (N_18339,N_11577,N_11301);
xor U18340 (N_18340,N_13309,N_12131);
or U18341 (N_18341,N_12823,N_10884);
xnor U18342 (N_18342,N_11233,N_13581);
xor U18343 (N_18343,N_12212,N_13862);
nand U18344 (N_18344,N_14564,N_13201);
and U18345 (N_18345,N_11417,N_13635);
or U18346 (N_18346,N_13521,N_13552);
and U18347 (N_18347,N_13606,N_13474);
nand U18348 (N_18348,N_12323,N_10146);
xnor U18349 (N_18349,N_12620,N_11649);
nand U18350 (N_18350,N_10622,N_10485);
and U18351 (N_18351,N_14775,N_11957);
nand U18352 (N_18352,N_13432,N_11638);
nand U18353 (N_18353,N_10402,N_13364);
nand U18354 (N_18354,N_14703,N_13446);
nand U18355 (N_18355,N_11171,N_12585);
xor U18356 (N_18356,N_14809,N_12205);
or U18357 (N_18357,N_12868,N_10345);
xor U18358 (N_18358,N_10208,N_12932);
nor U18359 (N_18359,N_13568,N_14535);
xor U18360 (N_18360,N_14450,N_12784);
nand U18361 (N_18361,N_10228,N_14283);
nand U18362 (N_18362,N_10873,N_14638);
nor U18363 (N_18363,N_13877,N_12997);
nor U18364 (N_18364,N_10481,N_13645);
and U18365 (N_18365,N_14905,N_14728);
and U18366 (N_18366,N_12835,N_12861);
or U18367 (N_18367,N_14138,N_10920);
nand U18368 (N_18368,N_11836,N_10916);
nor U18369 (N_18369,N_10608,N_12928);
xor U18370 (N_18370,N_13082,N_14278);
nand U18371 (N_18371,N_11181,N_10420);
or U18372 (N_18372,N_14747,N_12807);
xor U18373 (N_18373,N_11414,N_10387);
nor U18374 (N_18374,N_11986,N_12236);
and U18375 (N_18375,N_11608,N_10449);
nand U18376 (N_18376,N_14567,N_12490);
nor U18377 (N_18377,N_11258,N_10978);
xor U18378 (N_18378,N_10454,N_11915);
nand U18379 (N_18379,N_14199,N_10536);
xnor U18380 (N_18380,N_10799,N_14161);
nor U18381 (N_18381,N_13401,N_12842);
nand U18382 (N_18382,N_10886,N_10275);
nand U18383 (N_18383,N_11261,N_14323);
nor U18384 (N_18384,N_12490,N_12450);
xnor U18385 (N_18385,N_14560,N_13688);
or U18386 (N_18386,N_12619,N_13008);
and U18387 (N_18387,N_10186,N_14615);
nand U18388 (N_18388,N_13706,N_10033);
nand U18389 (N_18389,N_13734,N_11298);
nand U18390 (N_18390,N_11804,N_10677);
or U18391 (N_18391,N_10224,N_11344);
and U18392 (N_18392,N_14789,N_11837);
or U18393 (N_18393,N_14570,N_11399);
or U18394 (N_18394,N_10538,N_11104);
nand U18395 (N_18395,N_13551,N_12501);
or U18396 (N_18396,N_13597,N_10369);
or U18397 (N_18397,N_12280,N_10268);
and U18398 (N_18398,N_12637,N_14870);
xnor U18399 (N_18399,N_11732,N_11276);
nor U18400 (N_18400,N_13764,N_10037);
and U18401 (N_18401,N_11765,N_12014);
nand U18402 (N_18402,N_11919,N_12490);
nor U18403 (N_18403,N_12221,N_13126);
nand U18404 (N_18404,N_10931,N_14470);
or U18405 (N_18405,N_13794,N_13758);
xnor U18406 (N_18406,N_13073,N_14982);
or U18407 (N_18407,N_10347,N_13347);
or U18408 (N_18408,N_11686,N_12888);
or U18409 (N_18409,N_11795,N_13601);
and U18410 (N_18410,N_10314,N_13154);
nor U18411 (N_18411,N_11698,N_12513);
xnor U18412 (N_18412,N_10221,N_14651);
nor U18413 (N_18413,N_11915,N_10375);
xor U18414 (N_18414,N_10058,N_13122);
nand U18415 (N_18415,N_13393,N_14233);
nand U18416 (N_18416,N_14127,N_11912);
nor U18417 (N_18417,N_14389,N_14818);
nor U18418 (N_18418,N_13361,N_10532);
nand U18419 (N_18419,N_13067,N_11050);
and U18420 (N_18420,N_10634,N_12857);
nand U18421 (N_18421,N_14261,N_13321);
xnor U18422 (N_18422,N_13633,N_14712);
xnor U18423 (N_18423,N_10803,N_10147);
and U18424 (N_18424,N_12506,N_13030);
xnor U18425 (N_18425,N_10608,N_14607);
nand U18426 (N_18426,N_10312,N_14392);
nor U18427 (N_18427,N_10559,N_12867);
xor U18428 (N_18428,N_12033,N_11254);
or U18429 (N_18429,N_14274,N_13333);
or U18430 (N_18430,N_13458,N_10932);
xnor U18431 (N_18431,N_14724,N_14764);
xor U18432 (N_18432,N_11923,N_11982);
nor U18433 (N_18433,N_14746,N_12447);
nand U18434 (N_18434,N_14582,N_13567);
nand U18435 (N_18435,N_11711,N_12610);
or U18436 (N_18436,N_14163,N_10596);
xor U18437 (N_18437,N_13976,N_14428);
or U18438 (N_18438,N_14697,N_10467);
and U18439 (N_18439,N_11410,N_14550);
xor U18440 (N_18440,N_12318,N_10053);
nor U18441 (N_18441,N_12067,N_11874);
nor U18442 (N_18442,N_13057,N_11966);
nor U18443 (N_18443,N_11987,N_12310);
xnor U18444 (N_18444,N_10523,N_12322);
or U18445 (N_18445,N_14017,N_10360);
xnor U18446 (N_18446,N_10539,N_10164);
nor U18447 (N_18447,N_12113,N_13870);
xor U18448 (N_18448,N_11468,N_10978);
nor U18449 (N_18449,N_12420,N_11903);
or U18450 (N_18450,N_13213,N_12795);
and U18451 (N_18451,N_13299,N_11748);
nand U18452 (N_18452,N_14508,N_11237);
and U18453 (N_18453,N_11026,N_12335);
nor U18454 (N_18454,N_13244,N_13031);
nor U18455 (N_18455,N_13954,N_13142);
nor U18456 (N_18456,N_14740,N_11827);
nor U18457 (N_18457,N_12904,N_12240);
nor U18458 (N_18458,N_13787,N_11174);
or U18459 (N_18459,N_11197,N_14376);
nand U18460 (N_18460,N_11901,N_12171);
or U18461 (N_18461,N_11841,N_12011);
and U18462 (N_18462,N_13870,N_11138);
or U18463 (N_18463,N_14288,N_13695);
nor U18464 (N_18464,N_14508,N_14278);
and U18465 (N_18465,N_13700,N_14754);
and U18466 (N_18466,N_10459,N_10460);
or U18467 (N_18467,N_11038,N_14756);
nand U18468 (N_18468,N_13733,N_14497);
nor U18469 (N_18469,N_11162,N_12628);
and U18470 (N_18470,N_13721,N_13172);
and U18471 (N_18471,N_14394,N_13742);
nand U18472 (N_18472,N_10365,N_13454);
and U18473 (N_18473,N_13932,N_12695);
nor U18474 (N_18474,N_12258,N_10907);
or U18475 (N_18475,N_13362,N_12147);
and U18476 (N_18476,N_14013,N_12643);
nor U18477 (N_18477,N_11268,N_14108);
xnor U18478 (N_18478,N_12511,N_11768);
and U18479 (N_18479,N_11337,N_12949);
and U18480 (N_18480,N_12577,N_14651);
xnor U18481 (N_18481,N_13905,N_13151);
nand U18482 (N_18482,N_12996,N_13215);
and U18483 (N_18483,N_11352,N_12952);
nand U18484 (N_18484,N_12300,N_10081);
or U18485 (N_18485,N_14408,N_14105);
and U18486 (N_18486,N_14100,N_13705);
nor U18487 (N_18487,N_13821,N_11971);
nor U18488 (N_18488,N_11901,N_12725);
or U18489 (N_18489,N_12663,N_10830);
nor U18490 (N_18490,N_10507,N_14173);
nor U18491 (N_18491,N_11761,N_11312);
nand U18492 (N_18492,N_11488,N_11774);
xor U18493 (N_18493,N_12999,N_13843);
and U18494 (N_18494,N_13902,N_14876);
or U18495 (N_18495,N_11580,N_10864);
xor U18496 (N_18496,N_12803,N_11136);
and U18497 (N_18497,N_12417,N_14830);
xnor U18498 (N_18498,N_14366,N_10960);
xnor U18499 (N_18499,N_11940,N_14902);
and U18500 (N_18500,N_14964,N_13250);
xnor U18501 (N_18501,N_12366,N_14816);
xnor U18502 (N_18502,N_10174,N_14031);
nand U18503 (N_18503,N_12611,N_11043);
nand U18504 (N_18504,N_12533,N_14610);
nor U18505 (N_18505,N_13830,N_14791);
or U18506 (N_18506,N_10471,N_10668);
and U18507 (N_18507,N_10235,N_13922);
and U18508 (N_18508,N_10799,N_12648);
and U18509 (N_18509,N_13797,N_13125);
or U18510 (N_18510,N_13987,N_14002);
nand U18511 (N_18511,N_10064,N_13695);
or U18512 (N_18512,N_12714,N_14480);
or U18513 (N_18513,N_11272,N_14224);
and U18514 (N_18514,N_10512,N_10807);
or U18515 (N_18515,N_10383,N_14415);
xnor U18516 (N_18516,N_11612,N_10288);
and U18517 (N_18517,N_11264,N_13673);
xnor U18518 (N_18518,N_10079,N_12019);
and U18519 (N_18519,N_11441,N_10844);
nand U18520 (N_18520,N_11045,N_11660);
and U18521 (N_18521,N_10617,N_12273);
xor U18522 (N_18522,N_10805,N_12345);
or U18523 (N_18523,N_14545,N_12083);
or U18524 (N_18524,N_13133,N_13834);
xnor U18525 (N_18525,N_14492,N_13122);
xor U18526 (N_18526,N_10300,N_14724);
xor U18527 (N_18527,N_10181,N_12077);
xor U18528 (N_18528,N_10789,N_13953);
or U18529 (N_18529,N_10323,N_13780);
and U18530 (N_18530,N_13790,N_13483);
xnor U18531 (N_18531,N_13165,N_10252);
or U18532 (N_18532,N_13885,N_14618);
nand U18533 (N_18533,N_14638,N_12212);
or U18534 (N_18534,N_11899,N_13653);
or U18535 (N_18535,N_10959,N_10324);
and U18536 (N_18536,N_12318,N_10711);
nand U18537 (N_18537,N_14993,N_14629);
nand U18538 (N_18538,N_13599,N_13417);
nor U18539 (N_18539,N_13486,N_11253);
nand U18540 (N_18540,N_12085,N_12144);
or U18541 (N_18541,N_13469,N_10887);
xor U18542 (N_18542,N_12433,N_10956);
nor U18543 (N_18543,N_10544,N_14918);
nor U18544 (N_18544,N_11128,N_12954);
nand U18545 (N_18545,N_14752,N_13124);
or U18546 (N_18546,N_14619,N_14724);
or U18547 (N_18547,N_11112,N_12834);
nor U18548 (N_18548,N_13855,N_14342);
or U18549 (N_18549,N_12960,N_11317);
xor U18550 (N_18550,N_12130,N_13099);
and U18551 (N_18551,N_14620,N_10174);
or U18552 (N_18552,N_12551,N_11718);
nand U18553 (N_18553,N_10080,N_10611);
and U18554 (N_18554,N_12662,N_14912);
and U18555 (N_18555,N_14591,N_13867);
xnor U18556 (N_18556,N_13603,N_14205);
xor U18557 (N_18557,N_12376,N_13645);
xor U18558 (N_18558,N_10478,N_11232);
and U18559 (N_18559,N_14168,N_11965);
or U18560 (N_18560,N_13603,N_11626);
or U18561 (N_18561,N_11652,N_14900);
nor U18562 (N_18562,N_14228,N_12960);
and U18563 (N_18563,N_10399,N_11583);
or U18564 (N_18564,N_14968,N_10481);
nand U18565 (N_18565,N_10007,N_10423);
or U18566 (N_18566,N_13655,N_14098);
and U18567 (N_18567,N_14071,N_12619);
nor U18568 (N_18568,N_13896,N_11746);
nand U18569 (N_18569,N_11004,N_10953);
nor U18570 (N_18570,N_13233,N_12959);
or U18571 (N_18571,N_13123,N_14582);
or U18572 (N_18572,N_13922,N_14363);
nand U18573 (N_18573,N_10120,N_14796);
xnor U18574 (N_18574,N_14367,N_12619);
nand U18575 (N_18575,N_11692,N_10708);
or U18576 (N_18576,N_13816,N_12186);
nand U18577 (N_18577,N_13394,N_10313);
or U18578 (N_18578,N_12275,N_11801);
xor U18579 (N_18579,N_12849,N_11276);
xor U18580 (N_18580,N_12695,N_13955);
nand U18581 (N_18581,N_14973,N_13395);
xnor U18582 (N_18582,N_10046,N_13990);
nor U18583 (N_18583,N_10372,N_14812);
xnor U18584 (N_18584,N_11640,N_13817);
xor U18585 (N_18585,N_11525,N_13816);
xor U18586 (N_18586,N_10482,N_13775);
nand U18587 (N_18587,N_13669,N_10503);
or U18588 (N_18588,N_14939,N_11069);
nor U18589 (N_18589,N_14452,N_11271);
xor U18590 (N_18590,N_11558,N_12040);
or U18591 (N_18591,N_11662,N_14301);
nor U18592 (N_18592,N_12774,N_11495);
xor U18593 (N_18593,N_10794,N_10162);
and U18594 (N_18594,N_12503,N_12277);
or U18595 (N_18595,N_14173,N_12471);
or U18596 (N_18596,N_14973,N_14336);
nor U18597 (N_18597,N_11550,N_11718);
or U18598 (N_18598,N_14161,N_13036);
nand U18599 (N_18599,N_11715,N_10655);
xor U18600 (N_18600,N_11457,N_11297);
xor U18601 (N_18601,N_12390,N_13871);
nand U18602 (N_18602,N_13784,N_13704);
nor U18603 (N_18603,N_11041,N_10583);
xnor U18604 (N_18604,N_12136,N_10503);
or U18605 (N_18605,N_13559,N_11060);
or U18606 (N_18606,N_13081,N_10519);
or U18607 (N_18607,N_11772,N_10079);
nand U18608 (N_18608,N_10690,N_14427);
and U18609 (N_18609,N_10364,N_11705);
xnor U18610 (N_18610,N_14272,N_12866);
xor U18611 (N_18611,N_12118,N_11271);
nor U18612 (N_18612,N_12370,N_10151);
nand U18613 (N_18613,N_14552,N_11101);
nor U18614 (N_18614,N_13348,N_13624);
and U18615 (N_18615,N_12632,N_14358);
and U18616 (N_18616,N_14030,N_12186);
nor U18617 (N_18617,N_11311,N_14278);
nand U18618 (N_18618,N_11187,N_13292);
nor U18619 (N_18619,N_11174,N_13616);
or U18620 (N_18620,N_10467,N_13380);
nor U18621 (N_18621,N_11669,N_11644);
nor U18622 (N_18622,N_13317,N_13423);
nor U18623 (N_18623,N_14235,N_10396);
nand U18624 (N_18624,N_10923,N_11897);
nand U18625 (N_18625,N_11473,N_13907);
nor U18626 (N_18626,N_11883,N_12235);
and U18627 (N_18627,N_13862,N_13337);
or U18628 (N_18628,N_10420,N_11120);
and U18629 (N_18629,N_12904,N_13582);
or U18630 (N_18630,N_12470,N_10795);
nand U18631 (N_18631,N_10537,N_13340);
or U18632 (N_18632,N_14459,N_10498);
and U18633 (N_18633,N_14133,N_14906);
nand U18634 (N_18634,N_12370,N_11738);
xnor U18635 (N_18635,N_14295,N_10487);
xnor U18636 (N_18636,N_14025,N_10093);
nor U18637 (N_18637,N_12176,N_12375);
or U18638 (N_18638,N_14821,N_14547);
nor U18639 (N_18639,N_14145,N_10142);
and U18640 (N_18640,N_14350,N_14741);
or U18641 (N_18641,N_13502,N_10583);
nor U18642 (N_18642,N_12206,N_10195);
nor U18643 (N_18643,N_10252,N_11787);
or U18644 (N_18644,N_11346,N_10832);
nor U18645 (N_18645,N_13086,N_10354);
and U18646 (N_18646,N_13378,N_12111);
nand U18647 (N_18647,N_11437,N_10673);
or U18648 (N_18648,N_14004,N_14808);
or U18649 (N_18649,N_11856,N_11057);
xnor U18650 (N_18650,N_10559,N_11092);
and U18651 (N_18651,N_12591,N_10384);
xor U18652 (N_18652,N_13536,N_12078);
and U18653 (N_18653,N_14661,N_10998);
or U18654 (N_18654,N_12977,N_14605);
and U18655 (N_18655,N_10249,N_12687);
nor U18656 (N_18656,N_14542,N_14819);
or U18657 (N_18657,N_13637,N_10315);
nor U18658 (N_18658,N_11475,N_14588);
or U18659 (N_18659,N_13605,N_13816);
nor U18660 (N_18660,N_14766,N_11291);
nor U18661 (N_18661,N_12168,N_12831);
nand U18662 (N_18662,N_11008,N_13828);
xor U18663 (N_18663,N_14655,N_13154);
nor U18664 (N_18664,N_13170,N_13781);
nand U18665 (N_18665,N_14142,N_12861);
nand U18666 (N_18666,N_14007,N_14731);
nor U18667 (N_18667,N_10594,N_12966);
nand U18668 (N_18668,N_14602,N_13169);
nor U18669 (N_18669,N_13890,N_11053);
nand U18670 (N_18670,N_14566,N_12453);
or U18671 (N_18671,N_14556,N_12729);
or U18672 (N_18672,N_14187,N_10827);
and U18673 (N_18673,N_14583,N_10471);
or U18674 (N_18674,N_11018,N_13441);
or U18675 (N_18675,N_14296,N_10817);
or U18676 (N_18676,N_13661,N_11290);
nand U18677 (N_18677,N_10853,N_11541);
xnor U18678 (N_18678,N_10135,N_13607);
and U18679 (N_18679,N_10138,N_14973);
or U18680 (N_18680,N_13752,N_11867);
or U18681 (N_18681,N_12674,N_13045);
xnor U18682 (N_18682,N_10518,N_10384);
xor U18683 (N_18683,N_10522,N_14817);
nor U18684 (N_18684,N_11424,N_13717);
nor U18685 (N_18685,N_12424,N_14636);
nor U18686 (N_18686,N_11494,N_11878);
nor U18687 (N_18687,N_11833,N_11234);
or U18688 (N_18688,N_14222,N_14397);
or U18689 (N_18689,N_12082,N_11006);
nand U18690 (N_18690,N_10290,N_12491);
xor U18691 (N_18691,N_10903,N_10769);
nor U18692 (N_18692,N_12576,N_11517);
nor U18693 (N_18693,N_11952,N_12611);
and U18694 (N_18694,N_13181,N_10154);
or U18695 (N_18695,N_10714,N_12886);
or U18696 (N_18696,N_12803,N_14757);
nand U18697 (N_18697,N_14935,N_13785);
and U18698 (N_18698,N_10110,N_14447);
or U18699 (N_18699,N_14315,N_14113);
nand U18700 (N_18700,N_14156,N_10877);
nand U18701 (N_18701,N_14584,N_12538);
or U18702 (N_18702,N_12849,N_12083);
or U18703 (N_18703,N_11541,N_14392);
or U18704 (N_18704,N_10710,N_14768);
or U18705 (N_18705,N_13983,N_14204);
and U18706 (N_18706,N_10243,N_14767);
or U18707 (N_18707,N_11909,N_10276);
xor U18708 (N_18708,N_11061,N_10366);
nand U18709 (N_18709,N_10293,N_13490);
xnor U18710 (N_18710,N_14940,N_13756);
nand U18711 (N_18711,N_12242,N_14677);
and U18712 (N_18712,N_12625,N_12011);
and U18713 (N_18713,N_13153,N_14812);
nor U18714 (N_18714,N_11121,N_11565);
xnor U18715 (N_18715,N_10108,N_14907);
nand U18716 (N_18716,N_13845,N_12364);
nor U18717 (N_18717,N_10201,N_12224);
nor U18718 (N_18718,N_13209,N_11398);
xnor U18719 (N_18719,N_10146,N_10460);
or U18720 (N_18720,N_13436,N_13825);
and U18721 (N_18721,N_14120,N_13810);
nor U18722 (N_18722,N_14458,N_13419);
and U18723 (N_18723,N_12682,N_12845);
and U18724 (N_18724,N_11098,N_13299);
nand U18725 (N_18725,N_13815,N_12361);
nor U18726 (N_18726,N_12792,N_12244);
xnor U18727 (N_18727,N_10568,N_10950);
nor U18728 (N_18728,N_14056,N_10805);
xor U18729 (N_18729,N_13655,N_13629);
nor U18730 (N_18730,N_14805,N_10379);
nor U18731 (N_18731,N_13445,N_14247);
xor U18732 (N_18732,N_11428,N_11372);
nor U18733 (N_18733,N_10650,N_12857);
or U18734 (N_18734,N_14524,N_13239);
xnor U18735 (N_18735,N_11987,N_12162);
and U18736 (N_18736,N_13213,N_13456);
or U18737 (N_18737,N_13890,N_10161);
or U18738 (N_18738,N_10584,N_14557);
nand U18739 (N_18739,N_14865,N_10014);
and U18740 (N_18740,N_13063,N_12977);
and U18741 (N_18741,N_14314,N_14016);
and U18742 (N_18742,N_11587,N_12453);
xor U18743 (N_18743,N_12516,N_11982);
nand U18744 (N_18744,N_14846,N_13995);
nor U18745 (N_18745,N_11524,N_14652);
nor U18746 (N_18746,N_13075,N_13632);
and U18747 (N_18747,N_12665,N_12957);
nor U18748 (N_18748,N_11540,N_12171);
nand U18749 (N_18749,N_12301,N_13480);
nor U18750 (N_18750,N_11166,N_12200);
nand U18751 (N_18751,N_13757,N_11781);
nand U18752 (N_18752,N_14911,N_12068);
nand U18753 (N_18753,N_12726,N_13405);
xor U18754 (N_18754,N_13911,N_10154);
xnor U18755 (N_18755,N_10549,N_11323);
nand U18756 (N_18756,N_12089,N_11124);
nor U18757 (N_18757,N_11866,N_10957);
or U18758 (N_18758,N_14362,N_10565);
nand U18759 (N_18759,N_12101,N_14887);
xor U18760 (N_18760,N_11969,N_14910);
nand U18761 (N_18761,N_12359,N_12768);
and U18762 (N_18762,N_14696,N_13356);
xnor U18763 (N_18763,N_10127,N_12639);
and U18764 (N_18764,N_14193,N_13920);
nand U18765 (N_18765,N_14768,N_14397);
nor U18766 (N_18766,N_14892,N_10006);
xnor U18767 (N_18767,N_11356,N_12049);
nand U18768 (N_18768,N_14028,N_11952);
xnor U18769 (N_18769,N_10763,N_14204);
and U18770 (N_18770,N_10946,N_10835);
or U18771 (N_18771,N_11721,N_14201);
nor U18772 (N_18772,N_14237,N_14759);
and U18773 (N_18773,N_11443,N_12406);
or U18774 (N_18774,N_13788,N_12051);
nand U18775 (N_18775,N_12762,N_12526);
nand U18776 (N_18776,N_10307,N_11245);
and U18777 (N_18777,N_13728,N_10437);
xnor U18778 (N_18778,N_12366,N_11401);
and U18779 (N_18779,N_14888,N_14444);
or U18780 (N_18780,N_10099,N_14558);
or U18781 (N_18781,N_11766,N_11476);
xnor U18782 (N_18782,N_13761,N_12757);
nor U18783 (N_18783,N_10673,N_12651);
xor U18784 (N_18784,N_11020,N_10826);
xor U18785 (N_18785,N_11274,N_13263);
nand U18786 (N_18786,N_11426,N_10518);
or U18787 (N_18787,N_10420,N_11191);
nand U18788 (N_18788,N_12333,N_14157);
or U18789 (N_18789,N_11554,N_10839);
nand U18790 (N_18790,N_13019,N_13707);
or U18791 (N_18791,N_14615,N_12135);
nand U18792 (N_18792,N_14598,N_10329);
or U18793 (N_18793,N_14852,N_13469);
or U18794 (N_18794,N_10170,N_10231);
or U18795 (N_18795,N_11918,N_14770);
nand U18796 (N_18796,N_12061,N_12794);
or U18797 (N_18797,N_11360,N_10174);
nor U18798 (N_18798,N_12998,N_14820);
or U18799 (N_18799,N_10092,N_13460);
xnor U18800 (N_18800,N_10033,N_11029);
or U18801 (N_18801,N_11017,N_12036);
xor U18802 (N_18802,N_13558,N_14021);
and U18803 (N_18803,N_11230,N_12542);
nor U18804 (N_18804,N_11326,N_11559);
nor U18805 (N_18805,N_11461,N_12903);
nand U18806 (N_18806,N_13361,N_10758);
or U18807 (N_18807,N_12596,N_14573);
nand U18808 (N_18808,N_10980,N_14540);
nand U18809 (N_18809,N_11497,N_11433);
xnor U18810 (N_18810,N_10119,N_11381);
xor U18811 (N_18811,N_12026,N_12060);
nor U18812 (N_18812,N_12861,N_11526);
nor U18813 (N_18813,N_13424,N_11931);
nor U18814 (N_18814,N_12507,N_11047);
xnor U18815 (N_18815,N_11055,N_14906);
and U18816 (N_18816,N_10857,N_14262);
or U18817 (N_18817,N_12938,N_11982);
nand U18818 (N_18818,N_10241,N_12838);
xor U18819 (N_18819,N_13344,N_13478);
or U18820 (N_18820,N_14462,N_10708);
xor U18821 (N_18821,N_13782,N_12090);
and U18822 (N_18822,N_14585,N_14182);
nand U18823 (N_18823,N_11678,N_14051);
and U18824 (N_18824,N_14657,N_11164);
xor U18825 (N_18825,N_12203,N_14420);
nand U18826 (N_18826,N_11441,N_14231);
nor U18827 (N_18827,N_13428,N_13543);
nand U18828 (N_18828,N_12428,N_14562);
or U18829 (N_18829,N_14997,N_11620);
xor U18830 (N_18830,N_13165,N_14887);
nand U18831 (N_18831,N_13233,N_12400);
xnor U18832 (N_18832,N_13751,N_10625);
and U18833 (N_18833,N_10097,N_12564);
and U18834 (N_18834,N_14487,N_13744);
xnor U18835 (N_18835,N_14979,N_12645);
or U18836 (N_18836,N_14077,N_11226);
nand U18837 (N_18837,N_11691,N_14153);
xnor U18838 (N_18838,N_14336,N_14740);
and U18839 (N_18839,N_14914,N_14777);
xor U18840 (N_18840,N_14315,N_10046);
xor U18841 (N_18841,N_10404,N_11255);
and U18842 (N_18842,N_12952,N_11129);
nand U18843 (N_18843,N_10979,N_10660);
or U18844 (N_18844,N_12573,N_14844);
or U18845 (N_18845,N_14546,N_11334);
xor U18846 (N_18846,N_14026,N_13144);
nand U18847 (N_18847,N_14109,N_12707);
and U18848 (N_18848,N_11134,N_13872);
and U18849 (N_18849,N_13689,N_10431);
xnor U18850 (N_18850,N_11948,N_13035);
nand U18851 (N_18851,N_12021,N_13007);
nor U18852 (N_18852,N_10048,N_12938);
nand U18853 (N_18853,N_14187,N_11416);
nand U18854 (N_18854,N_14322,N_10581);
nor U18855 (N_18855,N_13166,N_13630);
nand U18856 (N_18856,N_13021,N_12893);
xor U18857 (N_18857,N_10176,N_13627);
nor U18858 (N_18858,N_10823,N_13265);
xnor U18859 (N_18859,N_14158,N_10405);
and U18860 (N_18860,N_11520,N_10907);
or U18861 (N_18861,N_13087,N_14906);
or U18862 (N_18862,N_13025,N_14781);
nor U18863 (N_18863,N_10947,N_12755);
and U18864 (N_18864,N_13346,N_14793);
or U18865 (N_18865,N_12045,N_12160);
and U18866 (N_18866,N_10076,N_12826);
or U18867 (N_18867,N_11599,N_13491);
or U18868 (N_18868,N_12281,N_11171);
nand U18869 (N_18869,N_12266,N_11207);
or U18870 (N_18870,N_14910,N_10085);
nor U18871 (N_18871,N_14326,N_14395);
and U18872 (N_18872,N_14824,N_12641);
nand U18873 (N_18873,N_14713,N_12858);
nand U18874 (N_18874,N_14914,N_11217);
and U18875 (N_18875,N_13343,N_13280);
xor U18876 (N_18876,N_13624,N_10607);
or U18877 (N_18877,N_12782,N_12319);
nand U18878 (N_18878,N_14582,N_10359);
or U18879 (N_18879,N_14256,N_13652);
and U18880 (N_18880,N_10796,N_11440);
nand U18881 (N_18881,N_14936,N_12265);
xor U18882 (N_18882,N_13062,N_10220);
nand U18883 (N_18883,N_14878,N_14536);
nor U18884 (N_18884,N_12968,N_10852);
or U18885 (N_18885,N_12059,N_11809);
xnor U18886 (N_18886,N_11942,N_14890);
xor U18887 (N_18887,N_14193,N_13278);
nor U18888 (N_18888,N_13508,N_10608);
xor U18889 (N_18889,N_12573,N_11396);
xor U18890 (N_18890,N_13016,N_11456);
and U18891 (N_18891,N_14043,N_10623);
nor U18892 (N_18892,N_12852,N_12952);
and U18893 (N_18893,N_13278,N_12686);
or U18894 (N_18894,N_12564,N_10942);
xnor U18895 (N_18895,N_12969,N_13025);
xnor U18896 (N_18896,N_13737,N_13453);
or U18897 (N_18897,N_14080,N_10508);
and U18898 (N_18898,N_10688,N_10896);
or U18899 (N_18899,N_11232,N_12717);
nand U18900 (N_18900,N_11012,N_11342);
and U18901 (N_18901,N_13114,N_12783);
nor U18902 (N_18902,N_12655,N_11336);
and U18903 (N_18903,N_12689,N_14529);
xor U18904 (N_18904,N_14946,N_13971);
nand U18905 (N_18905,N_12081,N_14095);
nand U18906 (N_18906,N_14237,N_13479);
and U18907 (N_18907,N_10074,N_10198);
or U18908 (N_18908,N_11568,N_11397);
nor U18909 (N_18909,N_11336,N_10594);
and U18910 (N_18910,N_12967,N_12644);
nand U18911 (N_18911,N_14403,N_10176);
nor U18912 (N_18912,N_10181,N_12775);
nand U18913 (N_18913,N_13686,N_11189);
and U18914 (N_18914,N_14057,N_14897);
nand U18915 (N_18915,N_10481,N_12464);
or U18916 (N_18916,N_13151,N_14995);
nand U18917 (N_18917,N_13819,N_10651);
xor U18918 (N_18918,N_12987,N_14460);
xor U18919 (N_18919,N_14850,N_12680);
or U18920 (N_18920,N_14387,N_13779);
nand U18921 (N_18921,N_12855,N_10882);
xnor U18922 (N_18922,N_11985,N_13496);
xor U18923 (N_18923,N_11054,N_13747);
xor U18924 (N_18924,N_11844,N_11981);
nand U18925 (N_18925,N_10628,N_12509);
xnor U18926 (N_18926,N_10810,N_13496);
nand U18927 (N_18927,N_12844,N_14788);
xnor U18928 (N_18928,N_11393,N_12677);
and U18929 (N_18929,N_10544,N_13550);
xor U18930 (N_18930,N_10334,N_12558);
xor U18931 (N_18931,N_14686,N_13354);
and U18932 (N_18932,N_10425,N_12611);
or U18933 (N_18933,N_10305,N_13559);
nand U18934 (N_18934,N_14147,N_14108);
xor U18935 (N_18935,N_12678,N_11234);
nor U18936 (N_18936,N_13145,N_12035);
and U18937 (N_18937,N_10108,N_14410);
or U18938 (N_18938,N_11045,N_13383);
nor U18939 (N_18939,N_13567,N_13808);
xor U18940 (N_18940,N_12056,N_14260);
nor U18941 (N_18941,N_10998,N_14858);
or U18942 (N_18942,N_14512,N_10440);
nand U18943 (N_18943,N_14933,N_13812);
and U18944 (N_18944,N_14904,N_11033);
and U18945 (N_18945,N_11524,N_10270);
nand U18946 (N_18946,N_13397,N_11267);
xnor U18947 (N_18947,N_13407,N_11251);
or U18948 (N_18948,N_12579,N_10368);
nor U18949 (N_18949,N_11454,N_14014);
or U18950 (N_18950,N_10927,N_13495);
or U18951 (N_18951,N_11491,N_11555);
nor U18952 (N_18952,N_10711,N_13091);
and U18953 (N_18953,N_13993,N_10866);
nand U18954 (N_18954,N_14158,N_12104);
nor U18955 (N_18955,N_12429,N_12222);
xor U18956 (N_18956,N_14942,N_11598);
xnor U18957 (N_18957,N_11215,N_14452);
nor U18958 (N_18958,N_10292,N_12663);
and U18959 (N_18959,N_14962,N_12194);
or U18960 (N_18960,N_10583,N_10507);
or U18961 (N_18961,N_13941,N_13308);
nand U18962 (N_18962,N_11438,N_11753);
nand U18963 (N_18963,N_13312,N_11544);
or U18964 (N_18964,N_14924,N_13640);
nand U18965 (N_18965,N_14458,N_13352);
and U18966 (N_18966,N_11170,N_11514);
nand U18967 (N_18967,N_12937,N_12784);
and U18968 (N_18968,N_12923,N_13237);
nor U18969 (N_18969,N_12802,N_11042);
xor U18970 (N_18970,N_10085,N_11915);
or U18971 (N_18971,N_13544,N_12325);
xnor U18972 (N_18972,N_11347,N_13015);
or U18973 (N_18973,N_12047,N_10920);
and U18974 (N_18974,N_10453,N_13044);
nor U18975 (N_18975,N_14303,N_12761);
and U18976 (N_18976,N_13130,N_10028);
nor U18977 (N_18977,N_12640,N_12475);
and U18978 (N_18978,N_14938,N_14843);
xor U18979 (N_18979,N_14409,N_11267);
xor U18980 (N_18980,N_10150,N_14219);
nand U18981 (N_18981,N_10101,N_12550);
nor U18982 (N_18982,N_11520,N_11642);
nor U18983 (N_18983,N_10019,N_13949);
nor U18984 (N_18984,N_11000,N_14079);
nor U18985 (N_18985,N_14224,N_14878);
and U18986 (N_18986,N_13247,N_11114);
and U18987 (N_18987,N_13044,N_10968);
nand U18988 (N_18988,N_10013,N_10651);
and U18989 (N_18989,N_12669,N_13105);
xor U18990 (N_18990,N_12216,N_13273);
and U18991 (N_18991,N_10543,N_13929);
xor U18992 (N_18992,N_14643,N_10418);
or U18993 (N_18993,N_14992,N_12716);
nand U18994 (N_18994,N_10125,N_12149);
nand U18995 (N_18995,N_11107,N_13405);
and U18996 (N_18996,N_13623,N_14883);
and U18997 (N_18997,N_14030,N_13178);
nor U18998 (N_18998,N_13488,N_14483);
or U18999 (N_18999,N_13878,N_13673);
or U19000 (N_19000,N_13019,N_11877);
xor U19001 (N_19001,N_12597,N_14008);
or U19002 (N_19002,N_11508,N_11094);
xor U19003 (N_19003,N_13665,N_13911);
nand U19004 (N_19004,N_11529,N_14176);
xnor U19005 (N_19005,N_13824,N_13254);
nand U19006 (N_19006,N_14738,N_11664);
or U19007 (N_19007,N_13050,N_13029);
nand U19008 (N_19008,N_12185,N_13691);
or U19009 (N_19009,N_13383,N_13765);
xnor U19010 (N_19010,N_13955,N_14966);
or U19011 (N_19011,N_11263,N_13537);
nand U19012 (N_19012,N_13068,N_12330);
or U19013 (N_19013,N_14421,N_13806);
nor U19014 (N_19014,N_10575,N_14627);
and U19015 (N_19015,N_11777,N_10960);
xor U19016 (N_19016,N_13019,N_12080);
nor U19017 (N_19017,N_14483,N_13975);
xor U19018 (N_19018,N_13851,N_12442);
nand U19019 (N_19019,N_14594,N_10958);
xnor U19020 (N_19020,N_12714,N_10426);
nor U19021 (N_19021,N_12922,N_12545);
and U19022 (N_19022,N_11294,N_13557);
and U19023 (N_19023,N_10668,N_10184);
nor U19024 (N_19024,N_12832,N_12006);
xnor U19025 (N_19025,N_14099,N_12699);
xor U19026 (N_19026,N_13344,N_10969);
and U19027 (N_19027,N_14538,N_13197);
nor U19028 (N_19028,N_13722,N_14965);
nand U19029 (N_19029,N_13553,N_11641);
and U19030 (N_19030,N_13968,N_10750);
nand U19031 (N_19031,N_12248,N_12654);
nand U19032 (N_19032,N_10862,N_10804);
and U19033 (N_19033,N_11723,N_13936);
and U19034 (N_19034,N_11347,N_10261);
and U19035 (N_19035,N_10377,N_12423);
nor U19036 (N_19036,N_14599,N_12233);
or U19037 (N_19037,N_13151,N_11740);
or U19038 (N_19038,N_14686,N_12239);
or U19039 (N_19039,N_11438,N_11974);
nand U19040 (N_19040,N_12408,N_12283);
nor U19041 (N_19041,N_10578,N_11475);
or U19042 (N_19042,N_14094,N_10027);
nand U19043 (N_19043,N_14672,N_10284);
or U19044 (N_19044,N_13066,N_11600);
xnor U19045 (N_19045,N_13926,N_14768);
nand U19046 (N_19046,N_13675,N_14743);
or U19047 (N_19047,N_10360,N_10901);
nand U19048 (N_19048,N_10058,N_14742);
and U19049 (N_19049,N_11261,N_11816);
or U19050 (N_19050,N_12819,N_11771);
nor U19051 (N_19051,N_10936,N_12591);
nor U19052 (N_19052,N_10169,N_14333);
xnor U19053 (N_19053,N_11026,N_12155);
or U19054 (N_19054,N_13302,N_12268);
nand U19055 (N_19055,N_12720,N_13239);
nand U19056 (N_19056,N_10406,N_12944);
and U19057 (N_19057,N_11768,N_10851);
or U19058 (N_19058,N_10444,N_14385);
or U19059 (N_19059,N_11865,N_13461);
or U19060 (N_19060,N_12196,N_13925);
nand U19061 (N_19061,N_10406,N_14010);
or U19062 (N_19062,N_13386,N_11101);
nor U19063 (N_19063,N_14040,N_14529);
nor U19064 (N_19064,N_10432,N_10484);
xor U19065 (N_19065,N_13795,N_14030);
nor U19066 (N_19066,N_11489,N_11865);
nand U19067 (N_19067,N_14453,N_13149);
nor U19068 (N_19068,N_14361,N_10509);
nand U19069 (N_19069,N_14027,N_10234);
nor U19070 (N_19070,N_12234,N_13941);
and U19071 (N_19071,N_12957,N_13057);
or U19072 (N_19072,N_12071,N_14370);
and U19073 (N_19073,N_12949,N_12675);
xnor U19074 (N_19074,N_12925,N_10441);
or U19075 (N_19075,N_12097,N_13182);
nand U19076 (N_19076,N_14374,N_13636);
nor U19077 (N_19077,N_11473,N_13293);
or U19078 (N_19078,N_10459,N_14328);
or U19079 (N_19079,N_14893,N_13998);
and U19080 (N_19080,N_12023,N_11688);
or U19081 (N_19081,N_14463,N_10903);
xor U19082 (N_19082,N_10079,N_13796);
nor U19083 (N_19083,N_11942,N_13276);
nor U19084 (N_19084,N_10028,N_14050);
and U19085 (N_19085,N_11148,N_10960);
and U19086 (N_19086,N_14447,N_10713);
xor U19087 (N_19087,N_12760,N_14807);
nor U19088 (N_19088,N_13198,N_13303);
xor U19089 (N_19089,N_13756,N_14917);
nand U19090 (N_19090,N_11431,N_12250);
xor U19091 (N_19091,N_14561,N_12901);
and U19092 (N_19092,N_11196,N_10504);
nand U19093 (N_19093,N_10086,N_14337);
or U19094 (N_19094,N_13039,N_14974);
and U19095 (N_19095,N_14911,N_12399);
xnor U19096 (N_19096,N_11997,N_11822);
nor U19097 (N_19097,N_11173,N_14478);
nand U19098 (N_19098,N_10115,N_11877);
or U19099 (N_19099,N_12392,N_13001);
nor U19100 (N_19100,N_14382,N_11105);
or U19101 (N_19101,N_12789,N_10461);
or U19102 (N_19102,N_11032,N_11502);
and U19103 (N_19103,N_12014,N_12100);
and U19104 (N_19104,N_14969,N_13668);
nand U19105 (N_19105,N_12977,N_12862);
and U19106 (N_19106,N_11195,N_14322);
nand U19107 (N_19107,N_13971,N_11180);
or U19108 (N_19108,N_12887,N_10297);
nor U19109 (N_19109,N_11877,N_14621);
nor U19110 (N_19110,N_12283,N_11404);
xor U19111 (N_19111,N_10226,N_13051);
or U19112 (N_19112,N_14852,N_12122);
nand U19113 (N_19113,N_14958,N_14231);
xnor U19114 (N_19114,N_11880,N_13169);
and U19115 (N_19115,N_10060,N_12248);
or U19116 (N_19116,N_11652,N_10979);
or U19117 (N_19117,N_11625,N_12604);
and U19118 (N_19118,N_13061,N_14791);
nand U19119 (N_19119,N_10060,N_11366);
and U19120 (N_19120,N_13956,N_13888);
nand U19121 (N_19121,N_12757,N_13429);
or U19122 (N_19122,N_14158,N_10087);
and U19123 (N_19123,N_14340,N_10235);
xnor U19124 (N_19124,N_12229,N_10555);
nor U19125 (N_19125,N_14051,N_12516);
and U19126 (N_19126,N_12867,N_14277);
nor U19127 (N_19127,N_12465,N_14579);
or U19128 (N_19128,N_13059,N_14486);
nor U19129 (N_19129,N_12724,N_13975);
nand U19130 (N_19130,N_14667,N_13128);
or U19131 (N_19131,N_10190,N_13027);
nor U19132 (N_19132,N_11297,N_13982);
or U19133 (N_19133,N_10118,N_13615);
nor U19134 (N_19134,N_14715,N_13896);
nand U19135 (N_19135,N_12155,N_12328);
nand U19136 (N_19136,N_13655,N_14966);
and U19137 (N_19137,N_12133,N_10400);
xnor U19138 (N_19138,N_14383,N_10749);
nor U19139 (N_19139,N_13847,N_11997);
or U19140 (N_19140,N_12177,N_12680);
or U19141 (N_19141,N_13924,N_14307);
xnor U19142 (N_19142,N_12976,N_13667);
xor U19143 (N_19143,N_10791,N_12889);
xnor U19144 (N_19144,N_11560,N_14188);
nor U19145 (N_19145,N_13180,N_10402);
and U19146 (N_19146,N_10576,N_14433);
xnor U19147 (N_19147,N_10536,N_11386);
nand U19148 (N_19148,N_14561,N_13413);
and U19149 (N_19149,N_13319,N_13050);
xnor U19150 (N_19150,N_13019,N_11250);
and U19151 (N_19151,N_13840,N_13312);
or U19152 (N_19152,N_11215,N_11910);
nand U19153 (N_19153,N_12239,N_10487);
nor U19154 (N_19154,N_14389,N_11878);
or U19155 (N_19155,N_13270,N_14201);
or U19156 (N_19156,N_14564,N_11197);
nor U19157 (N_19157,N_11569,N_11591);
nor U19158 (N_19158,N_13310,N_10742);
nor U19159 (N_19159,N_13947,N_13899);
nor U19160 (N_19160,N_13230,N_13410);
xor U19161 (N_19161,N_10030,N_13042);
xor U19162 (N_19162,N_14321,N_14723);
nand U19163 (N_19163,N_13247,N_14846);
nand U19164 (N_19164,N_12229,N_14032);
xor U19165 (N_19165,N_12452,N_13885);
xnor U19166 (N_19166,N_13774,N_11983);
and U19167 (N_19167,N_14753,N_12154);
and U19168 (N_19168,N_14179,N_13794);
or U19169 (N_19169,N_13379,N_10775);
and U19170 (N_19170,N_12457,N_14605);
or U19171 (N_19171,N_12175,N_12300);
xor U19172 (N_19172,N_12848,N_14193);
nand U19173 (N_19173,N_14232,N_11420);
nand U19174 (N_19174,N_13299,N_13497);
nand U19175 (N_19175,N_10933,N_14926);
and U19176 (N_19176,N_11816,N_14278);
nor U19177 (N_19177,N_12345,N_11077);
or U19178 (N_19178,N_12397,N_10790);
nand U19179 (N_19179,N_14194,N_13595);
and U19180 (N_19180,N_10730,N_14844);
nand U19181 (N_19181,N_11053,N_14045);
nor U19182 (N_19182,N_12641,N_13304);
or U19183 (N_19183,N_13056,N_13362);
and U19184 (N_19184,N_14427,N_13116);
or U19185 (N_19185,N_12237,N_10243);
xnor U19186 (N_19186,N_14288,N_14244);
xor U19187 (N_19187,N_12568,N_11510);
and U19188 (N_19188,N_10815,N_10864);
or U19189 (N_19189,N_10932,N_11842);
or U19190 (N_19190,N_10757,N_14178);
or U19191 (N_19191,N_12685,N_13491);
or U19192 (N_19192,N_11826,N_10559);
or U19193 (N_19193,N_11374,N_10209);
and U19194 (N_19194,N_14649,N_10464);
nor U19195 (N_19195,N_13476,N_11010);
or U19196 (N_19196,N_12547,N_11738);
nor U19197 (N_19197,N_10070,N_14095);
nor U19198 (N_19198,N_10451,N_13204);
xnor U19199 (N_19199,N_13760,N_14830);
nor U19200 (N_19200,N_14481,N_10642);
and U19201 (N_19201,N_10570,N_11617);
and U19202 (N_19202,N_11034,N_13458);
nor U19203 (N_19203,N_11043,N_13843);
xnor U19204 (N_19204,N_13280,N_10367);
or U19205 (N_19205,N_13211,N_12488);
or U19206 (N_19206,N_11098,N_10257);
and U19207 (N_19207,N_11849,N_11216);
and U19208 (N_19208,N_12619,N_12630);
and U19209 (N_19209,N_10749,N_13903);
xor U19210 (N_19210,N_11764,N_10818);
nand U19211 (N_19211,N_11602,N_12642);
xnor U19212 (N_19212,N_12854,N_12846);
nand U19213 (N_19213,N_13592,N_13761);
xnor U19214 (N_19214,N_13156,N_14861);
nor U19215 (N_19215,N_13779,N_11619);
nor U19216 (N_19216,N_10771,N_11585);
xor U19217 (N_19217,N_13292,N_13475);
nand U19218 (N_19218,N_14371,N_14141);
xnor U19219 (N_19219,N_12042,N_14376);
xnor U19220 (N_19220,N_11521,N_12426);
or U19221 (N_19221,N_12190,N_12945);
nor U19222 (N_19222,N_13174,N_12349);
xnor U19223 (N_19223,N_11192,N_12824);
xnor U19224 (N_19224,N_14312,N_11474);
and U19225 (N_19225,N_12958,N_10474);
xor U19226 (N_19226,N_10398,N_14236);
and U19227 (N_19227,N_11714,N_14079);
and U19228 (N_19228,N_10495,N_12356);
nand U19229 (N_19229,N_12343,N_12738);
nor U19230 (N_19230,N_12140,N_14933);
nand U19231 (N_19231,N_12921,N_10827);
nand U19232 (N_19232,N_12044,N_14407);
nor U19233 (N_19233,N_14171,N_14299);
and U19234 (N_19234,N_14952,N_10495);
xnor U19235 (N_19235,N_14711,N_10579);
nand U19236 (N_19236,N_13493,N_10040);
and U19237 (N_19237,N_13593,N_10174);
xnor U19238 (N_19238,N_10429,N_10530);
or U19239 (N_19239,N_10057,N_12436);
nand U19240 (N_19240,N_12774,N_12804);
or U19241 (N_19241,N_12045,N_11994);
xnor U19242 (N_19242,N_13326,N_13806);
xnor U19243 (N_19243,N_10786,N_10629);
xnor U19244 (N_19244,N_11935,N_13483);
or U19245 (N_19245,N_13076,N_13803);
nor U19246 (N_19246,N_13506,N_11879);
nand U19247 (N_19247,N_13628,N_11969);
nand U19248 (N_19248,N_13340,N_13783);
and U19249 (N_19249,N_13257,N_13034);
xor U19250 (N_19250,N_10571,N_13158);
and U19251 (N_19251,N_12425,N_11643);
xnor U19252 (N_19252,N_10994,N_12903);
nand U19253 (N_19253,N_12469,N_13010);
and U19254 (N_19254,N_10779,N_11403);
xnor U19255 (N_19255,N_11221,N_10257);
and U19256 (N_19256,N_10815,N_11779);
or U19257 (N_19257,N_14959,N_13983);
xor U19258 (N_19258,N_12998,N_14596);
nor U19259 (N_19259,N_11796,N_14086);
nor U19260 (N_19260,N_10643,N_11733);
nand U19261 (N_19261,N_10721,N_12500);
nand U19262 (N_19262,N_13314,N_14972);
and U19263 (N_19263,N_10935,N_10006);
or U19264 (N_19264,N_14519,N_14182);
xnor U19265 (N_19265,N_10935,N_13006);
xor U19266 (N_19266,N_11329,N_14658);
xnor U19267 (N_19267,N_11969,N_10325);
and U19268 (N_19268,N_12729,N_13475);
xnor U19269 (N_19269,N_14842,N_13472);
nor U19270 (N_19270,N_12197,N_10202);
nor U19271 (N_19271,N_13949,N_11019);
xor U19272 (N_19272,N_14567,N_12376);
or U19273 (N_19273,N_10620,N_11042);
nor U19274 (N_19274,N_12185,N_12108);
and U19275 (N_19275,N_13108,N_10319);
nand U19276 (N_19276,N_10025,N_12537);
or U19277 (N_19277,N_13497,N_10218);
nand U19278 (N_19278,N_14992,N_12355);
nor U19279 (N_19279,N_11265,N_14887);
or U19280 (N_19280,N_13723,N_11823);
xnor U19281 (N_19281,N_12282,N_10244);
and U19282 (N_19282,N_14997,N_14182);
xor U19283 (N_19283,N_11540,N_11961);
nor U19284 (N_19284,N_11541,N_14579);
and U19285 (N_19285,N_13372,N_12870);
and U19286 (N_19286,N_12412,N_13262);
and U19287 (N_19287,N_10682,N_12033);
nand U19288 (N_19288,N_11043,N_14578);
nor U19289 (N_19289,N_14284,N_11005);
nand U19290 (N_19290,N_11361,N_14292);
nor U19291 (N_19291,N_14298,N_12314);
or U19292 (N_19292,N_11331,N_11043);
and U19293 (N_19293,N_14850,N_12600);
xnor U19294 (N_19294,N_11971,N_14870);
nor U19295 (N_19295,N_10569,N_13640);
and U19296 (N_19296,N_11138,N_14035);
nand U19297 (N_19297,N_13576,N_13918);
nand U19298 (N_19298,N_11102,N_13181);
and U19299 (N_19299,N_12991,N_11936);
or U19300 (N_19300,N_11165,N_13119);
nor U19301 (N_19301,N_11820,N_13888);
and U19302 (N_19302,N_11081,N_12136);
or U19303 (N_19303,N_14921,N_11409);
nand U19304 (N_19304,N_11051,N_11006);
xnor U19305 (N_19305,N_10702,N_10009);
nand U19306 (N_19306,N_10659,N_14365);
nand U19307 (N_19307,N_14903,N_11509);
nand U19308 (N_19308,N_12730,N_12748);
or U19309 (N_19309,N_12386,N_13724);
xor U19310 (N_19310,N_12374,N_11632);
and U19311 (N_19311,N_10037,N_13247);
or U19312 (N_19312,N_14247,N_14579);
nand U19313 (N_19313,N_10476,N_14380);
and U19314 (N_19314,N_11552,N_14486);
xnor U19315 (N_19315,N_11247,N_11789);
or U19316 (N_19316,N_10763,N_10668);
nor U19317 (N_19317,N_10736,N_11361);
and U19318 (N_19318,N_11669,N_12100);
and U19319 (N_19319,N_11904,N_13549);
xnor U19320 (N_19320,N_10935,N_10645);
and U19321 (N_19321,N_11666,N_12241);
nor U19322 (N_19322,N_13240,N_12432);
nand U19323 (N_19323,N_11345,N_10846);
or U19324 (N_19324,N_13857,N_11852);
or U19325 (N_19325,N_10891,N_14385);
nor U19326 (N_19326,N_13651,N_14574);
and U19327 (N_19327,N_11946,N_14464);
xnor U19328 (N_19328,N_10039,N_14119);
nand U19329 (N_19329,N_13380,N_10362);
nand U19330 (N_19330,N_11431,N_10357);
or U19331 (N_19331,N_14272,N_10688);
nor U19332 (N_19332,N_14950,N_14834);
or U19333 (N_19333,N_13932,N_14095);
xor U19334 (N_19334,N_11633,N_14386);
xnor U19335 (N_19335,N_11692,N_10103);
nor U19336 (N_19336,N_12918,N_14165);
nand U19337 (N_19337,N_11407,N_10861);
xor U19338 (N_19338,N_14683,N_14842);
and U19339 (N_19339,N_10665,N_10556);
or U19340 (N_19340,N_12171,N_12493);
and U19341 (N_19341,N_12109,N_12114);
or U19342 (N_19342,N_13390,N_14488);
nor U19343 (N_19343,N_13692,N_12988);
nand U19344 (N_19344,N_10082,N_10936);
nand U19345 (N_19345,N_10686,N_10871);
nand U19346 (N_19346,N_13297,N_14335);
nand U19347 (N_19347,N_11816,N_13301);
xnor U19348 (N_19348,N_11073,N_12477);
nor U19349 (N_19349,N_11893,N_13110);
or U19350 (N_19350,N_10938,N_14310);
nor U19351 (N_19351,N_14370,N_11445);
or U19352 (N_19352,N_11401,N_11775);
or U19353 (N_19353,N_14938,N_11621);
nor U19354 (N_19354,N_14492,N_10281);
nand U19355 (N_19355,N_14542,N_12707);
xnor U19356 (N_19356,N_13913,N_10825);
nor U19357 (N_19357,N_11334,N_13053);
xor U19358 (N_19358,N_12403,N_14011);
xor U19359 (N_19359,N_10828,N_12871);
nand U19360 (N_19360,N_10017,N_14890);
nand U19361 (N_19361,N_14306,N_10804);
or U19362 (N_19362,N_10971,N_14688);
nor U19363 (N_19363,N_11018,N_10400);
and U19364 (N_19364,N_12056,N_11385);
or U19365 (N_19365,N_11584,N_10608);
or U19366 (N_19366,N_11518,N_11857);
nor U19367 (N_19367,N_13009,N_13751);
nor U19368 (N_19368,N_10043,N_12378);
nand U19369 (N_19369,N_12848,N_14475);
nor U19370 (N_19370,N_13376,N_12572);
xnor U19371 (N_19371,N_14534,N_12214);
or U19372 (N_19372,N_12086,N_12411);
or U19373 (N_19373,N_10200,N_12043);
nand U19374 (N_19374,N_13522,N_10554);
and U19375 (N_19375,N_11261,N_12779);
nor U19376 (N_19376,N_11130,N_10491);
nor U19377 (N_19377,N_10806,N_11474);
nor U19378 (N_19378,N_11377,N_10684);
nand U19379 (N_19379,N_11877,N_10442);
and U19380 (N_19380,N_12956,N_10734);
or U19381 (N_19381,N_13496,N_10606);
nand U19382 (N_19382,N_13758,N_10677);
nor U19383 (N_19383,N_12043,N_10736);
nand U19384 (N_19384,N_10760,N_14894);
nor U19385 (N_19385,N_14784,N_11832);
nor U19386 (N_19386,N_10304,N_13790);
nand U19387 (N_19387,N_14233,N_11267);
nand U19388 (N_19388,N_12698,N_13030);
nor U19389 (N_19389,N_14884,N_12675);
and U19390 (N_19390,N_11390,N_14941);
xnor U19391 (N_19391,N_14852,N_13902);
and U19392 (N_19392,N_12801,N_11450);
xnor U19393 (N_19393,N_14133,N_13537);
nor U19394 (N_19394,N_11033,N_11041);
xnor U19395 (N_19395,N_14156,N_12366);
xnor U19396 (N_19396,N_11857,N_10518);
nor U19397 (N_19397,N_12474,N_11917);
and U19398 (N_19398,N_10677,N_13802);
and U19399 (N_19399,N_11021,N_12789);
and U19400 (N_19400,N_12319,N_14537);
xor U19401 (N_19401,N_13890,N_14386);
nand U19402 (N_19402,N_13685,N_14901);
or U19403 (N_19403,N_14388,N_10015);
and U19404 (N_19404,N_12579,N_10499);
nand U19405 (N_19405,N_11846,N_11294);
nand U19406 (N_19406,N_13165,N_10176);
and U19407 (N_19407,N_14447,N_11754);
nor U19408 (N_19408,N_13160,N_10344);
xnor U19409 (N_19409,N_10568,N_12034);
and U19410 (N_19410,N_10166,N_10421);
nand U19411 (N_19411,N_14805,N_13519);
xor U19412 (N_19412,N_12807,N_12647);
nand U19413 (N_19413,N_12350,N_13913);
and U19414 (N_19414,N_10713,N_13532);
xor U19415 (N_19415,N_12787,N_13424);
nor U19416 (N_19416,N_10133,N_14099);
nor U19417 (N_19417,N_13775,N_13305);
xnor U19418 (N_19418,N_14183,N_10128);
xor U19419 (N_19419,N_12425,N_13796);
or U19420 (N_19420,N_10823,N_13624);
xor U19421 (N_19421,N_12735,N_11294);
nand U19422 (N_19422,N_11076,N_11640);
nand U19423 (N_19423,N_10052,N_14810);
xnor U19424 (N_19424,N_13152,N_12843);
nor U19425 (N_19425,N_13874,N_11013);
or U19426 (N_19426,N_14558,N_13372);
xnor U19427 (N_19427,N_14208,N_14356);
or U19428 (N_19428,N_10594,N_12171);
and U19429 (N_19429,N_13508,N_14594);
xnor U19430 (N_19430,N_13543,N_13721);
and U19431 (N_19431,N_14441,N_12492);
nand U19432 (N_19432,N_13561,N_12276);
nor U19433 (N_19433,N_10044,N_14365);
nor U19434 (N_19434,N_12287,N_14398);
nor U19435 (N_19435,N_12418,N_14426);
xnor U19436 (N_19436,N_14846,N_10379);
or U19437 (N_19437,N_13966,N_12987);
nor U19438 (N_19438,N_14943,N_13681);
or U19439 (N_19439,N_13265,N_14862);
or U19440 (N_19440,N_12262,N_10686);
nand U19441 (N_19441,N_11686,N_10930);
nor U19442 (N_19442,N_10047,N_11444);
nor U19443 (N_19443,N_14378,N_14658);
nor U19444 (N_19444,N_11307,N_12495);
nor U19445 (N_19445,N_10491,N_14053);
nor U19446 (N_19446,N_13548,N_12727);
nor U19447 (N_19447,N_13041,N_10066);
or U19448 (N_19448,N_10929,N_13045);
nor U19449 (N_19449,N_14131,N_14410);
nand U19450 (N_19450,N_12664,N_11795);
xnor U19451 (N_19451,N_14748,N_11097);
and U19452 (N_19452,N_12881,N_13779);
xor U19453 (N_19453,N_12993,N_12888);
nor U19454 (N_19454,N_10614,N_10116);
nor U19455 (N_19455,N_11303,N_13548);
and U19456 (N_19456,N_12273,N_10581);
or U19457 (N_19457,N_11351,N_12909);
xnor U19458 (N_19458,N_13979,N_11881);
and U19459 (N_19459,N_13223,N_12267);
and U19460 (N_19460,N_11140,N_10733);
nor U19461 (N_19461,N_12220,N_14079);
xor U19462 (N_19462,N_13637,N_12041);
nand U19463 (N_19463,N_10745,N_12284);
xor U19464 (N_19464,N_14845,N_14378);
nor U19465 (N_19465,N_14451,N_11204);
nand U19466 (N_19466,N_13203,N_10544);
or U19467 (N_19467,N_10170,N_14411);
nand U19468 (N_19468,N_10590,N_10917);
or U19469 (N_19469,N_13287,N_14164);
and U19470 (N_19470,N_13215,N_11245);
and U19471 (N_19471,N_10799,N_14421);
nor U19472 (N_19472,N_11992,N_13064);
nor U19473 (N_19473,N_12712,N_10047);
and U19474 (N_19474,N_14279,N_13292);
xnor U19475 (N_19475,N_12331,N_13218);
xor U19476 (N_19476,N_11843,N_11879);
xnor U19477 (N_19477,N_14566,N_10126);
nand U19478 (N_19478,N_13173,N_12692);
and U19479 (N_19479,N_13695,N_13311);
and U19480 (N_19480,N_14128,N_11303);
xnor U19481 (N_19481,N_11087,N_12009);
or U19482 (N_19482,N_13169,N_11001);
nand U19483 (N_19483,N_11305,N_10088);
or U19484 (N_19484,N_14324,N_10482);
xor U19485 (N_19485,N_12775,N_14386);
nor U19486 (N_19486,N_12552,N_10284);
xnor U19487 (N_19487,N_14408,N_14964);
or U19488 (N_19488,N_10131,N_10029);
and U19489 (N_19489,N_13508,N_10181);
or U19490 (N_19490,N_13966,N_13568);
nor U19491 (N_19491,N_11578,N_11165);
and U19492 (N_19492,N_12107,N_14786);
nand U19493 (N_19493,N_13109,N_12541);
and U19494 (N_19494,N_10642,N_12954);
xor U19495 (N_19495,N_10922,N_14382);
and U19496 (N_19496,N_12723,N_10131);
nand U19497 (N_19497,N_13955,N_10299);
nor U19498 (N_19498,N_11643,N_12043);
and U19499 (N_19499,N_14896,N_14319);
nand U19500 (N_19500,N_12885,N_12527);
nor U19501 (N_19501,N_14672,N_14099);
nor U19502 (N_19502,N_14251,N_13123);
nor U19503 (N_19503,N_12424,N_10706);
nor U19504 (N_19504,N_14370,N_12882);
or U19505 (N_19505,N_12048,N_13415);
nand U19506 (N_19506,N_11191,N_12503);
nand U19507 (N_19507,N_13269,N_11828);
and U19508 (N_19508,N_11921,N_14446);
or U19509 (N_19509,N_11452,N_11139);
and U19510 (N_19510,N_12804,N_13832);
or U19511 (N_19511,N_10435,N_12040);
and U19512 (N_19512,N_14347,N_11784);
xor U19513 (N_19513,N_13930,N_13856);
and U19514 (N_19514,N_14115,N_13690);
and U19515 (N_19515,N_12596,N_14203);
nor U19516 (N_19516,N_14003,N_12827);
xor U19517 (N_19517,N_10702,N_14465);
or U19518 (N_19518,N_11425,N_12560);
nor U19519 (N_19519,N_11889,N_13611);
or U19520 (N_19520,N_14097,N_14228);
nand U19521 (N_19521,N_10792,N_11732);
nand U19522 (N_19522,N_11393,N_12184);
nor U19523 (N_19523,N_13355,N_14647);
nand U19524 (N_19524,N_12493,N_11109);
nor U19525 (N_19525,N_11468,N_12713);
and U19526 (N_19526,N_13002,N_14926);
nand U19527 (N_19527,N_10674,N_13793);
and U19528 (N_19528,N_10253,N_10901);
and U19529 (N_19529,N_10020,N_14941);
nand U19530 (N_19530,N_10403,N_10289);
or U19531 (N_19531,N_11182,N_14225);
and U19532 (N_19532,N_10010,N_10281);
nand U19533 (N_19533,N_10464,N_14913);
and U19534 (N_19534,N_13190,N_12252);
and U19535 (N_19535,N_14505,N_10883);
or U19536 (N_19536,N_11186,N_14049);
nand U19537 (N_19537,N_12837,N_11626);
or U19538 (N_19538,N_10185,N_12288);
nor U19539 (N_19539,N_10879,N_11059);
nor U19540 (N_19540,N_10302,N_10543);
nand U19541 (N_19541,N_11039,N_11557);
xor U19542 (N_19542,N_10131,N_10227);
xor U19543 (N_19543,N_14931,N_12834);
and U19544 (N_19544,N_13215,N_11095);
and U19545 (N_19545,N_10631,N_10229);
xnor U19546 (N_19546,N_12638,N_14949);
xnor U19547 (N_19547,N_11183,N_11353);
or U19548 (N_19548,N_14548,N_10406);
nor U19549 (N_19549,N_12539,N_14162);
nor U19550 (N_19550,N_14286,N_10226);
or U19551 (N_19551,N_11732,N_10420);
and U19552 (N_19552,N_10712,N_11316);
nor U19553 (N_19553,N_10560,N_12562);
and U19554 (N_19554,N_14352,N_10788);
nor U19555 (N_19555,N_14933,N_10713);
and U19556 (N_19556,N_10485,N_10526);
and U19557 (N_19557,N_11640,N_12887);
and U19558 (N_19558,N_13870,N_13828);
or U19559 (N_19559,N_14717,N_13129);
nor U19560 (N_19560,N_13945,N_12209);
nand U19561 (N_19561,N_11488,N_13725);
nand U19562 (N_19562,N_14763,N_11108);
and U19563 (N_19563,N_10268,N_13562);
nand U19564 (N_19564,N_14826,N_11704);
xor U19565 (N_19565,N_13782,N_11519);
xor U19566 (N_19566,N_14395,N_11724);
nor U19567 (N_19567,N_11732,N_14961);
and U19568 (N_19568,N_10455,N_10400);
xor U19569 (N_19569,N_14364,N_12857);
or U19570 (N_19570,N_11540,N_10845);
xor U19571 (N_19571,N_14743,N_12548);
nand U19572 (N_19572,N_14717,N_11229);
or U19573 (N_19573,N_14809,N_10250);
nand U19574 (N_19574,N_13660,N_11730);
or U19575 (N_19575,N_14828,N_10123);
or U19576 (N_19576,N_14590,N_14663);
and U19577 (N_19577,N_14575,N_13637);
nand U19578 (N_19578,N_11826,N_13657);
and U19579 (N_19579,N_12611,N_12864);
and U19580 (N_19580,N_13823,N_10239);
xnor U19581 (N_19581,N_13111,N_10438);
nand U19582 (N_19582,N_14524,N_13007);
nor U19583 (N_19583,N_12714,N_14056);
xnor U19584 (N_19584,N_14628,N_11374);
or U19585 (N_19585,N_11400,N_13670);
nand U19586 (N_19586,N_14499,N_11316);
and U19587 (N_19587,N_13200,N_14158);
and U19588 (N_19588,N_14820,N_13000);
and U19589 (N_19589,N_12098,N_10793);
or U19590 (N_19590,N_11161,N_13064);
xor U19591 (N_19591,N_11498,N_11941);
nand U19592 (N_19592,N_11190,N_13716);
nand U19593 (N_19593,N_14427,N_14023);
nor U19594 (N_19594,N_12901,N_13992);
xnor U19595 (N_19595,N_10229,N_13971);
nor U19596 (N_19596,N_10200,N_13023);
or U19597 (N_19597,N_11818,N_12084);
and U19598 (N_19598,N_12970,N_11264);
and U19599 (N_19599,N_14375,N_12972);
nand U19600 (N_19600,N_11949,N_11870);
xor U19601 (N_19601,N_12988,N_12810);
or U19602 (N_19602,N_14249,N_14270);
xor U19603 (N_19603,N_11042,N_13264);
and U19604 (N_19604,N_14611,N_12563);
and U19605 (N_19605,N_12781,N_12918);
and U19606 (N_19606,N_11901,N_12392);
or U19607 (N_19607,N_10738,N_14081);
nor U19608 (N_19608,N_13875,N_10195);
xor U19609 (N_19609,N_13222,N_11647);
or U19610 (N_19610,N_11776,N_14806);
nor U19611 (N_19611,N_12963,N_14506);
or U19612 (N_19612,N_13614,N_11200);
nor U19613 (N_19613,N_13340,N_13976);
nand U19614 (N_19614,N_13291,N_11807);
and U19615 (N_19615,N_11646,N_14623);
nor U19616 (N_19616,N_10525,N_14618);
or U19617 (N_19617,N_12235,N_12367);
nor U19618 (N_19618,N_12315,N_11091);
nor U19619 (N_19619,N_10208,N_14595);
or U19620 (N_19620,N_11721,N_11802);
nor U19621 (N_19621,N_14081,N_12860);
or U19622 (N_19622,N_10572,N_13829);
and U19623 (N_19623,N_11209,N_12042);
nand U19624 (N_19624,N_10907,N_14736);
or U19625 (N_19625,N_12888,N_12309);
nor U19626 (N_19626,N_10515,N_14726);
or U19627 (N_19627,N_11813,N_13582);
xor U19628 (N_19628,N_11111,N_10560);
nor U19629 (N_19629,N_14467,N_10625);
or U19630 (N_19630,N_14704,N_14731);
xnor U19631 (N_19631,N_14353,N_12068);
nand U19632 (N_19632,N_12999,N_12250);
nand U19633 (N_19633,N_14456,N_12379);
or U19634 (N_19634,N_13163,N_11557);
and U19635 (N_19635,N_12252,N_14689);
nor U19636 (N_19636,N_10974,N_13964);
nand U19637 (N_19637,N_14471,N_10994);
nand U19638 (N_19638,N_11340,N_10969);
and U19639 (N_19639,N_12631,N_14020);
nand U19640 (N_19640,N_11241,N_14498);
nor U19641 (N_19641,N_10237,N_11118);
and U19642 (N_19642,N_12061,N_14578);
xnor U19643 (N_19643,N_10444,N_11877);
xor U19644 (N_19644,N_12882,N_10198);
or U19645 (N_19645,N_13149,N_10146);
or U19646 (N_19646,N_12308,N_13727);
nor U19647 (N_19647,N_10367,N_12737);
nor U19648 (N_19648,N_13222,N_11464);
or U19649 (N_19649,N_13618,N_13083);
nor U19650 (N_19650,N_11713,N_11221);
nand U19651 (N_19651,N_11265,N_11670);
xor U19652 (N_19652,N_11251,N_11832);
and U19653 (N_19653,N_11614,N_10819);
xnor U19654 (N_19654,N_12713,N_12108);
nor U19655 (N_19655,N_14593,N_14634);
or U19656 (N_19656,N_13661,N_13091);
xnor U19657 (N_19657,N_14821,N_10411);
or U19658 (N_19658,N_10625,N_13335);
and U19659 (N_19659,N_14292,N_14467);
or U19660 (N_19660,N_14770,N_10488);
nand U19661 (N_19661,N_12488,N_10774);
nor U19662 (N_19662,N_11339,N_10200);
xor U19663 (N_19663,N_13613,N_10730);
nand U19664 (N_19664,N_14894,N_11510);
xor U19665 (N_19665,N_13637,N_10139);
nand U19666 (N_19666,N_13955,N_13790);
xor U19667 (N_19667,N_12269,N_13114);
and U19668 (N_19668,N_11962,N_10555);
xor U19669 (N_19669,N_14233,N_14954);
and U19670 (N_19670,N_11330,N_14597);
xor U19671 (N_19671,N_11702,N_11475);
or U19672 (N_19672,N_10112,N_12649);
nand U19673 (N_19673,N_13719,N_10168);
nor U19674 (N_19674,N_10466,N_12274);
xor U19675 (N_19675,N_10919,N_10777);
nand U19676 (N_19676,N_10930,N_12749);
or U19677 (N_19677,N_14239,N_10845);
and U19678 (N_19678,N_14092,N_11210);
and U19679 (N_19679,N_11879,N_10931);
and U19680 (N_19680,N_13340,N_13336);
or U19681 (N_19681,N_11392,N_10273);
and U19682 (N_19682,N_14945,N_10090);
or U19683 (N_19683,N_10680,N_13381);
or U19684 (N_19684,N_12704,N_14735);
and U19685 (N_19685,N_10199,N_11063);
or U19686 (N_19686,N_14186,N_14774);
and U19687 (N_19687,N_14052,N_10207);
nor U19688 (N_19688,N_12515,N_12133);
nand U19689 (N_19689,N_14287,N_10215);
xnor U19690 (N_19690,N_12170,N_12192);
or U19691 (N_19691,N_10893,N_11422);
and U19692 (N_19692,N_11574,N_11948);
or U19693 (N_19693,N_14579,N_13831);
xor U19694 (N_19694,N_14158,N_13296);
xnor U19695 (N_19695,N_12104,N_14412);
xnor U19696 (N_19696,N_10947,N_10786);
and U19697 (N_19697,N_11457,N_13605);
and U19698 (N_19698,N_10162,N_12412);
xnor U19699 (N_19699,N_14190,N_12734);
and U19700 (N_19700,N_12387,N_14450);
nand U19701 (N_19701,N_10683,N_11084);
xnor U19702 (N_19702,N_14586,N_10498);
or U19703 (N_19703,N_14352,N_10162);
and U19704 (N_19704,N_13715,N_10783);
nand U19705 (N_19705,N_11731,N_14442);
or U19706 (N_19706,N_10664,N_14546);
nand U19707 (N_19707,N_10441,N_10594);
and U19708 (N_19708,N_14835,N_11599);
or U19709 (N_19709,N_14358,N_14569);
or U19710 (N_19710,N_11352,N_10654);
xor U19711 (N_19711,N_12399,N_12742);
nand U19712 (N_19712,N_10235,N_11865);
nor U19713 (N_19713,N_11834,N_11727);
xnor U19714 (N_19714,N_13840,N_12333);
nand U19715 (N_19715,N_12320,N_11985);
nor U19716 (N_19716,N_10140,N_11232);
nor U19717 (N_19717,N_14505,N_10360);
and U19718 (N_19718,N_13453,N_10105);
nor U19719 (N_19719,N_11656,N_11335);
and U19720 (N_19720,N_14512,N_13532);
nand U19721 (N_19721,N_11212,N_13189);
and U19722 (N_19722,N_12688,N_12806);
nand U19723 (N_19723,N_12047,N_10612);
nand U19724 (N_19724,N_12456,N_11441);
or U19725 (N_19725,N_11136,N_13375);
nand U19726 (N_19726,N_11433,N_11546);
nand U19727 (N_19727,N_10758,N_14808);
or U19728 (N_19728,N_12887,N_11038);
nor U19729 (N_19729,N_13391,N_12095);
or U19730 (N_19730,N_11119,N_12549);
nand U19731 (N_19731,N_13427,N_14957);
or U19732 (N_19732,N_11267,N_11061);
or U19733 (N_19733,N_13386,N_10027);
or U19734 (N_19734,N_10864,N_11093);
or U19735 (N_19735,N_14206,N_12773);
or U19736 (N_19736,N_10554,N_14881);
xor U19737 (N_19737,N_12326,N_11787);
and U19738 (N_19738,N_11886,N_13153);
or U19739 (N_19739,N_13157,N_11568);
or U19740 (N_19740,N_11532,N_13323);
nand U19741 (N_19741,N_14818,N_11112);
or U19742 (N_19742,N_14462,N_12971);
nand U19743 (N_19743,N_13721,N_10177);
nor U19744 (N_19744,N_14115,N_14029);
nor U19745 (N_19745,N_10636,N_14940);
nor U19746 (N_19746,N_13139,N_10035);
nand U19747 (N_19747,N_10579,N_14926);
nand U19748 (N_19748,N_13437,N_12902);
or U19749 (N_19749,N_14324,N_10579);
nand U19750 (N_19750,N_10731,N_10784);
or U19751 (N_19751,N_10772,N_11959);
xor U19752 (N_19752,N_12250,N_10203);
nand U19753 (N_19753,N_14108,N_11100);
nand U19754 (N_19754,N_13994,N_13276);
or U19755 (N_19755,N_12760,N_11037);
nor U19756 (N_19756,N_12350,N_10174);
xnor U19757 (N_19757,N_13687,N_10007);
nand U19758 (N_19758,N_11361,N_11558);
or U19759 (N_19759,N_13199,N_12333);
or U19760 (N_19760,N_12923,N_11601);
or U19761 (N_19761,N_14406,N_14858);
nor U19762 (N_19762,N_11766,N_12641);
xnor U19763 (N_19763,N_13989,N_13254);
or U19764 (N_19764,N_13359,N_14552);
xor U19765 (N_19765,N_13092,N_11248);
xor U19766 (N_19766,N_10639,N_13055);
xnor U19767 (N_19767,N_11534,N_12622);
nand U19768 (N_19768,N_14172,N_13250);
or U19769 (N_19769,N_11453,N_10733);
nor U19770 (N_19770,N_13680,N_14612);
xor U19771 (N_19771,N_12485,N_11829);
and U19772 (N_19772,N_13135,N_12876);
xor U19773 (N_19773,N_10204,N_14445);
xor U19774 (N_19774,N_12751,N_14630);
nand U19775 (N_19775,N_10973,N_12364);
or U19776 (N_19776,N_13290,N_14155);
xor U19777 (N_19777,N_10886,N_12902);
and U19778 (N_19778,N_14923,N_14335);
and U19779 (N_19779,N_10501,N_10487);
xor U19780 (N_19780,N_12346,N_10431);
nor U19781 (N_19781,N_14638,N_12792);
and U19782 (N_19782,N_12862,N_10482);
xor U19783 (N_19783,N_13745,N_14649);
nor U19784 (N_19784,N_10282,N_11133);
or U19785 (N_19785,N_13910,N_14718);
or U19786 (N_19786,N_12919,N_13134);
nor U19787 (N_19787,N_14498,N_11897);
xor U19788 (N_19788,N_14702,N_13425);
or U19789 (N_19789,N_11121,N_10694);
xnor U19790 (N_19790,N_12452,N_12103);
or U19791 (N_19791,N_12617,N_12145);
or U19792 (N_19792,N_12200,N_12920);
nor U19793 (N_19793,N_10680,N_10002);
or U19794 (N_19794,N_11012,N_14404);
xnor U19795 (N_19795,N_14182,N_14746);
and U19796 (N_19796,N_10788,N_12802);
and U19797 (N_19797,N_11559,N_11789);
or U19798 (N_19798,N_10564,N_10249);
nand U19799 (N_19799,N_11469,N_11891);
xnor U19800 (N_19800,N_11280,N_12872);
nor U19801 (N_19801,N_14677,N_11995);
or U19802 (N_19802,N_12193,N_11433);
or U19803 (N_19803,N_10917,N_13461);
or U19804 (N_19804,N_10551,N_12460);
xor U19805 (N_19805,N_12213,N_11588);
and U19806 (N_19806,N_13191,N_14371);
and U19807 (N_19807,N_11327,N_10163);
nor U19808 (N_19808,N_10030,N_13073);
or U19809 (N_19809,N_11708,N_12474);
xor U19810 (N_19810,N_13687,N_13277);
nor U19811 (N_19811,N_14776,N_12522);
xor U19812 (N_19812,N_11066,N_13344);
and U19813 (N_19813,N_12059,N_14599);
xor U19814 (N_19814,N_11421,N_11106);
or U19815 (N_19815,N_11347,N_12997);
and U19816 (N_19816,N_10930,N_14809);
or U19817 (N_19817,N_11298,N_13604);
nand U19818 (N_19818,N_14808,N_11437);
nor U19819 (N_19819,N_11998,N_14922);
and U19820 (N_19820,N_13137,N_11334);
and U19821 (N_19821,N_14146,N_13416);
nand U19822 (N_19822,N_10674,N_11113);
nor U19823 (N_19823,N_10754,N_14492);
xnor U19824 (N_19824,N_10775,N_10909);
and U19825 (N_19825,N_12412,N_13620);
nor U19826 (N_19826,N_14119,N_14002);
and U19827 (N_19827,N_12654,N_12898);
or U19828 (N_19828,N_10842,N_12854);
xnor U19829 (N_19829,N_10150,N_12604);
nor U19830 (N_19830,N_12342,N_10414);
or U19831 (N_19831,N_10866,N_13774);
nand U19832 (N_19832,N_14179,N_11029);
nor U19833 (N_19833,N_10199,N_10285);
or U19834 (N_19834,N_11384,N_12004);
xor U19835 (N_19835,N_11722,N_12224);
and U19836 (N_19836,N_12704,N_11629);
and U19837 (N_19837,N_13123,N_13089);
xor U19838 (N_19838,N_13436,N_10548);
and U19839 (N_19839,N_14397,N_11336);
xnor U19840 (N_19840,N_10447,N_12269);
nor U19841 (N_19841,N_12248,N_13823);
or U19842 (N_19842,N_12498,N_12189);
xnor U19843 (N_19843,N_12589,N_10168);
or U19844 (N_19844,N_11353,N_13949);
or U19845 (N_19845,N_14665,N_13720);
nor U19846 (N_19846,N_12747,N_13669);
and U19847 (N_19847,N_14208,N_11382);
nand U19848 (N_19848,N_10728,N_10221);
nand U19849 (N_19849,N_12148,N_12319);
xor U19850 (N_19850,N_11760,N_14300);
or U19851 (N_19851,N_14436,N_13906);
and U19852 (N_19852,N_12858,N_10518);
nor U19853 (N_19853,N_10087,N_12684);
xor U19854 (N_19854,N_10789,N_12854);
nor U19855 (N_19855,N_13722,N_11130);
nand U19856 (N_19856,N_14890,N_12639);
nor U19857 (N_19857,N_14451,N_13018);
and U19858 (N_19858,N_12406,N_12300);
nand U19859 (N_19859,N_13209,N_12991);
or U19860 (N_19860,N_12054,N_11177);
nand U19861 (N_19861,N_14305,N_13762);
and U19862 (N_19862,N_11496,N_13432);
and U19863 (N_19863,N_13731,N_14020);
and U19864 (N_19864,N_13868,N_10140);
and U19865 (N_19865,N_11182,N_10930);
nand U19866 (N_19866,N_11811,N_11490);
or U19867 (N_19867,N_11627,N_13187);
and U19868 (N_19868,N_11018,N_11375);
xor U19869 (N_19869,N_10939,N_12246);
or U19870 (N_19870,N_14552,N_11786);
nor U19871 (N_19871,N_12764,N_11457);
and U19872 (N_19872,N_14556,N_13070);
xnor U19873 (N_19873,N_10480,N_12744);
or U19874 (N_19874,N_10505,N_11399);
and U19875 (N_19875,N_11060,N_10340);
nor U19876 (N_19876,N_13516,N_11761);
nor U19877 (N_19877,N_10036,N_12489);
and U19878 (N_19878,N_10792,N_12687);
nand U19879 (N_19879,N_11954,N_13036);
or U19880 (N_19880,N_10909,N_11604);
nand U19881 (N_19881,N_12812,N_13545);
xor U19882 (N_19882,N_12898,N_12784);
nand U19883 (N_19883,N_14242,N_11986);
nor U19884 (N_19884,N_11404,N_12471);
and U19885 (N_19885,N_13447,N_13090);
or U19886 (N_19886,N_13107,N_12476);
or U19887 (N_19887,N_14771,N_14491);
xor U19888 (N_19888,N_13866,N_11054);
xor U19889 (N_19889,N_14122,N_12224);
xor U19890 (N_19890,N_11873,N_10126);
and U19891 (N_19891,N_10744,N_10388);
nor U19892 (N_19892,N_12256,N_12463);
or U19893 (N_19893,N_12871,N_12155);
and U19894 (N_19894,N_14064,N_10725);
and U19895 (N_19895,N_12571,N_14545);
and U19896 (N_19896,N_10198,N_14226);
or U19897 (N_19897,N_10097,N_11293);
nor U19898 (N_19898,N_13343,N_10796);
and U19899 (N_19899,N_12071,N_11437);
xnor U19900 (N_19900,N_11199,N_11054);
and U19901 (N_19901,N_12267,N_13448);
or U19902 (N_19902,N_10416,N_13662);
or U19903 (N_19903,N_13056,N_14383);
or U19904 (N_19904,N_13326,N_14944);
and U19905 (N_19905,N_11723,N_14023);
or U19906 (N_19906,N_13135,N_12631);
or U19907 (N_19907,N_12050,N_10995);
and U19908 (N_19908,N_10630,N_13233);
nand U19909 (N_19909,N_13521,N_13638);
nor U19910 (N_19910,N_11140,N_13127);
xor U19911 (N_19911,N_12620,N_13511);
xor U19912 (N_19912,N_14159,N_10430);
xor U19913 (N_19913,N_11923,N_13015);
and U19914 (N_19914,N_10808,N_12907);
nor U19915 (N_19915,N_14771,N_13952);
nor U19916 (N_19916,N_13650,N_13760);
xnor U19917 (N_19917,N_13146,N_14548);
xor U19918 (N_19918,N_14241,N_12104);
xnor U19919 (N_19919,N_11548,N_13043);
or U19920 (N_19920,N_13081,N_11955);
or U19921 (N_19921,N_13899,N_13616);
or U19922 (N_19922,N_13604,N_11477);
and U19923 (N_19923,N_14682,N_14004);
nand U19924 (N_19924,N_14890,N_12086);
nand U19925 (N_19925,N_14542,N_11820);
nand U19926 (N_19926,N_14977,N_14354);
xnor U19927 (N_19927,N_13275,N_11241);
or U19928 (N_19928,N_10922,N_12142);
and U19929 (N_19929,N_10019,N_11744);
xnor U19930 (N_19930,N_14327,N_10023);
xor U19931 (N_19931,N_14433,N_13961);
or U19932 (N_19932,N_10352,N_12567);
xor U19933 (N_19933,N_14551,N_14070);
and U19934 (N_19934,N_11028,N_12376);
xnor U19935 (N_19935,N_14342,N_14250);
nor U19936 (N_19936,N_10949,N_14159);
xnor U19937 (N_19937,N_14297,N_14696);
nand U19938 (N_19938,N_13448,N_10366);
xor U19939 (N_19939,N_11743,N_10119);
nor U19940 (N_19940,N_11463,N_14742);
or U19941 (N_19941,N_14066,N_13617);
nand U19942 (N_19942,N_14743,N_12028);
xnor U19943 (N_19943,N_12126,N_10689);
nand U19944 (N_19944,N_13380,N_11696);
and U19945 (N_19945,N_14849,N_13766);
xnor U19946 (N_19946,N_11750,N_13823);
nor U19947 (N_19947,N_13417,N_11798);
or U19948 (N_19948,N_11731,N_13472);
or U19949 (N_19949,N_12737,N_11648);
xor U19950 (N_19950,N_12769,N_14197);
and U19951 (N_19951,N_13162,N_12450);
xor U19952 (N_19952,N_12710,N_11122);
xnor U19953 (N_19953,N_10340,N_12768);
or U19954 (N_19954,N_11486,N_12896);
xnor U19955 (N_19955,N_10027,N_13290);
or U19956 (N_19956,N_14686,N_13214);
and U19957 (N_19957,N_11217,N_10013);
or U19958 (N_19958,N_11624,N_11809);
and U19959 (N_19959,N_14992,N_14132);
nor U19960 (N_19960,N_13432,N_14800);
and U19961 (N_19961,N_10868,N_12545);
xor U19962 (N_19962,N_13050,N_12021);
and U19963 (N_19963,N_13943,N_14328);
xor U19964 (N_19964,N_13823,N_14679);
or U19965 (N_19965,N_10449,N_12912);
nand U19966 (N_19966,N_11750,N_12067);
and U19967 (N_19967,N_14171,N_14941);
and U19968 (N_19968,N_14990,N_13318);
xnor U19969 (N_19969,N_10817,N_11919);
xnor U19970 (N_19970,N_13381,N_14752);
nor U19971 (N_19971,N_11257,N_13265);
nor U19972 (N_19972,N_12673,N_12916);
xor U19973 (N_19973,N_14986,N_14394);
xor U19974 (N_19974,N_12121,N_12099);
nand U19975 (N_19975,N_13473,N_10850);
or U19976 (N_19976,N_10725,N_14289);
xor U19977 (N_19977,N_12957,N_12858);
nand U19978 (N_19978,N_14271,N_11237);
or U19979 (N_19979,N_13071,N_13606);
and U19980 (N_19980,N_14835,N_13677);
xnor U19981 (N_19981,N_10184,N_12842);
nor U19982 (N_19982,N_11986,N_14331);
or U19983 (N_19983,N_11262,N_11705);
or U19984 (N_19984,N_13983,N_11759);
nand U19985 (N_19985,N_11390,N_11446);
and U19986 (N_19986,N_11292,N_10884);
xnor U19987 (N_19987,N_11946,N_11932);
xor U19988 (N_19988,N_14698,N_11931);
and U19989 (N_19989,N_10945,N_13191);
xor U19990 (N_19990,N_13771,N_13070);
and U19991 (N_19991,N_12216,N_10777);
or U19992 (N_19992,N_12371,N_10885);
nand U19993 (N_19993,N_14427,N_14141);
nor U19994 (N_19994,N_10292,N_11746);
nand U19995 (N_19995,N_11856,N_14202);
and U19996 (N_19996,N_14408,N_10231);
or U19997 (N_19997,N_14647,N_11030);
xor U19998 (N_19998,N_11616,N_10293);
xor U19999 (N_19999,N_11535,N_12394);
or U20000 (N_20000,N_17484,N_15555);
and U20001 (N_20001,N_15352,N_19351);
nor U20002 (N_20002,N_16343,N_19932);
nor U20003 (N_20003,N_16031,N_19274);
nand U20004 (N_20004,N_15663,N_18575);
xnor U20005 (N_20005,N_19070,N_18329);
or U20006 (N_20006,N_19815,N_15870);
xor U20007 (N_20007,N_18419,N_17227);
or U20008 (N_20008,N_19574,N_18499);
nand U20009 (N_20009,N_17667,N_17124);
nor U20010 (N_20010,N_19522,N_17017);
xnor U20011 (N_20011,N_16183,N_18551);
or U20012 (N_20012,N_16772,N_17783);
and U20013 (N_20013,N_18665,N_16602);
or U20014 (N_20014,N_19024,N_17800);
xor U20015 (N_20015,N_19993,N_16640);
nand U20016 (N_20016,N_17019,N_18463);
xnor U20017 (N_20017,N_19746,N_15368);
nand U20018 (N_20018,N_19558,N_15562);
nor U20019 (N_20019,N_17836,N_17307);
and U20020 (N_20020,N_15742,N_19719);
or U20021 (N_20021,N_17905,N_19144);
and U20022 (N_20022,N_18564,N_18642);
nor U20023 (N_20023,N_16252,N_15264);
xnor U20024 (N_20024,N_16756,N_17034);
xor U20025 (N_20025,N_17635,N_18236);
nor U20026 (N_20026,N_18561,N_16639);
nor U20027 (N_20027,N_16648,N_19565);
xor U20028 (N_20028,N_17389,N_18605);
nand U20029 (N_20029,N_18929,N_16040);
and U20030 (N_20030,N_16520,N_15575);
and U20031 (N_20031,N_16060,N_19515);
xor U20032 (N_20032,N_16903,N_15461);
or U20033 (N_20033,N_15434,N_16030);
xnor U20034 (N_20034,N_19092,N_17722);
xnor U20035 (N_20035,N_18442,N_16697);
nand U20036 (N_20036,N_15541,N_15448);
xor U20037 (N_20037,N_18336,N_18909);
or U20038 (N_20038,N_16306,N_19979);
nor U20039 (N_20039,N_19425,N_17180);
nand U20040 (N_20040,N_18550,N_15818);
and U20041 (N_20041,N_15805,N_17595);
nor U20042 (N_20042,N_15869,N_19026);
xnor U20043 (N_20043,N_19317,N_16690);
and U20044 (N_20044,N_18720,N_18973);
nor U20045 (N_20045,N_19588,N_19373);
xor U20046 (N_20046,N_15308,N_19028);
and U20047 (N_20047,N_17191,N_17195);
nor U20048 (N_20048,N_17750,N_18179);
nor U20049 (N_20049,N_18873,N_16975);
and U20050 (N_20050,N_15420,N_19275);
or U20051 (N_20051,N_15254,N_16416);
and U20052 (N_20052,N_15302,N_16966);
xor U20053 (N_20053,N_16887,N_17300);
and U20054 (N_20054,N_18826,N_15186);
xor U20055 (N_20055,N_19641,N_17039);
nor U20056 (N_20056,N_19450,N_19202);
and U20057 (N_20057,N_19777,N_16411);
nor U20058 (N_20058,N_15521,N_15674);
or U20059 (N_20059,N_19171,N_16522);
nand U20060 (N_20060,N_17182,N_17989);
xnor U20061 (N_20061,N_19420,N_18216);
nor U20062 (N_20062,N_19363,N_17707);
nand U20063 (N_20063,N_18253,N_17407);
and U20064 (N_20064,N_18633,N_18379);
or U20065 (N_20065,N_18144,N_15848);
nor U20066 (N_20066,N_15897,N_19455);
or U20067 (N_20067,N_15533,N_17062);
nor U20068 (N_20068,N_19090,N_18387);
nor U20069 (N_20069,N_16187,N_16022);
or U20070 (N_20070,N_18662,N_17700);
and U20071 (N_20071,N_19963,N_18680);
or U20072 (N_20072,N_17033,N_16382);
and U20073 (N_20073,N_18539,N_15898);
or U20074 (N_20074,N_19494,N_17310);
nand U20075 (N_20075,N_17998,N_19422);
or U20076 (N_20076,N_18765,N_19726);
nand U20077 (N_20077,N_17682,N_17961);
xor U20078 (N_20078,N_15202,N_16071);
and U20079 (N_20079,N_18712,N_17174);
or U20080 (N_20080,N_17398,N_19778);
xor U20081 (N_20081,N_18233,N_16097);
and U20082 (N_20082,N_19694,N_17984);
xor U20083 (N_20083,N_17817,N_16247);
and U20084 (N_20084,N_16625,N_17514);
and U20085 (N_20085,N_18975,N_18100);
and U20086 (N_20086,N_15179,N_18173);
nor U20087 (N_20087,N_15635,N_17952);
or U20088 (N_20088,N_18494,N_17141);
nor U20089 (N_20089,N_17269,N_18214);
nand U20090 (N_20090,N_16667,N_15907);
nor U20091 (N_20091,N_19985,N_15058);
or U20092 (N_20092,N_15799,N_16188);
nand U20093 (N_20093,N_17757,N_19721);
and U20094 (N_20094,N_15989,N_18604);
or U20095 (N_20095,N_17348,N_15713);
nand U20096 (N_20096,N_19811,N_19060);
nand U20097 (N_20097,N_18506,N_18485);
xnor U20098 (N_20098,N_16731,N_19414);
nor U20099 (N_20099,N_15846,N_19528);
xor U20100 (N_20100,N_17944,N_19232);
and U20101 (N_20101,N_19320,N_15084);
nor U20102 (N_20102,N_18952,N_16531);
or U20103 (N_20103,N_15594,N_15294);
nand U20104 (N_20104,N_16823,N_17327);
nor U20105 (N_20105,N_18113,N_15172);
and U20106 (N_20106,N_17705,N_16278);
nor U20107 (N_20107,N_18472,N_16855);
and U20108 (N_20108,N_16447,N_15191);
xnor U20109 (N_20109,N_16174,N_15245);
nor U20110 (N_20110,N_19483,N_15767);
nand U20111 (N_20111,N_19261,N_16897);
nor U20112 (N_20112,N_18710,N_17451);
nor U20113 (N_20113,N_17094,N_18822);
or U20114 (N_20114,N_18637,N_15388);
nor U20115 (N_20115,N_16563,N_17671);
and U20116 (N_20116,N_16679,N_17736);
and U20117 (N_20117,N_16961,N_15821);
or U20118 (N_20118,N_15291,N_16184);
and U20119 (N_20119,N_15181,N_18203);
nand U20120 (N_20120,N_19595,N_17012);
nand U20121 (N_20121,N_15085,N_17518);
and U20122 (N_20122,N_18423,N_15653);
xor U20123 (N_20123,N_15675,N_17409);
xnor U20124 (N_20124,N_19367,N_17250);
or U20125 (N_20125,N_18683,N_15959);
nand U20126 (N_20126,N_17354,N_18953);
or U20127 (N_20127,N_17274,N_16946);
nand U20128 (N_20128,N_19919,N_19032);
xor U20129 (N_20129,N_16718,N_18354);
nand U20130 (N_20130,N_17714,N_17555);
and U20131 (N_20131,N_19133,N_18139);
and U20132 (N_20132,N_16154,N_17218);
nand U20133 (N_20133,N_19710,N_16852);
xor U20134 (N_20134,N_17925,N_15692);
and U20135 (N_20135,N_18047,N_16319);
nor U20136 (N_20136,N_18502,N_15733);
nor U20137 (N_20137,N_17474,N_18478);
xor U20138 (N_20138,N_16970,N_15946);
xnor U20139 (N_20139,N_19017,N_15495);
xor U20140 (N_20140,N_19504,N_17365);
nand U20141 (N_20141,N_16711,N_18407);
and U20142 (N_20142,N_17076,N_19767);
xor U20143 (N_20143,N_18375,N_18532);
or U20144 (N_20144,N_16397,N_19552);
or U20145 (N_20145,N_18666,N_16534);
nand U20146 (N_20146,N_15396,N_18774);
xnor U20147 (N_20147,N_18938,N_15681);
nand U20148 (N_20148,N_19176,N_18092);
nand U20149 (N_20149,N_15778,N_17044);
nor U20150 (N_20150,N_17070,N_16923);
or U20151 (N_20151,N_17403,N_15343);
and U20152 (N_20152,N_15826,N_18837);
xor U20153 (N_20153,N_18793,N_18308);
nor U20154 (N_20154,N_18754,N_15101);
or U20155 (N_20155,N_18490,N_19946);
nor U20156 (N_20156,N_19853,N_16011);
nand U20157 (N_20157,N_15445,N_17534);
or U20158 (N_20158,N_18374,N_16387);
nand U20159 (N_20159,N_19696,N_15964);
and U20160 (N_20160,N_16224,N_18274);
and U20161 (N_20161,N_18220,N_18792);
and U20162 (N_20162,N_17129,N_15616);
or U20163 (N_20163,N_17346,N_17446);
or U20164 (N_20164,N_19897,N_15392);
or U20165 (N_20165,N_18381,N_19354);
xnor U20166 (N_20166,N_17460,N_15912);
nor U20167 (N_20167,N_19143,N_17367);
and U20168 (N_20168,N_18933,N_19905);
xnor U20169 (N_20169,N_19471,N_18635);
and U20170 (N_20170,N_19125,N_17316);
nand U20171 (N_20171,N_17099,N_15716);
or U20172 (N_20172,N_17261,N_15626);
or U20173 (N_20173,N_16332,N_18713);
nand U20174 (N_20174,N_18135,N_17976);
or U20175 (N_20175,N_18195,N_15809);
or U20176 (N_20176,N_19755,N_19251);
and U20177 (N_20177,N_16944,N_18342);
xnor U20178 (N_20178,N_17148,N_17499);
or U20179 (N_20179,N_18649,N_16094);
or U20180 (N_20180,N_19589,N_17030);
nor U20181 (N_20181,N_16485,N_18914);
and U20182 (N_20182,N_18142,N_16084);
xor U20183 (N_20183,N_18402,N_17536);
nor U20184 (N_20184,N_16118,N_19357);
nand U20185 (N_20185,N_15197,N_15487);
and U20186 (N_20186,N_16431,N_16902);
and U20187 (N_20187,N_17888,N_18185);
xor U20188 (N_20188,N_17724,N_19831);
nor U20189 (N_20189,N_15304,N_18722);
or U20190 (N_20190,N_16231,N_16845);
and U20191 (N_20191,N_19875,N_16034);
xnor U20192 (N_20192,N_17220,N_17073);
or U20193 (N_20193,N_19975,N_18303);
and U20194 (N_20194,N_19813,N_19272);
xor U20195 (N_20195,N_18225,N_15770);
nor U20196 (N_20196,N_16645,N_17337);
or U20197 (N_20197,N_17709,N_19240);
xnor U20198 (N_20198,N_18249,N_17100);
nor U20199 (N_20199,N_19680,N_19361);
nand U20200 (N_20200,N_19734,N_15173);
or U20201 (N_20201,N_15267,N_15646);
and U20202 (N_20202,N_16407,N_18339);
xnor U20203 (N_20203,N_17511,N_19447);
nor U20204 (N_20204,N_18291,N_15425);
nand U20205 (N_20205,N_16569,N_19517);
nand U20206 (N_20206,N_15225,N_19915);
xor U20207 (N_20207,N_17864,N_19200);
nor U20208 (N_20208,N_18698,N_18555);
xnor U20209 (N_20209,N_19702,N_15033);
nand U20210 (N_20210,N_19325,N_19646);
nor U20211 (N_20211,N_19224,N_15205);
or U20212 (N_20212,N_18739,N_17296);
xnor U20213 (N_20213,N_19663,N_19305);
nor U20214 (N_20214,N_19252,N_19645);
and U20215 (N_20215,N_18828,N_16559);
nor U20216 (N_20216,N_16781,N_16102);
xnor U20217 (N_20217,N_18153,N_16934);
nor U20218 (N_20218,N_16589,N_16585);
xor U20219 (N_20219,N_17929,N_16926);
nand U20220 (N_20220,N_18138,N_19713);
or U20221 (N_20221,N_15362,N_18756);
and U20222 (N_20222,N_17875,N_19923);
and U20223 (N_20223,N_16792,N_15330);
nand U20224 (N_20224,N_15451,N_17396);
xnor U20225 (N_20225,N_17320,N_15080);
nand U20226 (N_20226,N_15932,N_16186);
and U20227 (N_20227,N_17985,N_18706);
or U20228 (N_20228,N_19674,N_17428);
and U20229 (N_20229,N_16227,N_18278);
nand U20230 (N_20230,N_19877,N_19970);
nand U20231 (N_20231,N_17542,N_16225);
nand U20232 (N_20232,N_17262,N_15927);
and U20233 (N_20233,N_16012,N_19671);
or U20234 (N_20234,N_15542,N_16169);
xnor U20235 (N_20235,N_16738,N_18209);
nor U20236 (N_20236,N_16991,N_17416);
nand U20237 (N_20237,N_16873,N_18062);
nor U20238 (N_20238,N_16635,N_18037);
xnor U20239 (N_20239,N_19888,N_16010);
xnor U20240 (N_20240,N_16665,N_19010);
nand U20241 (N_20241,N_16208,N_18943);
nor U20242 (N_20242,N_19554,N_15129);
and U20243 (N_20243,N_17892,N_18513);
nand U20244 (N_20244,N_15170,N_19122);
or U20245 (N_20245,N_18071,N_17057);
nand U20246 (N_20246,N_16006,N_19188);
nand U20247 (N_20247,N_19748,N_18476);
nor U20248 (N_20248,N_16850,N_18978);
and U20249 (N_20249,N_15522,N_16391);
nand U20250 (N_20250,N_18987,N_19764);
nor U20251 (N_20251,N_15250,N_16253);
nand U20252 (N_20252,N_19747,N_19661);
nand U20253 (N_20253,N_19759,N_17489);
xor U20254 (N_20254,N_15666,N_17882);
or U20255 (N_20255,N_16583,N_19869);
xor U20256 (N_20256,N_17157,N_18385);
nand U20257 (N_20257,N_16308,N_19901);
and U20258 (N_20258,N_16777,N_17745);
xnor U20259 (N_20259,N_15365,N_16379);
nor U20260 (N_20260,N_16417,N_19986);
and U20261 (N_20261,N_17808,N_17498);
xor U20262 (N_20262,N_15473,N_19805);
and U20263 (N_20263,N_16784,N_17177);
and U20264 (N_20264,N_17924,N_19769);
or U20265 (N_20265,N_17936,N_16812);
or U20266 (N_20266,N_16920,N_16380);
and U20267 (N_20267,N_15501,N_19206);
nand U20268 (N_20268,N_16468,N_16594);
xnor U20269 (N_20269,N_17459,N_18076);
nand U20270 (N_20270,N_19794,N_17324);
nor U20271 (N_20271,N_19451,N_16650);
nand U20272 (N_20272,N_15615,N_15052);
nor U20273 (N_20273,N_16166,N_15293);
or U20274 (N_20274,N_18862,N_15856);
and U20275 (N_20275,N_18009,N_19005);
nor U20276 (N_20276,N_18883,N_19754);
nor U20277 (N_20277,N_16038,N_16787);
xnor U20278 (N_20278,N_18275,N_16462);
xor U20279 (N_20279,N_18001,N_17413);
nor U20280 (N_20280,N_17114,N_17247);
and U20281 (N_20281,N_15585,N_19104);
nor U20282 (N_20282,N_19925,N_16402);
and U20283 (N_20283,N_16013,N_19249);
or U20284 (N_20284,N_19538,N_19369);
nand U20285 (N_20285,N_19281,N_16835);
nand U20286 (N_20286,N_15842,N_17192);
nand U20287 (N_20287,N_15113,N_16547);
and U20288 (N_20288,N_19920,N_16950);
and U20289 (N_20289,N_16371,N_16212);
xor U20290 (N_20290,N_16694,N_19170);
nand U20291 (N_20291,N_15965,N_18194);
or U20292 (N_20292,N_16123,N_19947);
or U20293 (N_20293,N_18511,N_17756);
nand U20294 (N_20294,N_17948,N_15150);
nor U20295 (N_20295,N_19080,N_17265);
and U20296 (N_20296,N_15261,N_15447);
xnor U20297 (N_20297,N_18169,N_19983);
xor U20298 (N_20298,N_15061,N_18724);
nand U20299 (N_20299,N_16294,N_17663);
nor U20300 (N_20300,N_18729,N_17500);
nor U20301 (N_20301,N_16869,N_16846);
or U20302 (N_20302,N_17467,N_19793);
xor U20303 (N_20303,N_19536,N_16487);
or U20304 (N_20304,N_19291,N_15154);
nor U20305 (N_20305,N_17932,N_19207);
or U20306 (N_20306,N_19858,N_18921);
or U20307 (N_20307,N_16093,N_17580);
or U20308 (N_20308,N_17535,N_16956);
nor U20309 (N_20309,N_15960,N_16720);
nor U20310 (N_20310,N_16753,N_19259);
nor U20311 (N_20311,N_19198,N_19189);
nand U20312 (N_20312,N_17659,N_16331);
nand U20313 (N_20313,N_15109,N_17825);
nand U20314 (N_20314,N_17953,N_16958);
nor U20315 (N_20315,N_17377,N_18177);
xor U20316 (N_20316,N_15040,N_17922);
nand U20317 (N_20317,N_17287,N_19658);
and U20318 (N_20318,N_16825,N_16429);
or U20319 (N_20319,N_16538,N_16536);
xor U20320 (N_20320,N_19863,N_16647);
or U20321 (N_20321,N_15185,N_17856);
nor U20322 (N_20322,N_16088,N_15017);
and U20323 (N_20323,N_16143,N_19949);
nand U20324 (N_20324,N_15297,N_15403);
nand U20325 (N_20325,N_17268,N_15673);
or U20326 (N_20326,N_17977,N_16282);
or U20327 (N_20327,N_17438,N_15059);
nor U20328 (N_20328,N_18614,N_15055);
nor U20329 (N_20329,N_19806,N_19826);
xor U20330 (N_20330,N_19390,N_15399);
nor U20331 (N_20331,N_19049,N_15008);
xor U20332 (N_20332,N_17253,N_15119);
or U20333 (N_20333,N_19282,N_18147);
xor U20334 (N_20334,N_17118,N_16736);
or U20335 (N_20335,N_18180,N_18898);
or U20336 (N_20336,N_17490,N_16742);
or U20337 (N_20337,N_19157,N_17738);
or U20338 (N_20338,N_17732,N_18096);
nand U20339 (N_20339,N_19573,N_16483);
nor U20340 (N_20340,N_19638,N_18600);
and U20341 (N_20341,N_17110,N_17494);
nand U20342 (N_20342,N_19053,N_17031);
or U20343 (N_20343,N_18022,N_19604);
or U20344 (N_20344,N_19912,N_19128);
xor U20345 (N_20345,N_17318,N_15728);
or U20346 (N_20346,N_16156,N_18162);
and U20347 (N_20347,N_17799,N_16511);
and U20348 (N_20348,N_15421,N_15797);
nor U20349 (N_20349,N_16730,N_15108);
nand U20350 (N_20350,N_15679,N_18968);
and U20351 (N_20351,N_17450,N_17025);
xnor U20352 (N_20352,N_16372,N_17211);
or U20353 (N_20353,N_19059,N_18960);
or U20354 (N_20354,N_17102,N_17543);
or U20355 (N_20355,N_17630,N_17860);
and U20356 (N_20356,N_19715,N_17677);
nor U20357 (N_20357,N_19628,N_15717);
and U20358 (N_20358,N_16831,N_18824);
and U20359 (N_20359,N_17341,N_18029);
xnor U20360 (N_20360,N_16296,N_19845);
or U20361 (N_20361,N_18881,N_17257);
nand U20362 (N_20362,N_16042,N_16448);
xnor U20363 (N_20363,N_18825,N_16284);
xor U20364 (N_20364,N_17648,N_17956);
or U20365 (N_20365,N_19201,N_18200);
nand U20366 (N_20366,N_17909,N_16921);
and U20367 (N_20367,N_17035,N_17602);
nand U20368 (N_20368,N_18459,N_19677);
xor U20369 (N_20369,N_16307,N_15825);
or U20370 (N_20370,N_15775,N_19453);
xor U20371 (N_20371,N_19701,N_19506);
or U20372 (N_20372,N_17373,N_18251);
xnor U20373 (N_20373,N_15544,N_19954);
xor U20374 (N_20374,N_16827,N_19073);
or U20375 (N_20375,N_18204,N_19105);
or U20376 (N_20376,N_16693,N_19403);
and U20377 (N_20377,N_16895,N_18939);
nor U20378 (N_20378,N_18728,N_15872);
xnor U20379 (N_20379,N_18533,N_19197);
xor U20380 (N_20380,N_18726,N_17503);
xnor U20381 (N_20381,N_18202,N_15164);
xnor U20382 (N_20382,N_17997,N_17662);
nand U20383 (N_20383,N_15385,N_16159);
and U20384 (N_20384,N_15902,N_16421);
or U20385 (N_20385,N_15051,N_16026);
and U20386 (N_20386,N_15060,N_19727);
nand U20387 (N_20387,N_16479,N_19371);
or U20388 (N_20388,N_18884,N_15433);
nor U20389 (N_20389,N_17927,N_18227);
or U20390 (N_20390,N_15759,N_19194);
nor U20391 (N_20391,N_19173,N_17571);
and U20392 (N_20392,N_17355,N_17104);
nor U20393 (N_20393,N_17005,N_17149);
and U20394 (N_20394,N_17370,N_17780);
xor U20395 (N_20395,N_19347,N_19132);
xnor U20396 (N_20396,N_19387,N_19409);
nor U20397 (N_20397,N_15201,N_15086);
nand U20398 (N_20398,N_15953,N_19723);
xnor U20399 (N_20399,N_16894,N_19366);
xor U20400 (N_20400,N_18212,N_15702);
nand U20401 (N_20401,N_19564,N_17819);
xor U20402 (N_20402,N_17336,N_19810);
nand U20403 (N_20403,N_17769,N_15651);
or U20404 (N_20404,N_19219,N_18297);
xor U20405 (N_20405,N_18562,N_15391);
nand U20406 (N_20406,N_15331,N_16513);
or U20407 (N_20407,N_18025,N_17255);
nand U20408 (N_20408,N_16726,N_19116);
nand U20409 (N_20409,N_18007,N_16820);
or U20410 (N_20410,N_19339,N_15687);
nand U20411 (N_20411,N_15198,N_15395);
nand U20412 (N_20412,N_15310,N_19622);
and U20413 (N_20413,N_15701,N_19256);
nand U20414 (N_20414,N_15021,N_15161);
nor U20415 (N_20415,N_19166,N_17091);
xnor U20416 (N_20416,N_16963,N_15866);
or U20417 (N_20417,N_15335,N_17258);
xnor U20418 (N_20418,N_16053,N_18913);
xnor U20419 (N_20419,N_17639,N_18900);
and U20420 (N_20420,N_15075,N_15193);
or U20421 (N_20421,N_15836,N_16148);
xnor U20422 (N_20422,N_16363,N_18343);
xnor U20423 (N_20423,N_16676,N_16279);
and U20424 (N_20424,N_15613,N_15423);
and U20425 (N_20425,N_17541,N_17729);
or U20426 (N_20426,N_16057,N_17224);
nand U20427 (N_20427,N_17509,N_15148);
xor U20428 (N_20428,N_16604,N_16181);
xor U20429 (N_20429,N_16315,N_19928);
nor U20430 (N_20430,N_17381,N_18084);
nor U20431 (N_20431,N_17674,N_16525);
xnor U20432 (N_20432,N_17361,N_18206);
nor U20433 (N_20433,N_16430,N_15941);
nand U20434 (N_20434,N_18821,N_19956);
nand U20435 (N_20435,N_19030,N_17471);
and U20436 (N_20436,N_17937,N_17410);
xnor U20437 (N_20437,N_18963,N_19936);
nor U20438 (N_20438,N_16286,N_15873);
nor U20439 (N_20439,N_19650,N_19343);
nand U20440 (N_20440,N_17760,N_15527);
and U20441 (N_20441,N_19266,N_18368);
and U20442 (N_20442,N_18111,N_15576);
nor U20443 (N_20443,N_19935,N_17949);
or U20444 (N_20444,N_17421,N_16327);
xor U20445 (N_20445,N_16882,N_15642);
or U20446 (N_20446,N_19924,N_16770);
and U20447 (N_20447,N_16721,N_19878);
nand U20448 (N_20448,N_19750,N_16591);
nor U20449 (N_20449,N_17686,N_19337);
nand U20450 (N_20450,N_19434,N_17613);
and U20451 (N_20451,N_15621,N_15087);
xnor U20452 (N_20452,N_17371,N_17954);
xor U20453 (N_20453,N_16099,N_19697);
nand U20454 (N_20454,N_17751,N_18571);
and U20455 (N_20455,N_19236,N_18378);
or U20456 (N_20456,N_18493,N_16761);
xnor U20457 (N_20457,N_15921,N_17216);
or U20458 (N_20458,N_19185,N_16619);
xor U20459 (N_20459,N_17704,N_17779);
and U20460 (N_20460,N_16086,N_15844);
or U20461 (N_20461,N_17564,N_19585);
nand U20462 (N_20462,N_19728,N_15157);
nor U20463 (N_20463,N_17787,N_17228);
xor U20464 (N_20464,N_18905,N_19652);
xnor U20465 (N_20465,N_18391,N_19321);
xnor U20466 (N_20466,N_16443,N_19997);
xor U20467 (N_20467,N_15574,N_17721);
and U20468 (N_20468,N_19277,N_17951);
nand U20469 (N_20469,N_18507,N_16110);
nor U20470 (N_20470,N_18238,N_16129);
nor U20471 (N_20471,N_18045,N_15816);
nand U20472 (N_20472,N_17730,N_19740);
nand U20473 (N_20473,N_18155,N_15307);
or U20474 (N_20474,N_18860,N_18872);
nor U20475 (N_20475,N_15504,N_17179);
nand U20476 (N_20476,N_16117,N_17453);
and U20477 (N_20477,N_18468,N_19922);
nor U20478 (N_20478,N_15822,N_19846);
and U20479 (N_20479,N_15422,N_15439);
and U20480 (N_20480,N_15614,N_18210);
or U20481 (N_20481,N_18259,N_16695);
xor U20482 (N_20482,N_15804,N_17556);
xor U20483 (N_20483,N_18659,N_19636);
or U20484 (N_20484,N_19098,N_16698);
nand U20485 (N_20485,N_15436,N_17971);
nor U20486 (N_20486,N_17002,N_15512);
and U20487 (N_20487,N_15151,N_19115);
nor U20488 (N_20488,N_17831,N_16396);
xor U20489 (N_20489,N_17957,N_18330);
xnor U20490 (N_20490,N_17394,N_16087);
and U20491 (N_20491,N_16999,N_17282);
nand U20492 (N_20492,N_16990,N_16367);
nand U20493 (N_20493,N_16582,N_15380);
or U20494 (N_20494,N_16218,N_17788);
xnor U20495 (N_20495,N_17357,N_18805);
xnor U20496 (N_20496,N_16790,N_16424);
nand U20497 (N_20497,N_15712,N_15995);
and U20498 (N_20498,N_17766,N_15684);
xnor U20499 (N_20499,N_18365,N_15525);
or U20500 (N_20500,N_19452,N_17122);
xnor U20501 (N_20501,N_18440,N_16929);
nor U20502 (N_20502,N_17472,N_18912);
nor U20503 (N_20503,N_17640,N_17143);
nor U20504 (N_20504,N_15911,N_19180);
xor U20505 (N_20505,N_19957,N_17319);
or U20506 (N_20506,N_17933,N_15971);
nor U20507 (N_20507,N_16173,N_16116);
xnor U20508 (N_20508,N_15617,N_16955);
nand U20509 (N_20509,N_17213,N_19887);
nor U20510 (N_20510,N_19315,N_18432);
or U20511 (N_20511,N_16005,N_18803);
xnor U20512 (N_20512,N_18976,N_19958);
xor U20513 (N_20513,N_19823,N_17020);
nor U20514 (N_20514,N_15987,N_19749);
nor U20515 (N_20515,N_16194,N_16804);
and U20516 (N_20516,N_17899,N_19654);
xnor U20517 (N_20517,N_16004,N_19605);
nand U20518 (N_20518,N_17810,N_17189);
and U20519 (N_20519,N_16436,N_19868);
nor U20520 (N_20520,N_19865,N_15486);
xnor U20521 (N_20521,N_16158,N_19804);
nor U20522 (N_20522,N_15410,N_15599);
or U20523 (N_20523,N_18051,N_17137);
xnor U20524 (N_20524,N_16079,N_16617);
xor U20525 (N_20525,N_17702,N_16641);
nand U20526 (N_20526,N_19220,N_18027);
and U20527 (N_20527,N_15707,N_15864);
nand U20528 (N_20528,N_18063,N_17232);
xnor U20529 (N_20529,N_17790,N_19146);
xor U20530 (N_20530,N_17941,N_18986);
nand U20531 (N_20531,N_16621,N_15159);
and U20532 (N_20532,N_17085,N_19319);
nand U20533 (N_20533,N_19288,N_18226);
xnor U20534 (N_20534,N_16444,N_15233);
and U20535 (N_20535,N_18612,N_19439);
and U20536 (N_20536,N_16733,N_15139);
xor U20537 (N_20537,N_15875,N_16272);
nand U20538 (N_20538,N_19397,N_18082);
or U20539 (N_20539,N_16725,N_17151);
nand U20540 (N_20540,N_15056,N_16035);
and U20541 (N_20541,N_18703,N_16322);
or U20542 (N_20542,N_17607,N_17162);
nand U20543 (N_20543,N_19927,N_17468);
xor U20544 (N_20544,N_15513,N_15793);
nor U20545 (N_20545,N_18118,N_19916);
or U20546 (N_20546,N_15327,N_16204);
nor U20547 (N_20547,N_16505,N_18651);
xor U20548 (N_20548,N_19187,N_18088);
nand U20549 (N_20549,N_17222,N_15539);
nor U20550 (N_20550,N_16537,N_16931);
nor U20551 (N_20551,N_17631,N_16222);
nor U20552 (N_20552,N_18042,N_19276);
and U20553 (N_20553,N_17343,N_15023);
nand U20554 (N_20554,N_17540,N_15738);
or U20555 (N_20555,N_15498,N_17901);
xnor U20556 (N_20556,N_17507,N_18284);
nor U20557 (N_20557,N_15354,N_17150);
and U20558 (N_20558,N_17593,N_15039);
xnor U20559 (N_20559,N_19050,N_17749);
and U20560 (N_20560,N_18064,N_19426);
nor U20561 (N_20561,N_19511,N_15133);
and U20562 (N_20562,N_15531,N_17254);
and U20563 (N_20563,N_17891,N_18583);
or U20564 (N_20564,N_16653,N_18306);
xnor U20565 (N_20565,N_17942,N_17214);
nand U20566 (N_20566,N_16597,N_17975);
nor U20567 (N_20567,N_15449,N_16876);
xnor U20568 (N_20568,N_18397,N_18094);
xor U20569 (N_20569,N_16899,N_15857);
or U20570 (N_20570,N_18292,N_15007);
nand U20571 (N_20571,N_19257,N_19345);
nand U20572 (N_20572,N_18028,N_19248);
nand U20573 (N_20573,N_18193,N_19108);
and U20574 (N_20574,N_18097,N_15935);
or U20575 (N_20575,N_15360,N_17547);
or U20576 (N_20576,N_19890,N_15913);
nand U20577 (N_20577,N_15110,N_19825);
or U20578 (N_20578,N_18736,N_19472);
and U20579 (N_20579,N_16384,N_19088);
xor U20580 (N_20580,N_18807,N_16237);
and U20581 (N_20581,N_18106,N_19526);
nand U20582 (N_20582,N_18462,N_16283);
and U20583 (N_20583,N_19094,N_19933);
nand U20584 (N_20584,N_19460,N_19327);
or U20585 (N_20585,N_15710,N_15358);
and U20586 (N_20586,N_17171,N_18231);
or U20587 (N_20587,N_17890,N_16821);
or U20588 (N_20588,N_17299,N_16340);
nor U20589 (N_20589,N_15211,N_18151);
nand U20590 (N_20590,N_19678,N_18568);
or U20591 (N_20591,N_18741,N_15253);
xor U20592 (N_20592,N_19270,N_19074);
nor U20593 (N_20593,N_15379,N_17824);
nor U20594 (N_20594,N_18797,N_19174);
xnor U20595 (N_20595,N_18222,N_17868);
xor U20596 (N_20596,N_19885,N_16915);
and U20597 (N_20597,N_18964,N_15523);
xnor U20598 (N_20598,N_15697,N_16834);
xor U20599 (N_20599,N_18542,N_15916);
and U20600 (N_20600,N_15922,N_15833);
nand U20601 (N_20601,N_17670,N_19328);
and U20602 (N_20602,N_19642,N_17335);
nor U20603 (N_20603,N_18919,N_15862);
nor U20604 (N_20604,N_15565,N_18486);
and U20605 (N_20605,N_16715,N_19633);
and U20606 (N_20606,N_15275,N_19898);
and U20607 (N_20607,N_18289,N_16219);
and U20608 (N_20608,N_17866,N_16151);
nand U20609 (N_20609,N_18358,N_17281);
xnor U20610 (N_20610,N_16993,N_16015);
and U20611 (N_20611,N_17325,N_15994);
or U20612 (N_20612,N_17995,N_18078);
nand U20613 (N_20613,N_17350,N_16637);
xor U20614 (N_20614,N_16938,N_15752);
nor U20615 (N_20615,N_15606,N_15386);
and U20616 (N_20616,N_17627,N_15732);
and U20617 (N_20617,N_18035,N_16145);
xor U20618 (N_20618,N_17781,N_17392);
nand U20619 (N_20619,N_15915,N_16051);
nand U20620 (N_20620,N_15062,N_18798);
and U20621 (N_20621,N_18937,N_15672);
and U20622 (N_20622,N_16492,N_18870);
nand U20623 (N_20623,N_16532,N_16064);
and U20624 (N_20624,N_16313,N_17502);
nor U20625 (N_20625,N_18801,N_15442);
xor U20626 (N_20626,N_15776,N_17078);
nor U20627 (N_20627,N_15591,N_18972);
xnor U20628 (N_20628,N_16393,N_18957);
xor U20629 (N_20629,N_15859,N_17036);
nand U20630 (N_20630,N_15126,N_16919);
and U20631 (N_20631,N_16791,N_19314);
xnor U20632 (N_20632,N_16388,N_19953);
nor U20633 (N_20633,N_18951,N_18332);
or U20634 (N_20634,N_17419,N_18421);
or U20635 (N_20635,N_17420,N_15883);
nand U20636 (N_20636,N_19177,N_15102);
and U20637 (N_20637,N_18781,N_19725);
nand U20638 (N_20638,N_19700,N_16438);
or U20639 (N_20639,N_16815,N_17996);
nor U20640 (N_20640,N_18650,N_18832);
nor U20641 (N_20641,N_18775,N_15231);
nor U20642 (N_20642,N_18406,N_17399);
nor U20643 (N_20643,N_16334,N_17464);
nor U20644 (N_20644,N_16987,N_17442);
nor U20645 (N_20645,N_16056,N_19338);
xor U20646 (N_20646,N_19761,N_19738);
nand U20647 (N_20647,N_18116,N_19505);
and U20648 (N_20648,N_17965,N_17140);
nand U20649 (N_20649,N_15299,N_16364);
and U20650 (N_20650,N_15861,N_18229);
or U20651 (N_20651,N_17796,N_15740);
nand U20652 (N_20652,N_19995,N_17970);
nor U20653 (N_20653,N_16808,N_18080);
nor U20654 (N_20654,N_19103,N_16874);
and U20655 (N_20655,N_18508,N_17551);
nand U20656 (N_20656,N_18613,N_15477);
xnor U20657 (N_20657,N_15036,N_19161);
nor U20658 (N_20658,N_16127,N_17458);
or U20659 (N_20659,N_15983,N_19129);
nor U20660 (N_20660,N_19079,N_17622);
nand U20661 (N_20661,N_15924,N_15188);
nor U20662 (N_20662,N_18718,N_15194);
or U20663 (N_20663,N_15376,N_15508);
nor U20664 (N_20664,N_16959,N_16670);
nand U20665 (N_20665,N_17221,N_15366);
nand U20666 (N_20666,N_15041,N_15727);
xor U20667 (N_20667,N_17434,N_16972);
nor U20668 (N_20668,N_19559,N_19041);
nor U20669 (N_20669,N_18276,N_19608);
and U20670 (N_20670,N_15073,N_15781);
nor U20671 (N_20671,N_17513,N_18945);
nand U20672 (N_20672,N_17112,N_17519);
nor U20673 (N_20673,N_17574,N_16493);
nor U20674 (N_20674,N_17404,N_16101);
nand U20675 (N_20675,N_18171,N_15414);
and U20676 (N_20676,N_18436,N_16636);
or U20677 (N_20677,N_16339,N_15719);
xor U20678 (N_20678,N_16699,N_15598);
nor U20679 (N_20679,N_19616,N_17158);
and U20680 (N_20680,N_17042,N_17161);
nand U20681 (N_20681,N_19599,N_17339);
and U20682 (N_20682,N_19341,N_17798);
and U20683 (N_20683,N_16523,N_16664);
or U20684 (N_20684,N_19938,N_15344);
nor U20685 (N_20685,N_19156,N_19023);
nor U20686 (N_20686,N_19841,N_15070);
xor U20687 (N_20687,N_16612,N_16943);
or U20688 (N_20688,N_19556,N_19597);
xnor U20689 (N_20689,N_15782,N_19551);
xor U20690 (N_20690,N_15917,N_16263);
or U20691 (N_20691,N_18033,N_18897);
nand U20692 (N_20692,N_17009,N_16442);
nor U20693 (N_20693,N_18548,N_18577);
xnor U20694 (N_20694,N_18010,N_16277);
or U20695 (N_20695,N_19745,N_18757);
or U20696 (N_20696,N_15938,N_17988);
and U20697 (N_20697,N_19518,N_17136);
nand U20698 (N_20698,N_18624,N_15901);
and U20699 (N_20699,N_17146,N_16864);
nand U20700 (N_20700,N_18224,N_17986);
nand U20701 (N_20701,N_17955,N_18211);
and U20702 (N_20702,N_16274,N_17981);
xor U20703 (N_20703,N_18257,N_16623);
or U20704 (N_20704,N_17328,N_15237);
or U20705 (N_20705,N_15948,N_18091);
and U20706 (N_20706,N_19557,N_18780);
xor U20707 (N_20707,N_19686,N_16799);
xnor U20708 (N_20708,N_17040,N_15886);
nor U20709 (N_20709,N_15823,N_16729);
and U20710 (N_20710,N_18382,N_17835);
and U20711 (N_20711,N_18434,N_19492);
nor U20712 (N_20712,N_17848,N_17950);
nand U20713 (N_20713,N_19334,N_16489);
nand U20714 (N_20714,N_16318,N_17074);
or U20715 (N_20715,N_18733,N_16839);
xnor U20716 (N_20716,N_17069,N_18623);
nor U20717 (N_20717,N_18412,N_16517);
xnor U20718 (N_20718,N_18400,N_15803);
nor U20719 (N_20719,N_17426,N_15956);
xor U20720 (N_20720,N_16365,N_16744);
and U20721 (N_20721,N_17200,N_17207);
or U20722 (N_20722,N_17185,N_18740);
xor U20723 (N_20723,N_19442,N_15808);
and U20724 (N_20724,N_19833,N_15649);
nor U20725 (N_20725,N_15790,N_16691);
or U20726 (N_20726,N_18896,N_17958);
nor U20727 (N_20727,N_18015,N_16709);
or U20728 (N_20728,N_18126,N_19930);
nand U20729 (N_20729,N_15879,N_18791);
nand U20730 (N_20730,N_18580,N_19908);
and U20731 (N_20731,N_19617,N_19095);
xor U20732 (N_20732,N_16875,N_17378);
and U20733 (N_20733,N_18089,N_18535);
nor U20734 (N_20734,N_15528,N_18302);
xor U20735 (N_20735,N_17244,N_17225);
and U20736 (N_20736,N_15943,N_16316);
xnor U20737 (N_20737,N_18674,N_18386);
nand U20738 (N_20738,N_18667,N_19592);
and U20739 (N_20739,N_19703,N_16957);
xor U20740 (N_20740,N_15357,N_15025);
nand U20741 (N_20741,N_16638,N_19044);
and U20742 (N_20742,N_15003,N_19768);
xor U20743 (N_20743,N_15031,N_16163);
nand U20744 (N_20744,N_16518,N_15400);
nand U20745 (N_20745,N_15158,N_15455);
xor U20746 (N_20746,N_16764,N_17625);
or U20747 (N_20747,N_15634,N_15648);
or U20748 (N_20748,N_18867,N_16600);
nor U20749 (N_20749,N_18808,N_16215);
nor U20750 (N_20750,N_18176,N_18388);
nor U20751 (N_20751,N_15190,N_15572);
xor U20752 (N_20752,N_15394,N_18593);
nor U20753 (N_20753,N_16754,N_16007);
or U20754 (N_20754,N_15019,N_17011);
nand U20755 (N_20755,N_16927,N_15104);
or U20756 (N_20756,N_16806,N_18460);
nand U20757 (N_20757,N_15419,N_16270);
xor U20758 (N_20758,N_17415,N_17582);
or U20759 (N_20759,N_18020,N_16616);
nand U20760 (N_20760,N_15693,N_17550);
nor U20761 (N_20761,N_15115,N_18903);
and U20762 (N_20762,N_19286,N_18115);
nor U20763 (N_20763,N_15372,N_17245);
nand U20764 (N_20764,N_18607,N_18447);
or U20765 (N_20765,N_17007,N_17863);
xnor U20766 (N_20766,N_17923,N_15053);
nor U20767 (N_20767,N_16055,N_17617);
or U20768 (N_20768,N_19463,N_18906);
and U20769 (N_20769,N_18753,N_17621);
and U20770 (N_20770,N_16481,N_17363);
or U20771 (N_20771,N_19311,N_18002);
or U20772 (N_20772,N_19303,N_18285);
nand U20773 (N_20773,N_16146,N_19644);
xnor U20774 (N_20774,N_15078,N_15645);
or U20775 (N_20775,N_19627,N_17858);
or U20776 (N_20776,N_18917,N_16668);
xor U20777 (N_20777,N_16361,N_16112);
nor U20778 (N_20778,N_16047,N_18140);
and U20779 (N_20779,N_15050,N_19917);
and U20780 (N_20780,N_16666,N_18989);
and U20781 (N_20781,N_18280,N_16223);
or U20782 (N_20782,N_19469,N_19163);
nand U20783 (N_20783,N_16587,N_17510);
or U20784 (N_20784,N_16757,N_17095);
or U20785 (N_20785,N_15851,N_15999);
nand U20786 (N_20786,N_19532,N_18931);
or U20787 (N_20787,N_17673,N_19448);
xnor U20788 (N_20788,N_19051,N_18809);
nand U20789 (N_20789,N_19375,N_15227);
nor U20790 (N_20790,N_19687,N_15478);
or U20791 (N_20791,N_17604,N_18454);
and U20792 (N_20792,N_18759,N_17794);
xor U20793 (N_20793,N_15349,N_15802);
or U20794 (N_20794,N_18243,N_18617);
nor U20795 (N_20795,N_17877,N_16826);
nand U20796 (N_20796,N_19284,N_17567);
xnor U20797 (N_20797,N_18599,N_15996);
or U20798 (N_20798,N_15213,N_16063);
nor U20799 (N_20799,N_19577,N_19234);
nand U20800 (N_20800,N_16464,N_15934);
xor U20801 (N_20801,N_16473,N_19100);
nor U20802 (N_20802,N_15992,N_16748);
or U20803 (N_20803,N_15266,N_15855);
nor U20804 (N_20804,N_18991,N_19664);
and U20805 (N_20805,N_18510,N_15566);
or U20806 (N_20806,N_16009,N_19247);
nand U20807 (N_20807,N_15852,N_19822);
xor U20808 (N_20808,N_19164,N_18055);
or U20809 (N_20809,N_17531,N_18769);
nand U20810 (N_20810,N_18457,N_19698);
and U20811 (N_20811,N_17530,N_15320);
xor U20812 (N_20812,N_19117,N_18301);
nand U20813 (N_20813,N_18878,N_16075);
and U20814 (N_20814,N_19647,N_18428);
nor U20815 (N_20815,N_16644,N_17286);
xnor U20816 (N_20816,N_17353,N_16998);
nand U20817 (N_20817,N_19776,N_17773);
or U20818 (N_20818,N_16347,N_18248);
nor U20819 (N_20819,N_15092,N_17557);
and U20820 (N_20820,N_16392,N_17612);
nand U20821 (N_20821,N_17422,N_16375);
xnor U20822 (N_20822,N_16803,N_19431);
or U20823 (N_20823,N_18417,N_17235);
or U20824 (N_20824,N_15704,N_16276);
nand U20825 (N_20825,N_16651,N_18688);
or U20826 (N_20826,N_19716,N_15669);
xor U20827 (N_20827,N_17477,N_15874);
nand U20828 (N_20828,N_16717,N_16349);
and U20829 (N_20829,N_16971,N_18207);
or U20830 (N_20830,N_18999,N_15287);
xnor U20831 (N_20831,N_18974,N_15097);
and U20832 (N_20832,N_16478,N_16480);
and U20833 (N_20833,N_18578,N_18219);
and U20834 (N_20834,N_18165,N_19587);
or U20835 (N_20835,N_16701,N_15068);
and U20836 (N_20836,N_17097,N_18841);
nor U20837 (N_20837,N_18398,N_15127);
nor U20838 (N_20838,N_18990,N_18074);
xor U20839 (N_20839,N_16601,N_15316);
xnor U20840 (N_20840,N_19612,N_18671);
or U20841 (N_20841,N_17000,N_16702);
or U20842 (N_20842,N_16805,N_16789);
nor U20843 (N_20843,N_19061,N_19020);
xor U20844 (N_20844,N_16838,N_16552);
nand U20845 (N_20845,N_16273,N_17812);
xnor U20846 (N_20846,N_16649,N_17618);
nand U20847 (N_20847,N_17345,N_17006);
nor U20848 (N_20848,N_19741,N_18992);
or U20849 (N_20849,N_18818,N_17741);
and U20850 (N_20850,N_16100,N_16954);
and U20851 (N_20851,N_18504,N_15474);
nor U20852 (N_20852,N_18970,N_18656);
nor U20853 (N_20853,N_19799,N_16377);
xor U20854 (N_20854,N_19075,N_19609);
and U20855 (N_20855,N_15680,N_17679);
nor U20856 (N_20856,N_17298,N_19842);
nor U20857 (N_20857,N_16661,N_16024);
and U20858 (N_20858,N_18558,N_15698);
xor U20859 (N_20859,N_18643,N_16139);
and U20860 (N_20860,N_16841,N_19619);
or U20861 (N_20861,N_19244,N_18479);
nor U20862 (N_20862,N_15342,N_17963);
or U20863 (N_20863,N_16629,N_15296);
and U20864 (N_20864,N_15168,N_19540);
xor U20865 (N_20865,N_15632,N_18360);
or U20866 (N_20866,N_18307,N_15865);
and U20867 (N_20867,N_15800,N_19379);
nand U20868 (N_20868,N_19834,N_17959);
or U20869 (N_20869,N_17559,N_18217);
or U20870 (N_20870,N_19689,N_16951);
or U20871 (N_20871,N_18836,N_18755);
xnor U20872 (N_20872,N_17315,N_17387);
nand U20873 (N_20873,N_16271,N_19572);
xor U20874 (N_20874,N_19550,N_19297);
nor U20875 (N_20875,N_17238,N_16935);
and U20876 (N_20876,N_19847,N_19870);
nor U20877 (N_20877,N_17183,N_17821);
nand U20878 (N_20878,N_15564,N_15322);
and U20879 (N_20879,N_18172,N_16141);
xor U20880 (N_20880,N_18700,N_16255);
nor U20881 (N_20881,N_17940,N_17366);
nor U20882 (N_20882,N_19762,N_17164);
nor U20883 (N_20883,N_15428,N_15460);
xor U20884 (N_20884,N_19242,N_15440);
nor U20885 (N_20885,N_19904,N_17333);
xor U20886 (N_20886,N_15771,N_15502);
nand U20887 (N_20887,N_18586,N_17092);
and U20888 (N_20888,N_18823,N_15136);
nand U20889 (N_20889,N_16514,N_19153);
nand U20890 (N_20890,N_16541,N_15485);
nand U20891 (N_20891,N_16584,N_16216);
and U20892 (N_20892,N_17524,N_18293);
xor U20893 (N_20893,N_18152,N_15176);
nand U20894 (N_20894,N_16469,N_18527);
nor U20895 (N_20895,N_18488,N_19243);
and U20896 (N_20896,N_16061,N_17553);
nand U20897 (N_20897,N_19832,N_16266);
xor U20898 (N_20898,N_17424,N_18885);
nand U20899 (N_20899,N_19795,N_16039);
nor U20900 (N_20900,N_18058,N_19718);
xnor U20901 (N_20901,N_19861,N_19158);
and U20902 (N_20902,N_15945,N_15604);
or U20903 (N_20903,N_16497,N_17765);
nor U20904 (N_20904,N_16423,N_17271);
xnor U20905 (N_20905,N_19412,N_17696);
xor U20906 (N_20906,N_15177,N_16230);
xnor U20907 (N_20907,N_18966,N_16837);
nor U20908 (N_20908,N_17060,N_15072);
nand U20909 (N_20909,N_16540,N_16157);
or U20910 (N_20910,N_18902,N_17504);
and U20911 (N_20911,N_15660,N_16673);
or U20912 (N_20912,N_17052,N_15000);
nor U20913 (N_20913,N_17212,N_19362);
xnor U20914 (N_20914,N_17013,N_18121);
and U20915 (N_20915,N_15255,N_17113);
nor U20916 (N_20916,N_16774,N_15112);
or U20917 (N_20917,N_16548,N_19736);
nor U20918 (N_20918,N_16578,N_19123);
xor U20919 (N_20919,N_16368,N_17283);
and U20920 (N_20920,N_16091,N_17698);
and U20921 (N_20921,N_17762,N_15277);
nor U20922 (N_20922,N_17041,N_19415);
nor U20923 (N_20923,N_16847,N_16490);
or U20924 (N_20924,N_15510,N_18591);
and U20925 (N_20925,N_16355,N_16238);
and U20926 (N_20926,N_16672,N_17728);
xor U20927 (N_20927,N_18863,N_17352);
nand U20928 (N_20928,N_18777,N_15796);
xor U20929 (N_20929,N_15812,N_18286);
nand U20930 (N_20930,N_16221,N_19432);
and U20931 (N_20931,N_19033,N_18924);
nor U20932 (N_20932,N_19293,N_18467);
nor U20933 (N_20933,N_15974,N_17208);
or U20934 (N_20934,N_15393,N_16870);
or U20935 (N_20935,N_16904,N_16745);
xnor U20936 (N_20936,N_18829,N_17752);
and U20937 (N_20937,N_15235,N_19503);
nand U20938 (N_20938,N_19255,N_17990);
and U20939 (N_20939,N_16289,N_19481);
xnor U20940 (N_20940,N_15111,N_16455);
nand U20941 (N_20941,N_17437,N_18827);
xnor U20942 (N_20942,N_18901,N_18167);
or U20943 (N_20943,N_19214,N_15891);
nand U20944 (N_20944,N_16106,N_15656);
and U20945 (N_20945,N_18654,N_17497);
nor U20946 (N_20946,N_17408,N_17383);
or U20947 (N_20947,N_18340,N_16241);
xor U20948 (N_20948,N_16560,N_15970);
and U20949 (N_20949,N_18696,N_18526);
xor U20950 (N_20950,N_17276,N_19886);
and U20951 (N_20951,N_15784,N_18166);
or U20952 (N_20952,N_16342,N_15280);
nand U20953 (N_20953,N_18270,N_16872);
and U20954 (N_20954,N_19417,N_16453);
nor U20955 (N_20955,N_17087,N_17130);
and U20956 (N_20956,N_16692,N_18629);
or U20957 (N_20957,N_17684,N_18043);
nand U20958 (N_20958,N_18725,N_19063);
nand U20959 (N_20959,N_15069,N_16524);
nor U20960 (N_20960,N_18681,N_18461);
nand U20961 (N_20961,N_18416,N_17223);
and U20962 (N_20962,N_15807,N_17634);
xor U20963 (N_20963,N_15863,N_17943);
nor U20964 (N_20964,N_16000,N_18734);
nor U20965 (N_20965,N_16937,N_17289);
xnor U20966 (N_20966,N_15735,N_15519);
and U20967 (N_20967,N_18814,N_16317);
nand U20968 (N_20968,N_19208,N_19651);
xor U20969 (N_20969,N_18018,N_16539);
or U20970 (N_20970,N_18129,N_15251);
nor U20971 (N_20971,N_17646,N_16763);
nor U20972 (N_20972,N_16457,N_16357);
nand U20973 (N_20973,N_15026,N_18287);
xnor U20974 (N_20974,N_16862,N_17826);
and U20975 (N_20975,N_17059,N_15638);
and U20976 (N_20976,N_18429,N_19751);
nand U20977 (N_20977,N_15706,N_16575);
xnor U20978 (N_20978,N_16121,N_16369);
nor U20979 (N_20979,N_19660,N_18437);
or U20980 (N_20980,N_18146,N_18920);
xnor U20981 (N_20981,N_17376,N_18868);
xnor U20982 (N_20982,N_18751,N_17288);
and U20983 (N_20983,N_16287,N_19774);
nor U20984 (N_20984,N_17960,N_18882);
nand U20985 (N_20985,N_19394,N_16708);
xnor U20986 (N_20986,N_19884,N_18719);
or U20987 (N_20987,N_19488,N_16058);
nor U20988 (N_20988,N_18888,N_19964);
nor U20989 (N_20989,N_15636,N_17657);
nand U20990 (N_20990,N_15121,N_15593);
and U20991 (N_20991,N_18337,N_15757);
or U20992 (N_20992,N_17649,N_16994);
and U20993 (N_20993,N_19665,N_17874);
nor U20994 (N_20994,N_17256,N_16885);
and U20995 (N_20995,N_16983,N_17726);
nand U20996 (N_20996,N_17578,N_17470);
xor U20997 (N_20997,N_18349,N_18145);
or U20998 (N_20998,N_15076,N_17038);
nor U20999 (N_20999,N_15631,N_15694);
nand U21000 (N_21000,N_15083,N_17791);
nor U21001 (N_21001,N_17120,N_15561);
or U21002 (N_21002,N_18404,N_15841);
nor U21003 (N_21003,N_18239,N_16596);
xor U21004 (N_21004,N_19570,N_16203);
nor U21005 (N_21005,N_19008,N_17813);
and U21006 (N_21006,N_17338,N_17735);
and U21007 (N_21007,N_15579,N_19336);
xnor U21008 (N_21008,N_19940,N_18059);
and U21009 (N_21009,N_15124,N_19553);
or U21010 (N_21010,N_15187,N_15756);
xnor U21011 (N_21011,N_16705,N_17689);
xnor U21012 (N_21012,N_16866,N_18620);
or U21013 (N_21013,N_16706,N_18414);
and U21014 (N_21014,N_16484,N_15737);
xor U21015 (N_21015,N_17926,N_17884);
xnor U21016 (N_21016,N_19583,N_16164);
nand U21017 (N_21017,N_19977,N_16114);
or U21018 (N_21018,N_19568,N_17448);
nand U21019 (N_21019,N_16880,N_17515);
nand U21020 (N_21020,N_15288,N_15780);
nor U21021 (N_21021,N_19821,N_16985);
nor U21022 (N_21022,N_16814,N_16948);
or U21023 (N_21023,N_15274,N_18081);
nor U21024 (N_21024,N_16054,N_15088);
nor U21025 (N_21025,N_17175,N_16782);
nand U21026 (N_21026,N_19959,N_18005);
or U21027 (N_21027,N_17480,N_16267);
xor U21028 (N_21028,N_17417,N_16312);
xnor U21029 (N_21029,N_18738,N_15551);
nand U21030 (N_21030,N_15223,N_16798);
or U21031 (N_21031,N_15721,N_17710);
xnor U21032 (N_21032,N_17718,N_17193);
nor U21033 (N_21033,N_16134,N_17251);
nor U21034 (N_21034,N_18377,N_18852);
xnor U21035 (N_21035,N_16546,N_16562);
xor U21036 (N_21036,N_18016,N_18984);
or U21037 (N_21037,N_16346,N_18540);
and U21038 (N_21038,N_17865,N_19598);
or U21039 (N_21039,N_17945,N_15806);
nor U21040 (N_21040,N_17852,N_16633);
nor U21041 (N_21041,N_18636,N_19475);
or U21042 (N_21042,N_16992,N_19530);
nand U21043 (N_21043,N_15839,N_15469);
or U21044 (N_21044,N_15220,N_16328);
nand U21045 (N_21045,N_19630,N_17243);
nand U21046 (N_21046,N_15548,N_17629);
nor U21047 (N_21047,N_15029,N_19302);
and U21048 (N_21048,N_15145,N_16996);
or U21049 (N_21049,N_18709,N_16752);
or U21050 (N_21050,N_19210,N_15910);
nand U21051 (N_21051,N_19788,N_15270);
or U21052 (N_21052,N_15325,N_16586);
nand U21053 (N_21053,N_19203,N_17144);
nor U21054 (N_21054,N_19639,N_15885);
nand U21055 (N_21055,N_18424,N_16707);
or U21056 (N_21056,N_18735,N_17903);
xor U21057 (N_21057,N_19864,N_16968);
xnor U21058 (N_21058,N_16197,N_18547);
xnor U21059 (N_21059,N_18936,N_19545);
xor U21060 (N_21060,N_19848,N_16078);
nor U21061 (N_21061,N_15383,N_18157);
nand U21062 (N_21062,N_19895,N_15744);
nor U21063 (N_21063,N_19001,N_18859);
and U21064 (N_21064,N_15683,N_17217);
xor U21065 (N_21065,N_15832,N_17529);
nor U21066 (N_21066,N_18014,N_19112);
nand U21067 (N_21067,N_17433,N_18036);
and U21068 (N_21068,N_16737,N_15259);
xor U21069 (N_21069,N_15785,N_18969);
and U21070 (N_21070,N_16153,N_17620);
or U21071 (N_21071,N_19085,N_19025);
xor U21072 (N_21072,N_16809,N_17445);
nand U21073 (N_21073,N_17374,N_18288);
nor U21074 (N_21074,N_17001,N_18137);
or U21075 (N_21075,N_15925,N_15647);
nand U21076 (N_21076,N_17215,N_16750);
xor U21077 (N_21077,N_15281,N_18188);
and U21078 (N_21078,N_15207,N_19466);
nand U21079 (N_21079,N_17579,N_17126);
xor U21080 (N_21080,N_15165,N_17053);
xor U21081 (N_21081,N_16759,N_15415);
nor U21082 (N_21082,N_17772,N_15409);
xnor U21083 (N_21083,N_17280,N_18866);
nand U21084 (N_21084,N_19013,N_18104);
nand U21085 (N_21085,N_16571,N_18864);
or U21086 (N_21086,N_15064,N_19383);
or U21087 (N_21087,N_19066,N_15899);
and U21088 (N_21088,N_19855,N_19478);
nand U21089 (N_21089,N_18708,N_17930);
nand U21090 (N_21090,N_16995,N_18748);
and U21091 (N_21091,N_19418,N_17653);
nand U21092 (N_21092,N_19141,N_19235);
and U21093 (N_21093,N_19360,N_17917);
xor U21094 (N_21094,N_17037,N_18843);
nand U21095 (N_21095,N_16202,N_17576);
nor U21096 (N_21096,N_17716,N_17388);
and U21097 (N_21097,N_16390,N_16264);
or U21098 (N_21098,N_19118,N_19783);
or U21099 (N_21099,N_18907,N_19114);
nand U21100 (N_21100,N_17520,N_15741);
and U21101 (N_21101,N_17859,N_16234);
xor U21102 (N_21102,N_19596,N_18254);
nand U21103 (N_21103,N_19625,N_17443);
xor U21104 (N_21104,N_19332,N_15206);
and U21105 (N_21105,N_17978,N_17692);
or U21106 (N_21106,N_15536,N_16683);
or U21107 (N_21107,N_18154,N_19427);
nand U21108 (N_21108,N_17482,N_19871);
xor U21109 (N_21109,N_17139,N_19428);
nand U21110 (N_21110,N_16254,N_19892);
or U21111 (N_21111,N_15079,N_17740);
xnor U21112 (N_21112,N_17455,N_19195);
nor U21113 (N_21113,N_18850,N_18609);
or U21114 (N_21114,N_18618,N_17488);
nand U21115 (N_21115,N_17173,N_19186);
and U21116 (N_21116,N_18749,N_15609);
nand U21117 (N_21117,N_17685,N_15272);
or U21118 (N_21118,N_18072,N_16415);
nor U21119 (N_21119,N_15089,N_18465);
or U21120 (N_21120,N_16046,N_15550);
nand U21121 (N_21121,N_17236,N_16251);
xor U21122 (N_21122,N_19012,N_15208);
and U21123 (N_21123,N_19065,N_15276);
nor U21124 (N_21124,N_18536,N_16984);
nor U21125 (N_21125,N_17168,N_17661);
or U21126 (N_21126,N_19708,N_17125);
or U21127 (N_21127,N_15571,N_18451);
nand U21128 (N_21128,N_18834,N_18105);
xnor U21129 (N_21129,N_19730,N_16566);
and U21130 (N_21130,N_16350,N_17512);
xor U21131 (N_21131,N_19087,N_15612);
xor U21132 (N_21132,N_15982,N_16292);
nor U21133 (N_21133,N_19222,N_15312);
and U21134 (N_21134,N_16131,N_15547);
nand U21135 (N_21135,N_16811,N_18258);
xnor U21136 (N_21136,N_15726,N_18309);
nor U21137 (N_21137,N_19204,N_19484);
or U21138 (N_21138,N_18687,N_19712);
nor U21139 (N_21139,N_17527,N_17784);
nor U21140 (N_21140,N_19393,N_16413);
nand U21141 (N_21141,N_17439,N_18544);
and U21142 (N_21142,N_15792,N_19407);
and U21143 (N_21143,N_17521,N_19803);
or U21144 (N_21144,N_15313,N_17895);
nand U21145 (N_21145,N_19040,N_18876);
xor U21146 (N_21146,N_15830,N_16516);
nor U21147 (N_21147,N_19784,N_17569);
nand U21148 (N_21148,N_18861,N_19655);
nor U21149 (N_21149,N_19709,N_16291);
nand U21150 (N_21150,N_16883,N_15903);
xor U21151 (N_21151,N_16440,N_18410);
and U21152 (N_21152,N_19385,N_15954);
xor U21153 (N_21153,N_15608,N_18357);
and U21154 (N_21154,N_18877,N_16734);
and U21155 (N_21155,N_17776,N_15005);
nand U21156 (N_21156,N_15620,N_19857);
nor U21157 (N_21157,N_17522,N_15494);
xnor U21158 (N_21158,N_15369,N_15048);
nand U21159 (N_21159,N_19838,N_15535);
or U21160 (N_21160,N_15658,N_16905);
nand U21161 (N_21161,N_17277,N_18660);
and U21162 (N_21162,N_17202,N_17051);
or U21163 (N_21163,N_17043,N_15559);
nor U21164 (N_21164,N_17375,N_17633);
and U21165 (N_21165,N_19910,N_19942);
nor U21166 (N_21166,N_15764,N_19771);
nand U21167 (N_21167,N_16622,N_16580);
or U21168 (N_21168,N_17079,N_15690);
nor U21169 (N_21169,N_17294,N_16978);
nand U21170 (N_21170,N_18038,N_18887);
and U21171 (N_21171,N_18112,N_15843);
nor U21172 (N_21172,N_19381,N_17624);
xor U21173 (N_21173,N_19424,N_15560);
xnor U21174 (N_21174,N_16281,N_18744);
nand U21175 (N_21175,N_18731,N_18024);
nor U21176 (N_21176,N_19563,N_17071);
or U21177 (N_21177,N_19582,N_17811);
and U21178 (N_21178,N_19978,N_19068);
xor U21179 (N_21179,N_17436,N_17219);
nor U21180 (N_21180,N_17583,N_19896);
xor U21181 (N_21181,N_17797,N_17807);
xnor U21182 (N_21182,N_15622,N_19926);
and U21183 (N_21183,N_19395,N_19331);
xnor U21184 (N_21184,N_19047,N_16979);
and U21185 (N_21185,N_17802,N_15057);
and U21186 (N_21186,N_16193,N_15607);
nor U21187 (N_21187,N_19955,N_17727);
nand U21188 (N_21188,N_16947,N_19872);
nor U21189 (N_21189,N_17843,N_15453);
and U21190 (N_21190,N_15929,N_16981);
or U21191 (N_21191,N_18955,N_18344);
and U21192 (N_21192,N_18347,N_15878);
nand U21193 (N_21193,N_15966,N_19966);
nand U21194 (N_21194,N_18844,N_18075);
or U21195 (N_21195,N_16675,N_18255);
and U21196 (N_21196,N_19064,N_19693);
xnor U21197 (N_21197,N_19742,N_19724);
and U21198 (N_21198,N_17206,N_17190);
and U21199 (N_21199,N_15786,N_15131);
xor U21200 (N_21200,N_17132,N_15662);
nor U21201 (N_21201,N_17650,N_18537);
nor U21202 (N_21202,N_16977,N_19549);
nor U21203 (N_21203,N_17242,N_17606);
or U21204 (N_21204,N_19961,N_17178);
nor U21205 (N_21205,N_17628,N_16554);
and U21206 (N_21206,N_17093,N_18839);
and U21207 (N_21207,N_19828,N_16762);
xnor U21208 (N_21208,N_19626,N_17916);
nand U21209 (N_21209,N_17083,N_17233);
nand U21210 (N_21210,N_19690,N_15990);
nand U21211 (N_21211,N_16609,N_16778);
and U21212 (N_21212,N_16810,N_16710);
nor U21213 (N_21213,N_16595,N_17886);
nor U21214 (N_21214,N_16521,N_17850);
xor U21215 (N_21215,N_17611,N_18522);
xnor U21216 (N_21216,N_18061,N_17127);
nor U21217 (N_21217,N_19770,N_16816);
nor U21218 (N_21218,N_15980,N_17847);
nor U21219 (N_21219,N_16337,N_15958);
nor U21220 (N_21220,N_19003,N_17284);
nor U21221 (N_21221,N_18530,N_18052);
xor U21222 (N_21222,N_18840,N_18585);
nand U21223 (N_21223,N_19973,N_15600);
nand U21224 (N_21224,N_16304,N_19342);
nor U21225 (N_21225,N_17159,N_18223);
nor U21226 (N_21226,N_19495,N_17163);
or U21227 (N_21227,N_19851,N_16840);
or U21228 (N_21228,N_19704,N_16603);
xor U21229 (N_21229,N_16023,N_18835);
nand U21230 (N_21230,N_15149,N_18892);
nand U21231 (N_21231,N_19292,N_19683);
or U21232 (N_21232,N_17974,N_16918);
nor U21233 (N_21233,N_15045,N_16491);
or U21234 (N_21234,N_15914,N_18040);
xnor U21235 (N_21235,N_17014,N_17080);
or U21236 (N_21236,N_17526,N_17342);
or U21237 (N_21237,N_16871,N_16140);
and U21238 (N_21238,N_16506,N_16512);
nand U21239 (N_21239,N_17815,N_18483);
nor U21240 (N_21240,N_15506,N_16459);
xor U21241 (N_21241,N_15731,N_15114);
nand U21242 (N_21242,N_16495,N_17755);
and U21243 (N_21243,N_18471,N_16986);
and U21244 (N_21244,N_18766,N_15755);
or U21245 (N_21245,N_17291,N_16952);
nor U21246 (N_21246,N_15489,N_16135);
nand U21247 (N_21247,N_15063,N_19714);
or U21248 (N_21248,N_19706,N_19445);
and U21249 (N_21249,N_15214,N_18023);
nor U21250 (N_21250,N_17616,N_19830);
nor U21251 (N_21251,N_19019,N_15483);
or U21252 (N_21252,N_19190,N_16285);
or U21253 (N_21253,N_18773,N_18054);
and U21254 (N_21254,N_19894,N_19752);
xor U21255 (N_21255,N_15339,N_16663);
or U21256 (N_21256,N_15993,N_18579);
nor U21257 (N_21257,N_19790,N_17935);
nand U21258 (N_21258,N_15002,N_17809);
or U21259 (N_21259,N_15258,N_17478);
or U21260 (N_21260,N_16893,N_15814);
nand U21261 (N_21261,N_17934,N_16474);
or U21262 (N_21262,N_15209,N_17234);
nor U21263 (N_21263,N_17231,N_15500);
or U21264 (N_21264,N_18492,N_18678);
and U21265 (N_21265,N_16389,N_18595);
nand U21266 (N_21266,N_15493,N_19789);
or U21267 (N_21267,N_19399,N_18742);
xnor U21268 (N_21268,N_15482,N_19581);
xnor U21269 (N_21269,N_15774,N_19271);
xnor U21270 (N_21270,N_15278,N_18787);
and U21271 (N_21271,N_15027,N_17687);
xnor U21272 (N_21272,N_18433,N_17712);
nand U21273 (N_21273,N_15324,N_18455);
nand U21274 (N_21274,N_19436,N_16122);
xnor U21275 (N_21275,N_18646,N_18847);
nand U21276 (N_21276,N_16370,N_19525);
xor U21277 (N_21277,N_17548,N_16311);
nand U21278 (N_21278,N_17887,N_19145);
nand U21279 (N_21279,N_17946,N_17713);
nor U21280 (N_21280,N_15035,N_16660);
nor U21281 (N_21281,N_19350,N_17425);
xor U21282 (N_21282,N_15779,N_18997);
and U21283 (N_21283,N_15708,N_16066);
nand U21284 (N_21284,N_18283,N_16467);
xnor U21285 (N_21285,N_19330,N_15141);
xor U21286 (N_21286,N_18788,N_18186);
and U21287 (N_21287,N_16150,N_18743);
xor U21288 (N_21288,N_18021,N_18316);
nor U21289 (N_21289,N_17501,N_15100);
or U21290 (N_21290,N_16953,N_18640);
nor U21291 (N_21291,N_19477,N_18657);
and U21292 (N_21292,N_17194,N_18250);
or U21293 (N_21293,N_15067,N_15424);
nand U21294 (N_21294,N_17785,N_19230);
and U21295 (N_21295,N_18817,N_19996);
nand U21296 (N_21296,N_19547,N_18949);
or U21297 (N_21297,N_16428,N_19934);
or U21298 (N_21298,N_17210,N_19437);
nand U21299 (N_21299,N_15705,N_15238);
nor U21300 (N_21300,N_17441,N_18652);
nand U21301 (N_21301,N_16884,N_18464);
xnor U21302 (N_21302,N_19069,N_18049);
or U21303 (N_21303,N_15552,N_18355);
nor U21304 (N_21304,N_18148,N_15524);
xor U21305 (N_21305,N_16677,N_19430);
nor U21306 (N_21306,N_15269,N_16074);
nand U21307 (N_21307,N_17658,N_17027);
xnor U21308 (N_21308,N_15766,N_18247);
xnor U21309 (N_21309,N_18529,N_18394);
and U21310 (N_21310,N_16508,N_19389);
or U21311 (N_21311,N_18491,N_19519);
nand U21312 (N_21312,N_16766,N_19695);
nor U21313 (N_21313,N_16052,N_19939);
nor U21314 (N_21314,N_19514,N_17024);
or U21315 (N_21315,N_16630,N_19836);
xor U21316 (N_21316,N_18784,N_18528);
and U21317 (N_21317,N_19618,N_19533);
nor U21318 (N_21318,N_17303,N_15586);
xnor U21319 (N_21319,N_17572,N_19231);
or U21320 (N_21320,N_18857,N_15736);
xor U21321 (N_21321,N_19211,N_16849);
nor U21322 (N_21322,N_16045,N_18673);
nand U21323 (N_21323,N_18694,N_16549);
or U21324 (N_21324,N_16678,N_19067);
nand U21325 (N_21325,N_16743,N_16976);
nor U21326 (N_21326,N_19323,N_18370);
or U21327 (N_21327,N_16865,N_18450);
xnor U21328 (N_21328,N_17778,N_15905);
nor U21329 (N_21329,N_18923,N_17857);
and U21330 (N_21330,N_15587,N_16098);
or U21331 (N_21331,N_16410,N_19541);
xor U21332 (N_21332,N_16472,N_19135);
or U21333 (N_21333,N_18737,N_17188);
or U21334 (N_21334,N_16526,N_15722);
or U21335 (N_21335,N_15952,N_19531);
xor U21336 (N_21336,N_18778,N_16674);
or U21337 (N_21337,N_16631,N_17818);
or U21338 (N_21338,N_17623,N_17331);
nand U21339 (N_21339,N_19142,N_17045);
xor U21340 (N_21340,N_18158,N_18566);
and U21341 (N_21341,N_16848,N_16297);
xor U21342 (N_21342,N_15788,N_19459);
nor U21343 (N_21343,N_17347,N_17447);
nor U21344 (N_21344,N_15450,N_15789);
nand U21345 (N_21345,N_17098,N_18874);
nand U21346 (N_21346,N_17109,N_17596);
and U21347 (N_21347,N_15457,N_18763);
xor U21348 (N_21348,N_15762,N_16530);
nand U21349 (N_21349,N_17252,N_15248);
xor U21350 (N_21350,N_15468,N_16658);
and U21351 (N_21351,N_17681,N_18815);
and U21352 (N_21352,N_19520,N_19018);
xnor U21353 (N_21353,N_18120,N_17411);
xnor U21354 (N_21354,N_16626,N_16226);
nor U21355 (N_21355,N_17454,N_17533);
or U21356 (N_21356,N_16858,N_16189);
xor U21357 (N_21357,N_17088,N_16607);
or U21358 (N_21358,N_19691,N_19807);
and U21359 (N_21359,N_16300,N_16558);
nor U21360 (N_21360,N_15077,N_16072);
and U21361 (N_21361,N_15876,N_16949);
nand U21362 (N_21362,N_18697,N_15222);
xor U21363 (N_21363,N_18812,N_15881);
nor U21364 (N_21364,N_16356,N_16723);
or U21365 (N_21365,N_19250,N_19213);
nor U21366 (N_21366,N_17822,N_18312);
or U21367 (N_21367,N_17169,N_18592);
and U21368 (N_21368,N_16155,N_16449);
and U21369 (N_21369,N_15321,N_16018);
xor U21370 (N_21370,N_16341,N_15015);
xnor U21371 (N_21371,N_19468,N_17855);
and U21372 (N_21372,N_18262,N_15582);
nor U21373 (N_21373,N_16405,N_18944);
or U21374 (N_21374,N_15834,N_19512);
nand U21375 (N_21375,N_16941,N_18610);
xnor U21376 (N_21376,N_15279,N_16576);
nor U21377 (N_21377,N_16593,N_17665);
or U21378 (N_21378,N_16932,N_18670);
nor U21379 (N_21379,N_19278,N_18380);
nor U21380 (N_21380,N_17072,N_18908);
xnor U21381 (N_21381,N_15783,N_15246);
nand U21382 (N_21382,N_15570,N_19668);
or U21383 (N_21383,N_19152,N_16916);
nand U21384 (N_21384,N_15734,N_16851);
nor U21385 (N_21385,N_18606,N_18323);
or U21386 (N_21386,N_16824,N_16740);
and U21387 (N_21387,N_19265,N_19988);
or U21388 (N_21388,N_17293,N_19148);
xor U21389 (N_21389,N_19968,N_15054);
nor U21390 (N_21390,N_17549,N_18967);
xnor U21391 (N_21391,N_16177,N_19042);
and U21392 (N_21392,N_18030,N_17466);
and U21393 (N_21393,N_19800,N_17782);
and U21394 (N_21394,N_19444,N_19566);
nor U21395 (N_21395,N_16818,N_19167);
xor U21396 (N_21396,N_18954,N_16712);
or U21397 (N_21397,N_18644,N_18948);
nor U21398 (N_21398,N_15091,N_19258);
and U21399 (N_21399,N_16362,N_19962);
nor U21400 (N_21400,N_19365,N_18143);
nand U21401 (N_21401,N_17589,N_18653);
xor U21402 (N_21402,N_19035,N_15768);
and U21403 (N_21403,N_19082,N_17638);
or U21404 (N_21404,N_17914,N_17982);
or U21405 (N_21405,N_18932,N_18601);
xnor U21406 (N_21406,N_19909,N_18213);
or U21407 (N_21407,N_18985,N_17106);
nor U21408 (N_21408,N_16564,N_15286);
or U21409 (N_21409,N_18240,N_17429);
nor U21410 (N_21410,N_15868,N_15359);
xnor U21411 (N_21411,N_18524,N_16105);
nor U21412 (N_21412,N_17545,N_18184);
and U21413 (N_21413,N_16451,N_15044);
xor U21414 (N_21414,N_18031,N_17761);
and U21415 (N_21415,N_16083,N_15867);
nand U21416 (N_21416,N_19765,N_15252);
and U21417 (N_21417,N_19889,N_19245);
and U21418 (N_21418,N_16275,N_17931);
or U21419 (N_21419,N_19386,N_19078);
nor U21420 (N_21420,N_16786,N_17065);
xnor U21421 (N_21421,N_15580,N_19676);
xnor U21422 (N_21422,N_15353,N_18553);
nor U21423 (N_21423,N_18480,N_18099);
and U21424 (N_21424,N_19982,N_19263);
xnor U21425 (N_21425,N_18940,N_19461);
nand U21426 (N_21426,N_15838,N_17672);
and U21427 (N_21427,N_18875,N_15871);
and U21428 (N_21428,N_18541,N_19711);
nor U21429 (N_21429,N_15284,N_18013);
xnor U21430 (N_21430,N_19601,N_16190);
and U21431 (N_21431,N_16657,N_16867);
or U21432 (N_21432,N_18201,N_17435);
or U21433 (N_21433,N_17056,N_15337);
nand U21434 (N_21434,N_18466,N_17609);
or U21435 (N_21435,N_18692,N_17340);
nand U21436 (N_21436,N_18232,N_15556);
xnor U21437 (N_21437,N_19662,N_19457);
nand U21438 (N_21438,N_15038,N_19692);
xor U21439 (N_21439,N_17651,N_18811);
or U21440 (N_21440,N_15589,N_19780);
xor U21441 (N_21441,N_19670,N_18327);
nand U21442 (N_21442,N_15382,N_17691);
and U21443 (N_21443,N_15664,N_16077);
and U21444 (N_21444,N_18128,N_17495);
and U21445 (N_21445,N_18891,N_17015);
or U21446 (N_21446,N_15998,N_16179);
xnor U21447 (N_21447,N_19991,N_15441);
xnor U21448 (N_21448,N_15341,N_17594);
and U21449 (N_21449,N_16213,N_19623);
xor U21450 (N_21450,N_18242,N_19435);
nand U21451 (N_21451,N_18596,N_15210);
nand U21452 (N_21452,N_16860,N_18690);
or U21453 (N_21453,N_15978,N_15155);
and U21454 (N_21454,N_17308,N_17636);
or U21455 (N_21455,N_15584,N_15492);
nand U21456 (N_21456,N_18521,N_17117);
or U21457 (N_21457,N_18782,N_18520);
xor U21458 (N_21458,N_17577,N_17181);
nand U21459 (N_21459,N_19101,N_15811);
and U21460 (N_21460,N_15529,N_16930);
nand U21461 (N_21461,N_16567,N_18475);
or U21462 (N_21462,N_18281,N_17669);
and U21463 (N_21463,N_18584,N_16399);
xnor U21464 (N_21464,N_16906,N_18098);
nor U21465 (N_21465,N_19462,N_16588);
nand U21466 (N_21466,N_16886,N_16868);
nand U21467 (N_21467,N_18245,N_19782);
and U21468 (N_21468,N_18947,N_19981);
nand U21469 (N_21469,N_18717,N_18958);
and U21470 (N_21470,N_19669,N_18846);
nand U21471 (N_21471,N_16330,N_15920);
or U21472 (N_21472,N_16001,N_15623);
nor U21473 (N_21473,N_18364,N_18474);
or U21474 (N_21474,N_17966,N_18855);
and U21475 (N_21475,N_16655,N_15406);
xnor U21476 (N_21476,N_17068,N_19873);
and U21477 (N_21477,N_18234,N_16200);
nor U21478 (N_21478,N_15611,N_18804);
and U21479 (N_21479,N_17330,N_15979);
or U21480 (N_21480,N_18399,N_17805);
nor U21481 (N_21481,N_17910,N_18453);
nor U21482 (N_21482,N_15306,N_17008);
and U21483 (N_21483,N_18519,N_15643);
xnor U21484 (N_21484,N_15827,N_18443);
xnor U21485 (N_21485,N_19808,N_16133);
and U21486 (N_21486,N_15200,N_16167);
xor U21487 (N_21487,N_19260,N_15416);
nor U21488 (N_21488,N_19732,N_17734);
nor U21489 (N_21489,N_19307,N_16229);
and U21490 (N_21490,N_17295,N_16728);
and U21491 (N_21491,N_19681,N_18959);
or U21492 (N_21492,N_16239,N_19308);
nor U21493 (N_21493,N_15152,N_16768);
or U21494 (N_21494,N_15147,N_18981);
or U21495 (N_21495,N_16301,N_19744);
nand U21496 (N_21496,N_18363,N_15144);
and U21497 (N_21497,N_16735,N_19215);
nand U21498 (N_21498,N_16096,N_15986);
nand U21499 (N_21499,N_17050,N_17680);
xnor U21500 (N_21500,N_16624,N_16739);
xnor U21501 (N_21501,N_19797,N_19352);
xnor U21502 (N_21502,N_16120,N_15753);
xor U21503 (N_21503,N_18622,N_17199);
and U21504 (N_21504,N_15464,N_15387);
and U21505 (N_21505,N_18608,N_15928);
nand U21506 (N_21506,N_18192,N_15123);
or U21507 (N_21507,N_16196,N_17947);
xnor U21508 (N_21508,N_19843,N_17872);
nand U21509 (N_21509,N_15298,N_16111);
nand U21510 (N_21510,N_17753,N_15517);
nand U21511 (N_21511,N_16386,N_18318);
nor U21512 (N_21512,N_16618,N_18669);
xnor U21513 (N_21513,N_19902,N_16161);
xnor U21514 (N_21514,N_17829,N_16269);
xnor U21515 (N_21515,N_15024,N_15633);
nor U21516 (N_21516,N_16598,N_17018);
nand U21517 (N_21517,N_16610,N_16376);
nand U21518 (N_21518,N_18300,N_18230);
xnor U21519 (N_21519,N_15285,N_15668);
and U21520 (N_21520,N_19465,N_17656);
or U21521 (N_21521,N_16507,N_17391);
and U21522 (N_21522,N_17301,N_19911);
or U21523 (N_21523,N_19058,N_17197);
nand U21524 (N_21524,N_16746,N_15769);
or U21525 (N_21525,N_18109,N_15142);
and U21526 (N_21526,N_15143,N_15232);
and U21527 (N_21527,N_18770,N_16020);
nor U21528 (N_21528,N_15390,N_17105);
nand U21529 (N_21529,N_16819,N_18228);
xnor U21530 (N_21530,N_18880,N_15196);
or U21531 (N_21531,N_15398,N_15153);
or U21532 (N_21532,N_18361,N_15350);
or U21533 (N_21533,N_19377,N_17240);
or U21534 (N_21534,N_15659,N_15099);
xor U21535 (N_21535,N_17793,N_18573);
nand U21536 (N_21536,N_17525,N_16581);
and U21537 (N_21537,N_19312,N_18456);
nor U21538 (N_21538,N_19037,N_16614);
xnor U21539 (N_21539,N_17688,N_16830);
and U21540 (N_21540,N_18367,N_15689);
and U21541 (N_21541,N_16574,N_16988);
or U21542 (N_21542,N_18012,N_15467);
xor U21543 (N_21543,N_18420,N_18679);
and U21544 (N_21544,N_19529,N_17393);
or U21545 (N_21545,N_16555,N_15355);
or U21546 (N_21546,N_15163,N_16027);
nand U21547 (N_21547,N_16310,N_19527);
xnor U21548 (N_21548,N_16249,N_16452);
nand U21549 (N_21549,N_15860,N_16461);
or U21550 (N_21550,N_19456,N_18772);
and U21551 (N_21551,N_18602,N_15336);
nand U21552 (N_21552,N_15295,N_17321);
and U21553 (N_21553,N_17563,N_16228);
nand U21554 (N_21554,N_15429,N_17538);
nand U21555 (N_21555,N_18430,N_19998);
nor U21556 (N_21556,N_15505,N_19464);
and U21557 (N_21557,N_15283,N_18294);
nor U21558 (N_21558,N_16843,N_18324);
and U21559 (N_21559,N_18241,N_19613);
nor U21560 (N_21560,N_15629,N_19643);
or U21561 (N_21561,N_18102,N_18498);
or U21562 (N_21562,N_18362,N_17552);
xor U21563 (N_21563,N_17962,N_18487);
or U21564 (N_21564,N_19438,N_17715);
or U21565 (N_21565,N_18403,N_18107);
xor U21566 (N_21566,N_15627,N_17581);
or U21567 (N_21567,N_16577,N_15240);
nor U21568 (N_21568,N_17237,N_15725);
nor U21569 (N_21569,N_15081,N_18795);
xor U21570 (N_21570,N_19199,N_16460);
nor U21571 (N_21571,N_18458,N_18484);
nor U21572 (N_21572,N_17795,N_16515);
xor U21573 (N_21573,N_17880,N_18761);
and U21574 (N_21574,N_15877,N_15703);
nand U21575 (N_21575,N_17135,N_15329);
and U21576 (N_21576,N_15271,N_15583);
and U21577 (N_21577,N_17913,N_15723);
xor U21578 (N_21578,N_15215,N_19398);
nand U21579 (N_21579,N_15618,N_18925);
and U21580 (N_21580,N_17260,N_17166);
and U21581 (N_21581,N_18218,N_19913);
and U21582 (N_21582,N_18439,N_16732);
or U21583 (N_21583,N_19792,N_15071);
nand U21584 (N_21584,N_15203,N_15558);
and U21585 (N_21585,N_16176,N_18785);
and U21586 (N_21586,N_15171,N_18890);
nor U21587 (N_21587,N_17537,N_16290);
nand U21588 (N_21588,N_15377,N_19941);
or U21589 (N_21589,N_16209,N_16295);
xor U21590 (N_21590,N_18879,N_19401);
nor U21591 (N_21591,N_17587,N_16627);
xnor U21592 (N_21592,N_16767,N_19027);
or U21593 (N_21593,N_19610,N_17915);
xor U21594 (N_21594,N_17332,N_18215);
or U21595 (N_21595,N_18446,N_19818);
xor U21596 (N_21596,N_15037,N_15305);
nand U21597 (N_21597,N_16335,N_19542);
or U21598 (N_21598,N_15961,N_17089);
and U21599 (N_21599,N_17067,N_15431);
and U21600 (N_21600,N_18800,N_17851);
and U21601 (N_21601,N_18517,N_19883);
xor U21602 (N_21602,N_18164,N_19860);
xor U21603 (N_21603,N_15328,N_16366);
nor U21604 (N_21604,N_15125,N_16199);
and U21605 (N_21605,N_15363,N_19874);
nor U21606 (N_21606,N_15526,N_18070);
xnor U21607 (N_21607,N_18331,N_18934);
xnor U21608 (N_21608,N_18190,N_15476);
nand U21609 (N_21609,N_18685,N_16703);
and U21610 (N_21610,N_15204,N_16425);
or U21611 (N_21611,N_17908,N_18159);
and U21612 (N_21612,N_15122,N_16822);
xnor U21613 (N_21613,N_19561,N_17523);
nand U21614 (N_21614,N_19279,N_15968);
xnor U21615 (N_21615,N_19852,N_15887);
nand U21616 (N_21616,N_17134,N_17486);
and U21617 (N_21617,N_18714,N_16233);
xor U21618 (N_21618,N_19634,N_15824);
or U21619 (N_21619,N_18684,N_19672);
nand U21620 (N_21620,N_16813,N_18090);
and U21621 (N_21621,N_17285,N_16232);
nand U21622 (N_21622,N_15670,N_16765);
and U21623 (N_21623,N_15218,N_15367);
nor U21624 (N_21624,N_17305,N_17128);
nor U21625 (N_21625,N_18328,N_17597);
or U21626 (N_21626,N_18695,N_19467);
nor U21627 (N_21627,N_18971,N_17028);
or U21628 (N_21628,N_19110,N_15655);
and U21629 (N_21629,N_17575,N_16128);
and U21630 (N_21630,N_19624,N_18279);
and U21631 (N_21631,N_18631,N_17153);
and U21632 (N_21632,N_15685,N_17641);
and U21633 (N_21633,N_16288,N_18516);
nand U21634 (N_21634,N_15963,N_19722);
nor U21635 (N_21635,N_15228,N_17297);
or U21636 (N_21636,N_18418,N_16136);
nand U21637 (N_21637,N_19510,N_19318);
nand U21638 (N_21638,N_16908,N_19268);
nor U21639 (N_21639,N_15466,N_18256);
nand U21640 (N_21640,N_18197,N_15095);
and U21641 (N_21641,N_18689,N_16298);
or U21642 (N_21642,N_15748,N_17344);
and U21643 (N_21643,N_15569,N_19384);
nand U21644 (N_21644,N_15853,N_19850);
xnor U21645 (N_21645,N_17108,N_15520);
and U21646 (N_21646,N_17432,N_15967);
or U21647 (N_21647,N_18676,N_16080);
nand U21648 (N_21648,N_15105,N_17165);
nor U21649 (N_21649,N_15850,N_16048);
xnor U21650 (N_21650,N_16354,N_16323);
xnor U21651 (N_21651,N_19091,N_19083);
and U21652 (N_21652,N_17693,N_18641);
nand U21653 (N_21653,N_17938,N_17147);
and U21654 (N_21654,N_17003,N_17654);
and U21655 (N_21655,N_19138,N_18123);
and U21656 (N_21656,N_17719,N_15981);
xnor U21657 (N_21657,N_15408,N_17904);
nand U21658 (N_21658,N_18668,N_15475);
and U21659 (N_21659,N_19326,N_19760);
xor U21660 (N_21660,N_16456,N_19126);
and U21661 (N_21661,N_19675,N_16403);
xor U21662 (N_21662,N_15184,N_16669);
and U21663 (N_21663,N_15090,N_17356);
and U21664 (N_21664,N_15195,N_19029);
xor U21665 (N_21665,N_15650,N_19756);
and U21666 (N_21666,N_18915,N_16248);
xnor U21667 (N_21667,N_18170,N_16432);
nor U21668 (N_21668,N_19546,N_15904);
nand U21669 (N_21669,N_17010,N_19659);
or U21670 (N_21670,N_17465,N_17278);
and U21671 (N_21671,N_16152,N_18205);
nand U21672 (N_21672,N_15906,N_16025);
xor U21673 (N_21673,N_17401,N_15135);
or U21674 (N_21674,N_16853,N_16901);
and U21675 (N_21675,N_17440,N_16418);
nand U21676 (N_21676,N_16419,N_17814);
nor U21677 (N_21677,N_16414,N_17701);
nor U21678 (N_21678,N_18546,N_18282);
and U21679 (N_21679,N_19578,N_18704);
xor U21680 (N_21680,N_15432,N_19221);
and U21681 (N_21681,N_18338,N_15319);
nand U21682 (N_21682,N_17390,N_19006);
or U21683 (N_21683,N_17082,N_16727);
nand U21684 (N_21684,N_19301,N_17226);
nand U21685 (N_21685,N_19111,N_19372);
nor U21686 (N_21686,N_19579,N_18790);
and U21687 (N_21687,N_18603,N_17842);
and U21688 (N_21688,N_17668,N_16896);
nor U21689 (N_21689,N_15530,N_18993);
xor U21690 (N_21690,N_17879,N_15397);
nand U21691 (N_21691,N_17081,N_18321);
or U21692 (N_21692,N_15601,N_19593);
or U21693 (N_21693,N_15984,N_15471);
nand U21694 (N_21694,N_17774,N_16245);
and U21695 (N_21695,N_17364,N_17675);
nand U21696 (N_21696,N_18366,N_19022);
xor U21697 (N_21697,N_15849,N_15480);
xnor U21698 (N_21698,N_15132,N_17483);
nor U21699 (N_21699,N_19758,N_19606);
and U21700 (N_21700,N_17900,N_18500);
or U21701 (N_21701,N_19196,N_17457);
nor U21702 (N_21702,N_17290,N_17248);
xnor U21703 (N_21703,N_19835,N_15488);
xor U21704 (N_21704,N_16314,N_16528);
or U21705 (N_21705,N_16437,N_18290);
or U21706 (N_21706,N_16891,N_15034);
and U21707 (N_21707,N_16240,N_15962);
nand U21708 (N_21708,N_17695,N_19501);
or U21709 (N_21709,N_19004,N_18655);
or U21710 (N_21710,N_18422,N_18272);
nor U21711 (N_21711,N_15637,N_15006);
nor U21712 (N_21712,N_16201,N_15351);
xnor U21713 (N_21713,N_16373,N_16395);
and U21714 (N_21714,N_15951,N_17832);
xnor U21715 (N_21715,N_16069,N_15334);
or U21716 (N_21716,N_16309,N_16939);
nand U21717 (N_21717,N_18325,N_16125);
nor U21718 (N_21718,N_16925,N_18771);
nor U21719 (N_21719,N_15491,N_19179);
nor U21720 (N_21720,N_19900,N_17804);
nor U21721 (N_21721,N_19580,N_18831);
nand U21722 (N_21722,N_17869,N_18727);
or U21723 (N_21723,N_19666,N_19801);
xnor U21724 (N_21724,N_16962,N_19054);
and U21725 (N_21725,N_17264,N_19052);
or U21726 (N_21726,N_17152,N_16877);
nor U21727 (N_21727,N_18295,N_18961);
or U21728 (N_21728,N_19310,N_15743);
or U21729 (N_21729,N_19391,N_16488);
nand U21730 (N_21730,N_17449,N_18277);
or U21731 (N_21731,N_15543,N_16760);
nor U21732 (N_21732,N_19287,N_16162);
nand U21733 (N_21733,N_15326,N_18639);
xnor U21734 (N_21734,N_17610,N_15686);
nor U21735 (N_21735,N_16401,N_17406);
xnor U21736 (N_21736,N_16137,N_15370);
and U21737 (N_21737,N_15373,N_15810);
nor U21738 (N_21738,N_17239,N_17987);
xnor U21739 (N_21739,N_16779,N_19490);
and U21740 (N_21740,N_19421,N_15229);
xnor U21741 (N_21741,N_16477,N_17867);
and U21742 (N_21742,N_16422,N_15619);
xnor U21743 (N_21743,N_17967,N_17873);
or U21744 (N_21744,N_19571,N_19840);
and U21745 (N_21745,N_18946,N_17055);
xor U21746 (N_21746,N_16502,N_16458);
or U21747 (N_21747,N_19290,N_15817);
nand U21748 (N_21748,N_19513,N_18032);
xnor U21749 (N_21749,N_15456,N_18083);
nor U21750 (N_21750,N_15444,N_18675);
xnor U21751 (N_21751,N_19241,N_17894);
nor U21752 (N_21752,N_17456,N_18716);
xor U21753 (N_21753,N_17203,N_18512);
nor U21754 (N_21754,N_15918,N_19735);
xnor U21755 (N_21755,N_19172,N_16911);
nor U21756 (N_21756,N_18856,N_17979);
nor U21757 (N_21757,N_17167,N_19093);
nor U21758 (N_21758,N_19136,N_18922);
nand U21759 (N_21759,N_17921,N_19999);
and U21760 (N_21760,N_17046,N_18127);
xor U21761 (N_21761,N_17492,N_16544);
nor U21762 (N_21762,N_15348,N_18928);
nand U21763 (N_21763,N_16132,N_19491);
nand U21764 (N_21764,N_18838,N_15192);
xnor U21765 (N_21765,N_18501,N_15718);
and U21766 (N_21766,N_18598,N_15711);
xor U21767 (N_21767,N_19707,N_19849);
xnor U21768 (N_21768,N_16844,N_19216);
xor U21769 (N_21769,N_18514,N_18515);
xnor U21770 (N_21770,N_19147,N_17384);
nor U21771 (N_21771,N_19254,N_19656);
xor U21772 (N_21772,N_15553,N_18982);
xnor U21773 (N_21773,N_18369,N_17115);
nor U21774 (N_21774,N_18006,N_15577);
nand U21775 (N_21775,N_17803,N_18333);
nand U21776 (N_21776,N_15515,N_15976);
nand U21777 (N_21777,N_16326,N_15749);
and U21778 (N_21778,N_15407,N_16829);
nor U21779 (N_21779,N_15340,N_19562);
nand U21780 (N_21780,N_15605,N_19183);
nand U21781 (N_21781,N_16014,N_19280);
xnor U21782 (N_21782,N_15257,N_19876);
nor U21783 (N_21783,N_18721,N_15345);
xnor U21784 (N_21784,N_16909,N_17473);
nor U21785 (N_21785,N_17725,N_18849);
nand U21786 (N_21786,N_18103,N_15709);
nor U21787 (N_21787,N_19603,N_18050);
nor U21788 (N_21788,N_18746,N_15265);
xnor U21789 (N_21789,N_15244,N_19368);
nor U21790 (N_21790,N_16260,N_17599);
xor U21791 (N_21791,N_15462,N_19972);
xnor U21792 (N_21792,N_15667,N_19159);
nor U21793 (N_21793,N_16504,N_15895);
nor U21794 (N_21794,N_19353,N_16108);
and U21795 (N_21795,N_16967,N_17272);
xnor U21796 (N_21796,N_18445,N_19355);
and U21797 (N_21797,N_17077,N_18701);
nor U21798 (N_21798,N_16261,N_15239);
nor U21799 (N_21799,N_15107,N_19820);
nor U21800 (N_21800,N_16881,N_19238);
nor U21801 (N_21801,N_15230,N_16463);
nand U21802 (N_21802,N_15900,N_18965);
nand U21803 (N_21803,N_16470,N_15374);
or U21804 (N_21804,N_15020,N_17820);
nand U21805 (N_21805,N_18916,N_16268);
xnor U21806 (N_21806,N_18505,N_18557);
and U21807 (N_21807,N_16205,N_16494);
nand U21808 (N_21808,N_18265,N_16019);
nor U21809 (N_21809,N_16185,N_19757);
or U21810 (N_21810,N_15375,N_15314);
xor U21811 (N_21811,N_15160,N_15538);
and U21812 (N_21812,N_19340,N_15162);
nor U21813 (N_21813,N_19131,N_15747);
or U21814 (N_21814,N_16090,N_17666);
and U21815 (N_21815,N_17230,N_19034);
nor U21816 (N_21816,N_16557,N_19569);
or U21817 (N_21817,N_18796,N_16590);
nand U21818 (N_21818,N_15696,N_15940);
or U21819 (N_21819,N_18980,N_15347);
xnor U21820 (N_21820,N_19621,N_17881);
nor U21821 (N_21821,N_18334,N_19474);
or U21822 (N_21822,N_16836,N_17590);
xnor U21823 (N_21823,N_19987,N_16797);
and U21824 (N_21824,N_17385,N_19072);
nor U21825 (N_21825,N_18858,N_15459);
nor U21826 (N_21826,N_19169,N_19667);
nor U21827 (N_21827,N_15896,N_18431);
and U21828 (N_21828,N_19102,N_17816);
nor U21829 (N_21829,N_17004,N_17619);
or U21830 (N_21830,N_15729,N_16147);
and U21831 (N_21831,N_16089,N_16568);
and U21832 (N_21832,N_16033,N_19944);
nor U21833 (N_21833,N_17584,N_18638);
xnor U21834 (N_21834,N_15985,N_15262);
nor U21835 (N_21835,N_16656,N_18237);
and U21836 (N_21836,N_18384,N_19480);
nand U21837 (N_21837,N_19602,N_18048);
nor U21838 (N_21838,N_16989,N_18000);
or U21839 (N_21839,N_15699,N_15532);
nor U21840 (N_21840,N_18977,N_15094);
xor U21841 (N_21841,N_17176,N_15661);
and U21842 (N_21842,N_19400,N_16889);
xor U21843 (N_21843,N_16501,N_18830);
nor U21844 (N_21844,N_16119,N_17026);
nor U21845 (N_21845,N_17334,N_15290);
nor U21846 (N_21846,N_18590,N_18345);
nor U21847 (N_21847,N_18133,N_15578);
or U21848 (N_21848,N_15765,N_17476);
nor U21849 (N_21849,N_17586,N_18425);
xnor U21850 (N_21850,N_19839,N_17993);
and U21851 (N_21851,N_17229,N_19951);
xor U21852 (N_21852,N_15610,N_15588);
and U21853 (N_21853,N_19976,N_19162);
nor U21854 (N_21854,N_19476,N_19921);
nor U21855 (N_21855,N_17647,N_15496);
and U21856 (N_21856,N_17911,N_16751);
and U21857 (N_21857,N_17759,N_15371);
and U21858 (N_21858,N_16936,N_16198);
and U21859 (N_21859,N_18008,N_18711);
xnor U21860 (N_21860,N_19575,N_19165);
nand U21861 (N_21861,N_17786,N_17049);
or U21862 (N_21862,N_18077,N_17853);
nand U21863 (N_21863,N_17562,N_19411);
nand U21864 (N_21864,N_17209,N_16500);
xor U21865 (N_21865,N_17642,N_19971);
and U21866 (N_21866,N_19507,N_18819);
and U21867 (N_21867,N_19404,N_15972);
nand U21868 (N_21868,N_19151,N_18752);
or U21869 (N_21869,N_15167,N_18122);
and U21870 (N_21870,N_16776,N_18956);
nor U21871 (N_21871,N_17064,N_15404);
nor U21872 (N_21872,N_19509,N_17792);
and U21873 (N_21873,N_19498,N_17743);
nand U21874 (N_21874,N_15236,N_15472);
or U21875 (N_21875,N_19313,N_19785);
or U21876 (N_21876,N_19294,N_15096);
nand U21877 (N_21877,N_17747,N_19440);
nor U21878 (N_21878,N_18621,N_19635);
xnor U21879 (N_21879,N_18221,N_16257);
and U21880 (N_21880,N_18794,N_18672);
or U21881 (N_21881,N_19364,N_17382);
xnor U21882 (N_21882,N_15573,N_19984);
nand U21883 (N_21883,N_17591,N_15042);
nand U21884 (N_21884,N_15949,N_19048);
nand U21885 (N_21885,N_19433,N_16095);
or U21886 (N_21886,N_15937,N_17748);
and U21887 (N_21887,N_17306,N_18645);
nand U21888 (N_21888,N_16324,N_16172);
nor U21889 (N_21889,N_17764,N_19485);
nor U21890 (N_21890,N_16646,N_15361);
nor U21891 (N_21891,N_17172,N_16070);
and U21892 (N_21892,N_18543,N_18693);
nor U21893 (N_21893,N_19960,N_16828);
and U21894 (N_21894,N_18310,N_15923);
xor U21895 (N_21895,N_19139,N_16210);
nor U21896 (N_21896,N_19077,N_18767);
xor U21897 (N_21897,N_19009,N_18441);
nand U21898 (N_21898,N_17505,N_19931);
nand U21899 (N_21899,N_16685,N_16044);
nand U21900 (N_21900,N_16758,N_15249);
and U21901 (N_21901,N_15791,N_15936);
or U21902 (N_21902,N_16605,N_17479);
nand U21903 (N_21903,N_19120,N_18053);
xnor U21904 (N_21904,N_16085,N_16394);
and U21905 (N_21905,N_17096,N_19192);
and U21906 (N_21906,N_18373,N_17198);
or U21907 (N_21907,N_18187,N_18313);
or U21908 (N_21908,N_18065,N_18095);
nor U21909 (N_21909,N_18405,N_18802);
or U21910 (N_21910,N_16775,N_15997);
nand U21911 (N_21911,N_18570,N_17973);
or U21912 (N_21912,N_15247,N_16344);
xor U21913 (N_21913,N_17992,N_16997);
nand U21914 (N_21914,N_17107,N_19096);
xor U21915 (N_21915,N_19175,N_15908);
xnor U21916 (N_21916,N_19217,N_15518);
nor U21917 (N_21917,N_15346,N_18611);
or U21918 (N_21918,N_17561,N_17170);
xor U21919 (N_21919,N_19205,N_18383);
xnor U21920 (N_21920,N_19055,N_19487);
nand U21921 (N_21921,N_19388,N_16265);
nand U21922 (N_21922,N_18552,N_19879);
or U21923 (N_21923,N_15221,N_18503);
or U21924 (N_21924,N_16244,N_16180);
and U21925 (N_21925,N_16050,N_16385);
or U21926 (N_21926,N_17263,N_15470);
or U21927 (N_21927,N_16262,N_17883);
xor U21928 (N_21928,N_16910,N_15975);
and U21929 (N_21929,N_19980,N_16002);
nand U21930 (N_21930,N_19283,N_18842);
xor U21931 (N_21931,N_16236,N_17605);
xnor U21932 (N_21932,N_16659,N_16303);
nor U21933 (N_21933,N_17655,N_17485);
and U21934 (N_21934,N_15315,N_19374);
xnor U21935 (N_21935,N_15888,N_19907);
or U21936 (N_21936,N_16917,N_15130);
xor U21937 (N_21937,N_15507,N_17273);
and U21938 (N_21938,N_15364,N_19523);
nand U21939 (N_21939,N_15772,N_15443);
or U21940 (N_21940,N_17119,N_19057);
nand U21941 (N_21941,N_17870,N_16704);
xnor U21942 (N_21942,N_15819,N_18341);
nand U21943 (N_21943,N_15047,N_19267);
nand U21944 (N_21944,N_18093,N_17896);
nand U21945 (N_21945,N_16785,N_18348);
nand U21946 (N_21946,N_17906,N_17644);
and U21947 (N_21947,N_16211,N_18131);
nand U21948 (N_21948,N_19449,N_15592);
nor U21949 (N_21949,N_19106,N_19684);
and U21950 (N_21950,N_15942,N_17737);
nand U21951 (N_21951,N_16192,N_18927);
nor U21952 (N_21952,N_15720,N_16928);
nor U21953 (N_21953,N_16982,N_19150);
and U21954 (N_21954,N_16615,N_19225);
or U21955 (N_21955,N_18132,N_19945);
or U21956 (N_21956,N_18060,N_15678);
or U21957 (N_21957,N_17029,N_17196);
and U21958 (N_21958,N_15724,N_16879);
nor U21959 (N_21959,N_18572,N_16796);
nor U21960 (N_21960,N_17697,N_16681);
or U21961 (N_21961,N_18559,N_16036);
or U21962 (N_21962,N_18026,N_19615);
nor U21963 (N_21963,N_17386,N_19543);
nand U21964 (N_21964,N_16170,N_18531);
and U21965 (N_21965,N_18473,N_16016);
or U21966 (N_21966,N_18545,N_18085);
nand U21967 (N_21967,N_15503,N_16113);
or U21968 (N_21968,N_18647,N_16351);
nand U21969 (N_21969,N_19408,N_19812);
xnor U21970 (N_21970,N_17111,N_16191);
xnor U21971 (N_21971,N_18534,N_19002);
xnor U21972 (N_21972,N_19763,N_19309);
nor U21973 (N_21973,N_16606,N_16400);
and U21974 (N_21974,N_15957,N_15760);
nor U21975 (N_21975,N_17768,N_17418);
nand U21976 (N_21976,N_17823,N_16747);
and U21977 (N_21977,N_15268,N_17101);
and U21978 (N_21978,N_19458,N_16543);
and U21979 (N_21979,N_15889,N_15840);
nor U21980 (N_21980,N_17016,N_16144);
and U21981 (N_21981,N_19548,N_18630);
and U21982 (N_21982,N_19699,N_16408);
and U21983 (N_21983,N_17983,N_15761);
xor U21984 (N_21984,N_17907,N_19470);
xor U21985 (N_21985,N_18191,N_16642);
or U21986 (N_21986,N_16912,N_18175);
or U21987 (N_21987,N_15973,N_18851);
nor U21988 (N_21988,N_15417,N_18390);
nand U21989 (N_21989,N_15820,N_16529);
xor U21990 (N_21990,N_19881,N_17496);
or U21991 (N_21991,N_18658,N_16716);
nand U21992 (N_21992,N_19952,N_16795);
or U21993 (N_21993,N_17588,N_18615);
and U21994 (N_21994,N_16336,N_16974);
xor U21995 (N_21995,N_17806,N_17397);
or U21996 (N_21996,N_17827,N_17359);
xor U21997 (N_21997,N_18322,N_17683);
nor U21998 (N_21998,N_17643,N_17919);
nor U21999 (N_21999,N_19743,N_17360);
xnor U22000 (N_22000,N_18760,N_16550);
xnor U22001 (N_22001,N_18911,N_18549);
nor U22002 (N_22002,N_17201,N_18894);
nand U22003 (N_22003,N_16217,N_15323);
and U22004 (N_22004,N_18346,N_17312);
and U22005 (N_22005,N_15751,N_15049);
nor U22006 (N_22006,N_17664,N_18189);
and U22007 (N_22007,N_15217,N_19306);
and U22008 (N_22008,N_18261,N_15401);
xor U22009 (N_22009,N_16861,N_16933);
xnor U22010 (N_22010,N_18141,N_18686);
xor U22011 (N_22011,N_18304,N_18069);
nand U22012 (N_22012,N_18150,N_18268);
or U22013 (N_22013,N_17603,N_18497);
nor U22014 (N_22014,N_16454,N_18174);
xnor U22015 (N_22015,N_18904,N_17517);
nand U22016 (N_22016,N_15829,N_19948);
nor U22017 (N_22017,N_19295,N_19969);
xnor U22018 (N_22018,N_18699,N_18149);
nand U22019 (N_22019,N_18296,N_17920);
nor U22020 (N_22020,N_17544,N_15590);
and U22021 (N_22021,N_15676,N_15695);
nand U22022 (N_22022,N_19392,N_19322);
or U22023 (N_22023,N_16243,N_18563);
nand U22024 (N_22024,N_17266,N_16924);
nand U22025 (N_22025,N_15947,N_15452);
or U22026 (N_22026,N_17902,N_18762);
nor U22027 (N_22027,N_17022,N_19264);
nor U22028 (N_22028,N_15022,N_19827);
xor U22029 (N_22029,N_17566,N_19333);
and U22030 (N_22030,N_16076,N_17573);
or U22031 (N_22031,N_15815,N_18820);
and U22032 (N_22032,N_15146,N_15739);
xor U22033 (N_22033,N_16142,N_16922);
nor U22034 (N_22034,N_15787,N_17084);
xnor U22035 (N_22035,N_19499,N_18136);
xnor U22036 (N_22036,N_16029,N_19486);
and U22037 (N_22037,N_16028,N_16092);
xor U22038 (N_22038,N_18299,N_15540);
xor U22039 (N_22039,N_17918,N_17706);
nand U22040 (N_22040,N_17568,N_15093);
or U22041 (N_22041,N_19737,N_15004);
nand U22042 (N_22042,N_16103,N_19039);
nand U22043 (N_22043,N_17898,N_19516);
nor U22044 (N_22044,N_19097,N_15183);
and U22045 (N_22045,N_17767,N_15301);
nor U22046 (N_22046,N_19544,N_18086);
xor U22047 (N_22047,N_19637,N_15884);
nor U22048 (N_22048,N_16406,N_16067);
and U22049 (N_22049,N_19113,N_17871);
xor U22050 (N_22050,N_15950,N_19990);
xnor U22051 (N_22051,N_15944,N_16345);
xnor U22052 (N_22052,N_19036,N_15140);
and U22053 (N_22053,N_17154,N_15537);
nand U22054 (N_22054,N_15156,N_15509);
or U22055 (N_22055,N_15977,N_18648);
nand U22056 (N_22056,N_16857,N_17777);
xnor U22057 (N_22057,N_19893,N_19441);
nor U22058 (N_22058,N_15030,N_16305);
nand U22059 (N_22059,N_16149,N_19950);
and U22060 (N_22060,N_15384,N_17270);
nor U22061 (N_22061,N_15300,N_15835);
xnor U22062 (N_22062,N_16446,N_17155);
xnor U22063 (N_22063,N_19239,N_16246);
or U22064 (N_22064,N_18305,N_18594);
or U22065 (N_22065,N_16435,N_17086);
xnor U22066 (N_22066,N_16206,N_18319);
and U22067 (N_22067,N_16359,N_19648);
nand U22068 (N_22068,N_19837,N_16138);
or U22069 (N_22069,N_18926,N_15189);
nand U22070 (N_22070,N_16374,N_15463);
and U22071 (N_22071,N_18935,N_15292);
and U22072 (N_22072,N_16527,N_15427);
or U22073 (N_22073,N_18871,N_17632);
or U22074 (N_22074,N_16960,N_16802);
and U22075 (N_22075,N_17991,N_16235);
nand U22076 (N_22076,N_18730,N_18448);
nor U22077 (N_22077,N_17461,N_18413);
nand U22078 (N_22078,N_15628,N_15028);
nor U22079 (N_22079,N_16115,N_15484);
and U22080 (N_22080,N_15581,N_16353);
nand U22081 (N_22081,N_16378,N_19753);
or U22082 (N_22082,N_17145,N_19859);
nor U22083 (N_22083,N_16073,N_19405);
and U22084 (N_22084,N_16476,N_15777);
or U22085 (N_22085,N_17412,N_17075);
nand U22086 (N_22086,N_15356,N_17744);
nor U22087 (N_22087,N_19233,N_18747);
and U22088 (N_22088,N_16890,N_17414);
xor U22089 (N_22089,N_18677,N_18168);
xnor U22090 (N_22090,N_16358,N_16182);
nand U22091 (N_22091,N_19914,N_18854);
nand U22092 (N_22092,N_19273,N_16914);
and U22093 (N_22093,N_16551,N_16793);
or U22094 (N_22094,N_16722,N_16907);
and U22095 (N_22095,N_15241,N_17980);
and U22096 (N_22096,N_17608,N_19781);
xor U22097 (N_22097,N_19011,N_18124);
nand U22098 (N_22098,N_19359,N_16800);
xor U22099 (N_22099,N_17841,N_17349);
nand U22100 (N_22100,N_17763,N_17322);
nor U22101 (N_22101,N_15120,N_16832);
and U22102 (N_22102,N_15798,N_18664);
nand U22103 (N_22103,N_16654,N_17032);
nand U22104 (N_22104,N_17699,N_16486);
and U22105 (N_22105,N_17885,N_19086);
xor U22106 (N_22106,N_17565,N_16381);
and U22107 (N_22107,N_18057,N_19168);
and U22108 (N_22108,N_17708,N_18264);
nand U22109 (N_22109,N_19685,N_19649);
nor U22110 (N_22110,N_17379,N_15437);
xor U22111 (N_22111,N_16980,N_16898);
nor U22112 (N_22112,N_16553,N_16426);
nand U22113 (N_22113,N_18918,N_15180);
nand U22114 (N_22114,N_17720,N_17723);
and U22115 (N_22115,N_17047,N_19899);
nor U22116 (N_22116,N_16689,N_16611);
nand U22117 (N_22117,N_15746,N_17733);
and U22118 (N_22118,N_18017,N_19739);
nor U22119 (N_22119,N_18314,N_18950);
nand U22120 (N_22120,N_18482,N_18848);
nand U22121 (N_22121,N_17837,N_15175);
and U22122 (N_22122,N_16299,N_17241);
or U22123 (N_22123,N_17506,N_17690);
or U22124 (N_22124,N_15309,N_17061);
or U22125 (N_22125,N_15178,N_15043);
nand U22126 (N_22126,N_17423,N_18003);
or U22127 (N_22127,N_17066,N_15182);
or U22128 (N_22128,N_18046,N_16780);
nand U22129 (N_22129,N_15128,N_15242);
and U22130 (N_22130,N_18108,N_19212);
nor U22131 (N_22131,N_18438,N_19591);
or U22132 (N_22132,N_15224,N_15595);
xor U22133 (N_22133,N_19089,N_16856);
nor U22134 (N_22134,N_15435,N_19193);
nor U22135 (N_22135,N_15624,N_16817);
nand U22136 (N_22136,N_19218,N_17351);
and U22137 (N_22137,N_18705,N_18587);
or U22138 (N_22138,N_19994,N_16863);
xor U22139 (N_22139,N_15641,N_16572);
or U22140 (N_22140,N_16259,N_15933);
nand U22141 (N_22141,N_15137,N_18034);
or U22142 (N_22142,N_16433,N_18252);
xor U22143 (N_22143,N_15657,N_18910);
or U22144 (N_22144,N_19229,N_17528);
nor U22145 (N_22145,N_18865,N_19967);
and U22146 (N_22146,N_19611,N_17063);
xor U22147 (N_22147,N_15688,N_17546);
or U22148 (N_22148,N_18538,N_15858);
and U22149 (N_22149,N_18011,N_17999);
and U22150 (N_22150,N_18810,N_17834);
and U22151 (N_22151,N_15282,N_15166);
or U22152 (N_22152,N_17048,N_18067);
and U22153 (N_22153,N_19227,N_17532);
or U22154 (N_22154,N_19809,N_16783);
or U22155 (N_22155,N_16671,N_18260);
xnor U22156 (N_22156,N_19344,N_16168);
and U22157 (N_22157,N_16686,N_17131);
nand U22158 (N_22158,N_16465,N_19600);
nand U22159 (N_22159,N_19269,N_16065);
nand U22160 (N_22160,N_17928,N_18178);
or U22161 (N_22161,N_17626,N_16940);
or U22162 (N_22162,N_15758,N_15014);
or U22163 (N_22163,N_19370,N_19814);
and U22164 (N_22164,N_17317,N_15714);
xnor U22165 (N_22165,N_16043,N_18266);
nor U22166 (N_22166,N_16037,N_19705);
and U22167 (N_22167,N_18435,N_16427);
xor U22168 (N_22168,N_17862,N_17275);
nor U22169 (N_22169,N_18582,N_19482);
nand U22170 (N_22170,N_17400,N_18764);
nor U22171 (N_22171,N_16352,N_16620);
xnor U22172 (N_22172,N_18444,N_16032);
xor U22173 (N_22173,N_15554,N_16503);
nor U22174 (N_22174,N_15106,N_16329);
or U22175 (N_22175,N_15174,N_15289);
or U22176 (N_22176,N_17021,N_18845);
nand U22177 (N_22177,N_15260,N_17994);
nor U22178 (N_22178,N_16475,N_17186);
nor U22179 (N_22179,N_18556,N_19378);
xor U22180 (N_22180,N_17267,N_18359);
or U22181 (N_22181,N_18376,N_15479);
nand U22182 (N_22182,N_16124,N_19854);
nor U22183 (N_22183,N_19045,N_19154);
xor U22184 (N_22184,N_19209,N_18401);
nand U22185 (N_22185,N_18625,N_15481);
and U22186 (N_22186,N_19380,N_18806);
or U22187 (N_22187,N_15263,N_19586);
and U22188 (N_22188,N_18073,N_17058);
or U22189 (N_22189,N_16545,N_15303);
nor U22190 (N_22190,N_17592,N_16913);
nand U22191 (N_22191,N_16741,N_15066);
nand U22192 (N_22192,N_18353,N_15065);
nor U22193 (N_22193,N_15199,N_18588);
nand U22194 (N_22194,N_17558,N_15630);
xnor U22195 (N_22195,N_18395,N_18886);
xor U22196 (N_22196,N_17615,N_18134);
nand U22197 (N_22197,N_18619,N_18942);
and U22198 (N_22198,N_16682,N_17969);
xor U22199 (N_22199,N_16632,N_16684);
nor U22200 (N_22200,N_19819,N_16220);
or U22201 (N_22201,N_15499,N_18768);
or U22202 (N_22202,N_15682,N_18244);
nor U22203 (N_22203,N_16688,N_16859);
and U22204 (N_22204,N_18833,N_17570);
nand U22205 (N_22205,N_17838,N_19296);
xnor U22206 (N_22206,N_18869,N_15338);
or U22207 (N_22207,N_19396,N_17142);
xor U22208 (N_22208,N_17279,N_16608);
nand U22209 (N_22209,N_18182,N_16652);
or U22210 (N_22210,N_15801,N_18156);
or U22211 (N_22211,N_18899,N_17187);
nand U22212 (N_22212,N_18691,N_19918);
or U22213 (N_22213,N_15890,N_16662);
nand U22214 (N_22214,N_18449,N_18626);
and U22215 (N_22215,N_17758,N_19867);
nand U22216 (N_22216,N_19992,N_18996);
and U22217 (N_22217,N_16320,N_15603);
and U22218 (N_22218,N_18267,N_19014);
nor U22219 (N_22219,N_18576,N_19316);
and U22220 (N_22220,N_19237,N_16130);
nor U22221 (N_22221,N_16769,N_16561);
xor U22222 (N_22222,N_17742,N_16542);
nor U22223 (N_22223,N_18589,N_16104);
and U22224 (N_22224,N_19733,N_17481);
or U22225 (N_22225,N_19160,N_19560);
nand U22226 (N_22226,N_17801,N_16496);
and U22227 (N_22227,N_18199,N_19181);
nand U22228 (N_22228,N_19496,N_16482);
nand U22229 (N_22229,N_15514,N_16160);
xnor U22230 (N_22230,N_19632,N_18799);
nor U22231 (N_22231,N_16592,N_16634);
or U22232 (N_22232,N_15411,N_19076);
xor U22233 (N_22233,N_17601,N_19413);
nand U22234 (N_22234,N_19493,N_19304);
nor U22235 (N_22235,N_15691,N_18181);
xnor U22236 (N_22236,N_18995,N_16713);
and U22237 (N_22237,N_19640,N_18160);
xnor U22238 (N_22238,N_17912,N_19406);
xnor U22239 (N_22239,N_15671,N_19348);
xnor U22240 (N_22240,N_15402,N_17487);
xnor U22241 (N_22241,N_19299,N_19567);
nand U22242 (N_22242,N_17249,N_16510);
nor U22243 (N_22243,N_17972,N_18477);
nand U22244 (N_22244,N_18597,N_19155);
or U22245 (N_22245,N_19679,N_19119);
nor U22246 (N_22246,N_16333,N_18392);
and U22247 (N_22247,N_15652,N_15103);
xor U22248 (N_22248,N_15773,N_19787);
nor U22249 (N_22249,N_19772,N_19285);
or U22250 (N_22250,N_16807,N_15426);
or U22251 (N_22251,N_19688,N_19121);
nand U22252 (N_22252,N_19775,N_17402);
and U22253 (N_22253,N_15497,N_18426);
and U22254 (N_22254,N_18004,N_15018);
nor U22255 (N_22255,N_17358,N_19262);
xnor U22256 (N_22256,N_18119,N_17090);
xnor U22257 (N_22257,N_19084,N_17828);
nand U22258 (N_22258,N_16242,N_15256);
xor U22259 (N_22259,N_18125,N_15567);
or U22260 (N_22260,N_15639,N_18616);
nand U22261 (N_22261,N_17462,N_16171);
or U22262 (N_22262,N_19555,N_18998);
nand U22263 (N_22263,N_17889,N_15134);
nand U22264 (N_22264,N_19021,N_17845);
nand U22265 (N_22265,N_19937,N_19454);
and U22266 (N_22266,N_17600,N_18452);
nand U22267 (N_22267,N_16973,N_17939);
xnor U22268 (N_22268,N_16404,N_19346);
xnor U22269 (N_22269,N_16434,N_16892);
xor U22270 (N_22270,N_19007,N_19802);
or U22271 (N_22271,N_19989,N_17598);
and U22272 (N_22272,N_15381,N_16509);
and U22273 (N_22273,N_18661,N_19891);
nand U22274 (N_22274,N_16021,N_16773);
nor U22275 (N_22275,N_17156,N_17259);
nor U22276 (N_22276,N_15909,N_18994);
or U22277 (N_22277,N_16450,N_17830);
nor U22278 (N_22278,N_18163,N_18893);
and U22279 (N_22279,N_15412,N_15730);
or U22280 (N_22280,N_15454,N_15516);
nand U22281 (N_22281,N_17372,N_19335);
and U22282 (N_22282,N_18930,N_19539);
and U22283 (N_22283,N_18356,N_18235);
xor U22284 (N_22284,N_17554,N_19535);
or U22285 (N_22285,N_19182,N_19062);
nor U22286 (N_22286,N_16833,N_19226);
or U22287 (N_22287,N_17469,N_15640);
or U22288 (N_22288,N_18569,N_17313);
xor U22289 (N_22289,N_16195,N_19416);
nor U22290 (N_22290,N_17678,N_18117);
nand U22291 (N_22291,N_15939,N_19594);
nand U22292 (N_22292,N_17463,N_16175);
nand U22293 (N_22293,N_16964,N_15446);
or U22294 (N_22294,N_18813,N_18415);
xnor U22295 (N_22295,N_17614,N_19657);
xnor U22296 (N_22296,N_16888,N_18489);
nor U22297 (N_22297,N_16445,N_19016);
xnor U22298 (N_22298,N_16178,N_15138);
nor U22299 (N_22299,N_19191,N_17645);
nand U22300 (N_22300,N_17854,N_15568);
or U22301 (N_22301,N_18750,N_19298);
or U22302 (N_22302,N_15847,N_19046);
or U22303 (N_22303,N_15317,N_16466);
or U22304 (N_22304,N_15654,N_19137);
nand U22305 (N_22305,N_16788,N_16003);
nand U22306 (N_22306,N_15405,N_18723);
or U22307 (N_22307,N_18979,N_18574);
nor U22308 (N_22308,N_19423,N_17103);
xor U22309 (N_22309,N_17878,N_16499);
nor U22310 (N_22310,N_17770,N_16700);
and U22311 (N_22311,N_19134,N_16842);
and U22312 (N_22312,N_19038,N_18634);
nor U22313 (N_22313,N_18056,N_18183);
and U22314 (N_22314,N_19140,N_15438);
or U22315 (N_22315,N_17491,N_17362);
or U22316 (N_22316,N_18789,N_19500);
xnor U22317 (N_22317,N_15845,N_19773);
xnor U22318 (N_22318,N_19862,N_15715);
nor U22319 (N_22319,N_19786,N_18481);
and U22320 (N_22320,N_15226,N_16714);
or U22321 (N_22321,N_19729,N_16126);
nor U22322 (N_22322,N_17431,N_19473);
nand U22323 (N_22323,N_19974,N_16062);
or U22324 (N_22324,N_16570,N_17184);
and U22325 (N_22325,N_16049,N_16535);
or U22326 (N_22326,N_19508,N_17326);
xnor U22327 (N_22327,N_15892,N_17329);
xor U22328 (N_22328,N_18745,N_17746);
nor U22329 (N_22329,N_18317,N_19071);
nand U22330 (N_22330,N_15955,N_16696);
and U22331 (N_22331,N_15458,N_16107);
nand U22332 (N_22332,N_19429,N_18409);
or U22333 (N_22333,N_15010,N_19607);
nor U22334 (N_22334,N_17368,N_15813);
xnor U22335 (N_22335,N_15001,N_19929);
nand U22336 (N_22336,N_18068,N_19043);
nand U22337 (N_22337,N_18372,N_16471);
nor U22338 (N_22338,N_18315,N_16719);
nor U22339 (N_22339,N_18371,N_17138);
or U22340 (N_22340,N_16573,N_19731);
xor U22341 (N_22341,N_17637,N_15596);
xnor U22342 (N_22342,N_19446,N_18389);
xor U22343 (N_22343,N_17054,N_15318);
xor U22344 (N_22344,N_18732,N_15991);
xnor U22345 (N_22345,N_19376,N_18019);
or U22346 (N_22346,N_19107,N_18079);
and U22347 (N_22347,N_19149,N_15465);
and U22348 (N_22348,N_18525,N_15117);
and U22349 (N_22349,N_19631,N_19629);
nor U22350 (N_22350,N_16945,N_16771);
xnor U22351 (N_22351,N_16687,N_16398);
xnor U22352 (N_22352,N_18495,N_18263);
xnor U22353 (N_22353,N_18702,N_19443);
xor U22354 (N_22354,N_16207,N_16755);
nand U22355 (N_22355,N_17846,N_17427);
nand U22356 (N_22356,N_15333,N_18895);
nand U22357 (N_22357,N_15988,N_18044);
xnor U22358 (N_22358,N_17560,N_18208);
nand U22359 (N_22359,N_15216,N_16643);
nand U22360 (N_22360,N_15919,N_15012);
nor U22361 (N_22361,N_16383,N_18335);
nand U22362 (N_22362,N_17968,N_19127);
nand U22363 (N_22363,N_17323,N_16302);
nor U22364 (N_22364,N_15665,N_19015);
nand U22365 (N_22365,N_19324,N_15745);
nand U22366 (N_22366,N_18779,N_15116);
and U22367 (N_22367,N_16059,N_19402);
xnor U22368 (N_22368,N_16533,N_15169);
nor U22369 (N_22369,N_19576,N_19521);
nor U22370 (N_22370,N_15032,N_15234);
or U22371 (N_22371,N_18560,N_18411);
or U22372 (N_22372,N_18273,N_18988);
nor U22373 (N_22373,N_17893,N_17711);
xor U22374 (N_22374,N_16556,N_19866);
nor U22375 (N_22375,N_16749,N_15754);
and U22376 (N_22376,N_15677,N_17160);
nor U22377 (N_22377,N_18246,N_18682);
nor U22378 (N_22378,N_16724,N_19419);
nor U22379 (N_22379,N_18408,N_18470);
and U22380 (N_22380,N_18509,N_17116);
or U22381 (N_22381,N_17585,N_15413);
nand U22382 (N_22382,N_19791,N_17204);
nor U22383 (N_22383,N_19537,N_19223);
and U22384 (N_22384,N_18523,N_19903);
nor U22385 (N_22385,N_18114,N_18786);
nand U22386 (N_22386,N_18853,N_17789);
nand U22387 (N_22387,N_18518,N_15700);
xnor U22388 (N_22388,N_19124,N_15389);
nor U22389 (N_22389,N_16409,N_16942);
nor U22390 (N_22390,N_18776,N_16360);
or U22391 (N_22391,N_15831,N_18427);
nand U22392 (N_22392,N_19253,N_19130);
nor U22393 (N_22393,N_18311,N_16854);
nor U22394 (N_22394,N_16680,N_18783);
xnor U22395 (N_22395,N_19349,N_17771);
xor U22396 (N_22396,N_17452,N_19329);
and U22397 (N_22397,N_17775,N_19844);
nand U22398 (N_22398,N_19300,N_15882);
xnor U22399 (N_22399,N_16280,N_19682);
nor U22400 (N_22400,N_16214,N_15490);
and U22401 (N_22401,N_16878,N_17844);
xnor U22402 (N_22402,N_15828,N_18351);
or U22403 (N_22403,N_18628,N_19614);
and U22404 (N_22404,N_17023,N_17739);
xor U22405 (N_22405,N_15750,N_16293);
and U22406 (N_22406,N_18396,N_17395);
and U22407 (N_22407,N_19653,N_18758);
or U22408 (N_22408,N_15016,N_16965);
xor U22409 (N_22409,N_16325,N_19816);
xor U22410 (N_22410,N_17444,N_19590);
and U22411 (N_22411,N_18039,N_19356);
or U22412 (N_22412,N_19524,N_17849);
nor U22413 (N_22413,N_19000,N_16109);
nor U22414 (N_22414,N_18196,N_16565);
xnor U22415 (N_22415,N_15511,N_18962);
nand U22416 (N_22416,N_16794,N_18130);
nor U22417 (N_22417,N_18554,N_15931);
nand U22418 (N_22418,N_18041,N_17539);
nor U22419 (N_22419,N_17754,N_15837);
xor U22420 (N_22420,N_19246,N_17302);
or U22421 (N_22421,N_15378,N_17508);
nor U22422 (N_22422,N_15243,N_19410);
or U22423 (N_22423,N_15880,N_16348);
or U22424 (N_22424,N_15794,N_19184);
xor U22425 (N_22425,N_16082,N_17833);
and U22426 (N_22426,N_19824,N_17380);
nor U22427 (N_22427,N_15894,N_17694);
or U22428 (N_22428,N_18198,N_19289);
nor U22429 (N_22429,N_17369,N_15418);
or U22430 (N_22430,N_15557,N_18271);
or U22431 (N_22431,N_17311,N_18663);
xor U22432 (N_22432,N_19056,N_18941);
or U22433 (N_22433,N_16599,N_19534);
nand U22434 (N_22434,N_16321,N_15118);
xor U22435 (N_22435,N_19109,N_17292);
nand U22436 (N_22436,N_17314,N_19965);
nor U22437 (N_22437,N_18066,N_19906);
or U22438 (N_22438,N_19497,N_16008);
and U22439 (N_22439,N_19358,N_18581);
xor U22440 (N_22440,N_18298,N_19620);
and U22441 (N_22441,N_18496,N_15597);
xnor U22442 (N_22442,N_16801,N_19228);
or U22443 (N_22443,N_17121,N_17493);
and U22444 (N_22444,N_17246,N_19479);
nor U22445 (N_22445,N_17897,N_19081);
or U22446 (N_22446,N_15082,N_17876);
nor U22447 (N_22447,N_19829,N_17717);
or U22448 (N_22448,N_15011,N_15969);
nand U22449 (N_22449,N_19031,N_15545);
and U22450 (N_22450,N_18715,N_15098);
nor U22451 (N_22451,N_17676,N_19882);
and U22452 (N_22452,N_15074,N_15332);
or U22453 (N_22453,N_15763,N_19796);
nor U22454 (N_22454,N_18707,N_16441);
xor U22455 (N_22455,N_18352,N_15212);
nand U22456 (N_22456,N_19817,N_19798);
xnor U22457 (N_22457,N_16081,N_17405);
or U22458 (N_22458,N_19717,N_19766);
and U22459 (N_22459,N_19673,N_16900);
and U22460 (N_22460,N_18889,N_16338);
and U22461 (N_22461,N_15013,N_15046);
or U22462 (N_22462,N_15549,N_15534);
nor U22463 (N_22463,N_18320,N_18326);
nand U22464 (N_22464,N_16613,N_16068);
or U22465 (N_22465,N_17703,N_16250);
xor U22466 (N_22466,N_17964,N_16412);
and U22467 (N_22467,N_18632,N_15563);
or U22468 (N_22468,N_19720,N_18350);
nor U22469 (N_22469,N_15430,N_15546);
nor U22470 (N_22470,N_16165,N_15926);
and U22471 (N_22471,N_15273,N_18816);
nor U22472 (N_22472,N_18101,N_17731);
xor U22473 (N_22473,N_16439,N_17861);
xor U22474 (N_22474,N_15009,N_17839);
and U22475 (N_22475,N_17516,N_16969);
and U22476 (N_22476,N_15602,N_16041);
nor U22477 (N_22477,N_18269,N_19178);
xor U22478 (N_22478,N_17430,N_16258);
xnor U22479 (N_22479,N_18567,N_17309);
nand U22480 (N_22480,N_18161,N_18565);
nand U22481 (N_22481,N_19502,N_15625);
nand U22482 (N_22482,N_18983,N_15644);
nor U22483 (N_22483,N_16017,N_16420);
nand U22484 (N_22484,N_18087,N_17123);
nor U22485 (N_22485,N_18469,N_19880);
and U22486 (N_22486,N_17475,N_16579);
or U22487 (N_22487,N_16498,N_17660);
xor U22488 (N_22488,N_15311,N_19779);
nor U22489 (N_22489,N_16519,N_18627);
or U22490 (N_22490,N_17652,N_19943);
xnor U22491 (N_22491,N_17840,N_19099);
nor U22492 (N_22492,N_16628,N_15930);
or U22493 (N_22493,N_15854,N_18110);
nand U22494 (N_22494,N_19489,N_18393);
xnor U22495 (N_22495,N_17133,N_19382);
nor U22496 (N_22496,N_15893,N_15219);
xnor U22497 (N_22497,N_19584,N_19856);
xor U22498 (N_22498,N_15795,N_17205);
nand U22499 (N_22499,N_16256,N_17304);
and U22500 (N_22500,N_19206,N_19211);
or U22501 (N_22501,N_16317,N_16017);
or U22502 (N_22502,N_17919,N_15494);
nor U22503 (N_22503,N_17294,N_19766);
xor U22504 (N_22504,N_15696,N_19672);
xor U22505 (N_22505,N_17436,N_18872);
xor U22506 (N_22506,N_19625,N_19486);
nand U22507 (N_22507,N_18713,N_19816);
and U22508 (N_22508,N_17160,N_16414);
and U22509 (N_22509,N_19763,N_15892);
nor U22510 (N_22510,N_17163,N_17638);
nand U22511 (N_22511,N_17663,N_15579);
nand U22512 (N_22512,N_15683,N_15358);
xor U22513 (N_22513,N_16379,N_15988);
nand U22514 (N_22514,N_19246,N_17788);
and U22515 (N_22515,N_17642,N_16275);
or U22516 (N_22516,N_15024,N_15430);
nand U22517 (N_22517,N_19906,N_18006);
nor U22518 (N_22518,N_16735,N_18451);
nand U22519 (N_22519,N_15466,N_19494);
nor U22520 (N_22520,N_19023,N_15545);
nor U22521 (N_22521,N_18198,N_19207);
nand U22522 (N_22522,N_15948,N_15918);
nor U22523 (N_22523,N_15659,N_15262);
xor U22524 (N_22524,N_17028,N_16013);
and U22525 (N_22525,N_17088,N_15031);
xor U22526 (N_22526,N_16665,N_17323);
xor U22527 (N_22527,N_16337,N_16725);
nor U22528 (N_22528,N_18413,N_19555);
nand U22529 (N_22529,N_16367,N_16567);
nand U22530 (N_22530,N_16153,N_17087);
xnor U22531 (N_22531,N_18509,N_18715);
xor U22532 (N_22532,N_18792,N_15337);
nand U22533 (N_22533,N_16624,N_15903);
nor U22534 (N_22534,N_16216,N_16950);
nor U22535 (N_22535,N_18759,N_16959);
and U22536 (N_22536,N_19413,N_18376);
xnor U22537 (N_22537,N_16731,N_17399);
and U22538 (N_22538,N_16922,N_18492);
nand U22539 (N_22539,N_17996,N_16753);
or U22540 (N_22540,N_15927,N_15724);
xor U22541 (N_22541,N_17194,N_15369);
nor U22542 (N_22542,N_18577,N_15279);
xor U22543 (N_22543,N_16784,N_16849);
nand U22544 (N_22544,N_17018,N_18717);
and U22545 (N_22545,N_15810,N_19339);
nand U22546 (N_22546,N_17295,N_19594);
xor U22547 (N_22547,N_16176,N_18389);
or U22548 (N_22548,N_16514,N_19263);
nand U22549 (N_22549,N_18236,N_16139);
nand U22550 (N_22550,N_17051,N_17408);
nor U22551 (N_22551,N_15234,N_16998);
xor U22552 (N_22552,N_15798,N_19204);
nand U22553 (N_22553,N_17872,N_18422);
xor U22554 (N_22554,N_18596,N_17394);
or U22555 (N_22555,N_15012,N_18001);
xnor U22556 (N_22556,N_15878,N_19769);
xnor U22557 (N_22557,N_19821,N_16997);
nor U22558 (N_22558,N_15813,N_18821);
and U22559 (N_22559,N_16603,N_17110);
and U22560 (N_22560,N_18108,N_18481);
xor U22561 (N_22561,N_16181,N_15276);
or U22562 (N_22562,N_15387,N_18272);
and U22563 (N_22563,N_18588,N_17867);
or U22564 (N_22564,N_16317,N_19377);
nor U22565 (N_22565,N_19738,N_15320);
or U22566 (N_22566,N_16312,N_16571);
and U22567 (N_22567,N_15910,N_19364);
nand U22568 (N_22568,N_19243,N_18939);
xor U22569 (N_22569,N_16626,N_19646);
nand U22570 (N_22570,N_19229,N_18016);
nor U22571 (N_22571,N_17469,N_19879);
and U22572 (N_22572,N_15273,N_18205);
or U22573 (N_22573,N_16053,N_19973);
and U22574 (N_22574,N_15976,N_17213);
or U22575 (N_22575,N_19436,N_15262);
xnor U22576 (N_22576,N_17237,N_15964);
or U22577 (N_22577,N_18827,N_17179);
nand U22578 (N_22578,N_18881,N_15161);
xor U22579 (N_22579,N_19301,N_19095);
nor U22580 (N_22580,N_18195,N_15678);
nand U22581 (N_22581,N_17635,N_15170);
or U22582 (N_22582,N_16023,N_18837);
xnor U22583 (N_22583,N_18500,N_15211);
or U22584 (N_22584,N_18676,N_19188);
xnor U22585 (N_22585,N_15920,N_15768);
and U22586 (N_22586,N_16490,N_19848);
xnor U22587 (N_22587,N_18013,N_15835);
or U22588 (N_22588,N_19112,N_16319);
nand U22589 (N_22589,N_17508,N_17747);
nand U22590 (N_22590,N_15003,N_19544);
xnor U22591 (N_22591,N_17792,N_15867);
xnor U22592 (N_22592,N_15405,N_15508);
xnor U22593 (N_22593,N_19019,N_16316);
nor U22594 (N_22594,N_18463,N_16850);
and U22595 (N_22595,N_18273,N_18918);
nor U22596 (N_22596,N_18557,N_18655);
xor U22597 (N_22597,N_19995,N_17168);
and U22598 (N_22598,N_18356,N_19872);
nor U22599 (N_22599,N_16553,N_18528);
or U22600 (N_22600,N_16340,N_17788);
nand U22601 (N_22601,N_16876,N_19222);
or U22602 (N_22602,N_17868,N_18619);
nor U22603 (N_22603,N_19828,N_16760);
nor U22604 (N_22604,N_17425,N_15468);
and U22605 (N_22605,N_18428,N_16719);
or U22606 (N_22606,N_16445,N_16480);
and U22607 (N_22607,N_19327,N_18526);
nand U22608 (N_22608,N_15993,N_19007);
and U22609 (N_22609,N_18704,N_18500);
or U22610 (N_22610,N_15357,N_15884);
or U22611 (N_22611,N_15675,N_17686);
nand U22612 (N_22612,N_17317,N_17375);
nor U22613 (N_22613,N_18162,N_19764);
nand U22614 (N_22614,N_17051,N_17294);
or U22615 (N_22615,N_19997,N_18478);
nor U22616 (N_22616,N_17138,N_16804);
nor U22617 (N_22617,N_19103,N_18471);
xor U22618 (N_22618,N_18246,N_15725);
or U22619 (N_22619,N_15950,N_16891);
xor U22620 (N_22620,N_15058,N_15307);
nand U22621 (N_22621,N_19716,N_18568);
xor U22622 (N_22622,N_19782,N_18180);
nand U22623 (N_22623,N_15300,N_15980);
and U22624 (N_22624,N_19587,N_15456);
nand U22625 (N_22625,N_19001,N_18841);
xor U22626 (N_22626,N_16932,N_18337);
or U22627 (N_22627,N_15155,N_15935);
or U22628 (N_22628,N_16773,N_18016);
nor U22629 (N_22629,N_18880,N_15914);
nand U22630 (N_22630,N_19007,N_18585);
nand U22631 (N_22631,N_15096,N_16633);
xnor U22632 (N_22632,N_19759,N_16172);
and U22633 (N_22633,N_19015,N_16718);
or U22634 (N_22634,N_17583,N_18435);
and U22635 (N_22635,N_16707,N_15400);
nor U22636 (N_22636,N_19819,N_16343);
nand U22637 (N_22637,N_18172,N_17851);
or U22638 (N_22638,N_15555,N_15735);
nor U22639 (N_22639,N_16242,N_18624);
nand U22640 (N_22640,N_17090,N_17949);
xnor U22641 (N_22641,N_19656,N_18575);
and U22642 (N_22642,N_19664,N_18408);
and U22643 (N_22643,N_15731,N_16849);
and U22644 (N_22644,N_16377,N_18269);
nor U22645 (N_22645,N_16259,N_15589);
xor U22646 (N_22646,N_18961,N_19446);
nand U22647 (N_22647,N_15075,N_17389);
nand U22648 (N_22648,N_19496,N_19602);
or U22649 (N_22649,N_15090,N_17216);
or U22650 (N_22650,N_16191,N_16923);
xor U22651 (N_22651,N_16589,N_19646);
nand U22652 (N_22652,N_15076,N_18051);
or U22653 (N_22653,N_19740,N_18755);
xnor U22654 (N_22654,N_17354,N_19373);
or U22655 (N_22655,N_19227,N_15589);
or U22656 (N_22656,N_15735,N_18330);
and U22657 (N_22657,N_16751,N_17923);
nand U22658 (N_22658,N_15638,N_19171);
and U22659 (N_22659,N_19409,N_18526);
or U22660 (N_22660,N_18796,N_15014);
and U22661 (N_22661,N_18715,N_15736);
xor U22662 (N_22662,N_19578,N_15827);
nor U22663 (N_22663,N_17623,N_19119);
xor U22664 (N_22664,N_18479,N_15358);
and U22665 (N_22665,N_15612,N_17412);
xnor U22666 (N_22666,N_19549,N_17350);
xnor U22667 (N_22667,N_19604,N_19682);
nand U22668 (N_22668,N_16342,N_18491);
or U22669 (N_22669,N_16782,N_18405);
nand U22670 (N_22670,N_16561,N_18889);
or U22671 (N_22671,N_15479,N_17635);
xor U22672 (N_22672,N_18330,N_15141);
nand U22673 (N_22673,N_17561,N_15933);
nor U22674 (N_22674,N_15115,N_16652);
and U22675 (N_22675,N_17368,N_17934);
nor U22676 (N_22676,N_15219,N_19045);
xor U22677 (N_22677,N_18315,N_17711);
nor U22678 (N_22678,N_15946,N_16897);
nand U22679 (N_22679,N_19511,N_19569);
nor U22680 (N_22680,N_15014,N_19645);
and U22681 (N_22681,N_19557,N_16745);
or U22682 (N_22682,N_17926,N_18684);
nand U22683 (N_22683,N_18563,N_15544);
and U22684 (N_22684,N_17968,N_19437);
and U22685 (N_22685,N_19530,N_15128);
nand U22686 (N_22686,N_19028,N_16455);
nand U22687 (N_22687,N_17950,N_16294);
or U22688 (N_22688,N_18021,N_15243);
xnor U22689 (N_22689,N_15628,N_18469);
nand U22690 (N_22690,N_19259,N_18299);
nor U22691 (N_22691,N_16081,N_17168);
nor U22692 (N_22692,N_17937,N_15444);
nand U22693 (N_22693,N_19326,N_19670);
and U22694 (N_22694,N_17503,N_15338);
xnor U22695 (N_22695,N_17812,N_15559);
xnor U22696 (N_22696,N_15697,N_17882);
nor U22697 (N_22697,N_19891,N_18536);
nand U22698 (N_22698,N_17965,N_17798);
or U22699 (N_22699,N_18543,N_16037);
nor U22700 (N_22700,N_19788,N_18711);
xnor U22701 (N_22701,N_17342,N_16435);
nor U22702 (N_22702,N_19779,N_15411);
or U22703 (N_22703,N_16294,N_16567);
and U22704 (N_22704,N_19388,N_18205);
or U22705 (N_22705,N_15913,N_19337);
xor U22706 (N_22706,N_18032,N_18977);
nand U22707 (N_22707,N_15997,N_18726);
nand U22708 (N_22708,N_18355,N_16237);
and U22709 (N_22709,N_18135,N_15824);
nand U22710 (N_22710,N_16085,N_17229);
or U22711 (N_22711,N_16703,N_19591);
nor U22712 (N_22712,N_15068,N_17239);
nand U22713 (N_22713,N_19417,N_17363);
nor U22714 (N_22714,N_16827,N_18877);
nand U22715 (N_22715,N_18555,N_16483);
nand U22716 (N_22716,N_17395,N_18876);
or U22717 (N_22717,N_17676,N_19496);
xor U22718 (N_22718,N_19564,N_16095);
and U22719 (N_22719,N_16581,N_16371);
or U22720 (N_22720,N_17794,N_19319);
or U22721 (N_22721,N_17638,N_15915);
nor U22722 (N_22722,N_19005,N_18641);
xnor U22723 (N_22723,N_16311,N_19652);
xor U22724 (N_22724,N_15701,N_17235);
or U22725 (N_22725,N_15360,N_16146);
nor U22726 (N_22726,N_17487,N_16224);
xnor U22727 (N_22727,N_19229,N_19718);
nand U22728 (N_22728,N_17200,N_17307);
nor U22729 (N_22729,N_15338,N_17560);
nor U22730 (N_22730,N_19042,N_17150);
and U22731 (N_22731,N_18860,N_15871);
nor U22732 (N_22732,N_15295,N_18755);
nor U22733 (N_22733,N_17402,N_16459);
and U22734 (N_22734,N_18068,N_16502);
xnor U22735 (N_22735,N_19810,N_17433);
nand U22736 (N_22736,N_15023,N_19820);
xnor U22737 (N_22737,N_19168,N_17747);
nor U22738 (N_22738,N_15179,N_19097);
nand U22739 (N_22739,N_18720,N_19626);
nand U22740 (N_22740,N_15704,N_16527);
xor U22741 (N_22741,N_17018,N_19463);
nand U22742 (N_22742,N_18561,N_16860);
xor U22743 (N_22743,N_18829,N_18510);
and U22744 (N_22744,N_15922,N_19480);
xnor U22745 (N_22745,N_16490,N_18458);
or U22746 (N_22746,N_18482,N_17771);
nand U22747 (N_22747,N_19730,N_16281);
nand U22748 (N_22748,N_15504,N_18543);
nor U22749 (N_22749,N_17864,N_18459);
nand U22750 (N_22750,N_19909,N_19424);
xnor U22751 (N_22751,N_17675,N_15598);
xnor U22752 (N_22752,N_19212,N_16756);
xor U22753 (N_22753,N_16903,N_15380);
xnor U22754 (N_22754,N_15849,N_16437);
nand U22755 (N_22755,N_16670,N_16039);
and U22756 (N_22756,N_19755,N_16483);
or U22757 (N_22757,N_17482,N_16641);
nand U22758 (N_22758,N_16906,N_18507);
xnor U22759 (N_22759,N_17876,N_16397);
xnor U22760 (N_22760,N_17365,N_19213);
xnor U22761 (N_22761,N_19922,N_17837);
nor U22762 (N_22762,N_16736,N_18952);
nand U22763 (N_22763,N_17585,N_17327);
nor U22764 (N_22764,N_15290,N_18680);
and U22765 (N_22765,N_17959,N_15032);
xor U22766 (N_22766,N_18522,N_17069);
nand U22767 (N_22767,N_17676,N_17591);
xor U22768 (N_22768,N_17201,N_15921);
xnor U22769 (N_22769,N_18593,N_15410);
nor U22770 (N_22770,N_17824,N_17381);
or U22771 (N_22771,N_19139,N_17971);
nand U22772 (N_22772,N_17596,N_18482);
xnor U22773 (N_22773,N_18630,N_15549);
and U22774 (N_22774,N_16924,N_17021);
or U22775 (N_22775,N_18007,N_16312);
or U22776 (N_22776,N_16975,N_19001);
xnor U22777 (N_22777,N_15047,N_15642);
xnor U22778 (N_22778,N_18428,N_16244);
nand U22779 (N_22779,N_16554,N_15036);
xnor U22780 (N_22780,N_18817,N_15738);
nand U22781 (N_22781,N_17244,N_19824);
nand U22782 (N_22782,N_15486,N_17293);
and U22783 (N_22783,N_16842,N_19391);
and U22784 (N_22784,N_15960,N_15189);
nor U22785 (N_22785,N_17632,N_17094);
nand U22786 (N_22786,N_15869,N_18388);
and U22787 (N_22787,N_16562,N_17801);
nor U22788 (N_22788,N_16133,N_19004);
nand U22789 (N_22789,N_15575,N_19435);
or U22790 (N_22790,N_16339,N_19231);
nor U22791 (N_22791,N_18168,N_19391);
or U22792 (N_22792,N_16468,N_15127);
xnor U22793 (N_22793,N_19604,N_17038);
xor U22794 (N_22794,N_17436,N_15842);
nor U22795 (N_22795,N_17479,N_18334);
nor U22796 (N_22796,N_19251,N_16302);
xor U22797 (N_22797,N_18093,N_18986);
or U22798 (N_22798,N_17009,N_15071);
nand U22799 (N_22799,N_19423,N_15013);
xnor U22800 (N_22800,N_19329,N_16210);
xor U22801 (N_22801,N_16483,N_15369);
xnor U22802 (N_22802,N_15604,N_17346);
nand U22803 (N_22803,N_18841,N_15579);
or U22804 (N_22804,N_16442,N_18430);
xor U22805 (N_22805,N_16710,N_17565);
and U22806 (N_22806,N_16780,N_17335);
nor U22807 (N_22807,N_15492,N_16749);
nand U22808 (N_22808,N_15237,N_18949);
or U22809 (N_22809,N_19571,N_15486);
xnor U22810 (N_22810,N_16818,N_19363);
or U22811 (N_22811,N_19724,N_19604);
xor U22812 (N_22812,N_16848,N_18593);
xor U22813 (N_22813,N_17899,N_16742);
and U22814 (N_22814,N_18118,N_19184);
and U22815 (N_22815,N_18736,N_15580);
or U22816 (N_22816,N_16546,N_18096);
nor U22817 (N_22817,N_19606,N_17141);
and U22818 (N_22818,N_15372,N_17930);
xor U22819 (N_22819,N_19150,N_15779);
nand U22820 (N_22820,N_17907,N_16978);
nor U22821 (N_22821,N_17017,N_17241);
nor U22822 (N_22822,N_17197,N_17451);
xor U22823 (N_22823,N_18471,N_17076);
or U22824 (N_22824,N_19991,N_16656);
or U22825 (N_22825,N_17861,N_17606);
nand U22826 (N_22826,N_18951,N_16905);
and U22827 (N_22827,N_19561,N_16236);
nor U22828 (N_22828,N_17651,N_18446);
xor U22829 (N_22829,N_15467,N_19393);
xnor U22830 (N_22830,N_17181,N_18091);
or U22831 (N_22831,N_15926,N_19774);
or U22832 (N_22832,N_17057,N_18659);
nor U22833 (N_22833,N_18764,N_17336);
nor U22834 (N_22834,N_18040,N_15147);
nand U22835 (N_22835,N_19220,N_19764);
xnor U22836 (N_22836,N_17223,N_19924);
xnor U22837 (N_22837,N_16840,N_18352);
and U22838 (N_22838,N_17595,N_17875);
xor U22839 (N_22839,N_15296,N_18990);
or U22840 (N_22840,N_15743,N_17216);
or U22841 (N_22841,N_17102,N_19969);
xnor U22842 (N_22842,N_15164,N_19616);
xor U22843 (N_22843,N_17586,N_15924);
nand U22844 (N_22844,N_18302,N_18587);
nor U22845 (N_22845,N_16372,N_15010);
and U22846 (N_22846,N_15739,N_18745);
and U22847 (N_22847,N_16220,N_16768);
and U22848 (N_22848,N_16333,N_18944);
xnor U22849 (N_22849,N_17437,N_17136);
and U22850 (N_22850,N_16781,N_19221);
nor U22851 (N_22851,N_18634,N_19823);
or U22852 (N_22852,N_17756,N_19615);
nand U22853 (N_22853,N_18685,N_19072);
nand U22854 (N_22854,N_16481,N_19777);
nand U22855 (N_22855,N_18901,N_18872);
nor U22856 (N_22856,N_17451,N_19870);
and U22857 (N_22857,N_16909,N_17823);
nand U22858 (N_22858,N_17019,N_18336);
or U22859 (N_22859,N_19271,N_16262);
nand U22860 (N_22860,N_19639,N_16919);
xnor U22861 (N_22861,N_15840,N_19486);
nand U22862 (N_22862,N_18536,N_19247);
nor U22863 (N_22863,N_17494,N_19363);
xnor U22864 (N_22864,N_16294,N_15052);
or U22865 (N_22865,N_15784,N_17117);
or U22866 (N_22866,N_16722,N_18451);
or U22867 (N_22867,N_18980,N_18062);
nand U22868 (N_22868,N_16362,N_15412);
nand U22869 (N_22869,N_17696,N_19584);
and U22870 (N_22870,N_18600,N_15973);
nand U22871 (N_22871,N_18155,N_19603);
xor U22872 (N_22872,N_16048,N_17016);
nand U22873 (N_22873,N_17867,N_15526);
xnor U22874 (N_22874,N_19332,N_16909);
xor U22875 (N_22875,N_19625,N_19532);
or U22876 (N_22876,N_17778,N_17126);
and U22877 (N_22877,N_18648,N_15163);
nor U22878 (N_22878,N_16102,N_16920);
and U22879 (N_22879,N_18884,N_19501);
nor U22880 (N_22880,N_18969,N_16915);
and U22881 (N_22881,N_18299,N_16768);
and U22882 (N_22882,N_18157,N_15775);
xor U22883 (N_22883,N_17252,N_18402);
or U22884 (N_22884,N_17844,N_16076);
or U22885 (N_22885,N_15308,N_17051);
xnor U22886 (N_22886,N_19576,N_19630);
or U22887 (N_22887,N_17058,N_18392);
nor U22888 (N_22888,N_17982,N_19911);
xnor U22889 (N_22889,N_17490,N_19320);
nand U22890 (N_22890,N_16648,N_15450);
or U22891 (N_22891,N_16866,N_17098);
nor U22892 (N_22892,N_17226,N_17032);
nor U22893 (N_22893,N_17406,N_19005);
xnor U22894 (N_22894,N_15654,N_16775);
xor U22895 (N_22895,N_18089,N_19470);
and U22896 (N_22896,N_15433,N_17213);
nand U22897 (N_22897,N_17458,N_17350);
or U22898 (N_22898,N_16940,N_15647);
or U22899 (N_22899,N_16893,N_18280);
xnor U22900 (N_22900,N_17987,N_16668);
or U22901 (N_22901,N_18190,N_19076);
xor U22902 (N_22902,N_19674,N_16280);
xnor U22903 (N_22903,N_15398,N_15389);
xor U22904 (N_22904,N_19801,N_18317);
or U22905 (N_22905,N_17783,N_19988);
or U22906 (N_22906,N_16174,N_18470);
nor U22907 (N_22907,N_18172,N_15374);
or U22908 (N_22908,N_15184,N_19306);
or U22909 (N_22909,N_17581,N_15754);
and U22910 (N_22910,N_18194,N_19736);
and U22911 (N_22911,N_16408,N_18851);
or U22912 (N_22912,N_19933,N_16161);
nor U22913 (N_22913,N_15978,N_15281);
and U22914 (N_22914,N_16506,N_18352);
or U22915 (N_22915,N_15804,N_15363);
xor U22916 (N_22916,N_18711,N_15628);
nor U22917 (N_22917,N_16698,N_15287);
nand U22918 (N_22918,N_15383,N_17267);
or U22919 (N_22919,N_19247,N_18459);
nor U22920 (N_22920,N_15722,N_17846);
xor U22921 (N_22921,N_16574,N_18047);
and U22922 (N_22922,N_16330,N_19337);
or U22923 (N_22923,N_18709,N_16085);
xnor U22924 (N_22924,N_18230,N_16199);
nand U22925 (N_22925,N_16912,N_18840);
or U22926 (N_22926,N_15704,N_19167);
and U22927 (N_22927,N_16821,N_17389);
xor U22928 (N_22928,N_18468,N_18752);
nor U22929 (N_22929,N_18151,N_15470);
xnor U22930 (N_22930,N_17184,N_15223);
xnor U22931 (N_22931,N_15174,N_15762);
and U22932 (N_22932,N_17062,N_17804);
xor U22933 (N_22933,N_18604,N_18651);
nor U22934 (N_22934,N_17356,N_15408);
or U22935 (N_22935,N_18638,N_15930);
and U22936 (N_22936,N_15346,N_16435);
or U22937 (N_22937,N_15282,N_16241);
or U22938 (N_22938,N_17348,N_17061);
xor U22939 (N_22939,N_17206,N_15117);
nor U22940 (N_22940,N_17293,N_15472);
xnor U22941 (N_22941,N_17817,N_19347);
or U22942 (N_22942,N_17184,N_15935);
xnor U22943 (N_22943,N_19880,N_19052);
nor U22944 (N_22944,N_18777,N_16302);
or U22945 (N_22945,N_19786,N_17630);
or U22946 (N_22946,N_15291,N_16873);
or U22947 (N_22947,N_19694,N_19149);
xnor U22948 (N_22948,N_18595,N_19777);
or U22949 (N_22949,N_15960,N_19903);
nand U22950 (N_22950,N_17234,N_15896);
nand U22951 (N_22951,N_16323,N_18861);
or U22952 (N_22952,N_16829,N_16868);
or U22953 (N_22953,N_19103,N_16559);
nor U22954 (N_22954,N_19648,N_16469);
nand U22955 (N_22955,N_15631,N_15218);
xnor U22956 (N_22956,N_17354,N_19606);
xor U22957 (N_22957,N_15836,N_19540);
nand U22958 (N_22958,N_15620,N_16972);
or U22959 (N_22959,N_17452,N_18440);
and U22960 (N_22960,N_19768,N_18842);
xor U22961 (N_22961,N_15454,N_17006);
nand U22962 (N_22962,N_18195,N_17979);
xnor U22963 (N_22963,N_18856,N_19508);
nor U22964 (N_22964,N_18605,N_15136);
xnor U22965 (N_22965,N_16442,N_18528);
nand U22966 (N_22966,N_19508,N_18355);
nor U22967 (N_22967,N_18237,N_17315);
xnor U22968 (N_22968,N_17557,N_17226);
or U22969 (N_22969,N_17222,N_18946);
nor U22970 (N_22970,N_19702,N_17584);
or U22971 (N_22971,N_15308,N_15567);
or U22972 (N_22972,N_15820,N_16188);
nand U22973 (N_22973,N_15323,N_16100);
xor U22974 (N_22974,N_17916,N_15435);
or U22975 (N_22975,N_18724,N_16193);
xnor U22976 (N_22976,N_16645,N_17541);
nand U22977 (N_22977,N_19899,N_19559);
xnor U22978 (N_22978,N_18561,N_16641);
or U22979 (N_22979,N_15490,N_18269);
xor U22980 (N_22980,N_17182,N_19229);
nand U22981 (N_22981,N_18114,N_19910);
xnor U22982 (N_22982,N_19691,N_15010);
xnor U22983 (N_22983,N_16599,N_15237);
xor U22984 (N_22984,N_18229,N_18104);
or U22985 (N_22985,N_15962,N_19601);
xnor U22986 (N_22986,N_17509,N_17309);
or U22987 (N_22987,N_18462,N_17394);
xnor U22988 (N_22988,N_17927,N_17098);
xnor U22989 (N_22989,N_19275,N_18072);
xnor U22990 (N_22990,N_19504,N_18213);
nand U22991 (N_22991,N_16440,N_18717);
nand U22992 (N_22992,N_17307,N_17833);
nand U22993 (N_22993,N_18786,N_16417);
xor U22994 (N_22994,N_17896,N_16096);
nand U22995 (N_22995,N_17803,N_17741);
or U22996 (N_22996,N_15953,N_19953);
or U22997 (N_22997,N_18507,N_15047);
nor U22998 (N_22998,N_19842,N_19484);
and U22999 (N_22999,N_17141,N_19244);
or U23000 (N_23000,N_17914,N_16284);
and U23001 (N_23001,N_16255,N_18065);
or U23002 (N_23002,N_15545,N_19688);
nor U23003 (N_23003,N_15006,N_17955);
nand U23004 (N_23004,N_17073,N_17232);
nor U23005 (N_23005,N_15303,N_15119);
nand U23006 (N_23006,N_18124,N_16788);
nor U23007 (N_23007,N_17037,N_16310);
nand U23008 (N_23008,N_18291,N_18670);
nor U23009 (N_23009,N_18403,N_19081);
or U23010 (N_23010,N_15244,N_19851);
or U23011 (N_23011,N_16071,N_17307);
nor U23012 (N_23012,N_19740,N_19782);
xor U23013 (N_23013,N_19634,N_18723);
or U23014 (N_23014,N_19780,N_15683);
and U23015 (N_23015,N_15720,N_17550);
xnor U23016 (N_23016,N_19931,N_16169);
and U23017 (N_23017,N_17564,N_18354);
nand U23018 (N_23018,N_15891,N_15998);
nor U23019 (N_23019,N_17408,N_18483);
or U23020 (N_23020,N_19094,N_15358);
nand U23021 (N_23021,N_17314,N_19508);
nand U23022 (N_23022,N_17455,N_16261);
xor U23023 (N_23023,N_17794,N_17833);
and U23024 (N_23024,N_17213,N_19150);
or U23025 (N_23025,N_17038,N_17176);
nand U23026 (N_23026,N_15798,N_15411);
or U23027 (N_23027,N_17925,N_18785);
and U23028 (N_23028,N_19275,N_19705);
or U23029 (N_23029,N_16332,N_16146);
xor U23030 (N_23030,N_19036,N_17078);
nand U23031 (N_23031,N_16692,N_18892);
and U23032 (N_23032,N_16433,N_19741);
nor U23033 (N_23033,N_19646,N_17577);
nand U23034 (N_23034,N_16864,N_19588);
or U23035 (N_23035,N_18605,N_15805);
nor U23036 (N_23036,N_19016,N_18197);
xnor U23037 (N_23037,N_17704,N_16992);
and U23038 (N_23038,N_17809,N_18314);
and U23039 (N_23039,N_16591,N_18091);
or U23040 (N_23040,N_19137,N_16529);
nand U23041 (N_23041,N_15378,N_18066);
xnor U23042 (N_23042,N_19056,N_15921);
and U23043 (N_23043,N_17201,N_18759);
nor U23044 (N_23044,N_17943,N_18054);
or U23045 (N_23045,N_18137,N_17278);
nand U23046 (N_23046,N_19817,N_19345);
or U23047 (N_23047,N_18633,N_17267);
and U23048 (N_23048,N_18921,N_18453);
and U23049 (N_23049,N_17070,N_16766);
and U23050 (N_23050,N_16058,N_16578);
and U23051 (N_23051,N_18732,N_16793);
nor U23052 (N_23052,N_15239,N_16363);
or U23053 (N_23053,N_15463,N_15618);
and U23054 (N_23054,N_16698,N_15175);
nand U23055 (N_23055,N_17892,N_18308);
xnor U23056 (N_23056,N_16510,N_19161);
nand U23057 (N_23057,N_19576,N_16286);
and U23058 (N_23058,N_18732,N_18796);
xor U23059 (N_23059,N_18005,N_17514);
xnor U23060 (N_23060,N_19754,N_18871);
or U23061 (N_23061,N_19630,N_16414);
nor U23062 (N_23062,N_16690,N_15431);
and U23063 (N_23063,N_15124,N_16867);
xor U23064 (N_23064,N_18044,N_17577);
and U23065 (N_23065,N_18586,N_17181);
and U23066 (N_23066,N_19818,N_15596);
xnor U23067 (N_23067,N_16708,N_18883);
xnor U23068 (N_23068,N_17905,N_19155);
xnor U23069 (N_23069,N_18654,N_18857);
nor U23070 (N_23070,N_15384,N_15881);
nand U23071 (N_23071,N_15386,N_19490);
xor U23072 (N_23072,N_16265,N_19824);
xor U23073 (N_23073,N_19535,N_16459);
nor U23074 (N_23074,N_18444,N_18737);
xor U23075 (N_23075,N_18397,N_19333);
xor U23076 (N_23076,N_18794,N_17634);
and U23077 (N_23077,N_18799,N_18834);
or U23078 (N_23078,N_16586,N_18022);
and U23079 (N_23079,N_15023,N_17697);
and U23080 (N_23080,N_18946,N_17978);
and U23081 (N_23081,N_18499,N_19308);
nor U23082 (N_23082,N_16108,N_18165);
or U23083 (N_23083,N_16681,N_19197);
nand U23084 (N_23084,N_19695,N_19015);
and U23085 (N_23085,N_18610,N_16221);
and U23086 (N_23086,N_17151,N_17143);
xnor U23087 (N_23087,N_16064,N_17005);
nor U23088 (N_23088,N_18880,N_19548);
nand U23089 (N_23089,N_18854,N_15532);
or U23090 (N_23090,N_18866,N_16995);
xor U23091 (N_23091,N_18844,N_15508);
nand U23092 (N_23092,N_18996,N_16981);
xnor U23093 (N_23093,N_16797,N_17777);
or U23094 (N_23094,N_17022,N_18153);
nor U23095 (N_23095,N_16038,N_15863);
or U23096 (N_23096,N_16203,N_19682);
nand U23097 (N_23097,N_15137,N_16336);
xnor U23098 (N_23098,N_16455,N_19431);
or U23099 (N_23099,N_19073,N_16808);
and U23100 (N_23100,N_19435,N_17464);
xor U23101 (N_23101,N_17456,N_16742);
and U23102 (N_23102,N_19399,N_17241);
and U23103 (N_23103,N_19172,N_18489);
or U23104 (N_23104,N_15255,N_19299);
and U23105 (N_23105,N_18054,N_19549);
nor U23106 (N_23106,N_16709,N_19655);
or U23107 (N_23107,N_18136,N_16587);
and U23108 (N_23108,N_17976,N_15323);
nand U23109 (N_23109,N_18862,N_18845);
and U23110 (N_23110,N_16924,N_17140);
and U23111 (N_23111,N_18329,N_19291);
and U23112 (N_23112,N_18518,N_18212);
nor U23113 (N_23113,N_15417,N_16051);
or U23114 (N_23114,N_17347,N_15504);
nand U23115 (N_23115,N_17487,N_16918);
or U23116 (N_23116,N_16126,N_17409);
or U23117 (N_23117,N_16520,N_15850);
or U23118 (N_23118,N_16517,N_16261);
nand U23119 (N_23119,N_15249,N_19598);
nand U23120 (N_23120,N_19935,N_15343);
nand U23121 (N_23121,N_17464,N_17004);
or U23122 (N_23122,N_17073,N_16110);
xor U23123 (N_23123,N_15570,N_15188);
nand U23124 (N_23124,N_19482,N_16295);
or U23125 (N_23125,N_17918,N_17928);
and U23126 (N_23126,N_15836,N_18649);
nand U23127 (N_23127,N_16087,N_17637);
nor U23128 (N_23128,N_16921,N_18169);
or U23129 (N_23129,N_16917,N_17810);
nand U23130 (N_23130,N_15603,N_17700);
nand U23131 (N_23131,N_18725,N_15171);
and U23132 (N_23132,N_16979,N_19130);
nand U23133 (N_23133,N_19532,N_19529);
or U23134 (N_23134,N_19091,N_15173);
or U23135 (N_23135,N_16316,N_19875);
nor U23136 (N_23136,N_16342,N_19812);
and U23137 (N_23137,N_16448,N_19858);
xnor U23138 (N_23138,N_19197,N_16438);
nand U23139 (N_23139,N_16863,N_16309);
and U23140 (N_23140,N_17791,N_17272);
xor U23141 (N_23141,N_19315,N_18378);
nand U23142 (N_23142,N_17411,N_18347);
nor U23143 (N_23143,N_16598,N_18624);
and U23144 (N_23144,N_17765,N_18109);
xor U23145 (N_23145,N_18803,N_19354);
or U23146 (N_23146,N_18715,N_18747);
or U23147 (N_23147,N_15115,N_18069);
nand U23148 (N_23148,N_19921,N_15224);
nand U23149 (N_23149,N_15326,N_17926);
or U23150 (N_23150,N_16120,N_18713);
nor U23151 (N_23151,N_15715,N_18731);
nor U23152 (N_23152,N_19546,N_17634);
or U23153 (N_23153,N_18974,N_17737);
and U23154 (N_23154,N_15568,N_18554);
and U23155 (N_23155,N_18710,N_15038);
nor U23156 (N_23156,N_19930,N_18979);
and U23157 (N_23157,N_16656,N_19999);
xor U23158 (N_23158,N_15885,N_15975);
nor U23159 (N_23159,N_15306,N_18342);
or U23160 (N_23160,N_19921,N_18430);
nor U23161 (N_23161,N_16636,N_17030);
or U23162 (N_23162,N_16162,N_17964);
nand U23163 (N_23163,N_19881,N_19540);
and U23164 (N_23164,N_19005,N_17277);
or U23165 (N_23165,N_19208,N_15319);
and U23166 (N_23166,N_19561,N_18735);
nand U23167 (N_23167,N_16024,N_17571);
nand U23168 (N_23168,N_16627,N_15158);
or U23169 (N_23169,N_15326,N_16019);
xnor U23170 (N_23170,N_17136,N_18353);
xor U23171 (N_23171,N_18846,N_15584);
xnor U23172 (N_23172,N_16723,N_16551);
nand U23173 (N_23173,N_15211,N_17633);
or U23174 (N_23174,N_17675,N_18149);
nor U23175 (N_23175,N_17291,N_18760);
xnor U23176 (N_23176,N_18027,N_18442);
xor U23177 (N_23177,N_17313,N_16162);
nand U23178 (N_23178,N_15100,N_19174);
nor U23179 (N_23179,N_15737,N_18202);
nor U23180 (N_23180,N_15676,N_16466);
or U23181 (N_23181,N_15821,N_16312);
or U23182 (N_23182,N_17274,N_18934);
xnor U23183 (N_23183,N_15626,N_16769);
nand U23184 (N_23184,N_15692,N_19865);
xor U23185 (N_23185,N_18555,N_15673);
xor U23186 (N_23186,N_17036,N_19113);
and U23187 (N_23187,N_16957,N_18578);
nand U23188 (N_23188,N_18466,N_18536);
and U23189 (N_23189,N_17696,N_16538);
or U23190 (N_23190,N_17402,N_18985);
xor U23191 (N_23191,N_16636,N_19195);
or U23192 (N_23192,N_17813,N_18800);
nand U23193 (N_23193,N_17804,N_18832);
or U23194 (N_23194,N_15906,N_15661);
and U23195 (N_23195,N_18293,N_15738);
and U23196 (N_23196,N_18062,N_15557);
xnor U23197 (N_23197,N_17907,N_19338);
nor U23198 (N_23198,N_19893,N_16563);
nor U23199 (N_23199,N_17377,N_16731);
or U23200 (N_23200,N_19933,N_19040);
nor U23201 (N_23201,N_19492,N_17518);
nor U23202 (N_23202,N_16409,N_15171);
and U23203 (N_23203,N_15052,N_15209);
xnor U23204 (N_23204,N_17523,N_16491);
nor U23205 (N_23205,N_18667,N_15659);
xor U23206 (N_23206,N_19774,N_18231);
or U23207 (N_23207,N_18929,N_17009);
or U23208 (N_23208,N_18263,N_19588);
or U23209 (N_23209,N_18965,N_15235);
xor U23210 (N_23210,N_17220,N_17490);
and U23211 (N_23211,N_17696,N_18377);
nor U23212 (N_23212,N_19977,N_16800);
nand U23213 (N_23213,N_16680,N_16052);
or U23214 (N_23214,N_15528,N_17109);
xor U23215 (N_23215,N_17792,N_17767);
or U23216 (N_23216,N_16043,N_19913);
nor U23217 (N_23217,N_19073,N_18879);
xnor U23218 (N_23218,N_19304,N_19126);
nand U23219 (N_23219,N_17516,N_15125);
or U23220 (N_23220,N_17602,N_17495);
nand U23221 (N_23221,N_18086,N_19024);
and U23222 (N_23222,N_16774,N_18955);
xor U23223 (N_23223,N_17728,N_19298);
and U23224 (N_23224,N_15870,N_17553);
nand U23225 (N_23225,N_18973,N_16125);
nand U23226 (N_23226,N_19089,N_17119);
and U23227 (N_23227,N_16254,N_17007);
and U23228 (N_23228,N_17769,N_18395);
and U23229 (N_23229,N_16688,N_17616);
and U23230 (N_23230,N_17399,N_18697);
xor U23231 (N_23231,N_17248,N_16919);
and U23232 (N_23232,N_17129,N_17996);
nor U23233 (N_23233,N_18484,N_19305);
nor U23234 (N_23234,N_16061,N_17302);
or U23235 (N_23235,N_15161,N_17141);
nand U23236 (N_23236,N_17950,N_15629);
xor U23237 (N_23237,N_17238,N_17577);
and U23238 (N_23238,N_15983,N_15855);
nor U23239 (N_23239,N_19104,N_17170);
xnor U23240 (N_23240,N_16985,N_16277);
or U23241 (N_23241,N_19645,N_18172);
or U23242 (N_23242,N_15396,N_19278);
nor U23243 (N_23243,N_16649,N_19920);
nand U23244 (N_23244,N_15532,N_15806);
or U23245 (N_23245,N_15454,N_18879);
nor U23246 (N_23246,N_15190,N_15262);
and U23247 (N_23247,N_15729,N_19274);
or U23248 (N_23248,N_16661,N_16289);
nand U23249 (N_23249,N_19238,N_18346);
or U23250 (N_23250,N_15106,N_15937);
or U23251 (N_23251,N_19563,N_17092);
or U23252 (N_23252,N_17134,N_15293);
or U23253 (N_23253,N_18803,N_15757);
xor U23254 (N_23254,N_19408,N_18114);
and U23255 (N_23255,N_19078,N_16859);
nor U23256 (N_23256,N_15134,N_17270);
nor U23257 (N_23257,N_16999,N_15543);
or U23258 (N_23258,N_16730,N_18609);
and U23259 (N_23259,N_19745,N_16763);
and U23260 (N_23260,N_19150,N_15399);
nor U23261 (N_23261,N_17226,N_16448);
and U23262 (N_23262,N_17296,N_19108);
or U23263 (N_23263,N_17333,N_18306);
or U23264 (N_23264,N_17649,N_18120);
nand U23265 (N_23265,N_18849,N_17203);
nand U23266 (N_23266,N_15684,N_19769);
and U23267 (N_23267,N_19390,N_16484);
or U23268 (N_23268,N_18399,N_19469);
and U23269 (N_23269,N_19773,N_18147);
or U23270 (N_23270,N_17330,N_16469);
nand U23271 (N_23271,N_19488,N_19412);
or U23272 (N_23272,N_15876,N_19077);
nand U23273 (N_23273,N_18638,N_16310);
and U23274 (N_23274,N_17163,N_17588);
and U23275 (N_23275,N_18562,N_15770);
nor U23276 (N_23276,N_17881,N_16121);
nor U23277 (N_23277,N_17899,N_17856);
xnor U23278 (N_23278,N_16892,N_16575);
and U23279 (N_23279,N_16875,N_15446);
nor U23280 (N_23280,N_19879,N_15332);
or U23281 (N_23281,N_18647,N_17935);
and U23282 (N_23282,N_15221,N_16848);
and U23283 (N_23283,N_16940,N_15094);
nor U23284 (N_23284,N_19435,N_17407);
xor U23285 (N_23285,N_16658,N_18342);
or U23286 (N_23286,N_18738,N_18432);
nand U23287 (N_23287,N_15342,N_19440);
and U23288 (N_23288,N_19162,N_16673);
nand U23289 (N_23289,N_16046,N_19045);
xor U23290 (N_23290,N_18063,N_18175);
nand U23291 (N_23291,N_19403,N_19528);
and U23292 (N_23292,N_17742,N_15726);
or U23293 (N_23293,N_18010,N_15027);
or U23294 (N_23294,N_17223,N_19935);
xor U23295 (N_23295,N_17302,N_19734);
xor U23296 (N_23296,N_15612,N_17260);
xor U23297 (N_23297,N_17291,N_15638);
or U23298 (N_23298,N_15990,N_16843);
or U23299 (N_23299,N_19673,N_17180);
and U23300 (N_23300,N_18245,N_16287);
and U23301 (N_23301,N_17310,N_16132);
and U23302 (N_23302,N_19804,N_19575);
nor U23303 (N_23303,N_16990,N_19965);
nand U23304 (N_23304,N_18557,N_19170);
xnor U23305 (N_23305,N_15962,N_15129);
and U23306 (N_23306,N_17976,N_16907);
xnor U23307 (N_23307,N_17046,N_15347);
nand U23308 (N_23308,N_17051,N_17330);
nor U23309 (N_23309,N_16090,N_16483);
or U23310 (N_23310,N_16697,N_19340);
nand U23311 (N_23311,N_16664,N_15180);
nor U23312 (N_23312,N_15393,N_17622);
nand U23313 (N_23313,N_15936,N_15410);
and U23314 (N_23314,N_19548,N_19805);
and U23315 (N_23315,N_19086,N_18420);
nor U23316 (N_23316,N_15979,N_19182);
or U23317 (N_23317,N_15647,N_18057);
nand U23318 (N_23318,N_17177,N_17849);
xor U23319 (N_23319,N_17254,N_16938);
xor U23320 (N_23320,N_19943,N_17120);
nand U23321 (N_23321,N_16950,N_17319);
and U23322 (N_23322,N_17717,N_17089);
or U23323 (N_23323,N_15920,N_15672);
nand U23324 (N_23324,N_16652,N_18121);
and U23325 (N_23325,N_17113,N_18018);
and U23326 (N_23326,N_18314,N_17473);
xnor U23327 (N_23327,N_19815,N_16622);
nor U23328 (N_23328,N_16215,N_17734);
nand U23329 (N_23329,N_17974,N_17164);
xnor U23330 (N_23330,N_16438,N_15886);
nor U23331 (N_23331,N_15432,N_16541);
or U23332 (N_23332,N_17040,N_16784);
and U23333 (N_23333,N_15486,N_18035);
nand U23334 (N_23334,N_19353,N_15174);
nand U23335 (N_23335,N_18757,N_17148);
or U23336 (N_23336,N_19748,N_18793);
xor U23337 (N_23337,N_18974,N_19078);
or U23338 (N_23338,N_19449,N_16331);
xnor U23339 (N_23339,N_16452,N_19332);
nor U23340 (N_23340,N_16123,N_18268);
xor U23341 (N_23341,N_19966,N_19033);
xnor U23342 (N_23342,N_16438,N_15321);
or U23343 (N_23343,N_18207,N_17894);
and U23344 (N_23344,N_17853,N_15643);
xnor U23345 (N_23345,N_18705,N_17478);
xor U23346 (N_23346,N_19627,N_17420);
or U23347 (N_23347,N_17486,N_17126);
or U23348 (N_23348,N_15189,N_16702);
and U23349 (N_23349,N_16347,N_17691);
nand U23350 (N_23350,N_19909,N_16325);
and U23351 (N_23351,N_15726,N_15460);
nand U23352 (N_23352,N_16995,N_18027);
xor U23353 (N_23353,N_17718,N_17679);
and U23354 (N_23354,N_18650,N_19428);
nand U23355 (N_23355,N_19795,N_17296);
or U23356 (N_23356,N_17610,N_19728);
or U23357 (N_23357,N_15394,N_19281);
or U23358 (N_23358,N_19737,N_17749);
xor U23359 (N_23359,N_19322,N_19155);
nor U23360 (N_23360,N_15001,N_16229);
and U23361 (N_23361,N_17500,N_19681);
nand U23362 (N_23362,N_19633,N_16489);
or U23363 (N_23363,N_16931,N_19920);
or U23364 (N_23364,N_19180,N_19181);
nor U23365 (N_23365,N_15966,N_16717);
xor U23366 (N_23366,N_18103,N_19637);
nand U23367 (N_23367,N_19243,N_18498);
nand U23368 (N_23368,N_19056,N_19053);
nor U23369 (N_23369,N_15704,N_18662);
nor U23370 (N_23370,N_19687,N_16798);
nor U23371 (N_23371,N_18538,N_19632);
xor U23372 (N_23372,N_15646,N_16161);
xor U23373 (N_23373,N_19265,N_19239);
nand U23374 (N_23374,N_18982,N_19967);
or U23375 (N_23375,N_16896,N_15259);
nor U23376 (N_23376,N_18204,N_15980);
xor U23377 (N_23377,N_15533,N_17434);
nor U23378 (N_23378,N_15094,N_15767);
nand U23379 (N_23379,N_16699,N_19252);
and U23380 (N_23380,N_16758,N_19242);
and U23381 (N_23381,N_18337,N_18328);
and U23382 (N_23382,N_16287,N_15300);
nand U23383 (N_23383,N_18136,N_17765);
nand U23384 (N_23384,N_15294,N_17992);
and U23385 (N_23385,N_18050,N_19466);
or U23386 (N_23386,N_18173,N_17141);
or U23387 (N_23387,N_19142,N_17702);
and U23388 (N_23388,N_15987,N_16377);
nand U23389 (N_23389,N_19138,N_18809);
xnor U23390 (N_23390,N_17109,N_19629);
nor U23391 (N_23391,N_18387,N_18395);
xnor U23392 (N_23392,N_15042,N_18665);
and U23393 (N_23393,N_15920,N_19486);
and U23394 (N_23394,N_18581,N_18925);
or U23395 (N_23395,N_19019,N_15808);
or U23396 (N_23396,N_19649,N_19044);
and U23397 (N_23397,N_17100,N_15974);
or U23398 (N_23398,N_17106,N_16935);
xor U23399 (N_23399,N_19139,N_15084);
nor U23400 (N_23400,N_15149,N_17910);
or U23401 (N_23401,N_18454,N_17836);
nor U23402 (N_23402,N_16916,N_19696);
nor U23403 (N_23403,N_17537,N_18235);
nor U23404 (N_23404,N_19998,N_15160);
nand U23405 (N_23405,N_16531,N_15110);
or U23406 (N_23406,N_17791,N_18448);
nand U23407 (N_23407,N_16581,N_18749);
or U23408 (N_23408,N_15900,N_15522);
nor U23409 (N_23409,N_17942,N_19877);
nor U23410 (N_23410,N_16824,N_19307);
and U23411 (N_23411,N_18232,N_19832);
or U23412 (N_23412,N_16462,N_17263);
nor U23413 (N_23413,N_16066,N_15782);
or U23414 (N_23414,N_18142,N_17628);
nand U23415 (N_23415,N_19256,N_15457);
xor U23416 (N_23416,N_19311,N_19654);
nand U23417 (N_23417,N_15895,N_18767);
xor U23418 (N_23418,N_16957,N_15707);
and U23419 (N_23419,N_19555,N_15765);
and U23420 (N_23420,N_19882,N_15456);
or U23421 (N_23421,N_16885,N_18930);
nand U23422 (N_23422,N_17230,N_17482);
xor U23423 (N_23423,N_17600,N_18596);
xnor U23424 (N_23424,N_16512,N_16788);
or U23425 (N_23425,N_15595,N_17584);
nand U23426 (N_23426,N_15005,N_17730);
nor U23427 (N_23427,N_18534,N_19381);
or U23428 (N_23428,N_19315,N_18672);
and U23429 (N_23429,N_15638,N_18574);
and U23430 (N_23430,N_19676,N_15790);
and U23431 (N_23431,N_17591,N_15515);
nor U23432 (N_23432,N_15167,N_15097);
xor U23433 (N_23433,N_18508,N_15544);
nand U23434 (N_23434,N_15079,N_17662);
and U23435 (N_23435,N_16789,N_17995);
or U23436 (N_23436,N_17035,N_18626);
or U23437 (N_23437,N_16796,N_16734);
xor U23438 (N_23438,N_18616,N_15348);
nand U23439 (N_23439,N_19283,N_19863);
and U23440 (N_23440,N_16057,N_19097);
nor U23441 (N_23441,N_16942,N_19032);
nand U23442 (N_23442,N_17029,N_16626);
nand U23443 (N_23443,N_16835,N_19008);
xor U23444 (N_23444,N_15696,N_17633);
and U23445 (N_23445,N_18150,N_16350);
and U23446 (N_23446,N_18101,N_19231);
and U23447 (N_23447,N_16626,N_18738);
xnor U23448 (N_23448,N_16561,N_18581);
nand U23449 (N_23449,N_15645,N_17460);
nor U23450 (N_23450,N_19654,N_15299);
xor U23451 (N_23451,N_19886,N_15963);
and U23452 (N_23452,N_17153,N_19271);
xor U23453 (N_23453,N_18238,N_18277);
nand U23454 (N_23454,N_17949,N_18394);
xnor U23455 (N_23455,N_15638,N_19088);
or U23456 (N_23456,N_15266,N_15769);
xnor U23457 (N_23457,N_16115,N_17598);
nand U23458 (N_23458,N_16592,N_17504);
or U23459 (N_23459,N_16070,N_18609);
nand U23460 (N_23460,N_15445,N_16393);
nor U23461 (N_23461,N_19210,N_15258);
xnor U23462 (N_23462,N_18059,N_17610);
nor U23463 (N_23463,N_19567,N_19021);
and U23464 (N_23464,N_18027,N_15946);
nand U23465 (N_23465,N_16669,N_19256);
nor U23466 (N_23466,N_18308,N_15427);
nand U23467 (N_23467,N_18880,N_15779);
nand U23468 (N_23468,N_17443,N_17009);
nor U23469 (N_23469,N_15036,N_19669);
nor U23470 (N_23470,N_16269,N_18375);
nor U23471 (N_23471,N_15971,N_18449);
nand U23472 (N_23472,N_15634,N_15954);
xor U23473 (N_23473,N_16510,N_16334);
or U23474 (N_23474,N_15346,N_15155);
nand U23475 (N_23475,N_16585,N_17916);
nand U23476 (N_23476,N_19785,N_15519);
or U23477 (N_23477,N_18123,N_19951);
and U23478 (N_23478,N_19877,N_15170);
or U23479 (N_23479,N_15731,N_17271);
nand U23480 (N_23480,N_16781,N_19929);
xnor U23481 (N_23481,N_15876,N_18207);
nor U23482 (N_23482,N_19737,N_17014);
nor U23483 (N_23483,N_15477,N_19328);
and U23484 (N_23484,N_18846,N_17372);
nor U23485 (N_23485,N_18958,N_15903);
or U23486 (N_23486,N_19767,N_17908);
nand U23487 (N_23487,N_18570,N_18103);
nor U23488 (N_23488,N_16431,N_19439);
or U23489 (N_23489,N_16549,N_17752);
nor U23490 (N_23490,N_15023,N_18908);
nand U23491 (N_23491,N_19581,N_18255);
nor U23492 (N_23492,N_19154,N_16645);
or U23493 (N_23493,N_18629,N_16897);
or U23494 (N_23494,N_15521,N_15657);
xnor U23495 (N_23495,N_19248,N_17698);
nor U23496 (N_23496,N_16868,N_19456);
xnor U23497 (N_23497,N_19152,N_15928);
or U23498 (N_23498,N_19075,N_19394);
or U23499 (N_23499,N_17979,N_19937);
nand U23500 (N_23500,N_18868,N_18369);
nand U23501 (N_23501,N_18838,N_19767);
and U23502 (N_23502,N_18176,N_16389);
and U23503 (N_23503,N_19674,N_19408);
and U23504 (N_23504,N_18468,N_16734);
xor U23505 (N_23505,N_18545,N_17671);
nor U23506 (N_23506,N_18060,N_17935);
nor U23507 (N_23507,N_16390,N_17860);
and U23508 (N_23508,N_18666,N_17352);
and U23509 (N_23509,N_15195,N_18292);
or U23510 (N_23510,N_15730,N_19103);
and U23511 (N_23511,N_17160,N_17791);
nand U23512 (N_23512,N_17727,N_17363);
nand U23513 (N_23513,N_15131,N_16679);
xor U23514 (N_23514,N_18189,N_17481);
or U23515 (N_23515,N_18920,N_17530);
nor U23516 (N_23516,N_18711,N_18425);
nand U23517 (N_23517,N_18788,N_19530);
xor U23518 (N_23518,N_19166,N_17538);
nand U23519 (N_23519,N_18719,N_19434);
xnor U23520 (N_23520,N_18370,N_18350);
or U23521 (N_23521,N_18203,N_17660);
and U23522 (N_23522,N_15179,N_16692);
nor U23523 (N_23523,N_15006,N_17618);
nor U23524 (N_23524,N_17963,N_18466);
nand U23525 (N_23525,N_18677,N_17094);
xor U23526 (N_23526,N_16103,N_17525);
and U23527 (N_23527,N_16381,N_15424);
and U23528 (N_23528,N_19964,N_15794);
or U23529 (N_23529,N_15660,N_15401);
and U23530 (N_23530,N_16103,N_15669);
nand U23531 (N_23531,N_15640,N_17326);
xnor U23532 (N_23532,N_16425,N_15902);
nor U23533 (N_23533,N_18639,N_15376);
or U23534 (N_23534,N_19236,N_17039);
or U23535 (N_23535,N_17825,N_19547);
xnor U23536 (N_23536,N_16666,N_19407);
nand U23537 (N_23537,N_18929,N_19395);
and U23538 (N_23538,N_15374,N_17689);
or U23539 (N_23539,N_15657,N_17930);
and U23540 (N_23540,N_16020,N_16373);
nor U23541 (N_23541,N_17323,N_18718);
and U23542 (N_23542,N_15792,N_17743);
nor U23543 (N_23543,N_16831,N_16569);
nor U23544 (N_23544,N_15064,N_19355);
or U23545 (N_23545,N_16211,N_16601);
nor U23546 (N_23546,N_19495,N_16044);
nand U23547 (N_23547,N_19807,N_19132);
and U23548 (N_23548,N_18025,N_15408);
or U23549 (N_23549,N_17446,N_18672);
xor U23550 (N_23550,N_17371,N_18397);
and U23551 (N_23551,N_19842,N_17396);
nand U23552 (N_23552,N_15768,N_17901);
xor U23553 (N_23553,N_18332,N_16498);
nand U23554 (N_23554,N_19767,N_15948);
xnor U23555 (N_23555,N_17423,N_19852);
and U23556 (N_23556,N_19830,N_17665);
nand U23557 (N_23557,N_15940,N_15924);
and U23558 (N_23558,N_15355,N_19076);
xor U23559 (N_23559,N_18663,N_18259);
or U23560 (N_23560,N_18731,N_17029);
or U23561 (N_23561,N_15900,N_15848);
nor U23562 (N_23562,N_16489,N_17706);
and U23563 (N_23563,N_17519,N_17103);
nor U23564 (N_23564,N_16299,N_16234);
and U23565 (N_23565,N_16062,N_16592);
or U23566 (N_23566,N_19022,N_19193);
and U23567 (N_23567,N_18735,N_15160);
and U23568 (N_23568,N_15922,N_18920);
xor U23569 (N_23569,N_17998,N_15252);
nand U23570 (N_23570,N_17436,N_16661);
nor U23571 (N_23571,N_19255,N_18295);
xnor U23572 (N_23572,N_15039,N_17677);
nor U23573 (N_23573,N_15158,N_18363);
or U23574 (N_23574,N_19179,N_17804);
xor U23575 (N_23575,N_19861,N_17488);
or U23576 (N_23576,N_19067,N_18285);
xor U23577 (N_23577,N_17040,N_19645);
xnor U23578 (N_23578,N_19909,N_19877);
xor U23579 (N_23579,N_16968,N_16412);
and U23580 (N_23580,N_15439,N_15616);
nor U23581 (N_23581,N_17000,N_16570);
nand U23582 (N_23582,N_16622,N_16822);
and U23583 (N_23583,N_15399,N_19745);
and U23584 (N_23584,N_19693,N_19889);
nand U23585 (N_23585,N_19770,N_18658);
xnor U23586 (N_23586,N_16632,N_15266);
nand U23587 (N_23587,N_18915,N_16270);
nor U23588 (N_23588,N_15624,N_17584);
nand U23589 (N_23589,N_18772,N_17176);
nor U23590 (N_23590,N_17069,N_18477);
nand U23591 (N_23591,N_17321,N_17154);
xnor U23592 (N_23592,N_15095,N_18326);
nand U23593 (N_23593,N_16252,N_15994);
nand U23594 (N_23594,N_15588,N_19190);
and U23595 (N_23595,N_17589,N_18366);
nand U23596 (N_23596,N_19764,N_19887);
or U23597 (N_23597,N_18524,N_17003);
and U23598 (N_23598,N_17958,N_15185);
nand U23599 (N_23599,N_18162,N_19189);
nor U23600 (N_23600,N_19902,N_19275);
nand U23601 (N_23601,N_16509,N_18922);
nor U23602 (N_23602,N_18426,N_17070);
xnor U23603 (N_23603,N_16627,N_17140);
or U23604 (N_23604,N_16904,N_17255);
or U23605 (N_23605,N_15870,N_17081);
or U23606 (N_23606,N_17957,N_19510);
nor U23607 (N_23607,N_17934,N_17593);
nor U23608 (N_23608,N_19515,N_15129);
nand U23609 (N_23609,N_18182,N_17775);
nor U23610 (N_23610,N_18211,N_16717);
and U23611 (N_23611,N_15753,N_19250);
and U23612 (N_23612,N_17775,N_19720);
or U23613 (N_23613,N_16201,N_15352);
and U23614 (N_23614,N_19113,N_19383);
and U23615 (N_23615,N_17728,N_19210);
xor U23616 (N_23616,N_19337,N_17456);
and U23617 (N_23617,N_17727,N_17206);
nand U23618 (N_23618,N_17142,N_18313);
nand U23619 (N_23619,N_16003,N_17293);
nor U23620 (N_23620,N_17146,N_19590);
nand U23621 (N_23621,N_19983,N_17755);
nand U23622 (N_23622,N_16592,N_18542);
or U23623 (N_23623,N_17140,N_17758);
xnor U23624 (N_23624,N_15488,N_15739);
xor U23625 (N_23625,N_17194,N_15977);
and U23626 (N_23626,N_16094,N_16371);
nand U23627 (N_23627,N_18436,N_18610);
and U23628 (N_23628,N_19348,N_18054);
and U23629 (N_23629,N_15971,N_19528);
nand U23630 (N_23630,N_19900,N_16021);
nand U23631 (N_23631,N_18807,N_16626);
xnor U23632 (N_23632,N_17918,N_17739);
or U23633 (N_23633,N_18050,N_15145);
and U23634 (N_23634,N_15945,N_17550);
nor U23635 (N_23635,N_15316,N_17859);
nor U23636 (N_23636,N_17451,N_16214);
and U23637 (N_23637,N_16399,N_19089);
or U23638 (N_23638,N_19044,N_15779);
nor U23639 (N_23639,N_17602,N_18608);
and U23640 (N_23640,N_19179,N_16881);
and U23641 (N_23641,N_19920,N_18149);
or U23642 (N_23642,N_19605,N_15420);
xnor U23643 (N_23643,N_18596,N_15866);
or U23644 (N_23644,N_16380,N_16975);
and U23645 (N_23645,N_19588,N_16171);
nor U23646 (N_23646,N_17182,N_16239);
and U23647 (N_23647,N_16991,N_16023);
and U23648 (N_23648,N_19195,N_15514);
nor U23649 (N_23649,N_19527,N_17602);
and U23650 (N_23650,N_17736,N_19542);
or U23651 (N_23651,N_16278,N_15760);
nand U23652 (N_23652,N_16974,N_18840);
and U23653 (N_23653,N_15287,N_18478);
nand U23654 (N_23654,N_16828,N_17246);
or U23655 (N_23655,N_15295,N_17736);
xnor U23656 (N_23656,N_15557,N_18272);
nor U23657 (N_23657,N_16390,N_18566);
xor U23658 (N_23658,N_19771,N_17462);
nor U23659 (N_23659,N_19394,N_19220);
nor U23660 (N_23660,N_15394,N_19082);
and U23661 (N_23661,N_17953,N_18135);
or U23662 (N_23662,N_16919,N_17680);
nor U23663 (N_23663,N_18309,N_15509);
nor U23664 (N_23664,N_17603,N_19787);
nor U23665 (N_23665,N_17314,N_18373);
xnor U23666 (N_23666,N_16261,N_17609);
and U23667 (N_23667,N_15758,N_18486);
or U23668 (N_23668,N_19853,N_18682);
xor U23669 (N_23669,N_15972,N_18284);
and U23670 (N_23670,N_18615,N_16810);
xor U23671 (N_23671,N_19357,N_15946);
nor U23672 (N_23672,N_19121,N_16415);
nand U23673 (N_23673,N_18281,N_15904);
and U23674 (N_23674,N_17430,N_16043);
nand U23675 (N_23675,N_19278,N_18281);
xnor U23676 (N_23676,N_18997,N_19757);
and U23677 (N_23677,N_19775,N_18223);
nor U23678 (N_23678,N_19898,N_15897);
xor U23679 (N_23679,N_19781,N_16544);
nor U23680 (N_23680,N_15448,N_15872);
nor U23681 (N_23681,N_19770,N_19973);
and U23682 (N_23682,N_16845,N_15561);
xnor U23683 (N_23683,N_15865,N_15448);
nand U23684 (N_23684,N_19516,N_15952);
nand U23685 (N_23685,N_18843,N_17975);
xor U23686 (N_23686,N_18006,N_18402);
xnor U23687 (N_23687,N_19732,N_17979);
nor U23688 (N_23688,N_17351,N_15943);
nor U23689 (N_23689,N_16592,N_15754);
nor U23690 (N_23690,N_15117,N_15197);
and U23691 (N_23691,N_15917,N_16827);
or U23692 (N_23692,N_15611,N_19927);
nor U23693 (N_23693,N_18689,N_15791);
and U23694 (N_23694,N_15956,N_16342);
xor U23695 (N_23695,N_15199,N_19872);
nor U23696 (N_23696,N_17930,N_19780);
nor U23697 (N_23697,N_17896,N_15647);
xnor U23698 (N_23698,N_17720,N_16564);
xnor U23699 (N_23699,N_18911,N_15454);
nand U23700 (N_23700,N_16889,N_15459);
xor U23701 (N_23701,N_16456,N_15973);
nor U23702 (N_23702,N_16011,N_19738);
nand U23703 (N_23703,N_15937,N_16348);
nand U23704 (N_23704,N_16785,N_17215);
nor U23705 (N_23705,N_18097,N_19525);
xor U23706 (N_23706,N_16871,N_18127);
nor U23707 (N_23707,N_15992,N_17799);
nor U23708 (N_23708,N_18541,N_18011);
nand U23709 (N_23709,N_15058,N_19882);
or U23710 (N_23710,N_17477,N_17405);
and U23711 (N_23711,N_15453,N_15368);
nor U23712 (N_23712,N_18136,N_18449);
nor U23713 (N_23713,N_16472,N_16526);
or U23714 (N_23714,N_19488,N_19360);
nor U23715 (N_23715,N_16454,N_15982);
nor U23716 (N_23716,N_15631,N_19625);
or U23717 (N_23717,N_19797,N_16036);
or U23718 (N_23718,N_19966,N_17305);
and U23719 (N_23719,N_19048,N_19034);
nand U23720 (N_23720,N_18619,N_18282);
and U23721 (N_23721,N_19155,N_16728);
and U23722 (N_23722,N_17552,N_17951);
nand U23723 (N_23723,N_16017,N_15282);
nand U23724 (N_23724,N_19605,N_17036);
xnor U23725 (N_23725,N_18073,N_19053);
xor U23726 (N_23726,N_15632,N_19127);
xor U23727 (N_23727,N_17182,N_18220);
and U23728 (N_23728,N_16249,N_18645);
nor U23729 (N_23729,N_17485,N_15019);
or U23730 (N_23730,N_18414,N_15434);
or U23731 (N_23731,N_15582,N_16381);
and U23732 (N_23732,N_17949,N_15172);
and U23733 (N_23733,N_15133,N_16446);
nor U23734 (N_23734,N_19216,N_19115);
nor U23735 (N_23735,N_19181,N_17297);
nand U23736 (N_23736,N_17938,N_17780);
xor U23737 (N_23737,N_18508,N_19196);
xnor U23738 (N_23738,N_17417,N_18708);
nor U23739 (N_23739,N_19856,N_17014);
nand U23740 (N_23740,N_16788,N_17691);
nor U23741 (N_23741,N_16657,N_16767);
and U23742 (N_23742,N_19398,N_15131);
or U23743 (N_23743,N_16433,N_18381);
xnor U23744 (N_23744,N_15358,N_17857);
and U23745 (N_23745,N_16159,N_16199);
xnor U23746 (N_23746,N_18351,N_18243);
nand U23747 (N_23747,N_17172,N_17208);
or U23748 (N_23748,N_18445,N_18774);
or U23749 (N_23749,N_17401,N_17470);
nor U23750 (N_23750,N_15859,N_18685);
nor U23751 (N_23751,N_17578,N_15294);
nor U23752 (N_23752,N_16360,N_17524);
nand U23753 (N_23753,N_18751,N_17661);
nor U23754 (N_23754,N_15302,N_16787);
xnor U23755 (N_23755,N_17915,N_19524);
nor U23756 (N_23756,N_17359,N_18703);
and U23757 (N_23757,N_16745,N_17399);
xnor U23758 (N_23758,N_17230,N_18508);
xnor U23759 (N_23759,N_15811,N_19623);
xnor U23760 (N_23760,N_19477,N_15346);
nand U23761 (N_23761,N_18553,N_17865);
xnor U23762 (N_23762,N_19232,N_16060);
and U23763 (N_23763,N_19299,N_15497);
or U23764 (N_23764,N_16966,N_19198);
nor U23765 (N_23765,N_17745,N_19226);
nand U23766 (N_23766,N_15629,N_19767);
xnor U23767 (N_23767,N_17013,N_16049);
nand U23768 (N_23768,N_18140,N_15867);
nor U23769 (N_23769,N_18996,N_16676);
xor U23770 (N_23770,N_17932,N_19163);
or U23771 (N_23771,N_16265,N_19003);
and U23772 (N_23772,N_15938,N_15271);
nor U23773 (N_23773,N_16648,N_18125);
xor U23774 (N_23774,N_18450,N_16028);
and U23775 (N_23775,N_16635,N_18288);
and U23776 (N_23776,N_17358,N_19058);
xor U23777 (N_23777,N_17935,N_18216);
or U23778 (N_23778,N_17100,N_17217);
nand U23779 (N_23779,N_18361,N_15104);
nand U23780 (N_23780,N_16702,N_16609);
xor U23781 (N_23781,N_17038,N_18551);
or U23782 (N_23782,N_19173,N_17447);
nand U23783 (N_23783,N_19467,N_16796);
nor U23784 (N_23784,N_15562,N_19271);
xor U23785 (N_23785,N_18945,N_19404);
and U23786 (N_23786,N_15812,N_18163);
or U23787 (N_23787,N_15014,N_18964);
nor U23788 (N_23788,N_17603,N_16864);
or U23789 (N_23789,N_19599,N_19789);
or U23790 (N_23790,N_18258,N_18741);
and U23791 (N_23791,N_17093,N_15201);
nand U23792 (N_23792,N_16804,N_15511);
or U23793 (N_23793,N_15011,N_19226);
and U23794 (N_23794,N_17441,N_16170);
or U23795 (N_23795,N_18694,N_15473);
xnor U23796 (N_23796,N_16978,N_18377);
nand U23797 (N_23797,N_15749,N_16500);
xnor U23798 (N_23798,N_17379,N_16538);
xnor U23799 (N_23799,N_16261,N_16572);
nand U23800 (N_23800,N_19449,N_15973);
or U23801 (N_23801,N_18768,N_15899);
or U23802 (N_23802,N_19736,N_16157);
xor U23803 (N_23803,N_19695,N_15489);
xor U23804 (N_23804,N_18713,N_17024);
and U23805 (N_23805,N_19845,N_15791);
xor U23806 (N_23806,N_17604,N_18287);
and U23807 (N_23807,N_19498,N_17832);
nor U23808 (N_23808,N_17737,N_18877);
and U23809 (N_23809,N_16500,N_16306);
xnor U23810 (N_23810,N_15125,N_17698);
and U23811 (N_23811,N_16531,N_19425);
nand U23812 (N_23812,N_15801,N_17731);
and U23813 (N_23813,N_17811,N_17607);
or U23814 (N_23814,N_15548,N_15876);
nand U23815 (N_23815,N_18059,N_18846);
and U23816 (N_23816,N_17664,N_17430);
xnor U23817 (N_23817,N_18397,N_16427);
xnor U23818 (N_23818,N_15438,N_19900);
or U23819 (N_23819,N_15558,N_19649);
and U23820 (N_23820,N_19191,N_16944);
xnor U23821 (N_23821,N_16377,N_19350);
and U23822 (N_23822,N_16985,N_16697);
or U23823 (N_23823,N_18755,N_17235);
xor U23824 (N_23824,N_18268,N_17255);
nand U23825 (N_23825,N_16220,N_15973);
or U23826 (N_23826,N_17267,N_15055);
and U23827 (N_23827,N_19274,N_15179);
nand U23828 (N_23828,N_19134,N_16386);
nor U23829 (N_23829,N_18128,N_19757);
or U23830 (N_23830,N_15036,N_19739);
and U23831 (N_23831,N_16455,N_19852);
nor U23832 (N_23832,N_17574,N_17030);
nand U23833 (N_23833,N_15612,N_19139);
or U23834 (N_23834,N_17483,N_18073);
nor U23835 (N_23835,N_17037,N_17702);
and U23836 (N_23836,N_15522,N_16285);
or U23837 (N_23837,N_17319,N_16127);
or U23838 (N_23838,N_19733,N_18839);
nor U23839 (N_23839,N_18779,N_19710);
or U23840 (N_23840,N_15275,N_16256);
or U23841 (N_23841,N_18048,N_19468);
xnor U23842 (N_23842,N_15980,N_16107);
or U23843 (N_23843,N_19528,N_19418);
nand U23844 (N_23844,N_19727,N_16509);
xnor U23845 (N_23845,N_15431,N_16082);
nand U23846 (N_23846,N_17062,N_19322);
nor U23847 (N_23847,N_17457,N_15178);
xor U23848 (N_23848,N_16668,N_17652);
or U23849 (N_23849,N_19304,N_16485);
nand U23850 (N_23850,N_16185,N_17576);
nor U23851 (N_23851,N_18309,N_18527);
nor U23852 (N_23852,N_15163,N_16057);
xnor U23853 (N_23853,N_18489,N_16414);
nor U23854 (N_23854,N_19166,N_16440);
and U23855 (N_23855,N_16613,N_16605);
or U23856 (N_23856,N_19495,N_19289);
nor U23857 (N_23857,N_19005,N_19657);
xnor U23858 (N_23858,N_18379,N_15932);
or U23859 (N_23859,N_15898,N_18473);
or U23860 (N_23860,N_18804,N_19668);
nor U23861 (N_23861,N_18730,N_16405);
xnor U23862 (N_23862,N_18344,N_19994);
nor U23863 (N_23863,N_18120,N_15267);
or U23864 (N_23864,N_17054,N_16676);
xnor U23865 (N_23865,N_19595,N_15224);
nand U23866 (N_23866,N_18816,N_16545);
nand U23867 (N_23867,N_19143,N_19974);
or U23868 (N_23868,N_15379,N_17254);
nand U23869 (N_23869,N_18425,N_15121);
nor U23870 (N_23870,N_15168,N_15400);
and U23871 (N_23871,N_17311,N_15921);
xor U23872 (N_23872,N_15063,N_19548);
nand U23873 (N_23873,N_16847,N_19886);
nand U23874 (N_23874,N_16203,N_19796);
xor U23875 (N_23875,N_15700,N_18095);
nor U23876 (N_23876,N_15350,N_16145);
nor U23877 (N_23877,N_16544,N_16090);
or U23878 (N_23878,N_18604,N_18379);
xor U23879 (N_23879,N_19021,N_19443);
nor U23880 (N_23880,N_18120,N_16515);
nand U23881 (N_23881,N_15374,N_17709);
nand U23882 (N_23882,N_19173,N_15003);
and U23883 (N_23883,N_19418,N_16827);
nor U23884 (N_23884,N_18322,N_17439);
and U23885 (N_23885,N_15165,N_19722);
xor U23886 (N_23886,N_19711,N_15125);
nor U23887 (N_23887,N_15746,N_19254);
nand U23888 (N_23888,N_16023,N_18768);
or U23889 (N_23889,N_17284,N_18078);
nand U23890 (N_23890,N_15246,N_16442);
nand U23891 (N_23891,N_17756,N_18714);
nor U23892 (N_23892,N_16509,N_19458);
nand U23893 (N_23893,N_17030,N_17656);
or U23894 (N_23894,N_19815,N_18508);
nand U23895 (N_23895,N_18471,N_17065);
and U23896 (N_23896,N_15312,N_15939);
xnor U23897 (N_23897,N_19303,N_16774);
and U23898 (N_23898,N_15879,N_15899);
xor U23899 (N_23899,N_19635,N_15622);
or U23900 (N_23900,N_17059,N_19615);
nor U23901 (N_23901,N_15881,N_19611);
nor U23902 (N_23902,N_18729,N_16625);
nor U23903 (N_23903,N_19771,N_16679);
nor U23904 (N_23904,N_19338,N_18921);
xor U23905 (N_23905,N_17413,N_16675);
nor U23906 (N_23906,N_19497,N_18707);
nand U23907 (N_23907,N_15762,N_19501);
nor U23908 (N_23908,N_18014,N_19500);
and U23909 (N_23909,N_19765,N_18030);
nor U23910 (N_23910,N_16538,N_17631);
xor U23911 (N_23911,N_18493,N_16774);
nor U23912 (N_23912,N_17252,N_16227);
or U23913 (N_23913,N_19057,N_19337);
or U23914 (N_23914,N_16026,N_18562);
or U23915 (N_23915,N_15674,N_17635);
nor U23916 (N_23916,N_16209,N_18261);
nor U23917 (N_23917,N_19853,N_17887);
nor U23918 (N_23918,N_16502,N_16709);
or U23919 (N_23919,N_15648,N_15475);
xnor U23920 (N_23920,N_19692,N_19077);
and U23921 (N_23921,N_18063,N_16635);
and U23922 (N_23922,N_18295,N_17307);
xor U23923 (N_23923,N_16655,N_18061);
nor U23924 (N_23924,N_19242,N_15746);
xor U23925 (N_23925,N_15417,N_18440);
or U23926 (N_23926,N_19899,N_17244);
nor U23927 (N_23927,N_17070,N_18533);
nand U23928 (N_23928,N_16971,N_19873);
nand U23929 (N_23929,N_15245,N_17227);
xor U23930 (N_23930,N_18478,N_15958);
nor U23931 (N_23931,N_19093,N_15317);
or U23932 (N_23932,N_19999,N_16480);
nand U23933 (N_23933,N_15897,N_16229);
xnor U23934 (N_23934,N_16463,N_18364);
nor U23935 (N_23935,N_18006,N_19206);
and U23936 (N_23936,N_18527,N_17735);
or U23937 (N_23937,N_18573,N_15088);
or U23938 (N_23938,N_16039,N_16563);
xnor U23939 (N_23939,N_16454,N_15901);
nor U23940 (N_23940,N_19656,N_15906);
xnor U23941 (N_23941,N_19826,N_16265);
and U23942 (N_23942,N_16243,N_15872);
and U23943 (N_23943,N_17186,N_18570);
xor U23944 (N_23944,N_17893,N_19341);
nor U23945 (N_23945,N_18815,N_18346);
or U23946 (N_23946,N_16308,N_18670);
or U23947 (N_23947,N_17923,N_16437);
xnor U23948 (N_23948,N_18275,N_17887);
or U23949 (N_23949,N_18318,N_15574);
xor U23950 (N_23950,N_18912,N_19692);
and U23951 (N_23951,N_18651,N_19461);
or U23952 (N_23952,N_17807,N_15191);
xnor U23953 (N_23953,N_15108,N_18171);
nor U23954 (N_23954,N_19316,N_18188);
nor U23955 (N_23955,N_19949,N_19676);
nor U23956 (N_23956,N_17987,N_16212);
and U23957 (N_23957,N_16126,N_15375);
nand U23958 (N_23958,N_16761,N_16052);
nor U23959 (N_23959,N_18198,N_15804);
xnor U23960 (N_23960,N_17864,N_15954);
nand U23961 (N_23961,N_15080,N_17316);
or U23962 (N_23962,N_16695,N_15422);
nor U23963 (N_23963,N_17461,N_15107);
nor U23964 (N_23964,N_16896,N_19436);
nor U23965 (N_23965,N_18704,N_15517);
or U23966 (N_23966,N_19612,N_18750);
nor U23967 (N_23967,N_18380,N_16232);
or U23968 (N_23968,N_17517,N_18595);
nand U23969 (N_23969,N_16661,N_15873);
xnor U23970 (N_23970,N_19893,N_17251);
and U23971 (N_23971,N_18745,N_17714);
and U23972 (N_23972,N_17139,N_17521);
xnor U23973 (N_23973,N_15011,N_18666);
nor U23974 (N_23974,N_17416,N_15850);
and U23975 (N_23975,N_16375,N_17491);
or U23976 (N_23976,N_16567,N_19682);
and U23977 (N_23977,N_15893,N_19961);
nand U23978 (N_23978,N_16607,N_18269);
nand U23979 (N_23979,N_17425,N_16424);
nand U23980 (N_23980,N_18677,N_18653);
nand U23981 (N_23981,N_18030,N_18218);
or U23982 (N_23982,N_18399,N_16539);
or U23983 (N_23983,N_17050,N_17245);
xor U23984 (N_23984,N_17546,N_18766);
nand U23985 (N_23985,N_15504,N_16198);
nor U23986 (N_23986,N_17445,N_16527);
and U23987 (N_23987,N_17018,N_17068);
nand U23988 (N_23988,N_15270,N_15698);
nand U23989 (N_23989,N_17005,N_18218);
and U23990 (N_23990,N_16638,N_19116);
nand U23991 (N_23991,N_18188,N_17567);
or U23992 (N_23992,N_15075,N_16585);
nor U23993 (N_23993,N_17522,N_17242);
or U23994 (N_23994,N_16960,N_16740);
nand U23995 (N_23995,N_19776,N_17807);
nand U23996 (N_23996,N_16605,N_16429);
xor U23997 (N_23997,N_17645,N_15114);
nor U23998 (N_23998,N_15154,N_18671);
nor U23999 (N_23999,N_16017,N_19154);
nand U24000 (N_24000,N_15345,N_18061);
nand U24001 (N_24001,N_17566,N_19490);
nand U24002 (N_24002,N_15762,N_19684);
or U24003 (N_24003,N_15278,N_15743);
nor U24004 (N_24004,N_16948,N_19894);
or U24005 (N_24005,N_16426,N_19762);
or U24006 (N_24006,N_17496,N_17961);
nor U24007 (N_24007,N_19671,N_15076);
xor U24008 (N_24008,N_15137,N_16175);
xor U24009 (N_24009,N_19268,N_19697);
xnor U24010 (N_24010,N_15831,N_15528);
and U24011 (N_24011,N_18465,N_16048);
or U24012 (N_24012,N_15951,N_18072);
nor U24013 (N_24013,N_18100,N_17029);
or U24014 (N_24014,N_15152,N_17173);
or U24015 (N_24015,N_19578,N_15190);
or U24016 (N_24016,N_15645,N_19733);
nand U24017 (N_24017,N_16678,N_15665);
nor U24018 (N_24018,N_15394,N_16106);
or U24019 (N_24019,N_16130,N_16573);
xnor U24020 (N_24020,N_19958,N_19037);
nand U24021 (N_24021,N_19742,N_15599);
and U24022 (N_24022,N_18647,N_19492);
nand U24023 (N_24023,N_15753,N_17978);
and U24024 (N_24024,N_17891,N_16209);
xnor U24025 (N_24025,N_18273,N_19160);
nand U24026 (N_24026,N_15694,N_19819);
xor U24027 (N_24027,N_16424,N_15215);
xor U24028 (N_24028,N_19703,N_19334);
nor U24029 (N_24029,N_18140,N_16839);
nor U24030 (N_24030,N_17878,N_15607);
and U24031 (N_24031,N_15166,N_19796);
or U24032 (N_24032,N_16916,N_19367);
or U24033 (N_24033,N_17534,N_17645);
and U24034 (N_24034,N_19324,N_19506);
or U24035 (N_24035,N_15557,N_16358);
xnor U24036 (N_24036,N_18610,N_15844);
nand U24037 (N_24037,N_19600,N_19036);
and U24038 (N_24038,N_17028,N_17880);
and U24039 (N_24039,N_19795,N_15720);
nor U24040 (N_24040,N_19965,N_16452);
xor U24041 (N_24041,N_19855,N_17724);
and U24042 (N_24042,N_17060,N_15568);
xnor U24043 (N_24043,N_16216,N_17587);
nand U24044 (N_24044,N_17341,N_15633);
or U24045 (N_24045,N_17936,N_19487);
nor U24046 (N_24046,N_15679,N_16868);
xnor U24047 (N_24047,N_19888,N_15784);
xnor U24048 (N_24048,N_18972,N_19052);
or U24049 (N_24049,N_19448,N_18566);
nand U24050 (N_24050,N_16781,N_18791);
nor U24051 (N_24051,N_19254,N_16401);
xor U24052 (N_24052,N_15403,N_19763);
or U24053 (N_24053,N_18577,N_18682);
nor U24054 (N_24054,N_16942,N_16649);
nor U24055 (N_24055,N_17424,N_17006);
nor U24056 (N_24056,N_15093,N_15881);
nor U24057 (N_24057,N_15171,N_19076);
nor U24058 (N_24058,N_17502,N_18648);
nor U24059 (N_24059,N_17116,N_16548);
xnor U24060 (N_24060,N_17868,N_17587);
or U24061 (N_24061,N_17803,N_19464);
and U24062 (N_24062,N_15724,N_16393);
nand U24063 (N_24063,N_19708,N_18536);
and U24064 (N_24064,N_17709,N_18395);
or U24065 (N_24065,N_15896,N_17165);
nor U24066 (N_24066,N_18457,N_17642);
xor U24067 (N_24067,N_17818,N_17469);
nor U24068 (N_24068,N_17177,N_15049);
and U24069 (N_24069,N_16848,N_16888);
nor U24070 (N_24070,N_18037,N_19238);
xor U24071 (N_24071,N_15138,N_19281);
nor U24072 (N_24072,N_18195,N_17259);
or U24073 (N_24073,N_15314,N_16169);
xnor U24074 (N_24074,N_16281,N_18517);
xnor U24075 (N_24075,N_19903,N_15163);
or U24076 (N_24076,N_19985,N_17535);
nor U24077 (N_24077,N_15211,N_18895);
and U24078 (N_24078,N_18982,N_18803);
nor U24079 (N_24079,N_19974,N_18364);
nand U24080 (N_24080,N_19695,N_17377);
or U24081 (N_24081,N_18167,N_15669);
nor U24082 (N_24082,N_16265,N_15149);
xnor U24083 (N_24083,N_17401,N_17528);
nor U24084 (N_24084,N_17558,N_17658);
or U24085 (N_24085,N_18116,N_15106);
nor U24086 (N_24086,N_18061,N_15991);
xnor U24087 (N_24087,N_19827,N_19005);
nor U24088 (N_24088,N_19500,N_18646);
xor U24089 (N_24089,N_17041,N_15108);
nand U24090 (N_24090,N_15502,N_18971);
nor U24091 (N_24091,N_18905,N_17442);
nand U24092 (N_24092,N_15031,N_15896);
nand U24093 (N_24093,N_15250,N_15216);
nand U24094 (N_24094,N_17035,N_19593);
xnor U24095 (N_24095,N_15081,N_16107);
nor U24096 (N_24096,N_19612,N_17725);
nand U24097 (N_24097,N_18562,N_18416);
nand U24098 (N_24098,N_18111,N_16399);
and U24099 (N_24099,N_17276,N_17858);
xnor U24100 (N_24100,N_18902,N_17357);
or U24101 (N_24101,N_16822,N_18393);
xnor U24102 (N_24102,N_17988,N_19589);
or U24103 (N_24103,N_17283,N_19483);
and U24104 (N_24104,N_18580,N_15879);
nor U24105 (N_24105,N_18830,N_19059);
nand U24106 (N_24106,N_15449,N_17208);
nor U24107 (N_24107,N_18945,N_19443);
or U24108 (N_24108,N_19313,N_19404);
nor U24109 (N_24109,N_19804,N_18648);
nand U24110 (N_24110,N_16941,N_16407);
and U24111 (N_24111,N_17730,N_16067);
nand U24112 (N_24112,N_15231,N_17489);
and U24113 (N_24113,N_16907,N_17163);
nor U24114 (N_24114,N_15548,N_16873);
nor U24115 (N_24115,N_18012,N_17232);
nor U24116 (N_24116,N_18246,N_15618);
xnor U24117 (N_24117,N_16740,N_19469);
nor U24118 (N_24118,N_15473,N_18745);
and U24119 (N_24119,N_18663,N_19619);
nor U24120 (N_24120,N_18713,N_15785);
or U24121 (N_24121,N_18978,N_16624);
or U24122 (N_24122,N_16994,N_17796);
or U24123 (N_24123,N_16996,N_15319);
nor U24124 (N_24124,N_19970,N_15820);
xor U24125 (N_24125,N_17819,N_19403);
xnor U24126 (N_24126,N_18296,N_17987);
or U24127 (N_24127,N_15684,N_19095);
nor U24128 (N_24128,N_15963,N_19400);
nand U24129 (N_24129,N_18943,N_15223);
or U24130 (N_24130,N_18405,N_18207);
nor U24131 (N_24131,N_17537,N_17941);
nand U24132 (N_24132,N_15808,N_18574);
and U24133 (N_24133,N_16417,N_18741);
and U24134 (N_24134,N_18972,N_15371);
nand U24135 (N_24135,N_18387,N_18745);
nand U24136 (N_24136,N_16205,N_15957);
and U24137 (N_24137,N_15168,N_16764);
and U24138 (N_24138,N_16721,N_19391);
and U24139 (N_24139,N_19975,N_15452);
nand U24140 (N_24140,N_17278,N_19617);
nor U24141 (N_24141,N_18973,N_18404);
nand U24142 (N_24142,N_16206,N_16003);
and U24143 (N_24143,N_17885,N_17088);
and U24144 (N_24144,N_18833,N_17477);
xnor U24145 (N_24145,N_16593,N_18621);
nand U24146 (N_24146,N_18639,N_15243);
xnor U24147 (N_24147,N_15761,N_15231);
nor U24148 (N_24148,N_17767,N_19323);
or U24149 (N_24149,N_17842,N_17551);
and U24150 (N_24150,N_18086,N_18417);
nor U24151 (N_24151,N_15631,N_18744);
or U24152 (N_24152,N_18500,N_18592);
nand U24153 (N_24153,N_17900,N_19915);
and U24154 (N_24154,N_16172,N_19633);
nor U24155 (N_24155,N_16748,N_17842);
or U24156 (N_24156,N_18399,N_16179);
nor U24157 (N_24157,N_17891,N_18576);
or U24158 (N_24158,N_15820,N_16910);
and U24159 (N_24159,N_18378,N_17891);
and U24160 (N_24160,N_16601,N_19407);
and U24161 (N_24161,N_17609,N_19181);
nor U24162 (N_24162,N_15759,N_16443);
or U24163 (N_24163,N_15020,N_18936);
and U24164 (N_24164,N_19909,N_15884);
nand U24165 (N_24165,N_15790,N_18671);
xor U24166 (N_24166,N_15502,N_17298);
nand U24167 (N_24167,N_19985,N_15517);
and U24168 (N_24168,N_16298,N_17002);
nand U24169 (N_24169,N_15661,N_15633);
xnor U24170 (N_24170,N_18513,N_15127);
xor U24171 (N_24171,N_17452,N_16060);
nand U24172 (N_24172,N_15954,N_17228);
nor U24173 (N_24173,N_15853,N_15690);
or U24174 (N_24174,N_15539,N_16453);
nand U24175 (N_24175,N_15323,N_17441);
or U24176 (N_24176,N_16507,N_18089);
or U24177 (N_24177,N_18155,N_16507);
nor U24178 (N_24178,N_15788,N_17313);
nor U24179 (N_24179,N_16304,N_18247);
nor U24180 (N_24180,N_17377,N_19129);
and U24181 (N_24181,N_19811,N_19330);
or U24182 (N_24182,N_15146,N_17428);
and U24183 (N_24183,N_17789,N_18308);
and U24184 (N_24184,N_17564,N_18682);
nand U24185 (N_24185,N_15574,N_16569);
nand U24186 (N_24186,N_17865,N_15986);
xnor U24187 (N_24187,N_16397,N_16773);
xnor U24188 (N_24188,N_17881,N_16128);
nand U24189 (N_24189,N_15502,N_17290);
nor U24190 (N_24190,N_17720,N_15664);
and U24191 (N_24191,N_19238,N_18652);
nand U24192 (N_24192,N_17850,N_16790);
and U24193 (N_24193,N_16436,N_16641);
and U24194 (N_24194,N_19075,N_15443);
nor U24195 (N_24195,N_16694,N_16942);
nor U24196 (N_24196,N_17993,N_18966);
xnor U24197 (N_24197,N_17484,N_15199);
or U24198 (N_24198,N_16583,N_16821);
nand U24199 (N_24199,N_19122,N_19471);
nand U24200 (N_24200,N_17234,N_16509);
xnor U24201 (N_24201,N_18132,N_16975);
or U24202 (N_24202,N_19924,N_17645);
nor U24203 (N_24203,N_17740,N_15224);
or U24204 (N_24204,N_19324,N_19022);
and U24205 (N_24205,N_16858,N_19162);
xor U24206 (N_24206,N_18887,N_18155);
nand U24207 (N_24207,N_16061,N_16990);
and U24208 (N_24208,N_15747,N_19315);
or U24209 (N_24209,N_15132,N_16859);
xor U24210 (N_24210,N_15487,N_17086);
nor U24211 (N_24211,N_15288,N_19737);
nor U24212 (N_24212,N_16509,N_16478);
nor U24213 (N_24213,N_17450,N_18748);
nand U24214 (N_24214,N_18472,N_15668);
or U24215 (N_24215,N_17297,N_16418);
nand U24216 (N_24216,N_16267,N_19425);
nor U24217 (N_24217,N_15596,N_16441);
or U24218 (N_24218,N_17355,N_18967);
nor U24219 (N_24219,N_15338,N_19047);
xor U24220 (N_24220,N_16060,N_18267);
nand U24221 (N_24221,N_19674,N_17970);
nor U24222 (N_24222,N_19386,N_19826);
and U24223 (N_24223,N_15060,N_19019);
nor U24224 (N_24224,N_17278,N_15522);
xnor U24225 (N_24225,N_17628,N_16399);
and U24226 (N_24226,N_16344,N_18535);
and U24227 (N_24227,N_19681,N_17972);
xor U24228 (N_24228,N_18130,N_16316);
nand U24229 (N_24229,N_15508,N_19772);
nand U24230 (N_24230,N_18827,N_17023);
nor U24231 (N_24231,N_17752,N_16240);
nand U24232 (N_24232,N_19195,N_18800);
and U24233 (N_24233,N_17550,N_15267);
xor U24234 (N_24234,N_17572,N_16774);
and U24235 (N_24235,N_17645,N_15866);
and U24236 (N_24236,N_15935,N_16883);
nand U24237 (N_24237,N_15007,N_15162);
or U24238 (N_24238,N_19690,N_17901);
nand U24239 (N_24239,N_17893,N_15664);
and U24240 (N_24240,N_17974,N_15884);
nor U24241 (N_24241,N_19443,N_19601);
or U24242 (N_24242,N_19094,N_15137);
nand U24243 (N_24243,N_18054,N_16236);
or U24244 (N_24244,N_15544,N_18182);
xor U24245 (N_24245,N_19134,N_15394);
or U24246 (N_24246,N_17851,N_15961);
xor U24247 (N_24247,N_17156,N_18717);
xnor U24248 (N_24248,N_17297,N_16753);
nor U24249 (N_24249,N_15833,N_17107);
nor U24250 (N_24250,N_18348,N_15235);
nor U24251 (N_24251,N_16923,N_16018);
nor U24252 (N_24252,N_19490,N_15709);
or U24253 (N_24253,N_15828,N_19009);
and U24254 (N_24254,N_18683,N_19577);
xor U24255 (N_24255,N_16992,N_16312);
and U24256 (N_24256,N_15081,N_16744);
and U24257 (N_24257,N_15092,N_15769);
nand U24258 (N_24258,N_16571,N_16998);
or U24259 (N_24259,N_16145,N_15620);
or U24260 (N_24260,N_19308,N_17305);
or U24261 (N_24261,N_19564,N_19738);
xor U24262 (N_24262,N_15202,N_19071);
nand U24263 (N_24263,N_18594,N_15468);
nor U24264 (N_24264,N_17236,N_16445);
xor U24265 (N_24265,N_16359,N_17671);
xor U24266 (N_24266,N_17170,N_19615);
nor U24267 (N_24267,N_17549,N_19442);
or U24268 (N_24268,N_15819,N_18412);
xnor U24269 (N_24269,N_19921,N_17074);
or U24270 (N_24270,N_19047,N_16777);
and U24271 (N_24271,N_16105,N_19393);
xor U24272 (N_24272,N_16022,N_15873);
nand U24273 (N_24273,N_17857,N_18185);
nand U24274 (N_24274,N_18169,N_16695);
nor U24275 (N_24275,N_19183,N_15748);
and U24276 (N_24276,N_15052,N_15672);
nand U24277 (N_24277,N_15044,N_19737);
and U24278 (N_24278,N_15772,N_16070);
nand U24279 (N_24279,N_16822,N_19372);
nor U24280 (N_24280,N_16674,N_15680);
xnor U24281 (N_24281,N_19934,N_16208);
or U24282 (N_24282,N_19868,N_19702);
xnor U24283 (N_24283,N_15714,N_17666);
and U24284 (N_24284,N_19798,N_18661);
xor U24285 (N_24285,N_17011,N_15318);
xnor U24286 (N_24286,N_16040,N_17643);
and U24287 (N_24287,N_19977,N_17799);
or U24288 (N_24288,N_18007,N_15495);
nand U24289 (N_24289,N_16489,N_16019);
nand U24290 (N_24290,N_16492,N_17647);
or U24291 (N_24291,N_18971,N_19869);
xnor U24292 (N_24292,N_17622,N_19075);
and U24293 (N_24293,N_17189,N_19784);
nand U24294 (N_24294,N_19928,N_18508);
or U24295 (N_24295,N_19534,N_19739);
xor U24296 (N_24296,N_19707,N_18532);
xor U24297 (N_24297,N_19817,N_15808);
or U24298 (N_24298,N_19123,N_17849);
nor U24299 (N_24299,N_19080,N_18485);
nand U24300 (N_24300,N_16659,N_17485);
or U24301 (N_24301,N_15347,N_15727);
nor U24302 (N_24302,N_15842,N_15716);
nand U24303 (N_24303,N_16419,N_15195);
xor U24304 (N_24304,N_16693,N_17621);
or U24305 (N_24305,N_18752,N_18370);
nor U24306 (N_24306,N_15178,N_17770);
nor U24307 (N_24307,N_16665,N_15841);
xor U24308 (N_24308,N_15220,N_15445);
and U24309 (N_24309,N_16242,N_15828);
or U24310 (N_24310,N_16524,N_19854);
xnor U24311 (N_24311,N_18087,N_17227);
or U24312 (N_24312,N_16680,N_19511);
or U24313 (N_24313,N_19724,N_19254);
nor U24314 (N_24314,N_18806,N_16471);
nand U24315 (N_24315,N_15040,N_19603);
and U24316 (N_24316,N_17576,N_19084);
nand U24317 (N_24317,N_19794,N_19049);
and U24318 (N_24318,N_17593,N_16656);
nor U24319 (N_24319,N_17297,N_19345);
or U24320 (N_24320,N_16537,N_17022);
nor U24321 (N_24321,N_16760,N_15523);
nor U24322 (N_24322,N_15772,N_18103);
or U24323 (N_24323,N_16718,N_18570);
nand U24324 (N_24324,N_19080,N_19527);
xnor U24325 (N_24325,N_16675,N_15237);
nand U24326 (N_24326,N_15719,N_15534);
xor U24327 (N_24327,N_17645,N_15743);
xnor U24328 (N_24328,N_15780,N_19805);
xor U24329 (N_24329,N_17731,N_15835);
or U24330 (N_24330,N_17270,N_17941);
or U24331 (N_24331,N_19975,N_18927);
or U24332 (N_24332,N_15078,N_17764);
xnor U24333 (N_24333,N_19598,N_16374);
or U24334 (N_24334,N_19969,N_15086);
xnor U24335 (N_24335,N_15257,N_16008);
xnor U24336 (N_24336,N_16128,N_17227);
xnor U24337 (N_24337,N_16363,N_15130);
nor U24338 (N_24338,N_19480,N_17518);
and U24339 (N_24339,N_16678,N_15322);
nor U24340 (N_24340,N_15111,N_16978);
nand U24341 (N_24341,N_17515,N_16647);
nand U24342 (N_24342,N_17872,N_15723);
or U24343 (N_24343,N_18136,N_15513);
and U24344 (N_24344,N_18868,N_18866);
and U24345 (N_24345,N_19842,N_19273);
nand U24346 (N_24346,N_19383,N_16142);
and U24347 (N_24347,N_17741,N_19412);
nand U24348 (N_24348,N_19809,N_17397);
or U24349 (N_24349,N_18716,N_16298);
and U24350 (N_24350,N_16336,N_18891);
xnor U24351 (N_24351,N_15664,N_18410);
and U24352 (N_24352,N_17852,N_18504);
xnor U24353 (N_24353,N_19253,N_18618);
or U24354 (N_24354,N_19129,N_16748);
xor U24355 (N_24355,N_19495,N_19979);
nand U24356 (N_24356,N_19991,N_19087);
xor U24357 (N_24357,N_16512,N_16684);
or U24358 (N_24358,N_16411,N_15719);
and U24359 (N_24359,N_17388,N_19429);
xnor U24360 (N_24360,N_19219,N_15536);
nand U24361 (N_24361,N_17178,N_16925);
nand U24362 (N_24362,N_19081,N_18865);
xnor U24363 (N_24363,N_17003,N_18614);
or U24364 (N_24364,N_18745,N_15692);
nand U24365 (N_24365,N_19226,N_18120);
xnor U24366 (N_24366,N_16717,N_17012);
xnor U24367 (N_24367,N_18309,N_19972);
nor U24368 (N_24368,N_16814,N_19770);
nor U24369 (N_24369,N_15976,N_17010);
nand U24370 (N_24370,N_16483,N_16659);
xnor U24371 (N_24371,N_19863,N_19881);
nand U24372 (N_24372,N_15327,N_16445);
or U24373 (N_24373,N_16324,N_15844);
xor U24374 (N_24374,N_15962,N_19731);
or U24375 (N_24375,N_16149,N_17701);
or U24376 (N_24376,N_15137,N_15128);
and U24377 (N_24377,N_19573,N_16581);
and U24378 (N_24378,N_15609,N_15993);
nor U24379 (N_24379,N_15264,N_16367);
or U24380 (N_24380,N_16503,N_17464);
nor U24381 (N_24381,N_15630,N_18897);
or U24382 (N_24382,N_19579,N_19995);
and U24383 (N_24383,N_15785,N_17731);
xnor U24384 (N_24384,N_16447,N_16181);
and U24385 (N_24385,N_17119,N_19139);
nand U24386 (N_24386,N_19103,N_15276);
and U24387 (N_24387,N_17452,N_18005);
and U24388 (N_24388,N_15964,N_17842);
or U24389 (N_24389,N_16465,N_17553);
nor U24390 (N_24390,N_17602,N_17411);
nand U24391 (N_24391,N_16876,N_17487);
nor U24392 (N_24392,N_19292,N_17582);
xor U24393 (N_24393,N_15738,N_15068);
or U24394 (N_24394,N_15614,N_15918);
xnor U24395 (N_24395,N_19027,N_18991);
xnor U24396 (N_24396,N_18571,N_19837);
xor U24397 (N_24397,N_18909,N_16294);
nand U24398 (N_24398,N_15250,N_16359);
xor U24399 (N_24399,N_17186,N_18037);
or U24400 (N_24400,N_15288,N_18661);
nand U24401 (N_24401,N_18155,N_17183);
and U24402 (N_24402,N_18167,N_18328);
or U24403 (N_24403,N_19384,N_19160);
nor U24404 (N_24404,N_16113,N_19306);
xnor U24405 (N_24405,N_18754,N_19568);
xor U24406 (N_24406,N_15329,N_18613);
or U24407 (N_24407,N_18740,N_19007);
or U24408 (N_24408,N_16638,N_19969);
or U24409 (N_24409,N_16451,N_18689);
xnor U24410 (N_24410,N_17821,N_19624);
or U24411 (N_24411,N_15986,N_15009);
nand U24412 (N_24412,N_19151,N_16358);
nor U24413 (N_24413,N_15844,N_18645);
or U24414 (N_24414,N_19743,N_15230);
and U24415 (N_24415,N_18070,N_16970);
or U24416 (N_24416,N_17974,N_15092);
and U24417 (N_24417,N_15219,N_19197);
xnor U24418 (N_24418,N_17647,N_16400);
xor U24419 (N_24419,N_17983,N_15062);
nand U24420 (N_24420,N_15881,N_18646);
or U24421 (N_24421,N_18567,N_16467);
or U24422 (N_24422,N_19483,N_16647);
or U24423 (N_24423,N_17987,N_16300);
nand U24424 (N_24424,N_18066,N_15861);
and U24425 (N_24425,N_15014,N_16232);
and U24426 (N_24426,N_19179,N_19428);
or U24427 (N_24427,N_15883,N_17545);
nand U24428 (N_24428,N_18723,N_18343);
xor U24429 (N_24429,N_15987,N_19793);
and U24430 (N_24430,N_16223,N_19033);
and U24431 (N_24431,N_16751,N_19787);
and U24432 (N_24432,N_15428,N_17816);
nor U24433 (N_24433,N_17173,N_15924);
and U24434 (N_24434,N_15564,N_18521);
nor U24435 (N_24435,N_15068,N_17194);
or U24436 (N_24436,N_15850,N_17627);
nor U24437 (N_24437,N_19787,N_16953);
or U24438 (N_24438,N_17039,N_18763);
or U24439 (N_24439,N_16323,N_15490);
nand U24440 (N_24440,N_19283,N_16514);
xor U24441 (N_24441,N_19118,N_17144);
and U24442 (N_24442,N_18596,N_16909);
xnor U24443 (N_24443,N_17170,N_15298);
xor U24444 (N_24444,N_16173,N_15875);
nor U24445 (N_24445,N_17470,N_15301);
and U24446 (N_24446,N_16909,N_18348);
nand U24447 (N_24447,N_15342,N_15841);
or U24448 (N_24448,N_19951,N_19762);
xor U24449 (N_24449,N_18701,N_15605);
xor U24450 (N_24450,N_15145,N_19911);
and U24451 (N_24451,N_17225,N_19697);
and U24452 (N_24452,N_19754,N_15943);
nand U24453 (N_24453,N_19918,N_15397);
and U24454 (N_24454,N_17567,N_15292);
nand U24455 (N_24455,N_19913,N_15253);
xnor U24456 (N_24456,N_15951,N_19599);
nor U24457 (N_24457,N_19285,N_15996);
xor U24458 (N_24458,N_16856,N_19576);
nor U24459 (N_24459,N_15754,N_17246);
or U24460 (N_24460,N_17733,N_18536);
or U24461 (N_24461,N_17835,N_16462);
xnor U24462 (N_24462,N_15759,N_18620);
nand U24463 (N_24463,N_19614,N_19202);
or U24464 (N_24464,N_17590,N_15661);
or U24465 (N_24465,N_18880,N_16363);
nand U24466 (N_24466,N_19288,N_15930);
nand U24467 (N_24467,N_19306,N_15870);
and U24468 (N_24468,N_19567,N_17287);
or U24469 (N_24469,N_16429,N_16615);
xnor U24470 (N_24470,N_18184,N_19285);
nor U24471 (N_24471,N_18752,N_19533);
and U24472 (N_24472,N_19573,N_17494);
xor U24473 (N_24473,N_18990,N_19861);
or U24474 (N_24474,N_18656,N_18790);
xnor U24475 (N_24475,N_16255,N_19635);
xor U24476 (N_24476,N_16695,N_18583);
nor U24477 (N_24477,N_19998,N_16742);
or U24478 (N_24478,N_19619,N_15923);
nor U24479 (N_24479,N_16750,N_16197);
nor U24480 (N_24480,N_15046,N_15670);
or U24481 (N_24481,N_18637,N_15652);
xnor U24482 (N_24482,N_19680,N_17734);
or U24483 (N_24483,N_18423,N_19759);
xnor U24484 (N_24484,N_18954,N_16800);
nand U24485 (N_24485,N_19346,N_19875);
or U24486 (N_24486,N_17442,N_19293);
nand U24487 (N_24487,N_15293,N_19660);
and U24488 (N_24488,N_18575,N_15102);
nand U24489 (N_24489,N_17551,N_18128);
nor U24490 (N_24490,N_18821,N_17011);
xor U24491 (N_24491,N_18938,N_19737);
nor U24492 (N_24492,N_15294,N_17154);
nand U24493 (N_24493,N_18131,N_16906);
or U24494 (N_24494,N_15808,N_16711);
xnor U24495 (N_24495,N_16564,N_15267);
xor U24496 (N_24496,N_16836,N_17811);
nor U24497 (N_24497,N_16860,N_19817);
xnor U24498 (N_24498,N_17988,N_16994);
nand U24499 (N_24499,N_16571,N_19096);
xor U24500 (N_24500,N_15945,N_18739);
or U24501 (N_24501,N_18535,N_18242);
and U24502 (N_24502,N_17558,N_15800);
and U24503 (N_24503,N_18153,N_17600);
or U24504 (N_24504,N_15308,N_19235);
and U24505 (N_24505,N_19553,N_16290);
xnor U24506 (N_24506,N_16838,N_15169);
nor U24507 (N_24507,N_17779,N_18946);
or U24508 (N_24508,N_18565,N_19960);
or U24509 (N_24509,N_19354,N_15860);
nor U24510 (N_24510,N_16738,N_15373);
or U24511 (N_24511,N_16530,N_15286);
or U24512 (N_24512,N_18882,N_17208);
nor U24513 (N_24513,N_16058,N_17677);
and U24514 (N_24514,N_19374,N_18467);
nand U24515 (N_24515,N_19745,N_15519);
nor U24516 (N_24516,N_17882,N_16664);
and U24517 (N_24517,N_17437,N_16881);
nor U24518 (N_24518,N_18530,N_19458);
xor U24519 (N_24519,N_16780,N_17347);
nor U24520 (N_24520,N_18276,N_16901);
xnor U24521 (N_24521,N_17725,N_15525);
xnor U24522 (N_24522,N_18604,N_16367);
and U24523 (N_24523,N_15736,N_19101);
nand U24524 (N_24524,N_18254,N_15858);
or U24525 (N_24525,N_18201,N_18559);
xor U24526 (N_24526,N_15436,N_17172);
and U24527 (N_24527,N_16369,N_18396);
or U24528 (N_24528,N_15418,N_15896);
or U24529 (N_24529,N_19269,N_18958);
nor U24530 (N_24530,N_17346,N_18679);
nor U24531 (N_24531,N_17026,N_15360);
or U24532 (N_24532,N_17422,N_15957);
nand U24533 (N_24533,N_15174,N_16733);
nand U24534 (N_24534,N_16068,N_17518);
nor U24535 (N_24535,N_19863,N_15499);
nor U24536 (N_24536,N_19590,N_18833);
nor U24537 (N_24537,N_19802,N_17436);
or U24538 (N_24538,N_16222,N_17190);
nand U24539 (N_24539,N_18595,N_19992);
nand U24540 (N_24540,N_16151,N_17310);
and U24541 (N_24541,N_17866,N_19297);
and U24542 (N_24542,N_18786,N_18093);
nor U24543 (N_24543,N_19288,N_17218);
and U24544 (N_24544,N_17727,N_19002);
xor U24545 (N_24545,N_18191,N_17057);
nor U24546 (N_24546,N_15610,N_17281);
nand U24547 (N_24547,N_17351,N_16925);
nand U24548 (N_24548,N_18273,N_16696);
nor U24549 (N_24549,N_16376,N_16028);
nand U24550 (N_24550,N_17427,N_16093);
nand U24551 (N_24551,N_16506,N_19852);
and U24552 (N_24552,N_16869,N_16105);
and U24553 (N_24553,N_15871,N_16723);
xnor U24554 (N_24554,N_15986,N_16466);
nor U24555 (N_24555,N_18464,N_18784);
nor U24556 (N_24556,N_18116,N_18736);
nor U24557 (N_24557,N_16304,N_16403);
nand U24558 (N_24558,N_16267,N_19992);
xor U24559 (N_24559,N_18139,N_17021);
and U24560 (N_24560,N_19071,N_18780);
nor U24561 (N_24561,N_16171,N_15361);
nor U24562 (N_24562,N_16776,N_19872);
xor U24563 (N_24563,N_17388,N_15686);
xnor U24564 (N_24564,N_18109,N_18060);
nor U24565 (N_24565,N_16841,N_17260);
xor U24566 (N_24566,N_17016,N_17558);
nand U24567 (N_24567,N_15458,N_17315);
xnor U24568 (N_24568,N_17092,N_16355);
and U24569 (N_24569,N_15653,N_19347);
xnor U24570 (N_24570,N_16711,N_18406);
nor U24571 (N_24571,N_17291,N_19866);
xnor U24572 (N_24572,N_19447,N_16543);
nand U24573 (N_24573,N_17995,N_16504);
xnor U24574 (N_24574,N_16128,N_16179);
nor U24575 (N_24575,N_19960,N_15385);
xnor U24576 (N_24576,N_15752,N_18593);
or U24577 (N_24577,N_18299,N_15478);
or U24578 (N_24578,N_18811,N_16015);
or U24579 (N_24579,N_16346,N_17778);
and U24580 (N_24580,N_18193,N_15226);
nor U24581 (N_24581,N_19712,N_17081);
xor U24582 (N_24582,N_18465,N_17012);
nand U24583 (N_24583,N_15213,N_17172);
nor U24584 (N_24584,N_19411,N_16598);
and U24585 (N_24585,N_17097,N_19393);
nor U24586 (N_24586,N_19026,N_19475);
nor U24587 (N_24587,N_19366,N_17017);
xor U24588 (N_24588,N_16238,N_18997);
nor U24589 (N_24589,N_17506,N_19732);
xnor U24590 (N_24590,N_18348,N_19086);
nand U24591 (N_24591,N_18635,N_19596);
nor U24592 (N_24592,N_15709,N_18846);
nor U24593 (N_24593,N_16402,N_18019);
xor U24594 (N_24594,N_18238,N_17476);
nand U24595 (N_24595,N_17041,N_18249);
xnor U24596 (N_24596,N_17017,N_19487);
or U24597 (N_24597,N_18476,N_15198);
nand U24598 (N_24598,N_18883,N_15006);
or U24599 (N_24599,N_19222,N_18585);
or U24600 (N_24600,N_17267,N_16828);
or U24601 (N_24601,N_19794,N_18293);
or U24602 (N_24602,N_17406,N_16664);
nor U24603 (N_24603,N_17682,N_17023);
or U24604 (N_24604,N_15394,N_19512);
or U24605 (N_24605,N_19369,N_17536);
nand U24606 (N_24606,N_16030,N_15452);
xor U24607 (N_24607,N_18405,N_19822);
nand U24608 (N_24608,N_15424,N_16735);
xnor U24609 (N_24609,N_15341,N_19527);
and U24610 (N_24610,N_19023,N_18108);
xnor U24611 (N_24611,N_15631,N_17996);
nor U24612 (N_24612,N_15479,N_16554);
and U24613 (N_24613,N_18319,N_17411);
nor U24614 (N_24614,N_15260,N_18101);
xor U24615 (N_24615,N_15457,N_19105);
or U24616 (N_24616,N_19839,N_18164);
nor U24617 (N_24617,N_18817,N_18506);
or U24618 (N_24618,N_16877,N_18976);
or U24619 (N_24619,N_16499,N_17965);
nor U24620 (N_24620,N_17718,N_17736);
and U24621 (N_24621,N_15566,N_18085);
nand U24622 (N_24622,N_16986,N_18657);
and U24623 (N_24623,N_17549,N_17167);
nand U24624 (N_24624,N_16156,N_19768);
nor U24625 (N_24625,N_17565,N_15328);
nor U24626 (N_24626,N_19759,N_18984);
nand U24627 (N_24627,N_18887,N_16324);
or U24628 (N_24628,N_15083,N_18606);
and U24629 (N_24629,N_18560,N_17687);
xnor U24630 (N_24630,N_15340,N_15857);
xnor U24631 (N_24631,N_19842,N_15117);
nor U24632 (N_24632,N_19282,N_16067);
nor U24633 (N_24633,N_16597,N_17228);
nand U24634 (N_24634,N_19171,N_15932);
and U24635 (N_24635,N_15074,N_19542);
nor U24636 (N_24636,N_17047,N_16480);
nand U24637 (N_24637,N_18942,N_16538);
xnor U24638 (N_24638,N_18646,N_18788);
nor U24639 (N_24639,N_15032,N_18622);
and U24640 (N_24640,N_16937,N_18494);
nor U24641 (N_24641,N_19834,N_18880);
nor U24642 (N_24642,N_15455,N_18796);
nor U24643 (N_24643,N_18192,N_16329);
nor U24644 (N_24644,N_19483,N_19852);
nor U24645 (N_24645,N_19614,N_18324);
or U24646 (N_24646,N_16114,N_16369);
nor U24647 (N_24647,N_15475,N_15812);
nor U24648 (N_24648,N_18582,N_15840);
or U24649 (N_24649,N_18409,N_16939);
nand U24650 (N_24650,N_15740,N_17642);
xnor U24651 (N_24651,N_15182,N_17474);
xor U24652 (N_24652,N_17048,N_19251);
nor U24653 (N_24653,N_15318,N_17557);
or U24654 (N_24654,N_17963,N_18139);
nand U24655 (N_24655,N_15441,N_18316);
and U24656 (N_24656,N_17640,N_17538);
and U24657 (N_24657,N_19856,N_18550);
or U24658 (N_24658,N_16756,N_17945);
nor U24659 (N_24659,N_18091,N_19140);
and U24660 (N_24660,N_16827,N_16540);
nor U24661 (N_24661,N_15249,N_16894);
and U24662 (N_24662,N_17018,N_18936);
nor U24663 (N_24663,N_18074,N_19250);
nand U24664 (N_24664,N_17485,N_16952);
or U24665 (N_24665,N_17585,N_18937);
xnor U24666 (N_24666,N_19941,N_16702);
xnor U24667 (N_24667,N_19977,N_18394);
nand U24668 (N_24668,N_15718,N_16914);
or U24669 (N_24669,N_18223,N_17037);
nor U24670 (N_24670,N_19445,N_15109);
and U24671 (N_24671,N_16695,N_17775);
xnor U24672 (N_24672,N_18052,N_19650);
or U24673 (N_24673,N_16066,N_19537);
nor U24674 (N_24674,N_19723,N_16436);
nand U24675 (N_24675,N_15556,N_16755);
nor U24676 (N_24676,N_18389,N_17851);
xnor U24677 (N_24677,N_18210,N_16469);
nor U24678 (N_24678,N_18635,N_19401);
nor U24679 (N_24679,N_17226,N_18712);
nand U24680 (N_24680,N_19954,N_17985);
nand U24681 (N_24681,N_18526,N_15438);
nor U24682 (N_24682,N_19738,N_19666);
nand U24683 (N_24683,N_19061,N_17733);
nor U24684 (N_24684,N_18131,N_18839);
xor U24685 (N_24685,N_15050,N_19655);
nor U24686 (N_24686,N_15144,N_15589);
xnor U24687 (N_24687,N_19211,N_17117);
and U24688 (N_24688,N_15043,N_16684);
xor U24689 (N_24689,N_19964,N_16183);
nor U24690 (N_24690,N_19030,N_16465);
nand U24691 (N_24691,N_18196,N_19347);
nor U24692 (N_24692,N_19097,N_15949);
nand U24693 (N_24693,N_15772,N_19841);
nand U24694 (N_24694,N_18322,N_18585);
nor U24695 (N_24695,N_18394,N_15157);
xor U24696 (N_24696,N_18377,N_18583);
and U24697 (N_24697,N_15976,N_16222);
nand U24698 (N_24698,N_16049,N_19442);
xor U24699 (N_24699,N_16728,N_15502);
xnor U24700 (N_24700,N_17208,N_18455);
and U24701 (N_24701,N_15137,N_19883);
nor U24702 (N_24702,N_16914,N_18092);
and U24703 (N_24703,N_19460,N_18488);
xor U24704 (N_24704,N_17663,N_16805);
xor U24705 (N_24705,N_18809,N_17251);
nor U24706 (N_24706,N_19581,N_19976);
nand U24707 (N_24707,N_17944,N_18414);
nand U24708 (N_24708,N_19311,N_15275);
or U24709 (N_24709,N_15541,N_17271);
nand U24710 (N_24710,N_17020,N_19802);
or U24711 (N_24711,N_15478,N_17921);
xor U24712 (N_24712,N_18267,N_15925);
xnor U24713 (N_24713,N_19843,N_16405);
xnor U24714 (N_24714,N_15007,N_16370);
nand U24715 (N_24715,N_19527,N_16074);
or U24716 (N_24716,N_19205,N_15922);
xnor U24717 (N_24717,N_16181,N_18682);
or U24718 (N_24718,N_15220,N_18805);
and U24719 (N_24719,N_18497,N_17113);
or U24720 (N_24720,N_19206,N_16529);
nand U24721 (N_24721,N_17919,N_16748);
xnor U24722 (N_24722,N_16622,N_15181);
nor U24723 (N_24723,N_15808,N_19155);
xor U24724 (N_24724,N_17296,N_16711);
xnor U24725 (N_24725,N_17928,N_16572);
nand U24726 (N_24726,N_16326,N_18675);
and U24727 (N_24727,N_18232,N_16680);
xor U24728 (N_24728,N_18459,N_18938);
xnor U24729 (N_24729,N_17250,N_18789);
xor U24730 (N_24730,N_17785,N_16057);
nor U24731 (N_24731,N_18240,N_19992);
nand U24732 (N_24732,N_16595,N_15899);
and U24733 (N_24733,N_15491,N_15351);
and U24734 (N_24734,N_18012,N_18959);
or U24735 (N_24735,N_17953,N_15031);
nor U24736 (N_24736,N_19010,N_18470);
nand U24737 (N_24737,N_15722,N_18341);
nand U24738 (N_24738,N_18719,N_15180);
or U24739 (N_24739,N_19876,N_15474);
and U24740 (N_24740,N_15204,N_18389);
nand U24741 (N_24741,N_19007,N_19422);
nand U24742 (N_24742,N_17530,N_19633);
nor U24743 (N_24743,N_17191,N_16253);
nand U24744 (N_24744,N_18303,N_19960);
or U24745 (N_24745,N_15591,N_16077);
nor U24746 (N_24746,N_19511,N_19490);
nor U24747 (N_24747,N_16242,N_16673);
xnor U24748 (N_24748,N_15077,N_19411);
and U24749 (N_24749,N_15808,N_19457);
or U24750 (N_24750,N_17810,N_19507);
nand U24751 (N_24751,N_16220,N_16247);
nand U24752 (N_24752,N_16612,N_19662);
nor U24753 (N_24753,N_18244,N_18412);
nor U24754 (N_24754,N_15196,N_17053);
or U24755 (N_24755,N_18032,N_15606);
or U24756 (N_24756,N_16732,N_16365);
nand U24757 (N_24757,N_19969,N_16752);
xor U24758 (N_24758,N_19703,N_17989);
or U24759 (N_24759,N_17055,N_19730);
xor U24760 (N_24760,N_16254,N_18743);
xnor U24761 (N_24761,N_17943,N_19090);
nand U24762 (N_24762,N_18407,N_18263);
or U24763 (N_24763,N_17031,N_19494);
nor U24764 (N_24764,N_18891,N_19013);
nor U24765 (N_24765,N_15900,N_16601);
xor U24766 (N_24766,N_16905,N_18849);
and U24767 (N_24767,N_15356,N_18956);
nand U24768 (N_24768,N_15027,N_19801);
or U24769 (N_24769,N_17532,N_17543);
xor U24770 (N_24770,N_18031,N_18191);
nand U24771 (N_24771,N_16681,N_16987);
nand U24772 (N_24772,N_19359,N_19531);
xor U24773 (N_24773,N_17579,N_16380);
and U24774 (N_24774,N_15399,N_18024);
and U24775 (N_24775,N_18342,N_19035);
nor U24776 (N_24776,N_15641,N_18305);
xor U24777 (N_24777,N_18936,N_16596);
xnor U24778 (N_24778,N_19970,N_16503);
nand U24779 (N_24779,N_18505,N_15240);
nand U24780 (N_24780,N_17686,N_16217);
xor U24781 (N_24781,N_15036,N_18919);
xor U24782 (N_24782,N_19461,N_16909);
or U24783 (N_24783,N_15661,N_19815);
nor U24784 (N_24784,N_18847,N_17355);
xor U24785 (N_24785,N_16500,N_17446);
and U24786 (N_24786,N_19417,N_19695);
and U24787 (N_24787,N_19790,N_18822);
or U24788 (N_24788,N_15614,N_16231);
xnor U24789 (N_24789,N_18100,N_15452);
nor U24790 (N_24790,N_17258,N_16444);
nand U24791 (N_24791,N_17335,N_15159);
or U24792 (N_24792,N_19668,N_15967);
and U24793 (N_24793,N_15513,N_17765);
and U24794 (N_24794,N_19303,N_18638);
or U24795 (N_24795,N_17581,N_18132);
xnor U24796 (N_24796,N_17130,N_16295);
nor U24797 (N_24797,N_19167,N_15989);
nor U24798 (N_24798,N_18413,N_18294);
nand U24799 (N_24799,N_16806,N_17849);
xor U24800 (N_24800,N_19489,N_18233);
xnor U24801 (N_24801,N_16491,N_15549);
or U24802 (N_24802,N_19355,N_19064);
nor U24803 (N_24803,N_19499,N_17496);
xnor U24804 (N_24804,N_19882,N_17208);
xor U24805 (N_24805,N_17442,N_18829);
or U24806 (N_24806,N_17888,N_18796);
nand U24807 (N_24807,N_18459,N_17335);
nor U24808 (N_24808,N_16575,N_17608);
nor U24809 (N_24809,N_15348,N_19602);
nand U24810 (N_24810,N_19805,N_16367);
nand U24811 (N_24811,N_15662,N_19886);
nor U24812 (N_24812,N_19361,N_15069);
nand U24813 (N_24813,N_18100,N_17091);
or U24814 (N_24814,N_19983,N_17550);
xor U24815 (N_24815,N_17393,N_16941);
or U24816 (N_24816,N_18277,N_15551);
and U24817 (N_24817,N_15375,N_16814);
or U24818 (N_24818,N_19114,N_19780);
nand U24819 (N_24819,N_17554,N_18916);
xnor U24820 (N_24820,N_18662,N_16985);
or U24821 (N_24821,N_15031,N_18806);
nor U24822 (N_24822,N_17958,N_18692);
nor U24823 (N_24823,N_18115,N_17654);
xnor U24824 (N_24824,N_15990,N_16717);
and U24825 (N_24825,N_17890,N_19914);
and U24826 (N_24826,N_19148,N_15749);
or U24827 (N_24827,N_18348,N_18747);
xnor U24828 (N_24828,N_19839,N_16786);
xor U24829 (N_24829,N_17547,N_19071);
xor U24830 (N_24830,N_16201,N_17856);
xnor U24831 (N_24831,N_16902,N_17497);
xor U24832 (N_24832,N_16639,N_18451);
and U24833 (N_24833,N_18605,N_17503);
nand U24834 (N_24834,N_17948,N_17517);
or U24835 (N_24835,N_17183,N_19808);
or U24836 (N_24836,N_19921,N_17436);
xor U24837 (N_24837,N_15378,N_15237);
or U24838 (N_24838,N_16819,N_18557);
and U24839 (N_24839,N_16246,N_18497);
nand U24840 (N_24840,N_16438,N_15612);
xor U24841 (N_24841,N_19734,N_18025);
nand U24842 (N_24842,N_16272,N_15378);
or U24843 (N_24843,N_18085,N_18120);
xor U24844 (N_24844,N_15820,N_17271);
and U24845 (N_24845,N_18708,N_18541);
nor U24846 (N_24846,N_16618,N_15783);
nor U24847 (N_24847,N_17323,N_17796);
nand U24848 (N_24848,N_19722,N_18153);
nand U24849 (N_24849,N_19726,N_16608);
nor U24850 (N_24850,N_17936,N_16832);
and U24851 (N_24851,N_18638,N_19517);
or U24852 (N_24852,N_15113,N_16565);
nor U24853 (N_24853,N_19692,N_17000);
xor U24854 (N_24854,N_18304,N_17191);
or U24855 (N_24855,N_16810,N_17868);
nor U24856 (N_24856,N_18469,N_15853);
nor U24857 (N_24857,N_16257,N_17838);
xor U24858 (N_24858,N_17939,N_19879);
nor U24859 (N_24859,N_16817,N_15708);
or U24860 (N_24860,N_18809,N_19601);
nor U24861 (N_24861,N_16108,N_16404);
and U24862 (N_24862,N_18773,N_15474);
or U24863 (N_24863,N_16497,N_15508);
nand U24864 (N_24864,N_16758,N_17939);
xnor U24865 (N_24865,N_15046,N_15688);
xnor U24866 (N_24866,N_18901,N_18577);
nand U24867 (N_24867,N_16095,N_17567);
nor U24868 (N_24868,N_19068,N_15114);
xor U24869 (N_24869,N_18031,N_16341);
nand U24870 (N_24870,N_16971,N_19572);
or U24871 (N_24871,N_15778,N_19253);
nand U24872 (N_24872,N_17528,N_19822);
nand U24873 (N_24873,N_16624,N_17198);
nor U24874 (N_24874,N_16781,N_18620);
nand U24875 (N_24875,N_16421,N_17702);
and U24876 (N_24876,N_17757,N_17447);
nor U24877 (N_24877,N_17381,N_17494);
and U24878 (N_24878,N_16608,N_15216);
nand U24879 (N_24879,N_18499,N_15414);
xnor U24880 (N_24880,N_19506,N_15347);
xnor U24881 (N_24881,N_15989,N_16163);
nor U24882 (N_24882,N_15868,N_19454);
nor U24883 (N_24883,N_16275,N_18965);
or U24884 (N_24884,N_15948,N_18965);
nand U24885 (N_24885,N_19734,N_18532);
xnor U24886 (N_24886,N_17782,N_19962);
xor U24887 (N_24887,N_19773,N_18816);
or U24888 (N_24888,N_18773,N_16240);
nand U24889 (N_24889,N_15633,N_19467);
xnor U24890 (N_24890,N_19521,N_17058);
nor U24891 (N_24891,N_17725,N_16047);
xor U24892 (N_24892,N_17688,N_18718);
xor U24893 (N_24893,N_18051,N_16169);
nand U24894 (N_24894,N_17885,N_19294);
and U24895 (N_24895,N_19024,N_16986);
or U24896 (N_24896,N_15878,N_17585);
xor U24897 (N_24897,N_18093,N_17086);
and U24898 (N_24898,N_17341,N_16988);
nor U24899 (N_24899,N_15963,N_18248);
xor U24900 (N_24900,N_15352,N_15312);
nor U24901 (N_24901,N_15767,N_17301);
or U24902 (N_24902,N_15226,N_15551);
or U24903 (N_24903,N_16199,N_16521);
nor U24904 (N_24904,N_16845,N_16366);
nor U24905 (N_24905,N_18563,N_19216);
xor U24906 (N_24906,N_16027,N_15257);
nor U24907 (N_24907,N_18382,N_15731);
or U24908 (N_24908,N_18043,N_18571);
nand U24909 (N_24909,N_17074,N_19931);
nand U24910 (N_24910,N_19864,N_18101);
nor U24911 (N_24911,N_15040,N_19342);
nor U24912 (N_24912,N_15632,N_17717);
nor U24913 (N_24913,N_17190,N_16035);
or U24914 (N_24914,N_16329,N_19111);
nor U24915 (N_24915,N_17474,N_18145);
nor U24916 (N_24916,N_16143,N_16910);
xor U24917 (N_24917,N_15929,N_15746);
nor U24918 (N_24918,N_19909,N_18695);
nand U24919 (N_24919,N_19006,N_18128);
or U24920 (N_24920,N_17028,N_17475);
nand U24921 (N_24921,N_18885,N_16278);
nor U24922 (N_24922,N_16765,N_17701);
xnor U24923 (N_24923,N_18418,N_18639);
and U24924 (N_24924,N_15127,N_17628);
nand U24925 (N_24925,N_17458,N_15526);
or U24926 (N_24926,N_18348,N_15308);
nand U24927 (N_24927,N_15769,N_15737);
xor U24928 (N_24928,N_15775,N_15502);
nor U24929 (N_24929,N_17810,N_15524);
or U24930 (N_24930,N_18697,N_18187);
and U24931 (N_24931,N_15864,N_15563);
nor U24932 (N_24932,N_16297,N_19776);
or U24933 (N_24933,N_18291,N_19337);
or U24934 (N_24934,N_16231,N_18641);
nand U24935 (N_24935,N_18590,N_17153);
xor U24936 (N_24936,N_15060,N_19051);
and U24937 (N_24937,N_18698,N_16645);
or U24938 (N_24938,N_16572,N_17343);
xor U24939 (N_24939,N_18267,N_17832);
nand U24940 (N_24940,N_17378,N_18766);
and U24941 (N_24941,N_15255,N_19451);
nor U24942 (N_24942,N_17070,N_17151);
and U24943 (N_24943,N_17376,N_15823);
nand U24944 (N_24944,N_19575,N_16565);
nand U24945 (N_24945,N_15930,N_16236);
and U24946 (N_24946,N_19872,N_19720);
or U24947 (N_24947,N_16303,N_18569);
nand U24948 (N_24948,N_16092,N_19074);
nor U24949 (N_24949,N_16170,N_15392);
xnor U24950 (N_24950,N_15764,N_18595);
or U24951 (N_24951,N_19850,N_15032);
and U24952 (N_24952,N_16957,N_19733);
nand U24953 (N_24953,N_18622,N_16317);
nor U24954 (N_24954,N_16313,N_18795);
and U24955 (N_24955,N_17163,N_18613);
and U24956 (N_24956,N_19840,N_17371);
nor U24957 (N_24957,N_19931,N_16665);
nor U24958 (N_24958,N_16120,N_19756);
xnor U24959 (N_24959,N_15569,N_18020);
and U24960 (N_24960,N_16625,N_18247);
or U24961 (N_24961,N_15187,N_18103);
or U24962 (N_24962,N_18792,N_15695);
nand U24963 (N_24963,N_18055,N_19782);
xor U24964 (N_24964,N_18101,N_15518);
and U24965 (N_24965,N_18862,N_15678);
nor U24966 (N_24966,N_18288,N_15213);
or U24967 (N_24967,N_15839,N_19245);
xor U24968 (N_24968,N_18649,N_16950);
and U24969 (N_24969,N_18673,N_19618);
nor U24970 (N_24970,N_17425,N_16823);
xnor U24971 (N_24971,N_18738,N_18207);
or U24972 (N_24972,N_19214,N_15943);
xnor U24973 (N_24973,N_15978,N_16962);
xor U24974 (N_24974,N_17635,N_19491);
nor U24975 (N_24975,N_18045,N_18819);
nand U24976 (N_24976,N_18392,N_17393);
nand U24977 (N_24977,N_15387,N_16998);
or U24978 (N_24978,N_19901,N_16145);
nand U24979 (N_24979,N_17105,N_15918);
or U24980 (N_24980,N_18992,N_18073);
xor U24981 (N_24981,N_17482,N_17121);
xnor U24982 (N_24982,N_17139,N_18334);
or U24983 (N_24983,N_17687,N_18912);
xor U24984 (N_24984,N_15638,N_17569);
nand U24985 (N_24985,N_15839,N_18431);
or U24986 (N_24986,N_19572,N_15684);
xor U24987 (N_24987,N_16191,N_17344);
and U24988 (N_24988,N_19992,N_16250);
nand U24989 (N_24989,N_18843,N_16789);
xnor U24990 (N_24990,N_19582,N_17083);
and U24991 (N_24991,N_19912,N_17442);
xnor U24992 (N_24992,N_19185,N_15978);
nor U24993 (N_24993,N_17422,N_16358);
and U24994 (N_24994,N_17462,N_16796);
and U24995 (N_24995,N_17547,N_19996);
nor U24996 (N_24996,N_18028,N_18801);
xor U24997 (N_24997,N_19421,N_17203);
xor U24998 (N_24998,N_17958,N_15083);
nor U24999 (N_24999,N_19358,N_19180);
and UO_0 (O_0,N_22621,N_20007);
nor UO_1 (O_1,N_21920,N_22435);
or UO_2 (O_2,N_23170,N_23985);
nor UO_3 (O_3,N_20729,N_22750);
or UO_4 (O_4,N_23878,N_23447);
nand UO_5 (O_5,N_21830,N_23461);
nand UO_6 (O_6,N_24408,N_20706);
or UO_7 (O_7,N_24586,N_20659);
nand UO_8 (O_8,N_24920,N_22143);
and UO_9 (O_9,N_23250,N_21321);
nand UO_10 (O_10,N_24971,N_24674);
xnor UO_11 (O_11,N_22480,N_23981);
xnor UO_12 (O_12,N_22815,N_20159);
xnor UO_13 (O_13,N_23820,N_20409);
xor UO_14 (O_14,N_24344,N_21685);
or UO_15 (O_15,N_23754,N_22687);
nor UO_16 (O_16,N_22700,N_21174);
nor UO_17 (O_17,N_21940,N_21840);
nor UO_18 (O_18,N_21262,N_20910);
nand UO_19 (O_19,N_23464,N_20320);
nand UO_20 (O_20,N_21370,N_23612);
nand UO_21 (O_21,N_24595,N_21513);
and UO_22 (O_22,N_21154,N_24613);
or UO_23 (O_23,N_21866,N_24139);
nand UO_24 (O_24,N_24689,N_21613);
or UO_25 (O_25,N_23951,N_22804);
nand UO_26 (O_26,N_21228,N_24457);
and UO_27 (O_27,N_23284,N_23535);
and UO_28 (O_28,N_24077,N_24751);
xnor UO_29 (O_29,N_23716,N_23563);
nand UO_30 (O_30,N_21883,N_21646);
xor UO_31 (O_31,N_24225,N_21650);
or UO_32 (O_32,N_23101,N_20448);
and UO_33 (O_33,N_23694,N_24668);
xor UO_34 (O_34,N_23979,N_20335);
xor UO_35 (O_35,N_22604,N_22842);
and UO_36 (O_36,N_21582,N_22832);
nand UO_37 (O_37,N_23720,N_21778);
nand UO_38 (O_38,N_22839,N_20165);
or UO_39 (O_39,N_21602,N_24086);
nor UO_40 (O_40,N_21418,N_22572);
xnor UO_41 (O_41,N_20677,N_24900);
xnor UO_42 (O_42,N_22388,N_23301);
or UO_43 (O_43,N_24443,N_22860);
and UO_44 (O_44,N_23248,N_20507);
xor UO_45 (O_45,N_23160,N_24795);
and UO_46 (O_46,N_22620,N_20904);
or UO_47 (O_47,N_21201,N_22884);
xor UO_48 (O_48,N_23877,N_20351);
xnor UO_49 (O_49,N_20106,N_22879);
nand UO_50 (O_50,N_22564,N_24211);
xnor UO_51 (O_51,N_21786,N_24445);
or UO_52 (O_52,N_22780,N_24279);
or UO_53 (O_53,N_24927,N_23778);
or UO_54 (O_54,N_22182,N_22729);
nor UO_55 (O_55,N_21546,N_21320);
or UO_56 (O_56,N_24415,N_20275);
or UO_57 (O_57,N_24154,N_22658);
and UO_58 (O_58,N_20424,N_23347);
and UO_59 (O_59,N_22920,N_23448);
nand UO_60 (O_60,N_20143,N_20151);
or UO_61 (O_61,N_23411,N_23588);
nand UO_62 (O_62,N_20136,N_20191);
or UO_63 (O_63,N_21748,N_22481);
or UO_64 (O_64,N_22918,N_21294);
or UO_65 (O_65,N_22693,N_21302);
nand UO_66 (O_66,N_20011,N_22991);
nand UO_67 (O_67,N_24057,N_24039);
or UO_68 (O_68,N_20917,N_24126);
nor UO_69 (O_69,N_21383,N_20887);
xnor UO_70 (O_70,N_23927,N_23709);
xor UO_71 (O_71,N_20988,N_22233);
xnor UO_72 (O_72,N_22706,N_23683);
nor UO_73 (O_73,N_24204,N_23221);
nand UO_74 (O_74,N_24367,N_23199);
nand UO_75 (O_75,N_23868,N_22649);
nor UO_76 (O_76,N_20393,N_22033);
and UO_77 (O_77,N_21117,N_22577);
and UO_78 (O_78,N_22513,N_24609);
or UO_79 (O_79,N_20480,N_23648);
nand UO_80 (O_80,N_21015,N_22710);
xnor UO_81 (O_81,N_21637,N_21177);
nor UO_82 (O_82,N_21738,N_20438);
or UO_83 (O_83,N_22160,N_21851);
nand UO_84 (O_84,N_22339,N_22640);
nor UO_85 (O_85,N_24269,N_21491);
xor UO_86 (O_86,N_20337,N_21335);
and UO_87 (O_87,N_20831,N_21547);
xnor UO_88 (O_88,N_24250,N_24160);
and UO_89 (O_89,N_24429,N_21436);
or UO_90 (O_90,N_21938,N_20786);
nor UO_91 (O_91,N_20864,N_24635);
or UO_92 (O_92,N_20058,N_20533);
nand UO_93 (O_93,N_22323,N_23278);
nand UO_94 (O_94,N_20180,N_22811);
nor UO_95 (O_95,N_20052,N_23850);
nand UO_96 (O_96,N_23399,N_20281);
and UO_97 (O_97,N_20352,N_24738);
and UO_98 (O_98,N_20400,N_21087);
xor UO_99 (O_99,N_22568,N_22281);
xnor UO_100 (O_100,N_22555,N_23035);
and UO_101 (O_101,N_21809,N_21314);
nor UO_102 (O_102,N_22179,N_20751);
nand UO_103 (O_103,N_24376,N_23687);
and UO_104 (O_104,N_24251,N_20856);
nand UO_105 (O_105,N_21681,N_23750);
nand UO_106 (O_106,N_23988,N_22028);
xor UO_107 (O_107,N_24911,N_22615);
and UO_108 (O_108,N_21397,N_20416);
nor UO_109 (O_109,N_21250,N_22950);
and UO_110 (O_110,N_20031,N_22643);
nand UO_111 (O_111,N_24934,N_20763);
nand UO_112 (O_112,N_21910,N_22704);
nor UO_113 (O_113,N_23311,N_21743);
nor UO_114 (O_114,N_22016,N_23274);
nor UO_115 (O_115,N_22847,N_23304);
and UO_116 (O_116,N_23204,N_21163);
xor UO_117 (O_117,N_20899,N_21790);
nand UO_118 (O_118,N_24991,N_21726);
nand UO_119 (O_119,N_22773,N_21407);
and UO_120 (O_120,N_23320,N_23344);
nor UO_121 (O_121,N_20894,N_21917);
nor UO_122 (O_122,N_22347,N_23832);
or UO_123 (O_123,N_23336,N_24285);
nand UO_124 (O_124,N_21247,N_20370);
and UO_125 (O_125,N_24132,N_20877);
nor UO_126 (O_126,N_22512,N_22042);
and UO_127 (O_127,N_20230,N_22807);
nor UO_128 (O_128,N_20002,N_23355);
nor UO_129 (O_129,N_24584,N_24485);
nand UO_130 (O_130,N_21297,N_24277);
xnor UO_131 (O_131,N_22696,N_22414);
xor UO_132 (O_132,N_22048,N_21414);
nor UO_133 (O_133,N_21924,N_21212);
nor UO_134 (O_134,N_20360,N_22352);
nand UO_135 (O_135,N_20966,N_23911);
nor UO_136 (O_136,N_20436,N_23615);
nor UO_137 (O_137,N_23073,N_24284);
and UO_138 (O_138,N_21811,N_20692);
or UO_139 (O_139,N_21927,N_20719);
nand UO_140 (O_140,N_21240,N_22427);
and UO_141 (O_141,N_24929,N_20934);
nor UO_142 (O_142,N_21708,N_21588);
or UO_143 (O_143,N_21426,N_23958);
xor UO_144 (O_144,N_24133,N_21019);
xnor UO_145 (O_145,N_22191,N_22025);
xnor UO_146 (O_146,N_24252,N_23982);
nor UO_147 (O_147,N_23689,N_22765);
and UO_148 (O_148,N_20848,N_21120);
xnor UO_149 (O_149,N_21324,N_20774);
nand UO_150 (O_150,N_24603,N_21279);
and UO_151 (O_151,N_22008,N_24538);
nand UO_152 (O_152,N_20477,N_24757);
xnor UO_153 (O_153,N_24159,N_24213);
xnor UO_154 (O_154,N_23459,N_23150);
nand UO_155 (O_155,N_21260,N_24474);
xor UO_156 (O_156,N_23509,N_21025);
nand UO_157 (O_157,N_20100,N_22736);
and UO_158 (O_158,N_21231,N_20560);
nor UO_159 (O_159,N_20341,N_21978);
nand UO_160 (O_160,N_22968,N_21821);
nor UO_161 (O_161,N_22258,N_24069);
xor UO_162 (O_162,N_20897,N_24137);
xor UO_163 (O_163,N_23295,N_24106);
nor UO_164 (O_164,N_21275,N_23132);
and UO_165 (O_165,N_20549,N_24064);
nor UO_166 (O_166,N_20649,N_24328);
xor UO_167 (O_167,N_22456,N_24688);
or UO_168 (O_168,N_23436,N_21104);
nor UO_169 (O_169,N_21594,N_22189);
nand UO_170 (O_170,N_23650,N_21179);
nand UO_171 (O_171,N_23708,N_20911);
nand UO_172 (O_172,N_24628,N_21700);
or UO_173 (O_173,N_22669,N_24056);
nand UO_174 (O_174,N_22557,N_22911);
nand UO_175 (O_175,N_23034,N_23884);
nand UO_176 (O_176,N_20661,N_23993);
nand UO_177 (O_177,N_21736,N_20483);
or UO_178 (O_178,N_24568,N_24964);
nor UO_179 (O_179,N_20529,N_22685);
and UO_180 (O_180,N_20329,N_21099);
nand UO_181 (O_181,N_20365,N_20821);
nor UO_182 (O_182,N_23042,N_24536);
nand UO_183 (O_183,N_21661,N_21621);
xnor UO_184 (O_184,N_23256,N_24483);
nor UO_185 (O_185,N_24599,N_23460);
xnor UO_186 (O_186,N_23539,N_20739);
xor UO_187 (O_187,N_24303,N_23423);
and UO_188 (O_188,N_24870,N_23133);
nand UO_189 (O_189,N_24343,N_20025);
xnor UO_190 (O_190,N_23241,N_23099);
xnor UO_191 (O_191,N_22146,N_24841);
and UO_192 (O_192,N_20050,N_21574);
or UO_193 (O_193,N_23536,N_24111);
xor UO_194 (O_194,N_22275,N_20812);
nor UO_195 (O_195,N_20891,N_23482);
nand UO_196 (O_196,N_22056,N_23743);
nor UO_197 (O_197,N_21719,N_24007);
nand UO_198 (O_198,N_21632,N_20747);
or UO_199 (O_199,N_23242,N_21333);
and UO_200 (O_200,N_21007,N_24878);
xor UO_201 (O_201,N_20594,N_20305);
and UO_202 (O_202,N_23939,N_20947);
or UO_203 (O_203,N_23404,N_24329);
and UO_204 (O_204,N_23571,N_23548);
nor UO_205 (O_205,N_24661,N_22442);
or UO_206 (O_206,N_23790,N_24230);
nor UO_207 (O_207,N_20294,N_22045);
nor UO_208 (O_208,N_21276,N_20839);
nand UO_209 (O_209,N_20285,N_23151);
nand UO_210 (O_210,N_22924,N_21001);
xnor UO_211 (O_211,N_23185,N_24606);
and UO_212 (O_212,N_23007,N_20907);
nor UO_213 (O_213,N_21592,N_20005);
and UO_214 (O_214,N_21605,N_22629);
xnor UO_215 (O_215,N_20873,N_23352);
nand UO_216 (O_216,N_24995,N_21325);
nand UO_217 (O_217,N_22126,N_24905);
nor UO_218 (O_218,N_22495,N_23814);
xor UO_219 (O_219,N_20761,N_20123);
nor UO_220 (O_220,N_22415,N_24610);
xor UO_221 (O_221,N_23564,N_23283);
or UO_222 (O_222,N_20272,N_21593);
nand UO_223 (O_223,N_20362,N_24566);
nand UO_224 (O_224,N_21095,N_22366);
or UO_225 (O_225,N_23593,N_20000);
nand UO_226 (O_226,N_23033,N_20663);
nand UO_227 (O_227,N_24850,N_24231);
or UO_228 (O_228,N_20250,N_21429);
nand UO_229 (O_229,N_21941,N_23469);
or UO_230 (O_230,N_21449,N_22148);
nor UO_231 (O_231,N_22491,N_22128);
or UO_232 (O_232,N_24877,N_23236);
nor UO_233 (O_233,N_22987,N_21517);
xor UO_234 (O_234,N_20942,N_21774);
or UO_235 (O_235,N_20652,N_20845);
nor UO_236 (O_236,N_23124,N_20767);
nor UO_237 (O_237,N_24600,N_22406);
and UO_238 (O_238,N_22936,N_24021);
nand UO_239 (O_239,N_21717,N_20261);
nand UO_240 (O_240,N_20263,N_22834);
xor UO_241 (O_241,N_20323,N_20038);
nor UO_242 (O_242,N_21455,N_20183);
xnor UO_243 (O_243,N_20772,N_23675);
xnor UO_244 (O_244,N_23153,N_20125);
and UO_245 (O_245,N_20941,N_24540);
and UO_246 (O_246,N_22838,N_23439);
and UO_247 (O_247,N_20737,N_21504);
xnor UO_248 (O_248,N_20114,N_21051);
and UO_249 (O_249,N_20017,N_22975);
nor UO_250 (O_250,N_23126,N_21986);
nor UO_251 (O_251,N_21796,N_22720);
and UO_252 (O_252,N_23489,N_22945);
and UO_253 (O_253,N_22411,N_23656);
and UO_254 (O_254,N_24270,N_22170);
and UO_255 (O_255,N_21939,N_20334);
nand UO_256 (O_256,N_21295,N_20890);
nand UO_257 (O_257,N_21244,N_22398);
nand UO_258 (O_258,N_24008,N_22458);
nand UO_259 (O_259,N_20307,N_24531);
and UO_260 (O_260,N_22799,N_24105);
and UO_261 (O_261,N_22686,N_20544);
and UO_262 (O_262,N_22993,N_20475);
and UO_263 (O_263,N_23975,N_23473);
or UO_264 (O_264,N_24374,N_22180);
or UO_265 (O_265,N_20063,N_23051);
and UO_266 (O_266,N_22965,N_20804);
and UO_267 (O_267,N_20141,N_22650);
nor UO_268 (O_268,N_22881,N_22068);
nand UO_269 (O_269,N_21897,N_21447);
xnor UO_270 (O_270,N_20805,N_24027);
or UO_271 (O_271,N_22098,N_20656);
or UO_272 (O_272,N_20963,N_20803);
xnor UO_273 (O_273,N_24484,N_22348);
nor UO_274 (O_274,N_24972,N_22797);
nand UO_275 (O_275,N_22006,N_21690);
nand UO_276 (O_276,N_21783,N_23553);
nand UO_277 (O_277,N_21222,N_21848);
xor UO_278 (O_278,N_23599,N_20177);
nor UO_279 (O_279,N_20749,N_24138);
nor UO_280 (O_280,N_22484,N_23961);
nor UO_281 (O_281,N_24217,N_24977);
or UO_282 (O_282,N_24572,N_22431);
nor UO_283 (O_283,N_24393,N_21711);
or UO_284 (O_284,N_21289,N_23314);
xnor UO_285 (O_285,N_20004,N_22913);
nand UO_286 (O_286,N_21740,N_20233);
xor UO_287 (O_287,N_23560,N_20255);
xnor UO_288 (O_288,N_23235,N_23377);
nor UO_289 (O_289,N_20733,N_21996);
or UO_290 (O_290,N_22377,N_21310);
and UO_291 (O_291,N_22266,N_22074);
nand UO_292 (O_292,N_22009,N_21094);
xnor UO_293 (O_293,N_20931,N_23766);
or UO_294 (O_294,N_20008,N_22494);
nand UO_295 (O_295,N_24897,N_23366);
nand UO_296 (O_296,N_21864,N_23521);
or UO_297 (O_297,N_20811,N_24395);
nand UO_298 (O_298,N_23063,N_20976);
nor UO_299 (O_299,N_22997,N_21384);
nor UO_300 (O_300,N_23938,N_23629);
or UO_301 (O_301,N_21286,N_23259);
nand UO_302 (O_302,N_21387,N_24409);
and UO_303 (O_303,N_23614,N_20016);
or UO_304 (O_304,N_21727,N_22312);
xor UO_305 (O_305,N_21326,N_24206);
and UO_306 (O_306,N_23512,N_23086);
nor UO_307 (O_307,N_20762,N_21911);
or UO_308 (O_308,N_23357,N_20073);
and UO_309 (O_309,N_23093,N_22461);
nand UO_310 (O_310,N_20492,N_23880);
or UO_311 (O_311,N_24241,N_21899);
xnor UO_312 (O_312,N_24083,N_23807);
xnor UO_313 (O_313,N_20155,N_20420);
and UO_314 (O_314,N_24922,N_23004);
nor UO_315 (O_315,N_21338,N_24079);
xor UO_316 (O_316,N_24300,N_24493);
and UO_317 (O_317,N_24994,N_22558);
nand UO_318 (O_318,N_23704,N_24559);
nand UO_319 (O_319,N_23001,N_24743);
or UO_320 (O_320,N_23984,N_23742);
nand UO_321 (O_321,N_22344,N_24831);
xor UO_322 (O_322,N_20632,N_23827);
xnor UO_323 (O_323,N_20883,N_22283);
or UO_324 (O_324,N_23410,N_23928);
nor UO_325 (O_325,N_23478,N_20810);
nor UO_326 (O_326,N_23853,N_22420);
nand UO_327 (O_327,N_24107,N_22395);
or UO_328 (O_328,N_24098,N_24044);
nand UO_329 (O_329,N_24084,N_20216);
nor UO_330 (O_330,N_24399,N_20522);
or UO_331 (O_331,N_21113,N_22066);
nand UO_332 (O_332,N_23739,N_24459);
nor UO_333 (O_333,N_20595,N_24716);
or UO_334 (O_334,N_21600,N_24936);
nor UO_335 (O_335,N_20527,N_22809);
xnor UO_336 (O_336,N_24685,N_20296);
xnor UO_337 (O_337,N_21766,N_23251);
xor UO_338 (O_338,N_21890,N_23607);
and UO_339 (O_339,N_21011,N_20566);
and UO_340 (O_340,N_23503,N_22294);
or UO_341 (O_341,N_23799,N_20641);
nand UO_342 (O_342,N_20313,N_24188);
nor UO_343 (O_343,N_24565,N_23806);
xnor UO_344 (O_344,N_20037,N_21606);
xnor UO_345 (O_345,N_22562,N_23379);
or UO_346 (O_346,N_23918,N_21017);
nand UO_347 (O_347,N_22758,N_21686);
xnor UO_348 (O_348,N_21577,N_23608);
nor UO_349 (O_349,N_23657,N_24941);
xnor UO_350 (O_350,N_20056,N_20071);
nand UO_351 (O_351,N_23679,N_22313);
and UO_352 (O_352,N_22806,N_23934);
or UO_353 (O_353,N_20431,N_22752);
or UO_354 (O_354,N_21521,N_20557);
nor UO_355 (O_355,N_23498,N_24145);
or UO_356 (O_356,N_23839,N_20870);
or UO_357 (O_357,N_20363,N_23030);
or UO_358 (O_358,N_23430,N_24271);
nor UO_359 (O_359,N_22738,N_23723);
nand UO_360 (O_360,N_24460,N_20920);
xor UO_361 (O_361,N_21202,N_20771);
and UO_362 (O_362,N_23195,N_23722);
nand UO_363 (O_363,N_22209,N_22775);
or UO_364 (O_364,N_23135,N_24744);
nand UO_365 (O_365,N_22959,N_21443);
xnor UO_366 (O_366,N_22144,N_20430);
and UO_367 (O_367,N_23525,N_20510);
or UO_368 (O_368,N_20271,N_23475);
xor UO_369 (O_369,N_21124,N_20955);
nand UO_370 (O_370,N_24428,N_23176);
nor UO_371 (O_371,N_22177,N_24530);
or UO_372 (O_372,N_24156,N_20655);
nor UO_373 (O_373,N_20587,N_21208);
and UO_374 (O_374,N_22289,N_23788);
xor UO_375 (O_375,N_21266,N_23289);
nor UO_376 (O_376,N_24742,N_24551);
xnor UO_377 (O_377,N_21846,N_20978);
nor UO_378 (O_378,N_21770,N_21027);
xor UO_379 (O_379,N_23025,N_24434);
and UO_380 (O_380,N_22267,N_24984);
xnor UO_381 (O_381,N_24239,N_24490);
nor UO_382 (O_382,N_21501,N_21858);
xor UO_383 (O_383,N_24946,N_20109);
or UO_384 (O_384,N_22387,N_24268);
xor UO_385 (O_385,N_20023,N_22488);
xnor UO_386 (O_386,N_23881,N_23193);
nand UO_387 (O_387,N_22535,N_23692);
or UO_388 (O_388,N_20836,N_22631);
nand UO_389 (O_389,N_23089,N_20412);
or UO_390 (O_390,N_21049,N_22723);
nand UO_391 (O_391,N_23517,N_21789);
and UO_392 (O_392,N_24967,N_21833);
nor UO_393 (O_393,N_21351,N_22567);
xnor UO_394 (O_394,N_24807,N_22024);
and UO_395 (O_395,N_23332,N_21272);
nor UO_396 (O_396,N_20376,N_23960);
nor UO_397 (O_397,N_23661,N_23168);
nor UO_398 (O_398,N_24410,N_20354);
nor UO_399 (O_399,N_24371,N_22173);
xor UO_400 (O_400,N_21900,N_21567);
nor UO_401 (O_401,N_20019,N_23189);
nand UO_402 (O_402,N_23831,N_24604);
xor UO_403 (O_403,N_21510,N_24558);
xnor UO_404 (O_404,N_21614,N_23978);
xor UO_405 (O_405,N_24855,N_24687);
xnor UO_406 (O_406,N_20375,N_22376);
nor UO_407 (O_407,N_21963,N_22777);
xnor UO_408 (O_408,N_21536,N_23758);
and UO_409 (O_409,N_23600,N_24837);
or UO_410 (O_410,N_22211,N_20265);
xnor UO_411 (O_411,N_24264,N_23292);
nor UO_412 (O_412,N_22976,N_21946);
nor UO_413 (O_413,N_24914,N_24337);
and UO_414 (O_414,N_23549,N_21398);
xor UO_415 (O_415,N_20218,N_20918);
xnor UO_416 (O_416,N_24533,N_22930);
nor UO_417 (O_417,N_24049,N_20342);
nor UO_418 (O_418,N_22953,N_22482);
nor UO_419 (O_419,N_21009,N_20757);
and UO_420 (O_420,N_20417,N_24793);
xor UO_421 (O_421,N_20163,N_20040);
nor UO_422 (O_422,N_23625,N_22988);
nand UO_423 (O_423,N_24745,N_20078);
xnor UO_424 (O_424,N_21780,N_22836);
and UO_425 (O_425,N_22787,N_22525);
nor UO_426 (O_426,N_22971,N_23695);
and UO_427 (O_427,N_20208,N_21581);
nor UO_428 (O_428,N_21529,N_22537);
nand UO_429 (O_429,N_22759,N_24073);
xnor UO_430 (O_430,N_22397,N_22730);
nand UO_431 (O_431,N_20054,N_24425);
nand UO_432 (O_432,N_22129,N_20032);
nor UO_433 (O_433,N_22707,N_20173);
nand UO_434 (O_434,N_21016,N_21428);
and UO_435 (O_435,N_23010,N_22600);
nor UO_436 (O_436,N_24127,N_21484);
xor UO_437 (O_437,N_22138,N_22162);
and UO_438 (O_438,N_22751,N_20539);
or UO_439 (O_439,N_21578,N_21166);
or UO_440 (O_440,N_22372,N_21216);
nand UO_441 (O_441,N_22588,N_21149);
or UO_442 (O_442,N_24338,N_20833);
nor UO_443 (O_443,N_23462,N_24771);
nand UO_444 (O_444,N_21182,N_21097);
nor UO_445 (O_445,N_22301,N_22824);
xor UO_446 (O_446,N_21061,N_20224);
xnor UO_447 (O_447,N_20716,N_21550);
nor UO_448 (O_448,N_22746,N_23871);
nor UO_449 (O_449,N_21256,N_23944);
nor UO_450 (O_450,N_22589,N_24261);
and UO_451 (O_451,N_22770,N_20532);
or UO_452 (O_452,N_24085,N_21926);
or UO_453 (O_453,N_20860,N_21775);
nor UO_454 (O_454,N_20080,N_23577);
nor UO_455 (O_455,N_23119,N_24403);
nor UO_456 (O_456,N_21887,N_22188);
xor UO_457 (O_457,N_22900,N_21071);
xnor UO_458 (O_458,N_23114,N_23729);
or UO_459 (O_459,N_24396,N_21080);
nand UO_460 (O_460,N_22592,N_24889);
or UO_461 (O_461,N_24433,N_22114);
nor UO_462 (O_462,N_22212,N_21048);
and UO_463 (O_463,N_20473,N_22743);
or UO_464 (O_464,N_20267,N_21267);
nor UO_465 (O_465,N_22876,N_22390);
or UO_466 (O_466,N_24809,N_20443);
and UO_467 (O_467,N_24622,N_24117);
or UO_468 (O_468,N_24525,N_23203);
nand UO_469 (O_469,N_22329,N_22220);
xor UO_470 (O_470,N_20404,N_24605);
xnor UO_471 (O_471,N_24895,N_20482);
nor UO_472 (O_472,N_20053,N_20620);
nor UO_473 (O_473,N_21424,N_21710);
and UO_474 (O_474,N_23717,N_21677);
nor UO_475 (O_475,N_20730,N_23309);
or UO_476 (O_476,N_20189,N_21277);
nor UO_477 (O_477,N_22956,N_24948);
xor UO_478 (O_478,N_23935,N_24032);
xnor UO_479 (O_479,N_21597,N_20377);
or UO_480 (O_480,N_21507,N_20981);
nor UO_481 (O_481,N_24449,N_23817);
or UO_482 (O_482,N_20913,N_21406);
or UO_483 (O_483,N_20135,N_23245);
nand UO_484 (O_484,N_22697,N_23740);
or UO_485 (O_485,N_23865,N_22837);
or UO_486 (O_486,N_22053,N_21178);
nand UO_487 (O_487,N_20640,N_24013);
nor UO_488 (O_488,N_24259,N_21296);
nor UO_489 (O_489,N_21372,N_20682);
and UO_490 (O_490,N_22120,N_23415);
nand UO_491 (O_491,N_23899,N_22619);
or UO_492 (O_492,N_20432,N_20467);
and UO_493 (O_493,N_22576,N_24824);
nor UO_494 (O_494,N_24451,N_23217);
xnor UO_495 (O_495,N_20397,N_22291);
nor UO_496 (O_496,N_21872,N_21603);
nor UO_497 (O_497,N_20695,N_22475);
or UO_498 (O_498,N_22506,N_20210);
nand UO_499 (O_499,N_20014,N_21684);
xor UO_500 (O_500,N_23098,N_21865);
nand UO_501 (O_501,N_23169,N_20639);
and UO_502 (O_502,N_21667,N_24792);
and UO_503 (O_503,N_23127,N_24136);
nor UO_504 (O_504,N_21868,N_22087);
and UO_505 (O_505,N_22771,N_24509);
nor UO_506 (O_506,N_22928,N_24938);
or UO_507 (O_507,N_22460,N_21064);
xor UO_508 (O_508,N_20547,N_23940);
or UO_509 (O_509,N_21623,N_24177);
nor UO_510 (O_510,N_20914,N_20419);
nand UO_511 (O_511,N_22385,N_23414);
nor UO_512 (O_512,N_24869,N_21031);
nand UO_513 (O_513,N_21797,N_21674);
and UO_514 (O_514,N_23223,N_23578);
or UO_515 (O_515,N_22509,N_24790);
or UO_516 (O_516,N_20399,N_22310);
or UO_517 (O_517,N_23835,N_20555);
xor UO_518 (O_518,N_21959,N_20543);
and UO_519 (O_519,N_20124,N_24341);
xnor UO_520 (O_520,N_21634,N_20378);
and UO_521 (O_521,N_24149,N_22757);
xor UO_522 (O_522,N_21188,N_21850);
nand UO_523 (O_523,N_23520,N_21362);
nor UO_524 (O_524,N_22112,N_22216);
xnor UO_525 (O_525,N_20813,N_22904);
nand UO_526 (O_526,N_22019,N_22410);
nor UO_527 (O_527,N_21657,N_22280);
xnor UO_528 (O_528,N_20421,N_24621);
nor UO_529 (O_529,N_23392,N_24856);
nor UO_530 (O_530,N_24748,N_22614);
and UO_531 (O_531,N_23725,N_24390);
nor UO_532 (O_532,N_24947,N_22500);
and UO_533 (O_533,N_20201,N_23339);
or UO_534 (O_534,N_22812,N_22656);
nor UO_535 (O_535,N_21013,N_23942);
nand UO_536 (O_536,N_20708,N_22916);
xor UO_537 (O_537,N_20889,N_21672);
and UO_538 (O_538,N_20239,N_21288);
or UO_539 (O_539,N_22318,N_22311);
and UO_540 (O_540,N_21442,N_24335);
xnor UO_541 (O_541,N_21808,N_20277);
or UO_542 (O_542,N_21699,N_20946);
xor UO_543 (O_543,N_22864,N_22534);
and UO_544 (O_544,N_22337,N_21794);
or UO_545 (O_545,N_23895,N_24272);
nand UO_546 (O_546,N_23041,N_20886);
and UO_547 (O_547,N_21371,N_23644);
nand UO_548 (O_548,N_23646,N_21842);
and UO_549 (O_549,N_24081,N_23013);
or UO_550 (O_550,N_20010,N_23507);
xor UO_551 (O_551,N_23175,N_20170);
nor UO_552 (O_552,N_20447,N_24992);
or UO_553 (O_553,N_22116,N_21906);
nand UO_554 (O_554,N_20635,N_21722);
or UO_555 (O_555,N_20214,N_23308);
and UO_556 (O_556,N_21984,N_24293);
nand UO_557 (O_557,N_20030,N_21140);
and UO_558 (O_558,N_24851,N_24507);
or UO_559 (O_559,N_23121,N_21579);
xnor UO_560 (O_560,N_24707,N_23816);
nand UO_561 (O_561,N_24637,N_23523);
or UO_562 (O_562,N_22213,N_20735);
nand UO_563 (O_563,N_21885,N_24414);
xor UO_564 (O_564,N_22288,N_22067);
nand UO_565 (O_565,N_22873,N_20505);
nand UO_566 (O_566,N_21993,N_23047);
xor UO_567 (O_567,N_23580,N_20027);
xnor UO_568 (O_568,N_22073,N_22350);
and UO_569 (O_569,N_20121,N_24148);
and UO_570 (O_570,N_24496,N_22679);
xnor UO_571 (O_571,N_23201,N_24843);
nand UO_572 (O_572,N_21709,N_21194);
nor UO_573 (O_573,N_23313,N_24248);
nand UO_574 (O_574,N_20227,N_24351);
xor UO_575 (O_575,N_22268,N_22628);
nor UO_576 (O_576,N_20678,N_24113);
nor UO_577 (O_577,N_24253,N_22974);
xor UO_578 (O_578,N_21633,N_23952);
nor UO_579 (O_579,N_21213,N_20691);
xnor UO_580 (O_580,N_23470,N_21683);
and UO_581 (O_581,N_22441,N_22426);
and UO_582 (O_582,N_21664,N_21448);
nand UO_583 (O_583,N_22673,N_21209);
and UO_584 (O_584,N_20065,N_20160);
and UO_585 (O_585,N_21902,N_24491);
nand UO_586 (O_586,N_21891,N_21282);
nand UO_587 (O_587,N_21828,N_22662);
nor UO_588 (O_588,N_22552,N_23715);
and UO_589 (O_589,N_21423,N_21562);
xnor UO_590 (O_590,N_21160,N_23736);
nand UO_591 (O_591,N_20254,N_23394);
nor UO_592 (O_592,N_21367,N_21159);
xnor UO_593 (O_593,N_20336,N_23852);
nand UO_594 (O_594,N_23148,N_23882);
and UO_595 (O_595,N_22575,N_20386);
nor UO_596 (O_596,N_24278,N_24422);
xnor UO_597 (O_597,N_21107,N_21624);
xnor UO_598 (O_598,N_20321,N_24322);
nand UO_599 (O_599,N_24388,N_22020);
and UO_600 (O_600,N_23562,N_20605);
nor UO_601 (O_601,N_22915,N_21076);
and UO_602 (O_602,N_20696,N_20827);
nor UO_603 (O_603,N_24478,N_23872);
nor UO_604 (O_604,N_22470,N_24500);
or UO_605 (O_605,N_20454,N_23401);
and UO_606 (O_606,N_24960,N_22530);
xnor UO_607 (O_607,N_21759,N_20493);
or UO_608 (O_608,N_20583,N_22158);
xnor UO_609 (O_609,N_21217,N_22580);
xnor UO_610 (O_610,N_22413,N_20621);
xnor UO_611 (O_611,N_23325,N_22375);
and UO_612 (O_612,N_22651,N_22478);
and UO_613 (O_613,N_20815,N_24944);
nand UO_614 (O_614,N_23898,N_24072);
and UO_615 (O_615,N_21218,N_23212);
or UO_616 (O_616,N_24829,N_23690);
nand UO_617 (O_617,N_21524,N_23793);
xor UO_618 (O_618,N_21982,N_22247);
or UO_619 (O_619,N_21180,N_21976);
or UO_620 (O_620,N_24777,N_20959);
and UO_621 (O_621,N_21035,N_23340);
or UO_622 (O_622,N_21252,N_22051);
xor UO_623 (O_623,N_23487,N_23029);
xor UO_624 (O_624,N_24585,N_24140);
or UO_625 (O_625,N_23957,N_23810);
or UO_626 (O_626,N_24514,N_23365);
nor UO_627 (O_627,N_22159,N_21377);
xnor UO_628 (O_628,N_21143,N_21141);
xnor UO_629 (O_629,N_22901,N_23664);
or UO_630 (O_630,N_24535,N_21847);
xor UO_631 (O_631,N_24473,N_21434);
xnor UO_632 (O_632,N_24553,N_23744);
or UO_633 (O_633,N_22203,N_21004);
and UO_634 (O_634,N_22187,N_22496);
or UO_635 (O_635,N_23108,N_22763);
nor UO_636 (O_636,N_21041,N_24775);
xor UO_637 (O_637,N_24059,N_21867);
and UO_638 (O_638,N_23955,N_20670);
and UO_639 (O_639,N_23931,N_22075);
or UO_640 (O_640,N_21668,N_23732);
and UO_641 (O_641,N_20511,N_22293);
nand UO_642 (O_642,N_20538,N_23081);
nand UO_643 (O_643,N_23270,N_23647);
xor UO_644 (O_644,N_24708,N_21270);
nor UO_645 (O_645,N_21744,N_22972);
xor UO_646 (O_646,N_22260,N_24042);
or UO_647 (O_647,N_24028,N_24617);
or UO_648 (O_648,N_20958,N_24029);
xor UO_649 (O_649,N_23601,N_20693);
nor UO_650 (O_650,N_24426,N_23474);
or UO_651 (O_651,N_24346,N_21248);
xnor UO_652 (O_652,N_24614,N_24522);
xor UO_653 (O_653,N_23845,N_24715);
xor UO_654 (O_654,N_24169,N_23059);
and UO_655 (O_655,N_20554,N_20256);
or UO_656 (O_656,N_21478,N_24989);
xor UO_657 (O_657,N_21033,N_22553);
or UO_658 (O_658,N_20504,N_22231);
nand UO_659 (O_659,N_23534,N_21573);
nand UO_660 (O_660,N_24497,N_23894);
nand UO_661 (O_661,N_20961,N_24193);
and UO_662 (O_662,N_22418,N_24091);
xor UO_663 (O_663,N_22451,N_20036);
xnor UO_664 (O_664,N_21330,N_22657);
xor UO_665 (O_665,N_22748,N_24373);
nor UO_666 (O_666,N_21317,N_21884);
or UO_667 (O_667,N_20075,N_21929);
xor UO_668 (O_668,N_24968,N_22299);
nand UO_669 (O_669,N_22436,N_21755);
or UO_670 (O_670,N_23721,N_20559);
or UO_671 (O_671,N_20414,N_23855);
nor UO_672 (O_672,N_23905,N_22661);
and UO_673 (O_673,N_21274,N_23254);
nor UO_674 (O_674,N_24402,N_21378);
xor UO_675 (O_675,N_23310,N_22023);
nand UO_676 (O_676,N_21538,N_22825);
nor UO_677 (O_677,N_23103,N_23636);
nand UO_678 (O_678,N_20445,N_22463);
or UO_679 (O_679,N_23380,N_23491);
nor UO_680 (O_680,N_22088,N_21950);
nand UO_681 (O_681,N_21146,N_22219);
nand UO_682 (O_682,N_21760,N_20658);
nand UO_683 (O_683,N_22897,N_23454);
xnor UO_684 (O_684,N_24993,N_22598);
nand UO_685 (O_685,N_22421,N_20702);
nor UO_686 (O_686,N_24066,N_23050);
xor UO_687 (O_687,N_21527,N_21459);
xnor UO_688 (O_688,N_23929,N_24762);
or UO_689 (O_689,N_20983,N_21116);
xor UO_690 (O_690,N_23728,N_22566);
nor UO_691 (O_691,N_21913,N_23412);
or UO_692 (O_692,N_20312,N_20705);
and UO_693 (O_693,N_21653,N_24935);
xnor UO_694 (O_694,N_23917,N_23989);
and UO_695 (O_695,N_23862,N_24075);
xnor UO_696 (O_696,N_21958,N_24811);
nand UO_697 (O_697,N_23466,N_24981);
and UO_698 (O_698,N_22776,N_24280);
and UO_699 (O_699,N_20994,N_23798);
or UO_700 (O_700,N_21206,N_24952);
and UO_701 (O_701,N_22300,N_22499);
or UO_702 (O_702,N_22055,N_21565);
xor UO_703 (O_703,N_24389,N_20732);
nand UO_704 (O_704,N_23009,N_20850);
nand UO_705 (O_705,N_23229,N_23904);
or UO_706 (O_706,N_24273,N_21063);
nor UO_707 (O_707,N_20657,N_24220);
nand UO_708 (O_708,N_22039,N_24002);
nor UO_709 (O_709,N_22573,N_22914);
nand UO_710 (O_710,N_24578,N_24774);
nor UO_711 (O_711,N_24332,N_23000);
or UO_712 (O_712,N_20219,N_22474);
nand UO_713 (O_713,N_23569,N_23181);
or UO_714 (O_714,N_20584,N_24567);
or UO_715 (O_715,N_22226,N_21611);
xnor UO_716 (O_716,N_23206,N_23885);
xor UO_717 (O_717,N_24587,N_22184);
or UO_718 (O_718,N_20971,N_22476);
nor UO_719 (O_719,N_20350,N_20318);
or UO_720 (O_720,N_24235,N_24378);
nand UO_721 (O_721,N_22854,N_22910);
and UO_722 (O_722,N_23606,N_24937);
xnor UO_723 (O_723,N_23131,N_22032);
xor UO_724 (O_724,N_20535,N_21068);
nor UO_725 (O_725,N_24608,N_24472);
nor UO_726 (O_726,N_24794,N_24392);
nor UO_727 (O_727,N_22617,N_22943);
nand UO_728 (O_728,N_21590,N_20287);
nand UO_729 (O_729,N_21187,N_22140);
and UO_730 (O_730,N_22472,N_24468);
or UO_731 (O_731,N_20033,N_20190);
or UO_732 (O_732,N_20270,N_21220);
nor UO_733 (O_733,N_21359,N_22816);
or UO_734 (O_734,N_21280,N_20791);
and UO_735 (O_735,N_22102,N_24173);
or UO_736 (O_736,N_24080,N_21301);
and UO_737 (O_737,N_20346,N_20816);
xor UO_738 (O_738,N_21639,N_24733);
or UO_739 (O_739,N_20171,N_21724);
xor UO_740 (O_740,N_20576,N_22253);
nand UO_741 (O_741,N_21091,N_20450);
xor UO_742 (O_742,N_23936,N_21232);
nor UO_743 (O_743,N_23111,N_23922);
or UO_744 (O_744,N_22861,N_21843);
or UO_745 (O_745,N_20425,N_24184);
or UO_746 (O_746,N_24734,N_24945);
nand UO_747 (O_747,N_20884,N_24153);
nor UO_748 (O_748,N_23137,N_22425);
and UO_749 (O_749,N_20606,N_22541);
nor UO_750 (O_750,N_24910,N_24417);
or UO_751 (O_751,N_23912,N_20969);
nand UO_752 (O_752,N_23772,N_21468);
xnor UO_753 (O_753,N_23953,N_24386);
nor UO_754 (O_754,N_20688,N_21374);
nand UO_755 (O_755,N_24108,N_20968);
nor UO_756 (O_756,N_23805,N_24924);
nor UO_757 (O_757,N_21670,N_21254);
nor UO_758 (O_758,N_21981,N_24074);
xor UO_759 (O_759,N_23074,N_20319);
nand UO_760 (O_760,N_20669,N_22007);
and UO_761 (O_761,N_21136,N_21067);
nand UO_762 (O_762,N_21502,N_23144);
and UO_763 (O_763,N_23652,N_21659);
nor UO_764 (O_764,N_22694,N_23641);
and UO_765 (O_765,N_24170,N_24593);
or UO_766 (O_766,N_21128,N_22198);
or UO_767 (O_767,N_20146,N_24797);
or UO_768 (O_768,N_22817,N_23591);
nand UO_769 (O_769,N_20779,N_22358);
xor UO_770 (O_770,N_24723,N_23393);
nand UO_771 (O_771,N_21331,N_20193);
xor UO_772 (O_772,N_20368,N_21915);
nand UO_773 (O_773,N_20028,N_20875);
and UO_774 (O_774,N_20509,N_22094);
xnor UO_775 (O_775,N_23020,N_21284);
or UO_776 (O_776,N_23586,N_22416);
nor UO_777 (O_777,N_21390,N_21849);
nor UO_778 (O_778,N_21543,N_22563);
xnor UO_779 (O_779,N_22927,N_20753);
nor UO_780 (O_780,N_20650,N_22676);
and UO_781 (O_781,N_20916,N_22412);
nor UO_782 (O_782,N_22805,N_20865);
nor UO_783 (O_783,N_24765,N_24804);
nor UO_784 (O_784,N_20623,N_20161);
or UO_785 (O_785,N_23610,N_24955);
nand UO_786 (O_786,N_24017,N_22774);
or UO_787 (O_787,N_24065,N_24179);
nor UO_788 (O_788,N_22584,N_23054);
nand UO_789 (O_789,N_20018,N_20293);
nor UO_790 (O_790,N_24102,N_24237);
or UO_791 (O_791,N_22142,N_21381);
nor UO_792 (O_792,N_24045,N_23253);
or UO_793 (O_793,N_20069,N_22955);
or UO_794 (O_794,N_22852,N_23190);
nor UO_795 (O_795,N_20407,N_23232);
nor UO_796 (O_796,N_23329,N_21358);
xnor UO_797 (O_797,N_23724,N_22616);
xor UO_798 (O_798,N_23783,N_24162);
nor UO_799 (O_799,N_23627,N_20046);
nand UO_800 (O_800,N_24365,N_24656);
xnor UO_801 (O_801,N_23438,N_23085);
or UO_802 (O_802,N_23088,N_23747);
xnor UO_803 (O_803,N_20361,N_20317);
or UO_804 (O_804,N_23496,N_22501);
nor UO_805 (O_805,N_24699,N_24055);
nor UO_806 (O_806,N_22999,N_24642);
xor UO_807 (O_807,N_23626,N_22383);
and UO_808 (O_808,N_23432,N_22978);
nor UO_809 (O_809,N_24067,N_20238);
nand UO_810 (O_810,N_21554,N_20437);
xor UO_811 (O_811,N_20273,N_22005);
and UO_812 (O_812,N_24216,N_24325);
and UO_813 (O_813,N_22357,N_23453);
or UO_814 (O_814,N_22444,N_24778);
nand UO_815 (O_815,N_22342,N_20516);
nor UO_816 (O_816,N_22113,N_21416);
xnor UO_817 (O_817,N_23811,N_20009);
nor UO_818 (O_818,N_24331,N_22332);
and UO_819 (O_819,N_21077,N_21863);
and UO_820 (O_820,N_23848,N_23773);
xor UO_821 (O_821,N_23874,N_20588);
nand UO_822 (O_822,N_22274,N_20047);
nor UO_823 (O_823,N_22769,N_21876);
or UO_824 (O_824,N_22726,N_22942);
nand UO_825 (O_825,N_23655,N_20213);
or UO_826 (O_826,N_22201,N_21807);
xor UO_827 (O_827,N_21640,N_21761);
nand UO_828 (O_828,N_20823,N_21259);
or UO_829 (O_829,N_22346,N_24442);
or UO_830 (O_830,N_22221,N_24875);
or UO_831 (O_831,N_24963,N_20278);
xor UO_832 (O_832,N_24560,N_20276);
nand UO_833 (O_833,N_20837,N_21369);
or UO_834 (O_834,N_22671,N_20241);
nor UO_835 (O_835,N_20338,N_22404);
nand UO_836 (O_836,N_23762,N_20131);
xor UO_837 (O_837,N_23240,N_24246);
nand UO_838 (O_838,N_20970,N_22428);
and UO_839 (O_839,N_20902,N_24353);
xnor UO_840 (O_840,N_20840,N_23368);
and UO_841 (O_841,N_20624,N_20139);
nor UO_842 (O_842,N_20793,N_21995);
nor UO_843 (O_843,N_20900,N_24909);
xnor UO_844 (O_844,N_22870,N_20628);
nor UO_845 (O_845,N_24633,N_21388);
or UO_846 (O_846,N_20977,N_23105);
nor UO_847 (O_847,N_20503,N_20207);
xor UO_848 (O_848,N_24942,N_21654);
and UO_849 (O_849,N_21088,N_22919);
and UO_850 (O_850,N_22022,N_23207);
and UO_851 (O_851,N_20574,N_21454);
and UO_852 (O_852,N_21313,N_24333);
xnor UO_853 (O_853,N_23115,N_24755);
nor UO_854 (O_854,N_22734,N_23706);
nand UO_855 (O_855,N_24985,N_23426);
xor UO_856 (O_856,N_21292,N_23472);
nand UO_857 (O_857,N_21157,N_23501);
and UO_858 (O_858,N_24502,N_23471);
nor UO_859 (O_859,N_20087,N_24316);
xor UO_860 (O_860,N_20551,N_24431);
and UO_861 (O_861,N_20896,N_24238);
xor UO_862 (O_862,N_20434,N_24737);
nor UO_863 (O_863,N_22237,N_24359);
or UO_864 (O_864,N_22287,N_23505);
nor UO_865 (O_865,N_20921,N_22063);
nand UO_866 (O_866,N_22772,N_20745);
nor UO_867 (O_867,N_21703,N_20102);
nor UO_868 (O_868,N_21437,N_21446);
and UO_869 (O_869,N_24836,N_24110);
xnor UO_870 (O_870,N_21616,N_24590);
nand UO_871 (O_871,N_21183,N_21518);
or UO_872 (O_872,N_22026,N_20476);
and UO_873 (O_873,N_24503,N_24190);
or UO_874 (O_874,N_22896,N_23123);
and UO_875 (O_875,N_23522,N_24131);
xor UO_876 (O_876,N_21544,N_20357);
nor UO_877 (O_877,N_22449,N_20490);
xor UO_878 (O_878,N_22205,N_21357);
or UO_879 (O_879,N_24528,N_23261);
nand UO_880 (O_880,N_23431,N_20937);
xnor UO_881 (O_881,N_23420,N_24706);
xor UO_882 (O_882,N_20525,N_23866);
nor UO_883 (O_883,N_24171,N_22826);
nor UO_884 (O_884,N_22479,N_21070);
or UO_885 (O_885,N_23183,N_22324);
and UO_886 (O_886,N_21625,N_22384);
nor UO_887 (O_887,N_20508,N_22929);
nand UO_888 (O_888,N_22443,N_20681);
nor UO_889 (O_889,N_20498,N_24759);
nor UO_890 (O_890,N_22609,N_23897);
and UO_891 (O_891,N_21350,N_21511);
nand UO_892 (O_892,N_23971,N_23573);
or UO_893 (O_893,N_20150,N_23552);
or UO_894 (O_894,N_24495,N_21409);
and UO_895 (O_895,N_20194,N_20912);
xnor UO_896 (O_896,N_24966,N_23233);
nand UO_897 (O_897,N_23757,N_21968);
xor UO_898 (O_898,N_20589,N_20954);
or UO_899 (O_899,N_20269,N_21144);
or UO_900 (O_900,N_24959,N_22737);
nand UO_901 (O_901,N_21053,N_21746);
nand UO_902 (O_902,N_23618,N_21988);
and UO_903 (O_903,N_22240,N_23384);
nand UO_904 (O_904,N_21349,N_24596);
xnor UO_905 (O_905,N_21028,N_21591);
nor UO_906 (O_906,N_21430,N_23407);
or UO_907 (O_907,N_22095,N_23125);
or UO_908 (O_908,N_23467,N_20880);
or UO_909 (O_909,N_20722,N_24694);
xor UO_910 (O_910,N_23764,N_21229);
nor UO_911 (O_911,N_21781,N_24040);
or UO_912 (O_912,N_21909,N_23718);
nor UO_913 (O_913,N_21961,N_23282);
xor UO_914 (O_914,N_22962,N_20703);
or UO_915 (O_915,N_21059,N_20176);
nor UO_916 (O_916,N_23136,N_20925);
xnor UO_917 (O_917,N_23455,N_20781);
xnor UO_918 (O_918,N_23616,N_22400);
or UO_919 (O_919,N_24703,N_20463);
and UO_920 (O_920,N_23533,N_23022);
or UO_921 (O_921,N_21643,N_24048);
or UO_922 (O_922,N_22417,N_20264);
and UO_923 (O_923,N_22544,N_20653);
or UO_924 (O_924,N_21987,N_22549);
and UO_925 (O_925,N_23208,N_20251);
nand UO_926 (O_926,N_22249,N_23218);
nand UO_927 (O_927,N_22264,N_23045);
and UO_928 (O_928,N_21055,N_22595);
nor UO_929 (O_929,N_24022,N_23531);
nand UO_930 (O_930,N_20882,N_22271);
and UO_931 (O_931,N_22925,N_24772);
nor UO_932 (O_932,N_20742,N_20128);
and UO_933 (O_933,N_21989,N_21451);
xnor UO_934 (O_934,N_20236,N_24663);
nand UO_935 (O_935,N_24191,N_23997);
nand UO_936 (O_936,N_22907,N_20206);
and UO_937 (O_937,N_21965,N_21020);
xor UO_938 (O_938,N_22612,N_24527);
xor UO_939 (O_939,N_22419,N_22667);
xor UO_940 (O_940,N_20388,N_20521);
nand UO_941 (O_941,N_21608,N_22084);
nor UO_942 (O_942,N_20442,N_23524);
nand UO_943 (O_943,N_24939,N_22985);
nand UO_944 (O_944,N_23824,N_23052);
nor UO_945 (O_945,N_20091,N_23972);
xor UO_946 (O_946,N_21342,N_21283);
nor UO_947 (O_947,N_21085,N_23915);
or UO_948 (O_948,N_24978,N_21612);
or UO_949 (O_949,N_21747,N_22286);
nand UO_950 (O_950,N_22690,N_24078);
nand UO_951 (O_951,N_24659,N_24697);
xnor UO_952 (O_952,N_22990,N_24257);
xor UO_953 (O_953,N_20756,N_22498);
xnor UO_954 (O_954,N_22248,N_23246);
xnor UO_955 (O_955,N_24323,N_24873);
or UO_956 (O_956,N_21093,N_23483);
or UO_957 (O_957,N_22561,N_24658);
and UO_958 (O_958,N_20919,N_21966);
and UO_959 (O_959,N_21471,N_21130);
xor UO_960 (O_960,N_22702,N_24962);
xnor UO_961 (O_961,N_24999,N_24615);
xnor UO_962 (O_962,N_20972,N_22262);
or UO_963 (O_963,N_22235,N_23857);
nand UO_964 (O_964,N_22722,N_24210);
nand UO_965 (O_965,N_23299,N_21991);
and UO_966 (O_966,N_22229,N_23375);
xor UO_967 (O_967,N_20872,N_22610);
xor UO_968 (O_968,N_24263,N_21221);
nand UO_969 (O_969,N_24849,N_23446);
xnor UO_970 (O_970,N_23354,N_21304);
or UO_971 (O_971,N_24698,N_22001);
nor UO_972 (O_972,N_24223,N_20676);
nor UO_973 (O_973,N_22099,N_21931);
and UO_974 (O_974,N_24092,N_23429);
nor UO_975 (O_975,N_21779,N_21038);
and UO_976 (O_976,N_23513,N_23550);
nand UO_977 (O_977,N_22345,N_23830);
or UO_978 (O_978,N_21102,N_23667);
and UO_979 (O_979,N_20938,N_23901);
or UO_980 (O_980,N_20280,N_21551);
and UO_981 (O_981,N_23745,N_23686);
nand UO_982 (O_982,N_21857,N_20266);
nand UO_983 (O_983,N_23696,N_23843);
and UO_984 (O_984,N_21311,N_24319);
nor UO_985 (O_985,N_21812,N_21822);
xnor UO_986 (O_986,N_22031,N_24418);
xor UO_987 (O_987,N_21105,N_21992);
nor UO_988 (O_988,N_20097,N_22606);
xnor UO_989 (O_989,N_22326,N_21482);
and UO_990 (O_990,N_24853,N_20291);
nor UO_991 (O_991,N_23378,N_20853);
xnor UO_992 (O_992,N_23994,N_23711);
nor UO_993 (O_993,N_20486,N_21234);
or UO_994 (O_994,N_23748,N_20168);
and UO_995 (O_995,N_23592,N_24243);
and UO_996 (O_996,N_22872,N_21072);
nand UO_997 (O_997,N_20428,N_20406);
or UO_998 (O_998,N_20129,N_20074);
and UO_999 (O_999,N_24845,N_24921);
nor UO_1000 (O_1000,N_23002,N_24996);
nor UO_1001 (O_1001,N_20667,N_24988);
nor UO_1002 (O_1002,N_24063,N_23749);
nand UO_1003 (O_1003,N_22709,N_24800);
xnor UO_1004 (O_1004,N_22081,N_21151);
xnor UO_1005 (O_1005,N_23456,N_20862);
or UO_1006 (O_1006,N_22698,N_20789);
nor UO_1007 (O_1007,N_20237,N_23182);
nor UO_1008 (O_1008,N_24094,N_20096);
nand UO_1009 (O_1009,N_24728,N_24933);
nor UO_1010 (O_1010,N_21106,N_20866);
nor UO_1011 (O_1011,N_24494,N_22547);
and UO_1012 (O_1012,N_21737,N_23691);
or UO_1013 (O_1013,N_20211,N_24691);
nand UO_1014 (O_1014,N_24256,N_22091);
or UO_1015 (O_1015,N_23273,N_24115);
or UO_1016 (O_1016,N_21205,N_20590);
nor UO_1017 (O_1017,N_20427,N_21432);
or UO_1018 (O_1018,N_22801,N_21192);
xor UO_1019 (O_1019,N_24482,N_24655);
nor UO_1020 (O_1020,N_20932,N_23155);
nor UO_1021 (O_1021,N_22862,N_24652);
and UO_1022 (O_1022,N_23371,N_24842);
and UO_1023 (O_1023,N_20021,N_21494);
nor UO_1024 (O_1024,N_22680,N_22432);
nor UO_1025 (O_1025,N_20495,N_20802);
xor UO_1026 (O_1026,N_23024,N_23662);
or UO_1027 (O_1027,N_23211,N_23167);
xor UO_1028 (O_1028,N_21751,N_20039);
nor UO_1029 (O_1029,N_22471,N_21788);
nor UO_1030 (O_1030,N_21485,N_20854);
nand UO_1031 (O_1031,N_24354,N_24783);
nand UO_1032 (O_1032,N_23328,N_21990);
and UO_1033 (O_1033,N_21199,N_22659);
and UO_1034 (O_1034,N_20800,N_20245);
xor UO_1035 (O_1035,N_23480,N_20451);
nor UO_1036 (O_1036,N_21658,N_24155);
nor UO_1037 (O_1037,N_23032,N_20956);
nor UO_1038 (O_1038,N_24168,N_20095);
nand UO_1039 (O_1039,N_22228,N_21698);
or UO_1040 (O_1040,N_20531,N_24147);
and UO_1041 (O_1041,N_24255,N_21417);
nand UO_1042 (O_1042,N_22202,N_20715);
xnor UO_1043 (O_1043,N_23031,N_23005);
and UO_1044 (O_1044,N_22788,N_22433);
or UO_1045 (O_1045,N_22819,N_22906);
and UO_1046 (O_1046,N_21500,N_24479);
xor UO_1047 (O_1047,N_20660,N_21649);
nor UO_1048 (O_1048,N_23970,N_22278);
and UO_1049 (O_1049,N_24890,N_22134);
xor UO_1050 (O_1050,N_21879,N_20843);
or UO_1051 (O_1051,N_20646,N_21457);
and UO_1052 (O_1052,N_23490,N_23803);
nand UO_1053 (O_1053,N_20243,N_21211);
and UO_1054 (O_1054,N_22086,N_22934);
nand UO_1055 (O_1055,N_22276,N_24466);
nand UO_1056 (O_1056,N_24192,N_24511);
and UO_1057 (O_1057,N_21713,N_23291);
or UO_1058 (O_1058,N_21152,N_20965);
and UO_1059 (O_1059,N_23374,N_20472);
nor UO_1060 (O_1060,N_21045,N_21000);
xor UO_1061 (O_1061,N_23859,N_24582);
and UO_1062 (O_1062,N_22447,N_23038);
and UO_1063 (O_1063,N_24058,N_23145);
or UO_1064 (O_1064,N_21671,N_22627);
and UO_1065 (O_1065,N_23738,N_22605);
nor UO_1066 (O_1066,N_20460,N_23840);
or UO_1067 (O_1067,N_21826,N_23231);
nand UO_1068 (O_1068,N_23096,N_23977);
xnor UO_1069 (O_1069,N_22295,N_21896);
xnor UO_1070 (O_1070,N_24142,N_24695);
xnor UO_1071 (O_1071,N_24287,N_20068);
nor UO_1072 (O_1072,N_24887,N_21954);
xor UO_1073 (O_1073,N_21951,N_20936);
xnor UO_1074 (O_1074,N_21470,N_20563);
nor UO_1075 (O_1075,N_23822,N_22708);
or UO_1076 (O_1076,N_22466,N_24859);
nor UO_1077 (O_1077,N_21162,N_23973);
or UO_1078 (O_1078,N_21308,N_22587);
nor UO_1079 (O_1079,N_22716,N_24456);
and UO_1080 (O_1080,N_21707,N_21466);
nand UO_1081 (O_1081,N_22740,N_22889);
nand UO_1082 (O_1082,N_21595,N_23298);
or UO_1083 (O_1083,N_24761,N_24061);
nand UO_1084 (O_1084,N_20082,N_21147);
nor UO_1085 (O_1085,N_20540,N_22193);
nand UO_1086 (O_1086,N_20303,N_23353);
or UO_1087 (O_1087,N_22818,N_22853);
or UO_1088 (O_1088,N_24825,N_23237);
xnor UO_1089 (O_1089,N_24647,N_21732);
nor UO_1090 (O_1090,N_21693,N_23238);
nor UO_1091 (O_1091,N_22041,N_22732);
or UO_1092 (O_1092,N_23755,N_20174);
and UO_1093 (O_1093,N_20645,N_23084);
nor UO_1094 (O_1094,N_22284,N_23390);
or UO_1095 (O_1095,N_23106,N_22973);
xnor UO_1096 (O_1096,N_22998,N_22457);
or UO_1097 (O_1097,N_22367,N_21306);
nand UO_1098 (O_1098,N_22767,N_23358);
or UO_1099 (O_1099,N_23492,N_21119);
nor UO_1100 (O_1100,N_20665,N_20192);
xor UO_1101 (O_1101,N_24348,N_21586);
nand UO_1102 (O_1102,N_20825,N_21111);
and UO_1103 (O_1103,N_22711,N_23949);
or UO_1104 (O_1104,N_21904,N_22655);
nand UO_1105 (O_1105,N_20461,N_23903);
nor UO_1106 (O_1106,N_24872,N_24693);
xor UO_1107 (O_1107,N_20006,N_22963);
nand UO_1108 (O_1108,N_21555,N_24187);
nand UO_1109 (O_1109,N_24368,N_23741);
or UO_1110 (O_1110,N_21955,N_21557);
nand UO_1111 (O_1111,N_23776,N_20169);
and UO_1112 (O_1112,N_23703,N_22635);
nor UO_1113 (O_1113,N_22089,N_22894);
nor UO_1114 (O_1114,N_22515,N_24729);
or UO_1115 (O_1115,N_21816,N_20396);
or UO_1116 (O_1116,N_24926,N_20926);
or UO_1117 (O_1117,N_24030,N_22141);
and UO_1118 (O_1118,N_21319,N_22795);
nand UO_1119 (O_1119,N_24844,N_22829);
nand UO_1120 (O_1120,N_23638,N_20426);
and UO_1121 (O_1121,N_21721,N_23419);
or UO_1122 (O_1122,N_24222,N_20814);
xor UO_1123 (O_1123,N_23634,N_20158);
or UO_1124 (O_1124,N_20349,N_23012);
nand UO_1125 (O_1125,N_20090,N_24576);
or UO_1126 (O_1126,N_22784,N_20055);
nor UO_1127 (O_1127,N_22601,N_24275);
or UO_1128 (O_1128,N_24379,N_23067);
and UO_1129 (O_1129,N_22145,N_24557);
or UO_1130 (O_1130,N_21489,N_24629);
or UO_1131 (O_1131,N_22796,N_22322);
nor UO_1132 (O_1132,N_22440,N_23506);
and UO_1133 (O_1133,N_21413,N_21376);
or UO_1134 (O_1134,N_22485,N_24200);
xor UO_1135 (O_1135,N_20935,N_21115);
and UO_1136 (O_1136,N_22646,N_20685);
nor UO_1137 (O_1137,N_21323,N_21893);
nand UO_1138 (O_1138,N_24150,N_22705);
xor UO_1139 (O_1139,N_21682,N_20402);
nor UO_1140 (O_1140,N_22523,N_22683);
xor UO_1141 (O_1141,N_20759,N_23276);
nand UO_1142 (O_1142,N_23044,N_21395);
or UO_1143 (O_1143,N_20625,N_23797);
xor UO_1144 (O_1144,N_21953,N_21642);
xnor UO_1145 (O_1145,N_22077,N_24601);
nor UO_1146 (O_1146,N_21615,N_23056);
and UO_1147 (O_1147,N_21405,N_24326);
nand UO_1148 (O_1148,N_22511,N_21764);
nand UO_1149 (O_1149,N_24006,N_22798);
and UO_1150 (O_1150,N_21043,N_24423);
nand UO_1151 (O_1151,N_22047,N_22674);
nand UO_1152 (O_1152,N_22123,N_24768);
or UO_1153 (O_1153,N_22331,N_23363);
nand UO_1154 (O_1154,N_23838,N_23315);
nor UO_1155 (O_1155,N_20704,N_21241);
xnor UO_1156 (O_1156,N_23876,N_21126);
xnor UO_1157 (O_1157,N_20001,N_24036);
and UO_1158 (O_1158,N_22245,N_23809);
xor UO_1159 (O_1159,N_20600,N_21758);
or UO_1160 (O_1160,N_22951,N_22239);
nand UO_1161 (O_1161,N_21086,N_22320);
nor UO_1162 (O_1162,N_23118,N_23974);
and UO_1163 (O_1163,N_21575,N_23409);
nor UO_1164 (O_1164,N_24976,N_21584);
xnor UO_1165 (O_1165,N_20301,N_24548);
xor UO_1166 (O_1166,N_22230,N_20760);
or UO_1167 (O_1167,N_23528,N_24161);
xor UO_1168 (O_1168,N_22259,N_22583);
nand UO_1169 (O_1169,N_23678,N_23488);
nor UO_1170 (O_1170,N_20783,N_24247);
and UO_1171 (O_1171,N_24812,N_23609);
and UO_1172 (O_1172,N_22745,N_24499);
and UO_1173 (O_1173,N_23888,N_24520);
and UO_1174 (O_1174,N_23802,N_22049);
nor UO_1175 (O_1175,N_21777,N_23116);
or UO_1176 (O_1176,N_20686,N_21728);
nand UO_1177 (O_1177,N_20905,N_24221);
nor UO_1178 (O_1178,N_23632,N_24234);
nand UO_1179 (O_1179,N_21829,N_24035);
and UO_1180 (O_1180,N_20700,N_22626);
nor UO_1181 (O_1181,N_22131,N_20240);
or UO_1182 (O_1182,N_21082,N_24815);
nand UO_1183 (O_1183,N_20198,N_21534);
nand UO_1184 (O_1184,N_23021,N_20785);
nor UO_1185 (O_1185,N_20764,N_22371);
or UO_1186 (O_1186,N_24915,N_21638);
and UO_1187 (O_1187,N_20446,N_21729);
xnor UO_1188 (O_1188,N_24003,N_21411);
and UO_1189 (O_1189,N_24839,N_20283);
nor UO_1190 (O_1190,N_21420,N_20059);
and UO_1191 (O_1191,N_21207,N_21665);
or UO_1192 (O_1192,N_22107,N_22224);
xor UO_1193 (O_1193,N_23281,N_22903);
and UO_1194 (O_1194,N_24016,N_20515);
nor UO_1195 (O_1195,N_24861,N_22857);
xnor UO_1196 (O_1196,N_24281,N_21855);
nand UO_1197 (O_1197,N_20042,N_20308);
nand UO_1198 (O_1198,N_20949,N_23514);
and UO_1199 (O_1199,N_21916,N_23813);
nand UO_1200 (O_1200,N_22065,N_24397);
nand UO_1201 (O_1201,N_20268,N_22582);
and UO_1202 (O_1202,N_22361,N_20930);
nand UO_1203 (O_1203,N_21712,N_21010);
or UO_1204 (O_1204,N_23091,N_23200);
nand UO_1205 (O_1205,N_24440,N_20134);
nor UO_1206 (O_1206,N_21720,N_20332);
nor UO_1207 (O_1207,N_24447,N_21666);
or UO_1208 (O_1208,N_24453,N_22338);
xor UO_1209 (O_1209,N_20408,N_24229);
nor UO_1210 (O_1210,N_21631,N_22082);
nand UO_1211 (O_1211,N_24982,N_23590);
and UO_1212 (O_1212,N_22186,N_21191);
xnor UO_1213 (O_1213,N_23526,N_20132);
nand UO_1214 (O_1214,N_24508,N_22132);
nor UO_1215 (O_1215,N_21246,N_20863);
or UO_1216 (O_1216,N_24318,N_23828);
nor UO_1217 (O_1217,N_23710,N_21983);
or UO_1218 (O_1218,N_23705,N_22151);
nand UO_1219 (O_1219,N_23333,N_23500);
or UO_1220 (O_1220,N_20967,N_20980);
and UO_1221 (O_1221,N_20778,N_24226);
nand UO_1222 (O_1222,N_21552,N_20449);
nor UO_1223 (O_1223,N_21285,N_22691);
or UO_1224 (O_1224,N_22958,N_22970);
nor UO_1225 (O_1225,N_20292,N_21889);
xnor UO_1226 (O_1226,N_22438,N_21610);
xor UO_1227 (O_1227,N_22741,N_24589);
xnor UO_1228 (O_1228,N_22362,N_24163);
nand UO_1229 (O_1229,N_20410,N_24683);
nand UO_1230 (O_1230,N_22808,N_22393);
nor UO_1231 (O_1231,N_24954,N_23529);
nor UO_1232 (O_1232,N_21392,N_24907);
nand UO_1233 (O_1233,N_23557,N_22863);
or UO_1234 (O_1234,N_20530,N_21977);
or UO_1235 (O_1235,N_22252,N_20960);
nor UO_1236 (O_1236,N_21421,N_21410);
nor UO_1237 (O_1237,N_24611,N_20117);
and UO_1238 (O_1238,N_20598,N_20723);
nor UO_1239 (O_1239,N_23192,N_20462);
xor UO_1240 (O_1240,N_22317,N_20057);
xnor UO_1241 (O_1241,N_20455,N_23173);
and UO_1242 (O_1242,N_23846,N_23080);
nor UO_1243 (O_1243,N_24819,N_23999);
nand UO_1244 (O_1244,N_20290,N_23734);
nor UO_1245 (O_1245,N_21224,N_22195);
nand UO_1246 (O_1246,N_21526,N_23555);
or UO_1247 (O_1247,N_24401,N_23867);
nor UO_1248 (O_1248,N_23156,N_21300);
and UO_1249 (O_1249,N_22124,N_22354);
nand UO_1250 (O_1250,N_23457,N_22282);
or UO_1251 (O_1251,N_20948,N_24489);
and UO_1252 (O_1252,N_23015,N_23293);
nand UO_1253 (O_1253,N_23611,N_23296);
or UO_1254 (O_1254,N_22071,N_23666);
nand UO_1255 (O_1255,N_23364,N_22731);
nor UO_1256 (O_1256,N_24470,N_24832);
nor UO_1257 (O_1257,N_24228,N_21716);
or UO_1258 (O_1258,N_23532,N_23405);
and UO_1259 (O_1259,N_21754,N_20940);
xor UO_1260 (O_1260,N_22136,N_24321);
nand UO_1261 (O_1261,N_21225,N_23965);
or UO_1262 (O_1262,N_22849,N_24292);
and UO_1263 (O_1263,N_21170,N_23635);
nand UO_1264 (O_1264,N_21058,N_21553);
or UO_1265 (O_1265,N_20718,N_20111);
xnor UO_1266 (O_1266,N_22681,N_20689);
and UO_1267 (O_1267,N_23858,N_21934);
and UO_1268 (O_1268,N_20957,N_20558);
and UO_1269 (O_1269,N_20195,N_20728);
and UO_1270 (O_1270,N_21195,N_24336);
or UO_1271 (O_1271,N_24624,N_21856);
or UO_1272 (O_1272,N_24805,N_23152);
xnor UO_1273 (O_1273,N_21037,N_21921);
nand UO_1274 (O_1274,N_23818,N_20643);
nand UO_1275 (O_1275,N_21687,N_23510);
nand UO_1276 (O_1276,N_20358,N_21523);
nor UO_1277 (O_1277,N_22969,N_24513);
nand UO_1278 (O_1278,N_23620,N_23227);
and UO_1279 (O_1279,N_21477,N_24880);
and UO_1280 (O_1280,N_23992,N_20908);
and UO_1281 (O_1281,N_20668,N_23665);
xor UO_1282 (O_1282,N_20429,N_22744);
nor UO_1283 (O_1283,N_23078,N_24224);
nand UO_1284 (O_1284,N_20366,N_21264);
or UO_1285 (O_1285,N_20577,N_23244);
nand UO_1286 (O_1286,N_23066,N_24835);
or UO_1287 (O_1287,N_21444,N_21515);
xor UO_1288 (O_1288,N_20644,N_20888);
nor UO_1289 (O_1289,N_22452,N_23048);
and UO_1290 (O_1290,N_22297,N_21773);
or UO_1291 (O_1291,N_22218,N_21648);
or UO_1292 (O_1292,N_22109,N_23782);
nand UO_1293 (O_1293,N_22365,N_24822);
nand UO_1294 (O_1294,N_24244,N_23458);
or UO_1295 (O_1295,N_22672,N_23398);
nor UO_1296 (O_1296,N_22869,N_21464);
nor UO_1297 (O_1297,N_24808,N_21895);
nand UO_1298 (O_1298,N_24773,N_20229);
or UO_1299 (O_1299,N_23833,N_22949);
xor UO_1300 (O_1300,N_21460,N_21347);
xor UO_1301 (O_1301,N_23849,N_23547);
nor UO_1302 (O_1302,N_23785,N_20382);
nor UO_1303 (O_1303,N_23567,N_21481);
nand UO_1304 (O_1304,N_24427,N_24214);
nand UO_1305 (O_1305,N_23427,N_20149);
and UO_1306 (O_1306,N_20901,N_24212);
nand UO_1307 (O_1307,N_23202,N_24471);
and UO_1308 (O_1308,N_20221,N_23680);
and UO_1309 (O_1309,N_22402,N_21021);
or UO_1310 (O_1310,N_20599,N_20950);
and UO_1311 (O_1311,N_24258,N_23623);
or UO_1312 (O_1312,N_24764,N_23639);
or UO_1313 (O_1313,N_21799,N_21925);
and UO_1314 (O_1314,N_24347,N_23306);
or UO_1315 (O_1315,N_21108,N_22898);
nor UO_1316 (O_1316,N_22570,N_20322);
nand UO_1317 (O_1317,N_22522,N_21475);
and UO_1318 (O_1318,N_24151,N_21235);
nor UO_1319 (O_1319,N_20452,N_21198);
and UO_1320 (O_1320,N_22521,N_22423);
nor UO_1321 (O_1321,N_20247,N_23900);
xnor UO_1322 (O_1322,N_20330,N_21483);
and UO_1323 (O_1323,N_22011,N_21805);
nand UO_1324 (O_1324,N_24579,N_22161);
nand UO_1325 (O_1325,N_22273,N_21960);
nand UO_1326 (O_1326,N_24785,N_20820);
or UO_1327 (O_1327,N_23037,N_21636);
nor UO_1328 (O_1328,N_20231,N_23445);
nand UO_1329 (O_1329,N_24010,N_23887);
and UO_1330 (O_1330,N_21249,N_21050);
or UO_1331 (O_1331,N_21520,N_22238);
or UO_1332 (O_1332,N_20545,N_20973);
and UO_1333 (O_1333,N_24342,N_22296);
nor UO_1334 (O_1334,N_23418,N_21571);
xor UO_1335 (O_1335,N_24700,N_24124);
nand UO_1336 (O_1336,N_20878,N_24088);
and UO_1337 (O_1337,N_24638,N_20608);
nor UO_1338 (O_1338,N_22392,N_21261);
and UO_1339 (O_1339,N_22017,N_24144);
and UO_1340 (O_1340,N_21506,N_20982);
xnor UO_1341 (O_1341,N_23220,N_23633);
nand UO_1342 (O_1342,N_22181,N_22793);
nor UO_1343 (O_1343,N_23424,N_22139);
or UO_1344 (O_1344,N_23481,N_22540);
xor UO_1345 (O_1345,N_22887,N_22497);
xnor UO_1346 (O_1346,N_23285,N_21057);
xnor UO_1347 (O_1347,N_20142,N_20858);
or UO_1348 (O_1348,N_22227,N_23572);
nor UO_1349 (O_1349,N_22871,N_24492);
and UO_1350 (O_1350,N_20697,N_23019);
xor UO_1351 (O_1351,N_21824,N_21190);
xnor UO_1352 (O_1352,N_20258,N_23444);
or UO_1353 (O_1353,N_21619,N_20441);
or UO_1354 (O_1354,N_20077,N_20552);
or UO_1355 (O_1355,N_21742,N_20162);
xnor UO_1356 (O_1356,N_23230,N_21560);
xor UO_1357 (O_1357,N_20103,N_23969);
and UO_1358 (O_1358,N_24038,N_20514);
and UO_1359 (O_1359,N_20184,N_23926);
and UO_1360 (O_1360,N_21172,N_24973);
or UO_1361 (O_1361,N_22340,N_20371);
or UO_1362 (O_1362,N_21609,N_24464);
or UO_1363 (O_1363,N_22996,N_20612);
nor UO_1364 (O_1364,N_23326,N_22096);
nor UO_1365 (O_1365,N_23079,N_20769);
or UO_1366 (O_1366,N_24290,N_20257);
nor UO_1367 (O_1367,N_22206,N_24050);
and UO_1368 (O_1368,N_21765,N_21340);
nor UO_1369 (O_1369,N_21008,N_23987);
and UO_1370 (O_1370,N_21952,N_21480);
nor UO_1371 (O_1371,N_23574,N_23076);
xnor UO_1372 (O_1372,N_20398,N_23541);
xnor UO_1373 (O_1373,N_20740,N_21305);
or UO_1374 (O_1374,N_24854,N_20457);
nand UO_1375 (O_1375,N_20721,N_23663);
xnor UO_1376 (O_1376,N_23883,N_24564);
and UO_1377 (O_1377,N_24420,N_23733);
nor UO_1378 (O_1378,N_22083,N_21979);
or UO_1379 (O_1379,N_20326,N_22642);
nand UO_1380 (O_1380,N_22546,N_22370);
nand UO_1381 (O_1381,N_23216,N_23947);
or UO_1382 (O_1382,N_21542,N_24504);
and UO_1383 (O_1383,N_24898,N_24625);
or UO_1384 (O_1384,N_22125,N_20344);
and UO_1385 (O_1385,N_22185,N_21114);
xor UO_1386 (O_1386,N_22891,N_22935);
and UO_1387 (O_1387,N_21985,N_23913);
nor UO_1388 (O_1388,N_20794,N_23350);
xor UO_1389 (O_1389,N_24833,N_24416);
and UO_1390 (O_1390,N_22660,N_20572);
nor UO_1391 (O_1391,N_24682,N_20299);
and UO_1392 (O_1392,N_22315,N_23891);
xor UO_1393 (O_1393,N_24634,N_23515);
nor UO_1394 (O_1394,N_24990,N_21361);
or UO_1395 (O_1395,N_20512,N_20613);
xor UO_1396 (O_1396,N_21353,N_21731);
xor UO_1397 (O_1397,N_24400,N_24753);
nor UO_1398 (O_1398,N_22058,N_21957);
nor UO_1399 (O_1399,N_24575,N_20553);
nand UO_1400 (O_1400,N_20379,N_20415);
and UO_1401 (O_1401,N_20484,N_23197);
or UO_1402 (O_1402,N_23812,N_23497);
xnor UO_1403 (O_1403,N_21176,N_20325);
and UO_1404 (O_1404,N_22090,N_23205);
xnor UO_1405 (O_1405,N_23643,N_20801);
nand UO_1406 (O_1406,N_24384,N_20300);
and UO_1407 (O_1407,N_21572,N_21026);
nor UO_1408 (O_1408,N_24304,N_24189);
xor UO_1409 (O_1409,N_21834,N_24100);
xor UO_1410 (O_1410,N_24419,N_22256);
and UO_1411 (O_1411,N_21641,N_22992);
xor UO_1412 (O_1412,N_21332,N_21463);
nor UO_1413 (O_1413,N_23980,N_24632);
and UO_1414 (O_1414,N_24983,N_20673);
and UO_1415 (O_1415,N_24879,N_22307);
or UO_1416 (O_1416,N_23134,N_22835);
nand UO_1417 (O_1417,N_21165,N_23493);
or UO_1418 (O_1418,N_22085,N_22103);
nor UO_1419 (O_1419,N_20093,N_24481);
or UO_1420 (O_1420,N_24288,N_20627);
and UO_1421 (O_1421,N_20561,N_20765);
nand UO_1422 (O_1422,N_22895,N_22196);
or UO_1423 (O_1423,N_20435,N_22369);
xor UO_1424 (O_1424,N_24262,N_22954);
and UO_1425 (O_1425,N_24512,N_20246);
nor UO_1426 (O_1426,N_22802,N_24314);
xnor UO_1427 (O_1427,N_24597,N_21937);
nand UO_1428 (O_1428,N_22487,N_23396);
or UO_1429 (O_1429,N_22137,N_22062);
nor UO_1430 (O_1430,N_24791,N_21404);
and UO_1431 (O_1431,N_24004,N_21622);
nor UO_1432 (O_1432,N_20200,N_24709);
nor UO_1433 (O_1433,N_24469,N_21837);
nand UO_1434 (O_1434,N_24208,N_20105);
nor UO_1435 (O_1435,N_24782,N_22038);
and UO_1436 (O_1436,N_20578,N_24120);
nand UO_1437 (O_1437,N_21679,N_20796);
and UO_1438 (O_1438,N_22199,N_24546);
xnor UO_1439 (O_1439,N_20927,N_21336);
xnor UO_1440 (O_1440,N_21725,N_22848);
nor UO_1441 (O_1441,N_21715,N_22559);
xnor UO_1442 (O_1442,N_21644,N_21768);
or UO_1443 (O_1443,N_21030,N_20797);
or UO_1444 (O_1444,N_21839,N_23869);
or UO_1445 (O_1445,N_23434,N_20440);
nor UO_1446 (O_1446,N_21908,N_23349);
nor UO_1447 (O_1447,N_23433,N_21704);
nand UO_1448 (O_1448,N_22844,N_23057);
or UO_1449 (O_1449,N_24330,N_22052);
and UO_1450 (O_1450,N_24291,N_24041);
or UO_1451 (O_1451,N_24891,N_24324);
nand UO_1452 (O_1452,N_22507,N_22989);
nand UO_1453 (O_1453,N_20045,N_22810);
nand UO_1454 (O_1454,N_23387,N_24205);
or UO_1455 (O_1455,N_20088,N_24232);
nand UO_1456 (O_1456,N_23441,N_24011);
and UO_1457 (O_1457,N_21559,N_22855);
nor UO_1458 (O_1458,N_20485,N_21253);
or UO_1459 (O_1459,N_23053,N_24630);
xor UO_1460 (O_1460,N_21525,N_21923);
xnor UO_1461 (O_1461,N_20401,N_21078);
xor UO_1462 (O_1462,N_22316,N_21861);
and UO_1463 (O_1463,N_21888,N_21745);
xnor UO_1464 (O_1464,N_22351,N_23956);
nand UO_1465 (O_1465,N_21516,N_20654);
and UO_1466 (O_1466,N_22183,N_22603);
and UO_1467 (O_1467,N_24076,N_24254);
nand UO_1468 (O_1468,N_24195,N_24970);
xor UO_1469 (O_1469,N_21905,N_23468);
xor UO_1470 (O_1470,N_23300,N_21688);
and UO_1471 (O_1471,N_22437,N_20881);
or UO_1472 (O_1472,N_22703,N_20564);
xor UO_1473 (O_1473,N_20339,N_22429);
xor UO_1474 (O_1474,N_23554,N_24001);
xor UO_1475 (O_1475,N_23323,N_21859);
nor UO_1476 (O_1476,N_24340,N_22192);
nor UO_1477 (O_1477,N_22594,N_23886);
nor UO_1478 (O_1478,N_21427,N_20015);
or UO_1479 (O_1479,N_21243,N_23272);
and UO_1480 (O_1480,N_20524,N_20604);
nand UO_1481 (O_1481,N_23581,N_23693);
and UO_1482 (O_1482,N_20683,N_24681);
nand UO_1483 (O_1483,N_22455,N_24701);
or UO_1484 (O_1484,N_24769,N_20196);
and UO_1485 (O_1485,N_20274,N_21322);
and UO_1486 (O_1486,N_24432,N_21798);
or UO_1487 (O_1487,N_24876,N_24014);
nor UO_1488 (O_1488,N_24727,N_21024);
xor UO_1489 (O_1489,N_21549,N_24758);
nor UO_1490 (O_1490,N_20387,N_24009);
or UO_1491 (O_1491,N_23719,N_20110);
nand UO_1492 (O_1492,N_21680,N_23945);
and UO_1493 (O_1493,N_23014,N_24012);
and UO_1494 (O_1494,N_24731,N_23875);
or UO_1495 (O_1495,N_24616,N_22150);
nor UO_1496 (O_1496,N_22543,N_21073);
or UO_1497 (O_1497,N_20629,N_22639);
and UO_1498 (O_1498,N_22156,N_23027);
or UO_1499 (O_1499,N_24283,N_21509);
xnor UO_1500 (O_1500,N_20372,N_21079);
xnor UO_1501 (O_1501,N_20784,N_22349);
or UO_1502 (O_1502,N_22396,N_22747);
nand UO_1503 (O_1503,N_23651,N_22070);
or UO_1504 (O_1504,N_23442,N_20672);
xor UO_1505 (O_1505,N_23753,N_24789);
nor UO_1506 (O_1506,N_24653,N_21214);
or UO_1507 (O_1507,N_23342,N_20809);
nor UO_1508 (O_1508,N_23909,N_22754);
and UO_1509 (O_1509,N_22030,N_22684);
and UO_1510 (O_1510,N_21467,N_22994);
or UO_1511 (O_1511,N_20999,N_24207);
nor UO_1512 (O_1512,N_23924,N_24141);
nand UO_1513 (O_1513,N_24308,N_20945);
xor UO_1514 (O_1514,N_23255,N_23568);
or UO_1515 (O_1515,N_23391,N_22171);
and UO_1516 (O_1516,N_21694,N_20601);
or UO_1517 (O_1517,N_24806,N_24803);
and UO_1518 (O_1518,N_22625,N_24364);
or UO_1519 (O_1519,N_21389,N_21439);
nand UO_1520 (O_1520,N_21873,N_24185);
nand UO_1521 (O_1521,N_22015,N_22092);
or UO_1522 (O_1522,N_21948,N_20701);
and UO_1523 (O_1523,N_21291,N_21795);
and UO_1524 (O_1524,N_22760,N_22764);
xor UO_1525 (O_1525,N_21903,N_22586);
xor UO_1526 (O_1526,N_24840,N_20909);
xor UO_1527 (O_1527,N_20086,N_23109);
and UO_1528 (O_1528,N_23605,N_23082);
nor UO_1529 (O_1529,N_24860,N_20849);
nor UO_1530 (O_1530,N_20602,N_21930);
xor UO_1531 (O_1531,N_22394,N_23258);
nand UO_1532 (O_1532,N_22492,N_21566);
nor UO_1533 (O_1533,N_21734,N_22503);
xnor UO_1534 (O_1534,N_24577,N_24598);
or UO_1535 (O_1535,N_24902,N_24786);
nand UO_1536 (O_1536,N_21318,N_24462);
or UO_1537 (O_1537,N_21769,N_24054);
nor UO_1538 (O_1538,N_24931,N_21673);
nor UO_1539 (O_1539,N_21576,N_20345);
and UO_1540 (O_1540,N_20385,N_21184);
nand UO_1541 (O_1541,N_21832,N_21936);
xnor UO_1542 (O_1542,N_20029,N_22790);
or UO_1543 (O_1543,N_23337,N_22578);
nand UO_1544 (O_1544,N_21570,N_24961);
xor UO_1545 (O_1545,N_20939,N_20727);
or UO_1546 (O_1546,N_22880,N_22637);
nor UO_1547 (O_1547,N_23933,N_21023);
nand UO_1548 (O_1548,N_23003,N_21299);
nor UO_1549 (O_1549,N_20792,N_21110);
nand UO_1550 (O_1550,N_21854,N_24802);
nor UO_1551 (O_1551,N_24874,N_21169);
nor UO_1552 (O_1552,N_22303,N_23963);
nand UO_1553 (O_1553,N_24750,N_23243);
or UO_1554 (O_1554,N_23213,N_24196);
or UO_1555 (O_1555,N_22678,N_23660);
nor UO_1556 (O_1556,N_23925,N_22465);
nand UO_1557 (O_1557,N_22467,N_22786);
nor UO_1558 (O_1558,N_22856,N_24301);
xor UO_1559 (O_1559,N_23449,N_20717);
nor UO_1560 (O_1560,N_23759,N_24643);
and UO_1561 (O_1561,N_22223,N_23307);
nor UO_1562 (O_1562,N_24517,N_20212);
and UO_1563 (O_1563,N_21772,N_21701);
xnor UO_1564 (O_1564,N_22018,N_23386);
or UO_1565 (O_1565,N_23146,N_24657);
xnor UO_1566 (O_1566,N_23967,N_21994);
and UO_1567 (O_1567,N_22119,N_24356);
and UO_1568 (O_1568,N_23964,N_20491);
nand UO_1569 (O_1569,N_24667,N_23631);
nand UO_1570 (O_1570,N_23359,N_22486);
nor UO_1571 (O_1571,N_23346,N_22302);
and UO_1572 (O_1572,N_24313,N_21399);
nor UO_1573 (O_1573,N_24516,N_20315);
nor UO_1574 (O_1574,N_21675,N_23107);
nor UO_1575 (O_1575,N_20648,N_21382);
or UO_1576 (O_1576,N_24675,N_24233);
or UO_1577 (O_1577,N_24826,N_22477);
and UO_1578 (O_1578,N_21074,N_21181);
nor UO_1579 (O_1579,N_22243,N_22304);
and UO_1580 (O_1580,N_20923,N_21271);
or UO_1581 (O_1581,N_21307,N_22840);
nor UO_1582 (O_1582,N_20127,N_22493);
nand UO_1583 (O_1583,N_23286,N_23893);
or UO_1584 (O_1584,N_23584,N_22029);
nand UO_1585 (O_1585,N_20603,N_20636);
or UO_1586 (O_1586,N_23906,N_20741);
xor UO_1587 (O_1587,N_24908,N_23781);
or UO_1588 (O_1588,N_21836,N_20962);
nor UO_1589 (O_1589,N_20944,N_23194);
nor UO_1590 (O_1590,N_21062,N_20048);
and UO_1591 (O_1591,N_23421,N_20083);
or UO_1592 (O_1592,N_23761,N_20651);
xor UO_1593 (O_1593,N_21776,N_23804);
and UO_1594 (O_1594,N_23266,N_20773);
nand UO_1595 (O_1595,N_23110,N_22335);
and UO_1596 (O_1596,N_22664,N_21245);
and UO_1597 (O_1597,N_23249,N_21750);
nor UO_1598 (O_1598,N_21563,N_24883);
nor UO_1599 (O_1599,N_24943,N_22888);
nor UO_1600 (O_1600,N_20674,N_24770);
nand UO_1601 (O_1601,N_24801,N_24369);
nand UO_1602 (O_1602,N_22550,N_24438);
xnor UO_1603 (O_1603,N_20089,N_23998);
and UO_1604 (O_1604,N_20675,N_20537);
or UO_1605 (O_1605,N_24372,N_20327);
and UO_1606 (O_1606,N_24202,N_21352);
nor UO_1607 (O_1607,N_21161,N_20470);
nand UO_1608 (O_1608,N_23559,N_20466);
xnor UO_1609 (O_1609,N_20915,N_24799);
nand UO_1610 (O_1610,N_22149,N_23921);
or UO_1611 (O_1611,N_20232,N_23594);
nand UO_1612 (O_1612,N_20895,N_23794);
or UO_1613 (O_1613,N_24543,N_24588);
and UO_1614 (O_1614,N_20534,N_24476);
and UO_1615 (O_1615,N_20637,N_21838);
nand UO_1616 (O_1616,N_20680,N_20489);
and UO_1617 (O_1617,N_21561,N_24096);
nor UO_1618 (O_1618,N_20182,N_24573);
xor UO_1619 (O_1619,N_24104,N_23566);
xor UO_1620 (O_1620,N_24412,N_22314);
xnor UO_1621 (O_1621,N_21932,N_23976);
nor UO_1622 (O_1622,N_22768,N_22623);
or UO_1623 (O_1623,N_24450,N_22554);
nand UO_1624 (O_1624,N_24940,N_20731);
and UO_1625 (O_1625,N_20471,N_23737);
nand UO_1626 (O_1626,N_24648,N_22719);
nor UO_1627 (O_1627,N_20126,N_21278);
or UO_1628 (O_1628,N_20026,N_23265);
or UO_1629 (O_1629,N_22246,N_23699);
xnor UO_1630 (O_1630,N_21257,N_20710);
or UO_1631 (O_1631,N_21312,N_22519);
and UO_1632 (O_1632,N_21465,N_21871);
and UO_1633 (O_1633,N_22076,N_23792);
xor UO_1634 (O_1634,N_23165,N_21425);
xor UO_1635 (O_1635,N_20279,N_24767);
nor UO_1636 (O_1636,N_22157,N_24382);
nand UO_1637 (O_1637,N_20885,N_23837);
nor UO_1638 (O_1638,N_20013,N_23943);
or UO_1639 (O_1639,N_23422,N_20413);
or UO_1640 (O_1640,N_20518,N_23351);
or UO_1641 (O_1641,N_22874,N_21153);
or UO_1642 (O_1642,N_21749,N_24581);
or UO_1643 (O_1643,N_23700,N_21065);
nor UO_1644 (O_1644,N_21503,N_21496);
nand UO_1645 (O_1645,N_24545,N_21892);
xnor UO_1646 (O_1646,N_23765,N_22938);
and UO_1647 (O_1647,N_20311,N_21419);
and UO_1648 (O_1648,N_20369,N_23287);
nor UO_1649 (O_1649,N_22236,N_22677);
nor UO_1650 (O_1650,N_24201,N_20582);
xor UO_1651 (O_1651,N_22215,N_24641);
or UO_1652 (O_1652,N_23842,N_22040);
nand UO_1653 (O_1653,N_21341,N_21290);
and UO_1654 (O_1654,N_21098,N_21348);
and UO_1655 (O_1655,N_24480,N_23225);
or UO_1656 (O_1656,N_22866,N_24580);
xnor UO_1657 (O_1657,N_23746,N_23688);
and UO_1658 (O_1658,N_24315,N_21973);
or UO_1659 (O_1659,N_22078,N_24562);
xor UO_1660 (O_1660,N_23184,N_22794);
or UO_1661 (O_1661,N_23406,N_21488);
and UO_1662 (O_1662,N_24838,N_20041);
and UO_1663 (O_1663,N_20768,N_21942);
and UO_1664 (O_1664,N_20298,N_22292);
or UO_1665 (O_1665,N_23770,N_21997);
or UO_1666 (O_1666,N_22822,N_21137);
nor UO_1667 (O_1667,N_22960,N_24125);
xnor UO_1668 (O_1668,N_21239,N_21771);
nor UO_1669 (O_1669,N_21039,N_23122);
and UO_1670 (O_1670,N_24714,N_21733);
and UO_1671 (O_1671,N_20726,N_24787);
or UO_1672 (O_1672,N_24245,N_24730);
nand UO_1673 (O_1673,N_21912,N_22163);
nor UO_1674 (O_1674,N_24747,N_21569);
xor UO_1675 (O_1675,N_24953,N_22858);
xnor UO_1676 (O_1676,N_24087,N_20750);
nor UO_1677 (O_1677,N_22531,N_20242);
nor UO_1678 (O_1678,N_24441,N_21164);
or UO_1679 (O_1679,N_23334,N_23330);
nand UO_1680 (O_1680,N_20614,N_22341);
and UO_1681 (O_1681,N_21974,N_21393);
xnor UO_1682 (O_1682,N_24327,N_22742);
or UO_1683 (O_1683,N_23946,N_24312);
and UO_1684 (O_1684,N_20076,N_20144);
nor UO_1685 (O_1685,N_22072,N_20662);
and UO_1686 (O_1686,N_23617,N_23162);
nor UO_1687 (O_1687,N_24477,N_22638);
xnor UO_1688 (O_1688,N_21125,N_22755);
or UO_1689 (O_1689,N_24754,N_23659);
or UO_1690 (O_1690,N_23317,N_24702);
or UO_1691 (O_1691,N_23575,N_21118);
nand UO_1692 (O_1692,N_20324,N_21006);
or UO_1693 (O_1693,N_22514,N_22459);
nor UO_1694 (O_1694,N_22165,N_24711);
nor UO_1695 (O_1695,N_23851,N_24680);
nand UO_1696 (O_1696,N_20787,N_20569);
or UO_1697 (O_1697,N_24752,N_21784);
and UO_1698 (O_1698,N_24618,N_23018);
xnor UO_1699 (O_1699,N_23143,N_22290);
or UO_1700 (O_1700,N_22538,N_21422);
or UO_1701 (O_1701,N_22172,N_23130);
xnor UO_1702 (O_1702,N_22714,N_23011);
or UO_1703 (O_1703,N_22403,N_20684);
nand UO_1704 (O_1704,N_23402,N_20690);
and UO_1705 (O_1705,N_24383,N_20284);
nor UO_1706 (O_1706,N_23369,N_20874);
nor UO_1707 (O_1707,N_24411,N_21596);
and UO_1708 (O_1708,N_23452,N_23288);
nand UO_1709 (O_1709,N_21044,N_22556);
xor UO_1710 (O_1710,N_24660,N_20309);
and UO_1711 (O_1711,N_23826,N_21090);
and UO_1712 (O_1712,N_24998,N_22373);
nand UO_1713 (O_1713,N_23621,N_20244);
xnor UO_1714 (O_1714,N_23075,N_20154);
xor UO_1715 (O_1715,N_22155,N_22517);
or UO_1716 (O_1716,N_21823,N_21408);
xor UO_1717 (O_1717,N_21103,N_24357);
xor UO_1718 (O_1718,N_21651,N_24339);
and UO_1719 (O_1719,N_22766,N_21803);
xnor UO_1720 (O_1720,N_21519,N_23360);
nand UO_1721 (O_1721,N_20618,N_20343);
xor UO_1722 (O_1722,N_23297,N_23701);
or UO_1723 (O_1723,N_22727,N_23210);
and UO_1724 (O_1724,N_24370,N_21663);
xnor UO_1725 (O_1725,N_21100,N_20356);
and UO_1726 (O_1726,N_23294,N_22214);
xnor UO_1727 (O_1727,N_22241,N_23324);
and UO_1728 (O_1728,N_21462,N_24719);
nor UO_1729 (O_1729,N_20178,N_22204);
xnor UO_1730 (O_1730,N_24366,N_20084);
nor UO_1731 (O_1731,N_23907,N_24864);
or UO_1732 (O_1732,N_21472,N_21535);
xor UO_1733 (O_1733,N_20367,N_22867);
nor UO_1734 (O_1734,N_24135,N_21356);
and UO_1735 (O_1735,N_23403,N_22827);
nand UO_1736 (O_1736,N_20453,N_20611);
or UO_1737 (O_1737,N_24949,N_21487);
nor UO_1738 (O_1738,N_24645,N_20439);
or UO_1739 (O_1739,N_23090,N_22845);
and UO_1740 (O_1740,N_20392,N_22933);
xnor UO_1741 (O_1741,N_22044,N_21052);
and UO_1742 (O_1742,N_22305,N_24097);
nand UO_1743 (O_1743,N_21380,N_22689);
nand UO_1744 (O_1744,N_21528,N_23138);
nand UO_1745 (O_1745,N_22263,N_22012);
xor UO_1746 (O_1746,N_21752,N_22330);
nand UO_1747 (O_1747,N_21696,N_24670);
nand UO_1748 (O_1748,N_22654,N_21735);
nor UO_1749 (O_1749,N_21898,N_22424);
xor UO_1750 (O_1750,N_22721,N_21943);
and UO_1751 (O_1751,N_20707,N_21122);
nand UO_1752 (O_1752,N_22828,N_23504);
and UO_1753 (O_1753,N_20807,N_24679);
and UO_1754 (O_1754,N_21548,N_21089);
and UO_1755 (O_1755,N_23763,N_22961);
nor UO_1756 (O_1756,N_23072,N_23966);
nor UO_1757 (O_1757,N_20202,N_21787);
xor UO_1758 (O_1758,N_20714,N_24506);
or UO_1759 (O_1759,N_20575,N_21386);
and UO_1760 (O_1760,N_24060,N_21645);
nor UO_1761 (O_1761,N_22560,N_22607);
nand UO_1762 (O_1762,N_24541,N_22574);
xnor UO_1763 (O_1763,N_24542,N_20548);
xor UO_1764 (O_1764,N_24969,N_23598);
or UO_1765 (O_1765,N_22106,N_24570);
or UO_1766 (O_1766,N_24882,N_22265);
xnor UO_1767 (O_1767,N_20523,N_20647);
nand UO_1768 (O_1768,N_24180,N_24607);
or UO_1769 (O_1769,N_20990,N_20295);
xnor UO_1770 (O_1770,N_21265,N_24602);
xnor UO_1771 (O_1771,N_20694,N_23065);
nor UO_1772 (O_1772,N_21852,N_20034);
and UO_1773 (O_1773,N_20709,N_20235);
nand UO_1774 (O_1774,N_21479,N_20353);
xor UO_1775 (O_1775,N_20570,N_24524);
and UO_1776 (O_1776,N_22565,N_23932);
or UO_1777 (O_1777,N_22251,N_23654);
or UO_1778 (O_1778,N_24355,N_23100);
nand UO_1779 (O_1779,N_21458,N_22176);
and UO_1780 (O_1780,N_21242,N_21599);
nand UO_1781 (O_1781,N_24165,N_21002);
or UO_1782 (O_1782,N_24309,N_22624);
nand UO_1783 (O_1783,N_22309,N_21473);
nor UO_1784 (O_1784,N_20422,N_23787);
or UO_1785 (O_1785,N_21741,N_24928);
nand UO_1786 (O_1786,N_21492,N_24118);
nand UO_1787 (O_1787,N_22632,N_22152);
nor UO_1788 (O_1788,N_24930,N_22272);
nor UO_1789 (O_1789,N_22939,N_24763);
nand UO_1790 (O_1790,N_20556,N_22883);
or UO_1791 (O_1791,N_21368,N_23948);
xor UO_1792 (O_1792,N_21604,N_23178);
or UO_1793 (O_1793,N_24266,N_24260);
and UO_1794 (O_1794,N_24037,N_22453);
xor UO_1795 (O_1795,N_21075,N_21880);
and UO_1796 (O_1796,N_21792,N_22069);
and UO_1797 (O_1797,N_24881,N_24183);
or UO_1798 (O_1798,N_23990,N_23923);
or UO_1799 (O_1799,N_22483,N_24821);
xnor UO_1800 (O_1800,N_23120,N_23322);
nand UO_1801 (O_1801,N_20893,N_23435);
nand UO_1802 (O_1802,N_20687,N_20234);
nand UO_1803 (O_1803,N_24112,N_23373);
and UO_1804 (O_1804,N_23919,N_21069);
and UO_1805 (O_1805,N_24646,N_23319);
nand UO_1806 (O_1806,N_20991,N_22966);
xnor UO_1807 (O_1807,N_20799,N_23585);
xnor UO_1808 (O_1808,N_21514,N_24662);
nor UO_1809 (O_1809,N_23570,N_22379);
xnor UO_1810 (O_1810,N_21373,N_22054);
and UO_1811 (O_1811,N_20871,N_24286);
xnor UO_1812 (O_1812,N_21601,N_21134);
or UO_1813 (O_1813,N_22336,N_23698);
nand UO_1814 (O_1814,N_24721,N_24090);
and UO_1815 (O_1815,N_23443,N_20798);
and UO_1816 (O_1816,N_22800,N_21964);
nand UO_1817 (O_1817,N_24436,N_23544);
nand UO_1818 (O_1818,N_20304,N_20481);
or UO_1819 (O_1819,N_24363,N_24518);
nor UO_1820 (O_1820,N_20928,N_21825);
xor UO_1821 (O_1821,N_24834,N_20085);
or UO_1822 (O_1822,N_22715,N_23275);
nor UO_1823 (O_1823,N_20119,N_22590);
xor UO_1824 (O_1824,N_24665,N_22833);
nand UO_1825 (O_1825,N_22469,N_21412);
xnor UO_1826 (O_1826,N_20374,N_22923);
xnor UO_1827 (O_1827,N_23864,N_20585);
nor UO_1828 (O_1828,N_22353,N_23844);
or UO_1829 (O_1829,N_23260,N_20469);
and UO_1830 (O_1830,N_22652,N_22820);
or UO_1831 (O_1831,N_24664,N_24846);
or UO_1832 (O_1832,N_24899,N_23395);
nand UO_1833 (O_1833,N_21226,N_21580);
or UO_1834 (O_1834,N_24152,N_20851);
nor UO_1835 (O_1835,N_24549,N_21379);
nand UO_1836 (O_1836,N_21585,N_20776);
nor UO_1837 (O_1837,N_20616,N_23069);
xnor UO_1838 (O_1838,N_24649,N_21767);
xnor UO_1839 (O_1839,N_20738,N_20122);
nor UO_1840 (O_1840,N_24640,N_24350);
nand UO_1841 (O_1841,N_22473,N_21474);
nand UO_1842 (O_1842,N_20204,N_23061);
nand UO_1843 (O_1843,N_21054,N_20137);
nand UO_1844 (O_1844,N_20092,N_23821);
nand UO_1845 (O_1845,N_22516,N_23731);
xnor UO_1846 (O_1846,N_23149,N_20248);
and UO_1847 (O_1847,N_24398,N_23986);
nor UO_1848 (O_1848,N_22952,N_22279);
xor UO_1849 (O_1849,N_24865,N_22803);
or UO_1850 (O_1850,N_21337,N_24863);
or UO_1851 (O_1851,N_22675,N_23416);
or UO_1852 (O_1852,N_21499,N_22663);
or UO_1853 (O_1853,N_21193,N_22713);
nor UO_1854 (O_1854,N_23271,N_22147);
nor UO_1855 (O_1855,N_20289,N_23879);
nor UO_1856 (O_1856,N_21450,N_23234);
nand UO_1857 (O_1857,N_21452,N_24718);
nand UO_1858 (O_1858,N_20526,N_21813);
xnor UO_1859 (O_1859,N_21014,N_23920);
nor UO_1860 (O_1860,N_23583,N_23463);
nor UO_1861 (O_1861,N_20857,N_20164);
or UO_1862 (O_1862,N_24361,N_22325);
nand UO_1863 (O_1863,N_23546,N_21607);
and UO_1864 (O_1864,N_24529,N_20607);
nand UO_1865 (O_1865,N_21139,N_22814);
and UO_1866 (O_1866,N_20355,N_24823);
nor UO_1867 (O_1867,N_24544,N_24867);
nor UO_1868 (O_1868,N_24498,N_22850);
nor UO_1869 (O_1869,N_23622,N_24956);
nand UO_1870 (O_1870,N_24671,N_20380);
nor UO_1871 (O_1871,N_20550,N_21541);
and UO_1872 (O_1872,N_22334,N_24448);
or UO_1873 (O_1873,N_21210,N_24198);
or UO_1874 (O_1874,N_20465,N_24710);
nor UO_1875 (O_1875,N_21227,N_22725);
or UO_1876 (O_1876,N_22585,N_23335);
nand UO_1877 (O_1877,N_24178,N_24654);
nor UO_1878 (O_1878,N_23642,N_24109);
nand UO_1879 (O_1879,N_23280,N_21476);
nand UO_1880 (O_1880,N_23712,N_21928);
and UO_1881 (O_1881,N_22778,N_24722);
or UO_1882 (O_1882,N_23494,N_22105);
nand UO_1883 (O_1883,N_24455,N_24563);
nor UO_1884 (O_1884,N_24019,N_24047);
or UO_1885 (O_1885,N_23388,N_21327);
nand UO_1886 (O_1886,N_22608,N_21999);
and UO_1887 (O_1887,N_22520,N_24053);
nand UO_1888 (O_1888,N_23995,N_23479);
and UO_1889 (O_1889,N_22043,N_22941);
nor UO_1890 (O_1890,N_24847,N_23542);
or UO_1891 (O_1891,N_20094,N_24167);
or UO_1892 (O_1892,N_20933,N_22634);
nand UO_1893 (O_1893,N_20979,N_20197);
xnor UO_1894 (O_1894,N_21189,N_21391);
nand UO_1895 (O_1895,N_23645,N_23247);
nor UO_1896 (O_1896,N_20567,N_22244);
and UO_1897 (O_1897,N_21706,N_24358);
nand UO_1898 (O_1898,N_24031,N_23768);
nand UO_1899 (O_1899,N_22168,N_24736);
and UO_1900 (O_1900,N_24639,N_21022);
xor UO_1901 (O_1901,N_22912,N_21366);
and UO_1902 (O_1902,N_21629,N_21972);
and UO_1903 (O_1903,N_20501,N_20468);
nand UO_1904 (O_1904,N_24444,N_22446);
and UO_1905 (O_1905,N_23502,N_23428);
and UO_1906 (O_1906,N_20022,N_20340);
and UO_1907 (O_1907,N_21628,N_22613);
nor UO_1908 (O_1908,N_22036,N_22382);
or UO_1909 (O_1909,N_22979,N_22133);
and UO_1910 (O_1910,N_20964,N_23540);
nor UO_1911 (O_1911,N_24523,N_21344);
nor UO_1912 (O_1912,N_21142,N_24025);
xnor UO_1913 (O_1913,N_21441,N_23222);
and UO_1914 (O_1914,N_20766,N_21375);
or UO_1915 (O_1915,N_23916,N_20536);
nor UO_1916 (O_1916,N_21495,N_23361);
nand UO_1917 (O_1917,N_24612,N_21158);
and UO_1918 (O_1918,N_24986,N_24919);
xor UO_1919 (O_1919,N_20876,N_24780);
and UO_1920 (O_1920,N_24896,N_23312);
or UO_1921 (O_1921,N_23179,N_24095);
and UO_1922 (O_1922,N_24817,N_22097);
nor UO_1923 (O_1923,N_20788,N_20528);
nor UO_1924 (O_1924,N_21817,N_23870);
or UO_1925 (O_1925,N_21365,N_20282);
nor UO_1926 (O_1926,N_20609,N_20829);
and UO_1927 (O_1927,N_22977,N_24404);
or UO_1928 (O_1928,N_21530,N_24119);
xnor UO_1929 (O_1929,N_23267,N_20943);
xnor UO_1930 (O_1930,N_20081,N_24172);
and UO_1931 (O_1931,N_21723,N_22782);
nand UO_1932 (O_1932,N_24827,N_21564);
nand UO_1933 (O_1933,N_23808,N_23450);
nor UO_1934 (O_1934,N_23188,N_21155);
nand UO_1935 (O_1935,N_22422,N_20043);
and UO_1936 (O_1936,N_23669,N_21907);
xor UO_1937 (O_1937,N_23341,N_23735);
xnor UO_1938 (O_1938,N_20541,N_24296);
nand UO_1939 (O_1939,N_21268,N_24932);
nor UO_1940 (O_1940,N_20383,N_24725);
nor UO_1941 (O_1941,N_24164,N_23823);
xor UO_1942 (O_1942,N_20101,N_21233);
or UO_1943 (O_1943,N_22682,N_24276);
xnor UO_1944 (O_1944,N_23372,N_21364);
and UO_1945 (O_1945,N_22781,N_22490);
xor UO_1946 (O_1946,N_22728,N_20062);
xnor UO_1947 (O_1947,N_21129,N_21969);
nand UO_1948 (O_1948,N_20517,N_23129);
nand UO_1949 (O_1949,N_21801,N_24380);
nor UO_1950 (O_1950,N_24796,N_20892);
nand UO_1951 (O_1951,N_23587,N_20615);
nand UO_1952 (O_1952,N_23198,N_24788);
xnor UO_1953 (O_1953,N_21869,N_21486);
nor UO_1954 (O_1954,N_24218,N_24672);
or UO_1955 (O_1955,N_23582,N_20634);
xnor UO_1956 (O_1956,N_23902,N_23668);
or UO_1957 (O_1957,N_21512,N_20989);
and UO_1958 (O_1958,N_22079,N_20995);
or UO_1959 (O_1959,N_22524,N_23172);
nor UO_1960 (O_1960,N_23440,N_24776);
or UO_1961 (O_1961,N_21656,N_24862);
and UO_1962 (O_1962,N_24122,N_20148);
or UO_1963 (O_1963,N_20847,N_21820);
or UO_1964 (O_1964,N_23795,N_22666);
nor UO_1965 (O_1965,N_21329,N_22885);
nand UO_1966 (O_1966,N_24501,N_24892);
nand UO_1967 (O_1967,N_21998,N_21131);
or UO_1968 (O_1968,N_24289,N_24176);
xor UO_1969 (O_1969,N_22175,N_21935);
and UO_1970 (O_1970,N_24334,N_22948);
nor UO_1971 (O_1971,N_22208,N_23164);
xor UO_1972 (O_1972,N_22865,N_23962);
and UO_1973 (O_1973,N_23676,N_20819);
nor UO_1974 (O_1974,N_24724,N_20384);
nor UO_1975 (O_1975,N_22321,N_22050);
xor UO_1976 (O_1976,N_22783,N_20975);
and UO_1977 (O_1977,N_23726,N_24720);
and UO_1978 (O_1978,N_21853,N_23801);
xor UO_1979 (O_1979,N_24051,N_24958);
nand UO_1980 (O_1980,N_20167,N_20824);
and UO_1981 (O_1981,N_24294,N_21056);
xor UO_1982 (O_1982,N_21186,N_21757);
and UO_1983 (O_1983,N_20758,N_23561);
and UO_1984 (O_1984,N_20592,N_22899);
xnor UO_1985 (O_1985,N_23376,N_20795);
and UO_1986 (O_1986,N_22035,N_24925);
nand UO_1987 (O_1987,N_23268,N_21886);
nor UO_1988 (O_1988,N_22450,N_22222);
nor UO_1989 (O_1989,N_21531,N_20188);
nor UO_1990 (O_1990,N_23834,N_21841);
nor UO_1991 (O_1991,N_24951,N_21415);
xnor UO_1992 (O_1992,N_22207,N_21691);
and UO_1993 (O_1993,N_23264,N_20924);
or UO_1994 (O_1994,N_24099,N_21922);
or UO_1995 (O_1995,N_20147,N_23815);
nor UO_1996 (O_1996,N_20222,N_20828);
and UO_1997 (O_1997,N_21012,N_23277);
xor UO_1998 (O_1998,N_22932,N_23187);
nand UO_1999 (O_1999,N_20049,N_23174);
nor UO_2000 (O_2000,N_23856,N_21346);
or UO_2001 (O_2001,N_23556,N_22984);
nand UO_2002 (O_2002,N_22724,N_21537);
nand UO_2003 (O_2003,N_24974,N_23713);
xnor UO_2004 (O_2004,N_22695,N_24158);
xor UO_2005 (O_2005,N_23484,N_20619);
nand UO_2006 (O_2006,N_21705,N_22121);
nor UO_2007 (O_2007,N_24394,N_21676);
nand UO_2008 (O_2008,N_23140,N_21815);
nor UO_2009 (O_2009,N_22527,N_24650);
and UO_2010 (O_2010,N_20752,N_21334);
or UO_2011 (O_2011,N_22061,N_20217);
nor UO_2012 (O_2012,N_24116,N_22877);
or UO_2013 (O_2013,N_24488,N_22946);
xnor UO_2014 (O_2014,N_24756,N_24458);
nand UO_2015 (O_2015,N_22882,N_21881);
nand UO_2016 (O_2016,N_24571,N_23389);
nand UO_2017 (O_2017,N_20712,N_20260);
xnor UO_2018 (O_2018,N_22909,N_21400);
nand UO_2019 (O_2019,N_20562,N_21354);
nand UO_2020 (O_2020,N_20286,N_23767);
and UO_2021 (O_2021,N_20306,N_23290);
nor UO_2022 (O_2022,N_20859,N_21762);
or UO_2023 (O_2023,N_23937,N_24475);
nor UO_2024 (O_2024,N_24128,N_24717);
nor UO_2025 (O_2025,N_24487,N_23417);
and UO_2026 (O_2026,N_21533,N_23062);
nor UO_2027 (O_2027,N_22957,N_22922);
and UO_2028 (O_2028,N_20423,N_21251);
or UO_2029 (O_2029,N_20199,N_21238);
nor UO_2030 (O_2030,N_24950,N_24979);
nand UO_2031 (O_2031,N_23890,N_20003);
nand UO_2032 (O_2032,N_21445,N_23861);
xnor UO_2033 (O_2033,N_24561,N_22762);
nand UO_2034 (O_2034,N_21167,N_21689);
nand UO_2035 (O_2035,N_21084,N_20107);
and UO_2036 (O_2036,N_23070,N_24732);
or UO_2037 (O_2037,N_24532,N_24858);
nand UO_2038 (O_2038,N_22735,N_23437);
nor UO_2039 (O_2039,N_23910,N_22539);
nor UO_2040 (O_2040,N_23485,N_20108);
or UO_2041 (O_2041,N_22688,N_20631);
xor UO_2042 (O_2042,N_20952,N_22135);
nor UO_2043 (O_2043,N_22593,N_20586);
or UO_2044 (O_2044,N_24311,N_23771);
xor UO_2045 (O_2045,N_23385,N_21396);
or UO_2046 (O_2046,N_20456,N_24302);
xor UO_2047 (O_2047,N_21835,N_24134);
nor UO_2048 (O_2048,N_23147,N_24848);
nor UO_2049 (O_2049,N_20777,N_20868);
nand UO_2050 (O_2050,N_22059,N_22533);
xor UO_2051 (O_2051,N_24345,N_20869);
or UO_2052 (O_2052,N_20987,N_21309);
xor UO_2053 (O_2053,N_20571,N_20433);
and UO_2054 (O_2054,N_23215,N_21402);
xor UO_2055 (O_2055,N_22947,N_21508);
nor UO_2056 (O_2056,N_22374,N_20755);
or UO_2057 (O_2057,N_21498,N_23527);
nand UO_2058 (O_2058,N_20359,N_21433);
and UO_2059 (O_2059,N_23516,N_21627);
nand UO_2060 (O_2060,N_20373,N_24349);
nand UO_2061 (O_2061,N_22010,N_20138);
and UO_2062 (O_2062,N_22255,N_23697);
xor UO_2063 (O_2063,N_24298,N_23685);
nor UO_2064 (O_2064,N_21219,N_23653);
nand UO_2065 (O_2065,N_20993,N_23499);
and UO_2066 (O_2066,N_23829,N_22399);
and UO_2067 (O_2067,N_21112,N_24552);
xor UO_2068 (O_2068,N_21556,N_20736);
and UO_2069 (O_2069,N_23996,N_20444);
xor UO_2070 (O_2070,N_22234,N_23841);
xnor UO_2071 (O_2071,N_20568,N_21109);
xor UO_2072 (O_2072,N_22831,N_22823);
nor UO_2073 (O_2073,N_22813,N_21355);
or UO_2074 (O_2074,N_21558,N_22454);
nor UO_2075 (O_2075,N_21532,N_24274);
and UO_2076 (O_2076,N_24070,N_22448);
or UO_2077 (O_2077,N_23558,N_24052);
nand UO_2078 (O_2078,N_24421,N_22210);
xor UO_2079 (O_2079,N_23097,N_21753);
or UO_2080 (O_2080,N_20806,N_23670);
nor UO_2081 (O_2081,N_24046,N_23959);
nor UO_2082 (O_2082,N_22571,N_23157);
nand UO_2083 (O_2083,N_23889,N_22579);
or UO_2084 (O_2084,N_21281,N_22944);
xnor UO_2085 (O_2085,N_21756,N_21258);
and UO_2086 (O_2086,N_21652,N_21894);
or UO_2087 (O_2087,N_21339,N_20215);
nor UO_2088 (O_2088,N_20098,N_23303);
and UO_2089 (O_2089,N_23756,N_20035);
and UO_2090 (O_2090,N_21101,N_20679);
nor UO_2091 (O_2091,N_22841,N_22518);
or UO_2092 (O_2092,N_20699,N_24018);
nor UO_2093 (O_2093,N_21714,N_23046);
and UO_2094 (O_2094,N_23262,N_24215);
nand UO_2095 (O_2095,N_23613,N_21718);
xnor UO_2096 (O_2096,N_24816,N_20855);
and UO_2097 (O_2097,N_22905,N_20302);
nand UO_2098 (O_2098,N_22599,N_22926);
and UO_2099 (O_2099,N_21203,N_21127);
and UO_2100 (O_2100,N_23039,N_20314);
nand UO_2101 (O_2101,N_22596,N_22328);
nand UO_2102 (O_2102,N_24884,N_24375);
nand UO_2103 (O_2103,N_22670,N_24240);
and UO_2104 (O_2104,N_23730,N_23316);
xor UO_2105 (O_2105,N_22581,N_22434);
nand UO_2106 (O_2106,N_21493,N_24362);
xor UO_2107 (O_2107,N_22360,N_22389);
and UO_2108 (O_2108,N_24868,N_24923);
or UO_2109 (O_2109,N_24023,N_24556);
xor UO_2110 (O_2110,N_24413,N_23847);
xnor UO_2111 (O_2111,N_24387,N_20209);
nand UO_2112 (O_2112,N_21123,N_23451);
or UO_2113 (O_2113,N_21435,N_21032);
or UO_2114 (O_2114,N_21818,N_21135);
nand UO_2115 (O_2115,N_23930,N_22489);
nand UO_2116 (O_2116,N_22060,N_22127);
nor UO_2117 (O_2117,N_23383,N_24182);
xor UO_2118 (O_2118,N_23345,N_24454);
and UO_2119 (O_2119,N_20061,N_20381);
and UO_2120 (O_2120,N_22779,N_23511);
and UO_2121 (O_2121,N_21204,N_23684);
and UO_2122 (O_2122,N_24917,N_23263);
nor UO_2123 (O_2123,N_24209,N_23196);
or UO_2124 (O_2124,N_24712,N_20817);
xor UO_2125 (O_2125,N_24713,N_24043);
xor UO_2126 (O_2126,N_20288,N_20565);
nand UO_2127 (O_2127,N_24779,N_21438);
nand UO_2128 (O_2128,N_20992,N_22749);
nor UO_2129 (O_2129,N_24857,N_24975);
and UO_2130 (O_2130,N_24310,N_21263);
and UO_2131 (O_2131,N_21669,N_23425);
nand UO_2132 (O_2132,N_20998,N_22037);
nor UO_2133 (O_2133,N_20259,N_20711);
xnor UO_2134 (O_2134,N_21877,N_23382);
nand UO_2135 (O_2135,N_22917,N_20591);
nor UO_2136 (O_2136,N_24547,N_22217);
xor UO_2137 (O_2137,N_22154,N_21040);
nand UO_2138 (O_2138,N_22363,N_22526);
or UO_2139 (O_2139,N_23775,N_21223);
xor UO_2140 (O_2140,N_21793,N_20120);
or UO_2141 (O_2141,N_23682,N_21156);
or UO_2142 (O_2142,N_23602,N_24906);
xnor UO_2143 (O_2143,N_24676,N_22232);
and UO_2144 (O_2144,N_24627,N_20622);
nand UO_2145 (O_2145,N_20513,N_24219);
xor UO_2146 (O_2146,N_23860,N_21587);
nand UO_2147 (O_2147,N_23537,N_23800);
and UO_2148 (O_2148,N_20633,N_22364);
nand UO_2149 (O_2149,N_21345,N_22739);
or UO_2150 (O_2150,N_24636,N_20985);
or UO_2151 (O_2151,N_22445,N_23348);
and UO_2152 (O_2152,N_23064,N_23777);
nand UO_2153 (O_2153,N_24439,N_23780);
and UO_2154 (O_2154,N_24686,N_22057);
xor UO_2155 (O_2155,N_22381,N_24677);
or UO_2156 (O_2156,N_21933,N_21185);
nand UO_2157 (O_2157,N_20152,N_20852);
nor UO_2158 (O_2158,N_22641,N_23023);
nor UO_2159 (O_2159,N_21692,N_22064);
or UO_2160 (O_2160,N_23983,N_22536);
and UO_2161 (O_2161,N_23343,N_22890);
xor UO_2162 (O_2162,N_22618,N_20390);
nor UO_2163 (O_2163,N_21545,N_20579);
and UO_2164 (O_2164,N_20519,N_23327);
or UO_2165 (O_2165,N_20743,N_22122);
and UO_2166 (O_2166,N_22242,N_24830);
and UO_2167 (O_2167,N_22718,N_23083);
nor UO_2168 (O_2168,N_23413,N_20179);
xor UO_2169 (O_2169,N_21678,N_24760);
xor UO_2170 (O_2170,N_20403,N_24550);
or UO_2171 (O_2171,N_22830,N_22753);
xnor UO_2172 (O_2172,N_22359,N_23228);
nand UO_2173 (O_2173,N_21967,N_24068);
nor UO_2174 (O_2174,N_23318,N_24510);
or UO_2175 (O_2175,N_24871,N_21878);
or UO_2176 (O_2176,N_24705,N_23596);
and UO_2177 (O_2177,N_21315,N_21005);
or UO_2178 (O_2178,N_24918,N_22921);
or UO_2179 (O_2179,N_22118,N_20974);
nor UO_2180 (O_2180,N_22981,N_24987);
and UO_2181 (O_2181,N_20842,N_21298);
xor UO_2182 (O_2182,N_20617,N_23214);
xnor UO_2183 (O_2183,N_23914,N_24157);
and UO_2184 (O_2184,N_24446,N_23026);
nand UO_2185 (O_2185,N_20024,N_23177);
and UO_2186 (O_2186,N_22983,N_22622);
nand UO_2187 (O_2187,N_20546,N_23892);
nor UO_2188 (O_2188,N_21583,N_23049);
xor UO_2189 (O_2189,N_20112,N_24381);
nand UO_2190 (O_2190,N_20157,N_22597);
and UO_2191 (O_2191,N_23854,N_22306);
and UO_2192 (O_2192,N_21034,N_20790);
nand UO_2193 (O_2193,N_20205,N_21874);
and UO_2194 (O_2194,N_20906,N_20113);
xor UO_2195 (O_2195,N_24569,N_20130);
xnor UO_2196 (O_2196,N_20405,N_22548);
nand UO_2197 (O_2197,N_20596,N_23954);
xnor UO_2198 (O_2198,N_20903,N_22386);
and UO_2199 (O_2199,N_21046,N_22319);
nand UO_2200 (O_2200,N_21662,N_21630);
nand UO_2201 (O_2201,N_23674,N_22644);
and UO_2202 (O_2202,N_22257,N_22843);
nor UO_2203 (O_2203,N_21522,N_22569);
and UO_2204 (O_2204,N_22937,N_23640);
xor UO_2205 (O_2205,N_20698,N_24888);
nand UO_2206 (O_2206,N_23658,N_20834);
or UO_2207 (O_2207,N_20226,N_21200);
nand UO_2208 (O_2208,N_20746,N_22717);
and UO_2209 (O_2209,N_24000,N_21785);
xnor UO_2210 (O_2210,N_21230,N_21293);
xor UO_2211 (O_2211,N_24666,N_20626);
xor UO_2212 (O_2212,N_20389,N_21802);
xnor UO_2213 (O_2213,N_23530,N_23219);
nor UO_2214 (O_2214,N_21440,N_23226);
nand UO_2215 (O_2215,N_23576,N_24669);
nand UO_2216 (O_2216,N_21695,N_20488);
nor UO_2217 (O_2217,N_23154,N_22166);
nand UO_2218 (O_2218,N_22529,N_22602);
nor UO_2219 (O_2219,N_22298,N_23139);
nand UO_2220 (O_2220,N_23252,N_21539);
nand UO_2221 (O_2221,N_23538,N_21237);
or UO_2222 (O_2222,N_23159,N_21806);
nor UO_2223 (O_2223,N_24197,N_24620);
nand UO_2224 (O_2224,N_20479,N_24199);
and UO_2225 (O_2225,N_20253,N_21791);
and UO_2226 (O_2226,N_20458,N_21456);
xnor UO_2227 (O_2227,N_24521,N_23477);
and UO_2228 (O_2228,N_23991,N_24194);
nand UO_2229 (O_2229,N_20744,N_21042);
nor UO_2230 (O_2230,N_23604,N_21810);
xor UO_2231 (O_2231,N_22908,N_20838);
nor UO_2232 (O_2232,N_24123,N_22502);
and UO_2233 (O_2233,N_22510,N_24297);
or UO_2234 (O_2234,N_23751,N_20861);
nor UO_2235 (O_2235,N_22285,N_24623);
or UO_2236 (O_2236,N_20832,N_20720);
nor UO_2237 (O_2237,N_22046,N_22636);
nor UO_2238 (O_2238,N_21882,N_23112);
xnor UO_2239 (O_2239,N_21827,N_20328);
xnor UO_2240 (O_2240,N_24885,N_24385);
and UO_2241 (O_2241,N_24465,N_20725);
and UO_2242 (O_2242,N_24305,N_22701);
or UO_2243 (O_2243,N_22982,N_20664);
nand UO_2244 (O_2244,N_21018,N_20391);
or UO_2245 (O_2245,N_22115,N_24684);
nor UO_2246 (O_2246,N_24024,N_23784);
nand UO_2247 (O_2247,N_20066,N_24746);
nor UO_2248 (O_2248,N_22528,N_21138);
and UO_2249 (O_2249,N_21800,N_22439);
and UO_2250 (O_2250,N_21029,N_22355);
nor UO_2251 (O_2251,N_20630,N_24574);
or UO_2252 (O_2252,N_24424,N_21036);
and UO_2253 (O_2253,N_21403,N_20494);
xor UO_2254 (O_2254,N_23397,N_23968);
nor UO_2255 (O_2255,N_23789,N_24814);
nand UO_2256 (O_2256,N_22405,N_23077);
or UO_2257 (O_2257,N_23209,N_24997);
xnor UO_2258 (O_2258,N_21197,N_24739);
nor UO_2259 (O_2259,N_21947,N_24405);
nor UO_2260 (O_2260,N_23779,N_21540);
and UO_2261 (O_2261,N_22391,N_23305);
nor UO_2262 (O_2262,N_22093,N_21620);
or UO_2263 (O_2263,N_22153,N_21589);
or UO_2264 (O_2264,N_20573,N_23008);
nor UO_2265 (O_2265,N_23370,N_20225);
xnor UO_2266 (O_2266,N_21269,N_23630);
nand UO_2267 (O_2267,N_20316,N_24852);
nor UO_2268 (O_2268,N_24690,N_24784);
nand UO_2269 (O_2269,N_23186,N_23908);
and UO_2270 (O_2270,N_22343,N_20153);
nor UO_2271 (O_2271,N_24901,N_23551);
and UO_2272 (O_2272,N_22027,N_22167);
and UO_2273 (O_2273,N_23673,N_22591);
or UO_2274 (O_2274,N_21918,N_23518);
xnor UO_2275 (O_2275,N_24406,N_20118);
or UO_2276 (O_2276,N_24203,N_21635);
nor UO_2277 (O_2277,N_22791,N_24913);
nand UO_2278 (O_2278,N_23040,N_24912);
and UO_2279 (O_2279,N_23400,N_24093);
or UO_2280 (O_2280,N_22542,N_22505);
xnor UO_2281 (O_2281,N_24267,N_20487);
and UO_2282 (O_2282,N_22250,N_23791);
xnor UO_2283 (O_2283,N_24678,N_23095);
nand UO_2284 (O_2284,N_23760,N_23163);
nor UO_2285 (O_2285,N_21003,N_20223);
and UO_2286 (O_2286,N_23068,N_24486);
or UO_2287 (O_2287,N_21568,N_23092);
and UO_2288 (O_2288,N_20830,N_20020);
or UO_2289 (O_2289,N_22665,N_22468);
xor UO_2290 (O_2290,N_22792,N_21919);
and UO_2291 (O_2291,N_22327,N_24903);
xor UO_2292 (O_2292,N_24813,N_24820);
xnor UO_2293 (O_2293,N_24957,N_22014);
or UO_2294 (O_2294,N_21505,N_23941);
and UO_2295 (O_2295,N_23158,N_22508);
and UO_2296 (O_2296,N_21287,N_20364);
xnor UO_2297 (O_2297,N_21975,N_23543);
nor UO_2298 (O_2298,N_22859,N_21763);
nand UO_2299 (O_2299,N_21702,N_20520);
or UO_2300 (O_2300,N_23104,N_20203);
or UO_2301 (O_2301,N_21092,N_24810);
or UO_2302 (O_2302,N_20496,N_21945);
and UO_2303 (O_2303,N_23476,N_23058);
and UO_2304 (O_2304,N_22000,N_24452);
or UO_2305 (O_2305,N_22789,N_22964);
and UO_2306 (O_2306,N_21385,N_20297);
nor UO_2307 (O_2307,N_24594,N_23836);
nor UO_2308 (O_2308,N_23036,N_22021);
nand UO_2309 (O_2309,N_24894,N_20597);
nor UO_2310 (O_2310,N_24174,N_23094);
nor UO_2311 (O_2311,N_24146,N_22104);
or UO_2312 (O_2312,N_20808,N_20079);
nand UO_2313 (O_2313,N_24114,N_24034);
xnor UO_2314 (O_2314,N_20542,N_22269);
nand UO_2315 (O_2315,N_20996,N_22013);
nor UO_2316 (O_2316,N_22380,N_20826);
and UO_2317 (O_2317,N_22004,N_21490);
or UO_2318 (O_2318,N_22878,N_23191);
nor UO_2319 (O_2319,N_24166,N_23239);
xnor UO_2320 (O_2320,N_20186,N_20070);
nand UO_2321 (O_2321,N_23637,N_23180);
nor UO_2322 (O_2322,N_22333,N_24735);
and UO_2323 (O_2323,N_24886,N_23166);
xor UO_2324 (O_2324,N_23017,N_21956);
nor UO_2325 (O_2325,N_24121,N_20638);
nand UO_2326 (O_2326,N_24101,N_24435);
and UO_2327 (O_2327,N_20929,N_21730);
nand UO_2328 (O_2328,N_24505,N_20060);
and UO_2329 (O_2329,N_21343,N_23628);
and UO_2330 (O_2330,N_20474,N_24539);
and UO_2331 (O_2331,N_22886,N_24020);
xor UO_2332 (O_2332,N_20347,N_22653);
nor UO_2333 (O_2333,N_21328,N_23028);
nand UO_2334 (O_2334,N_21316,N_24965);
nor UO_2335 (O_2335,N_24781,N_22851);
or UO_2336 (O_2336,N_20581,N_20953);
nor UO_2337 (O_2337,N_24904,N_21944);
nand UO_2338 (O_2338,N_20348,N_21363);
nand UO_2339 (O_2339,N_23224,N_20394);
nor UO_2340 (O_2340,N_24980,N_24282);
or UO_2341 (O_2341,N_23043,N_22225);
nor UO_2342 (O_2342,N_20262,N_23142);
xnor UO_2343 (O_2343,N_23006,N_21255);
xor UO_2344 (O_2344,N_24692,N_24306);
xor UO_2345 (O_2345,N_21196,N_21148);
or UO_2346 (O_2346,N_23769,N_22668);
or UO_2347 (O_2347,N_24071,N_20867);
and UO_2348 (O_2348,N_22356,N_24818);
or UO_2349 (O_2349,N_20984,N_23128);
and UO_2350 (O_2350,N_22401,N_21626);
nor UO_2351 (O_2351,N_22504,N_24740);
and UO_2352 (O_2352,N_22761,N_23331);
nor UO_2353 (O_2353,N_22821,N_21431);
or UO_2354 (O_2354,N_20228,N_24186);
nand UO_2355 (O_2355,N_24828,N_22462);
nor UO_2356 (O_2356,N_24352,N_23672);
nor UO_2357 (O_2357,N_23714,N_22034);
xnor UO_2358 (O_2358,N_22931,N_20879);
nand UO_2359 (O_2359,N_24519,N_23362);
nor UO_2360 (O_2360,N_21461,N_20844);
nor UO_2361 (O_2361,N_24299,N_24181);
and UO_2362 (O_2362,N_22111,N_23707);
or UO_2363 (O_2363,N_20145,N_20770);
or UO_2364 (O_2364,N_23269,N_23873);
and UO_2365 (O_2365,N_22003,N_23381);
or UO_2366 (O_2366,N_23589,N_20187);
nor UO_2367 (O_2367,N_24320,N_23141);
and UO_2368 (O_2368,N_22101,N_20782);
nand UO_2369 (O_2369,N_22110,N_22980);
and UO_2370 (O_2370,N_24555,N_22378);
xor UO_2371 (O_2371,N_21360,N_24726);
nand UO_2372 (O_2372,N_24130,N_21171);
nor UO_2373 (O_2373,N_23545,N_21145);
nand UO_2374 (O_2374,N_24026,N_21121);
nor UO_2375 (O_2375,N_22995,N_22100);
nor UO_2376 (O_2376,N_21980,N_23321);
nor UO_2377 (O_2377,N_24005,N_22368);
nor UO_2378 (O_2378,N_20671,N_20734);
nor UO_2379 (O_2379,N_22645,N_20331);
xnor UO_2380 (O_2380,N_21083,N_22407);
nand UO_2381 (O_2381,N_20846,N_22190);
nand UO_2382 (O_2382,N_24591,N_21598);
or UO_2383 (O_2383,N_20044,N_21860);
nand UO_2384 (O_2384,N_21150,N_21804);
and UO_2385 (O_2385,N_22756,N_21819);
or UO_2386 (O_2386,N_22648,N_22551);
xnor UO_2387 (O_2387,N_20115,N_24143);
or UO_2388 (O_2388,N_23408,N_24526);
xnor UO_2389 (O_2389,N_20249,N_22308);
and UO_2390 (O_2390,N_24696,N_24916);
nor UO_2391 (O_2391,N_23367,N_24515);
nand UO_2392 (O_2392,N_23117,N_24704);
nand UO_2393 (O_2393,N_22108,N_23087);
xnor UO_2394 (O_2394,N_23619,N_21168);
nor UO_2395 (O_2395,N_23055,N_23624);
xnor UO_2396 (O_2396,N_23595,N_22986);
or UO_2397 (O_2397,N_22002,N_20459);
nor UO_2398 (O_2398,N_21215,N_21845);
nand UO_2399 (O_2399,N_24461,N_23495);
or UO_2400 (O_2400,N_24295,N_22967);
and UO_2401 (O_2401,N_21655,N_20072);
or UO_2402 (O_2402,N_21401,N_21394);
nand UO_2403 (O_2403,N_20133,N_24626);
nand UO_2404 (O_2404,N_23786,N_23465);
nor UO_2405 (O_2405,N_23950,N_23519);
or UO_2406 (O_2406,N_24236,N_24377);
or UO_2407 (O_2407,N_24033,N_22630);
or UO_2408 (O_2408,N_22130,N_23071);
xor UO_2409 (O_2409,N_20395,N_20012);
or UO_2410 (O_2410,N_23356,N_21617);
nand UO_2411 (O_2411,N_23161,N_24407);
and UO_2412 (O_2412,N_22875,N_20497);
nand UO_2413 (O_2413,N_24554,N_24534);
nor UO_2414 (O_2414,N_24089,N_21949);
xor UO_2415 (O_2415,N_20748,N_21273);
nor UO_2416 (O_2416,N_22692,N_22545);
nor UO_2417 (O_2417,N_21236,N_20610);
nand UO_2418 (O_2418,N_20822,N_22868);
nand UO_2419 (O_2419,N_23649,N_23257);
or UO_2420 (O_2420,N_20418,N_23671);
and UO_2421 (O_2421,N_20499,N_21970);
nand UO_2422 (O_2422,N_24227,N_24265);
xor UO_2423 (O_2423,N_24175,N_21047);
or UO_2424 (O_2424,N_20841,N_20411);
nor UO_2425 (O_2425,N_24673,N_21133);
and UO_2426 (O_2426,N_24307,N_20067);
or UO_2427 (O_2427,N_23752,N_22174);
xnor UO_2428 (O_2428,N_24741,N_20478);
nand UO_2429 (O_2429,N_23603,N_21901);
and UO_2430 (O_2430,N_20156,N_22430);
or UO_2431 (O_2431,N_20172,N_22409);
xor UO_2432 (O_2432,N_20464,N_22178);
or UO_2433 (O_2433,N_20116,N_23677);
xor UO_2434 (O_2434,N_22699,N_21739);
xnor UO_2435 (O_2435,N_24360,N_20898);
and UO_2436 (O_2436,N_20051,N_22902);
or UO_2437 (O_2437,N_22464,N_22194);
xor UO_2438 (O_2438,N_23681,N_21081);
or UO_2439 (O_2439,N_24242,N_20140);
nor UO_2440 (O_2440,N_24062,N_21497);
xnor UO_2441 (O_2441,N_21469,N_20252);
nor UO_2442 (O_2442,N_21962,N_20099);
nand UO_2443 (O_2443,N_23565,N_22197);
nand UO_2444 (O_2444,N_20310,N_24015);
nand UO_2445 (O_2445,N_21173,N_23279);
nand UO_2446 (O_2446,N_24103,N_20780);
or UO_2447 (O_2447,N_22532,N_23302);
xor UO_2448 (O_2448,N_24631,N_22611);
nor UO_2449 (O_2449,N_21831,N_20922);
and UO_2450 (O_2450,N_24583,N_24391);
nand UO_2451 (O_2451,N_20997,N_20175);
nor UO_2452 (O_2452,N_20713,N_21814);
xnor UO_2453 (O_2453,N_20986,N_21647);
nand UO_2454 (O_2454,N_22169,N_24467);
nor UO_2455 (O_2455,N_22277,N_22893);
nand UO_2456 (O_2456,N_22785,N_21697);
nand UO_2457 (O_2457,N_21875,N_20775);
nor UO_2458 (O_2458,N_21453,N_23825);
xnor UO_2459 (O_2459,N_22846,N_24317);
or UO_2460 (O_2460,N_21132,N_24749);
nor UO_2461 (O_2461,N_22633,N_24619);
nor UO_2462 (O_2462,N_22254,N_21660);
and UO_2463 (O_2463,N_22712,N_24082);
nor UO_2464 (O_2464,N_24651,N_20181);
xor UO_2465 (O_2465,N_23016,N_22647);
xor UO_2466 (O_2466,N_20333,N_20220);
nor UO_2467 (O_2467,N_20818,N_24463);
xnor UO_2468 (O_2468,N_24866,N_23338);
nand UO_2469 (O_2469,N_20500,N_22408);
nand UO_2470 (O_2470,N_24129,N_21870);
nand UO_2471 (O_2471,N_24644,N_20185);
xor UO_2472 (O_2472,N_24249,N_23113);
xnor UO_2473 (O_2473,N_23508,N_23727);
xnor UO_2474 (O_2474,N_20166,N_23597);
or UO_2475 (O_2475,N_21303,N_22940);
and UO_2476 (O_2476,N_23774,N_22733);
nand UO_2477 (O_2477,N_22117,N_20502);
nor UO_2478 (O_2478,N_21066,N_20064);
nor UO_2479 (O_2479,N_23796,N_23702);
and UO_2480 (O_2480,N_22270,N_21782);
nand UO_2481 (O_2481,N_22261,N_23486);
xor UO_2482 (O_2482,N_24893,N_24437);
and UO_2483 (O_2483,N_20666,N_21914);
xnor UO_2484 (O_2484,N_21618,N_23819);
and UO_2485 (O_2485,N_20835,N_21175);
and UO_2486 (O_2486,N_22200,N_23102);
or UO_2487 (O_2487,N_20642,N_23171);
nand UO_2488 (O_2488,N_24798,N_20724);
nor UO_2489 (O_2489,N_21096,N_23060);
nand UO_2490 (O_2490,N_20754,N_22080);
xor UO_2491 (O_2491,N_21060,N_24537);
xor UO_2492 (O_2492,N_21971,N_24592);
xor UO_2493 (O_2493,N_23896,N_20104);
nor UO_2494 (O_2494,N_20580,N_22892);
or UO_2495 (O_2495,N_21862,N_23863);
nand UO_2496 (O_2496,N_20593,N_22164);
nor UO_2497 (O_2497,N_20506,N_24430);
nand UO_2498 (O_2498,N_24766,N_21844);
xnor UO_2499 (O_2499,N_20951,N_23579);
and UO_2500 (O_2500,N_22091,N_20405);
and UO_2501 (O_2501,N_24265,N_21096);
nand UO_2502 (O_2502,N_21388,N_23863);
and UO_2503 (O_2503,N_22647,N_24518);
nor UO_2504 (O_2504,N_24222,N_20217);
xnor UO_2505 (O_2505,N_24038,N_20516);
and UO_2506 (O_2506,N_24960,N_24408);
xnor UO_2507 (O_2507,N_21545,N_22304);
xor UO_2508 (O_2508,N_23618,N_24186);
xnor UO_2509 (O_2509,N_22073,N_22815);
and UO_2510 (O_2510,N_21238,N_22951);
and UO_2511 (O_2511,N_23965,N_24983);
nand UO_2512 (O_2512,N_24524,N_22941);
nand UO_2513 (O_2513,N_22329,N_24533);
nor UO_2514 (O_2514,N_21745,N_23719);
or UO_2515 (O_2515,N_21747,N_20221);
xor UO_2516 (O_2516,N_22617,N_22114);
nand UO_2517 (O_2517,N_23422,N_20302);
nor UO_2518 (O_2518,N_21142,N_24726);
and UO_2519 (O_2519,N_24422,N_24023);
nor UO_2520 (O_2520,N_20103,N_24642);
nand UO_2521 (O_2521,N_22012,N_21338);
or UO_2522 (O_2522,N_22117,N_23272);
and UO_2523 (O_2523,N_24102,N_24459);
nor UO_2524 (O_2524,N_20806,N_22657);
and UO_2525 (O_2525,N_24085,N_23165);
or UO_2526 (O_2526,N_22235,N_24136);
or UO_2527 (O_2527,N_20034,N_23828);
xnor UO_2528 (O_2528,N_22667,N_21833);
and UO_2529 (O_2529,N_20586,N_21863);
nand UO_2530 (O_2530,N_20533,N_22566);
nor UO_2531 (O_2531,N_23894,N_20271);
xnor UO_2532 (O_2532,N_24105,N_23633);
nand UO_2533 (O_2533,N_23161,N_21901);
or UO_2534 (O_2534,N_23441,N_21300);
and UO_2535 (O_2535,N_22648,N_20342);
and UO_2536 (O_2536,N_22902,N_22227);
nand UO_2537 (O_2537,N_20584,N_21285);
xnor UO_2538 (O_2538,N_21121,N_22778);
and UO_2539 (O_2539,N_20303,N_20817);
nor UO_2540 (O_2540,N_24492,N_23448);
nor UO_2541 (O_2541,N_21339,N_22859);
and UO_2542 (O_2542,N_20692,N_23329);
nand UO_2543 (O_2543,N_21402,N_22423);
xor UO_2544 (O_2544,N_24723,N_24380);
nand UO_2545 (O_2545,N_20236,N_20850);
nor UO_2546 (O_2546,N_21566,N_23953);
nand UO_2547 (O_2547,N_20242,N_22513);
or UO_2548 (O_2548,N_21397,N_23849);
xor UO_2549 (O_2549,N_20426,N_21384);
nand UO_2550 (O_2550,N_20951,N_21471);
nand UO_2551 (O_2551,N_21481,N_24584);
nor UO_2552 (O_2552,N_21730,N_23018);
nand UO_2553 (O_2553,N_22086,N_22608);
nand UO_2554 (O_2554,N_24603,N_22584);
nand UO_2555 (O_2555,N_21037,N_22608);
xor UO_2556 (O_2556,N_23371,N_21382);
and UO_2557 (O_2557,N_22029,N_20351);
and UO_2558 (O_2558,N_21916,N_20195);
xor UO_2559 (O_2559,N_21503,N_23962);
or UO_2560 (O_2560,N_20315,N_20255);
and UO_2561 (O_2561,N_23894,N_23020);
and UO_2562 (O_2562,N_21851,N_24966);
nand UO_2563 (O_2563,N_22914,N_24517);
nor UO_2564 (O_2564,N_22371,N_24644);
or UO_2565 (O_2565,N_22875,N_23715);
nor UO_2566 (O_2566,N_21855,N_22297);
or UO_2567 (O_2567,N_23592,N_22727);
xnor UO_2568 (O_2568,N_23413,N_20327);
nor UO_2569 (O_2569,N_23833,N_22628);
xor UO_2570 (O_2570,N_24378,N_20997);
nor UO_2571 (O_2571,N_24627,N_23863);
xor UO_2572 (O_2572,N_24208,N_23579);
or UO_2573 (O_2573,N_23298,N_20370);
or UO_2574 (O_2574,N_22218,N_24973);
nand UO_2575 (O_2575,N_24730,N_24045);
xor UO_2576 (O_2576,N_24502,N_22249);
and UO_2577 (O_2577,N_24148,N_21316);
nor UO_2578 (O_2578,N_21211,N_24515);
nand UO_2579 (O_2579,N_23852,N_22910);
nand UO_2580 (O_2580,N_20541,N_20720);
xnor UO_2581 (O_2581,N_21700,N_22327);
nand UO_2582 (O_2582,N_21529,N_23009);
and UO_2583 (O_2583,N_24470,N_24738);
nand UO_2584 (O_2584,N_23590,N_23176);
or UO_2585 (O_2585,N_21273,N_24415);
nor UO_2586 (O_2586,N_21966,N_24781);
and UO_2587 (O_2587,N_20722,N_23103);
xor UO_2588 (O_2588,N_20519,N_20665);
and UO_2589 (O_2589,N_21777,N_20302);
or UO_2590 (O_2590,N_24627,N_20816);
and UO_2591 (O_2591,N_22381,N_22802);
and UO_2592 (O_2592,N_24259,N_24567);
nor UO_2593 (O_2593,N_20304,N_23493);
and UO_2594 (O_2594,N_21448,N_21528);
xor UO_2595 (O_2595,N_21835,N_24621);
nand UO_2596 (O_2596,N_22511,N_22071);
nand UO_2597 (O_2597,N_20567,N_20975);
or UO_2598 (O_2598,N_22689,N_22123);
nand UO_2599 (O_2599,N_23629,N_21228);
xnor UO_2600 (O_2600,N_20162,N_23745);
xnor UO_2601 (O_2601,N_20496,N_22989);
or UO_2602 (O_2602,N_24047,N_23240);
and UO_2603 (O_2603,N_24551,N_20045);
xnor UO_2604 (O_2604,N_21887,N_22088);
nand UO_2605 (O_2605,N_20917,N_21921);
xor UO_2606 (O_2606,N_20808,N_23212);
and UO_2607 (O_2607,N_22057,N_21455);
nand UO_2608 (O_2608,N_20777,N_22008);
nand UO_2609 (O_2609,N_24161,N_21616);
nand UO_2610 (O_2610,N_21393,N_20537);
nor UO_2611 (O_2611,N_24965,N_24430);
nand UO_2612 (O_2612,N_22101,N_24998);
and UO_2613 (O_2613,N_21047,N_24315);
or UO_2614 (O_2614,N_20154,N_22299);
nor UO_2615 (O_2615,N_22628,N_23456);
or UO_2616 (O_2616,N_22779,N_20467);
nand UO_2617 (O_2617,N_20461,N_24166);
and UO_2618 (O_2618,N_24904,N_21536);
nand UO_2619 (O_2619,N_20358,N_22410);
or UO_2620 (O_2620,N_20675,N_20878);
nor UO_2621 (O_2621,N_23395,N_24249);
nor UO_2622 (O_2622,N_22072,N_20217);
nand UO_2623 (O_2623,N_20778,N_20387);
nand UO_2624 (O_2624,N_21731,N_21545);
and UO_2625 (O_2625,N_20237,N_24483);
xnor UO_2626 (O_2626,N_23795,N_24963);
xnor UO_2627 (O_2627,N_21439,N_23325);
and UO_2628 (O_2628,N_20525,N_23616);
nand UO_2629 (O_2629,N_23749,N_21435);
and UO_2630 (O_2630,N_20935,N_24298);
and UO_2631 (O_2631,N_21432,N_20126);
xnor UO_2632 (O_2632,N_22326,N_23773);
nand UO_2633 (O_2633,N_24388,N_22385);
xor UO_2634 (O_2634,N_21112,N_23729);
or UO_2635 (O_2635,N_21960,N_24334);
xor UO_2636 (O_2636,N_24233,N_24986);
and UO_2637 (O_2637,N_21881,N_22130);
and UO_2638 (O_2638,N_20729,N_22301);
nor UO_2639 (O_2639,N_20283,N_20534);
nor UO_2640 (O_2640,N_23373,N_20735);
or UO_2641 (O_2641,N_22732,N_23372);
or UO_2642 (O_2642,N_23339,N_24819);
and UO_2643 (O_2643,N_24860,N_24310);
nand UO_2644 (O_2644,N_21085,N_24377);
or UO_2645 (O_2645,N_23591,N_22055);
or UO_2646 (O_2646,N_21460,N_23980);
and UO_2647 (O_2647,N_20025,N_24722);
xor UO_2648 (O_2648,N_23286,N_21025);
nand UO_2649 (O_2649,N_23625,N_20318);
and UO_2650 (O_2650,N_22821,N_21844);
nor UO_2651 (O_2651,N_20108,N_20264);
or UO_2652 (O_2652,N_21041,N_24285);
or UO_2653 (O_2653,N_23204,N_21894);
and UO_2654 (O_2654,N_20281,N_21842);
nor UO_2655 (O_2655,N_20712,N_24016);
nand UO_2656 (O_2656,N_23784,N_23515);
or UO_2657 (O_2657,N_23483,N_22462);
or UO_2658 (O_2658,N_24680,N_20457);
xor UO_2659 (O_2659,N_20465,N_21867);
xor UO_2660 (O_2660,N_24017,N_21346);
or UO_2661 (O_2661,N_22375,N_22268);
nor UO_2662 (O_2662,N_21768,N_23836);
nand UO_2663 (O_2663,N_20419,N_22563);
or UO_2664 (O_2664,N_20521,N_23920);
nand UO_2665 (O_2665,N_21099,N_22400);
or UO_2666 (O_2666,N_23800,N_21896);
or UO_2667 (O_2667,N_21076,N_20167);
nand UO_2668 (O_2668,N_24673,N_22157);
nor UO_2669 (O_2669,N_20951,N_22815);
xor UO_2670 (O_2670,N_23132,N_24543);
nor UO_2671 (O_2671,N_21682,N_22168);
xnor UO_2672 (O_2672,N_22238,N_21152);
and UO_2673 (O_2673,N_22630,N_22078);
nand UO_2674 (O_2674,N_23683,N_23180);
nand UO_2675 (O_2675,N_23799,N_23278);
nand UO_2676 (O_2676,N_21888,N_21279);
xnor UO_2677 (O_2677,N_24794,N_22058);
and UO_2678 (O_2678,N_21792,N_22082);
or UO_2679 (O_2679,N_24244,N_24530);
and UO_2680 (O_2680,N_22566,N_22833);
nand UO_2681 (O_2681,N_21377,N_23475);
xnor UO_2682 (O_2682,N_23657,N_22717);
xnor UO_2683 (O_2683,N_21008,N_21913);
or UO_2684 (O_2684,N_21133,N_21927);
or UO_2685 (O_2685,N_22419,N_22337);
xnor UO_2686 (O_2686,N_23165,N_23851);
nor UO_2687 (O_2687,N_20345,N_23074);
nand UO_2688 (O_2688,N_23449,N_20909);
nor UO_2689 (O_2689,N_20278,N_23604);
xor UO_2690 (O_2690,N_22764,N_23739);
and UO_2691 (O_2691,N_22808,N_21470);
nor UO_2692 (O_2692,N_20141,N_21940);
or UO_2693 (O_2693,N_20768,N_23882);
and UO_2694 (O_2694,N_24966,N_24613);
xnor UO_2695 (O_2695,N_20442,N_21459);
nor UO_2696 (O_2696,N_21141,N_23569);
nand UO_2697 (O_2697,N_23040,N_20942);
and UO_2698 (O_2698,N_24136,N_21036);
nand UO_2699 (O_2699,N_20646,N_23944);
and UO_2700 (O_2700,N_20245,N_24890);
nor UO_2701 (O_2701,N_20029,N_20788);
xnor UO_2702 (O_2702,N_22834,N_23107);
or UO_2703 (O_2703,N_21840,N_20330);
nand UO_2704 (O_2704,N_21817,N_24189);
nor UO_2705 (O_2705,N_24738,N_24453);
xor UO_2706 (O_2706,N_23396,N_21052);
nand UO_2707 (O_2707,N_23963,N_20913);
or UO_2708 (O_2708,N_24580,N_22764);
or UO_2709 (O_2709,N_24350,N_21611);
xor UO_2710 (O_2710,N_22687,N_23824);
nor UO_2711 (O_2711,N_21883,N_21431);
nand UO_2712 (O_2712,N_22950,N_20853);
and UO_2713 (O_2713,N_23142,N_23229);
or UO_2714 (O_2714,N_21632,N_21020);
nand UO_2715 (O_2715,N_24916,N_21650);
nor UO_2716 (O_2716,N_23102,N_24827);
nor UO_2717 (O_2717,N_20545,N_20121);
and UO_2718 (O_2718,N_22180,N_22426);
nand UO_2719 (O_2719,N_24090,N_23437);
or UO_2720 (O_2720,N_21062,N_23129);
and UO_2721 (O_2721,N_24041,N_22310);
xnor UO_2722 (O_2722,N_23947,N_21867);
xnor UO_2723 (O_2723,N_20457,N_20899);
and UO_2724 (O_2724,N_24105,N_24539);
or UO_2725 (O_2725,N_22852,N_22753);
and UO_2726 (O_2726,N_22051,N_20757);
or UO_2727 (O_2727,N_20864,N_22070);
nand UO_2728 (O_2728,N_20232,N_22909);
nor UO_2729 (O_2729,N_21337,N_21043);
nand UO_2730 (O_2730,N_24635,N_23707);
nand UO_2731 (O_2731,N_22101,N_24876);
and UO_2732 (O_2732,N_23427,N_24762);
xor UO_2733 (O_2733,N_20468,N_23119);
xor UO_2734 (O_2734,N_23291,N_24792);
nor UO_2735 (O_2735,N_24836,N_22496);
xor UO_2736 (O_2736,N_24435,N_24717);
or UO_2737 (O_2737,N_24498,N_20047);
nand UO_2738 (O_2738,N_24278,N_22121);
and UO_2739 (O_2739,N_22422,N_21988);
nand UO_2740 (O_2740,N_21944,N_23088);
nor UO_2741 (O_2741,N_23467,N_24145);
nand UO_2742 (O_2742,N_24030,N_23001);
and UO_2743 (O_2743,N_20040,N_21609);
nor UO_2744 (O_2744,N_20262,N_24965);
nand UO_2745 (O_2745,N_22160,N_23950);
nand UO_2746 (O_2746,N_23468,N_21809);
nor UO_2747 (O_2747,N_24075,N_23051);
nor UO_2748 (O_2748,N_24701,N_21320);
nor UO_2749 (O_2749,N_20457,N_23062);
nor UO_2750 (O_2750,N_22630,N_21308);
and UO_2751 (O_2751,N_24672,N_20346);
or UO_2752 (O_2752,N_24292,N_22179);
nand UO_2753 (O_2753,N_24711,N_23404);
xnor UO_2754 (O_2754,N_20284,N_20052);
nor UO_2755 (O_2755,N_23538,N_21961);
nor UO_2756 (O_2756,N_22791,N_22913);
nand UO_2757 (O_2757,N_21815,N_21478);
xnor UO_2758 (O_2758,N_21644,N_24982);
nand UO_2759 (O_2759,N_20710,N_21574);
or UO_2760 (O_2760,N_21735,N_20891);
xor UO_2761 (O_2761,N_22416,N_24632);
xnor UO_2762 (O_2762,N_20628,N_24490);
nor UO_2763 (O_2763,N_21574,N_20278);
xor UO_2764 (O_2764,N_23070,N_23059);
xnor UO_2765 (O_2765,N_20132,N_22927);
or UO_2766 (O_2766,N_21173,N_20136);
nor UO_2767 (O_2767,N_22062,N_20994);
nor UO_2768 (O_2768,N_21727,N_21376);
and UO_2769 (O_2769,N_20917,N_22035);
or UO_2770 (O_2770,N_22176,N_20925);
nor UO_2771 (O_2771,N_23113,N_20431);
and UO_2772 (O_2772,N_24175,N_22893);
nand UO_2773 (O_2773,N_21658,N_20752);
xor UO_2774 (O_2774,N_20895,N_20077);
nor UO_2775 (O_2775,N_24427,N_20205);
xnor UO_2776 (O_2776,N_23488,N_22265);
or UO_2777 (O_2777,N_22857,N_22019);
and UO_2778 (O_2778,N_22364,N_24446);
or UO_2779 (O_2779,N_20308,N_22485);
or UO_2780 (O_2780,N_20633,N_21199);
or UO_2781 (O_2781,N_21804,N_21501);
nor UO_2782 (O_2782,N_22315,N_21221);
nand UO_2783 (O_2783,N_22399,N_21674);
and UO_2784 (O_2784,N_21656,N_21903);
or UO_2785 (O_2785,N_20015,N_20104);
xor UO_2786 (O_2786,N_23230,N_23369);
xnor UO_2787 (O_2787,N_21146,N_21543);
or UO_2788 (O_2788,N_22535,N_20308);
nand UO_2789 (O_2789,N_24223,N_20291);
or UO_2790 (O_2790,N_23159,N_20235);
or UO_2791 (O_2791,N_22242,N_20641);
or UO_2792 (O_2792,N_22201,N_21654);
nor UO_2793 (O_2793,N_23368,N_21109);
nand UO_2794 (O_2794,N_20465,N_20352);
nand UO_2795 (O_2795,N_24066,N_21924);
xnor UO_2796 (O_2796,N_23413,N_23656);
nor UO_2797 (O_2797,N_24583,N_23036);
nor UO_2798 (O_2798,N_21146,N_21953);
and UO_2799 (O_2799,N_22698,N_21867);
xnor UO_2800 (O_2800,N_23451,N_24162);
nor UO_2801 (O_2801,N_20381,N_20364);
nor UO_2802 (O_2802,N_20557,N_22687);
xor UO_2803 (O_2803,N_24173,N_22842);
xnor UO_2804 (O_2804,N_21500,N_23207);
or UO_2805 (O_2805,N_20196,N_22300);
nand UO_2806 (O_2806,N_21442,N_24170);
or UO_2807 (O_2807,N_21712,N_22090);
and UO_2808 (O_2808,N_24611,N_23197);
nor UO_2809 (O_2809,N_24178,N_23284);
or UO_2810 (O_2810,N_22969,N_22375);
xnor UO_2811 (O_2811,N_20514,N_23828);
nor UO_2812 (O_2812,N_22900,N_22673);
xnor UO_2813 (O_2813,N_22335,N_21333);
and UO_2814 (O_2814,N_22164,N_20174);
nor UO_2815 (O_2815,N_20674,N_22829);
or UO_2816 (O_2816,N_23128,N_20560);
and UO_2817 (O_2817,N_24612,N_22502);
nor UO_2818 (O_2818,N_22296,N_20935);
nor UO_2819 (O_2819,N_21531,N_20561);
nand UO_2820 (O_2820,N_20893,N_21351);
xor UO_2821 (O_2821,N_21619,N_22636);
nor UO_2822 (O_2822,N_22717,N_20408);
nor UO_2823 (O_2823,N_22482,N_21979);
xor UO_2824 (O_2824,N_21950,N_20525);
xor UO_2825 (O_2825,N_23162,N_20815);
and UO_2826 (O_2826,N_20651,N_21237);
xor UO_2827 (O_2827,N_20227,N_24443);
xor UO_2828 (O_2828,N_22054,N_23845);
nand UO_2829 (O_2829,N_24124,N_20102);
and UO_2830 (O_2830,N_22892,N_20556);
nor UO_2831 (O_2831,N_20847,N_22058);
or UO_2832 (O_2832,N_24443,N_20417);
xor UO_2833 (O_2833,N_24399,N_23003);
or UO_2834 (O_2834,N_22050,N_21526);
and UO_2835 (O_2835,N_24600,N_20186);
or UO_2836 (O_2836,N_22508,N_20762);
and UO_2837 (O_2837,N_24234,N_21224);
nand UO_2838 (O_2838,N_21424,N_22780);
nand UO_2839 (O_2839,N_21727,N_22038);
and UO_2840 (O_2840,N_24822,N_23273);
nand UO_2841 (O_2841,N_24070,N_23234);
and UO_2842 (O_2842,N_22011,N_22905);
and UO_2843 (O_2843,N_21147,N_21478);
and UO_2844 (O_2844,N_23674,N_23699);
xnor UO_2845 (O_2845,N_24865,N_23427);
and UO_2846 (O_2846,N_21002,N_23553);
or UO_2847 (O_2847,N_24383,N_24586);
xor UO_2848 (O_2848,N_23413,N_23906);
nor UO_2849 (O_2849,N_22019,N_23795);
and UO_2850 (O_2850,N_24342,N_21482);
and UO_2851 (O_2851,N_23612,N_21119);
xnor UO_2852 (O_2852,N_22032,N_22931);
xnor UO_2853 (O_2853,N_22785,N_22005);
or UO_2854 (O_2854,N_21035,N_22080);
or UO_2855 (O_2855,N_21564,N_20799);
nand UO_2856 (O_2856,N_21159,N_22683);
nand UO_2857 (O_2857,N_22693,N_21948);
or UO_2858 (O_2858,N_24729,N_22006);
xor UO_2859 (O_2859,N_23831,N_22468);
nand UO_2860 (O_2860,N_21630,N_20193);
or UO_2861 (O_2861,N_20807,N_21522);
nor UO_2862 (O_2862,N_21612,N_21866);
and UO_2863 (O_2863,N_23417,N_21289);
nand UO_2864 (O_2864,N_23763,N_20365);
and UO_2865 (O_2865,N_20272,N_22114);
xor UO_2866 (O_2866,N_24729,N_20507);
or UO_2867 (O_2867,N_22897,N_24126);
nand UO_2868 (O_2868,N_22802,N_24845);
nor UO_2869 (O_2869,N_22679,N_21249);
or UO_2870 (O_2870,N_24080,N_24670);
or UO_2871 (O_2871,N_24205,N_23948);
nor UO_2872 (O_2872,N_24146,N_23947);
nand UO_2873 (O_2873,N_20873,N_23079);
xnor UO_2874 (O_2874,N_24249,N_20029);
or UO_2875 (O_2875,N_20256,N_22865);
nor UO_2876 (O_2876,N_20289,N_20830);
nor UO_2877 (O_2877,N_23983,N_22251);
nor UO_2878 (O_2878,N_24945,N_20011);
nor UO_2879 (O_2879,N_24368,N_21751);
nand UO_2880 (O_2880,N_24085,N_22576);
nand UO_2881 (O_2881,N_23566,N_22214);
or UO_2882 (O_2882,N_21227,N_20038);
or UO_2883 (O_2883,N_20137,N_24243);
xor UO_2884 (O_2884,N_24963,N_20192);
nand UO_2885 (O_2885,N_20273,N_23541);
nand UO_2886 (O_2886,N_24536,N_22093);
nor UO_2887 (O_2887,N_24087,N_24415);
nand UO_2888 (O_2888,N_22955,N_20980);
or UO_2889 (O_2889,N_21746,N_24652);
and UO_2890 (O_2890,N_20286,N_21503);
nand UO_2891 (O_2891,N_22135,N_24070);
xor UO_2892 (O_2892,N_24128,N_22285);
nor UO_2893 (O_2893,N_24558,N_21146);
nand UO_2894 (O_2894,N_23568,N_20184);
and UO_2895 (O_2895,N_22812,N_21138);
or UO_2896 (O_2896,N_21306,N_20059);
xnor UO_2897 (O_2897,N_21795,N_23540);
or UO_2898 (O_2898,N_20981,N_24550);
nand UO_2899 (O_2899,N_22967,N_20914);
and UO_2900 (O_2900,N_21960,N_24018);
xor UO_2901 (O_2901,N_20305,N_22766);
nor UO_2902 (O_2902,N_23562,N_20510);
xnor UO_2903 (O_2903,N_21683,N_20926);
nor UO_2904 (O_2904,N_20620,N_20348);
or UO_2905 (O_2905,N_20693,N_22585);
nor UO_2906 (O_2906,N_21748,N_24421);
nor UO_2907 (O_2907,N_21654,N_23148);
xor UO_2908 (O_2908,N_22530,N_22631);
xnor UO_2909 (O_2909,N_24585,N_22119);
xor UO_2910 (O_2910,N_23601,N_20157);
or UO_2911 (O_2911,N_23607,N_22590);
nand UO_2912 (O_2912,N_22727,N_20378);
nor UO_2913 (O_2913,N_21139,N_22865);
and UO_2914 (O_2914,N_21227,N_21462);
nand UO_2915 (O_2915,N_24359,N_23422);
nand UO_2916 (O_2916,N_24289,N_23918);
or UO_2917 (O_2917,N_22403,N_24324);
xnor UO_2918 (O_2918,N_23469,N_23192);
or UO_2919 (O_2919,N_24077,N_20589);
xnor UO_2920 (O_2920,N_20705,N_23737);
or UO_2921 (O_2921,N_23510,N_22315);
or UO_2922 (O_2922,N_21888,N_20661);
nor UO_2923 (O_2923,N_22113,N_24109);
xnor UO_2924 (O_2924,N_24466,N_23736);
xnor UO_2925 (O_2925,N_23220,N_22833);
nor UO_2926 (O_2926,N_23104,N_24075);
and UO_2927 (O_2927,N_24818,N_21590);
or UO_2928 (O_2928,N_24573,N_22938);
nand UO_2929 (O_2929,N_21487,N_23652);
nor UO_2930 (O_2930,N_21585,N_20951);
xor UO_2931 (O_2931,N_22069,N_24800);
nor UO_2932 (O_2932,N_22908,N_22370);
nand UO_2933 (O_2933,N_20447,N_20136);
nand UO_2934 (O_2934,N_22358,N_23165);
nor UO_2935 (O_2935,N_21237,N_24368);
xnor UO_2936 (O_2936,N_24261,N_24124);
or UO_2937 (O_2937,N_23295,N_21022);
nor UO_2938 (O_2938,N_20800,N_24628);
nor UO_2939 (O_2939,N_24212,N_23812);
nor UO_2940 (O_2940,N_21371,N_22939);
or UO_2941 (O_2941,N_23316,N_23646);
xor UO_2942 (O_2942,N_24191,N_24018);
or UO_2943 (O_2943,N_24849,N_24795);
nor UO_2944 (O_2944,N_22005,N_21687);
or UO_2945 (O_2945,N_22606,N_22977);
or UO_2946 (O_2946,N_23700,N_21548);
nor UO_2947 (O_2947,N_24263,N_21721);
xor UO_2948 (O_2948,N_21452,N_21784);
xnor UO_2949 (O_2949,N_23993,N_21800);
or UO_2950 (O_2950,N_23498,N_24722);
xnor UO_2951 (O_2951,N_24416,N_20002);
or UO_2952 (O_2952,N_22650,N_20607);
nand UO_2953 (O_2953,N_22603,N_23306);
nand UO_2954 (O_2954,N_24776,N_23775);
nand UO_2955 (O_2955,N_22807,N_23961);
xor UO_2956 (O_2956,N_22583,N_24743);
xnor UO_2957 (O_2957,N_20654,N_21210);
and UO_2958 (O_2958,N_24984,N_20696);
or UO_2959 (O_2959,N_21748,N_24092);
and UO_2960 (O_2960,N_23169,N_24156);
nor UO_2961 (O_2961,N_24091,N_22390);
xor UO_2962 (O_2962,N_20729,N_20212);
and UO_2963 (O_2963,N_23169,N_23961);
nor UO_2964 (O_2964,N_23611,N_24360);
or UO_2965 (O_2965,N_22848,N_23421);
and UO_2966 (O_2966,N_22104,N_21070);
xor UO_2967 (O_2967,N_22788,N_20459);
and UO_2968 (O_2968,N_23475,N_23393);
or UO_2969 (O_2969,N_23430,N_23728);
nor UO_2970 (O_2970,N_21182,N_21390);
xnor UO_2971 (O_2971,N_20535,N_24037);
nor UO_2972 (O_2972,N_21849,N_22932);
nand UO_2973 (O_2973,N_21583,N_24481);
nor UO_2974 (O_2974,N_23229,N_22099);
nor UO_2975 (O_2975,N_22949,N_23065);
nand UO_2976 (O_2976,N_24532,N_22018);
nand UO_2977 (O_2977,N_24518,N_22739);
nor UO_2978 (O_2978,N_21720,N_24113);
or UO_2979 (O_2979,N_21333,N_22541);
nand UO_2980 (O_2980,N_24395,N_21217);
and UO_2981 (O_2981,N_23090,N_24498);
xor UO_2982 (O_2982,N_23510,N_21728);
xnor UO_2983 (O_2983,N_20196,N_24878);
xnor UO_2984 (O_2984,N_24588,N_24669);
and UO_2985 (O_2985,N_22919,N_22466);
nand UO_2986 (O_2986,N_22601,N_22387);
nand UO_2987 (O_2987,N_22402,N_23864);
or UO_2988 (O_2988,N_21737,N_22591);
or UO_2989 (O_2989,N_24180,N_23756);
and UO_2990 (O_2990,N_20260,N_24625);
and UO_2991 (O_2991,N_22424,N_21817);
and UO_2992 (O_2992,N_23689,N_23786);
nor UO_2993 (O_2993,N_23212,N_23385);
nand UO_2994 (O_2994,N_22462,N_20682);
and UO_2995 (O_2995,N_20321,N_22998);
nand UO_2996 (O_2996,N_20669,N_21765);
nand UO_2997 (O_2997,N_20313,N_20246);
and UO_2998 (O_2998,N_20846,N_22926);
or UO_2999 (O_2999,N_22746,N_21834);
endmodule