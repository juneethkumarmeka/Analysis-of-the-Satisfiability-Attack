module basic_500_3000_500_50_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_72,In_453);
or U1 (N_1,In_442,In_329);
nand U2 (N_2,In_263,In_154);
nand U3 (N_3,In_308,In_368);
nor U4 (N_4,In_87,In_491);
nand U5 (N_5,In_279,In_365);
xor U6 (N_6,In_255,In_425);
xnor U7 (N_7,In_139,In_466);
nand U8 (N_8,In_307,In_15);
nand U9 (N_9,In_496,In_495);
or U10 (N_10,In_124,In_483);
nand U11 (N_11,In_82,In_347);
xor U12 (N_12,In_437,In_353);
or U13 (N_13,In_311,In_249);
or U14 (N_14,In_235,In_81);
nand U15 (N_15,In_53,In_444);
nor U16 (N_16,In_273,In_141);
xor U17 (N_17,In_216,In_56);
and U18 (N_18,In_169,In_332);
or U19 (N_19,In_184,In_327);
nand U20 (N_20,In_193,In_383);
or U21 (N_21,In_423,In_277);
nand U22 (N_22,In_232,In_73);
xnor U23 (N_23,In_213,In_486);
nor U24 (N_24,In_3,In_92);
and U25 (N_25,In_234,In_497);
or U26 (N_26,In_11,In_5);
xor U27 (N_27,In_421,In_320);
xnor U28 (N_28,In_465,In_138);
nand U29 (N_29,In_168,In_121);
xor U30 (N_30,In_108,In_0);
and U31 (N_31,In_284,In_116);
nor U32 (N_32,In_50,In_155);
or U33 (N_33,In_104,In_162);
xor U34 (N_34,In_387,In_258);
and U35 (N_35,In_191,In_370);
nor U36 (N_36,In_412,In_343);
xnor U37 (N_37,In_474,In_44);
or U38 (N_38,In_23,In_315);
nand U39 (N_39,In_71,In_183);
nor U40 (N_40,In_489,In_254);
xnor U41 (N_41,In_237,In_51);
xor U42 (N_42,In_174,In_276);
nor U43 (N_43,In_460,In_159);
xor U44 (N_44,In_221,In_268);
and U45 (N_45,In_170,In_84);
nor U46 (N_46,In_404,In_328);
xnor U47 (N_47,In_222,In_274);
xor U48 (N_48,In_59,In_76);
nand U49 (N_49,In_269,In_122);
or U50 (N_50,In_402,In_107);
nand U51 (N_51,In_61,In_231);
xor U52 (N_52,In_24,In_285);
nand U53 (N_53,In_78,In_94);
or U54 (N_54,In_450,In_325);
or U55 (N_55,In_447,In_27);
nand U56 (N_56,In_409,In_481);
and U57 (N_57,In_334,In_54);
or U58 (N_58,In_103,In_242);
nand U59 (N_59,In_98,In_380);
nand U60 (N_60,In_93,In_131);
or U61 (N_61,In_397,N_31);
nor U62 (N_62,In_123,In_405);
nand U63 (N_63,In_386,In_462);
nand U64 (N_64,In_22,N_23);
and U65 (N_65,In_185,In_323);
and U66 (N_66,In_128,In_469);
or U67 (N_67,In_270,In_135);
nor U68 (N_68,In_105,N_55);
xor U69 (N_69,In_314,In_398);
xor U70 (N_70,In_58,In_459);
xnor U71 (N_71,In_291,In_424);
or U72 (N_72,In_228,In_297);
and U73 (N_73,In_223,In_403);
and U74 (N_74,In_245,In_261);
nand U75 (N_75,In_326,In_449);
or U76 (N_76,In_161,N_39);
and U77 (N_77,N_14,In_182);
or U78 (N_78,In_375,In_195);
nor U79 (N_79,In_211,In_472);
nor U80 (N_80,In_256,In_2);
xnor U81 (N_81,In_417,In_363);
and U82 (N_82,In_248,N_32);
xnor U83 (N_83,N_42,In_374);
nor U84 (N_84,In_118,In_149);
xnor U85 (N_85,N_41,In_25);
xnor U86 (N_86,In_257,N_17);
and U87 (N_87,In_392,In_341);
and U88 (N_88,In_172,In_319);
and U89 (N_89,N_11,In_280);
nor U90 (N_90,In_8,In_371);
nor U91 (N_91,In_321,In_342);
and U92 (N_92,In_492,In_42);
nand U93 (N_93,In_90,In_125);
and U94 (N_94,In_391,In_385);
nor U95 (N_95,In_160,In_439);
and U96 (N_96,N_47,In_306);
nand U97 (N_97,In_494,In_146);
or U98 (N_98,N_12,In_362);
or U99 (N_99,In_384,In_83);
nor U100 (N_100,In_215,In_113);
and U101 (N_101,In_441,In_173);
xor U102 (N_102,In_477,In_432);
xor U103 (N_103,In_150,N_16);
xnor U104 (N_104,In_251,In_37);
nor U105 (N_105,In_230,In_85);
or U106 (N_106,In_318,N_19);
or U107 (N_107,N_36,N_37);
nor U108 (N_108,In_74,In_243);
nand U109 (N_109,In_357,N_20);
nor U110 (N_110,N_38,In_281);
and U111 (N_111,In_14,In_229);
nor U112 (N_112,In_140,In_18);
nand U113 (N_113,In_132,In_322);
or U114 (N_114,In_1,In_266);
nor U115 (N_115,In_80,In_227);
xnor U116 (N_116,In_298,In_356);
or U117 (N_117,In_448,In_331);
and U118 (N_118,In_264,N_27);
xor U119 (N_119,In_130,N_51);
nor U120 (N_120,In_272,In_36);
or U121 (N_121,In_79,In_147);
nand U122 (N_122,In_426,In_354);
or U123 (N_123,In_236,In_247);
nand U124 (N_124,In_389,In_422);
nand U125 (N_125,In_286,N_8);
or U126 (N_126,In_420,In_260);
nand U127 (N_127,In_88,In_373);
or U128 (N_128,N_100,In_351);
or U129 (N_129,In_144,In_180);
nand U130 (N_130,In_46,N_2);
nor U131 (N_131,In_259,In_464);
or U132 (N_132,N_113,In_438);
or U133 (N_133,In_119,N_4);
nor U134 (N_134,N_109,In_241);
xor U135 (N_135,In_200,In_152);
xor U136 (N_136,In_451,In_299);
nand U137 (N_137,In_153,In_359);
and U138 (N_138,N_48,In_394);
nor U139 (N_139,N_3,N_34);
nand U140 (N_140,N_43,In_488);
xnor U141 (N_141,In_456,In_339);
nor U142 (N_142,In_64,In_69);
xor U143 (N_143,In_369,In_115);
and U144 (N_144,N_6,In_324);
nor U145 (N_145,N_116,N_102);
and U146 (N_146,In_114,In_35);
nand U147 (N_147,In_9,N_26);
xor U148 (N_148,In_10,In_177);
nor U149 (N_149,In_151,In_95);
nand U150 (N_150,In_209,In_210);
xnor U151 (N_151,In_109,In_303);
nor U152 (N_152,In_480,In_262);
xor U153 (N_153,In_396,N_62);
and U154 (N_154,In_330,In_436);
nand U155 (N_155,In_454,N_108);
xor U156 (N_156,N_35,In_360);
nor U157 (N_157,In_337,In_302);
nand U158 (N_158,In_290,In_293);
nor U159 (N_159,In_187,In_77);
and U160 (N_160,In_400,In_47);
nand U161 (N_161,In_296,In_431);
nand U162 (N_162,In_156,In_295);
xnor U163 (N_163,In_34,In_41);
xnor U164 (N_164,In_30,In_443);
and U165 (N_165,In_127,In_294);
or U166 (N_166,In_67,N_65);
xnor U167 (N_167,In_493,N_117);
nor U168 (N_168,In_350,N_13);
nand U169 (N_169,In_129,In_445);
and U170 (N_170,In_393,N_106);
or U171 (N_171,In_345,N_1);
xnor U172 (N_172,In_317,N_71);
xor U173 (N_173,In_240,In_112);
and U174 (N_174,In_188,In_461);
and U175 (N_175,In_457,In_134);
and U176 (N_176,N_79,N_90);
nand U177 (N_177,In_239,In_26);
xor U178 (N_178,In_120,N_87);
nor U179 (N_179,In_189,N_98);
xor U180 (N_180,N_9,N_174);
nor U181 (N_181,In_309,In_143);
or U182 (N_182,In_287,In_68);
nor U183 (N_183,N_58,N_129);
or U184 (N_184,In_48,N_85);
and U185 (N_185,In_142,In_205);
or U186 (N_186,In_300,In_406);
or U187 (N_187,In_304,In_246);
nand U188 (N_188,In_60,N_22);
nor U189 (N_189,In_194,In_275);
xor U190 (N_190,In_207,In_99);
nor U191 (N_191,In_446,In_479);
and U192 (N_192,In_111,In_201);
and U193 (N_193,N_89,In_6);
nor U194 (N_194,N_5,N_103);
or U195 (N_195,N_165,In_43);
and U196 (N_196,In_490,In_401);
nand U197 (N_197,In_358,In_196);
nand U198 (N_198,N_30,In_28);
nand U199 (N_199,In_250,N_119);
nand U200 (N_200,N_125,In_407);
nand U201 (N_201,N_91,In_433);
xnor U202 (N_202,N_145,In_219);
nor U203 (N_203,In_166,N_104);
nor U204 (N_204,In_366,In_411);
xnor U205 (N_205,N_82,In_413);
or U206 (N_206,N_175,N_50);
nand U207 (N_207,In_190,N_136);
nand U208 (N_208,In_267,In_333);
xor U209 (N_209,In_499,In_55);
and U210 (N_210,N_146,In_430);
or U211 (N_211,In_137,In_70);
and U212 (N_212,In_212,In_225);
nor U213 (N_213,In_468,In_157);
or U214 (N_214,N_69,In_89);
or U215 (N_215,In_305,In_416);
nor U216 (N_216,In_313,In_399);
and U217 (N_217,N_101,N_149);
nand U218 (N_218,N_44,In_158);
and U219 (N_219,In_289,N_124);
xnor U220 (N_220,In_301,N_63);
or U221 (N_221,In_288,In_19);
and U222 (N_222,N_141,In_388);
xnor U223 (N_223,N_95,N_83);
xor U224 (N_224,N_176,In_163);
nand U225 (N_225,In_473,In_164);
or U226 (N_226,In_471,N_142);
and U227 (N_227,In_45,In_16);
and U228 (N_228,In_38,In_126);
or U229 (N_229,N_156,In_271);
and U230 (N_230,N_172,N_92);
and U231 (N_231,In_265,N_123);
or U232 (N_232,N_52,In_348);
or U233 (N_233,N_178,N_53);
nand U234 (N_234,N_153,In_336);
or U235 (N_235,In_349,N_107);
and U236 (N_236,In_382,In_4);
nor U237 (N_237,In_206,N_167);
nor U238 (N_238,In_428,In_352);
xnor U239 (N_239,In_204,N_60);
nand U240 (N_240,N_207,N_203);
and U241 (N_241,N_64,N_206);
and U242 (N_242,N_81,N_194);
nor U243 (N_243,In_203,N_202);
nand U244 (N_244,N_205,N_171);
nor U245 (N_245,In_179,N_111);
nor U246 (N_246,N_179,N_216);
xor U247 (N_247,N_127,N_147);
nand U248 (N_248,In_376,N_0);
xor U249 (N_249,N_130,N_164);
xor U250 (N_250,In_198,In_427);
nand U251 (N_251,N_120,N_219);
or U252 (N_252,In_452,In_485);
or U253 (N_253,N_121,N_7);
and U254 (N_254,In_136,N_234);
or U255 (N_255,N_223,N_239);
xnor U256 (N_256,In_419,N_134);
and U257 (N_257,In_176,In_335);
or U258 (N_258,In_252,In_57);
or U259 (N_259,N_230,N_139);
or U260 (N_260,N_187,In_364);
nand U261 (N_261,In_310,N_162);
and U262 (N_262,N_168,N_18);
nand U263 (N_263,In_475,In_467);
nor U264 (N_264,N_118,N_232);
and U265 (N_265,In_102,N_192);
and U266 (N_266,N_40,N_169);
nor U267 (N_267,In_312,N_222);
nor U268 (N_268,In_7,N_152);
nor U269 (N_269,N_137,In_482);
xnor U270 (N_270,N_233,N_229);
nor U271 (N_271,In_414,In_29);
nor U272 (N_272,N_200,In_282);
or U273 (N_273,In_226,N_224);
and U274 (N_274,In_244,N_211);
or U275 (N_275,N_84,In_145);
nor U276 (N_276,In_253,N_46);
nand U277 (N_277,In_415,In_197);
xnor U278 (N_278,In_101,In_435);
nor U279 (N_279,In_429,In_316);
and U280 (N_280,N_218,In_49);
xnor U281 (N_281,In_233,In_278);
nor U282 (N_282,N_143,In_478);
nor U283 (N_283,In_208,In_181);
nor U284 (N_284,In_338,N_10);
or U285 (N_285,N_54,N_140);
nor U286 (N_286,N_73,N_221);
or U287 (N_287,In_378,N_197);
and U288 (N_288,N_99,In_66);
xor U289 (N_289,In_476,In_40);
nor U290 (N_290,N_28,N_128);
nor U291 (N_291,N_184,In_220);
and U292 (N_292,In_458,In_148);
nand U293 (N_293,In_418,In_75);
or U294 (N_294,N_56,In_202);
nand U295 (N_295,In_165,N_220);
xor U296 (N_296,N_191,In_379);
nand U297 (N_297,N_110,N_231);
and U298 (N_298,In_100,N_235);
or U299 (N_299,N_195,N_144);
and U300 (N_300,In_17,N_77);
nand U301 (N_301,In_346,In_13);
or U302 (N_302,N_183,In_367);
nor U303 (N_303,N_273,N_198);
nor U304 (N_304,N_228,N_157);
nor U305 (N_305,N_59,N_68);
nand U306 (N_306,N_122,N_265);
or U307 (N_307,N_131,N_188);
nor U308 (N_308,N_281,N_236);
or U309 (N_309,N_282,In_214);
and U310 (N_310,N_253,N_155);
or U311 (N_311,N_185,In_86);
nand U312 (N_312,In_340,N_249);
nand U313 (N_313,N_268,N_214);
or U314 (N_314,N_240,N_180);
or U315 (N_315,In_12,N_264);
nand U316 (N_316,N_250,N_193);
nand U317 (N_317,N_263,N_213);
or U318 (N_318,N_29,In_463);
and U319 (N_319,N_74,N_33);
nor U320 (N_320,In_487,In_20);
or U321 (N_321,N_93,In_52);
or U322 (N_322,In_484,N_288);
and U323 (N_323,In_32,N_259);
or U324 (N_324,N_159,N_258);
xnor U325 (N_325,N_208,In_395);
nand U326 (N_326,N_247,N_244);
nand U327 (N_327,N_278,In_238);
and U328 (N_328,N_21,In_344);
or U329 (N_329,N_266,N_210);
nor U330 (N_330,In_434,N_291);
nor U331 (N_331,N_126,N_170);
or U332 (N_332,In_224,N_61);
and U333 (N_333,In_377,In_175);
and U334 (N_334,N_25,N_163);
nand U335 (N_335,N_270,N_275);
or U336 (N_336,In_62,N_57);
nor U337 (N_337,In_217,N_212);
or U338 (N_338,In_63,In_283);
xor U339 (N_339,N_114,N_279);
or U340 (N_340,In_390,N_72);
and U341 (N_341,N_67,N_112);
xnor U342 (N_342,N_15,N_225);
or U343 (N_343,N_257,In_381);
and U344 (N_344,N_227,N_161);
and U345 (N_345,N_286,N_260);
and U346 (N_346,N_173,N_243);
nand U347 (N_347,N_105,In_106);
nor U348 (N_348,N_76,N_287);
and U349 (N_349,In_110,N_135);
and U350 (N_350,In_97,In_292);
and U351 (N_351,N_276,N_75);
or U352 (N_352,N_271,N_277);
and U353 (N_353,N_166,N_283);
or U354 (N_354,In_218,N_133);
xnor U355 (N_355,N_66,In_171);
and U356 (N_356,N_255,In_91);
xnor U357 (N_357,N_251,In_372);
or U358 (N_358,N_189,N_154);
nor U359 (N_359,N_262,In_440);
xnor U360 (N_360,N_318,N_305);
nor U361 (N_361,N_350,N_274);
xnor U362 (N_362,N_352,N_284);
nand U363 (N_363,In_410,N_310);
xor U364 (N_364,N_302,N_340);
or U365 (N_365,N_86,N_343);
or U366 (N_366,In_21,N_80);
or U367 (N_367,N_325,N_94);
and U368 (N_368,N_349,N_267);
nand U369 (N_369,In_470,N_215);
or U370 (N_370,N_217,N_345);
nand U371 (N_371,N_150,N_196);
nand U372 (N_372,N_158,N_272);
or U373 (N_373,N_115,N_181);
xnor U374 (N_374,N_182,N_313);
or U375 (N_375,N_256,N_320);
xor U376 (N_376,In_39,N_280);
nor U377 (N_377,N_242,N_307);
nand U378 (N_378,N_151,N_88);
nor U379 (N_379,N_331,N_45);
nand U380 (N_380,N_312,N_348);
or U381 (N_381,N_328,N_321);
or U382 (N_382,N_356,N_358);
or U383 (N_383,In_199,N_248);
nand U384 (N_384,In_133,N_355);
nor U385 (N_385,N_327,N_357);
nor U386 (N_386,N_252,N_317);
nor U387 (N_387,N_298,N_308);
xnor U388 (N_388,N_346,N_344);
or U389 (N_389,N_226,N_245);
and U390 (N_390,N_160,N_347);
and U391 (N_391,N_148,In_167);
and U392 (N_392,In_33,N_292);
xor U393 (N_393,In_96,N_296);
xnor U394 (N_394,N_314,N_201);
xnor U395 (N_395,N_285,N_315);
nand U396 (N_396,N_329,N_186);
nor U397 (N_397,In_178,N_290);
nand U398 (N_398,N_269,N_204);
xnor U399 (N_399,N_330,N_334);
nor U400 (N_400,N_303,In_455);
or U401 (N_401,N_319,N_138);
nor U402 (N_402,N_351,N_261);
xnor U403 (N_403,N_78,N_254);
nand U404 (N_404,N_354,In_355);
or U405 (N_405,N_24,N_316);
and U406 (N_406,N_336,In_361);
xnor U407 (N_407,N_294,N_237);
nor U408 (N_408,N_338,N_339);
xor U409 (N_409,N_324,N_342);
xnor U410 (N_410,N_289,N_70);
xor U411 (N_411,N_306,N_96);
nand U412 (N_412,N_322,N_209);
nor U413 (N_413,N_49,N_337);
nand U414 (N_414,N_359,In_65);
nor U415 (N_415,N_190,N_333);
xor U416 (N_416,N_177,N_311);
and U417 (N_417,N_335,In_117);
and U418 (N_418,N_309,N_300);
nor U419 (N_419,N_341,N_199);
nor U420 (N_420,In_31,N_379);
nand U421 (N_421,N_361,N_382);
xnor U422 (N_422,N_295,N_392);
nand U423 (N_423,N_380,N_370);
nand U424 (N_424,N_394,N_299);
xnor U425 (N_425,N_387,In_498);
or U426 (N_426,N_407,N_398);
nor U427 (N_427,N_301,N_384);
nand U428 (N_428,N_366,N_323);
or U429 (N_429,N_293,N_389);
nor U430 (N_430,N_406,N_381);
or U431 (N_431,N_395,N_332);
and U432 (N_432,N_403,N_365);
xnor U433 (N_433,N_416,N_238);
and U434 (N_434,N_418,N_399);
and U435 (N_435,In_186,N_368);
nand U436 (N_436,N_376,N_363);
or U437 (N_437,N_362,N_404);
nand U438 (N_438,N_419,N_326);
or U439 (N_439,N_408,N_375);
nor U440 (N_440,N_297,N_383);
nor U441 (N_441,N_378,N_246);
nand U442 (N_442,N_97,N_377);
nor U443 (N_443,N_413,N_415);
or U444 (N_444,N_304,N_353);
nand U445 (N_445,N_396,In_408);
or U446 (N_446,N_371,N_412);
and U447 (N_447,N_132,N_417);
nand U448 (N_448,N_390,N_386);
or U449 (N_449,N_397,N_374);
and U450 (N_450,N_364,N_393);
and U451 (N_451,In_192,N_409);
nor U452 (N_452,N_401,N_405);
xnor U453 (N_453,N_411,N_367);
and U454 (N_454,N_410,N_360);
and U455 (N_455,N_391,N_400);
nand U456 (N_456,N_369,N_388);
or U457 (N_457,N_373,N_414);
or U458 (N_458,N_241,N_385);
nor U459 (N_459,N_372,N_402);
or U460 (N_460,N_408,N_403);
and U461 (N_461,N_375,N_419);
and U462 (N_462,N_390,N_301);
xnor U463 (N_463,N_301,N_401);
nand U464 (N_464,N_295,N_363);
and U465 (N_465,N_246,N_401);
and U466 (N_466,In_186,N_416);
xnor U467 (N_467,N_364,N_403);
nand U468 (N_468,N_385,N_364);
nand U469 (N_469,N_372,N_375);
xnor U470 (N_470,N_378,N_406);
xnor U471 (N_471,N_362,N_377);
xor U472 (N_472,N_360,N_398);
nor U473 (N_473,N_381,N_412);
nand U474 (N_474,N_391,N_370);
xnor U475 (N_475,N_374,N_332);
or U476 (N_476,N_241,N_401);
nor U477 (N_477,N_391,N_373);
nand U478 (N_478,N_360,N_361);
nand U479 (N_479,N_401,In_186);
xor U480 (N_480,N_442,N_443);
and U481 (N_481,N_460,N_421);
or U482 (N_482,N_436,N_438);
xnor U483 (N_483,N_464,N_479);
xor U484 (N_484,N_462,N_452);
nor U485 (N_485,N_475,N_447);
and U486 (N_486,N_432,N_444);
or U487 (N_487,N_477,N_430);
xor U488 (N_488,N_472,N_453);
or U489 (N_489,N_433,N_478);
xor U490 (N_490,N_471,N_476);
xor U491 (N_491,N_468,N_423);
nor U492 (N_492,N_450,N_454);
and U493 (N_493,N_420,N_463);
xnor U494 (N_494,N_455,N_466);
or U495 (N_495,N_473,N_422);
nand U496 (N_496,N_439,N_437);
or U497 (N_497,N_459,N_429);
and U498 (N_498,N_469,N_435);
nand U499 (N_499,N_474,N_428);
nand U500 (N_500,N_446,N_461);
and U501 (N_501,N_425,N_426);
or U502 (N_502,N_449,N_431);
nand U503 (N_503,N_424,N_467);
or U504 (N_504,N_448,N_465);
nor U505 (N_505,N_434,N_457);
and U506 (N_506,N_451,N_470);
nand U507 (N_507,N_445,N_441);
xor U508 (N_508,N_427,N_456);
or U509 (N_509,N_458,N_440);
and U510 (N_510,N_443,N_438);
and U511 (N_511,N_426,N_469);
or U512 (N_512,N_447,N_437);
nand U513 (N_513,N_449,N_441);
or U514 (N_514,N_423,N_458);
xnor U515 (N_515,N_425,N_451);
nand U516 (N_516,N_421,N_434);
or U517 (N_517,N_449,N_435);
xnor U518 (N_518,N_455,N_433);
or U519 (N_519,N_468,N_446);
xor U520 (N_520,N_451,N_455);
xor U521 (N_521,N_472,N_446);
or U522 (N_522,N_423,N_469);
nand U523 (N_523,N_471,N_464);
and U524 (N_524,N_476,N_454);
nor U525 (N_525,N_470,N_452);
and U526 (N_526,N_431,N_464);
xnor U527 (N_527,N_430,N_437);
nor U528 (N_528,N_473,N_478);
or U529 (N_529,N_420,N_476);
nor U530 (N_530,N_422,N_453);
nor U531 (N_531,N_459,N_464);
xor U532 (N_532,N_476,N_468);
and U533 (N_533,N_467,N_471);
xor U534 (N_534,N_461,N_422);
or U535 (N_535,N_436,N_442);
nand U536 (N_536,N_452,N_427);
nand U537 (N_537,N_445,N_423);
nor U538 (N_538,N_436,N_473);
xor U539 (N_539,N_470,N_427);
nor U540 (N_540,N_512,N_525);
nand U541 (N_541,N_481,N_507);
xnor U542 (N_542,N_485,N_532);
and U543 (N_543,N_503,N_516);
or U544 (N_544,N_498,N_502);
or U545 (N_545,N_505,N_486);
nor U546 (N_546,N_514,N_500);
nor U547 (N_547,N_494,N_526);
xnor U548 (N_548,N_488,N_497);
nand U549 (N_549,N_538,N_517);
and U550 (N_550,N_499,N_492);
xor U551 (N_551,N_521,N_511);
and U552 (N_552,N_491,N_487);
xor U553 (N_553,N_509,N_480);
or U554 (N_554,N_508,N_496);
nand U555 (N_555,N_537,N_483);
nor U556 (N_556,N_531,N_495);
and U557 (N_557,N_518,N_520);
nand U558 (N_558,N_489,N_493);
or U559 (N_559,N_510,N_529);
nand U560 (N_560,N_534,N_515);
xor U561 (N_561,N_484,N_535);
xnor U562 (N_562,N_490,N_519);
nor U563 (N_563,N_536,N_539);
nand U564 (N_564,N_504,N_482);
or U565 (N_565,N_528,N_501);
or U566 (N_566,N_513,N_533);
nand U567 (N_567,N_506,N_530);
nor U568 (N_568,N_527,N_522);
and U569 (N_569,N_523,N_524);
nand U570 (N_570,N_514,N_482);
and U571 (N_571,N_525,N_504);
nor U572 (N_572,N_532,N_514);
or U573 (N_573,N_538,N_515);
xnor U574 (N_574,N_518,N_525);
nand U575 (N_575,N_503,N_532);
nor U576 (N_576,N_497,N_518);
or U577 (N_577,N_492,N_513);
nand U578 (N_578,N_528,N_487);
nand U579 (N_579,N_528,N_524);
and U580 (N_580,N_516,N_482);
nand U581 (N_581,N_486,N_515);
nor U582 (N_582,N_511,N_481);
nand U583 (N_583,N_534,N_520);
nand U584 (N_584,N_504,N_535);
or U585 (N_585,N_518,N_481);
xor U586 (N_586,N_510,N_496);
nor U587 (N_587,N_518,N_522);
and U588 (N_588,N_531,N_504);
nor U589 (N_589,N_527,N_503);
and U590 (N_590,N_483,N_517);
or U591 (N_591,N_514,N_537);
nor U592 (N_592,N_525,N_493);
or U593 (N_593,N_538,N_527);
or U594 (N_594,N_509,N_499);
or U595 (N_595,N_514,N_497);
nor U596 (N_596,N_496,N_502);
or U597 (N_597,N_505,N_499);
xnor U598 (N_598,N_496,N_507);
xnor U599 (N_599,N_533,N_526);
or U600 (N_600,N_553,N_577);
xnor U601 (N_601,N_579,N_582);
or U602 (N_602,N_566,N_590);
xor U603 (N_603,N_576,N_595);
or U604 (N_604,N_587,N_567);
nor U605 (N_605,N_546,N_547);
or U606 (N_606,N_593,N_588);
or U607 (N_607,N_568,N_562);
xnor U608 (N_608,N_541,N_592);
xor U609 (N_609,N_570,N_555);
xnor U610 (N_610,N_597,N_554);
or U611 (N_611,N_544,N_540);
xnor U612 (N_612,N_575,N_550);
or U613 (N_613,N_564,N_551);
or U614 (N_614,N_543,N_594);
nor U615 (N_615,N_558,N_589);
or U616 (N_616,N_557,N_599);
nand U617 (N_617,N_552,N_585);
nand U618 (N_618,N_581,N_583);
nor U619 (N_619,N_559,N_545);
nor U620 (N_620,N_571,N_556);
nand U621 (N_621,N_584,N_548);
nand U622 (N_622,N_560,N_572);
and U623 (N_623,N_580,N_549);
or U624 (N_624,N_569,N_586);
or U625 (N_625,N_596,N_591);
and U626 (N_626,N_542,N_578);
nor U627 (N_627,N_561,N_598);
xnor U628 (N_628,N_574,N_565);
nand U629 (N_629,N_563,N_573);
or U630 (N_630,N_548,N_579);
and U631 (N_631,N_579,N_567);
nor U632 (N_632,N_593,N_586);
and U633 (N_633,N_557,N_597);
nor U634 (N_634,N_556,N_574);
xnor U635 (N_635,N_555,N_596);
and U636 (N_636,N_542,N_560);
xor U637 (N_637,N_594,N_553);
or U638 (N_638,N_598,N_557);
xnor U639 (N_639,N_541,N_561);
nor U640 (N_640,N_553,N_566);
or U641 (N_641,N_578,N_566);
nor U642 (N_642,N_571,N_555);
xnor U643 (N_643,N_591,N_594);
xnor U644 (N_644,N_587,N_545);
nor U645 (N_645,N_549,N_595);
xor U646 (N_646,N_547,N_586);
or U647 (N_647,N_579,N_549);
nor U648 (N_648,N_549,N_567);
nor U649 (N_649,N_579,N_592);
and U650 (N_650,N_588,N_560);
nand U651 (N_651,N_549,N_573);
or U652 (N_652,N_581,N_554);
and U653 (N_653,N_591,N_573);
and U654 (N_654,N_583,N_559);
or U655 (N_655,N_596,N_595);
nor U656 (N_656,N_577,N_556);
nand U657 (N_657,N_553,N_551);
nor U658 (N_658,N_595,N_579);
or U659 (N_659,N_551,N_577);
nand U660 (N_660,N_605,N_636);
and U661 (N_661,N_658,N_651);
nor U662 (N_662,N_626,N_654);
and U663 (N_663,N_615,N_655);
xnor U664 (N_664,N_645,N_601);
xnor U665 (N_665,N_618,N_607);
nand U666 (N_666,N_652,N_604);
nor U667 (N_667,N_621,N_627);
nand U668 (N_668,N_632,N_629);
nand U669 (N_669,N_617,N_634);
nand U670 (N_670,N_659,N_606);
and U671 (N_671,N_613,N_638);
and U672 (N_672,N_609,N_608);
xnor U673 (N_673,N_639,N_643);
and U674 (N_674,N_637,N_622);
xor U675 (N_675,N_653,N_624);
and U676 (N_676,N_640,N_642);
and U677 (N_677,N_603,N_631);
and U678 (N_678,N_628,N_648);
nor U679 (N_679,N_614,N_610);
nand U680 (N_680,N_641,N_616);
xnor U681 (N_681,N_623,N_656);
nor U682 (N_682,N_611,N_647);
and U683 (N_683,N_602,N_635);
or U684 (N_684,N_644,N_612);
xnor U685 (N_685,N_657,N_600);
nand U686 (N_686,N_619,N_630);
and U687 (N_687,N_650,N_620);
nor U688 (N_688,N_633,N_646);
nand U689 (N_689,N_649,N_625);
nand U690 (N_690,N_615,N_610);
and U691 (N_691,N_605,N_602);
nor U692 (N_692,N_639,N_652);
xnor U693 (N_693,N_604,N_631);
or U694 (N_694,N_614,N_640);
xnor U695 (N_695,N_655,N_625);
xnor U696 (N_696,N_622,N_651);
or U697 (N_697,N_625,N_653);
nor U698 (N_698,N_624,N_629);
xor U699 (N_699,N_614,N_649);
nand U700 (N_700,N_645,N_620);
nand U701 (N_701,N_600,N_642);
or U702 (N_702,N_635,N_625);
or U703 (N_703,N_619,N_621);
nand U704 (N_704,N_642,N_623);
or U705 (N_705,N_659,N_640);
and U706 (N_706,N_600,N_643);
xor U707 (N_707,N_622,N_623);
nand U708 (N_708,N_621,N_647);
xnor U709 (N_709,N_658,N_608);
nand U710 (N_710,N_632,N_649);
and U711 (N_711,N_624,N_613);
xnor U712 (N_712,N_604,N_623);
or U713 (N_713,N_603,N_604);
and U714 (N_714,N_604,N_644);
and U715 (N_715,N_633,N_652);
nor U716 (N_716,N_627,N_646);
xnor U717 (N_717,N_608,N_633);
and U718 (N_718,N_638,N_623);
nor U719 (N_719,N_636,N_634);
and U720 (N_720,N_682,N_694);
or U721 (N_721,N_679,N_688);
and U722 (N_722,N_665,N_713);
nor U723 (N_723,N_669,N_711);
or U724 (N_724,N_674,N_695);
or U725 (N_725,N_705,N_691);
or U726 (N_726,N_704,N_718);
or U727 (N_727,N_677,N_710);
or U728 (N_728,N_683,N_696);
nor U729 (N_729,N_701,N_703);
nor U730 (N_730,N_709,N_671);
or U731 (N_731,N_690,N_707);
xor U732 (N_732,N_667,N_708);
nand U733 (N_733,N_715,N_689);
or U734 (N_734,N_670,N_719);
nor U735 (N_735,N_684,N_716);
xnor U736 (N_736,N_706,N_676);
nand U737 (N_737,N_712,N_698);
or U738 (N_738,N_662,N_686);
nor U739 (N_739,N_660,N_664);
nand U740 (N_740,N_675,N_693);
xor U741 (N_741,N_697,N_681);
xor U742 (N_742,N_700,N_685);
or U743 (N_743,N_714,N_692);
or U744 (N_744,N_699,N_687);
nand U745 (N_745,N_666,N_680);
nor U746 (N_746,N_661,N_672);
nand U747 (N_747,N_663,N_668);
xnor U748 (N_748,N_678,N_702);
and U749 (N_749,N_673,N_717);
and U750 (N_750,N_697,N_717);
or U751 (N_751,N_710,N_664);
nor U752 (N_752,N_663,N_664);
nand U753 (N_753,N_694,N_677);
nor U754 (N_754,N_683,N_692);
nand U755 (N_755,N_719,N_672);
or U756 (N_756,N_668,N_696);
or U757 (N_757,N_712,N_681);
xor U758 (N_758,N_688,N_696);
xnor U759 (N_759,N_684,N_719);
or U760 (N_760,N_680,N_698);
or U761 (N_761,N_702,N_667);
or U762 (N_762,N_718,N_678);
xnor U763 (N_763,N_688,N_676);
and U764 (N_764,N_695,N_669);
nand U765 (N_765,N_665,N_691);
nor U766 (N_766,N_699,N_714);
xnor U767 (N_767,N_682,N_717);
nand U768 (N_768,N_675,N_716);
nand U769 (N_769,N_666,N_661);
or U770 (N_770,N_697,N_698);
nand U771 (N_771,N_679,N_665);
and U772 (N_772,N_666,N_698);
or U773 (N_773,N_684,N_691);
and U774 (N_774,N_680,N_707);
or U775 (N_775,N_694,N_712);
nor U776 (N_776,N_694,N_667);
or U777 (N_777,N_700,N_680);
nand U778 (N_778,N_719,N_680);
nor U779 (N_779,N_717,N_709);
nand U780 (N_780,N_759,N_756);
xor U781 (N_781,N_732,N_770);
and U782 (N_782,N_755,N_757);
or U783 (N_783,N_744,N_738);
and U784 (N_784,N_751,N_777);
nor U785 (N_785,N_735,N_749);
xor U786 (N_786,N_760,N_773);
xor U787 (N_787,N_771,N_731);
or U788 (N_788,N_778,N_763);
and U789 (N_789,N_758,N_723);
xnor U790 (N_790,N_721,N_727);
or U791 (N_791,N_753,N_747);
xnor U792 (N_792,N_737,N_724);
or U793 (N_793,N_761,N_746);
nor U794 (N_794,N_743,N_769);
and U795 (N_795,N_765,N_739);
nand U796 (N_796,N_776,N_775);
xnor U797 (N_797,N_734,N_766);
nor U798 (N_798,N_722,N_720);
or U799 (N_799,N_772,N_736);
xor U800 (N_800,N_725,N_748);
xnor U801 (N_801,N_752,N_764);
xor U802 (N_802,N_741,N_767);
and U803 (N_803,N_733,N_754);
xnor U804 (N_804,N_745,N_726);
and U805 (N_805,N_740,N_730);
and U806 (N_806,N_742,N_779);
or U807 (N_807,N_728,N_774);
nor U808 (N_808,N_768,N_762);
nor U809 (N_809,N_729,N_750);
and U810 (N_810,N_746,N_777);
nand U811 (N_811,N_737,N_749);
and U812 (N_812,N_754,N_752);
nor U813 (N_813,N_758,N_759);
nand U814 (N_814,N_725,N_765);
nand U815 (N_815,N_733,N_743);
nor U816 (N_816,N_722,N_768);
and U817 (N_817,N_768,N_726);
and U818 (N_818,N_773,N_737);
nor U819 (N_819,N_747,N_774);
and U820 (N_820,N_767,N_744);
xor U821 (N_821,N_773,N_755);
or U822 (N_822,N_736,N_743);
xnor U823 (N_823,N_741,N_770);
xor U824 (N_824,N_760,N_730);
or U825 (N_825,N_726,N_733);
and U826 (N_826,N_776,N_758);
nor U827 (N_827,N_754,N_759);
or U828 (N_828,N_757,N_747);
xor U829 (N_829,N_743,N_759);
nand U830 (N_830,N_778,N_769);
nand U831 (N_831,N_765,N_741);
nor U832 (N_832,N_770,N_726);
and U833 (N_833,N_760,N_744);
nor U834 (N_834,N_771,N_746);
nor U835 (N_835,N_728,N_754);
nand U836 (N_836,N_738,N_727);
nor U837 (N_837,N_726,N_753);
and U838 (N_838,N_749,N_757);
xnor U839 (N_839,N_760,N_778);
nand U840 (N_840,N_814,N_824);
or U841 (N_841,N_788,N_785);
nand U842 (N_842,N_825,N_795);
xnor U843 (N_843,N_830,N_823);
nor U844 (N_844,N_831,N_838);
or U845 (N_845,N_822,N_790);
nor U846 (N_846,N_819,N_832);
nor U847 (N_847,N_809,N_784);
or U848 (N_848,N_792,N_800);
and U849 (N_849,N_794,N_783);
nand U850 (N_850,N_837,N_839);
or U851 (N_851,N_812,N_789);
or U852 (N_852,N_793,N_816);
nand U853 (N_853,N_796,N_781);
and U854 (N_854,N_806,N_829);
nor U855 (N_855,N_780,N_786);
or U856 (N_856,N_802,N_798);
nand U857 (N_857,N_801,N_818);
or U858 (N_858,N_826,N_787);
nand U859 (N_859,N_815,N_807);
and U860 (N_860,N_782,N_799);
nand U861 (N_861,N_803,N_791);
or U862 (N_862,N_810,N_820);
nand U863 (N_863,N_808,N_821);
nor U864 (N_864,N_836,N_817);
nand U865 (N_865,N_797,N_813);
or U866 (N_866,N_804,N_835);
and U867 (N_867,N_834,N_828);
or U868 (N_868,N_827,N_805);
xor U869 (N_869,N_833,N_811);
or U870 (N_870,N_788,N_824);
or U871 (N_871,N_821,N_834);
or U872 (N_872,N_838,N_837);
xor U873 (N_873,N_797,N_819);
or U874 (N_874,N_784,N_791);
nor U875 (N_875,N_811,N_800);
nor U876 (N_876,N_811,N_837);
or U877 (N_877,N_798,N_816);
nor U878 (N_878,N_795,N_814);
nor U879 (N_879,N_809,N_804);
and U880 (N_880,N_822,N_834);
or U881 (N_881,N_839,N_814);
xor U882 (N_882,N_816,N_827);
nor U883 (N_883,N_836,N_807);
or U884 (N_884,N_802,N_805);
nand U885 (N_885,N_790,N_828);
nor U886 (N_886,N_796,N_787);
and U887 (N_887,N_814,N_796);
and U888 (N_888,N_791,N_800);
or U889 (N_889,N_808,N_813);
xnor U890 (N_890,N_828,N_813);
or U891 (N_891,N_803,N_809);
nor U892 (N_892,N_799,N_809);
or U893 (N_893,N_824,N_818);
nor U894 (N_894,N_837,N_830);
or U895 (N_895,N_828,N_789);
xor U896 (N_896,N_788,N_814);
or U897 (N_897,N_805,N_808);
or U898 (N_898,N_793,N_839);
nand U899 (N_899,N_801,N_839);
nand U900 (N_900,N_873,N_853);
xnor U901 (N_901,N_879,N_870);
and U902 (N_902,N_895,N_848);
nand U903 (N_903,N_890,N_866);
nor U904 (N_904,N_847,N_849);
or U905 (N_905,N_869,N_844);
nor U906 (N_906,N_843,N_868);
nor U907 (N_907,N_886,N_856);
xnor U908 (N_908,N_878,N_887);
nand U909 (N_909,N_855,N_851);
xnor U910 (N_910,N_889,N_841);
xnor U911 (N_911,N_884,N_876);
and U912 (N_912,N_891,N_842);
or U913 (N_913,N_854,N_877);
xnor U914 (N_914,N_885,N_894);
nand U915 (N_915,N_882,N_898);
or U916 (N_916,N_845,N_883);
nand U917 (N_917,N_874,N_871);
and U918 (N_918,N_865,N_896);
and U919 (N_919,N_892,N_861);
nand U920 (N_920,N_840,N_867);
and U921 (N_921,N_875,N_863);
or U922 (N_922,N_850,N_888);
and U923 (N_923,N_864,N_899);
nand U924 (N_924,N_860,N_893);
xor U925 (N_925,N_858,N_852);
and U926 (N_926,N_881,N_897);
or U927 (N_927,N_857,N_872);
or U928 (N_928,N_862,N_880);
or U929 (N_929,N_846,N_859);
nand U930 (N_930,N_892,N_876);
nor U931 (N_931,N_863,N_883);
or U932 (N_932,N_883,N_894);
nor U933 (N_933,N_872,N_868);
or U934 (N_934,N_848,N_866);
or U935 (N_935,N_895,N_876);
xor U936 (N_936,N_855,N_867);
nand U937 (N_937,N_893,N_888);
xnor U938 (N_938,N_844,N_897);
and U939 (N_939,N_867,N_886);
nor U940 (N_940,N_892,N_855);
and U941 (N_941,N_864,N_884);
nor U942 (N_942,N_882,N_883);
nand U943 (N_943,N_889,N_884);
and U944 (N_944,N_858,N_847);
or U945 (N_945,N_860,N_885);
nand U946 (N_946,N_855,N_876);
and U947 (N_947,N_890,N_859);
xor U948 (N_948,N_897,N_849);
nor U949 (N_949,N_859,N_843);
or U950 (N_950,N_856,N_857);
nor U951 (N_951,N_884,N_886);
xor U952 (N_952,N_843,N_889);
and U953 (N_953,N_881,N_862);
nand U954 (N_954,N_898,N_861);
and U955 (N_955,N_857,N_890);
nand U956 (N_956,N_854,N_850);
xnor U957 (N_957,N_852,N_894);
xor U958 (N_958,N_861,N_884);
nor U959 (N_959,N_865,N_840);
nand U960 (N_960,N_939,N_912);
or U961 (N_961,N_954,N_946);
xor U962 (N_962,N_900,N_933);
nor U963 (N_963,N_908,N_903);
nor U964 (N_964,N_910,N_959);
nor U965 (N_965,N_914,N_924);
or U966 (N_966,N_955,N_943);
and U967 (N_967,N_938,N_905);
and U968 (N_968,N_901,N_929);
xor U969 (N_969,N_934,N_949);
or U970 (N_970,N_928,N_948);
xor U971 (N_971,N_952,N_931);
nand U972 (N_972,N_925,N_958);
nand U973 (N_973,N_906,N_935);
or U974 (N_974,N_940,N_913);
and U975 (N_975,N_941,N_956);
nor U976 (N_976,N_942,N_915);
or U977 (N_977,N_911,N_921);
nand U978 (N_978,N_951,N_918);
nand U979 (N_979,N_922,N_904);
and U980 (N_980,N_916,N_909);
or U981 (N_981,N_937,N_927);
nand U982 (N_982,N_957,N_944);
xor U983 (N_983,N_917,N_923);
nand U984 (N_984,N_902,N_907);
or U985 (N_985,N_950,N_945);
nand U986 (N_986,N_930,N_947);
or U987 (N_987,N_936,N_953);
xor U988 (N_988,N_920,N_926);
and U989 (N_989,N_932,N_919);
xnor U990 (N_990,N_940,N_941);
and U991 (N_991,N_916,N_925);
nor U992 (N_992,N_949,N_906);
nand U993 (N_993,N_941,N_904);
and U994 (N_994,N_944,N_933);
nor U995 (N_995,N_951,N_915);
and U996 (N_996,N_918,N_904);
nor U997 (N_997,N_956,N_942);
nand U998 (N_998,N_911,N_914);
nor U999 (N_999,N_916,N_936);
nor U1000 (N_1000,N_937,N_906);
xor U1001 (N_1001,N_937,N_941);
xnor U1002 (N_1002,N_936,N_923);
nand U1003 (N_1003,N_946,N_914);
and U1004 (N_1004,N_935,N_944);
xor U1005 (N_1005,N_944,N_926);
nand U1006 (N_1006,N_930,N_923);
or U1007 (N_1007,N_922,N_926);
or U1008 (N_1008,N_923,N_955);
xor U1009 (N_1009,N_902,N_918);
and U1010 (N_1010,N_925,N_926);
nor U1011 (N_1011,N_902,N_931);
and U1012 (N_1012,N_913,N_921);
nand U1013 (N_1013,N_931,N_921);
and U1014 (N_1014,N_954,N_922);
xor U1015 (N_1015,N_936,N_920);
xnor U1016 (N_1016,N_909,N_924);
nand U1017 (N_1017,N_931,N_920);
xor U1018 (N_1018,N_908,N_920);
and U1019 (N_1019,N_905,N_906);
xnor U1020 (N_1020,N_983,N_989);
and U1021 (N_1021,N_981,N_993);
or U1022 (N_1022,N_966,N_985);
nand U1023 (N_1023,N_1001,N_970);
nor U1024 (N_1024,N_996,N_1002);
xor U1025 (N_1025,N_1017,N_972);
nor U1026 (N_1026,N_964,N_1019);
xor U1027 (N_1027,N_967,N_998);
nor U1028 (N_1028,N_1012,N_988);
nand U1029 (N_1029,N_1011,N_994);
and U1030 (N_1030,N_1013,N_969);
nor U1031 (N_1031,N_968,N_1000);
nor U1032 (N_1032,N_963,N_990);
and U1033 (N_1033,N_979,N_982);
or U1034 (N_1034,N_980,N_984);
and U1035 (N_1035,N_1004,N_992);
and U1036 (N_1036,N_987,N_1010);
nand U1037 (N_1037,N_962,N_1015);
and U1038 (N_1038,N_1018,N_975);
or U1039 (N_1039,N_1007,N_1003);
and U1040 (N_1040,N_960,N_1006);
and U1041 (N_1041,N_1016,N_1008);
or U1042 (N_1042,N_997,N_976);
nor U1043 (N_1043,N_965,N_971);
or U1044 (N_1044,N_961,N_973);
nand U1045 (N_1045,N_974,N_977);
nand U1046 (N_1046,N_978,N_1009);
nand U1047 (N_1047,N_999,N_991);
nor U1048 (N_1048,N_986,N_1014);
and U1049 (N_1049,N_995,N_1005);
nand U1050 (N_1050,N_1018,N_1011);
nand U1051 (N_1051,N_1012,N_1015);
or U1052 (N_1052,N_1000,N_1014);
xor U1053 (N_1053,N_965,N_990);
xor U1054 (N_1054,N_1002,N_993);
nand U1055 (N_1055,N_981,N_1013);
and U1056 (N_1056,N_995,N_1002);
and U1057 (N_1057,N_988,N_984);
nand U1058 (N_1058,N_969,N_1009);
nand U1059 (N_1059,N_973,N_984);
nand U1060 (N_1060,N_975,N_1007);
and U1061 (N_1061,N_984,N_1013);
nor U1062 (N_1062,N_962,N_966);
xnor U1063 (N_1063,N_1001,N_982);
xor U1064 (N_1064,N_984,N_999);
nand U1065 (N_1065,N_994,N_1002);
xnor U1066 (N_1066,N_999,N_996);
nand U1067 (N_1067,N_972,N_973);
nor U1068 (N_1068,N_991,N_1003);
nor U1069 (N_1069,N_989,N_980);
or U1070 (N_1070,N_990,N_971);
xor U1071 (N_1071,N_989,N_1007);
nand U1072 (N_1072,N_1011,N_972);
or U1073 (N_1073,N_1012,N_977);
nor U1074 (N_1074,N_965,N_980);
nor U1075 (N_1075,N_988,N_1002);
or U1076 (N_1076,N_974,N_1004);
and U1077 (N_1077,N_967,N_985);
xor U1078 (N_1078,N_995,N_991);
or U1079 (N_1079,N_996,N_973);
or U1080 (N_1080,N_1063,N_1066);
xor U1081 (N_1081,N_1035,N_1077);
nand U1082 (N_1082,N_1034,N_1045);
xnor U1083 (N_1083,N_1057,N_1067);
and U1084 (N_1084,N_1056,N_1028);
or U1085 (N_1085,N_1049,N_1076);
xor U1086 (N_1086,N_1029,N_1043);
or U1087 (N_1087,N_1041,N_1052);
and U1088 (N_1088,N_1072,N_1037);
or U1089 (N_1089,N_1046,N_1055);
xor U1090 (N_1090,N_1044,N_1059);
and U1091 (N_1091,N_1075,N_1062);
and U1092 (N_1092,N_1068,N_1050);
or U1093 (N_1093,N_1048,N_1073);
and U1094 (N_1094,N_1031,N_1033);
nor U1095 (N_1095,N_1032,N_1064);
xor U1096 (N_1096,N_1038,N_1039);
nor U1097 (N_1097,N_1023,N_1022);
nor U1098 (N_1098,N_1065,N_1054);
nor U1099 (N_1099,N_1061,N_1051);
nor U1100 (N_1100,N_1027,N_1036);
and U1101 (N_1101,N_1060,N_1020);
and U1102 (N_1102,N_1070,N_1047);
nor U1103 (N_1103,N_1025,N_1040);
and U1104 (N_1104,N_1074,N_1030);
and U1105 (N_1105,N_1021,N_1053);
nor U1106 (N_1106,N_1069,N_1024);
nand U1107 (N_1107,N_1078,N_1079);
nor U1108 (N_1108,N_1058,N_1042);
or U1109 (N_1109,N_1071,N_1026);
or U1110 (N_1110,N_1028,N_1057);
nor U1111 (N_1111,N_1029,N_1047);
and U1112 (N_1112,N_1063,N_1021);
nand U1113 (N_1113,N_1068,N_1037);
or U1114 (N_1114,N_1027,N_1060);
nor U1115 (N_1115,N_1036,N_1058);
nor U1116 (N_1116,N_1023,N_1069);
or U1117 (N_1117,N_1025,N_1034);
nor U1118 (N_1118,N_1069,N_1020);
nand U1119 (N_1119,N_1066,N_1044);
or U1120 (N_1120,N_1068,N_1032);
and U1121 (N_1121,N_1023,N_1044);
or U1122 (N_1122,N_1073,N_1023);
nand U1123 (N_1123,N_1025,N_1066);
or U1124 (N_1124,N_1064,N_1075);
and U1125 (N_1125,N_1020,N_1063);
and U1126 (N_1126,N_1021,N_1075);
nand U1127 (N_1127,N_1076,N_1070);
xnor U1128 (N_1128,N_1020,N_1058);
nor U1129 (N_1129,N_1071,N_1040);
nor U1130 (N_1130,N_1023,N_1058);
or U1131 (N_1131,N_1065,N_1071);
xnor U1132 (N_1132,N_1076,N_1042);
nand U1133 (N_1133,N_1026,N_1055);
and U1134 (N_1134,N_1033,N_1075);
or U1135 (N_1135,N_1074,N_1063);
or U1136 (N_1136,N_1053,N_1073);
and U1137 (N_1137,N_1051,N_1055);
nor U1138 (N_1138,N_1074,N_1077);
and U1139 (N_1139,N_1076,N_1050);
nand U1140 (N_1140,N_1134,N_1099);
xnor U1141 (N_1141,N_1123,N_1091);
and U1142 (N_1142,N_1121,N_1100);
or U1143 (N_1143,N_1116,N_1102);
xor U1144 (N_1144,N_1095,N_1101);
and U1145 (N_1145,N_1103,N_1084);
nor U1146 (N_1146,N_1119,N_1125);
or U1147 (N_1147,N_1089,N_1096);
and U1148 (N_1148,N_1085,N_1136);
nor U1149 (N_1149,N_1120,N_1087);
or U1150 (N_1150,N_1131,N_1113);
or U1151 (N_1151,N_1132,N_1088);
nor U1152 (N_1152,N_1092,N_1093);
and U1153 (N_1153,N_1137,N_1129);
xor U1154 (N_1154,N_1090,N_1107);
xor U1155 (N_1155,N_1104,N_1138);
xnor U1156 (N_1156,N_1108,N_1094);
nor U1157 (N_1157,N_1122,N_1115);
or U1158 (N_1158,N_1118,N_1109);
and U1159 (N_1159,N_1127,N_1135);
xor U1160 (N_1160,N_1110,N_1117);
or U1161 (N_1161,N_1097,N_1130);
nand U1162 (N_1162,N_1081,N_1083);
nand U1163 (N_1163,N_1106,N_1111);
nor U1164 (N_1164,N_1105,N_1080);
nand U1165 (N_1165,N_1098,N_1126);
nand U1166 (N_1166,N_1114,N_1086);
xnor U1167 (N_1167,N_1139,N_1124);
or U1168 (N_1168,N_1112,N_1133);
nand U1169 (N_1169,N_1082,N_1128);
nor U1170 (N_1170,N_1112,N_1124);
xnor U1171 (N_1171,N_1134,N_1114);
xor U1172 (N_1172,N_1121,N_1128);
or U1173 (N_1173,N_1132,N_1080);
nor U1174 (N_1174,N_1138,N_1118);
and U1175 (N_1175,N_1136,N_1088);
and U1176 (N_1176,N_1104,N_1110);
or U1177 (N_1177,N_1107,N_1132);
nor U1178 (N_1178,N_1114,N_1104);
xor U1179 (N_1179,N_1137,N_1119);
xnor U1180 (N_1180,N_1093,N_1111);
nand U1181 (N_1181,N_1121,N_1081);
and U1182 (N_1182,N_1129,N_1089);
xor U1183 (N_1183,N_1133,N_1134);
or U1184 (N_1184,N_1095,N_1124);
and U1185 (N_1185,N_1124,N_1105);
and U1186 (N_1186,N_1091,N_1139);
nor U1187 (N_1187,N_1085,N_1103);
nand U1188 (N_1188,N_1086,N_1109);
and U1189 (N_1189,N_1112,N_1109);
and U1190 (N_1190,N_1086,N_1110);
nor U1191 (N_1191,N_1094,N_1091);
xnor U1192 (N_1192,N_1131,N_1094);
or U1193 (N_1193,N_1137,N_1093);
or U1194 (N_1194,N_1138,N_1101);
and U1195 (N_1195,N_1139,N_1112);
nand U1196 (N_1196,N_1082,N_1120);
nand U1197 (N_1197,N_1136,N_1115);
nor U1198 (N_1198,N_1098,N_1117);
xor U1199 (N_1199,N_1110,N_1085);
nand U1200 (N_1200,N_1194,N_1190);
nand U1201 (N_1201,N_1168,N_1147);
and U1202 (N_1202,N_1178,N_1170);
or U1203 (N_1203,N_1154,N_1182);
nand U1204 (N_1204,N_1157,N_1188);
xnor U1205 (N_1205,N_1149,N_1172);
nand U1206 (N_1206,N_1158,N_1173);
or U1207 (N_1207,N_1144,N_1192);
nand U1208 (N_1208,N_1151,N_1169);
nor U1209 (N_1209,N_1153,N_1191);
nor U1210 (N_1210,N_1166,N_1165);
and U1211 (N_1211,N_1183,N_1160);
nand U1212 (N_1212,N_1142,N_1186);
nand U1213 (N_1213,N_1167,N_1141);
or U1214 (N_1214,N_1159,N_1187);
xor U1215 (N_1215,N_1152,N_1185);
nor U1216 (N_1216,N_1196,N_1179);
nand U1217 (N_1217,N_1143,N_1180);
or U1218 (N_1218,N_1181,N_1163);
and U1219 (N_1219,N_1174,N_1184);
nand U1220 (N_1220,N_1156,N_1197);
xnor U1221 (N_1221,N_1164,N_1150);
or U1222 (N_1222,N_1148,N_1171);
and U1223 (N_1223,N_1176,N_1198);
and U1224 (N_1224,N_1177,N_1155);
or U1225 (N_1225,N_1189,N_1193);
nor U1226 (N_1226,N_1140,N_1195);
nand U1227 (N_1227,N_1175,N_1199);
xnor U1228 (N_1228,N_1146,N_1162);
and U1229 (N_1229,N_1145,N_1161);
nor U1230 (N_1230,N_1146,N_1192);
and U1231 (N_1231,N_1155,N_1145);
nand U1232 (N_1232,N_1181,N_1159);
nand U1233 (N_1233,N_1166,N_1153);
xor U1234 (N_1234,N_1185,N_1145);
nor U1235 (N_1235,N_1163,N_1140);
nor U1236 (N_1236,N_1147,N_1196);
or U1237 (N_1237,N_1159,N_1158);
and U1238 (N_1238,N_1156,N_1190);
nor U1239 (N_1239,N_1177,N_1173);
xor U1240 (N_1240,N_1182,N_1174);
and U1241 (N_1241,N_1182,N_1167);
nor U1242 (N_1242,N_1193,N_1150);
or U1243 (N_1243,N_1161,N_1180);
or U1244 (N_1244,N_1179,N_1180);
xor U1245 (N_1245,N_1182,N_1152);
and U1246 (N_1246,N_1184,N_1167);
and U1247 (N_1247,N_1194,N_1178);
nor U1248 (N_1248,N_1165,N_1161);
xor U1249 (N_1249,N_1151,N_1156);
nand U1250 (N_1250,N_1185,N_1179);
and U1251 (N_1251,N_1147,N_1156);
nor U1252 (N_1252,N_1162,N_1153);
nor U1253 (N_1253,N_1145,N_1156);
or U1254 (N_1254,N_1166,N_1170);
or U1255 (N_1255,N_1140,N_1178);
or U1256 (N_1256,N_1140,N_1161);
xor U1257 (N_1257,N_1196,N_1152);
nor U1258 (N_1258,N_1195,N_1176);
xor U1259 (N_1259,N_1195,N_1193);
xnor U1260 (N_1260,N_1217,N_1208);
nand U1261 (N_1261,N_1238,N_1228);
nand U1262 (N_1262,N_1224,N_1246);
nand U1263 (N_1263,N_1241,N_1225);
and U1264 (N_1264,N_1230,N_1251);
nor U1265 (N_1265,N_1215,N_1232);
or U1266 (N_1266,N_1221,N_1209);
xor U1267 (N_1267,N_1214,N_1236);
nor U1268 (N_1268,N_1250,N_1245);
and U1269 (N_1269,N_1239,N_1212);
nor U1270 (N_1270,N_1242,N_1243);
or U1271 (N_1271,N_1255,N_1223);
xnor U1272 (N_1272,N_1220,N_1258);
and U1273 (N_1273,N_1216,N_1226);
and U1274 (N_1274,N_1253,N_1252);
and U1275 (N_1275,N_1218,N_1234);
or U1276 (N_1276,N_1207,N_1237);
or U1277 (N_1277,N_1244,N_1249);
nor U1278 (N_1278,N_1248,N_1259);
or U1279 (N_1279,N_1200,N_1213);
nand U1280 (N_1280,N_1256,N_1206);
xor U1281 (N_1281,N_1222,N_1254);
nor U1282 (N_1282,N_1210,N_1247);
nor U1283 (N_1283,N_1235,N_1229);
or U1284 (N_1284,N_1205,N_1203);
and U1285 (N_1285,N_1231,N_1257);
or U1286 (N_1286,N_1204,N_1240);
xor U1287 (N_1287,N_1219,N_1233);
nand U1288 (N_1288,N_1201,N_1202);
or U1289 (N_1289,N_1227,N_1211);
nor U1290 (N_1290,N_1218,N_1246);
nand U1291 (N_1291,N_1202,N_1218);
nor U1292 (N_1292,N_1235,N_1200);
and U1293 (N_1293,N_1248,N_1255);
xor U1294 (N_1294,N_1240,N_1213);
or U1295 (N_1295,N_1218,N_1200);
and U1296 (N_1296,N_1253,N_1223);
xnor U1297 (N_1297,N_1215,N_1245);
or U1298 (N_1298,N_1202,N_1242);
nand U1299 (N_1299,N_1241,N_1254);
nor U1300 (N_1300,N_1214,N_1212);
nor U1301 (N_1301,N_1212,N_1240);
nor U1302 (N_1302,N_1256,N_1250);
nor U1303 (N_1303,N_1256,N_1229);
nor U1304 (N_1304,N_1219,N_1240);
or U1305 (N_1305,N_1243,N_1227);
xnor U1306 (N_1306,N_1232,N_1243);
or U1307 (N_1307,N_1227,N_1221);
and U1308 (N_1308,N_1246,N_1232);
nor U1309 (N_1309,N_1201,N_1224);
nand U1310 (N_1310,N_1250,N_1213);
and U1311 (N_1311,N_1249,N_1224);
or U1312 (N_1312,N_1204,N_1206);
xor U1313 (N_1313,N_1242,N_1205);
nand U1314 (N_1314,N_1221,N_1231);
and U1315 (N_1315,N_1236,N_1211);
nand U1316 (N_1316,N_1232,N_1238);
xnor U1317 (N_1317,N_1201,N_1248);
xor U1318 (N_1318,N_1228,N_1239);
xor U1319 (N_1319,N_1240,N_1249);
and U1320 (N_1320,N_1281,N_1307);
nor U1321 (N_1321,N_1272,N_1314);
nand U1322 (N_1322,N_1296,N_1288);
xor U1323 (N_1323,N_1295,N_1306);
xnor U1324 (N_1324,N_1270,N_1278);
nand U1325 (N_1325,N_1319,N_1279);
xor U1326 (N_1326,N_1268,N_1299);
xnor U1327 (N_1327,N_1305,N_1289);
nor U1328 (N_1328,N_1318,N_1266);
xnor U1329 (N_1329,N_1264,N_1308);
nand U1330 (N_1330,N_1302,N_1277);
and U1331 (N_1331,N_1301,N_1276);
or U1332 (N_1332,N_1269,N_1315);
nand U1333 (N_1333,N_1311,N_1282);
or U1334 (N_1334,N_1316,N_1291);
and U1335 (N_1335,N_1303,N_1285);
xor U1336 (N_1336,N_1300,N_1263);
nand U1337 (N_1337,N_1283,N_1286);
or U1338 (N_1338,N_1292,N_1297);
and U1339 (N_1339,N_1312,N_1280);
and U1340 (N_1340,N_1293,N_1274);
xnor U1341 (N_1341,N_1287,N_1275);
and U1342 (N_1342,N_1294,N_1317);
xnor U1343 (N_1343,N_1273,N_1265);
nor U1344 (N_1344,N_1284,N_1310);
and U1345 (N_1345,N_1271,N_1309);
or U1346 (N_1346,N_1267,N_1304);
nor U1347 (N_1347,N_1260,N_1290);
or U1348 (N_1348,N_1261,N_1313);
xnor U1349 (N_1349,N_1298,N_1262);
or U1350 (N_1350,N_1269,N_1286);
nand U1351 (N_1351,N_1319,N_1263);
nor U1352 (N_1352,N_1262,N_1278);
xnor U1353 (N_1353,N_1302,N_1310);
nand U1354 (N_1354,N_1262,N_1282);
nand U1355 (N_1355,N_1291,N_1318);
or U1356 (N_1356,N_1292,N_1268);
or U1357 (N_1357,N_1315,N_1316);
nor U1358 (N_1358,N_1262,N_1311);
and U1359 (N_1359,N_1279,N_1288);
nand U1360 (N_1360,N_1308,N_1305);
nand U1361 (N_1361,N_1300,N_1271);
nand U1362 (N_1362,N_1310,N_1319);
xor U1363 (N_1363,N_1306,N_1303);
and U1364 (N_1364,N_1299,N_1293);
nand U1365 (N_1365,N_1264,N_1303);
nor U1366 (N_1366,N_1293,N_1308);
or U1367 (N_1367,N_1270,N_1312);
nor U1368 (N_1368,N_1302,N_1272);
or U1369 (N_1369,N_1286,N_1305);
nor U1370 (N_1370,N_1304,N_1289);
or U1371 (N_1371,N_1305,N_1317);
xor U1372 (N_1372,N_1267,N_1297);
or U1373 (N_1373,N_1288,N_1309);
xor U1374 (N_1374,N_1302,N_1316);
or U1375 (N_1375,N_1271,N_1297);
nand U1376 (N_1376,N_1293,N_1285);
or U1377 (N_1377,N_1315,N_1287);
nor U1378 (N_1378,N_1274,N_1263);
and U1379 (N_1379,N_1298,N_1272);
nand U1380 (N_1380,N_1329,N_1345);
nand U1381 (N_1381,N_1373,N_1374);
nand U1382 (N_1382,N_1356,N_1333);
xor U1383 (N_1383,N_1342,N_1353);
xor U1384 (N_1384,N_1322,N_1339);
or U1385 (N_1385,N_1320,N_1341);
xor U1386 (N_1386,N_1351,N_1344);
nand U1387 (N_1387,N_1375,N_1334);
or U1388 (N_1388,N_1323,N_1324);
nand U1389 (N_1389,N_1364,N_1348);
nor U1390 (N_1390,N_1365,N_1368);
nor U1391 (N_1391,N_1369,N_1378);
and U1392 (N_1392,N_1326,N_1360);
nand U1393 (N_1393,N_1371,N_1338);
and U1394 (N_1394,N_1367,N_1332);
nand U1395 (N_1395,N_1328,N_1346);
or U1396 (N_1396,N_1379,N_1327);
and U1397 (N_1397,N_1330,N_1336);
and U1398 (N_1398,N_1370,N_1335);
or U1399 (N_1399,N_1337,N_1361);
or U1400 (N_1400,N_1376,N_1366);
or U1401 (N_1401,N_1362,N_1377);
nand U1402 (N_1402,N_1357,N_1372);
nor U1403 (N_1403,N_1331,N_1343);
nand U1404 (N_1404,N_1363,N_1321);
or U1405 (N_1405,N_1354,N_1340);
and U1406 (N_1406,N_1349,N_1359);
nand U1407 (N_1407,N_1352,N_1355);
or U1408 (N_1408,N_1358,N_1350);
nor U1409 (N_1409,N_1347,N_1325);
and U1410 (N_1410,N_1365,N_1355);
and U1411 (N_1411,N_1331,N_1351);
nand U1412 (N_1412,N_1345,N_1363);
xor U1413 (N_1413,N_1322,N_1374);
nor U1414 (N_1414,N_1352,N_1322);
or U1415 (N_1415,N_1336,N_1374);
xor U1416 (N_1416,N_1345,N_1339);
or U1417 (N_1417,N_1369,N_1350);
or U1418 (N_1418,N_1352,N_1363);
nor U1419 (N_1419,N_1331,N_1340);
nor U1420 (N_1420,N_1338,N_1350);
nand U1421 (N_1421,N_1334,N_1341);
xor U1422 (N_1422,N_1349,N_1343);
and U1423 (N_1423,N_1359,N_1322);
nor U1424 (N_1424,N_1358,N_1328);
nand U1425 (N_1425,N_1377,N_1330);
and U1426 (N_1426,N_1379,N_1373);
and U1427 (N_1427,N_1369,N_1365);
and U1428 (N_1428,N_1324,N_1325);
nand U1429 (N_1429,N_1337,N_1351);
xnor U1430 (N_1430,N_1322,N_1325);
and U1431 (N_1431,N_1358,N_1376);
xor U1432 (N_1432,N_1372,N_1343);
and U1433 (N_1433,N_1352,N_1376);
nand U1434 (N_1434,N_1359,N_1372);
nor U1435 (N_1435,N_1329,N_1339);
nor U1436 (N_1436,N_1343,N_1358);
or U1437 (N_1437,N_1333,N_1360);
or U1438 (N_1438,N_1335,N_1377);
and U1439 (N_1439,N_1356,N_1350);
nand U1440 (N_1440,N_1381,N_1422);
nor U1441 (N_1441,N_1394,N_1424);
nor U1442 (N_1442,N_1415,N_1399);
and U1443 (N_1443,N_1433,N_1404);
nor U1444 (N_1444,N_1421,N_1416);
or U1445 (N_1445,N_1438,N_1405);
nand U1446 (N_1446,N_1393,N_1407);
and U1447 (N_1447,N_1382,N_1401);
and U1448 (N_1448,N_1423,N_1396);
xor U1449 (N_1449,N_1386,N_1437);
nor U1450 (N_1450,N_1380,N_1390);
xnor U1451 (N_1451,N_1431,N_1419);
and U1452 (N_1452,N_1397,N_1383);
and U1453 (N_1453,N_1414,N_1395);
xor U1454 (N_1454,N_1426,N_1406);
xnor U1455 (N_1455,N_1411,N_1418);
or U1456 (N_1456,N_1435,N_1417);
nor U1457 (N_1457,N_1409,N_1408);
nor U1458 (N_1458,N_1402,N_1432);
nor U1459 (N_1459,N_1420,N_1388);
or U1460 (N_1460,N_1439,N_1410);
and U1461 (N_1461,N_1392,N_1429);
nand U1462 (N_1462,N_1384,N_1430);
nand U1463 (N_1463,N_1427,N_1436);
or U1464 (N_1464,N_1403,N_1413);
xnor U1465 (N_1465,N_1400,N_1398);
and U1466 (N_1466,N_1389,N_1434);
nand U1467 (N_1467,N_1385,N_1412);
and U1468 (N_1468,N_1391,N_1428);
nand U1469 (N_1469,N_1425,N_1387);
nand U1470 (N_1470,N_1398,N_1380);
or U1471 (N_1471,N_1384,N_1394);
and U1472 (N_1472,N_1433,N_1438);
nor U1473 (N_1473,N_1394,N_1405);
or U1474 (N_1474,N_1381,N_1426);
nand U1475 (N_1475,N_1413,N_1401);
nor U1476 (N_1476,N_1389,N_1394);
or U1477 (N_1477,N_1395,N_1396);
nor U1478 (N_1478,N_1385,N_1425);
xor U1479 (N_1479,N_1403,N_1412);
xnor U1480 (N_1480,N_1410,N_1399);
xor U1481 (N_1481,N_1426,N_1407);
nand U1482 (N_1482,N_1382,N_1407);
nand U1483 (N_1483,N_1437,N_1436);
nor U1484 (N_1484,N_1384,N_1393);
nand U1485 (N_1485,N_1427,N_1385);
nand U1486 (N_1486,N_1382,N_1391);
or U1487 (N_1487,N_1381,N_1424);
and U1488 (N_1488,N_1428,N_1407);
nand U1489 (N_1489,N_1423,N_1439);
and U1490 (N_1490,N_1422,N_1438);
xor U1491 (N_1491,N_1415,N_1405);
and U1492 (N_1492,N_1390,N_1425);
nor U1493 (N_1493,N_1380,N_1404);
and U1494 (N_1494,N_1397,N_1401);
or U1495 (N_1495,N_1388,N_1404);
nor U1496 (N_1496,N_1400,N_1381);
xor U1497 (N_1497,N_1416,N_1411);
nor U1498 (N_1498,N_1398,N_1439);
and U1499 (N_1499,N_1395,N_1389);
or U1500 (N_1500,N_1479,N_1471);
nor U1501 (N_1501,N_1470,N_1454);
nor U1502 (N_1502,N_1467,N_1457);
and U1503 (N_1503,N_1477,N_1494);
or U1504 (N_1504,N_1469,N_1492);
and U1505 (N_1505,N_1476,N_1495);
xor U1506 (N_1506,N_1450,N_1486);
xor U1507 (N_1507,N_1498,N_1466);
and U1508 (N_1508,N_1488,N_1474);
nor U1509 (N_1509,N_1484,N_1458);
or U1510 (N_1510,N_1460,N_1455);
and U1511 (N_1511,N_1480,N_1489);
or U1512 (N_1512,N_1468,N_1440);
or U1513 (N_1513,N_1445,N_1473);
nand U1514 (N_1514,N_1478,N_1463);
nand U1515 (N_1515,N_1496,N_1491);
nor U1516 (N_1516,N_1487,N_1448);
and U1517 (N_1517,N_1446,N_1485);
and U1518 (N_1518,N_1482,N_1441);
or U1519 (N_1519,N_1456,N_1447);
xnor U1520 (N_1520,N_1483,N_1499);
nand U1521 (N_1521,N_1451,N_1472);
xor U1522 (N_1522,N_1490,N_1453);
or U1523 (N_1523,N_1443,N_1462);
and U1524 (N_1524,N_1465,N_1461);
xnor U1525 (N_1525,N_1459,N_1444);
and U1526 (N_1526,N_1449,N_1442);
nand U1527 (N_1527,N_1475,N_1493);
nor U1528 (N_1528,N_1497,N_1464);
xnor U1529 (N_1529,N_1481,N_1452);
and U1530 (N_1530,N_1450,N_1442);
xnor U1531 (N_1531,N_1463,N_1441);
and U1532 (N_1532,N_1464,N_1490);
nand U1533 (N_1533,N_1457,N_1481);
and U1534 (N_1534,N_1475,N_1457);
nand U1535 (N_1535,N_1493,N_1490);
xnor U1536 (N_1536,N_1452,N_1485);
and U1537 (N_1537,N_1441,N_1495);
nor U1538 (N_1538,N_1471,N_1490);
and U1539 (N_1539,N_1476,N_1491);
or U1540 (N_1540,N_1497,N_1443);
and U1541 (N_1541,N_1490,N_1462);
and U1542 (N_1542,N_1451,N_1454);
nand U1543 (N_1543,N_1478,N_1454);
or U1544 (N_1544,N_1471,N_1448);
and U1545 (N_1545,N_1498,N_1453);
nor U1546 (N_1546,N_1457,N_1451);
or U1547 (N_1547,N_1479,N_1483);
nor U1548 (N_1548,N_1486,N_1443);
nor U1549 (N_1549,N_1496,N_1456);
xor U1550 (N_1550,N_1445,N_1484);
or U1551 (N_1551,N_1487,N_1454);
nor U1552 (N_1552,N_1441,N_1473);
nor U1553 (N_1553,N_1486,N_1470);
and U1554 (N_1554,N_1476,N_1498);
xor U1555 (N_1555,N_1492,N_1462);
nor U1556 (N_1556,N_1495,N_1497);
nand U1557 (N_1557,N_1462,N_1450);
xor U1558 (N_1558,N_1472,N_1488);
nand U1559 (N_1559,N_1456,N_1444);
and U1560 (N_1560,N_1521,N_1544);
or U1561 (N_1561,N_1530,N_1519);
or U1562 (N_1562,N_1547,N_1503);
xor U1563 (N_1563,N_1552,N_1558);
nand U1564 (N_1564,N_1505,N_1548);
nand U1565 (N_1565,N_1529,N_1536);
xor U1566 (N_1566,N_1534,N_1516);
nand U1567 (N_1567,N_1540,N_1538);
nand U1568 (N_1568,N_1506,N_1512);
nand U1569 (N_1569,N_1518,N_1510);
or U1570 (N_1570,N_1556,N_1522);
nor U1571 (N_1571,N_1524,N_1500);
nand U1572 (N_1572,N_1541,N_1502);
and U1573 (N_1573,N_1511,N_1537);
nand U1574 (N_1574,N_1520,N_1532);
nor U1575 (N_1575,N_1555,N_1514);
xnor U1576 (N_1576,N_1523,N_1554);
nor U1577 (N_1577,N_1531,N_1528);
nand U1578 (N_1578,N_1517,N_1549);
xnor U1579 (N_1579,N_1553,N_1539);
and U1580 (N_1580,N_1545,N_1546);
nand U1581 (N_1581,N_1501,N_1504);
nor U1582 (N_1582,N_1526,N_1515);
or U1583 (N_1583,N_1527,N_1525);
nand U1584 (N_1584,N_1513,N_1535);
xnor U1585 (N_1585,N_1508,N_1533);
xor U1586 (N_1586,N_1543,N_1559);
and U1587 (N_1587,N_1509,N_1557);
nor U1588 (N_1588,N_1551,N_1507);
or U1589 (N_1589,N_1550,N_1542);
and U1590 (N_1590,N_1511,N_1541);
nand U1591 (N_1591,N_1514,N_1527);
xnor U1592 (N_1592,N_1505,N_1518);
nand U1593 (N_1593,N_1506,N_1534);
or U1594 (N_1594,N_1557,N_1508);
xnor U1595 (N_1595,N_1533,N_1507);
nand U1596 (N_1596,N_1500,N_1557);
or U1597 (N_1597,N_1523,N_1525);
nand U1598 (N_1598,N_1541,N_1559);
and U1599 (N_1599,N_1552,N_1500);
xnor U1600 (N_1600,N_1522,N_1524);
xor U1601 (N_1601,N_1552,N_1550);
nand U1602 (N_1602,N_1541,N_1530);
or U1603 (N_1603,N_1537,N_1512);
nand U1604 (N_1604,N_1505,N_1553);
and U1605 (N_1605,N_1507,N_1557);
xor U1606 (N_1606,N_1505,N_1552);
or U1607 (N_1607,N_1531,N_1548);
or U1608 (N_1608,N_1527,N_1532);
and U1609 (N_1609,N_1542,N_1546);
and U1610 (N_1610,N_1527,N_1543);
xor U1611 (N_1611,N_1502,N_1519);
or U1612 (N_1612,N_1532,N_1547);
nand U1613 (N_1613,N_1506,N_1547);
xnor U1614 (N_1614,N_1512,N_1528);
and U1615 (N_1615,N_1503,N_1544);
nor U1616 (N_1616,N_1558,N_1506);
nor U1617 (N_1617,N_1546,N_1541);
xor U1618 (N_1618,N_1556,N_1534);
nand U1619 (N_1619,N_1512,N_1543);
nand U1620 (N_1620,N_1599,N_1575);
and U1621 (N_1621,N_1563,N_1617);
nor U1622 (N_1622,N_1614,N_1576);
and U1623 (N_1623,N_1562,N_1596);
nor U1624 (N_1624,N_1604,N_1593);
nand U1625 (N_1625,N_1589,N_1588);
nand U1626 (N_1626,N_1597,N_1608);
xor U1627 (N_1627,N_1618,N_1602);
and U1628 (N_1628,N_1610,N_1619);
or U1629 (N_1629,N_1565,N_1587);
or U1630 (N_1630,N_1571,N_1598);
or U1631 (N_1631,N_1564,N_1581);
nor U1632 (N_1632,N_1573,N_1560);
nand U1633 (N_1633,N_1561,N_1594);
and U1634 (N_1634,N_1591,N_1605);
or U1635 (N_1635,N_1580,N_1612);
and U1636 (N_1636,N_1574,N_1567);
or U1637 (N_1637,N_1582,N_1600);
and U1638 (N_1638,N_1577,N_1585);
and U1639 (N_1639,N_1616,N_1568);
nand U1640 (N_1640,N_1613,N_1603);
nor U1641 (N_1641,N_1578,N_1606);
nor U1642 (N_1642,N_1609,N_1584);
or U1643 (N_1643,N_1579,N_1572);
and U1644 (N_1644,N_1566,N_1583);
or U1645 (N_1645,N_1601,N_1570);
or U1646 (N_1646,N_1615,N_1569);
nor U1647 (N_1647,N_1586,N_1595);
and U1648 (N_1648,N_1592,N_1590);
nor U1649 (N_1649,N_1607,N_1611);
and U1650 (N_1650,N_1618,N_1614);
xnor U1651 (N_1651,N_1593,N_1565);
nor U1652 (N_1652,N_1611,N_1610);
xnor U1653 (N_1653,N_1614,N_1560);
nor U1654 (N_1654,N_1573,N_1592);
and U1655 (N_1655,N_1561,N_1603);
xnor U1656 (N_1656,N_1614,N_1602);
or U1657 (N_1657,N_1575,N_1613);
nor U1658 (N_1658,N_1612,N_1588);
and U1659 (N_1659,N_1567,N_1569);
or U1660 (N_1660,N_1579,N_1610);
nor U1661 (N_1661,N_1610,N_1572);
nand U1662 (N_1662,N_1576,N_1607);
nor U1663 (N_1663,N_1615,N_1575);
xor U1664 (N_1664,N_1591,N_1600);
or U1665 (N_1665,N_1586,N_1577);
and U1666 (N_1666,N_1592,N_1601);
xor U1667 (N_1667,N_1585,N_1590);
and U1668 (N_1668,N_1613,N_1605);
or U1669 (N_1669,N_1565,N_1603);
nor U1670 (N_1670,N_1583,N_1613);
nor U1671 (N_1671,N_1575,N_1611);
xnor U1672 (N_1672,N_1569,N_1587);
nor U1673 (N_1673,N_1597,N_1561);
xnor U1674 (N_1674,N_1574,N_1595);
nor U1675 (N_1675,N_1583,N_1594);
or U1676 (N_1676,N_1571,N_1604);
xor U1677 (N_1677,N_1576,N_1596);
nor U1678 (N_1678,N_1567,N_1607);
xnor U1679 (N_1679,N_1572,N_1560);
nand U1680 (N_1680,N_1677,N_1627);
xor U1681 (N_1681,N_1629,N_1660);
nor U1682 (N_1682,N_1626,N_1650);
or U1683 (N_1683,N_1645,N_1663);
or U1684 (N_1684,N_1621,N_1678);
or U1685 (N_1685,N_1649,N_1679);
or U1686 (N_1686,N_1671,N_1638);
or U1687 (N_1687,N_1632,N_1653);
and U1688 (N_1688,N_1672,N_1646);
xor U1689 (N_1689,N_1659,N_1637);
and U1690 (N_1690,N_1652,N_1647);
xor U1691 (N_1691,N_1639,N_1658);
and U1692 (N_1692,N_1676,N_1623);
nand U1693 (N_1693,N_1664,N_1643);
or U1694 (N_1694,N_1675,N_1670);
and U1695 (N_1695,N_1674,N_1642);
nand U1696 (N_1696,N_1655,N_1636);
or U1697 (N_1697,N_1631,N_1641);
and U1698 (N_1698,N_1662,N_1668);
xnor U1699 (N_1699,N_1644,N_1656);
nand U1700 (N_1700,N_1657,N_1635);
nor U1701 (N_1701,N_1673,N_1628);
xnor U1702 (N_1702,N_1624,N_1648);
nand U1703 (N_1703,N_1661,N_1634);
nand U1704 (N_1704,N_1625,N_1622);
or U1705 (N_1705,N_1630,N_1666);
and U1706 (N_1706,N_1620,N_1669);
nand U1707 (N_1707,N_1633,N_1651);
nand U1708 (N_1708,N_1665,N_1667);
xnor U1709 (N_1709,N_1654,N_1640);
or U1710 (N_1710,N_1655,N_1633);
nor U1711 (N_1711,N_1641,N_1665);
and U1712 (N_1712,N_1639,N_1666);
and U1713 (N_1713,N_1657,N_1636);
and U1714 (N_1714,N_1678,N_1648);
xnor U1715 (N_1715,N_1626,N_1636);
nand U1716 (N_1716,N_1666,N_1636);
nand U1717 (N_1717,N_1633,N_1670);
nor U1718 (N_1718,N_1659,N_1668);
nor U1719 (N_1719,N_1677,N_1651);
or U1720 (N_1720,N_1668,N_1673);
and U1721 (N_1721,N_1670,N_1664);
xnor U1722 (N_1722,N_1632,N_1645);
xor U1723 (N_1723,N_1675,N_1674);
xor U1724 (N_1724,N_1633,N_1632);
nor U1725 (N_1725,N_1637,N_1669);
or U1726 (N_1726,N_1637,N_1643);
xor U1727 (N_1727,N_1652,N_1649);
or U1728 (N_1728,N_1620,N_1628);
and U1729 (N_1729,N_1671,N_1627);
or U1730 (N_1730,N_1678,N_1620);
and U1731 (N_1731,N_1643,N_1634);
and U1732 (N_1732,N_1629,N_1651);
xor U1733 (N_1733,N_1637,N_1672);
and U1734 (N_1734,N_1673,N_1622);
and U1735 (N_1735,N_1642,N_1630);
or U1736 (N_1736,N_1678,N_1643);
xor U1737 (N_1737,N_1641,N_1643);
and U1738 (N_1738,N_1679,N_1620);
or U1739 (N_1739,N_1642,N_1671);
or U1740 (N_1740,N_1719,N_1704);
nor U1741 (N_1741,N_1705,N_1710);
and U1742 (N_1742,N_1688,N_1696);
and U1743 (N_1743,N_1715,N_1697);
or U1744 (N_1744,N_1707,N_1702);
xnor U1745 (N_1745,N_1722,N_1725);
or U1746 (N_1746,N_1735,N_1689);
and U1747 (N_1747,N_1712,N_1723);
nand U1748 (N_1748,N_1701,N_1693);
or U1749 (N_1749,N_1730,N_1734);
nand U1750 (N_1750,N_1739,N_1721);
nand U1751 (N_1751,N_1681,N_1720);
nor U1752 (N_1752,N_1709,N_1718);
or U1753 (N_1753,N_1727,N_1713);
xor U1754 (N_1754,N_1683,N_1711);
xor U1755 (N_1755,N_1690,N_1698);
or U1756 (N_1756,N_1724,N_1694);
xor U1757 (N_1757,N_1680,N_1706);
and U1758 (N_1758,N_1717,N_1708);
nor U1759 (N_1759,N_1728,N_1733);
xnor U1760 (N_1760,N_1691,N_1737);
and U1761 (N_1761,N_1686,N_1687);
xnor U1762 (N_1762,N_1736,N_1703);
nand U1763 (N_1763,N_1738,N_1684);
and U1764 (N_1764,N_1714,N_1699);
and U1765 (N_1765,N_1685,N_1729);
and U1766 (N_1766,N_1731,N_1732);
and U1767 (N_1767,N_1700,N_1682);
xnor U1768 (N_1768,N_1692,N_1726);
nand U1769 (N_1769,N_1716,N_1695);
nor U1770 (N_1770,N_1694,N_1692);
or U1771 (N_1771,N_1727,N_1711);
and U1772 (N_1772,N_1730,N_1720);
and U1773 (N_1773,N_1703,N_1729);
or U1774 (N_1774,N_1710,N_1685);
and U1775 (N_1775,N_1725,N_1697);
nor U1776 (N_1776,N_1709,N_1686);
or U1777 (N_1777,N_1726,N_1709);
and U1778 (N_1778,N_1718,N_1729);
and U1779 (N_1779,N_1720,N_1698);
nor U1780 (N_1780,N_1715,N_1681);
nor U1781 (N_1781,N_1705,N_1691);
xnor U1782 (N_1782,N_1684,N_1698);
and U1783 (N_1783,N_1698,N_1722);
and U1784 (N_1784,N_1695,N_1688);
nor U1785 (N_1785,N_1684,N_1680);
and U1786 (N_1786,N_1715,N_1710);
and U1787 (N_1787,N_1734,N_1719);
and U1788 (N_1788,N_1697,N_1732);
nor U1789 (N_1789,N_1729,N_1698);
and U1790 (N_1790,N_1708,N_1709);
and U1791 (N_1791,N_1709,N_1724);
and U1792 (N_1792,N_1726,N_1719);
nor U1793 (N_1793,N_1732,N_1700);
nor U1794 (N_1794,N_1733,N_1720);
xnor U1795 (N_1795,N_1722,N_1690);
nand U1796 (N_1796,N_1701,N_1681);
xnor U1797 (N_1797,N_1715,N_1692);
xor U1798 (N_1798,N_1723,N_1683);
or U1799 (N_1799,N_1719,N_1681);
nand U1800 (N_1800,N_1761,N_1799);
and U1801 (N_1801,N_1775,N_1780);
nand U1802 (N_1802,N_1789,N_1753);
nor U1803 (N_1803,N_1765,N_1746);
nand U1804 (N_1804,N_1791,N_1741);
nor U1805 (N_1805,N_1792,N_1784);
xor U1806 (N_1806,N_1759,N_1794);
or U1807 (N_1807,N_1755,N_1785);
xor U1808 (N_1808,N_1787,N_1773);
nor U1809 (N_1809,N_1790,N_1786);
or U1810 (N_1810,N_1772,N_1793);
xor U1811 (N_1811,N_1744,N_1742);
or U1812 (N_1812,N_1764,N_1779);
or U1813 (N_1813,N_1781,N_1777);
and U1814 (N_1814,N_1783,N_1796);
and U1815 (N_1815,N_1747,N_1776);
nor U1816 (N_1816,N_1743,N_1752);
nand U1817 (N_1817,N_1757,N_1750);
nor U1818 (N_1818,N_1751,N_1762);
or U1819 (N_1819,N_1740,N_1748);
and U1820 (N_1820,N_1778,N_1758);
nor U1821 (N_1821,N_1770,N_1771);
or U1822 (N_1822,N_1745,N_1756);
nor U1823 (N_1823,N_1766,N_1795);
or U1824 (N_1824,N_1763,N_1769);
or U1825 (N_1825,N_1754,N_1798);
xor U1826 (N_1826,N_1774,N_1760);
xor U1827 (N_1827,N_1788,N_1767);
and U1828 (N_1828,N_1797,N_1782);
xor U1829 (N_1829,N_1749,N_1768);
nor U1830 (N_1830,N_1761,N_1765);
and U1831 (N_1831,N_1786,N_1772);
nand U1832 (N_1832,N_1791,N_1788);
nand U1833 (N_1833,N_1783,N_1759);
and U1834 (N_1834,N_1750,N_1793);
or U1835 (N_1835,N_1754,N_1783);
or U1836 (N_1836,N_1789,N_1761);
nand U1837 (N_1837,N_1792,N_1787);
nand U1838 (N_1838,N_1795,N_1785);
xnor U1839 (N_1839,N_1774,N_1799);
or U1840 (N_1840,N_1767,N_1773);
nand U1841 (N_1841,N_1758,N_1763);
xor U1842 (N_1842,N_1741,N_1783);
or U1843 (N_1843,N_1773,N_1782);
nand U1844 (N_1844,N_1794,N_1792);
and U1845 (N_1845,N_1763,N_1783);
or U1846 (N_1846,N_1779,N_1752);
nand U1847 (N_1847,N_1743,N_1751);
xor U1848 (N_1848,N_1751,N_1775);
and U1849 (N_1849,N_1792,N_1765);
xnor U1850 (N_1850,N_1780,N_1779);
nand U1851 (N_1851,N_1763,N_1748);
and U1852 (N_1852,N_1754,N_1794);
xnor U1853 (N_1853,N_1764,N_1760);
nand U1854 (N_1854,N_1757,N_1794);
or U1855 (N_1855,N_1758,N_1745);
xnor U1856 (N_1856,N_1760,N_1770);
or U1857 (N_1857,N_1776,N_1755);
and U1858 (N_1858,N_1755,N_1798);
or U1859 (N_1859,N_1786,N_1751);
and U1860 (N_1860,N_1833,N_1832);
nor U1861 (N_1861,N_1807,N_1853);
nor U1862 (N_1862,N_1835,N_1851);
nand U1863 (N_1863,N_1803,N_1849);
nand U1864 (N_1864,N_1815,N_1800);
nand U1865 (N_1865,N_1856,N_1822);
xor U1866 (N_1866,N_1852,N_1841);
nor U1867 (N_1867,N_1823,N_1811);
nor U1868 (N_1868,N_1837,N_1844);
xnor U1869 (N_1869,N_1812,N_1810);
nand U1870 (N_1870,N_1805,N_1829);
nand U1871 (N_1871,N_1821,N_1806);
or U1872 (N_1872,N_1834,N_1857);
and U1873 (N_1873,N_1858,N_1839);
nand U1874 (N_1874,N_1859,N_1828);
nor U1875 (N_1875,N_1814,N_1850);
nor U1876 (N_1876,N_1840,N_1820);
nand U1877 (N_1877,N_1804,N_1831);
and U1878 (N_1878,N_1826,N_1842);
or U1879 (N_1879,N_1830,N_1854);
or U1880 (N_1880,N_1845,N_1809);
nand U1881 (N_1881,N_1813,N_1843);
and U1882 (N_1882,N_1817,N_1846);
nor U1883 (N_1883,N_1836,N_1801);
nand U1884 (N_1884,N_1816,N_1802);
nand U1885 (N_1885,N_1825,N_1847);
nand U1886 (N_1886,N_1808,N_1838);
and U1887 (N_1887,N_1824,N_1819);
or U1888 (N_1888,N_1818,N_1827);
or U1889 (N_1889,N_1848,N_1855);
or U1890 (N_1890,N_1845,N_1814);
nand U1891 (N_1891,N_1850,N_1842);
xnor U1892 (N_1892,N_1831,N_1809);
or U1893 (N_1893,N_1814,N_1811);
or U1894 (N_1894,N_1836,N_1857);
nand U1895 (N_1895,N_1802,N_1851);
nor U1896 (N_1896,N_1807,N_1834);
xnor U1897 (N_1897,N_1827,N_1821);
xor U1898 (N_1898,N_1804,N_1849);
nand U1899 (N_1899,N_1809,N_1815);
and U1900 (N_1900,N_1829,N_1841);
or U1901 (N_1901,N_1826,N_1808);
nor U1902 (N_1902,N_1849,N_1855);
nand U1903 (N_1903,N_1830,N_1829);
nand U1904 (N_1904,N_1855,N_1836);
nand U1905 (N_1905,N_1849,N_1856);
nand U1906 (N_1906,N_1830,N_1832);
nand U1907 (N_1907,N_1811,N_1810);
or U1908 (N_1908,N_1855,N_1830);
or U1909 (N_1909,N_1844,N_1811);
xnor U1910 (N_1910,N_1806,N_1812);
xnor U1911 (N_1911,N_1802,N_1846);
and U1912 (N_1912,N_1807,N_1830);
xnor U1913 (N_1913,N_1831,N_1843);
and U1914 (N_1914,N_1815,N_1822);
nand U1915 (N_1915,N_1831,N_1855);
nand U1916 (N_1916,N_1856,N_1830);
nor U1917 (N_1917,N_1843,N_1851);
or U1918 (N_1918,N_1811,N_1834);
and U1919 (N_1919,N_1839,N_1856);
or U1920 (N_1920,N_1885,N_1877);
xnor U1921 (N_1921,N_1887,N_1881);
nor U1922 (N_1922,N_1916,N_1914);
nand U1923 (N_1923,N_1893,N_1898);
or U1924 (N_1924,N_1876,N_1896);
nor U1925 (N_1925,N_1913,N_1905);
nor U1926 (N_1926,N_1908,N_1912);
nand U1927 (N_1927,N_1875,N_1904);
nor U1928 (N_1928,N_1910,N_1889);
and U1929 (N_1929,N_1918,N_1907);
nor U1930 (N_1930,N_1892,N_1873);
xnor U1931 (N_1931,N_1872,N_1891);
or U1932 (N_1932,N_1878,N_1864);
or U1933 (N_1933,N_1894,N_1915);
and U1934 (N_1934,N_1874,N_1902);
xor U1935 (N_1935,N_1862,N_1884);
and U1936 (N_1936,N_1897,N_1900);
or U1937 (N_1937,N_1906,N_1870);
and U1938 (N_1938,N_1890,N_1865);
nor U1939 (N_1939,N_1903,N_1860);
nor U1940 (N_1940,N_1919,N_1868);
and U1941 (N_1941,N_1917,N_1879);
xor U1942 (N_1942,N_1883,N_1869);
nand U1943 (N_1943,N_1895,N_1911);
or U1944 (N_1944,N_1886,N_1861);
nand U1945 (N_1945,N_1888,N_1867);
xnor U1946 (N_1946,N_1880,N_1863);
xor U1947 (N_1947,N_1866,N_1871);
xnor U1948 (N_1948,N_1882,N_1909);
nand U1949 (N_1949,N_1899,N_1901);
or U1950 (N_1950,N_1911,N_1903);
nor U1951 (N_1951,N_1873,N_1886);
nand U1952 (N_1952,N_1902,N_1897);
and U1953 (N_1953,N_1884,N_1865);
or U1954 (N_1954,N_1877,N_1864);
or U1955 (N_1955,N_1881,N_1902);
nand U1956 (N_1956,N_1878,N_1906);
nor U1957 (N_1957,N_1901,N_1893);
or U1958 (N_1958,N_1901,N_1881);
or U1959 (N_1959,N_1874,N_1861);
xor U1960 (N_1960,N_1915,N_1916);
nor U1961 (N_1961,N_1895,N_1901);
xor U1962 (N_1962,N_1886,N_1868);
nand U1963 (N_1963,N_1912,N_1895);
nand U1964 (N_1964,N_1887,N_1873);
xor U1965 (N_1965,N_1917,N_1906);
or U1966 (N_1966,N_1904,N_1880);
and U1967 (N_1967,N_1881,N_1873);
nor U1968 (N_1968,N_1871,N_1902);
nor U1969 (N_1969,N_1900,N_1871);
nor U1970 (N_1970,N_1862,N_1900);
nand U1971 (N_1971,N_1908,N_1888);
xnor U1972 (N_1972,N_1874,N_1888);
and U1973 (N_1973,N_1916,N_1902);
nand U1974 (N_1974,N_1891,N_1886);
nand U1975 (N_1975,N_1902,N_1878);
or U1976 (N_1976,N_1910,N_1919);
nand U1977 (N_1977,N_1904,N_1906);
or U1978 (N_1978,N_1915,N_1913);
or U1979 (N_1979,N_1915,N_1869);
nor U1980 (N_1980,N_1939,N_1930);
nand U1981 (N_1981,N_1948,N_1977);
nor U1982 (N_1982,N_1945,N_1972);
xor U1983 (N_1983,N_1965,N_1973);
and U1984 (N_1984,N_1958,N_1951);
xnor U1985 (N_1985,N_1924,N_1969);
nand U1986 (N_1986,N_1956,N_1940);
and U1987 (N_1987,N_1921,N_1937);
and U1988 (N_1988,N_1960,N_1935);
nand U1989 (N_1989,N_1941,N_1950);
or U1990 (N_1990,N_1959,N_1963);
xor U1991 (N_1991,N_1967,N_1923);
or U1992 (N_1992,N_1952,N_1954);
or U1993 (N_1993,N_1949,N_1979);
and U1994 (N_1994,N_1975,N_1957);
nor U1995 (N_1995,N_1938,N_1961);
or U1996 (N_1996,N_1927,N_1974);
and U1997 (N_1997,N_1942,N_1925);
nand U1998 (N_1998,N_1932,N_1978);
or U1999 (N_1999,N_1970,N_1920);
or U2000 (N_2000,N_1922,N_1944);
nor U2001 (N_2001,N_1962,N_1936);
xnor U2002 (N_2002,N_1933,N_1953);
nor U2003 (N_2003,N_1964,N_1926);
and U2004 (N_2004,N_1943,N_1966);
and U2005 (N_2005,N_1976,N_1947);
nand U2006 (N_2006,N_1928,N_1971);
nor U2007 (N_2007,N_1931,N_1946);
xnor U2008 (N_2008,N_1968,N_1934);
nand U2009 (N_2009,N_1929,N_1955);
or U2010 (N_2010,N_1956,N_1974);
and U2011 (N_2011,N_1972,N_1931);
or U2012 (N_2012,N_1929,N_1953);
nor U2013 (N_2013,N_1929,N_1960);
and U2014 (N_2014,N_1961,N_1963);
or U2015 (N_2015,N_1961,N_1954);
nor U2016 (N_2016,N_1934,N_1958);
and U2017 (N_2017,N_1952,N_1921);
nor U2018 (N_2018,N_1963,N_1958);
nor U2019 (N_2019,N_1926,N_1962);
nand U2020 (N_2020,N_1948,N_1936);
and U2021 (N_2021,N_1963,N_1976);
xor U2022 (N_2022,N_1978,N_1938);
xor U2023 (N_2023,N_1944,N_1942);
nor U2024 (N_2024,N_1935,N_1940);
and U2025 (N_2025,N_1941,N_1943);
nor U2026 (N_2026,N_1963,N_1939);
and U2027 (N_2027,N_1932,N_1977);
xor U2028 (N_2028,N_1924,N_1927);
nor U2029 (N_2029,N_1941,N_1934);
or U2030 (N_2030,N_1951,N_1971);
nand U2031 (N_2031,N_1936,N_1928);
nand U2032 (N_2032,N_1945,N_1926);
nand U2033 (N_2033,N_1923,N_1927);
nor U2034 (N_2034,N_1975,N_1926);
xor U2035 (N_2035,N_1967,N_1961);
nor U2036 (N_2036,N_1928,N_1958);
and U2037 (N_2037,N_1962,N_1940);
or U2038 (N_2038,N_1937,N_1938);
nor U2039 (N_2039,N_1978,N_1951);
nor U2040 (N_2040,N_2037,N_1983);
nor U2041 (N_2041,N_1987,N_1993);
and U2042 (N_2042,N_1994,N_1999);
and U2043 (N_2043,N_1981,N_2018);
nand U2044 (N_2044,N_2014,N_2031);
nor U2045 (N_2045,N_2001,N_1988);
or U2046 (N_2046,N_1995,N_2028);
nand U2047 (N_2047,N_2006,N_1989);
nand U2048 (N_2048,N_2011,N_2005);
xor U2049 (N_2049,N_2016,N_2009);
and U2050 (N_2050,N_2034,N_1997);
or U2051 (N_2051,N_2004,N_1984);
nand U2052 (N_2052,N_2007,N_2002);
and U2053 (N_2053,N_2013,N_2000);
and U2054 (N_2054,N_2008,N_2015);
and U2055 (N_2055,N_2021,N_2024);
or U2056 (N_2056,N_2017,N_2039);
and U2057 (N_2057,N_2012,N_2026);
xor U2058 (N_2058,N_2010,N_1991);
nor U2059 (N_2059,N_1990,N_2036);
nand U2060 (N_2060,N_1986,N_2003);
or U2061 (N_2061,N_1992,N_2023);
nand U2062 (N_2062,N_2038,N_1998);
nand U2063 (N_2063,N_2019,N_1996);
and U2064 (N_2064,N_1980,N_1982);
and U2065 (N_2065,N_2020,N_2030);
xnor U2066 (N_2066,N_1985,N_2029);
or U2067 (N_2067,N_2035,N_2025);
or U2068 (N_2068,N_2027,N_2022);
nand U2069 (N_2069,N_2032,N_2033);
and U2070 (N_2070,N_1986,N_1998);
nor U2071 (N_2071,N_1992,N_1982);
xor U2072 (N_2072,N_1991,N_2029);
or U2073 (N_2073,N_2024,N_2006);
nor U2074 (N_2074,N_1989,N_1987);
nor U2075 (N_2075,N_2023,N_2017);
xnor U2076 (N_2076,N_1991,N_2027);
xnor U2077 (N_2077,N_1996,N_2021);
xor U2078 (N_2078,N_2000,N_2017);
and U2079 (N_2079,N_2014,N_1996);
xor U2080 (N_2080,N_2030,N_2010);
nand U2081 (N_2081,N_2022,N_1990);
or U2082 (N_2082,N_1985,N_2028);
or U2083 (N_2083,N_1990,N_2008);
nand U2084 (N_2084,N_1991,N_2016);
and U2085 (N_2085,N_2031,N_2026);
nand U2086 (N_2086,N_2037,N_1980);
xnor U2087 (N_2087,N_1983,N_2010);
nand U2088 (N_2088,N_2015,N_2014);
or U2089 (N_2089,N_1981,N_2032);
xor U2090 (N_2090,N_1980,N_2008);
nand U2091 (N_2091,N_1996,N_2029);
or U2092 (N_2092,N_2039,N_1982);
nand U2093 (N_2093,N_2006,N_1983);
nand U2094 (N_2094,N_1998,N_1996);
nand U2095 (N_2095,N_2025,N_2015);
nor U2096 (N_2096,N_1980,N_1997);
xnor U2097 (N_2097,N_2007,N_2038);
and U2098 (N_2098,N_2039,N_2004);
or U2099 (N_2099,N_1986,N_1992);
and U2100 (N_2100,N_2046,N_2041);
nor U2101 (N_2101,N_2075,N_2040);
nand U2102 (N_2102,N_2080,N_2089);
xnor U2103 (N_2103,N_2073,N_2091);
nor U2104 (N_2104,N_2074,N_2081);
and U2105 (N_2105,N_2054,N_2063);
xor U2106 (N_2106,N_2070,N_2042);
and U2107 (N_2107,N_2062,N_2085);
or U2108 (N_2108,N_2076,N_2088);
xnor U2109 (N_2109,N_2078,N_2060);
or U2110 (N_2110,N_2096,N_2045);
nand U2111 (N_2111,N_2084,N_2068);
or U2112 (N_2112,N_2067,N_2053);
and U2113 (N_2113,N_2065,N_2095);
or U2114 (N_2114,N_2079,N_2047);
nand U2115 (N_2115,N_2083,N_2052);
nor U2116 (N_2116,N_2071,N_2061);
or U2117 (N_2117,N_2048,N_2094);
nor U2118 (N_2118,N_2099,N_2082);
or U2119 (N_2119,N_2044,N_2072);
nor U2120 (N_2120,N_2050,N_2049);
or U2121 (N_2121,N_2086,N_2066);
or U2122 (N_2122,N_2098,N_2064);
and U2123 (N_2123,N_2093,N_2043);
nand U2124 (N_2124,N_2051,N_2097);
xnor U2125 (N_2125,N_2058,N_2087);
or U2126 (N_2126,N_2055,N_2057);
and U2127 (N_2127,N_2090,N_2069);
nand U2128 (N_2128,N_2077,N_2056);
and U2129 (N_2129,N_2092,N_2059);
nor U2130 (N_2130,N_2082,N_2072);
nand U2131 (N_2131,N_2049,N_2080);
and U2132 (N_2132,N_2058,N_2069);
xor U2133 (N_2133,N_2093,N_2086);
nor U2134 (N_2134,N_2081,N_2065);
or U2135 (N_2135,N_2051,N_2083);
xnor U2136 (N_2136,N_2088,N_2074);
or U2137 (N_2137,N_2089,N_2097);
nand U2138 (N_2138,N_2082,N_2069);
or U2139 (N_2139,N_2070,N_2049);
xnor U2140 (N_2140,N_2080,N_2052);
xor U2141 (N_2141,N_2055,N_2069);
or U2142 (N_2142,N_2098,N_2046);
nand U2143 (N_2143,N_2070,N_2067);
nand U2144 (N_2144,N_2064,N_2054);
xor U2145 (N_2145,N_2097,N_2050);
and U2146 (N_2146,N_2056,N_2091);
or U2147 (N_2147,N_2087,N_2077);
nand U2148 (N_2148,N_2057,N_2067);
and U2149 (N_2149,N_2052,N_2088);
and U2150 (N_2150,N_2075,N_2049);
or U2151 (N_2151,N_2092,N_2049);
nand U2152 (N_2152,N_2085,N_2042);
or U2153 (N_2153,N_2045,N_2086);
xor U2154 (N_2154,N_2060,N_2075);
or U2155 (N_2155,N_2041,N_2072);
nand U2156 (N_2156,N_2087,N_2051);
xor U2157 (N_2157,N_2060,N_2042);
nand U2158 (N_2158,N_2098,N_2085);
xor U2159 (N_2159,N_2097,N_2049);
and U2160 (N_2160,N_2112,N_2159);
nand U2161 (N_2161,N_2119,N_2149);
xnor U2162 (N_2162,N_2148,N_2110);
and U2163 (N_2163,N_2121,N_2145);
nand U2164 (N_2164,N_2105,N_2158);
or U2165 (N_2165,N_2133,N_2152);
xor U2166 (N_2166,N_2153,N_2106);
nand U2167 (N_2167,N_2132,N_2129);
nor U2168 (N_2168,N_2130,N_2115);
or U2169 (N_2169,N_2151,N_2107);
xnor U2170 (N_2170,N_2142,N_2116);
and U2171 (N_2171,N_2118,N_2103);
nor U2172 (N_2172,N_2143,N_2155);
or U2173 (N_2173,N_2135,N_2147);
nand U2174 (N_2174,N_2104,N_2127);
or U2175 (N_2175,N_2100,N_2124);
nand U2176 (N_2176,N_2111,N_2150);
nand U2177 (N_2177,N_2154,N_2136);
and U2178 (N_2178,N_2125,N_2139);
xnor U2179 (N_2179,N_2102,N_2128);
or U2180 (N_2180,N_2126,N_2109);
xor U2181 (N_2181,N_2137,N_2114);
nand U2182 (N_2182,N_2108,N_2146);
or U2183 (N_2183,N_2141,N_2138);
nand U2184 (N_2184,N_2122,N_2156);
nand U2185 (N_2185,N_2117,N_2101);
nand U2186 (N_2186,N_2120,N_2144);
nand U2187 (N_2187,N_2131,N_2123);
xnor U2188 (N_2188,N_2157,N_2134);
nand U2189 (N_2189,N_2140,N_2113);
nand U2190 (N_2190,N_2132,N_2116);
or U2191 (N_2191,N_2105,N_2100);
nand U2192 (N_2192,N_2103,N_2158);
nand U2193 (N_2193,N_2139,N_2112);
or U2194 (N_2194,N_2121,N_2147);
and U2195 (N_2195,N_2110,N_2134);
xor U2196 (N_2196,N_2140,N_2131);
or U2197 (N_2197,N_2132,N_2110);
or U2198 (N_2198,N_2110,N_2119);
xnor U2199 (N_2199,N_2141,N_2101);
xnor U2200 (N_2200,N_2150,N_2154);
and U2201 (N_2201,N_2132,N_2158);
or U2202 (N_2202,N_2149,N_2155);
xor U2203 (N_2203,N_2146,N_2154);
nor U2204 (N_2204,N_2158,N_2102);
or U2205 (N_2205,N_2146,N_2156);
or U2206 (N_2206,N_2159,N_2124);
xor U2207 (N_2207,N_2147,N_2120);
and U2208 (N_2208,N_2115,N_2112);
xor U2209 (N_2209,N_2137,N_2100);
and U2210 (N_2210,N_2120,N_2122);
nor U2211 (N_2211,N_2147,N_2125);
and U2212 (N_2212,N_2129,N_2121);
and U2213 (N_2213,N_2147,N_2126);
xnor U2214 (N_2214,N_2138,N_2116);
xor U2215 (N_2215,N_2108,N_2157);
and U2216 (N_2216,N_2131,N_2135);
nand U2217 (N_2217,N_2107,N_2114);
nand U2218 (N_2218,N_2127,N_2158);
nand U2219 (N_2219,N_2132,N_2131);
and U2220 (N_2220,N_2173,N_2172);
and U2221 (N_2221,N_2176,N_2186);
nor U2222 (N_2222,N_2165,N_2175);
nor U2223 (N_2223,N_2218,N_2182);
xor U2224 (N_2224,N_2177,N_2181);
nor U2225 (N_2225,N_2211,N_2203);
and U2226 (N_2226,N_2194,N_2187);
nand U2227 (N_2227,N_2202,N_2196);
nor U2228 (N_2228,N_2189,N_2208);
or U2229 (N_2229,N_2167,N_2213);
xnor U2230 (N_2230,N_2188,N_2178);
xnor U2231 (N_2231,N_2180,N_2219);
xor U2232 (N_2232,N_2174,N_2169);
and U2233 (N_2233,N_2201,N_2197);
or U2234 (N_2234,N_2210,N_2191);
or U2235 (N_2235,N_2184,N_2214);
and U2236 (N_2236,N_2198,N_2160);
xor U2237 (N_2237,N_2163,N_2192);
or U2238 (N_2238,N_2168,N_2216);
nor U2239 (N_2239,N_2166,N_2170);
and U2240 (N_2240,N_2190,N_2204);
nand U2241 (N_2241,N_2215,N_2206);
nand U2242 (N_2242,N_2207,N_2162);
xnor U2243 (N_2243,N_2199,N_2193);
xnor U2244 (N_2244,N_2209,N_2212);
nor U2245 (N_2245,N_2205,N_2171);
xnor U2246 (N_2246,N_2195,N_2179);
nand U2247 (N_2247,N_2161,N_2183);
or U2248 (N_2248,N_2185,N_2200);
or U2249 (N_2249,N_2164,N_2217);
and U2250 (N_2250,N_2186,N_2188);
and U2251 (N_2251,N_2160,N_2197);
and U2252 (N_2252,N_2183,N_2199);
and U2253 (N_2253,N_2174,N_2191);
and U2254 (N_2254,N_2197,N_2206);
nor U2255 (N_2255,N_2204,N_2164);
and U2256 (N_2256,N_2199,N_2198);
xnor U2257 (N_2257,N_2213,N_2168);
or U2258 (N_2258,N_2196,N_2173);
xor U2259 (N_2259,N_2204,N_2216);
nand U2260 (N_2260,N_2215,N_2186);
nor U2261 (N_2261,N_2214,N_2182);
and U2262 (N_2262,N_2176,N_2170);
or U2263 (N_2263,N_2212,N_2201);
nand U2264 (N_2264,N_2181,N_2213);
nand U2265 (N_2265,N_2188,N_2196);
nor U2266 (N_2266,N_2215,N_2209);
or U2267 (N_2267,N_2201,N_2189);
nor U2268 (N_2268,N_2193,N_2211);
xnor U2269 (N_2269,N_2188,N_2202);
or U2270 (N_2270,N_2192,N_2217);
or U2271 (N_2271,N_2185,N_2182);
and U2272 (N_2272,N_2213,N_2191);
and U2273 (N_2273,N_2180,N_2202);
or U2274 (N_2274,N_2190,N_2206);
or U2275 (N_2275,N_2211,N_2186);
nand U2276 (N_2276,N_2191,N_2181);
nor U2277 (N_2277,N_2175,N_2196);
or U2278 (N_2278,N_2179,N_2199);
and U2279 (N_2279,N_2198,N_2176);
nand U2280 (N_2280,N_2236,N_2225);
nor U2281 (N_2281,N_2229,N_2254);
xnor U2282 (N_2282,N_2248,N_2265);
and U2283 (N_2283,N_2232,N_2223);
nand U2284 (N_2284,N_2252,N_2228);
and U2285 (N_2285,N_2230,N_2250);
xor U2286 (N_2286,N_2243,N_2257);
or U2287 (N_2287,N_2255,N_2260);
or U2288 (N_2288,N_2259,N_2221);
nor U2289 (N_2289,N_2244,N_2267);
or U2290 (N_2290,N_2234,N_2273);
and U2291 (N_2291,N_2277,N_2274);
and U2292 (N_2292,N_2275,N_2269);
or U2293 (N_2293,N_2235,N_2246);
and U2294 (N_2294,N_2237,N_2271);
nand U2295 (N_2295,N_2231,N_2222);
nor U2296 (N_2296,N_2233,N_2245);
xor U2297 (N_2297,N_2226,N_2239);
nor U2298 (N_2298,N_2278,N_2270);
and U2299 (N_2299,N_2258,N_2276);
nand U2300 (N_2300,N_2227,N_2240);
or U2301 (N_2301,N_2251,N_2238);
xor U2302 (N_2302,N_2262,N_2264);
nor U2303 (N_2303,N_2256,N_2253);
xnor U2304 (N_2304,N_2279,N_2224);
xor U2305 (N_2305,N_2268,N_2247);
xor U2306 (N_2306,N_2242,N_2241);
xnor U2307 (N_2307,N_2220,N_2261);
or U2308 (N_2308,N_2272,N_2266);
xor U2309 (N_2309,N_2249,N_2263);
or U2310 (N_2310,N_2250,N_2274);
nand U2311 (N_2311,N_2279,N_2245);
or U2312 (N_2312,N_2227,N_2232);
nand U2313 (N_2313,N_2237,N_2262);
and U2314 (N_2314,N_2279,N_2278);
nand U2315 (N_2315,N_2227,N_2245);
nor U2316 (N_2316,N_2230,N_2247);
nand U2317 (N_2317,N_2234,N_2251);
xor U2318 (N_2318,N_2255,N_2265);
xnor U2319 (N_2319,N_2276,N_2256);
and U2320 (N_2320,N_2263,N_2221);
nand U2321 (N_2321,N_2244,N_2235);
and U2322 (N_2322,N_2229,N_2267);
xnor U2323 (N_2323,N_2272,N_2257);
and U2324 (N_2324,N_2251,N_2241);
and U2325 (N_2325,N_2242,N_2262);
or U2326 (N_2326,N_2224,N_2265);
xnor U2327 (N_2327,N_2251,N_2233);
xnor U2328 (N_2328,N_2223,N_2249);
nor U2329 (N_2329,N_2223,N_2237);
or U2330 (N_2330,N_2230,N_2254);
or U2331 (N_2331,N_2237,N_2249);
nand U2332 (N_2332,N_2243,N_2263);
nand U2333 (N_2333,N_2244,N_2230);
and U2334 (N_2334,N_2263,N_2259);
nand U2335 (N_2335,N_2273,N_2257);
xor U2336 (N_2336,N_2250,N_2271);
xnor U2337 (N_2337,N_2269,N_2270);
xnor U2338 (N_2338,N_2231,N_2225);
or U2339 (N_2339,N_2274,N_2262);
nor U2340 (N_2340,N_2281,N_2317);
nor U2341 (N_2341,N_2287,N_2313);
nor U2342 (N_2342,N_2293,N_2304);
xnor U2343 (N_2343,N_2300,N_2305);
nand U2344 (N_2344,N_2329,N_2292);
or U2345 (N_2345,N_2327,N_2315);
nand U2346 (N_2346,N_2320,N_2309);
and U2347 (N_2347,N_2323,N_2310);
or U2348 (N_2348,N_2330,N_2326);
and U2349 (N_2349,N_2299,N_2335);
nor U2350 (N_2350,N_2302,N_2321);
nand U2351 (N_2351,N_2322,N_2290);
nand U2352 (N_2352,N_2297,N_2339);
nor U2353 (N_2353,N_2284,N_2286);
xnor U2354 (N_2354,N_2285,N_2314);
or U2355 (N_2355,N_2318,N_2303);
and U2356 (N_2356,N_2331,N_2338);
nor U2357 (N_2357,N_2301,N_2280);
or U2358 (N_2358,N_2294,N_2283);
nor U2359 (N_2359,N_2316,N_2336);
and U2360 (N_2360,N_2311,N_2334);
xnor U2361 (N_2361,N_2337,N_2333);
xnor U2362 (N_2362,N_2298,N_2324);
nand U2363 (N_2363,N_2288,N_2307);
nor U2364 (N_2364,N_2328,N_2308);
xnor U2365 (N_2365,N_2295,N_2319);
xor U2366 (N_2366,N_2296,N_2282);
nor U2367 (N_2367,N_2289,N_2332);
nor U2368 (N_2368,N_2291,N_2306);
nand U2369 (N_2369,N_2325,N_2312);
or U2370 (N_2370,N_2332,N_2288);
xor U2371 (N_2371,N_2325,N_2329);
nand U2372 (N_2372,N_2318,N_2295);
xnor U2373 (N_2373,N_2289,N_2321);
and U2374 (N_2374,N_2285,N_2323);
or U2375 (N_2375,N_2286,N_2305);
and U2376 (N_2376,N_2298,N_2323);
or U2377 (N_2377,N_2301,N_2311);
and U2378 (N_2378,N_2285,N_2326);
xnor U2379 (N_2379,N_2288,N_2328);
nand U2380 (N_2380,N_2294,N_2286);
xor U2381 (N_2381,N_2298,N_2293);
xnor U2382 (N_2382,N_2310,N_2309);
or U2383 (N_2383,N_2292,N_2325);
or U2384 (N_2384,N_2318,N_2323);
nor U2385 (N_2385,N_2300,N_2330);
nand U2386 (N_2386,N_2286,N_2316);
xor U2387 (N_2387,N_2308,N_2327);
xnor U2388 (N_2388,N_2284,N_2309);
or U2389 (N_2389,N_2333,N_2287);
xor U2390 (N_2390,N_2309,N_2317);
xor U2391 (N_2391,N_2291,N_2339);
xor U2392 (N_2392,N_2286,N_2314);
xnor U2393 (N_2393,N_2314,N_2302);
nand U2394 (N_2394,N_2292,N_2326);
or U2395 (N_2395,N_2313,N_2321);
nand U2396 (N_2396,N_2339,N_2329);
and U2397 (N_2397,N_2326,N_2291);
xor U2398 (N_2398,N_2285,N_2336);
or U2399 (N_2399,N_2302,N_2329);
nor U2400 (N_2400,N_2360,N_2370);
nand U2401 (N_2401,N_2342,N_2393);
xor U2402 (N_2402,N_2389,N_2386);
and U2403 (N_2403,N_2384,N_2345);
and U2404 (N_2404,N_2387,N_2383);
nor U2405 (N_2405,N_2361,N_2375);
nand U2406 (N_2406,N_2371,N_2349);
or U2407 (N_2407,N_2344,N_2346);
xnor U2408 (N_2408,N_2390,N_2395);
and U2409 (N_2409,N_2362,N_2354);
xor U2410 (N_2410,N_2380,N_2357);
nand U2411 (N_2411,N_2379,N_2373);
nor U2412 (N_2412,N_2396,N_2356);
or U2413 (N_2413,N_2381,N_2385);
or U2414 (N_2414,N_2369,N_2394);
nor U2415 (N_2415,N_2378,N_2351);
xnor U2416 (N_2416,N_2358,N_2348);
xor U2417 (N_2417,N_2377,N_2363);
and U2418 (N_2418,N_2398,N_2341);
and U2419 (N_2419,N_2367,N_2352);
nor U2420 (N_2420,N_2399,N_2392);
nand U2421 (N_2421,N_2368,N_2347);
nand U2422 (N_2422,N_2365,N_2397);
nand U2423 (N_2423,N_2350,N_2391);
nor U2424 (N_2424,N_2388,N_2374);
nor U2425 (N_2425,N_2372,N_2359);
nand U2426 (N_2426,N_2343,N_2382);
or U2427 (N_2427,N_2366,N_2364);
nand U2428 (N_2428,N_2340,N_2355);
and U2429 (N_2429,N_2376,N_2353);
and U2430 (N_2430,N_2394,N_2361);
and U2431 (N_2431,N_2392,N_2372);
and U2432 (N_2432,N_2345,N_2399);
or U2433 (N_2433,N_2351,N_2399);
or U2434 (N_2434,N_2349,N_2391);
and U2435 (N_2435,N_2398,N_2392);
nor U2436 (N_2436,N_2379,N_2370);
xnor U2437 (N_2437,N_2359,N_2365);
or U2438 (N_2438,N_2373,N_2382);
xor U2439 (N_2439,N_2352,N_2394);
nand U2440 (N_2440,N_2361,N_2341);
nand U2441 (N_2441,N_2384,N_2389);
or U2442 (N_2442,N_2396,N_2381);
xor U2443 (N_2443,N_2368,N_2392);
or U2444 (N_2444,N_2352,N_2391);
nand U2445 (N_2445,N_2393,N_2397);
nor U2446 (N_2446,N_2379,N_2363);
or U2447 (N_2447,N_2370,N_2392);
xor U2448 (N_2448,N_2355,N_2398);
and U2449 (N_2449,N_2353,N_2391);
nand U2450 (N_2450,N_2347,N_2369);
xnor U2451 (N_2451,N_2387,N_2384);
nand U2452 (N_2452,N_2345,N_2351);
and U2453 (N_2453,N_2356,N_2397);
or U2454 (N_2454,N_2375,N_2370);
nor U2455 (N_2455,N_2359,N_2345);
nor U2456 (N_2456,N_2349,N_2358);
and U2457 (N_2457,N_2356,N_2361);
or U2458 (N_2458,N_2359,N_2383);
nand U2459 (N_2459,N_2355,N_2360);
and U2460 (N_2460,N_2410,N_2425);
and U2461 (N_2461,N_2432,N_2400);
nor U2462 (N_2462,N_2429,N_2457);
xor U2463 (N_2463,N_2428,N_2422);
nor U2464 (N_2464,N_2440,N_2442);
xor U2465 (N_2465,N_2446,N_2437);
xnor U2466 (N_2466,N_2443,N_2419);
or U2467 (N_2467,N_2412,N_2450);
xnor U2468 (N_2468,N_2416,N_2421);
and U2469 (N_2469,N_2445,N_2407);
nor U2470 (N_2470,N_2431,N_2434);
or U2471 (N_2471,N_2453,N_2411);
xor U2472 (N_2472,N_2424,N_2427);
nor U2473 (N_2473,N_2409,N_2403);
xnor U2474 (N_2474,N_2418,N_2451);
nor U2475 (N_2475,N_2447,N_2402);
nor U2476 (N_2476,N_2406,N_2458);
nor U2477 (N_2477,N_2404,N_2430);
nand U2478 (N_2478,N_2439,N_2454);
xnor U2479 (N_2479,N_2438,N_2449);
or U2480 (N_2480,N_2417,N_2414);
or U2481 (N_2481,N_2459,N_2456);
xor U2482 (N_2482,N_2448,N_2444);
nand U2483 (N_2483,N_2433,N_2415);
nor U2484 (N_2484,N_2408,N_2420);
nand U2485 (N_2485,N_2455,N_2436);
nand U2486 (N_2486,N_2441,N_2401);
or U2487 (N_2487,N_2405,N_2435);
and U2488 (N_2488,N_2452,N_2413);
or U2489 (N_2489,N_2426,N_2423);
or U2490 (N_2490,N_2419,N_2441);
and U2491 (N_2491,N_2427,N_2438);
nand U2492 (N_2492,N_2408,N_2449);
or U2493 (N_2493,N_2455,N_2432);
or U2494 (N_2494,N_2447,N_2413);
nor U2495 (N_2495,N_2402,N_2428);
nand U2496 (N_2496,N_2427,N_2448);
and U2497 (N_2497,N_2414,N_2444);
or U2498 (N_2498,N_2408,N_2416);
or U2499 (N_2499,N_2429,N_2448);
and U2500 (N_2500,N_2450,N_2404);
or U2501 (N_2501,N_2419,N_2424);
xnor U2502 (N_2502,N_2425,N_2458);
nand U2503 (N_2503,N_2415,N_2401);
xnor U2504 (N_2504,N_2412,N_2438);
or U2505 (N_2505,N_2405,N_2408);
nand U2506 (N_2506,N_2423,N_2458);
and U2507 (N_2507,N_2412,N_2439);
xnor U2508 (N_2508,N_2416,N_2403);
and U2509 (N_2509,N_2409,N_2400);
nor U2510 (N_2510,N_2417,N_2456);
and U2511 (N_2511,N_2453,N_2425);
and U2512 (N_2512,N_2419,N_2458);
xnor U2513 (N_2513,N_2444,N_2458);
and U2514 (N_2514,N_2453,N_2406);
or U2515 (N_2515,N_2443,N_2438);
nor U2516 (N_2516,N_2418,N_2403);
nand U2517 (N_2517,N_2418,N_2424);
nor U2518 (N_2518,N_2413,N_2429);
nor U2519 (N_2519,N_2407,N_2406);
nand U2520 (N_2520,N_2489,N_2468);
or U2521 (N_2521,N_2502,N_2462);
nand U2522 (N_2522,N_2478,N_2463);
xor U2523 (N_2523,N_2474,N_2498);
xor U2524 (N_2524,N_2499,N_2479);
and U2525 (N_2525,N_2461,N_2484);
or U2526 (N_2526,N_2492,N_2482);
nand U2527 (N_2527,N_2494,N_2510);
nand U2528 (N_2528,N_2466,N_2505);
or U2529 (N_2529,N_2469,N_2497);
and U2530 (N_2530,N_2515,N_2475);
and U2531 (N_2531,N_2471,N_2517);
and U2532 (N_2532,N_2512,N_2467);
or U2533 (N_2533,N_2501,N_2514);
or U2534 (N_2534,N_2493,N_2496);
or U2535 (N_2535,N_2511,N_2506);
nor U2536 (N_2536,N_2488,N_2465);
nor U2537 (N_2537,N_2508,N_2477);
and U2538 (N_2538,N_2507,N_2481);
and U2539 (N_2539,N_2460,N_2500);
nand U2540 (N_2540,N_2480,N_2486);
or U2541 (N_2541,N_2518,N_2464);
nor U2542 (N_2542,N_2504,N_2491);
and U2543 (N_2543,N_2472,N_2519);
nand U2544 (N_2544,N_2490,N_2483);
nor U2545 (N_2545,N_2509,N_2476);
xor U2546 (N_2546,N_2473,N_2513);
nor U2547 (N_2547,N_2495,N_2470);
nor U2548 (N_2548,N_2485,N_2487);
or U2549 (N_2549,N_2503,N_2516);
or U2550 (N_2550,N_2489,N_2509);
nor U2551 (N_2551,N_2489,N_2463);
nor U2552 (N_2552,N_2503,N_2504);
and U2553 (N_2553,N_2483,N_2460);
nand U2554 (N_2554,N_2490,N_2513);
nand U2555 (N_2555,N_2477,N_2463);
xor U2556 (N_2556,N_2509,N_2511);
xor U2557 (N_2557,N_2460,N_2510);
nor U2558 (N_2558,N_2513,N_2510);
and U2559 (N_2559,N_2467,N_2485);
and U2560 (N_2560,N_2474,N_2483);
xnor U2561 (N_2561,N_2508,N_2518);
and U2562 (N_2562,N_2503,N_2467);
nand U2563 (N_2563,N_2504,N_2487);
nand U2564 (N_2564,N_2497,N_2477);
xnor U2565 (N_2565,N_2506,N_2485);
nand U2566 (N_2566,N_2483,N_2487);
nor U2567 (N_2567,N_2502,N_2478);
nor U2568 (N_2568,N_2514,N_2509);
nor U2569 (N_2569,N_2496,N_2460);
or U2570 (N_2570,N_2475,N_2462);
and U2571 (N_2571,N_2461,N_2462);
and U2572 (N_2572,N_2468,N_2484);
nand U2573 (N_2573,N_2502,N_2517);
nand U2574 (N_2574,N_2484,N_2518);
nor U2575 (N_2575,N_2502,N_2503);
or U2576 (N_2576,N_2517,N_2494);
xnor U2577 (N_2577,N_2470,N_2491);
xor U2578 (N_2578,N_2491,N_2519);
or U2579 (N_2579,N_2504,N_2516);
nand U2580 (N_2580,N_2557,N_2540);
or U2581 (N_2581,N_2579,N_2560);
or U2582 (N_2582,N_2546,N_2524);
xor U2583 (N_2583,N_2539,N_2561);
xnor U2584 (N_2584,N_2542,N_2553);
and U2585 (N_2585,N_2572,N_2554);
xor U2586 (N_2586,N_2567,N_2522);
nand U2587 (N_2587,N_2574,N_2547);
xnor U2588 (N_2588,N_2575,N_2569);
nor U2589 (N_2589,N_2571,N_2576);
or U2590 (N_2590,N_2573,N_2535);
and U2591 (N_2591,N_2544,N_2564);
nand U2592 (N_2592,N_2577,N_2552);
or U2593 (N_2593,N_2558,N_2531);
or U2594 (N_2594,N_2570,N_2551);
and U2595 (N_2595,N_2566,N_2556);
nand U2596 (N_2596,N_2549,N_2559);
or U2597 (N_2597,N_2562,N_2550);
nor U2598 (N_2598,N_2538,N_2529);
and U2599 (N_2599,N_2543,N_2523);
or U2600 (N_2600,N_2530,N_2533);
nor U2601 (N_2601,N_2565,N_2520);
nor U2602 (N_2602,N_2537,N_2528);
xor U2603 (N_2603,N_2548,N_2521);
nand U2604 (N_2604,N_2532,N_2527);
and U2605 (N_2605,N_2534,N_2563);
nand U2606 (N_2606,N_2541,N_2545);
or U2607 (N_2607,N_2536,N_2525);
nand U2608 (N_2608,N_2526,N_2568);
nand U2609 (N_2609,N_2578,N_2555);
nor U2610 (N_2610,N_2571,N_2545);
or U2611 (N_2611,N_2531,N_2560);
nor U2612 (N_2612,N_2559,N_2523);
xnor U2613 (N_2613,N_2551,N_2556);
nand U2614 (N_2614,N_2556,N_2549);
xor U2615 (N_2615,N_2554,N_2568);
and U2616 (N_2616,N_2552,N_2562);
nand U2617 (N_2617,N_2530,N_2558);
and U2618 (N_2618,N_2526,N_2528);
or U2619 (N_2619,N_2561,N_2534);
nor U2620 (N_2620,N_2574,N_2572);
nor U2621 (N_2621,N_2537,N_2551);
or U2622 (N_2622,N_2542,N_2563);
and U2623 (N_2623,N_2536,N_2520);
xnor U2624 (N_2624,N_2553,N_2541);
nor U2625 (N_2625,N_2524,N_2531);
nor U2626 (N_2626,N_2571,N_2573);
nor U2627 (N_2627,N_2566,N_2550);
nand U2628 (N_2628,N_2562,N_2557);
xnor U2629 (N_2629,N_2530,N_2565);
nand U2630 (N_2630,N_2525,N_2539);
nand U2631 (N_2631,N_2553,N_2565);
and U2632 (N_2632,N_2548,N_2574);
nor U2633 (N_2633,N_2566,N_2520);
and U2634 (N_2634,N_2564,N_2548);
and U2635 (N_2635,N_2525,N_2559);
nor U2636 (N_2636,N_2571,N_2540);
nor U2637 (N_2637,N_2533,N_2575);
nand U2638 (N_2638,N_2571,N_2541);
xnor U2639 (N_2639,N_2520,N_2546);
xor U2640 (N_2640,N_2636,N_2631);
nand U2641 (N_2641,N_2614,N_2592);
xor U2642 (N_2642,N_2616,N_2625);
nand U2643 (N_2643,N_2582,N_2591);
or U2644 (N_2644,N_2624,N_2620);
or U2645 (N_2645,N_2623,N_2603);
or U2646 (N_2646,N_2617,N_2605);
xnor U2647 (N_2647,N_2587,N_2607);
or U2648 (N_2648,N_2597,N_2633);
nor U2649 (N_2649,N_2581,N_2598);
and U2650 (N_2650,N_2601,N_2622);
xor U2651 (N_2651,N_2637,N_2621);
and U2652 (N_2652,N_2612,N_2585);
nor U2653 (N_2653,N_2615,N_2609);
and U2654 (N_2654,N_2628,N_2596);
xnor U2655 (N_2655,N_2638,N_2639);
or U2656 (N_2656,N_2600,N_2593);
nor U2657 (N_2657,N_2586,N_2613);
nor U2658 (N_2658,N_2626,N_2630);
and U2659 (N_2659,N_2602,N_2618);
nand U2660 (N_2660,N_2611,N_2584);
nor U2661 (N_2661,N_2580,N_2632);
nand U2662 (N_2662,N_2606,N_2604);
and U2663 (N_2663,N_2599,N_2588);
nand U2664 (N_2664,N_2629,N_2619);
nor U2665 (N_2665,N_2590,N_2589);
xnor U2666 (N_2666,N_2595,N_2583);
nor U2667 (N_2667,N_2610,N_2634);
or U2668 (N_2668,N_2627,N_2608);
xnor U2669 (N_2669,N_2635,N_2594);
xnor U2670 (N_2670,N_2582,N_2627);
xor U2671 (N_2671,N_2595,N_2639);
nand U2672 (N_2672,N_2615,N_2607);
nor U2673 (N_2673,N_2639,N_2617);
xor U2674 (N_2674,N_2618,N_2591);
and U2675 (N_2675,N_2592,N_2608);
and U2676 (N_2676,N_2628,N_2638);
nor U2677 (N_2677,N_2615,N_2608);
nor U2678 (N_2678,N_2632,N_2622);
xor U2679 (N_2679,N_2588,N_2636);
and U2680 (N_2680,N_2596,N_2597);
nor U2681 (N_2681,N_2604,N_2585);
nand U2682 (N_2682,N_2588,N_2602);
or U2683 (N_2683,N_2622,N_2594);
and U2684 (N_2684,N_2595,N_2608);
xor U2685 (N_2685,N_2622,N_2627);
xnor U2686 (N_2686,N_2605,N_2602);
and U2687 (N_2687,N_2621,N_2627);
or U2688 (N_2688,N_2607,N_2612);
and U2689 (N_2689,N_2629,N_2610);
nor U2690 (N_2690,N_2582,N_2602);
nand U2691 (N_2691,N_2609,N_2623);
xor U2692 (N_2692,N_2600,N_2625);
xnor U2693 (N_2693,N_2595,N_2589);
and U2694 (N_2694,N_2621,N_2617);
nand U2695 (N_2695,N_2590,N_2609);
or U2696 (N_2696,N_2604,N_2607);
nand U2697 (N_2697,N_2594,N_2600);
or U2698 (N_2698,N_2601,N_2603);
or U2699 (N_2699,N_2602,N_2587);
or U2700 (N_2700,N_2659,N_2690);
or U2701 (N_2701,N_2640,N_2646);
nor U2702 (N_2702,N_2681,N_2699);
nand U2703 (N_2703,N_2647,N_2674);
xnor U2704 (N_2704,N_2662,N_2687);
xor U2705 (N_2705,N_2650,N_2658);
xor U2706 (N_2706,N_2693,N_2692);
xnor U2707 (N_2707,N_2654,N_2657);
and U2708 (N_2708,N_2648,N_2664);
nor U2709 (N_2709,N_2697,N_2684);
or U2710 (N_2710,N_2691,N_2644);
and U2711 (N_2711,N_2677,N_2645);
nor U2712 (N_2712,N_2670,N_2696);
or U2713 (N_2713,N_2686,N_2665);
xor U2714 (N_2714,N_2655,N_2652);
or U2715 (N_2715,N_2685,N_2643);
and U2716 (N_2716,N_2668,N_2656);
xnor U2717 (N_2717,N_2688,N_2653);
nand U2718 (N_2718,N_2663,N_2679);
nor U2719 (N_2719,N_2678,N_2641);
and U2720 (N_2720,N_2671,N_2667);
nand U2721 (N_2721,N_2661,N_2669);
and U2722 (N_2722,N_2660,N_2666);
nand U2723 (N_2723,N_2683,N_2680);
and U2724 (N_2724,N_2642,N_2694);
nand U2725 (N_2725,N_2651,N_2675);
nor U2726 (N_2726,N_2672,N_2695);
and U2727 (N_2727,N_2676,N_2682);
and U2728 (N_2728,N_2673,N_2689);
nand U2729 (N_2729,N_2649,N_2698);
nor U2730 (N_2730,N_2646,N_2654);
or U2731 (N_2731,N_2641,N_2642);
and U2732 (N_2732,N_2699,N_2690);
nand U2733 (N_2733,N_2679,N_2681);
or U2734 (N_2734,N_2685,N_2691);
xnor U2735 (N_2735,N_2647,N_2656);
or U2736 (N_2736,N_2661,N_2689);
nor U2737 (N_2737,N_2646,N_2671);
nand U2738 (N_2738,N_2673,N_2690);
nand U2739 (N_2739,N_2649,N_2668);
xnor U2740 (N_2740,N_2667,N_2656);
nand U2741 (N_2741,N_2645,N_2676);
and U2742 (N_2742,N_2656,N_2671);
xor U2743 (N_2743,N_2656,N_2681);
xor U2744 (N_2744,N_2692,N_2642);
and U2745 (N_2745,N_2696,N_2665);
nand U2746 (N_2746,N_2650,N_2655);
or U2747 (N_2747,N_2656,N_2696);
xnor U2748 (N_2748,N_2669,N_2663);
or U2749 (N_2749,N_2687,N_2644);
nand U2750 (N_2750,N_2699,N_2684);
nand U2751 (N_2751,N_2654,N_2691);
xnor U2752 (N_2752,N_2696,N_2658);
and U2753 (N_2753,N_2654,N_2648);
nor U2754 (N_2754,N_2649,N_2677);
nor U2755 (N_2755,N_2681,N_2676);
xnor U2756 (N_2756,N_2672,N_2699);
or U2757 (N_2757,N_2660,N_2645);
or U2758 (N_2758,N_2651,N_2693);
nand U2759 (N_2759,N_2685,N_2640);
nand U2760 (N_2760,N_2703,N_2731);
or U2761 (N_2761,N_2721,N_2733);
or U2762 (N_2762,N_2746,N_2700);
and U2763 (N_2763,N_2719,N_2756);
and U2764 (N_2764,N_2704,N_2749);
nand U2765 (N_2765,N_2711,N_2739);
or U2766 (N_2766,N_2715,N_2747);
or U2767 (N_2767,N_2741,N_2743);
or U2768 (N_2768,N_2717,N_2724);
nand U2769 (N_2769,N_2748,N_2742);
and U2770 (N_2770,N_2732,N_2726);
and U2771 (N_2771,N_2754,N_2736);
nand U2772 (N_2772,N_2758,N_2716);
xor U2773 (N_2773,N_2701,N_2707);
or U2774 (N_2774,N_2718,N_2757);
nor U2775 (N_2775,N_2713,N_2750);
and U2776 (N_2776,N_2753,N_2752);
and U2777 (N_2777,N_2729,N_2737);
and U2778 (N_2778,N_2734,N_2710);
and U2779 (N_2779,N_2728,N_2740);
xnor U2780 (N_2780,N_2712,N_2745);
or U2781 (N_2781,N_2708,N_2720);
or U2782 (N_2782,N_2727,N_2709);
nor U2783 (N_2783,N_2735,N_2725);
or U2784 (N_2784,N_2751,N_2722);
or U2785 (N_2785,N_2723,N_2706);
nor U2786 (N_2786,N_2755,N_2705);
and U2787 (N_2787,N_2759,N_2744);
xnor U2788 (N_2788,N_2738,N_2702);
nor U2789 (N_2789,N_2730,N_2714);
or U2790 (N_2790,N_2726,N_2749);
and U2791 (N_2791,N_2742,N_2707);
nor U2792 (N_2792,N_2732,N_2748);
nor U2793 (N_2793,N_2742,N_2713);
xor U2794 (N_2794,N_2740,N_2730);
xor U2795 (N_2795,N_2754,N_2717);
nand U2796 (N_2796,N_2718,N_2744);
or U2797 (N_2797,N_2740,N_2751);
nand U2798 (N_2798,N_2705,N_2726);
xor U2799 (N_2799,N_2721,N_2720);
nor U2800 (N_2800,N_2734,N_2756);
nand U2801 (N_2801,N_2754,N_2733);
nand U2802 (N_2802,N_2755,N_2706);
or U2803 (N_2803,N_2750,N_2753);
xnor U2804 (N_2804,N_2740,N_2723);
and U2805 (N_2805,N_2735,N_2724);
xor U2806 (N_2806,N_2707,N_2717);
nand U2807 (N_2807,N_2756,N_2722);
nor U2808 (N_2808,N_2741,N_2755);
and U2809 (N_2809,N_2718,N_2752);
nand U2810 (N_2810,N_2725,N_2711);
or U2811 (N_2811,N_2757,N_2730);
or U2812 (N_2812,N_2749,N_2717);
or U2813 (N_2813,N_2731,N_2726);
or U2814 (N_2814,N_2722,N_2718);
or U2815 (N_2815,N_2750,N_2717);
nand U2816 (N_2816,N_2729,N_2718);
and U2817 (N_2817,N_2758,N_2747);
or U2818 (N_2818,N_2740,N_2747);
nor U2819 (N_2819,N_2710,N_2737);
nand U2820 (N_2820,N_2781,N_2771);
and U2821 (N_2821,N_2812,N_2792);
or U2822 (N_2822,N_2778,N_2760);
xnor U2823 (N_2823,N_2811,N_2813);
nor U2824 (N_2824,N_2818,N_2805);
nor U2825 (N_2825,N_2769,N_2785);
and U2826 (N_2826,N_2763,N_2795);
xor U2827 (N_2827,N_2782,N_2774);
and U2828 (N_2828,N_2762,N_2793);
nor U2829 (N_2829,N_2804,N_2780);
xor U2830 (N_2830,N_2790,N_2773);
nor U2831 (N_2831,N_2766,N_2794);
nand U2832 (N_2832,N_2789,N_2802);
nor U2833 (N_2833,N_2808,N_2799);
xnor U2834 (N_2834,N_2772,N_2770);
and U2835 (N_2835,N_2779,N_2810);
nand U2836 (N_2836,N_2797,N_2784);
nor U2837 (N_2837,N_2798,N_2800);
and U2838 (N_2838,N_2761,N_2788);
nor U2839 (N_2839,N_2775,N_2814);
or U2840 (N_2840,N_2816,N_2807);
nand U2841 (N_2841,N_2786,N_2767);
xor U2842 (N_2842,N_2817,N_2776);
and U2843 (N_2843,N_2809,N_2765);
or U2844 (N_2844,N_2815,N_2791);
nor U2845 (N_2845,N_2806,N_2783);
xnor U2846 (N_2846,N_2801,N_2768);
xor U2847 (N_2847,N_2777,N_2796);
nand U2848 (N_2848,N_2819,N_2764);
nor U2849 (N_2849,N_2787,N_2803);
nor U2850 (N_2850,N_2809,N_2781);
nand U2851 (N_2851,N_2806,N_2796);
nand U2852 (N_2852,N_2800,N_2781);
or U2853 (N_2853,N_2765,N_2767);
xor U2854 (N_2854,N_2796,N_2785);
nor U2855 (N_2855,N_2789,N_2777);
nor U2856 (N_2856,N_2766,N_2769);
or U2857 (N_2857,N_2811,N_2792);
and U2858 (N_2858,N_2780,N_2805);
and U2859 (N_2859,N_2807,N_2792);
nor U2860 (N_2860,N_2763,N_2768);
or U2861 (N_2861,N_2765,N_2797);
nor U2862 (N_2862,N_2800,N_2809);
nor U2863 (N_2863,N_2776,N_2764);
or U2864 (N_2864,N_2799,N_2777);
and U2865 (N_2865,N_2794,N_2762);
and U2866 (N_2866,N_2802,N_2803);
and U2867 (N_2867,N_2767,N_2781);
and U2868 (N_2868,N_2767,N_2762);
nor U2869 (N_2869,N_2765,N_2772);
and U2870 (N_2870,N_2775,N_2786);
nor U2871 (N_2871,N_2783,N_2781);
and U2872 (N_2872,N_2774,N_2809);
or U2873 (N_2873,N_2784,N_2815);
nand U2874 (N_2874,N_2805,N_2797);
nand U2875 (N_2875,N_2776,N_2809);
nor U2876 (N_2876,N_2800,N_2783);
or U2877 (N_2877,N_2780,N_2768);
nor U2878 (N_2878,N_2785,N_2770);
xor U2879 (N_2879,N_2761,N_2779);
nand U2880 (N_2880,N_2853,N_2864);
and U2881 (N_2881,N_2860,N_2827);
nor U2882 (N_2882,N_2839,N_2873);
nand U2883 (N_2883,N_2867,N_2856);
and U2884 (N_2884,N_2859,N_2837);
and U2885 (N_2885,N_2830,N_2842);
xor U2886 (N_2886,N_2863,N_2878);
nor U2887 (N_2887,N_2861,N_2870);
and U2888 (N_2888,N_2840,N_2828);
or U2889 (N_2889,N_2824,N_2854);
or U2890 (N_2890,N_2826,N_2844);
xor U2891 (N_2891,N_2868,N_2848);
and U2892 (N_2892,N_2841,N_2850);
or U2893 (N_2893,N_2862,N_2834);
nor U2894 (N_2894,N_2869,N_2829);
nand U2895 (N_2895,N_2876,N_2852);
and U2896 (N_2896,N_2872,N_2821);
and U2897 (N_2897,N_2831,N_2875);
xnor U2898 (N_2898,N_2836,N_2846);
nor U2899 (N_2899,N_2845,N_2833);
or U2900 (N_2900,N_2866,N_2823);
and U2901 (N_2901,N_2849,N_2822);
and U2902 (N_2902,N_2838,N_2855);
xor U2903 (N_2903,N_2851,N_2877);
xnor U2904 (N_2904,N_2832,N_2825);
nor U2905 (N_2905,N_2871,N_2857);
and U2906 (N_2906,N_2835,N_2879);
and U2907 (N_2907,N_2858,N_2865);
nor U2908 (N_2908,N_2847,N_2874);
xor U2909 (N_2909,N_2843,N_2820);
or U2910 (N_2910,N_2878,N_2867);
nor U2911 (N_2911,N_2851,N_2822);
xnor U2912 (N_2912,N_2859,N_2870);
xnor U2913 (N_2913,N_2851,N_2821);
xor U2914 (N_2914,N_2872,N_2860);
or U2915 (N_2915,N_2879,N_2834);
xnor U2916 (N_2916,N_2854,N_2852);
and U2917 (N_2917,N_2865,N_2837);
nor U2918 (N_2918,N_2827,N_2856);
xor U2919 (N_2919,N_2873,N_2833);
and U2920 (N_2920,N_2820,N_2845);
or U2921 (N_2921,N_2845,N_2838);
xnor U2922 (N_2922,N_2840,N_2864);
xnor U2923 (N_2923,N_2870,N_2835);
and U2924 (N_2924,N_2823,N_2867);
and U2925 (N_2925,N_2854,N_2834);
nand U2926 (N_2926,N_2868,N_2852);
and U2927 (N_2927,N_2840,N_2835);
and U2928 (N_2928,N_2820,N_2856);
nand U2929 (N_2929,N_2856,N_2824);
xnor U2930 (N_2930,N_2879,N_2855);
nor U2931 (N_2931,N_2879,N_2836);
xnor U2932 (N_2932,N_2865,N_2868);
xnor U2933 (N_2933,N_2836,N_2839);
or U2934 (N_2934,N_2847,N_2821);
or U2935 (N_2935,N_2847,N_2868);
and U2936 (N_2936,N_2823,N_2879);
or U2937 (N_2937,N_2822,N_2844);
and U2938 (N_2938,N_2865,N_2842);
nor U2939 (N_2939,N_2825,N_2849);
and U2940 (N_2940,N_2895,N_2902);
nand U2941 (N_2941,N_2886,N_2914);
nor U2942 (N_2942,N_2898,N_2912);
nand U2943 (N_2943,N_2913,N_2891);
nand U2944 (N_2944,N_2910,N_2893);
nand U2945 (N_2945,N_2882,N_2924);
and U2946 (N_2946,N_2896,N_2925);
xor U2947 (N_2947,N_2915,N_2908);
xnor U2948 (N_2948,N_2919,N_2918);
nand U2949 (N_2949,N_2926,N_2937);
or U2950 (N_2950,N_2887,N_2881);
xor U2951 (N_2951,N_2880,N_2911);
xor U2952 (N_2952,N_2905,N_2923);
and U2953 (N_2953,N_2888,N_2936);
nor U2954 (N_2954,N_2897,N_2935);
nand U2955 (N_2955,N_2916,N_2907);
nand U2956 (N_2956,N_2903,N_2885);
nand U2957 (N_2957,N_2931,N_2922);
and U2958 (N_2958,N_2939,N_2906);
nand U2959 (N_2959,N_2889,N_2938);
or U2960 (N_2960,N_2930,N_2892);
nor U2961 (N_2961,N_2900,N_2932);
xnor U2962 (N_2962,N_2909,N_2928);
or U2963 (N_2963,N_2933,N_2934);
nand U2964 (N_2964,N_2929,N_2927);
nor U2965 (N_2965,N_2920,N_2890);
nor U2966 (N_2966,N_2883,N_2904);
xnor U2967 (N_2967,N_2894,N_2921);
xnor U2968 (N_2968,N_2901,N_2899);
and U2969 (N_2969,N_2917,N_2884);
and U2970 (N_2970,N_2902,N_2939);
nand U2971 (N_2971,N_2903,N_2928);
and U2972 (N_2972,N_2883,N_2903);
and U2973 (N_2973,N_2902,N_2917);
or U2974 (N_2974,N_2924,N_2928);
or U2975 (N_2975,N_2932,N_2914);
nand U2976 (N_2976,N_2934,N_2919);
nor U2977 (N_2977,N_2882,N_2923);
nand U2978 (N_2978,N_2921,N_2888);
nor U2979 (N_2979,N_2893,N_2896);
or U2980 (N_2980,N_2936,N_2921);
nand U2981 (N_2981,N_2923,N_2897);
nand U2982 (N_2982,N_2921,N_2905);
nor U2983 (N_2983,N_2917,N_2906);
nand U2984 (N_2984,N_2937,N_2906);
and U2985 (N_2985,N_2895,N_2931);
xor U2986 (N_2986,N_2924,N_2930);
nor U2987 (N_2987,N_2926,N_2934);
nand U2988 (N_2988,N_2920,N_2885);
nor U2989 (N_2989,N_2891,N_2906);
or U2990 (N_2990,N_2906,N_2885);
nor U2991 (N_2991,N_2901,N_2885);
and U2992 (N_2992,N_2932,N_2909);
or U2993 (N_2993,N_2938,N_2904);
nor U2994 (N_2994,N_2919,N_2928);
and U2995 (N_2995,N_2891,N_2927);
or U2996 (N_2996,N_2928,N_2889);
or U2997 (N_2997,N_2893,N_2935);
and U2998 (N_2998,N_2899,N_2926);
and U2999 (N_2999,N_2887,N_2892);
nand UO_0 (O_0,N_2954,N_2984);
nor UO_1 (O_1,N_2948,N_2958);
or UO_2 (O_2,N_2988,N_2949);
xor UO_3 (O_3,N_2998,N_2980);
or UO_4 (O_4,N_2943,N_2950);
xnor UO_5 (O_5,N_2978,N_2963);
xor UO_6 (O_6,N_2955,N_2983);
or UO_7 (O_7,N_2969,N_2942);
xnor UO_8 (O_8,N_2953,N_2973);
or UO_9 (O_9,N_2986,N_2981);
nor UO_10 (O_10,N_2965,N_2974);
and UO_11 (O_11,N_2992,N_2995);
and UO_12 (O_12,N_2956,N_2993);
nor UO_13 (O_13,N_2985,N_2945);
nor UO_14 (O_14,N_2996,N_2941);
nand UO_15 (O_15,N_2999,N_2989);
nand UO_16 (O_16,N_2975,N_2987);
or UO_17 (O_17,N_2944,N_2964);
nor UO_18 (O_18,N_2994,N_2972);
or UO_19 (O_19,N_2947,N_2970);
and UO_20 (O_20,N_2962,N_2946);
nand UO_21 (O_21,N_2982,N_2940);
nor UO_22 (O_22,N_2997,N_2951);
nor UO_23 (O_23,N_2959,N_2990);
and UO_24 (O_24,N_2968,N_2961);
nor UO_25 (O_25,N_2952,N_2991);
nand UO_26 (O_26,N_2976,N_2971);
xor UO_27 (O_27,N_2960,N_2977);
or UO_28 (O_28,N_2979,N_2967);
xor UO_29 (O_29,N_2966,N_2957);
nor UO_30 (O_30,N_2956,N_2969);
nor UO_31 (O_31,N_2983,N_2999);
nor UO_32 (O_32,N_2989,N_2997);
xnor UO_33 (O_33,N_2983,N_2952);
and UO_34 (O_34,N_2992,N_2953);
and UO_35 (O_35,N_2972,N_2983);
xnor UO_36 (O_36,N_2948,N_2984);
and UO_37 (O_37,N_2960,N_2996);
or UO_38 (O_38,N_2956,N_2957);
and UO_39 (O_39,N_2968,N_2981);
nand UO_40 (O_40,N_2978,N_2973);
nand UO_41 (O_41,N_2945,N_2997);
nor UO_42 (O_42,N_2964,N_2995);
nor UO_43 (O_43,N_2994,N_2969);
and UO_44 (O_44,N_2957,N_2958);
and UO_45 (O_45,N_2998,N_2974);
and UO_46 (O_46,N_2991,N_2994);
nand UO_47 (O_47,N_2978,N_2994);
nor UO_48 (O_48,N_2979,N_2985);
and UO_49 (O_49,N_2943,N_2940);
xnor UO_50 (O_50,N_2955,N_2979);
xor UO_51 (O_51,N_2949,N_2995);
or UO_52 (O_52,N_2956,N_2986);
xnor UO_53 (O_53,N_2948,N_2974);
nand UO_54 (O_54,N_2994,N_2985);
nor UO_55 (O_55,N_2989,N_2972);
and UO_56 (O_56,N_2955,N_2946);
nand UO_57 (O_57,N_2966,N_2988);
and UO_58 (O_58,N_2987,N_2993);
and UO_59 (O_59,N_2980,N_2995);
or UO_60 (O_60,N_2964,N_2972);
nand UO_61 (O_61,N_2991,N_2953);
xnor UO_62 (O_62,N_2962,N_2967);
xnor UO_63 (O_63,N_2989,N_2973);
or UO_64 (O_64,N_2981,N_2984);
or UO_65 (O_65,N_2954,N_2995);
or UO_66 (O_66,N_2962,N_2942);
or UO_67 (O_67,N_2990,N_2993);
and UO_68 (O_68,N_2995,N_2948);
nand UO_69 (O_69,N_2947,N_2944);
or UO_70 (O_70,N_2951,N_2989);
nor UO_71 (O_71,N_2978,N_2954);
xnor UO_72 (O_72,N_2969,N_2999);
and UO_73 (O_73,N_2961,N_2977);
nor UO_74 (O_74,N_2988,N_2986);
and UO_75 (O_75,N_2944,N_2997);
or UO_76 (O_76,N_2991,N_2990);
xnor UO_77 (O_77,N_2951,N_2949);
nand UO_78 (O_78,N_2977,N_2965);
or UO_79 (O_79,N_2967,N_2995);
xnor UO_80 (O_80,N_2947,N_2950);
and UO_81 (O_81,N_2998,N_2943);
and UO_82 (O_82,N_2947,N_2981);
or UO_83 (O_83,N_2988,N_2980);
xnor UO_84 (O_84,N_2977,N_2987);
or UO_85 (O_85,N_2948,N_2973);
or UO_86 (O_86,N_2991,N_2985);
or UO_87 (O_87,N_2951,N_2978);
nand UO_88 (O_88,N_2978,N_2967);
nand UO_89 (O_89,N_2950,N_2976);
and UO_90 (O_90,N_2999,N_2957);
nor UO_91 (O_91,N_2969,N_2958);
xor UO_92 (O_92,N_2970,N_2979);
nor UO_93 (O_93,N_2944,N_2963);
nor UO_94 (O_94,N_2995,N_2941);
xnor UO_95 (O_95,N_2955,N_2970);
and UO_96 (O_96,N_2985,N_2949);
nor UO_97 (O_97,N_2967,N_2961);
xor UO_98 (O_98,N_2940,N_2978);
and UO_99 (O_99,N_2979,N_2994);
xnor UO_100 (O_100,N_2948,N_2949);
xor UO_101 (O_101,N_2940,N_2997);
xnor UO_102 (O_102,N_2980,N_2957);
nor UO_103 (O_103,N_2961,N_2976);
and UO_104 (O_104,N_2973,N_2960);
nor UO_105 (O_105,N_2964,N_2975);
nand UO_106 (O_106,N_2960,N_2991);
nand UO_107 (O_107,N_2993,N_2997);
xor UO_108 (O_108,N_2950,N_2992);
nand UO_109 (O_109,N_2979,N_2957);
xor UO_110 (O_110,N_2956,N_2981);
or UO_111 (O_111,N_2987,N_2942);
or UO_112 (O_112,N_2986,N_2963);
nand UO_113 (O_113,N_2941,N_2954);
nand UO_114 (O_114,N_2974,N_2982);
or UO_115 (O_115,N_2996,N_2976);
and UO_116 (O_116,N_2984,N_2994);
or UO_117 (O_117,N_2974,N_2985);
nor UO_118 (O_118,N_2943,N_2973);
xnor UO_119 (O_119,N_2970,N_2941);
nand UO_120 (O_120,N_2967,N_2945);
and UO_121 (O_121,N_2997,N_2996);
or UO_122 (O_122,N_2961,N_2955);
nand UO_123 (O_123,N_2945,N_2970);
nand UO_124 (O_124,N_2957,N_2992);
or UO_125 (O_125,N_2966,N_2983);
nor UO_126 (O_126,N_2960,N_2992);
or UO_127 (O_127,N_2997,N_2954);
xnor UO_128 (O_128,N_2956,N_2992);
xnor UO_129 (O_129,N_2953,N_2975);
or UO_130 (O_130,N_2955,N_2999);
xor UO_131 (O_131,N_2995,N_2959);
nor UO_132 (O_132,N_2982,N_2994);
nand UO_133 (O_133,N_2997,N_2973);
nand UO_134 (O_134,N_2944,N_2993);
xnor UO_135 (O_135,N_2951,N_2963);
or UO_136 (O_136,N_2960,N_2943);
and UO_137 (O_137,N_2961,N_2966);
or UO_138 (O_138,N_2942,N_2958);
or UO_139 (O_139,N_2955,N_2969);
and UO_140 (O_140,N_2990,N_2953);
and UO_141 (O_141,N_2964,N_2974);
nand UO_142 (O_142,N_2998,N_2958);
nor UO_143 (O_143,N_2953,N_2997);
nand UO_144 (O_144,N_2980,N_2943);
nor UO_145 (O_145,N_2944,N_2971);
xor UO_146 (O_146,N_2966,N_2996);
or UO_147 (O_147,N_2989,N_2958);
nor UO_148 (O_148,N_2951,N_2975);
xor UO_149 (O_149,N_2940,N_2966);
nor UO_150 (O_150,N_2945,N_2980);
xor UO_151 (O_151,N_2947,N_2997);
or UO_152 (O_152,N_2998,N_2992);
nand UO_153 (O_153,N_2981,N_2944);
nand UO_154 (O_154,N_2964,N_2994);
or UO_155 (O_155,N_2948,N_2963);
nand UO_156 (O_156,N_2981,N_2998);
nand UO_157 (O_157,N_2944,N_2956);
nor UO_158 (O_158,N_2974,N_2943);
and UO_159 (O_159,N_2994,N_2971);
or UO_160 (O_160,N_2951,N_2962);
nand UO_161 (O_161,N_2974,N_2949);
nand UO_162 (O_162,N_2990,N_2955);
xnor UO_163 (O_163,N_2995,N_2987);
xor UO_164 (O_164,N_2973,N_2967);
nand UO_165 (O_165,N_2961,N_2972);
or UO_166 (O_166,N_2974,N_2991);
nor UO_167 (O_167,N_2947,N_2976);
xnor UO_168 (O_168,N_2980,N_2955);
xor UO_169 (O_169,N_2993,N_2943);
or UO_170 (O_170,N_2955,N_2943);
or UO_171 (O_171,N_2982,N_2990);
and UO_172 (O_172,N_2997,N_2970);
xnor UO_173 (O_173,N_2995,N_2975);
or UO_174 (O_174,N_2968,N_2959);
or UO_175 (O_175,N_2994,N_2956);
and UO_176 (O_176,N_2996,N_2956);
nand UO_177 (O_177,N_2986,N_2970);
and UO_178 (O_178,N_2963,N_2997);
xor UO_179 (O_179,N_2972,N_2976);
and UO_180 (O_180,N_2974,N_2961);
nor UO_181 (O_181,N_2975,N_2989);
nand UO_182 (O_182,N_2942,N_2957);
and UO_183 (O_183,N_2998,N_2991);
nand UO_184 (O_184,N_2988,N_2971);
or UO_185 (O_185,N_2989,N_2980);
and UO_186 (O_186,N_2980,N_2950);
nor UO_187 (O_187,N_2940,N_2944);
nand UO_188 (O_188,N_2951,N_2943);
nand UO_189 (O_189,N_2977,N_2951);
and UO_190 (O_190,N_2977,N_2976);
xnor UO_191 (O_191,N_2984,N_2993);
and UO_192 (O_192,N_2966,N_2986);
or UO_193 (O_193,N_2982,N_2961);
xor UO_194 (O_194,N_2987,N_2978);
nor UO_195 (O_195,N_2942,N_2960);
xor UO_196 (O_196,N_2943,N_2981);
nand UO_197 (O_197,N_2966,N_2971);
and UO_198 (O_198,N_2969,N_2944);
or UO_199 (O_199,N_2989,N_2955);
and UO_200 (O_200,N_2999,N_2968);
and UO_201 (O_201,N_2984,N_2956);
nand UO_202 (O_202,N_2947,N_2969);
and UO_203 (O_203,N_2972,N_2948);
nor UO_204 (O_204,N_2954,N_2961);
and UO_205 (O_205,N_2940,N_2951);
nor UO_206 (O_206,N_2944,N_2960);
or UO_207 (O_207,N_2965,N_2958);
and UO_208 (O_208,N_2992,N_2952);
xnor UO_209 (O_209,N_2969,N_2948);
xnor UO_210 (O_210,N_2974,N_2950);
nor UO_211 (O_211,N_2972,N_2992);
or UO_212 (O_212,N_2950,N_2962);
or UO_213 (O_213,N_2983,N_2967);
and UO_214 (O_214,N_2975,N_2970);
xnor UO_215 (O_215,N_2972,N_2975);
xor UO_216 (O_216,N_2973,N_2966);
nor UO_217 (O_217,N_2976,N_2979);
and UO_218 (O_218,N_2981,N_2995);
or UO_219 (O_219,N_2999,N_2965);
or UO_220 (O_220,N_2954,N_2974);
xnor UO_221 (O_221,N_2986,N_2984);
xnor UO_222 (O_222,N_2985,N_2980);
nor UO_223 (O_223,N_2984,N_2988);
and UO_224 (O_224,N_2997,N_2986);
xor UO_225 (O_225,N_2967,N_2974);
nor UO_226 (O_226,N_2976,N_2967);
xor UO_227 (O_227,N_2944,N_2945);
or UO_228 (O_228,N_2971,N_2973);
and UO_229 (O_229,N_2949,N_2964);
xnor UO_230 (O_230,N_2980,N_2959);
or UO_231 (O_231,N_2976,N_2957);
nand UO_232 (O_232,N_2962,N_2966);
or UO_233 (O_233,N_2945,N_2969);
nor UO_234 (O_234,N_2969,N_2957);
or UO_235 (O_235,N_2963,N_2981);
and UO_236 (O_236,N_2961,N_2971);
and UO_237 (O_237,N_2985,N_2964);
nand UO_238 (O_238,N_2947,N_2978);
xnor UO_239 (O_239,N_2949,N_2960);
nor UO_240 (O_240,N_2995,N_2985);
nand UO_241 (O_241,N_2962,N_2943);
and UO_242 (O_242,N_2992,N_2993);
nand UO_243 (O_243,N_2999,N_2991);
nand UO_244 (O_244,N_2979,N_2962);
nand UO_245 (O_245,N_2973,N_2968);
xor UO_246 (O_246,N_2957,N_2963);
nand UO_247 (O_247,N_2940,N_2964);
xnor UO_248 (O_248,N_2968,N_2948);
nor UO_249 (O_249,N_2954,N_2967);
nor UO_250 (O_250,N_2960,N_2972);
nor UO_251 (O_251,N_2942,N_2970);
and UO_252 (O_252,N_2946,N_2957);
or UO_253 (O_253,N_2963,N_2964);
and UO_254 (O_254,N_2965,N_2981);
or UO_255 (O_255,N_2990,N_2981);
or UO_256 (O_256,N_2999,N_2960);
or UO_257 (O_257,N_2944,N_2984);
xnor UO_258 (O_258,N_2964,N_2942);
nand UO_259 (O_259,N_2988,N_2969);
xnor UO_260 (O_260,N_2959,N_2963);
or UO_261 (O_261,N_2975,N_2957);
nand UO_262 (O_262,N_2944,N_2982);
xnor UO_263 (O_263,N_2989,N_2957);
nand UO_264 (O_264,N_2990,N_2986);
and UO_265 (O_265,N_2955,N_2996);
xnor UO_266 (O_266,N_2944,N_2999);
or UO_267 (O_267,N_2990,N_2985);
xor UO_268 (O_268,N_2947,N_2989);
nand UO_269 (O_269,N_2967,N_2964);
or UO_270 (O_270,N_2942,N_2980);
nor UO_271 (O_271,N_2992,N_2963);
nor UO_272 (O_272,N_2993,N_2982);
xor UO_273 (O_273,N_2961,N_2950);
xnor UO_274 (O_274,N_2967,N_2947);
nor UO_275 (O_275,N_2996,N_2994);
and UO_276 (O_276,N_2971,N_2967);
and UO_277 (O_277,N_2952,N_2980);
or UO_278 (O_278,N_2991,N_2973);
or UO_279 (O_279,N_2993,N_2965);
nand UO_280 (O_280,N_2981,N_2969);
nor UO_281 (O_281,N_2965,N_2970);
nand UO_282 (O_282,N_2981,N_2992);
and UO_283 (O_283,N_2995,N_2982);
xor UO_284 (O_284,N_2971,N_2965);
and UO_285 (O_285,N_2968,N_2950);
and UO_286 (O_286,N_2981,N_2993);
nor UO_287 (O_287,N_2960,N_2978);
xnor UO_288 (O_288,N_2999,N_2954);
nand UO_289 (O_289,N_2960,N_2990);
xor UO_290 (O_290,N_2949,N_2950);
nand UO_291 (O_291,N_2949,N_2980);
xnor UO_292 (O_292,N_2960,N_2959);
nand UO_293 (O_293,N_2973,N_2982);
and UO_294 (O_294,N_2981,N_2975);
xnor UO_295 (O_295,N_2995,N_2976);
and UO_296 (O_296,N_2996,N_2982);
xor UO_297 (O_297,N_2950,N_2953);
nand UO_298 (O_298,N_2967,N_2948);
xor UO_299 (O_299,N_2956,N_2975);
nand UO_300 (O_300,N_2982,N_2958);
nor UO_301 (O_301,N_2964,N_2957);
xnor UO_302 (O_302,N_2973,N_2992);
xnor UO_303 (O_303,N_2962,N_2948);
nand UO_304 (O_304,N_2999,N_2980);
nand UO_305 (O_305,N_2993,N_2955);
or UO_306 (O_306,N_2971,N_2964);
nand UO_307 (O_307,N_2974,N_2980);
nand UO_308 (O_308,N_2968,N_2975);
nor UO_309 (O_309,N_2966,N_2981);
xor UO_310 (O_310,N_2984,N_2950);
nor UO_311 (O_311,N_2953,N_2977);
nor UO_312 (O_312,N_2949,N_2978);
xnor UO_313 (O_313,N_2988,N_2962);
and UO_314 (O_314,N_2949,N_2957);
or UO_315 (O_315,N_2941,N_2952);
nand UO_316 (O_316,N_2942,N_2977);
nand UO_317 (O_317,N_2985,N_2975);
nor UO_318 (O_318,N_2976,N_2958);
xnor UO_319 (O_319,N_2968,N_2952);
and UO_320 (O_320,N_2984,N_2989);
or UO_321 (O_321,N_2978,N_2995);
xnor UO_322 (O_322,N_2981,N_2953);
and UO_323 (O_323,N_2989,N_2967);
and UO_324 (O_324,N_2970,N_2961);
and UO_325 (O_325,N_2965,N_2942);
and UO_326 (O_326,N_2947,N_2958);
nand UO_327 (O_327,N_2962,N_2978);
xor UO_328 (O_328,N_2946,N_2945);
nand UO_329 (O_329,N_2975,N_2954);
xnor UO_330 (O_330,N_2963,N_2958);
and UO_331 (O_331,N_2950,N_2993);
xor UO_332 (O_332,N_2957,N_2997);
and UO_333 (O_333,N_2980,N_2967);
and UO_334 (O_334,N_2976,N_2981);
and UO_335 (O_335,N_2957,N_2993);
and UO_336 (O_336,N_2973,N_2984);
nor UO_337 (O_337,N_2972,N_2969);
nand UO_338 (O_338,N_2982,N_2954);
nor UO_339 (O_339,N_2975,N_2962);
nand UO_340 (O_340,N_2962,N_2981);
and UO_341 (O_341,N_2951,N_2945);
nand UO_342 (O_342,N_2963,N_2977);
nand UO_343 (O_343,N_2957,N_2972);
nor UO_344 (O_344,N_2999,N_2946);
and UO_345 (O_345,N_2945,N_2961);
or UO_346 (O_346,N_2999,N_2974);
and UO_347 (O_347,N_2958,N_2951);
xor UO_348 (O_348,N_2946,N_2974);
and UO_349 (O_349,N_2984,N_2947);
nor UO_350 (O_350,N_2972,N_2980);
nand UO_351 (O_351,N_2950,N_2982);
or UO_352 (O_352,N_2988,N_2982);
or UO_353 (O_353,N_2940,N_2948);
xnor UO_354 (O_354,N_2959,N_2983);
nor UO_355 (O_355,N_2997,N_2991);
or UO_356 (O_356,N_2943,N_2952);
xor UO_357 (O_357,N_2963,N_2941);
or UO_358 (O_358,N_2942,N_2953);
nor UO_359 (O_359,N_2988,N_2942);
and UO_360 (O_360,N_2990,N_2974);
or UO_361 (O_361,N_2947,N_2963);
nor UO_362 (O_362,N_2954,N_2994);
and UO_363 (O_363,N_2986,N_2998);
nand UO_364 (O_364,N_2942,N_2990);
nand UO_365 (O_365,N_2951,N_2979);
or UO_366 (O_366,N_2982,N_2963);
and UO_367 (O_367,N_2997,N_2981);
xnor UO_368 (O_368,N_2970,N_2964);
and UO_369 (O_369,N_2945,N_2975);
nor UO_370 (O_370,N_2964,N_2945);
nand UO_371 (O_371,N_2963,N_2983);
xnor UO_372 (O_372,N_2998,N_2940);
nor UO_373 (O_373,N_2977,N_2971);
xnor UO_374 (O_374,N_2986,N_2964);
nor UO_375 (O_375,N_2980,N_2944);
nand UO_376 (O_376,N_2973,N_2974);
or UO_377 (O_377,N_2988,N_2953);
nor UO_378 (O_378,N_2955,N_2973);
xor UO_379 (O_379,N_2992,N_2979);
nor UO_380 (O_380,N_2951,N_2972);
nor UO_381 (O_381,N_2958,N_2996);
nor UO_382 (O_382,N_2969,N_2962);
and UO_383 (O_383,N_2978,N_2970);
xnor UO_384 (O_384,N_2940,N_2977);
xnor UO_385 (O_385,N_2992,N_2989);
nand UO_386 (O_386,N_2974,N_2970);
xor UO_387 (O_387,N_2983,N_2992);
nand UO_388 (O_388,N_2970,N_2976);
and UO_389 (O_389,N_2963,N_2994);
nor UO_390 (O_390,N_2977,N_2962);
nor UO_391 (O_391,N_2968,N_2989);
and UO_392 (O_392,N_2962,N_2983);
and UO_393 (O_393,N_2990,N_2980);
or UO_394 (O_394,N_2985,N_2978);
and UO_395 (O_395,N_2950,N_2946);
nor UO_396 (O_396,N_2994,N_2989);
and UO_397 (O_397,N_2967,N_2984);
nor UO_398 (O_398,N_2971,N_2960);
xnor UO_399 (O_399,N_2984,N_2966);
nor UO_400 (O_400,N_2969,N_2979);
xnor UO_401 (O_401,N_2956,N_2962);
xor UO_402 (O_402,N_2940,N_2945);
nor UO_403 (O_403,N_2970,N_2949);
and UO_404 (O_404,N_2957,N_2971);
nor UO_405 (O_405,N_2972,N_2966);
or UO_406 (O_406,N_2970,N_2995);
nand UO_407 (O_407,N_2959,N_2993);
or UO_408 (O_408,N_2970,N_2962);
xnor UO_409 (O_409,N_2978,N_2966);
or UO_410 (O_410,N_2989,N_2959);
xor UO_411 (O_411,N_2954,N_2947);
nor UO_412 (O_412,N_2979,N_2940);
and UO_413 (O_413,N_2997,N_2968);
nand UO_414 (O_414,N_2991,N_2945);
or UO_415 (O_415,N_2988,N_2991);
and UO_416 (O_416,N_2984,N_2975);
nor UO_417 (O_417,N_2956,N_2985);
nor UO_418 (O_418,N_2967,N_2943);
xor UO_419 (O_419,N_2999,N_2943);
nor UO_420 (O_420,N_2958,N_2960);
or UO_421 (O_421,N_2999,N_2966);
nand UO_422 (O_422,N_2977,N_2956);
or UO_423 (O_423,N_2969,N_2966);
nor UO_424 (O_424,N_2953,N_2955);
and UO_425 (O_425,N_2970,N_2989);
nand UO_426 (O_426,N_2976,N_2959);
nand UO_427 (O_427,N_2940,N_2956);
and UO_428 (O_428,N_2998,N_2968);
nand UO_429 (O_429,N_2999,N_2976);
or UO_430 (O_430,N_2956,N_2941);
or UO_431 (O_431,N_2969,N_2959);
xnor UO_432 (O_432,N_2999,N_2940);
nor UO_433 (O_433,N_2947,N_2961);
or UO_434 (O_434,N_2940,N_2955);
nand UO_435 (O_435,N_2963,N_2962);
nand UO_436 (O_436,N_2952,N_2994);
nand UO_437 (O_437,N_2982,N_2969);
or UO_438 (O_438,N_2968,N_2956);
and UO_439 (O_439,N_2998,N_2954);
nand UO_440 (O_440,N_2982,N_2975);
and UO_441 (O_441,N_2959,N_2987);
or UO_442 (O_442,N_2970,N_2993);
or UO_443 (O_443,N_2990,N_2966);
or UO_444 (O_444,N_2964,N_2999);
or UO_445 (O_445,N_2969,N_2943);
and UO_446 (O_446,N_2981,N_2954);
and UO_447 (O_447,N_2960,N_2997);
nor UO_448 (O_448,N_2990,N_2950);
or UO_449 (O_449,N_2988,N_2961);
and UO_450 (O_450,N_2970,N_2987);
xnor UO_451 (O_451,N_2951,N_2967);
and UO_452 (O_452,N_2961,N_2941);
and UO_453 (O_453,N_2959,N_2945);
nand UO_454 (O_454,N_2955,N_2967);
or UO_455 (O_455,N_2941,N_2965);
nor UO_456 (O_456,N_2989,N_2981);
nand UO_457 (O_457,N_2992,N_2943);
nor UO_458 (O_458,N_2967,N_2959);
nor UO_459 (O_459,N_2982,N_2997);
nand UO_460 (O_460,N_2964,N_2979);
and UO_461 (O_461,N_2963,N_2953);
or UO_462 (O_462,N_2940,N_2958);
and UO_463 (O_463,N_2972,N_2962);
nand UO_464 (O_464,N_2986,N_2957);
and UO_465 (O_465,N_2940,N_2990);
or UO_466 (O_466,N_2961,N_2958);
nor UO_467 (O_467,N_2962,N_2990);
xor UO_468 (O_468,N_2956,N_2963);
or UO_469 (O_469,N_2966,N_2991);
nand UO_470 (O_470,N_2952,N_2976);
or UO_471 (O_471,N_2958,N_2988);
or UO_472 (O_472,N_2953,N_2969);
nand UO_473 (O_473,N_2977,N_2952);
and UO_474 (O_474,N_2952,N_2962);
or UO_475 (O_475,N_2963,N_2949);
xor UO_476 (O_476,N_2949,N_2982);
xnor UO_477 (O_477,N_2998,N_2951);
nand UO_478 (O_478,N_2951,N_2982);
nor UO_479 (O_479,N_2960,N_2945);
or UO_480 (O_480,N_2941,N_2981);
nand UO_481 (O_481,N_2974,N_2994);
nand UO_482 (O_482,N_2942,N_2974);
xor UO_483 (O_483,N_2996,N_2963);
nor UO_484 (O_484,N_2991,N_2941);
or UO_485 (O_485,N_2989,N_2953);
nand UO_486 (O_486,N_2961,N_2948);
nor UO_487 (O_487,N_2969,N_2954);
nor UO_488 (O_488,N_2949,N_2946);
xnor UO_489 (O_489,N_2961,N_2996);
or UO_490 (O_490,N_2946,N_2968);
xnor UO_491 (O_491,N_2968,N_2980);
nor UO_492 (O_492,N_2986,N_2950);
nand UO_493 (O_493,N_2959,N_2946);
xor UO_494 (O_494,N_2980,N_2940);
xor UO_495 (O_495,N_2992,N_2948);
nand UO_496 (O_496,N_2996,N_2978);
and UO_497 (O_497,N_2964,N_2950);
xnor UO_498 (O_498,N_2973,N_2987);
or UO_499 (O_499,N_2962,N_2960);
endmodule